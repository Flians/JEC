// Benchmark "c7552" written by ABC on Wed May 27 22:07:51 2020

module rf_c7552 ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496,
    G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253,
    G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743,
    G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432,
    G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire n317, n318, n319, n320, n321, n322, n324, n325, n326, n327, n328,
    n329, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342,
    n343, n345, n347, n348, n349, n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1127,
    n1128, n1129, n1130, n1131, n1132, n1134, n1136, n1137, n1139, n1140,
    n1142, n1143, n1144, n1146, n1148, n1149, n1150, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1387, n1388, n1389,
    n1390, n1391, n1392, n1394, n1395, n1396, n1397, n1398, n1399, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1410, n1412, n1413,
    n1414, n1415, n1417, n1418, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1429, n1430, n1432, n1433, n1435, n1436, n1438, n1439,
    n1440, n1441, n1442, n1444, n1445, n1446, n1447, n1448, n1449, n1451,
    n1453, n1454, n1455, n1456, n1460, n1461, n1462, n1463, n1464, n1465,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1477, n1479,
    n1480, n1482, n1483, n1484, n1486, n1487, n1488, n1490, n1492, n1493,
    n1494, n1495, n1496, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
  jnot g0000(.din(G15), .dout(G279));
  jor  g0001(.dina(G57), .dinb(G5), .dout(G402));
  jnot g0002(.din(G184), .dout(n317));
  jnot g0003(.din(G228), .dout(n318));
  jor  g0004(.dina(n318), .dinb(n317), .dout(n319));
  jnot g0005(.din(G150), .dout(n320));
  jnot g0006(.din(G240), .dout(n321));
  jor  g0007(.dina(n321), .dinb(n320), .dout(n322));
  jor  g0008(.dina(n322), .dinb(n319), .dout(G404));
  jnot g0009(.din(G210), .dout(n324));
  jnot g0010(.din(G218), .dout(n325));
  jor  g0011(.dina(n325), .dinb(n324), .dout(n326));
  jnot g0012(.din(G152), .dout(n327));
  jnot g0013(.din(G230), .dout(n328));
  jor  g0014(.dina(n328), .dinb(n327), .dout(n329));
  jor  g0015(.dina(n329), .dinb(n326), .dout(G406));
  jnot g0016(.din(G183), .dout(n331));
  jnot g0017(.din(G185), .dout(n332));
  jor  g0018(.dina(n332), .dinb(n331), .dout(n333));
  jnot g0019(.din(G182), .dout(n334));
  jnot g0020(.din(G186), .dout(n335));
  jor  g0021(.dina(n335), .dinb(n334), .dout(n336));
  jor  g0022(.dina(n336), .dinb(n333), .dout(G408));
  jnot g0023(.din(G172), .dout(n338));
  jnot g0024(.din(G188), .dout(n339));
  jor  g0025(.dina(n339), .dinb(n338), .dout(n340));
  jnot g0026(.din(G162), .dout(n341));
  jnot g0027(.din(G199), .dout(n342));
  jor  g0028(.dina(n342), .dinb(n341), .dout(n343));
  jor  g0029(.dina(n343), .dinb(n340), .dout(G410));
  jnot g0030(.din(G1197), .dout(n345));
  jor  g0031(.dina(n345), .dinb(G5), .dout(G284));
  jnot g0032(.din(G133), .dout(n347));
  jnot g0033(.din(G134), .dout(n348));
  jor  g0034(.dina(n348), .dinb(n347), .dout(n349));
  jor  g0035(.dina(n349), .dinb(G5), .dout(G292));
  jand g0036(.dina(G163), .dinb(G1), .dout(G278));
  jnot g0037(.din(G41), .dout(n352));
  jor  g0038(.dina(n352), .dinb(G18), .dout(n353));
  jor  g0039(.dina(n353), .dinb(G3701), .dout(n354));
  jnot g0040(.din(G18), .dout(n355));
  jand g0041(.dina(G41), .dinb(n355), .dout(n356));
  jand g0042(.dina(G229), .dinb(G18), .dout(n357));
  jor  g0043(.dina(n357), .dinb(n356), .dout(n358));
  jand g0044(.dina(G3701), .dinb(n355), .dout(n359));
  jnot g0045(.din(n359), .dout(n360));
  jor  g0046(.dina(n360), .dinb(n358), .dout(n361));
  jand g0047(.dina(n361), .dinb(n354), .dout(n362));
  jxor g0048(.dina(n362), .dinb(G4526), .dout(G373));
  jand g0049(.dina(G4528), .dinb(G1496), .dout(n364));
  jxor g0050(.dina(n364), .dinb(G38), .dout(n365));
  jnot g0051(.din(G3723), .dout(n366));
  jand g0052(.dina(G235), .dinb(G18), .dout(n367));
  jnot g0053(.din(n367), .dout(n368));
  jnot g0054(.din(G103), .dout(n369));
  jor  g0055(.dina(n369), .dinb(G18), .dout(n370));
  jand g0056(.dina(n370), .dinb(n368), .dout(n371));
  jxor g0057(.dina(n371), .dinb(n366), .dout(n372));
  jand g0058(.dina(G236), .dinb(G18), .dout(n373));
  jnot g0059(.din(n373), .dout(n374));
  jnot g0060(.din(G23), .dout(n375));
  jor  g0061(.dina(n375), .dinb(G18), .dout(n376));
  jand g0062(.dina(n376), .dinb(n374), .dout(n377));
  jnot g0063(.din(n377), .dout(n378));
  jxor g0064(.dina(n378), .dinb(G3717), .dout(n379));
  jor  g0065(.dina(n379), .dinb(n372), .dout(n380));
  jnot g0066(.din(G3711), .dout(n381));
  jand g0067(.dina(G237), .dinb(G18), .dout(n382));
  jnot g0068(.din(n382), .dout(n383));
  jnot g0069(.din(G26), .dout(n384));
  jor  g0070(.dina(n384), .dinb(G18), .dout(n385));
  jand g0071(.dina(n385), .dinb(n383), .dout(n386));
  jxor g0072(.dina(n386), .dinb(n381), .dout(n387));
  jnot g0073(.din(G4526), .dout(n388));
  jnot g0074(.din(G3701), .dout(n389));
  jand g0075(.dina(n356), .dinb(n389), .dout(n390));
  jnot g0076(.din(G229), .dout(n391));
  jor  g0077(.dina(n391), .dinb(n355), .dout(n392));
  jand g0078(.dina(n392), .dinb(n353), .dout(n393));
  jand g0079(.dina(n359), .dinb(n393), .dout(n394));
  jor  g0080(.dina(n394), .dinb(n390), .dout(n395));
  jnot g0081(.din(G3705), .dout(n396));
  jnot g0082(.din(G238), .dout(n397));
  jor  g0083(.dina(n397), .dinb(n355), .dout(n398));
  jnot g0084(.din(G29), .dout(n399));
  jor  g0085(.dina(n399), .dinb(G18), .dout(n400));
  jand g0086(.dina(n400), .dinb(n398), .dout(n401));
  jxor g0087(.dina(n401), .dinb(n396), .dout(n402));
  jor  g0088(.dina(n402), .dinb(n395), .dout(n403));
  jor  g0089(.dina(n403), .dinb(n388), .dout(n404));
  jor  g0090(.dina(n404), .dinb(n387), .dout(n405));
  jor  g0091(.dina(n405), .dinb(n380), .dout(n406));
  jor  g0092(.dina(n386), .dinb(G3711), .dout(n407));
  jor  g0093(.dina(n402), .dinb(n354), .dout(n408));
  jor  g0094(.dina(n408), .dinb(n387), .dout(n409));
  jand g0095(.dina(n409), .dinb(n407), .dout(n410));
  jor  g0096(.dina(n410), .dinb(n380), .dout(n411));
  jor  g0097(.dina(n401), .dinb(G3705), .dout(n412));
  jor  g0098(.dina(n412), .dinb(n387), .dout(n413));
  jor  g0099(.dina(n413), .dinb(n380), .dout(n414));
  jor  g0100(.dina(n371), .dinb(G3723), .dout(n415));
  jand g0101(.dina(n371), .dinb(G3723), .dout(n416));
  jor  g0102(.dina(n377), .dinb(G3717), .dout(n417));
  jor  g0103(.dina(n417), .dinb(n416), .dout(n418));
  jand g0104(.dina(n418), .dinb(n415), .dout(n419));
  jand g0105(.dina(n419), .dinb(n414), .dout(n420));
  jand g0106(.dina(n420), .dinb(n411), .dout(n421));
  jand g0107(.dina(n421), .dinb(n406), .dout(n422));
  jnot g0108(.din(G3737), .dout(n423));
  jand g0109(.dina(G233), .dinb(G18), .dout(n424));
  jnot g0110(.din(n424), .dout(n425));
  jnot g0111(.din(G127), .dout(n426));
  jor  g0112(.dina(n426), .dinb(G18), .dout(n427));
  jand g0113(.dina(n427), .dinb(n425), .dout(n428));
  jxor g0114(.dina(n428), .dinb(n423), .dout(n429));
  jnot g0115(.din(G3729), .dout(n430));
  jand g0116(.dina(G234), .dinb(G18), .dout(n431));
  jnot g0117(.din(n431), .dout(n432));
  jnot g0118(.din(G130), .dout(n433));
  jor  g0119(.dina(n433), .dinb(G18), .dout(n434));
  jand g0120(.dina(n434), .dinb(n432), .dout(n435));
  jxor g0121(.dina(n435), .dinb(n430), .dout(n436));
  jor  g0122(.dina(n436), .dinb(n429), .dout(n437));
  jand g0123(.dina(G231), .dinb(G18), .dout(n438));
  jnot g0124(.din(n438), .dout(n439));
  jnot g0125(.din(G100), .dout(n440));
  jor  g0126(.dina(n440), .dinb(G18), .dout(n441));
  jand g0127(.dina(n441), .dinb(n439), .dout(n442));
  jor  g0128(.dina(n442), .dinb(G3749), .dout(n443));
  jnot g0129(.din(n443), .dout(n444));
  jand g0130(.dina(n442), .dinb(G3749), .dout(n445));
  jor  g0131(.dina(n445), .dinb(n444), .dout(n446));
  jand g0132(.dina(G232), .dinb(G18), .dout(n447));
  jand g0133(.dina(G124), .dinb(n355), .dout(n448));
  jor  g0134(.dina(n448), .dinb(n447), .dout(n449));
  jxor g0135(.dina(n449), .dinb(G3743), .dout(n450));
  jor  g0136(.dina(n450), .dinb(n446), .dout(n451));
  jor  g0137(.dina(n451), .dinb(n437), .dout(n452));
  jor  g0138(.dina(n452), .dinb(n422), .dout(n453));
  jnot g0139(.din(n449), .dout(n454));
  jor  g0140(.dina(n454), .dinb(G3743), .dout(n455));
  jand g0141(.dina(n454), .dinb(G3743), .dout(n456));
  jor  g0142(.dina(n428), .dinb(G3737), .dout(n457));
  jor  g0143(.dina(n435), .dinb(G3729), .dout(n458));
  jor  g0144(.dina(n458), .dinb(n429), .dout(n459));
  jand g0145(.dina(n459), .dinb(n457), .dout(n460));
  jor  g0146(.dina(n460), .dinb(n456), .dout(n461));
  jand g0147(.dina(n461), .dinb(n455), .dout(n462));
  jand g0148(.dina(n462), .dinb(n443), .dout(n463));
  jor  g0149(.dina(n463), .dinb(n445), .dout(n464));
  jand g0150(.dina(n464), .dinb(n453), .dout(n465));
  jnot g0151(.din(G4415), .dout(n466));
  jand g0152(.dina(G223), .dinb(G18), .dout(n467));
  jand g0153(.dina(G47), .dinb(n355), .dout(n468));
  jor  g0154(.dina(n468), .dinb(n467), .dout(n469));
  jxor g0155(.dina(n469), .dinb(n466), .dout(n470));
  jnot g0156(.din(G4400), .dout(n471));
  jand g0157(.dina(G226), .dinb(G18), .dout(n472));
  jand g0158(.dina(G97), .dinb(n355), .dout(n473));
  jor  g0159(.dina(n473), .dinb(n472), .dout(n474));
  jxor g0160(.dina(n474), .dinb(n471), .dout(n475));
  jand g0161(.dina(G217), .dinb(G18), .dout(n476));
  jand g0162(.dina(G118), .dinb(n355), .dout(n477));
  jor  g0163(.dina(n477), .dinb(n476), .dout(n478));
  jnot g0164(.din(n478), .dout(n479));
  jxor g0165(.dina(n479), .dinb(G4394), .dout(n480));
  jand g0166(.dina(n480), .dinb(n475), .dout(n481));
  jnot g0167(.din(G4410), .dout(n482));
  jand g0168(.dina(G224), .dinb(G18), .dout(n483));
  jand g0169(.dina(G121), .dinb(n355), .dout(n484));
  jor  g0170(.dina(n484), .dinb(n483), .dout(n485));
  jxor g0171(.dina(n485), .dinb(n482), .dout(n486));
  jand g0172(.dina(G225), .dinb(G18), .dout(n487));
  jand g0173(.dina(G94), .dinb(n355), .dout(n488));
  jor  g0174(.dina(n488), .dinb(n487), .dout(n489));
  jnot g0175(.din(n489), .dout(n490));
  jxor g0176(.dina(n490), .dinb(G4405), .dout(n491));
  jand g0177(.dina(n491), .dinb(n486), .dout(n492));
  jand g0178(.dina(n492), .dinb(n481), .dout(n493));
  jand g0179(.dina(n493), .dinb(n470), .dout(n494));
  jnot g0180(.din(n494), .dout(n495));
  jor  g0181(.dina(n495), .dinb(n465), .dout(n496));
  jnot g0182(.din(n469), .dout(n497));
  jand g0183(.dina(n497), .dinb(G4415), .dout(n498));
  jand g0184(.dina(n469), .dinb(n466), .dout(n499));
  jnot g0185(.din(n499), .dout(n500));
  jand g0186(.dina(n485), .dinb(n482), .dout(n501));
  jnot g0187(.din(n501), .dout(n502));
  jnot g0188(.din(n485), .dout(n503));
  jand g0189(.dina(n503), .dinb(G4410), .dout(n504));
  jand g0190(.dina(n490), .dinb(G4405), .dout(n505));
  jnot g0191(.din(n475), .dout(n506));
  jor  g0192(.dina(n479), .dinb(G4394), .dout(n507));
  jor  g0193(.dina(n507), .dinb(n506), .dout(n508));
  jand g0194(.dina(n474), .dinb(n471), .dout(n509));
  jnot g0195(.din(n509), .dout(n510));
  jor  g0196(.dina(n490), .dinb(G4405), .dout(n511));
  jand g0197(.dina(n511), .dinb(n510), .dout(n512));
  jand g0198(.dina(n512), .dinb(n508), .dout(n513));
  jor  g0199(.dina(n513), .dinb(n505), .dout(n514));
  jor  g0200(.dina(n514), .dinb(n504), .dout(n515));
  jand g0201(.dina(n515), .dinb(n502), .dout(n516));
  jand g0202(.dina(n516), .dinb(n500), .dout(n517));
  jor  g0203(.dina(n517), .dinb(n498), .dout(n518));
  jand g0204(.dina(n518), .dinb(n496), .dout(n519));
  jnot g0205(.din(G4427), .dout(n520));
  jand g0206(.dina(G221), .dinb(G18), .dout(n521));
  jand g0207(.dina(G32), .dinb(n355), .dout(n522));
  jor  g0208(.dina(n522), .dinb(n521), .dout(n523));
  jxor g0209(.dina(n523), .dinb(n520), .dout(n524));
  jnot g0210(.din(G4420), .dout(n525));
  jand g0211(.dina(G222), .dinb(G18), .dout(n526));
  jand g0212(.dina(G35), .dinb(n355), .dout(n527));
  jor  g0213(.dina(n527), .dinb(n526), .dout(n528));
  jxor g0214(.dina(n528), .dinb(n525), .dout(n529));
  jand g0215(.dina(n529), .dinb(n524), .dout(n530));
  jnot g0216(.din(G4437), .dout(n531));
  jand g0217(.dina(G219), .dinb(G18), .dout(n532));
  jand g0218(.dina(G66), .dinb(n355), .dout(n533));
  jor  g0219(.dina(n533), .dinb(n532), .dout(n534));
  jxor g0220(.dina(n534), .dinb(n531), .dout(n535));
  jnot g0221(.din(G4432), .dout(n536));
  jand g0222(.dina(G220), .dinb(G18), .dout(n537));
  jand g0223(.dina(G50), .dinb(n355), .dout(n538));
  jor  g0224(.dina(n538), .dinb(n537), .dout(n539));
  jxor g0225(.dina(n539), .dinb(n536), .dout(n540));
  jand g0226(.dina(n540), .dinb(n535), .dout(n541));
  jand g0227(.dina(n541), .dinb(n530), .dout(n542));
  jnot g0228(.din(n542), .dout(n543));
  jor  g0229(.dina(n543), .dinb(n519), .dout(n544));
  jnot g0230(.din(n534), .dout(n545));
  jand g0231(.dina(n545), .dinb(G4437), .dout(n546));
  jnot g0232(.din(n546), .dout(n547));
  jand g0233(.dina(n534), .dinb(n531), .dout(n548));
  jand g0234(.dina(n539), .dinb(n536), .dout(n549));
  jnot g0235(.din(n539), .dout(n550));
  jand g0236(.dina(n550), .dinb(G4432), .dout(n551));
  jnot g0237(.din(n551), .dout(n552));
  jand g0238(.dina(n523), .dinb(n520), .dout(n553));
  jand g0239(.dina(n528), .dinb(n525), .dout(n554));
  jand g0240(.dina(n554), .dinb(n524), .dout(n555));
  jor  g0241(.dina(n555), .dinb(n553), .dout(n556));
  jand g0242(.dina(n556), .dinb(n552), .dout(n557));
  jor  g0243(.dina(n557), .dinb(n549), .dout(n558));
  jor  g0244(.dina(n558), .dinb(n548), .dout(n559));
  jand g0245(.dina(n559), .dinb(n547), .dout(n560));
  jnot g0246(.din(n560), .dout(n561));
  jand g0247(.dina(n561), .dinb(n544), .dout(n562));
  jnot g0248(.din(G2236), .dout(n563));
  jand g0249(.dina(G12), .dinb(G9), .dout(n564));
  jnot g0250(.din(n564), .dout(n565));
  jor  g0251(.dina(G157), .dinb(n355), .dout(n566));
  jand g0252(.dina(n566), .dinb(n565), .dout(n567));
  jxor g0253(.dina(n567), .dinb(n563), .dout(n568));
  jnot g0254(.din(G2218), .dout(n569));
  jand g0255(.dina(G138), .dinb(n355), .dout(n570));
  jand g0256(.dina(G160), .dinb(G18), .dout(n571));
  jor  g0257(.dina(n571), .dinb(n570), .dout(n572));
  jxor g0258(.dina(n572), .dinb(n569), .dout(n573));
  jnot g0259(.din(G2211), .dout(n574));
  jand g0260(.dina(G147), .dinb(n355), .dout(n575));
  jand g0261(.dina(G151), .dinb(G18), .dout(n576));
  jor  g0262(.dina(n576), .dinb(n575), .dout(n577));
  jxor g0263(.dina(n577), .dinb(n574), .dout(n578));
  jand g0264(.dina(n578), .dinb(n573), .dout(n579));
  jnot g0265(.din(G2230), .dout(n580));
  jand g0266(.dina(G135), .dinb(n355), .dout(n581));
  jand g0267(.dina(G158), .dinb(G18), .dout(n582));
  jor  g0268(.dina(n582), .dinb(n581), .dout(n583));
  jxor g0269(.dina(n583), .dinb(n580), .dout(n584));
  jnot g0270(.din(G2224), .dout(n585));
  jand g0271(.dina(G144), .dinb(n355), .dout(n586));
  jand g0272(.dina(G159), .dinb(G18), .dout(n587));
  jor  g0273(.dina(n587), .dinb(n586), .dout(n588));
  jxor g0274(.dina(n588), .dinb(n585), .dout(n589));
  jand g0275(.dina(n589), .dinb(n584), .dout(n590));
  jand g0276(.dina(n590), .dinb(n579), .dout(n591));
  jand g0277(.dina(n591), .dinb(n568), .dout(n592));
  jnot g0278(.din(n592), .dout(n593));
  jor  g0279(.dina(n593), .dinb(n562), .dout(n594));
  jand g0280(.dina(n567), .dinb(n563), .dout(n595));
  jnot g0281(.din(n595), .dout(n596));
  jnot g0282(.din(n567), .dout(n597));
  jand g0283(.dina(n597), .dinb(G2236), .dout(n598));
  jand g0284(.dina(n583), .dinb(n580), .dout(n599));
  jnot g0285(.din(n599), .dout(n600));
  jnot g0286(.din(n583), .dout(n601));
  jand g0287(.dina(n601), .dinb(G2230), .dout(n602));
  jnot g0288(.din(n588), .dout(n603));
  jand g0289(.dina(n603), .dinb(G2224), .dout(n604));
  jnot g0290(.din(n604), .dout(n605));
  jand g0291(.dina(n577), .dinb(n574), .dout(n606));
  jand g0292(.dina(n606), .dinb(n573), .dout(n607));
  jand g0293(.dina(n572), .dinb(n569), .dout(n608));
  jand g0294(.dina(n588), .dinb(n585), .dout(n609));
  jor  g0295(.dina(n609), .dinb(n608), .dout(n610));
  jor  g0296(.dina(n610), .dinb(n607), .dout(n611));
  jand g0297(.dina(n611), .dinb(n605), .dout(n612));
  jnot g0298(.din(n612), .dout(n613));
  jor  g0299(.dina(n613), .dinb(n602), .dout(n614));
  jand g0300(.dina(n614), .dinb(n600), .dout(n615));
  jor  g0301(.dina(n615), .dinb(n598), .dout(n616));
  jand g0302(.dina(n616), .dinb(n596), .dout(n617));
  jand g0303(.dina(n617), .dinb(n594), .dout(n618));
  jnot g0304(.din(G2247), .dout(n619));
  jor  g0305(.dina(G155), .dinb(n355), .dout(n620));
  jand g0306(.dina(n620), .dinb(n565), .dout(n621));
  jxor g0307(.dina(n621), .dinb(n619), .dout(n622));
  jnot g0308(.din(G2239), .dout(n623));
  jor  g0309(.dina(G156), .dinb(n355), .dout(n624));
  jand g0310(.dina(n624), .dinb(n565), .dout(n625));
  jxor g0311(.dina(n625), .dinb(n623), .dout(n626));
  jand g0312(.dina(n626), .dinb(n622), .dout(n627));
  jnot g0313(.din(G2256), .dout(n628));
  jor  g0314(.dina(G153), .dinb(n355), .dout(n629));
  jand g0315(.dina(n629), .dinb(n565), .dout(n630));
  jxor g0316(.dina(n630), .dinb(n628), .dout(n631));
  jnot g0317(.din(G2253), .dout(n632));
  jor  g0318(.dina(G154), .dinb(n355), .dout(n633));
  jand g0319(.dina(n633), .dinb(n565), .dout(n634));
  jxor g0320(.dina(n634), .dinb(n632), .dout(n635));
  jand g0321(.dina(n635), .dinb(n631), .dout(n636));
  jand g0322(.dina(n636), .dinb(n627), .dout(n637));
  jnot g0323(.din(n637), .dout(n638));
  jor  g0324(.dina(n638), .dinb(n618), .dout(n639));
  jand g0325(.dina(n630), .dinb(n628), .dout(n640));
  jnot g0326(.din(n640), .dout(n641));
  jand g0327(.dina(n634), .dinb(n632), .dout(n642));
  jnot g0328(.din(n642), .dout(n643));
  jand g0329(.dina(n621), .dinb(n619), .dout(n644));
  jand g0330(.dina(n625), .dinb(n623), .dout(n645));
  jand g0331(.dina(n645), .dinb(n622), .dout(n646));
  jor  g0332(.dina(n646), .dinb(n644), .dout(n647));
  jnot g0333(.din(n647), .dout(n648));
  jand g0334(.dina(n648), .dinb(n643), .dout(n649));
  jnot g0335(.din(n630), .dout(n650));
  jand g0336(.dina(n650), .dinb(G2256), .dout(n651));
  jnot g0337(.din(n634), .dout(n652));
  jand g0338(.dina(n652), .dinb(G2253), .dout(n653));
  jor  g0339(.dina(n653), .dinb(n651), .dout(n654));
  jor  g0340(.dina(n654), .dinb(n649), .dout(n655));
  jand g0341(.dina(n655), .dinb(n641), .dout(n656));
  jand g0342(.dina(n656), .dinb(n639), .dout(n657));
  jnot g0343(.din(G1486), .dout(n658));
  jor  g0344(.dina(G213), .dinb(n355), .dout(n659));
  jand g0345(.dina(n659), .dinb(n565), .dout(n660));
  jxor g0346(.dina(n660), .dinb(n658), .dout(n661));
  jnot g0347(.din(G1480), .dout(n662));
  jor  g0348(.dina(G214), .dinb(n355), .dout(n663));
  jand g0349(.dina(n663), .dinb(n565), .dout(n664));
  jxor g0350(.dina(n664), .dinb(n662), .dout(n665));
  jnot g0351(.din(G106), .dout(n666));
  jor  g0352(.dina(G215), .dinb(n355), .dout(n667));
  jand g0353(.dina(n667), .dinb(n565), .dout(n668));
  jxor g0354(.dina(n668), .dinb(n666), .dout(n669));
  jand g0355(.dina(n669), .dinb(n665), .dout(n670));
  jnot g0356(.din(G1469), .dout(n671));
  jor  g0357(.dina(G216), .dinb(n355), .dout(n672));
  jand g0358(.dina(n672), .dinb(n565), .dout(n673));
  jxor g0359(.dina(n673), .dinb(n671), .dout(n674));
  jnot g0360(.din(G1462), .dout(n675));
  jor  g0361(.dina(G209), .dinb(n355), .dout(n676));
  jand g0362(.dina(n676), .dinb(n565), .dout(n677));
  jxor g0363(.dina(n677), .dinb(n675), .dout(n678));
  jand g0364(.dina(n678), .dinb(n674), .dout(n679));
  jand g0365(.dina(n679), .dinb(n670), .dout(n680));
  jand g0366(.dina(n680), .dinb(n661), .dout(n681));
  jnot g0367(.din(n681), .dout(n682));
  jor  g0368(.dina(n682), .dinb(n657), .dout(n683));
  jand g0369(.dina(n660), .dinb(n658), .dout(n684));
  jor  g0370(.dina(n660), .dinb(n658), .dout(n685));
  jand g0371(.dina(n664), .dinb(n662), .dout(n686));
  jnot g0372(.din(n686), .dout(n687));
  jor  g0373(.dina(n664), .dinb(n662), .dout(n688));
  jand g0374(.dina(n668), .dinb(n666), .dout(n689));
  jnot g0375(.din(n668), .dout(n690));
  jand g0376(.dina(n690), .dinb(G106), .dout(n691));
  jnot g0377(.din(n691), .dout(n692));
  jnot g0378(.din(n673), .dout(n693));
  jand g0379(.dina(n693), .dinb(G1469), .dout(n694));
  jnot g0380(.din(n694), .dout(n695));
  jand g0381(.dina(n673), .dinb(n671), .dout(n696));
  jand g0382(.dina(n677), .dinb(n675), .dout(n697));
  jor  g0383(.dina(n697), .dinb(n696), .dout(n698));
  jand g0384(.dina(n698), .dinb(n695), .dout(n699));
  jand g0385(.dina(n699), .dinb(n692), .dout(n700));
  jor  g0386(.dina(n700), .dinb(n689), .dout(n701));
  jand g0387(.dina(n701), .dinb(n688), .dout(n702));
  jnot g0388(.din(n702), .dout(n703));
  jand g0389(.dina(n703), .dinb(n687), .dout(n704));
  jnot g0390(.din(n704), .dout(n705));
  jand g0391(.dina(n705), .dinb(n685), .dout(n706));
  jor  g0392(.dina(n706), .dinb(n684), .dout(n707));
  jnot g0393(.din(n707), .dout(n708));
  jand g0394(.dina(n708), .dinb(n683), .dout(n709));
  jnot g0395(.din(G38), .dout(n710));
  jand g0396(.dina(G4528), .dinb(G1492), .dout(n711));
  jxor g0397(.dina(n711), .dinb(n710), .dout(n712));
  jnot g0398(.din(n712), .dout(n713));
  jor  g0399(.dina(n713), .dinb(n709), .dout(n714));
  jor  g0400(.dina(n714), .dinb(n365), .dout(n715));
  jnot g0401(.din(n715), .dout(n716));
  jnot g0402(.din(G1492), .dout(n717));
  jnot g0403(.din(n364), .dout(n718));
  jor  g0404(.dina(n718), .dinb(n717), .dout(n719));
  jand g0405(.dina(n719), .dinb(G38), .dout(n720));
  jor  g0406(.dina(n720), .dinb(n716), .dout(G246));
  jor  g0407(.dina(G177), .dinb(n355), .dout(n722));
  jand g0408(.dina(n722), .dinb(n565), .dout(n723));
  jand g0409(.dina(G2236), .dinb(G18), .dout(n724));
  jnot g0410(.din(n724), .dout(n725));
  jor  g0411(.dina(G64), .dinb(G18), .dout(n726));
  jand g0412(.dina(n726), .dinb(n725), .dout(n727));
  jor  g0413(.dina(n727), .dinb(n723), .dout(n728));
  jand g0414(.dina(G178), .dinb(G18), .dout(n729));
  jor  g0415(.dina(n729), .dinb(n581), .dout(n730));
  jand g0416(.dina(G2230), .dinb(G18), .dout(n731));
  jnot g0417(.din(n731), .dout(n732));
  jor  g0418(.dina(G85), .dinb(G18), .dout(n733));
  jand g0419(.dina(n733), .dinb(n732), .dout(n734));
  jor  g0420(.dina(n734), .dinb(n730), .dout(n735));
  jand g0421(.dina(G179), .dinb(G18), .dout(n736));
  jor  g0422(.dina(n736), .dinb(n586), .dout(n737));
  jand g0423(.dina(G2224), .dinb(G18), .dout(n738));
  jnot g0424(.din(n738), .dout(n739));
  jor  g0425(.dina(G84), .dinb(G18), .dout(n740));
  jand g0426(.dina(n740), .dinb(n739), .dout(n741));
  jand g0427(.dina(n741), .dinb(n737), .dout(n742));
  jand g0428(.dina(G180), .dinb(G18), .dout(n743));
  jor  g0429(.dina(n743), .dinb(n570), .dout(n744));
  jand g0430(.dina(G2218), .dinb(G18), .dout(n745));
  jnot g0431(.din(n745), .dout(n746));
  jor  g0432(.dina(G83), .dinb(G18), .dout(n747));
  jand g0433(.dina(n747), .dinb(n746), .dout(n748));
  jor  g0434(.dina(n748), .dinb(n744), .dout(n749));
  jor  g0435(.dina(n741), .dinb(n737), .dout(n750));
  jand g0436(.dina(n750), .dinb(n749), .dout(n751));
  jand g0437(.dina(n748), .dinb(n744), .dout(n752));
  jand g0438(.dina(G171), .dinb(G18), .dout(n753));
  jor  g0439(.dina(n753), .dinb(n575), .dout(n754));
  jand g0440(.dina(G2211), .dinb(G18), .dout(n755));
  jnot g0441(.din(n755), .dout(n756));
  jor  g0442(.dina(G65), .dinb(G18), .dout(n757));
  jand g0443(.dina(n757), .dinb(n756), .dout(n758));
  jand g0444(.dina(n758), .dinb(n754), .dout(n759));
  jor  g0445(.dina(n759), .dinb(n752), .dout(n760));
  jand g0446(.dina(n760), .dinb(n751), .dout(n761));
  jor  g0447(.dina(n761), .dinb(n742), .dout(n762));
  jand g0448(.dina(n762), .dinb(n735), .dout(n763));
  jand g0449(.dina(n734), .dinb(n730), .dout(n764));
  jand g0450(.dina(n727), .dinb(n723), .dout(n765));
  jor  g0451(.dina(n765), .dinb(n764), .dout(n766));
  jor  g0452(.dina(n766), .dinb(n763), .dout(n767));
  jand g0453(.dina(n767), .dinb(n728), .dout(n768));
  jnot g0454(.din(n752), .dout(n769));
  jand g0455(.dina(n769), .dinb(n735), .dout(n770));
  jnot g0456(.din(n742), .dout(n771));
  jnot g0457(.din(n759), .dout(n772));
  jand g0458(.dina(n772), .dinb(n771), .dout(n773));
  jand g0459(.dina(n773), .dinb(n770), .dout(n774));
  jnot g0460(.din(n765), .dout(n775));
  jor  g0461(.dina(n758), .dinb(n754), .dout(n776));
  jand g0462(.dina(n776), .dinb(n775), .dout(n777));
  jnot g0463(.din(n764), .dout(n778));
  jand g0464(.dina(n778), .dinb(n728), .dout(n779));
  jand g0465(.dina(n779), .dinb(n777), .dout(n780));
  jand g0466(.dina(n780), .dinb(n751), .dout(n781));
  jand g0467(.dina(n781), .dinb(n774), .dout(n782));
  jand g0468(.dina(G191), .dinb(G18), .dout(n783));
  jor  g0469(.dina(n783), .dinb(n522), .dout(n784));
  jor  g0470(.dina(G60), .dinb(G18), .dout(n785));
  jor  g0471(.dina(n520), .dinb(n355), .dout(n786));
  jand g0472(.dina(n786), .dinb(n785), .dout(n787));
  jxor g0473(.dina(n787), .dinb(n784), .dout(n788));
  jand g0474(.dina(G189), .dinb(G18), .dout(n789));
  jor  g0475(.dina(n789), .dinb(n533), .dout(n790));
  jor  g0476(.dina(G62), .dinb(G18), .dout(n791));
  jor  g0477(.dina(n531), .dinb(n355), .dout(n792));
  jand g0478(.dina(n792), .dinb(n791), .dout(n793));
  jxor g0479(.dina(n793), .dinb(n790), .dout(n794));
  jand g0480(.dina(n794), .dinb(n788), .dout(n795));
  jand g0481(.dina(G190), .dinb(G18), .dout(n796));
  jor  g0482(.dina(n796), .dinb(n538), .dout(n797));
  jor  g0483(.dina(G61), .dinb(G18), .dout(n798));
  jand g0484(.dina(G4432), .dinb(G18), .dout(n799));
  jnot g0485(.din(n799), .dout(n800));
  jand g0486(.dina(n800), .dinb(n798), .dout(n801));
  jxor g0487(.dina(n801), .dinb(n797), .dout(n802));
  jand g0488(.dina(G192), .dinb(G18), .dout(n803));
  jor  g0489(.dina(n803), .dinb(n527), .dout(n804));
  jor  g0490(.dina(G79), .dinb(G18), .dout(n805));
  jor  g0491(.dina(n525), .dinb(n355), .dout(n806));
  jand g0492(.dina(n806), .dinb(n805), .dout(n807));
  jxor g0493(.dina(n807), .dinb(n804), .dout(n808));
  jand g0494(.dina(n808), .dinb(n802), .dout(n809));
  jand g0495(.dina(n809), .dinb(n795), .dout(n810));
  jand g0496(.dina(G196), .dinb(G18), .dout(n811));
  jor  g0497(.dina(n811), .dinb(n473), .dout(n812));
  jor  g0498(.dina(G78), .dinb(G18), .dout(n813));
  jand g0499(.dina(G4400), .dinb(G18), .dout(n814));
  jnot g0500(.din(n814), .dout(n815));
  jand g0501(.dina(n815), .dinb(n813), .dout(n816));
  jor  g0502(.dina(n816), .dinb(n812), .dout(n817));
  jand g0503(.dina(G195), .dinb(G18), .dout(n818));
  jor  g0504(.dina(n818), .dinb(n488), .dout(n819));
  jor  g0505(.dina(G59), .dinb(G18), .dout(n820));
  jand g0506(.dina(G4405), .dinb(G18), .dout(n821));
  jnot g0507(.din(n821), .dout(n822));
  jand g0508(.dina(n822), .dinb(n820), .dout(n823));
  jor  g0509(.dina(n823), .dinb(n819), .dout(n824));
  jand g0510(.dina(n824), .dinb(n817), .dout(n825));
  jand g0511(.dina(G187), .dinb(G18), .dout(n826));
  jor  g0512(.dina(n826), .dinb(n477), .dout(n827));
  jor  g0513(.dina(G77), .dinb(G18), .dout(n828));
  jand g0514(.dina(G4394), .dinb(G18), .dout(n829));
  jnot g0515(.din(n829), .dout(n830));
  jand g0516(.dina(n830), .dinb(n828), .dout(n831));
  jand g0517(.dina(n831), .dinb(n827), .dout(n832));
  jnot g0518(.din(n832), .dout(n833));
  jand g0519(.dina(n823), .dinb(n819), .dout(n834));
  jnot g0520(.din(n834), .dout(n835));
  jand g0521(.dina(n835), .dinb(n833), .dout(n836));
  jand g0522(.dina(n836), .dinb(n825), .dout(n837));
  jand g0523(.dina(n816), .dinb(n812), .dout(n838));
  jnot g0524(.din(n838), .dout(n839));
  jor  g0525(.dina(n831), .dinb(n827), .dout(n840));
  jand g0526(.dina(n840), .dinb(n839), .dout(n841));
  jand g0527(.dina(G193), .dinb(G18), .dout(n842));
  jor  g0528(.dina(n842), .dinb(n468), .dout(n843));
  jor  g0529(.dina(G80), .dinb(G18), .dout(n844));
  jand g0530(.dina(G4415), .dinb(G18), .dout(n845));
  jnot g0531(.din(n845), .dout(n846));
  jand g0532(.dina(n846), .dinb(n844), .dout(n847));
  jand g0533(.dina(n847), .dinb(n843), .dout(n848));
  jnot g0534(.din(n848), .dout(n849));
  jand g0535(.dina(G194), .dinb(G18), .dout(n850));
  jor  g0536(.dina(n850), .dinb(n484), .dout(n851));
  jor  g0537(.dina(G81), .dinb(G18), .dout(n852));
  jand g0538(.dina(G4410), .dinb(G18), .dout(n853));
  jnot g0539(.din(n853), .dout(n854));
  jand g0540(.dina(n854), .dinb(n852), .dout(n855));
  jor  g0541(.dina(n855), .dinb(n851), .dout(n856));
  jand g0542(.dina(n856), .dinb(n849), .dout(n857));
  jor  g0543(.dina(n847), .dinb(n843), .dout(n858));
  jand g0544(.dina(n855), .dinb(n851), .dout(n859));
  jnot g0545(.din(n859), .dout(n860));
  jand g0546(.dina(n860), .dinb(n858), .dout(n861));
  jand g0547(.dina(n861), .dinb(n857), .dout(n862));
  jand g0548(.dina(n862), .dinb(n841), .dout(n863));
  jand g0549(.dina(n863), .dinb(n837), .dout(n864));
  jand g0550(.dina(n864), .dinb(n810), .dout(n865));
  jand g0551(.dina(G200), .dinb(G18), .dout(n866));
  jnot g0552(.din(n866), .dout(n867));
  jand g0553(.dina(n867), .dinb(n441), .dout(n868));
  jnot g0554(.din(n868), .dout(n869));
  jor  g0555(.dina(G56), .dinb(G18), .dout(n870));
  jand g0556(.dina(G3749), .dinb(G18), .dout(n871));
  jnot g0557(.din(n871), .dout(n872));
  jand g0558(.dina(n872), .dinb(n870), .dout(n873));
  jand g0559(.dina(n873), .dinb(n869), .dout(n874));
  jnot g0560(.din(n874), .dout(n875));
  jnot g0561(.din(n427), .dout(n876));
  jand g0562(.dina(G202), .dinb(G18), .dout(n877));
  jor  g0563(.dina(n877), .dinb(n876), .dout(n878));
  jor  g0564(.dina(G54), .dinb(G18), .dout(n879));
  jand g0565(.dina(G3737), .dinb(G18), .dout(n880));
  jnot g0566(.din(n880), .dout(n881));
  jand g0567(.dina(n881), .dinb(n879), .dout(n882));
  jor  g0568(.dina(n882), .dinb(n878), .dout(n883));
  jand g0569(.dina(n883), .dinb(n875), .dout(n884));
  jand g0570(.dina(n882), .dinb(n878), .dout(n885));
  jnot g0571(.din(n885), .dout(n886));
  jor  g0572(.dina(n873), .dinb(n869), .dout(n887));
  jand g0573(.dina(n887), .dinb(n886), .dout(n888));
  jand g0574(.dina(n888), .dinb(n884), .dout(n889));
  jand g0575(.dina(G201), .dinb(G18), .dout(n890));
  jor  g0576(.dina(n890), .dinb(n448), .dout(n891));
  jor  g0577(.dina(G55), .dinb(G18), .dout(n892));
  jand g0578(.dina(G3743), .dinb(G18), .dout(n893));
  jnot g0579(.din(n893), .dout(n894));
  jand g0580(.dina(n894), .dinb(n892), .dout(n895));
  jxor g0581(.dina(n895), .dinb(n891), .dout(n896));
  jnot g0582(.din(n434), .dout(n897));
  jand g0583(.dina(G203), .dinb(G18), .dout(n898));
  jor  g0584(.dina(n898), .dinb(n897), .dout(n899));
  jor  g0585(.dina(G53), .dinb(G18), .dout(n900));
  jor  g0586(.dina(n430), .dinb(n355), .dout(n901));
  jand g0587(.dina(n901), .dinb(n900), .dout(n902));
  jxor g0588(.dina(n902), .dinb(n899), .dout(n903));
  jand g0589(.dina(n903), .dinb(n896), .dout(n904));
  jand g0590(.dina(n904), .dinb(n889), .dout(n905));
  jnot g0591(.din(n400), .dout(n906));
  jand g0592(.dina(G207), .dinb(G18), .dout(n907));
  jor  g0593(.dina(n907), .dinb(n906), .dout(n908));
  jor  g0594(.dina(G74), .dinb(G18), .dout(n909));
  jand g0595(.dina(G3705), .dinb(G18), .dout(n910));
  jnot g0596(.din(n910), .dout(n911));
  jand g0597(.dina(n911), .dinb(n909), .dout(n912));
  jor  g0598(.dina(n912), .dinb(n908), .dout(n913));
  jnot g0599(.din(n376), .dout(n914));
  jand g0600(.dina(G205), .dinb(G18), .dout(n915));
  jor  g0601(.dina(n915), .dinb(n914), .dout(n916));
  jor  g0602(.dina(G75), .dinb(G18), .dout(n917));
  jand g0603(.dina(G3717), .dinb(G18), .dout(n918));
  jnot g0604(.din(n918), .dout(n919));
  jand g0605(.dina(n919), .dinb(n917), .dout(n920));
  jor  g0606(.dina(n920), .dinb(n916), .dout(n921));
  jand g0607(.dina(n921), .dinb(n913), .dout(n922));
  jand g0608(.dina(n920), .dinb(n916), .dout(n923));
  jnot g0609(.din(n923), .dout(n924));
  jnot g0610(.din(n385), .dout(n925));
  jand g0611(.dina(G206), .dinb(G18), .dout(n926));
  jor  g0612(.dina(n926), .dinb(n925), .dout(n927));
  jor  g0613(.dina(G76), .dinb(G18), .dout(n928));
  jand g0614(.dina(G3711), .dinb(G18), .dout(n929));
  jnot g0615(.din(n929), .dout(n930));
  jand g0616(.dina(n930), .dinb(n928), .dout(n931));
  jor  g0617(.dina(n931), .dinb(n927), .dout(n932));
  jand g0618(.dina(n932), .dinb(n924), .dout(n933));
  jand g0619(.dina(n933), .dinb(n922), .dout(n934));
  jnot g0620(.din(G70), .dout(n935));
  jand g0621(.dina(n935), .dinb(n355), .dout(n936));
  jnot g0622(.din(n936), .dout(n937));
  jor  g0623(.dina(n937), .dinb(G41), .dout(n938));
  jand g0624(.dina(n937), .dinb(n356), .dout(n939));
  jnot g0625(.din(n939), .dout(n940));
  jand g0626(.dina(n940), .dinb(G89), .dout(n941));
  jand g0627(.dina(n941), .dinb(n938), .dout(n942));
  jnot g0628(.din(n370), .dout(n943));
  jand g0629(.dina(G204), .dinb(G18), .dout(n944));
  jor  g0630(.dina(n944), .dinb(n943), .dout(n945));
  jor  g0631(.dina(G73), .dinb(G18), .dout(n946));
  jor  g0632(.dina(n366), .dinb(n355), .dout(n947));
  jand g0633(.dina(n947), .dinb(n946), .dout(n948));
  jxor g0634(.dina(n948), .dinb(n945), .dout(n949));
  jand g0635(.dina(n912), .dinb(n908), .dout(n950));
  jnot g0636(.din(n950), .dout(n951));
  jand g0637(.dina(n931), .dinb(n927), .dout(n952));
  jnot g0638(.din(n952), .dout(n953));
  jand g0639(.dina(n953), .dinb(n951), .dout(n954));
  jand g0640(.dina(n954), .dinb(n949), .dout(n955));
  jand g0641(.dina(n955), .dinb(n942), .dout(n956));
  jand g0642(.dina(n956), .dinb(n934), .dout(n957));
  jand g0643(.dina(n957), .dinb(n905), .dout(n958));
  jand g0644(.dina(n958), .dinb(n865), .dout(n959));
  jand g0645(.dina(n807), .dinb(n804), .dout(n960));
  jand g0646(.dina(n960), .dinb(n802), .dout(n961));
  jand g0647(.dina(n961), .dinb(n795), .dout(n962));
  jand g0648(.dina(n793), .dinb(n790), .dout(n963));
  jand g0649(.dina(n787), .dinb(n784), .dout(n964));
  jand g0650(.dina(n801), .dinb(n797), .dout(n965));
  jor  g0651(.dina(n965), .dinb(n964), .dout(n966));
  jor  g0652(.dina(n793), .dinb(n790), .dout(n967));
  jor  g0653(.dina(n801), .dinb(n797), .dout(n968));
  jand g0654(.dina(n968), .dinb(n967), .dout(n969));
  jand g0655(.dina(n969), .dinb(n966), .dout(n970));
  jor  g0656(.dina(n970), .dinb(n963), .dout(n971));
  jor  g0657(.dina(n971), .dinb(n962), .dout(n972));
  jand g0658(.dina(n832), .dinb(n817), .dout(n973));
  jor  g0659(.dina(n838), .dinb(n834), .dout(n974));
  jor  g0660(.dina(n974), .dinb(n973), .dout(n975));
  jand g0661(.dina(n858), .dinb(n856), .dout(n976));
  jand g0662(.dina(n976), .dinb(n824), .dout(n977));
  jand g0663(.dina(n977), .dinb(n975), .dout(n978));
  jand g0664(.dina(n859), .dinb(n858), .dout(n979));
  jor  g0665(.dina(n979), .dinb(n848), .dout(n980));
  jor  g0666(.dina(n980), .dinb(n978), .dout(n981));
  jand g0667(.dina(n981), .dinb(n810), .dout(n982));
  jor  g0668(.dina(n982), .dinb(n972), .dout(n983));
  jor  g0669(.dina(n983), .dinb(n959), .dout(n984));
  jand g0670(.dina(n984), .dinb(n782), .dout(n985));
  jor  g0671(.dina(n985), .dinb(n768), .dout(n986));
  jor  g0672(.dina(G173), .dinb(n355), .dout(n987));
  jand g0673(.dina(n987), .dinb(n565), .dout(n988));
  jand g0674(.dina(G2256), .dinb(G18), .dout(n989));
  jnot g0675(.din(n989), .dout(n990));
  jor  g0676(.dina(G110), .dinb(G18), .dout(n991));
  jand g0677(.dina(n991), .dinb(n990), .dout(n992));
  jor  g0678(.dina(n992), .dinb(n988), .dout(n993));
  jor  g0679(.dina(G175), .dinb(n355), .dout(n994));
  jand g0680(.dina(n994), .dinb(n565), .dout(n995));
  jand g0681(.dina(G2247), .dinb(G18), .dout(n996));
  jnot g0682(.din(n996), .dout(n997));
  jor  g0683(.dina(G86), .dinb(G18), .dout(n998));
  jand g0684(.dina(n998), .dinb(n997), .dout(n999));
  jand g0685(.dina(n999), .dinb(n995), .dout(n1000));
  jnot g0686(.din(n1000), .dout(n1001));
  jand g0687(.dina(n1001), .dinb(n993), .dout(n1002));
  jand g0688(.dina(n992), .dinb(n988), .dout(n1003));
  jnot g0689(.din(n1003), .dout(n1004));
  jor  g0690(.dina(n999), .dinb(n995), .dout(n1005));
  jand g0691(.dina(n1005), .dinb(n1004), .dout(n1006));
  jand g0692(.dina(n1006), .dinb(n1002), .dout(n1007));
  jor  g0693(.dina(G174), .dinb(n355), .dout(n1008));
  jand g0694(.dina(n1008), .dinb(n565), .dout(n1009));
  jand g0695(.dina(G2253), .dinb(G18), .dout(n1010));
  jnot g0696(.din(n1010), .dout(n1011));
  jor  g0697(.dina(G109), .dinb(G18), .dout(n1012));
  jand g0698(.dina(n1012), .dinb(n1011), .dout(n1013));
  jxor g0699(.dina(n1013), .dinb(n1009), .dout(n1014));
  jor  g0700(.dina(G176), .dinb(n355), .dout(n1015));
  jand g0701(.dina(n1015), .dinb(n565), .dout(n1016));
  jor  g0702(.dina(n623), .dinb(n355), .dout(n1017));
  jor  g0703(.dina(G63), .dinb(G18), .dout(n1018));
  jand g0704(.dina(n1018), .dinb(n1017), .dout(n1019));
  jxor g0705(.dina(n1019), .dinb(n1016), .dout(n1020));
  jand g0706(.dina(n1020), .dinb(n1014), .dout(n1021));
  jand g0707(.dina(n1021), .dinb(n1007), .dout(n1022));
  jand g0708(.dina(n1022), .dinb(n986), .dout(n1023));
  jand g0709(.dina(n948), .dinb(n945), .dout(n1024));
  jor  g0710(.dina(n950), .dinb(n939), .dout(n1025));
  jand g0711(.dina(n932), .dinb(n913), .dout(n1026));
  jand g0712(.dina(n1026), .dinb(n1025), .dout(n1027));
  jor  g0713(.dina(n952), .dinb(n923), .dout(n1028));
  jor  g0714(.dina(n1028), .dinb(n1027), .dout(n1029));
  jor  g0715(.dina(n948), .dinb(n945), .dout(n1030));
  jand g0716(.dina(n1030), .dinb(n921), .dout(n1031));
  jand g0717(.dina(n1031), .dinb(n1029), .dout(n1032));
  jor  g0718(.dina(n1032), .dinb(n1024), .dout(n1033));
  jand g0719(.dina(n1033), .dinb(n905), .dout(n1034));
  jand g0720(.dina(n902), .dinb(n899), .dout(n1035));
  jand g0721(.dina(n1035), .dinb(n896), .dout(n1036));
  jand g0722(.dina(n1036), .dinb(n889), .dout(n1037));
  jand g0723(.dina(n895), .dinb(n891), .dout(n1038));
  jor  g0724(.dina(n1038), .dinb(n885), .dout(n1039));
  jor  g0725(.dina(n895), .dinb(n891), .dout(n1040));
  jand g0726(.dina(n1040), .dinb(n887), .dout(n1041));
  jand g0727(.dina(n1041), .dinb(n1039), .dout(n1042));
  jor  g0728(.dina(n1042), .dinb(n874), .dout(n1043));
  jor  g0729(.dina(n1043), .dinb(n1037), .dout(n1044));
  jor  g0730(.dina(n1044), .dinb(n1034), .dout(n1045));
  jand g0731(.dina(n1022), .dinb(n782), .dout(n1046));
  jand g0732(.dina(n1046), .dinb(n865), .dout(n1047));
  jand g0733(.dina(n1047), .dinb(n1045), .dout(n1048));
  jand g0734(.dina(n1019), .dinb(n1016), .dout(n1049));
  jand g0735(.dina(n1049), .dinb(n1014), .dout(n1050));
  jand g0736(.dina(n1050), .dinb(n1007), .dout(n1051));
  jand g0737(.dina(n1013), .dinb(n1009), .dout(n1052));
  jor  g0738(.dina(n1052), .dinb(n1000), .dout(n1053));
  jor  g0739(.dina(n1013), .dinb(n1009), .dout(n1054));
  jand g0740(.dina(n1054), .dinb(n993), .dout(n1055));
  jand g0741(.dina(n1055), .dinb(n1053), .dout(n1056));
  jor  g0742(.dina(n1056), .dinb(n1003), .dout(n1057));
  jor  g0743(.dina(n1057), .dinb(n1051), .dout(n1058));
  jor  g0744(.dina(n1058), .dinb(n1048), .dout(n1059));
  jor  g0745(.dina(n1059), .dinb(n1023), .dout(n1060));
  jor  g0746(.dina(G167), .dinb(n355), .dout(n1061));
  jand g0747(.dina(n1061), .dinb(n565), .dout(n1062));
  jand g0748(.dina(G1480), .dinb(G18), .dout(n1063));
  jnot g0749(.din(n1063), .dout(n1064));
  jor  g0750(.dina(G112), .dinb(G18), .dout(n1065));
  jand g0751(.dina(n1065), .dinb(n1064), .dout(n1066));
  jor  g0752(.dina(n1066), .dinb(n1062), .dout(n1067));
  jor  g0753(.dina(G166), .dinb(n355), .dout(n1068));
  jand g0754(.dina(n1068), .dinb(n565), .dout(n1069));
  jand g0755(.dina(G1486), .dinb(G18), .dout(n1070));
  jnot g0756(.din(n1070), .dout(n1071));
  jor  g0757(.dina(G88), .dinb(G18), .dout(n1072));
  jand g0758(.dina(n1072), .dinb(n1071), .dout(n1073));
  jor  g0759(.dina(n1073), .dinb(n1069), .dout(n1074));
  jand g0760(.dina(n1074), .dinb(n1067), .dout(n1075));
  jor  g0761(.dina(G169), .dinb(n355), .dout(n1076));
  jand g0762(.dina(n1076), .dinb(n565), .dout(n1077));
  jand g0763(.dina(G1469), .dinb(G18), .dout(n1078));
  jnot g0764(.din(n1078), .dout(n1079));
  jor  g0765(.dina(G111), .dinb(G18), .dout(n1080));
  jand g0766(.dina(n1080), .dinb(n1079), .dout(n1081));
  jor  g0767(.dina(n1081), .dinb(n1077), .dout(n1082));
  jand g0768(.dina(G1462), .dinb(G18), .dout(n1083));
  jnot g0769(.din(n1083), .dout(n1084));
  jor  g0770(.dina(G113), .dinb(G18), .dout(n1085));
  jand g0771(.dina(n1085), .dinb(n1084), .dout(n1086));
  jor  g0772(.dina(n1086), .dinb(n565), .dout(n1087));
  jand g0773(.dina(n1087), .dinb(n1082), .dout(n1088));
  jand g0774(.dina(n1088), .dinb(n1075), .dout(n1089));
  jand g0775(.dina(n1081), .dinb(n1077), .dout(n1090));
  jand g0776(.dina(n1086), .dinb(n565), .dout(n1091));
  jor  g0777(.dina(n1091), .dinb(n1090), .dout(n1092));
  jnot g0778(.din(n1092), .dout(n1093));
  jand g0779(.dina(n1066), .dinb(n1062), .dout(n1094));
  jor  g0780(.dina(G168), .dinb(n355), .dout(n1095));
  jand g0781(.dina(n1095), .dinb(n565), .dout(n1096));
  jand g0782(.dina(G106), .dinb(G18), .dout(n1097));
  jnot g0783(.din(n1097), .dout(n1098));
  jor  g0784(.dina(G87), .dinb(G18), .dout(n1099));
  jand g0785(.dina(n1099), .dinb(n1098), .dout(n1100));
  jand g0786(.dina(n1100), .dinb(n1096), .dout(n1101));
  jor  g0787(.dina(n1101), .dinb(n1094), .dout(n1102));
  jnot g0788(.din(n1102), .dout(n1103));
  jor  g0789(.dina(n1100), .dinb(n1096), .dout(n1104));
  jand g0790(.dina(n1073), .dinb(n1069), .dout(n1105));
  jnot g0791(.din(n1105), .dout(n1106));
  jand g0792(.dina(n1106), .dinb(n1104), .dout(n1107));
  jand g0793(.dina(n1107), .dinb(n1103), .dout(n1108));
  jand g0794(.dina(n1108), .dinb(n1093), .dout(n1109));
  jand g0795(.dina(n1109), .dinb(n1089), .dout(n1110));
  jand g0796(.dina(n1110), .dinb(n1060), .dout(n1111));
  jand g0797(.dina(n1104), .dinb(n1082), .dout(n1112));
  jand g0798(.dina(n1112), .dinb(n1092), .dout(n1113));
  jor  g0799(.dina(n1113), .dinb(n1102), .dout(n1114));
  jand g0800(.dina(n1114), .dinb(n1075), .dout(n1115));
  jnot g0801(.din(G4528), .dout(n1116));
  jor  g0802(.dina(G2204), .dinb(G1455), .dout(n1117));
  jor  g0803(.dina(n1117), .dinb(n1116), .dout(n1118));
  jand g0804(.dina(n1118), .dinb(G38), .dout(n1119));
  jor  g0805(.dina(n1119), .dinb(n1105), .dout(n1120));
  jor  g0806(.dina(n1120), .dinb(n1115), .dout(n1121));
  jor  g0807(.dina(n1121), .dinb(n1111), .dout(n1122));
  jand g0808(.dina(G2204), .dinb(G1455), .dout(n1123));
  jor  g0809(.dina(n1116), .dinb(G38), .dout(n1124));
  jor  g0810(.dina(n1124), .dinb(n1123), .dout(n1125));
  jand g0811(.dina(n1125), .dinb(n1122), .dout(G258));
  jand g0812(.dina(n377), .dinb(G3717), .dout(n1127));
  jand g0813(.dina(n413), .dinb(n410), .dout(n1128));
  jor  g0814(.dina(n1128), .dinb(n1127), .dout(n1129));
  jand g0815(.dina(n1129), .dinb(n417), .dout(n1130));
  jor  g0816(.dina(n405), .dinb(n379), .dout(n1131));
  jand g0817(.dina(n1131), .dinb(n1130), .dout(n1132));
  jxor g0818(.dina(n1132), .dinb(n372), .dout(G388));
  jand g0819(.dina(n1128), .dinb(n405), .dout(n1134));
  jxor g0820(.dina(n1134), .dinb(n379), .dout(G391));
  jand g0821(.dina(n408), .dinb(n412), .dout(n1136));
  jand g0822(.dina(n1136), .dinb(n404), .dout(n1137));
  jxor g0823(.dina(n1137), .dinb(n387), .dout(G394));
  jor  g0824(.dina(n395), .dinb(n388), .dout(n1139));
  jand g0825(.dina(n1139), .dinb(n354), .dout(n1140));
  jxor g0826(.dina(n1140), .dinb(n402), .dout(G397));
  jor  g0827(.dina(n437), .dinb(n422), .dout(n1142));
  jor  g0828(.dina(n1142), .dinb(n456), .dout(n1143));
  jand g0829(.dina(n1143), .dinb(n462), .dout(n1144));
  jxor g0830(.dina(n1144), .dinb(n446), .dout(G376));
  jand g0831(.dina(n1142), .dinb(n460), .dout(n1146));
  jxor g0832(.dina(n1146), .dinb(n450), .dout(G379));
  jand g0833(.dina(n435), .dinb(G3729), .dout(n1148));
  jor  g0834(.dina(n1148), .dinb(n422), .dout(n1149));
  jand g0835(.dina(n1149), .dinb(n458), .dout(n1150));
  jxor g0836(.dina(n1150), .dinb(n429), .dout(G382));
  jxor g0837(.dina(n436), .dinb(n422), .dout(G385));
  jxor g0838(.dina(n583), .dinb(n577), .dout(n1153));
  jxor g0839(.dina(n588), .dinb(n567), .dout(n1154));
  jxor g0840(.dina(n1154), .dinb(n572), .dout(n1155));
  jnot g0841(.din(n625), .dout(n1156));
  jor  g0842(.dina(n1156), .dinb(n620), .dout(n1157));
  jnot g0843(.din(n621), .dout(n1158));
  jor  g0844(.dina(n624), .dinb(n1158), .dout(n1159));
  jand g0845(.dina(n1159), .dinb(n1157), .dout(n1160));
  jor  g0846(.dina(n652), .dinb(n629), .dout(n1161));
  jor  g0847(.dina(n633), .dinb(n650), .dout(n1162));
  jand g0848(.dina(n1162), .dinb(n1161), .dout(n1163));
  jxor g0849(.dina(n1163), .dinb(n1160), .dout(n1164));
  jnot g0850(.din(G141), .dout(n1165));
  jor  g0851(.dina(n1165), .dinb(G18), .dout(n1166));
  jnot g0852(.din(G161), .dout(n1167));
  jor  g0853(.dina(n1167), .dinb(n355), .dout(n1168));
  jand g0854(.dina(n1168), .dinb(n1166), .dout(n1169));
  jxor g0855(.dina(n1169), .dinb(n1164), .dout(n1170));
  jxor g0856(.dina(n1170), .dinb(n1155), .dout(n1171));
  jxor g0857(.dina(n1171), .dinb(n1153), .dout(n1172));
  jand g0858(.dina(n565), .dinb(G18), .dout(n1173));
  jxor g0859(.dina(G212), .dinb(G211), .dout(n1174));
  jand g0860(.dina(n1174), .dinb(n1173), .dout(n1175));
  jor  g0861(.dina(n676), .dinb(n564), .dout(n1176));
  jnot g0862(.din(n659), .dout(n1177));
  jand g0863(.dina(n664), .dinb(n1177), .dout(n1178));
  jnot g0864(.din(n663), .dout(n1179));
  jand g0865(.dina(n1179), .dinb(n660), .dout(n1180));
  jor  g0866(.dina(n1180), .dinb(n1178), .dout(n1181));
  jor  g0867(.dina(n693), .dinb(n667), .dout(n1182));
  jor  g0868(.dina(n672), .dinb(n690), .dout(n1183));
  jand g0869(.dina(n1183), .dinb(n1182), .dout(n1184));
  jxor g0870(.dina(n1184), .dinb(n1181), .dout(n1185));
  jxor g0871(.dina(n1185), .dinb(n1176), .dout(n1186));
  jxor g0872(.dina(n1186), .dinb(n1175), .dout(n1187));
  jand g0873(.dina(G239), .dinb(G18), .dout(n1188));
  jand g0874(.dina(G44), .dinb(n355), .dout(n1189));
  jor  g0875(.dina(n1189), .dinb(n1188), .dout(n1190));
  jxor g0876(.dina(n442), .dinb(n428), .dout(n1191));
  jxor g0877(.dina(n449), .dinb(n435), .dout(n1192));
  jxor g0878(.dina(n1192), .dinb(n1191), .dout(n1193));
  jxor g0879(.dina(n1193), .dinb(n1190), .dout(n1194));
  jxor g0880(.dina(n401), .dinb(n371), .dout(n1195));
  jxor g0881(.dina(n1195), .dinb(n377), .dout(n1196));
  jxor g0882(.dina(n386), .dinb(n358), .dout(n1197));
  jxor g0883(.dina(n1197), .dinb(n1196), .dout(n1198));
  jxor g0884(.dina(n1198), .dinb(n1194), .dout(n1199));
  jxor g0885(.dina(n534), .dinb(n523), .dout(n1200));
  jxor g0886(.dina(n539), .dinb(n528), .dout(n1201));
  jxor g0887(.dina(n1201), .dinb(n1200), .dout(n1202));
  jxor g0888(.dina(n1202), .dinb(n503), .dout(n1203));
  jand g0889(.dina(G227), .dinb(G18), .dout(n1204));
  jand g0890(.dina(G115), .dinb(n355), .dout(n1205));
  jor  g0891(.dina(n1205), .dinb(n1204), .dout(n1206));
  jxor g0892(.dina(n489), .dinb(n478), .dout(n1207));
  jxor g0893(.dina(n1207), .dinb(n1206), .dout(n1208));
  jxor g0894(.dina(n474), .dinb(n469), .dout(n1209));
  jxor g0895(.dina(n1209), .dinb(n1208), .dout(n1210));
  jxor g0896(.dina(n1210), .dinb(n1203), .dout(n1211));
  jor  g0897(.dina(n1211), .dinb(n1199), .dout(n1212));
  jor  g0898(.dina(n1212), .dinb(n1187), .dout(n1213));
  jor  g0899(.dina(n1213), .dinb(n1172), .dout(G412));
  jxor g0900(.dina(n831), .dinb(n823), .dout(n1215));
  jxor g0901(.dina(n847), .dinb(n816), .dout(n1216));
  jxor g0902(.dina(n1216), .dinb(n855), .dout(n1217));
  jxor g0903(.dina(n793), .dinb(n787), .dout(n1218));
  jxor g0904(.dina(n807), .dinb(n801), .dout(n1219));
  jxor g0905(.dina(n1219), .dinb(n1218), .dout(n1220));
  jor  g0906(.dina(G4393), .dinb(n355), .dout(n1221));
  jnot g0907(.din(G58), .dout(n1222));
  jor  g0908(.dina(n1222), .dinb(G18), .dout(n1223));
  jand g0909(.dina(n1223), .dinb(n1221), .dout(n1224));
  jxor g0910(.dina(n1224), .dinb(n1220), .dout(n1225));
  jxor g0911(.dina(n1225), .dinb(n1217), .dout(n1226));
  jxor g0912(.dina(n1226), .dinb(n1215), .dout(n1227));
  jxor g0913(.dina(n389), .dinb(G3698), .dout(n1228));
  jor  g0914(.dina(n1228), .dinb(n355), .dout(n1229));
  jnot g0915(.din(G69), .dout(n1230));
  jand g0916(.dina(n935), .dinb(n1230), .dout(n1231));
  jand g0917(.dina(G70), .dinb(G69), .dout(n1232));
  jor  g0918(.dina(n1232), .dinb(G18), .dout(n1233));
  jor  g0919(.dina(n1233), .dinb(n1231), .dout(n1234));
  jand g0920(.dina(n1234), .dinb(n1229), .dout(n1235));
  jxor g0921(.dina(n1235), .dinb(n912), .dout(n1236));
  jnot g0922(.din(n1236), .dout(n1237));
  jxor g0923(.dina(n948), .dinb(n931), .dout(n1238));
  jnot g0924(.din(n920), .dout(n1239));
  jxor g0925(.dina(n882), .dinb(n873), .dout(n1240));
  jxor g0926(.dina(n902), .dinb(n895), .dout(n1241));
  jxor g0927(.dina(n1241), .dinb(n1240), .dout(n1242));
  jxor g0928(.dina(n1242), .dinb(n1239), .dout(n1243));
  jxor g0929(.dina(n1243), .dinb(n1238), .dout(n1244));
  jnot g0930(.din(n1244), .dout(n1245));
  jand g0931(.dina(n1245), .dinb(n1237), .dout(n1246));
  jand g0932(.dina(n1244), .dinb(n1236), .dout(n1247));
  jor  g0933(.dina(G1459), .dinb(n355), .dout(n1248));
  jnot g0934(.din(G114), .dout(n1249));
  jor  g0935(.dina(n1249), .dinb(G18), .dout(n1250));
  jand g0936(.dina(n1250), .dinb(n1248), .dout(n1251));
  jxor g0937(.dina(n1086), .dinb(n1081), .dout(n1252));
  jxor g0938(.dina(n1252), .dinb(n1251), .dout(n1253));
  jxor g0939(.dina(n1100), .dinb(n1073), .dout(n1254));
  jxor g0940(.dina(n1254), .dinb(n1066), .dout(n1255));
  jxor g0941(.dina(G1496), .dinb(G1492), .dout(n1256));
  jor  g0942(.dina(n1256), .dinb(n355), .dout(n1257));
  jxor g0943(.dina(G2204), .dinb(G1455), .dout(n1258));
  jor  g0944(.dina(n1258), .dinb(G18), .dout(n1259));
  jand g0945(.dina(n1259), .dinb(n1257), .dout(n1260));
  jxor g0946(.dina(n1260), .dinb(n1255), .dout(n1261));
  jxor g0947(.dina(n1261), .dinb(n1253), .dout(n1262));
  jxor g0948(.dina(n999), .dinb(n992), .dout(n1263));
  jxor g0949(.dina(n1019), .dinb(n1013), .dout(n1264));
  jxor g0950(.dina(n1264), .dinb(n1263), .dout(n1265));
  jxor g0951(.dina(n1265), .dinb(n727), .dout(n1266));
  jor  g0952(.dina(G2208), .dinb(n355), .dout(n1267));
  jnot g0953(.din(G82), .dout(n1268));
  jor  g0954(.dina(n1268), .dinb(G18), .dout(n1269));
  jand g0955(.dina(n1269), .dinb(n1267), .dout(n1270));
  jxor g0956(.dina(n758), .dinb(n748), .dout(n1271));
  jxor g0957(.dina(n1271), .dinb(n1270), .dout(n1272));
  jxor g0958(.dina(n741), .dinb(n734), .dout(n1273));
  jxor g0959(.dina(n1273), .dinb(n1272), .dout(n1274));
  jxor g0960(.dina(n1274), .dinb(n1266), .dout(n1275));
  jor  g0961(.dina(n1275), .dinb(n1262), .dout(n1276));
  jor  g0962(.dina(n1276), .dinb(n1247), .dout(n1277));
  jor  g0963(.dina(n1277), .dinb(n1246), .dout(n1278));
  jor  g0964(.dina(n1278), .dinb(n1227), .dout(G414));
  jnot g0965(.din(n1061), .dout(n1280));
  jnot g0966(.din(G170), .dout(n1281));
  jand g0967(.dina(n1281), .dinb(G18), .dout(n1282));
  jxor g0968(.dina(n1282), .dinb(n1068), .dout(n1283));
  jnot g0969(.din(n1283), .dout(n1284));
  jand g0970(.dina(n1284), .dinb(n1280), .dout(n1285));
  jand g0971(.dina(n1283), .dinb(n1061), .dout(n1286));
  jor  g0972(.dina(n1286), .dinb(n564), .dout(n1287));
  jor  g0973(.dina(n1287), .dinb(n1285), .dout(n1288));
  jnot g0974(.din(n1077), .dout(n1289));
  jor  g0975(.dina(n1095), .dinb(n1289), .dout(n1290));
  jnot g0976(.din(n1096), .dout(n1291));
  jor  g0977(.dina(n1291), .dinb(n1076), .dout(n1292));
  jand g0978(.dina(n1292), .dinb(n1290), .dout(n1293));
  jxor g0979(.dina(G165), .dinb(G164), .dout(n1294));
  jand g0980(.dina(n1294), .dinb(n1173), .dout(n1295));
  jxor g0981(.dina(n1295), .dinb(n1293), .dout(n1296));
  jxor g0982(.dina(n1296), .dinb(n1288), .dout(n1297));
  jxor g0983(.dina(n790), .dinb(n784), .dout(n1298));
  jxor g0984(.dina(n804), .dinb(n797), .dout(n1299));
  jxor g0985(.dina(n1299), .dinb(n1298), .dout(n1300));
  jxor g0986(.dina(n1300), .dinb(n851), .dout(n1301));
  jand g0987(.dina(G197), .dinb(G18), .dout(n1302));
  jor  g0988(.dina(n1302), .dinb(n1205), .dout(n1303));
  jnot g0989(.din(n1303), .dout(n1304));
  jxor g0990(.dina(n827), .dinb(n819), .dout(n1305));
  jxor g0991(.dina(n1305), .dinb(n1304), .dout(n1306));
  jnot g0992(.din(n1306), .dout(n1307));
  jxor g0993(.dina(n843), .dinb(n812), .dout(n1308));
  jxor g0994(.dina(n1308), .dinb(n1307), .dout(n1309));
  jand g0995(.dina(n1309), .dinb(n1301), .dout(n1310));
  jor  g0996(.dina(n1310), .dinb(n1297), .dout(n1311));
  jand g0997(.dina(G208), .dinb(G18), .dout(n1312));
  jor  g0998(.dina(n1312), .dinb(n1189), .dout(n1313));
  jxor g0999(.dina(n878), .dinb(n869), .dout(n1314));
  jxor g1000(.dina(n899), .dinb(n891), .dout(n1315));
  jxor g1001(.dina(n1315), .dinb(n1314), .dout(n1316));
  jxor g1002(.dina(n1316), .dinb(n1313), .dout(n1317));
  jnot g1003(.din(n916), .dout(n1318));
  jxor g1004(.dina(n945), .dinb(n927), .dout(n1319));
  jxor g1005(.dina(n1319), .dinb(n1318), .dout(n1320));
  jnot g1006(.din(G198), .dout(n1321));
  jor  g1007(.dina(n1321), .dinb(n355), .dout(n1322));
  jand g1008(.dina(n1322), .dinb(n353), .dout(n1323));
  jxor g1009(.dina(n1323), .dinb(n908), .dout(n1324));
  jxor g1010(.dina(n1324), .dinb(n1320), .dout(n1325));
  jand g1011(.dina(n1325), .dinb(n1317), .dout(n1326));
  jnot g1012(.din(n1301), .dout(n1327));
  jnot g1013(.din(n1309), .dout(n1328));
  jand g1014(.dina(n1328), .dinb(n1327), .dout(n1329));
  jnot g1015(.din(n1317), .dout(n1330));
  jnot g1016(.din(n1325), .dout(n1331));
  jand g1017(.dina(n1331), .dinb(n1330), .dout(n1332));
  jor  g1018(.dina(n1332), .dinb(n1329), .dout(n1333));
  jor  g1019(.dina(n1333), .dinb(n1326), .dout(n1334));
  jor  g1020(.dina(n1334), .dinb(n1311), .dout(n1335));
  jxor g1021(.dina(n744), .dinb(n730), .dout(n1336));
  jxor g1022(.dina(n1336), .dinb(n737), .dout(n1337));
  jxor g1023(.dina(n754), .dinb(n723), .dout(n1338));
  jnot g1024(.din(n994), .dout(n1339));
  jand g1025(.dina(n1016), .dinb(n1339), .dout(n1340));
  jnot g1026(.din(n1015), .dout(n1341));
  jand g1027(.dina(n1341), .dinb(n995), .dout(n1342));
  jor  g1028(.dina(n1342), .dinb(n1340), .dout(n1343));
  jnot g1029(.din(n987), .dout(n1344));
  jand g1030(.dina(n1009), .dinb(n1344), .dout(n1345));
  jnot g1031(.din(n1008), .dout(n1346));
  jand g1032(.dina(n1346), .dinb(n988), .dout(n1347));
  jor  g1033(.dina(n1347), .dinb(n1345), .dout(n1348));
  jxor g1034(.dina(n1348), .dinb(n1343), .dout(n1349));
  jnot g1035(.din(G181), .dout(n1350));
  jor  g1036(.dina(n1350), .dinb(n355), .dout(n1351));
  jand g1037(.dina(n1351), .dinb(n1166), .dout(n1352));
  jxor g1038(.dina(n1352), .dinb(n1349), .dout(n1353));
  jxor g1039(.dina(n1353), .dinb(n1338), .dout(n1354));
  jxor g1040(.dina(n1354), .dinb(n1337), .dout(n1355));
  jor  g1041(.dina(n1355), .dinb(n1335), .dout(G416));
  jnot g1042(.din(n372), .dout(n1357));
  jxor g1043(.dina(n377), .dinb(G3717), .dout(n1358));
  jand g1044(.dina(n1358), .dinb(n1357), .dout(n1359));
  jnot g1045(.din(n387), .dout(n1360));
  jxor g1046(.dina(n401), .dinb(G3705), .dout(n1361));
  jand g1047(.dina(n1361), .dinb(n362), .dout(n1362));
  jand g1048(.dina(n1362), .dinb(G4526), .dout(n1363));
  jand g1049(.dina(n1363), .dinb(n1360), .dout(n1364));
  jand g1050(.dina(n1364), .dinb(n1359), .dout(n1365));
  jnot g1051(.din(n407), .dout(n1366));
  jand g1052(.dina(n1361), .dinb(n390), .dout(n1367));
  jand g1053(.dina(n1367), .dinb(n1360), .dout(n1368));
  jor  g1054(.dina(n1368), .dinb(n1366), .dout(n1369));
  jand g1055(.dina(n1369), .dinb(n1359), .dout(n1370));
  jnot g1056(.din(n413), .dout(n1371));
  jand g1057(.dina(n1371), .dinb(n1359), .dout(n1372));
  jnot g1058(.din(n419), .dout(n1373));
  jor  g1059(.dina(n1373), .dinb(n1372), .dout(n1374));
  jor  g1060(.dina(n1374), .dinb(n1370), .dout(n1375));
  jor  g1061(.dina(n1375), .dinb(n1365), .dout(n1376));
  jnot g1062(.din(n452), .dout(n1377));
  jand g1063(.dina(n1377), .dinb(n1376), .dout(n1378));
  jnot g1064(.din(n464), .dout(n1379));
  jor  g1065(.dina(n1379), .dinb(n1378), .dout(n1380));
  jand g1066(.dina(n494), .dinb(n1380), .dout(n1381));
  jnot g1067(.din(n518), .dout(n1382));
  jor  g1068(.dina(n1382), .dinb(n1381), .dout(n1383));
  jand g1069(.dina(n542), .dinb(n1383), .dout(n1384));
  jor  g1070(.dina(n560), .dinb(n1384), .dout(n1385));
  jxor g1071(.dina(n578), .dinb(n1385), .dout(G295));
  jand g1072(.dina(n592), .dinb(n1385), .dout(n1387));
  jnot g1073(.din(n617), .dout(n1388));
  jor  g1074(.dina(n1388), .dinb(n1387), .dout(n1389));
  jand g1075(.dina(n637), .dinb(n1389), .dout(n1390));
  jnot g1076(.din(n656), .dout(n1391));
  jor  g1077(.dina(n1391), .dinb(n1390), .dout(n1392));
  jxor g1078(.dina(n678), .dinb(n1392), .dout(G324));
  jor  g1079(.dina(n1033), .dinb(n957), .dout(n1394));
  jand g1080(.dina(n1394), .dinb(n905), .dout(n1395));
  jor  g1081(.dina(n1395), .dinb(n1044), .dout(n1396));
  jand g1082(.dina(n1396), .dinb(n864), .dout(n1397));
  jor  g1083(.dina(n1397), .dinb(n981), .dout(n1398));
  jand g1084(.dina(n1398), .dinb(n810), .dout(n1399));
  jor  g1085(.dina(n1399), .dinb(n972), .dout(G252));
  jnot g1086(.din(n568), .dout(n1401));
  jnot g1087(.din(n584), .dout(n1402));
  jnot g1088(.din(n589), .dout(n1403));
  jnot g1089(.din(n579), .dout(n1404));
  jor  g1090(.dina(n1404), .dinb(n562), .dout(n1405));
  jor  g1091(.dina(n1405), .dinb(n1403), .dout(n1406));
  jor  g1092(.dina(n1406), .dinb(n1402), .dout(n1407));
  jand g1093(.dina(n1407), .dinb(n615), .dout(n1408));
  jxor g1094(.dina(n1408), .dinb(n1401), .dout(G310));
  jand g1095(.dina(n1406), .dinb(n613), .dout(n1410));
  jxor g1096(.dina(n1410), .dinb(n1402), .dout(G313));
  jnot g1097(.din(n608), .dout(n1412));
  jnot g1098(.din(n607), .dout(n1413));
  jand g1099(.dina(n1413), .dinb(n1412), .dout(n1414));
  jand g1100(.dina(n1414), .dinb(n1405), .dout(n1415));
  jxor g1101(.dina(n1415), .dinb(n1403), .dout(G316));
  jand g1102(.dina(n578), .dinb(n1385), .dout(n1417));
  jor  g1103(.dina(n1417), .dinb(n606), .dout(n1418));
  jxor g1104(.dina(n1418), .dinb(n573), .dout(G319));
  jnot g1105(.din(n661), .dout(n1420));
  jnot g1106(.din(n665), .dout(n1421));
  jnot g1107(.din(n669), .dout(n1422));
  jnot g1108(.din(n679), .dout(n1423));
  jor  g1109(.dina(n1423), .dinb(n657), .dout(n1424));
  jor  g1110(.dina(n1424), .dinb(n1422), .dout(n1425));
  jor  g1111(.dina(n1425), .dinb(n1421), .dout(n1426));
  jand g1112(.dina(n1426), .dinb(n704), .dout(n1427));
  jxor g1113(.dina(n1427), .dinb(n1420), .dout(G327));
  jnot g1114(.din(n701), .dout(n1429));
  jand g1115(.dina(n1425), .dinb(n1429), .dout(n1430));
  jxor g1116(.dina(n1430), .dinb(n1421), .dout(G330));
  jnot g1117(.din(n699), .dout(n1432));
  jand g1118(.dina(n1424), .dinb(n1432), .dout(n1433));
  jxor g1119(.dina(n1433), .dinb(n1422), .dout(G333));
  jand g1120(.dina(n678), .dinb(n1392), .dout(n1435));
  jor  g1121(.dina(n1435), .dinb(n697), .dout(n1436));
  jxor g1122(.dina(n1436), .dinb(n674), .dout(G336));
  jor  g1123(.dina(G408), .dinb(G404), .dout(n1438));
  jor  g1124(.dina(G410), .dinb(G406), .dout(n1439));
  jor  g1125(.dina(n1439), .dinb(n1438), .dout(n1440));
  jor  g1126(.dina(n1440), .dinb(G412), .dout(n1441));
  jor  g1127(.dina(n1441), .dinb(G416), .dout(n1442));
  jor  g1128(.dina(n1442), .dinb(G414), .dout(G418));
  jnot g1129(.din(n631), .dout(n1444));
  jnot g1130(.din(n627), .dout(n1445));
  jor  g1131(.dina(n1445), .dinb(n618), .dout(n1446));
  jand g1132(.dina(n1446), .dinb(n648), .dout(n1447));
  jor  g1133(.dina(n1447), .dinb(n653), .dout(n1448));
  jand g1134(.dina(n1448), .dinb(n643), .dout(n1449));
  jxor g1135(.dina(n1449), .dinb(n1444), .dout(G298));
  jnot g1136(.din(n635), .dout(n1451));
  jxor g1137(.dina(n1447), .dinb(n1451), .dout(G301));
  jand g1138(.dina(n1156), .dinb(G2239), .dout(n1453));
  jnot g1139(.din(n1453), .dout(n1454));
  jand g1140(.dina(n1454), .dinb(n1389), .dout(n1455));
  jor  g1141(.dina(n1455), .dinb(n645), .dout(n1456));
  jxor g1142(.dina(n1456), .dinb(n622), .dout(G304));
  jxor g1143(.dina(n626), .dinb(n1389), .dout(G307));
  jxor g1144(.dina(n480), .dinb(n1380), .dout(G344));
  jnot g1145(.din(n714), .dout(n1460));
  jnot g1146(.din(n365), .dout(n1461));
  jor  g1147(.dina(n711), .dinb(n710), .dout(n1462));
  jxor g1148(.dina(n1462), .dinb(n1461), .dout(n1463));
  jnot g1149(.din(n1463), .dout(n1464));
  jor  g1150(.dina(n1464), .dinb(n1460), .dout(n1465));
  jand g1151(.dina(n1465), .dinb(n715), .dout(G422));
  jxor g1152(.dina(n713), .dinb(n709), .dout(G419));
  jnot g1153(.din(n470), .dout(n1468));
  jnot g1154(.din(n486), .dout(n1469));
  jnot g1155(.din(n491), .dout(n1470));
  jnot g1156(.din(n481), .dout(n1471));
  jor  g1157(.dina(n1471), .dinb(n465), .dout(n1472));
  jor  g1158(.dina(n1472), .dinb(n1470), .dout(n1473));
  jor  g1159(.dina(n1473), .dinb(n1469), .dout(n1474));
  jand g1160(.dina(n1474), .dinb(n516), .dout(n1475));
  jxor g1161(.dina(n1475), .dinb(n1468), .dout(G359));
  jand g1162(.dina(n1473), .dinb(n514), .dout(n1477));
  jxor g1163(.dina(n1477), .dinb(n1469), .dout(G362));
  jand g1164(.dina(n508), .dinb(n510), .dout(n1479));
  jand g1165(.dina(n1479), .dinb(n1472), .dout(n1480));
  jxor g1166(.dina(n1480), .dinb(n1470), .dout(G365));
  jnot g1167(.din(n507), .dout(n1482));
  jand g1168(.dina(n480), .dinb(n1380), .dout(n1483));
  jor  g1169(.dina(n1483), .dinb(n1482), .dout(n1484));
  jxor g1170(.dina(n1484), .dinb(n475), .dout(G368));
  jand g1171(.dina(n530), .dinb(n1383), .dout(n1486));
  jand g1172(.dina(n1486), .dinb(n552), .dout(n1487));
  jor  g1173(.dina(n1487), .dinb(n558), .dout(n1488));
  jxor g1174(.dina(n1488), .dinb(n535), .dout(G347));
  jor  g1175(.dina(n1486), .dinb(n556), .dout(n1490));
  jxor g1176(.dina(n1490), .dinb(n540), .dout(G350));
  jnot g1177(.din(n528), .dout(n1492));
  jand g1178(.dina(n1492), .dinb(G4420), .dout(n1493));
  jnot g1179(.din(n1493), .dout(n1494));
  jand g1180(.dina(n1494), .dinb(n1383), .dout(n1495));
  jor  g1181(.dina(n1495), .dinb(n554), .dout(n1496));
  jxor g1182(.dina(n1496), .dinb(n524), .dout(G353));
  jxor g1183(.dina(n529), .dinb(n1383), .dout(G356));
  jxor g1184(.dina(n589), .dinb(n584), .dout(n1499));
  jxor g1185(.dina(n1499), .dinb(n635), .dout(n1500));
  jnot g1186(.din(n622), .dout(n1501));
  jnot g1187(.din(n653), .dout(n1502));
  jand g1188(.dina(n647), .dinb(n1502), .dout(n1503));
  jor  g1189(.dina(n1503), .dinb(n649), .dout(n1504));
  jxor g1190(.dina(n1504), .dinb(n1444), .dout(n1505));
  jxor g1191(.dina(n1505), .dinb(n1501), .dout(n1506));
  jxor g1192(.dina(n1506), .dinb(n1454), .dout(n1507));
  jand g1193(.dina(n1507), .dinb(n618), .dout(n1508));
  jxor g1194(.dina(n645), .dinb(n1501), .dout(n1509));
  jand g1195(.dina(n648), .dinb(n1445), .dout(n1510));
  jnot g1196(.din(n1510), .dout(n1511));
  jor  g1197(.dina(n1511), .dinb(n642), .dout(n1512));
  jor  g1198(.dina(n1510), .dinb(n653), .dout(n1513));
  jand g1199(.dina(n1513), .dinb(n1512), .dout(n1514));
  jxor g1200(.dina(n1514), .dinb(n1444), .dout(n1515));
  jxor g1201(.dina(n1515), .dinb(n1509), .dout(n1516));
  jand g1202(.dina(n1516), .dinb(n1389), .dout(n1517));
  jor  g1203(.dina(n1517), .dinb(n1508), .dout(n1518));
  jand g1204(.dina(n613), .dinb(n606), .dout(n1519));
  jnot g1205(.din(n606), .dout(n1520));
  jand g1206(.dina(n605), .dinb(n1520), .dout(n1521));
  jand g1207(.dina(n1521), .dinb(n610), .dout(n1522));
  jxor g1208(.dina(n1522), .dinb(n578), .dout(n1523));
  jor  g1209(.dina(n1523), .dinb(n1519), .dout(n1524));
  jor  g1210(.dina(n572), .dinb(n569), .dout(n1525));
  jand g1211(.dina(n1520), .dinb(n1525), .dout(n1526));
  jor  g1212(.dina(n1526), .dinb(n608), .dout(n1527));
  jxor g1213(.dina(n1527), .dinb(n615), .dout(n1528));
  jxor g1214(.dina(n1528), .dinb(n1401), .dout(n1529));
  jxor g1215(.dina(n1529), .dinb(n1524), .dout(n1530));
  jor  g1216(.dina(n1530), .dinb(n1385), .dout(n1531));
  jand g1217(.dina(n1414), .dinb(n1404), .dout(n1532));
  jxor g1218(.dina(n1532), .dinb(n568), .dout(n1533));
  jxor g1219(.dina(n606), .dinb(n573), .dout(n1534));
  jand g1220(.dina(n589), .dinb(n579), .dout(n1535));
  jor  g1221(.dina(n1535), .dinb(n612), .dout(n1536));
  jnot g1222(.din(n1536), .dout(n1537));
  jand g1223(.dina(n1537), .dinb(n599), .dout(n1538));
  jnot g1224(.din(n591), .dout(n1539));
  jand g1225(.dina(n1536), .dinb(n1539), .dout(n1540));
  jand g1226(.dina(n1540), .dinb(n615), .dout(n1541));
  jor  g1227(.dina(n1541), .dinb(n1538), .dout(n1542));
  jxor g1228(.dina(n1542), .dinb(n1534), .dout(n1543));
  jxor g1229(.dina(n1543), .dinb(n1533), .dout(n1544));
  jor  g1230(.dina(n1544), .dinb(n562), .dout(n1545));
  jand g1231(.dina(n1545), .dinb(n1531), .dout(n1546));
  jxor g1232(.dina(n1546), .dinb(n1518), .dout(n1547));
  jxor g1233(.dina(n1547), .dinb(n1500), .dout(G321));
  jand g1234(.dina(n713), .dinb(n709), .dout(n1549));
  jor  g1235(.dina(n1549), .dinb(n1463), .dout(n1550));
  jnot g1236(.din(n683), .dout(n1551));
  jand g1237(.dina(n707), .dinb(n1392), .dout(n1552));
  jand g1238(.dina(n712), .dinb(n708), .dout(n1553));
  jor  g1239(.dina(n1553), .dinb(n1464), .dout(n1554));
  jor  g1240(.dina(n1554), .dinb(n1552), .dout(n1555));
  jor  g1241(.dina(n1555), .dinb(n1551), .dout(n1556));
  jand g1242(.dina(n1556), .dinb(n1550), .dout(n1557));
  jand g1243(.dina(n1463), .dinb(n707), .dout(n1558));
  jand g1244(.dina(n1558), .dinb(n657), .dout(n1559));
  jor  g1245(.dina(n1559), .dinb(n1557), .dout(n1560));
  jxor g1246(.dina(n669), .dinb(n665), .dout(n1561));
  jor  g1247(.dina(n701), .dinb(n686), .dout(n1562));
  jand g1248(.dina(n1562), .dinb(n703), .dout(n1563));
  jxor g1249(.dina(n1563), .dinb(n1420), .dout(n1564));
  jor  g1250(.dina(n677), .dinb(n675), .dout(n1565));
  jxor g1251(.dina(n1565), .dinb(n674), .dout(n1566));
  jxor g1252(.dina(n1566), .dinb(n699), .dout(n1567));
  jxor g1253(.dina(n1567), .dinb(n1564), .dout(n1568));
  jand g1254(.dina(n1568), .dinb(n657), .dout(n1569));
  jand g1255(.dina(n679), .dinb(n692), .dout(n1570));
  jor  g1256(.dina(n1570), .dinb(n701), .dout(n1571));
  jor  g1257(.dina(n1571), .dinb(n687), .dout(n1572));
  jnot g1258(.din(n1571), .dout(n1573));
  jor  g1259(.dina(n1573), .dinb(n680), .dout(n1574));
  jor  g1260(.dina(n1574), .dinb(n705), .dout(n1575));
  jand g1261(.dina(n1575), .dinb(n1572), .dout(n1576));
  jor  g1262(.dina(n699), .dinb(n679), .dout(n1577));
  jxor g1263(.dina(n1577), .dinb(n1420), .dout(n1578));
  jxor g1264(.dina(n1578), .dinb(n1576), .dout(n1579));
  jxor g1265(.dina(n1579), .dinb(n697), .dout(n1580));
  jxor g1266(.dina(n1580), .dinb(n674), .dout(n1581));
  jand g1267(.dina(n1581), .dinb(n1392), .dout(n1582));
  jor  g1268(.dina(n1582), .dinb(n1569), .dout(n1583));
  jxor g1269(.dina(n1583), .dinb(n1561), .dout(n1584));
  jxor g1270(.dina(n1584), .dinb(n1560), .dout(G338));
  jxor g1271(.dina(n491), .dinb(n486), .dout(n1586));
  jxor g1272(.dina(n1586), .dinb(n540), .dout(n1587));
  jnot g1273(.din(n535), .dout(n1588));
  jnot g1274(.din(n557), .dout(n1589));
  jor  g1275(.dina(n556), .dinb(n549), .dout(n1590));
  jand g1276(.dina(n1590), .dinb(n1589), .dout(n1591));
  jxor g1277(.dina(n1591), .dinb(n1588), .dout(n1592));
  jxor g1278(.dina(n1494), .dinb(n524), .dout(n1593));
  jxor g1279(.dina(n1593), .dinb(n1592), .dout(n1594));
  jand g1280(.dina(n1594), .dinb(n519), .dout(n1595));
  jxor g1281(.dina(n554), .dinb(n524), .dout(n1596));
  jxor g1282(.dina(n1596), .dinb(n535), .dout(n1597));
  jand g1283(.dina(n1494), .dinb(n524), .dout(n1598));
  jor  g1284(.dina(n1598), .dinb(n553), .dout(n1599));
  jnot g1285(.din(n1599), .dout(n1600));
  jand g1286(.dina(n1600), .dinb(n558), .dout(n1601));
  jand g1287(.dina(n1599), .dinb(n551), .dout(n1602));
  jor  g1288(.dina(n1602), .dinb(n1601), .dout(n1603));
  jxor g1289(.dina(n1603), .dinb(n1597), .dout(n1604));
  jand g1290(.dina(n1604), .dinb(n1383), .dout(n1605));
  jor  g1291(.dina(n1605), .dinb(n1595), .dout(n1606));
  jor  g1292(.dina(n474), .dinb(n471), .dout(n1607));
  jand g1293(.dina(n507), .dinb(n1607), .dout(n1608));
  jor  g1294(.dina(n1608), .dinb(n509), .dout(n1609));
  jnot g1295(.din(n516), .dout(n1610));
  jnot g1296(.din(n514), .dout(n1611));
  jor  g1297(.dina(n1611), .dinb(n507), .dout(n1612));
  jor  g1298(.dina(n505), .dinb(n1482), .dout(n1613));
  jor  g1299(.dina(n1613), .dinb(n512), .dout(n1614));
  jxor g1300(.dina(n1614), .dinb(n480), .dout(n1615));
  jand g1301(.dina(n1615), .dinb(n1612), .dout(n1616));
  jxor g1302(.dina(n1616), .dinb(n1468), .dout(n1617));
  jxor g1303(.dina(n1617), .dinb(n1610), .dout(n1618));
  jxor g1304(.dina(n1618), .dinb(n1609), .dout(n1619));
  jor  g1305(.dina(n1619), .dinb(n1380), .dout(n1620));
  jand g1306(.dina(n1479), .dinb(n1471), .dout(n1621));
  jxor g1307(.dina(n1621), .dinb(n470), .dout(n1622));
  jxor g1308(.dina(n507), .dinb(n475), .dout(n1623));
  jand g1309(.dina(n491), .dinb(n481), .dout(n1624));
  jor  g1310(.dina(n1624), .dinb(n1611), .dout(n1625));
  jor  g1311(.dina(n1625), .dinb(n502), .dout(n1626));
  jnot g1312(.din(n1625), .dout(n1627));
  jor  g1313(.dina(n1627), .dinb(n493), .dout(n1628));
  jor  g1314(.dina(n1628), .dinb(n1610), .dout(n1629));
  jand g1315(.dina(n1629), .dinb(n1626), .dout(n1630));
  jxor g1316(.dina(n1630), .dinb(n1623), .dout(n1631));
  jxor g1317(.dina(n1631), .dinb(n1622), .dout(n1632));
  jor  g1318(.dina(n1632), .dinb(n465), .dout(n1633));
  jand g1319(.dina(n1633), .dinb(n1620), .dout(n1634));
  jxor g1320(.dina(n1634), .dinb(n1606), .dout(n1635));
  jxor g1321(.dina(n1635), .dinb(n1587), .dout(G370));
  jxor g1322(.dina(n450), .dinb(n1360), .dout(n1637));
  jnot g1323(.din(n455), .dout(n1638));
  jnot g1324(.din(n460), .dout(n1639));
  jor  g1325(.dina(n1639), .dinb(n1638), .dout(n1640));
  jand g1326(.dina(n1640), .dinb(n461), .dout(n1641));
  jxor g1327(.dina(n1641), .dinb(n446), .dout(n1642));
  jnot g1328(.din(n1642), .dout(n1643));
  jxor g1329(.dina(n1148), .dinb(n429), .dout(n1644));
  jnot g1330(.din(n1644), .dout(n1645));
  jor  g1331(.dina(n1645), .dinb(n1643), .dout(n1646));
  jor  g1332(.dina(n1644), .dinb(n1642), .dout(n1647));
  jand g1333(.dina(n1647), .dinb(n422), .dout(n1648));
  jand g1334(.dina(n1648), .dinb(n1646), .dout(n1649));
  jxor g1335(.dina(n458), .dinb(n429), .dout(n1650));
  jxor g1336(.dina(n1650), .dinb(n446), .dout(n1651));
  jnot g1337(.din(n462), .dout(n1652));
  jor  g1338(.dina(n1148), .dinb(n429), .dout(n1653));
  jand g1339(.dina(n1653), .dinb(n457), .dout(n1654));
  jand g1340(.dina(n1654), .dinb(n1652), .dout(n1655));
  jnot g1341(.din(n1655), .dout(n1656));
  jnot g1342(.din(n456), .dout(n1657));
  jor  g1343(.dina(n1654), .dinb(n1657), .dout(n1658));
  jand g1344(.dina(n1658), .dinb(n1656), .dout(n1659));
  jor  g1345(.dina(n1659), .dinb(n1651), .dout(n1660));
  jnot g1346(.din(n1651), .dout(n1661));
  jnot g1347(.din(n1659), .dout(n1662));
  jor  g1348(.dina(n1662), .dinb(n1661), .dout(n1663));
  jand g1349(.dina(n1663), .dinb(n1376), .dout(n1664));
  jand g1350(.dina(n1664), .dinb(n1660), .dout(n1665));
  jor  g1351(.dina(n1665), .dinb(n1649), .dout(n1666));
  jand g1352(.dina(n1136), .dinb(n403), .dout(n1667));
  jnot g1353(.din(n1667), .dout(n1668));
  jor  g1354(.dina(n1668), .dinb(n1128), .dout(n1669));
  jnot g1355(.din(n1128), .dout(n1670));
  jand g1356(.dina(n1362), .dinb(n1360), .dout(n1671));
  jor  g1357(.dina(n1671), .dinb(n1670), .dout(n1672));
  jor  g1358(.dina(n1672), .dinb(n1667), .dout(n1673));
  jand g1359(.dina(n1673), .dinb(n1669), .dout(n1674));
  jxor g1360(.dina(n1674), .dinb(n372), .dout(n1675));
  jnot g1361(.din(n1672), .dout(n1676));
  jor  g1362(.dina(n1676), .dinb(n1127), .dout(n1677));
  jand g1363(.dina(n1677), .dinb(n417), .dout(n1678));
  jxor g1364(.dina(n1678), .dinb(n402), .dout(n1679));
  jxor g1365(.dina(n1679), .dinb(n354), .dout(n1680));
  jnot g1366(.din(n1680), .dout(n1681));
  jand g1367(.dina(n1681), .dinb(n1675), .dout(n1682));
  jnot g1368(.din(n1675), .dout(n1683));
  jand g1369(.dina(n1680), .dinb(n1683), .dout(n1684));
  jor  g1370(.dina(n1684), .dinb(n388), .dout(n1685));
  jor  g1371(.dina(n1685), .dinb(n1682), .dout(n1686));
  jxor g1372(.dina(n1130), .dinb(n372), .dout(n1687));
  jand g1373(.dina(n407), .dinb(n354), .dout(n1688));
  jand g1374(.dina(n1688), .dinb(n413), .dout(n1689));
  jand g1375(.dina(n1689), .dinb(n395), .dout(n1690));
  jnot g1376(.din(n1689), .dout(n1691));
  jand g1377(.dina(n1670), .dinb(n390), .dout(n1692));
  jor  g1378(.dina(n1692), .dinb(n362), .dout(n1693));
  jand g1379(.dina(n1693), .dinb(n1691), .dout(n1694));
  jor  g1380(.dina(n1694), .dinb(n1690), .dout(n1695));
  jand g1381(.dina(n401), .dinb(G3705), .dout(n1696));
  jor  g1382(.dina(n1696), .dinb(n390), .dout(n1697));
  jand g1383(.dina(n1697), .dinb(n412), .dout(n1698));
  jxor g1384(.dina(n1698), .dinb(n1695), .dout(n1699));
  jnot g1385(.din(n1699), .dout(n1700));
  jand g1386(.dina(n1700), .dinb(n1687), .dout(n1701));
  jnot g1387(.din(n1687), .dout(n1702));
  jand g1388(.dina(n1699), .dinb(n1702), .dout(n1703));
  jor  g1389(.dina(n1703), .dinb(G4526), .dout(n1704));
  jor  g1390(.dina(n1704), .dinb(n1701), .dout(n1705));
  jand g1391(.dina(n1705), .dinb(n1686), .dout(n1706));
  jxor g1392(.dina(n1706), .dinb(n379), .dout(n1707));
  jxor g1393(.dina(n1707), .dinb(n1666), .dout(n1708));
  jxor g1394(.dina(n1708), .dinb(n1637), .dout(G399));
  jdff  g1395(.din(G1), .dout(G2));
  jdff  g1396(.din(G1), .dout(G3));
  jdff  g1397(.din(G1459), .dout(G450));
  jdff  g1398(.din(G1469), .dout(G448));
  jdff  g1399(.din(G1480), .dout(G444));
  jdff  g1400(.din(G1486), .dout(G442));
  jdff  g1401(.din(G1492), .dout(G440));
  jdff  g1402(.din(G1496), .dout(G438));
  jdff  g1403(.din(G2208), .dout(G496));
  jdff  g1404(.din(G2218), .dout(G494));
  jdff  g1405(.din(G2224), .dout(G492));
  jdff  g1406(.din(G2230), .dout(G490));
  jdff  g1407(.din(G2236), .dout(G488));
  jdff  g1408(.din(G2239), .dout(G486));
  jdff  g1409(.din(G2247), .dout(G484));
  jdff  g1410(.din(G2253), .dout(G482));
  jdff  g1411(.din(G2256), .dout(G480));
  jdff  g1412(.din(G3698), .dout(G560));
  jdff  g1413(.din(G3701), .dout(G542));
  jdff  g1414(.din(G3705), .dout(G558));
  jdff  g1415(.din(G3711), .dout(G556));
  jdff  g1416(.din(G3717), .dout(G554));
  jdff  g1417(.din(G3723), .dout(G552));
  jdff  g1418(.din(G3729), .dout(G550));
  jdff  g1419(.din(G3737), .dout(G548));
  jdff  g1420(.din(G3743), .dout(G546));
  jdff  g1421(.din(G3749), .dout(G544));
  jdff  g1422(.din(G4393), .dout(G540));
  jdff  g1423(.din(G4400), .dout(G538));
  jdff  g1424(.din(G4405), .dout(G536));
  jdff  g1425(.din(G4410), .dout(G534));
  jdff  g1426(.din(G4415), .dout(G532));
  jdff  g1427(.din(G4420), .dout(G530));
  jdff  g1428(.din(G4427), .dout(G528));
  jdff  g1429(.din(G4432), .dout(G526));
  jdff  g1430(.din(G4437), .dout(G524));
  jdff  g1431(.din(G1462), .dout(G436));
  jdff  g1432(.din(G2211), .dout(G478));
  jdff  g1433(.din(G4394), .dout(G522));
  jdff  g1434(.din(G1), .dout(G432));
  jdff  g1435(.din(G106), .dout(G446));
  jnot g1436(.din(G15), .dout(G286));
  jor  g1437(.dina(n345), .dinb(G5), .dout(G289));
  jnot g1438(.din(G15), .dout(G341));
  jor  g1439(.dina(n349), .dinb(G5), .dout(G281));
  jdff  g1440(.din(G1), .dout(G453));
  jand g1441(.dina(n1125), .dinb(n1122), .dout(G264));
  jor  g1442(.dina(n720), .dinb(n716), .dout(G270));
  jand g1443(.dina(n1125), .dinb(n1122), .dout(G249));
  jor  g1444(.dina(n720), .dinb(n716), .dout(G276));
  jor  g1445(.dina(n720), .dinb(n716), .dout(G273));
  jand g1446(.dina(n1465), .dinb(n715), .dout(G469));
  jxor g1447(.dina(n713), .dinb(n709), .dout(G471));
endmodule


