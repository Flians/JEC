/*

c432:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 1154
	jand: 104
	jor: 104

Summary:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 1154
	jand: 104
	jor: 104
*/

module c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G4gat_0;
	wire[2:0] w_G8gat_0;
	wire[2:0] w_G11gat_0;
	wire[2:0] w_G14gat_0;
	wire[2:0] w_G17gat_0;
	wire[2:0] w_G21gat_0;
	wire[2:0] w_G24gat_0;
	wire[1:0] w_G27gat_0;
	wire[2:0] w_G30gat_0;
	wire[2:0] w_G34gat_0;
	wire[1:0] w_G40gat_0;
	wire[1:0] w_G43gat_0;
	wire[2:0] w_G47gat_0;
	wire[1:0] w_G50gat_0;
	wire[1:0] w_G53gat_0;
	wire[2:0] w_G56gat_0;
	wire[1:0] w_G56gat_1;
	wire[1:0] w_G60gat_0;
	wire[2:0] w_G63gat_0;
	wire[2:0] w_G66gat_0;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G73gat_0;
	wire[2:0] w_G76gat_0;
	wire[1:0] w_G79gat_0;
	wire[2:0] w_G82gat_0;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G89gat_0;
	wire[2:0] w_G92gat_0;
	wire[2:0] w_G95gat_0;
	wire[2:0] w_G99gat_0;
	wire[1:0] w_G102gat_0;
	wire[1:0] w_G105gat_0;
	wire[2:0] w_G108gat_0;
	wire[2:0] w_G112gat_0;
	wire[1:0] w_G115gat_0;
	wire[2:0] w_G223gat_0;
	wire[2:0] w_G223gat_1;
	wire[2:0] w_G223gat_2;
	wire[2:0] w_G223gat_3;
	wire w_G223gat_4;
	wire G223gat_fa_;
	wire[2:0] w_G329gat_0;
	wire[2:0] w_G329gat_1;
	wire[2:0] w_G329gat_2;
	wire[2:0] w_G329gat_3;
	wire w_G329gat_4;
	wire G329gat_fa_;
	wire[2:0] w_G370gat_0;
	wire[1:0] w_G370gat_1;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire[1:0] w_n43_0;
	wire[1:0] w_n44_0;
	wire[1:0] w_n45_0;
	wire[2:0] w_n46_0;
	wire[1:0] w_n47_0;
	wire[1:0] w_n49_0;
	wire[1:0] w_n51_0;
	wire[1:0] w_n54_0;
	wire[1:0] w_n57_0;
	wire[1:0] w_n60_0;
	wire[1:0] w_n62_0;
	wire[1:0] w_n64_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n73_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n78_0;
	wire[1:0] w_n80_0;
	wire[1:0] w_n81_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n88_0;
	wire[2:0] w_n93_0;
	wire[2:0] w_n93_1;
	wire[2:0] w_n93_2;
	wire[2:0] w_n93_3;
	wire[1:0] w_n95_0;
	wire[1:0] w_n102_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n106_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n111_0;
	wire[1:0] w_n113_0;
	wire[1:0] w_n117_0;
	wire[2:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n123_0;
	wire[1:0] w_n125_0;
	wire[1:0] w_n127_0;
	wire[2:0] w_n131_0;
	wire[1:0] w_n138_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n141_0;
	wire[1:0] w_n144_0;
	wire[1:0] w_n145_0;
	wire[1:0] w_n147_0;
	wire[1:0] w_n149_0;
	wire[1:0] w_n151_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n159_0;
	wire[1:0] w_n164_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n173_0;
	wire[2:0] w_n181_0;
	wire[2:0] w_n181_1;
	wire[2:0] w_n181_2;
	wire[1:0] w_n183_0;
	wire[1:0] w_n185_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n202_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n209_0;
	wire[1:0] w_n211_0;
	wire[1:0] w_n222_0;
	wire[1:0] w_n227_0;
	wire[1:0] w_n230_0;
	wire[2:0] w_n246_0;
	wire[2:0] w_n246_1;
	wire[2:0] w_n246_2;
	wire[1:0] w_n248_0;
	wire[1:0] w_n250_0;
	wire[1:0] w_n251_0;
	wire[1:0] w_n253_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n257_0;
	wire[1:0] w_n264_0;
	wire[1:0] w_n265_0;
	wire[1:0] w_n269_0;
	wire[1:0] w_n271_0;
	wire[1:0] w_n281_0;
	wire[1:0] w_n288_0;
	wire[1:0] w_n290_0;
	wire w_dff_B_bPjHBH3h8_0;
	wire w_dff_B_yl2terfh9_0;
	wire w_dff_B_nMZ6D5Dx3_0;
	wire w_dff_B_mm8gENSW7_0;
	wire w_dff_B_VtDiiVvS3_0;
	wire w_dff_B_QyI9FYcT2_0;
	wire w_dff_B_UDYFs09n4_0;
	wire w_dff_B_6cLSZGCT2_0;
	wire w_dff_B_haira9qa2_0;
	wire w_dff_B_Xk0lJJfU6_2;
	wire w_dff_A_ecMX45fI9_0;
	wire w_dff_B_3lorr8c26_2;
	wire w_dff_A_5PGDgAJZ2_1;
	wire w_dff_B_arOPje5Y0_1;
	wire w_dff_B_wMWas1jf9_1;
	wire w_dff_B_gwwz2dgp4_1;
	wire w_dff_B_UTeYUHQH9_1;
	wire w_dff_B_4YKhSSsa8_1;
	wire w_dff_B_KwnugGjf3_1;
	wire w_dff_B_zFq2nHU27_1;
	wire w_dff_B_swwBgBw02_1;
	wire w_dff_B_9WkdFLZQ5_1;
	wire w_dff_B_WzV5yZLZ4_1;
	wire w_dff_B_pocnB0Ie0_1;
	wire w_dff_B_gNmCbR4p6_1;
	wire w_dff_B_UVX5Q52q3_1;
	wire w_dff_B_mFrxlkXZ5_1;
	wire w_dff_B_bhNwvLJR9_1;
	wire w_dff_B_NwEF1kHj0_1;
	wire w_dff_B_hNun5WHj5_1;
	wire w_dff_B_m3FlmHAJ4_1;
	wire w_dff_B_3rIGQKTy5_1;
	wire w_dff_B_oZQrNMZb0_1;
	wire w_dff_B_YQ88Mjss7_1;
	wire w_dff_B_qmBZId8f7_1;
	wire w_dff_B_MqXRGYB47_1;
	wire w_dff_B_sWI2zR2Z2_1;
	wire w_dff_B_L6dqpViB0_2;
	wire w_dff_A_lk5oN2Px8_0;
	wire w_dff_A_YmGPrnxB0_0;
	wire w_dff_A_sQdHh1n37_0;
	wire w_dff_B_T4nIGQqQ2_1;
	wire w_dff_A_pLGLSxkP3_0;
	wire w_dff_A_6Feo5qj86_0;
	wire w_dff_A_VufXFsyk5_0;
	wire w_dff_A_lDO0LMfw6_0;
	wire w_dff_A_w6gnDch55_0;
	wire w_dff_A_K4aNRt418_0;
	wire w_dff_B_2uLaRsxG9_1;
	wire w_dff_B_1sNgVaS14_1;
	wire w_dff_B_C2r8BW9j4_1;
	wire w_dff_B_CyXqCiNp0_1;
	wire w_dff_B_ybIFUs8m1_1;
	wire w_dff_B_K7INepNu6_1;
	wire w_dff_B_sm8nqeof3_1;
	wire w_dff_B_Gt05Sxcy8_0;
	wire w_dff_B_F5NQ7doP6_0;
	wire w_dff_B_1DnC2YYM8_0;
	wire w_dff_B_Ia4EvD1F4_0;
	wire w_dff_A_y06fDyTX5_1;
	wire w_dff_A_00iMpKMO8_1;
	wire w_dff_A_kw7p7WYb9_1;
	wire w_dff_A_n5gMisvx6_1;
	wire w_dff_A_clcYDvzU5_1;
	wire w_dff_B_YYPEZ8R58_1;
	wire w_dff_B_qSKNWnMq2_0;
	wire w_dff_A_ZeHLK5Up7_0;
	wire w_dff_A_RLuC4rbH2_0;
	wire w_dff_A_KjzGsVNx1_0;
	wire w_dff_A_45igkSop1_0;
	wire w_dff_A_xBPB0U0t7_0;
	wire w_dff_A_RLkBIp1p8_0;
	wire w_dff_A_RolMB63E2_0;
	wire w_dff_A_e2DkesIj1_0;
	wire w_dff_A_VLqdQm978_0;
	wire w_dff_A_Cit0T6vd5_0;
	wire w_dff_A_1IQXxtG49_0;
	wire w_dff_B_5QBn9vwG9_2;
	wire w_dff_B_UvZaV2l65_2;
	wire w_dff_B_Jcb2xc3Y9_2;
	wire w_dff_B_IPfJvSUz0_2;
	wire w_dff_B_lKj5Z0wb7_2;
	wire w_dff_B_GsCLyO7a6_2;
	wire w_dff_B_ckcbK40t4_2;
	wire w_dff_B_zbMJB66E0_2;
	wire w_dff_B_pBv53cVB3_2;
	wire w_dff_B_u1gy6WZq5_2;
	wire w_dff_B_JK1MxHSR1_2;
	wire w_dff_B_wxTuSRiP1_2;
	wire w_dff_B_Y5QRsITF6_2;
	wire w_dff_B_ZpqHa7210_2;
	wire w_dff_A_Twl7KQTI4_0;
	wire w_dff_A_2AwORB5l2_0;
	wire w_dff_A_NRKkQU364_0;
	wire w_dff_A_YW6uijQe5_0;
	wire w_dff_A_keTKdMYW4_0;
	wire w_dff_A_xvjiRNkU4_0;
	wire w_dff_A_zFeo3qiT8_0;
	wire w_dff_A_KYaFkvxH3_0;
	wire w_dff_A_AQs67B543_0;
	wire w_dff_A_GCx0MWnl7_0;
	wire w_dff_A_FkjMFXXK7_0;
	wire w_dff_B_pyvjmihX0_2;
	wire w_dff_B_Rqoa51le1_2;
	wire w_dff_B_FVRNWe4T3_2;
	wire w_dff_B_2aIldgDc7_2;
	wire w_dff_B_3MW6ahhJ6_2;
	wire w_dff_B_JN560gq67_2;
	wire w_dff_B_JiWso3Dt5_2;
	wire w_dff_B_aoExucFl0_2;
	wire w_dff_B_aUO21Keg9_2;
	wire w_dff_B_D9Qw4Dr58_2;
	wire w_dff_B_Ctc46mOx3_2;
	wire w_dff_B_oPIgScKF0_2;
	wire w_dff_B_x2nzTAyz6_2;
	wire w_dff_B_11kHvXQO6_2;
	wire w_dff_B_EWMUwY8D6_1;
	wire w_dff_B_NoK4utvG1_1;
	wire w_dff_B_dWPghv9I9_1;
	wire w_dff_B_dt9IvtXm4_1;
	wire w_dff_B_9lW2wGo79_1;
	wire w_dff_B_NZTeA8Qx8_1;
	wire w_dff_B_YcQdMbcb1_1;
	wire w_dff_B_REjk8CP10_1;
	wire w_dff_B_4qvRdGYB5_1;
	wire w_dff_B_3wJs1hff5_1;
	wire w_dff_B_JsbSEA9S6_1;
	wire w_dff_B_cHIierqT4_1;
	wire w_dff_B_fuA4Pupk1_1;
	wire w_dff_B_V6kzopNN6_1;
	wire w_dff_B_q7cwNexr6_1;
	wire w_dff_B_23izKn4C8_1;
	wire w_dff_B_ASLHyAfW8_1;
	wire w_dff_B_idwTemFi1_1;
	wire w_dff_B_5Ugyj6ki2_1;
	wire w_dff_B_ls6Ys0ht3_1;
	wire w_dff_B_rnRxmECU0_1;
	wire w_dff_B_8XewBiFj9_1;
	wire w_dff_B_Fk3MAnap5_1;
	wire w_dff_B_w2tuWnAq2_1;
	wire w_dff_B_MQS63P3w3_1;
	wire w_dff_B_2rjG9oEl4_1;
	wire w_dff_B_M3IeiHw62_1;
	wire w_dff_B_1ab0SRD63_1;
	wire w_dff_A_qEHxUWUw7_0;
	wire w_dff_A_nmowiDWS1_0;
	wire w_dff_A_wtAqk43u5_0;
	wire w_dff_A_o5aZb5hM7_0;
	wire w_dff_A_KfpRo5LZ4_0;
	wire w_dff_B_w3nCi8Ca7_2;
	wire w_dff_B_X9S9FndA7_2;
	wire w_dff_B_Poaye4d59_2;
	wire w_dff_B_aqUtM0TL6_2;
	wire w_dff_B_BrvhUVLZ7_2;
	wire w_dff_B_pjjIQtIO9_2;
	wire w_dff_B_cU2FmDGn3_2;
	wire w_dff_B_L2vDqohC6_2;
	wire w_dff_B_Q7kbfaUg1_2;
	wire w_dff_B_63kkTZgB6_2;
	wire w_dff_B_ggr7m1UT8_2;
	wire w_dff_B_SOcydkLC5_2;
	wire w_dff_B_7yBeHPJ67_2;
	wire w_dff_B_8zFPGK4q8_2;
	wire w_dff_B_Dxuofd8Z2_2;
	wire w_dff_A_T9mV3NnG5_0;
	wire w_dff_A_OZYfqWzk6_0;
	wire w_dff_A_aUFXydqr0_0;
	wire w_dff_A_iyzUq9O70_0;
	wire w_dff_A_xQpPy1Km9_0;
	wire w_dff_B_4HDTrH7R5_2;
	wire w_dff_B_u1Yo01bb8_2;
	wire w_dff_B_G8MiyEs00_2;
	wire w_dff_B_H31XRr0r0_2;
	wire w_dff_B_G5dnU2xU5_2;
	wire w_dff_B_sMGCvCnC6_2;
	wire w_dff_B_OEi3EvXT8_2;
	wire w_dff_B_hUJnCLyW7_2;
	wire w_dff_B_jxfeYicl8_2;
	wire w_dff_B_htpEslNe9_2;
	wire w_dff_B_8Hw6z0XB2_2;
	wire w_dff_B_FNTAziHu9_2;
	wire w_dff_B_urenHQeE1_2;
	wire w_dff_B_Ao6Eg4Y10_2;
	wire w_dff_A_PbtSaNKS8_0;
	wire w_dff_A_u0WAQt203_0;
	wire w_dff_A_crKpqWTZ5_0;
	wire w_dff_A_ls0Xmgj72_0;
	wire w_dff_A_BHv2sUzV1_0;
	wire w_dff_A_npMJPdxG5_0;
	wire w_dff_A_2cuzIc1f9_0;
	wire w_dff_A_HkdP4Wa46_0;
	wire w_dff_A_re46KwVH6_0;
	wire w_dff_B_LR9dAh5R7_1;
	wire w_dff_B_B7W15AHw3_0;
	wire w_dff_A_XrnIk4bn8_0;
	wire w_dff_A_2ot3g6Jk2_0;
	wire w_dff_A_X3C8Pmc37_0;
	wire w_dff_A_xQdhGddt2_0;
	wire w_dff_A_XWQsult97_0;
	wire w_dff_A_Q6oFFsFn8_0;
	wire w_dff_A_bW5LykPj5_0;
	wire w_dff_A_JXKToiTb4_0;
	wire w_dff_A_PXdvU1ov1_0;
	wire w_dff_A_em0haHZN6_0;
	wire w_dff_A_2e6k5BFq9_0;
	wire w_dff_A_tdukIwAy8_0;
	wire w_dff_A_M29Fgj9d8_0;
	wire w_dff_A_xTlXDaKf3_0;
	wire w_dff_A_t1lvHTWN3_0;
	wire w_dff_A_gQ4GPX5n4_0;
	wire w_dff_A_bcu8cZWX0_0;
	wire w_dff_A_HozFfQbX4_0;
	wire w_dff_A_5Y8CGgZd9_0;
	wire w_dff_A_9dtdvi1f9_0;
	wire w_dff_A_OPd7hUjC2_0;
	wire w_dff_A_fdKUXmEi0_0;
	wire w_dff_A_ZzhT5Luj8_0;
	wire w_dff_A_FeSuzuR20_0;
	wire w_dff_A_Bk0xriSz6_0;
	wire w_dff_A_pSUpvoc61_0;
	wire w_dff_A_TeHHmgXQ8_0;
	wire w_dff_A_c897qPZX6_0;
	wire w_dff_A_m2FxBFAN5_0;
	wire w_dff_A_BrB88TYv0_0;
	wire w_dff_A_TE5ZFhsM0_0;
	wire w_dff_A_B8wPd7556_0;
	wire w_dff_A_gxksOdZQ9_0;
	wire w_dff_A_SUSk2GZb9_0;
	wire w_dff_A_w9cGeVtq8_0;
	wire w_dff_A_MYdu8TrK4_0;
	wire w_dff_A_XPwPzKIp6_0;
	wire w_dff_A_9IRuOFH21_0;
	wire w_dff_A_IUafJYUi9_0;
	wire w_dff_A_k7Ha5SNK8_0;
	wire w_dff_A_EC2q37lL9_0;
	wire w_dff_A_77MK1I3v7_0;
	wire w_dff_A_mSy5WXBu8_0;
	wire w_dff_A_EQPuw4Xx8_0;
	wire w_dff_A_ZEM7Owvf2_0;
	wire w_dff_A_3jxfSrxU6_0;
	wire w_dff_A_4vCTaY2l7_0;
	wire w_dff_A_ge7cvY329_0;
	wire w_dff_A_nKvyGjSi1_0;
	wire w_dff_A_s80YZnEh9_0;
	wire w_dff_A_2tdWEtSC8_0;
	wire w_dff_A_B20RmEEi8_0;
	wire w_dff_A_ul9HRwnU4_0;
	wire w_dff_A_A0eZaJkW1_0;
	wire w_dff_A_Htdhkaoi2_0;
	wire w_dff_A_sHVhMF8S9_0;
	wire w_dff_A_mnRhacPx5_1;
	wire w_dff_A_zP7Ve7Rj5_1;
	wire w_dff_A_9WgDQZaW4_1;
	wire w_dff_A_rH22nS0W6_1;
	wire w_dff_A_FVBT3PBs0_1;
	wire w_dff_A_UcHNbOBb1_1;
	wire w_dff_A_a4uJBmZA5_1;
	wire w_dff_A_McnMWF4i8_1;
	wire w_dff_A_kh3xpoMR7_1;
	wire w_dff_A_FSe6SYPE6_1;
	wire w_dff_A_AHjkNldU9_1;
	wire w_dff_A_DkAf5t1k3_1;
	wire w_dff_A_6JHxCAyW2_1;
	wire w_dff_A_4LA2JJJp0_1;
	wire w_dff_A_YT8iWFLb1_1;
	wire w_dff_A_5YFQazP93_0;
	wire w_dff_A_nPCNiFv90_0;
	wire w_dff_A_fCmm0Yfz5_0;
	wire w_dff_A_R2rr5sTk3_0;
	wire w_dff_A_iXbJSuJB2_0;
	wire w_dff_A_URiQhGSh9_0;
	wire w_dff_A_omBVryHd6_0;
	wire w_dff_A_rdeVdRNz3_0;
	wire w_dff_A_9oXFHW0V8_0;
	wire w_dff_A_b6jPoXU51_0;
	wire w_dff_A_LsBEZ58d8_0;
	wire w_dff_A_ggeOITuZ3_0;
	wire w_dff_A_6xg5YICe5_0;
	wire w_dff_A_0fZNLKVp9_0;
	wire w_dff_A_3rxHug5I6_0;
	wire w_dff_A_SmMkBNte8_0;
	wire w_dff_A_7oKWTgbK1_0;
	wire w_dff_A_8c7QOeGs8_0;
	wire w_dff_A_qNYUmA6T4_0;
	wire w_dff_A_oYrNu0tu8_0;
	wire w_dff_A_0uYgz50H6_0;
	wire w_dff_A_t1Pd64y51_0;
	wire w_dff_A_uQBwZtPd6_0;
	wire w_dff_A_Ffetb79U9_0;
	wire w_dff_A_XLIG9Ewp3_0;
	wire w_dff_A_B9LX9zz21_0;
	wire w_dff_A_oWXfa6Cc4_1;
	wire w_dff_A_rdmP5a6T0_1;
	wire w_dff_A_RzYyp0Ox5_1;
	wire w_dff_A_ZMBjp6Q04_1;
	wire w_dff_A_nYGzuNUw7_1;
	wire w_dff_A_u10Rjnzn5_1;
	wire w_dff_A_xDbOsd0l1_1;
	wire w_dff_A_fdyWZa240_1;
	wire w_dff_A_0Y0QXG8n4_1;
	wire w_dff_A_AQjnpTW43_1;
	wire w_dff_A_pTR124rD5_1;
	wire w_dff_A_RNUZXDNp4_1;
	wire w_dff_A_NKQ4mBEE9_1;
	wire w_dff_A_RXeTVk6A3_1;
	wire w_dff_A_iA559QVq3_1;
	wire w_dff_B_TSGJYjC88_1;
	wire w_dff_B_Vor8q6b36_1;
	wire w_dff_B_t1m9d1w16_1;
	wire w_dff_B_h1iPyZE83_1;
	wire w_dff_B_0zhaWSMg6_1;
	wire w_dff_A_YA4T75yo6_0;
	wire w_dff_A_hodyrOoN8_0;
	wire w_dff_A_7QvCauur8_0;
	wire w_dff_A_D0tRt7ml1_0;
	wire w_dff_A_DGCf7jsN3_0;
	wire w_dff_A_L4RaDarK3_0;
	wire w_dff_A_fMGEdRT69_0;
	wire w_dff_A_k5vx8KWr9_0;
	wire w_dff_A_iKdmFnYb9_0;
	wire w_dff_A_HfdzV5iC9_0;
	wire w_dff_A_aLG49hB42_0;
	wire w_dff_A_ueuykuks7_0;
	wire w_dff_A_ZhVJwpZO3_0;
	wire w_dff_A_YJBSrbur9_0;
	wire w_dff_A_iWhog36v9_0;
	wire w_dff_A_M2OIffg29_0;
	wire w_dff_A_u07h95AP6_0;
	wire w_dff_A_4T3hAL9z2_0;
	wire w_dff_A_LoBPcUcI0_0;
	wire w_dff_A_40SG9CPg4_0;
	wire w_dff_A_NMf0EbFR5_1;
	wire w_dff_A_9XnP4ArK7_1;
	wire w_dff_A_tJAVIllD3_1;
	wire w_dff_A_NMUZW6aA8_1;
	wire w_dff_A_ajNIy8Tk0_1;
	wire w_dff_A_4X8tPYDK9_1;
	wire w_dff_A_kwZueTpZ6_1;
	wire w_dff_A_GYzVYy4W4_1;
	wire w_dff_A_ICeUlMas8_1;
	wire w_dff_A_G1YXUitm2_1;
	wire w_dff_A_UbNZK9ix3_1;
	wire w_dff_A_k1WU7RTL7_1;
	wire w_dff_A_K2oUXlZz3_1;
	wire w_dff_A_A1DlU1gM0_1;
	wire w_dff_A_0ARvSZ8F9_1;
	wire w_dff_A_GqUV8JKA9_0;
	wire w_dff_A_48eaq5Ir5_0;
	wire w_dff_A_NvyiPqS37_0;
	wire w_dff_A_wuz6Fc069_0;
	wire w_dff_A_B9lTBLGU4_0;
	wire w_dff_A_r0oD3pQw5_0;
	wire w_dff_A_TXKiECU73_0;
	wire w_dff_A_mp9hLhBg7_0;
	wire w_dff_A_RhnNqOOW1_0;
	wire w_dff_A_sottCIB02_0;
	wire w_dff_A_rwc6q2dn2_0;
	wire w_dff_A_gxtiFyyH8_0;
	wire w_dff_A_xbnXnNeJ5_0;
	wire w_dff_A_3vOkVf0c5_0;
	wire w_dff_A_S9Y8jeJ59_0;
	wire w_dff_A_2nMf8lIr9_1;
	wire w_dff_B_hgRNJLr90_0;
	wire w_dff_B_8toNLRwD6_0;
	wire w_dff_B_YrCFl0P75_0;
	wire w_dff_B_TXJwmJs32_0;
	wire w_dff_B_T6Rc6Deo2_0;
	wire w_dff_B_paiVXyJb5_0;
	wire w_dff_A_VDhjwMVA7_0;
	wire w_dff_A_HCaIh7oj7_0;
	wire w_dff_A_N8jagXYC1_0;
	wire w_dff_A_GCm9gLmv1_0;
	wire w_dff_A_H3at82mu6_0;
	wire w_dff_A_pPnQxv1e3_0;
	wire w_dff_A_WDJJMe4c4_0;
	wire w_dff_A_zEsNOJXv9_0;
	wire w_dff_A_iajL2Dnv6_0;
	wire w_dff_A_ti2L8lQ49_0;
	wire w_dff_A_fy2ss3vq8_0;
	wire w_dff_A_O0wQlBzA7_0;
	wire w_dff_B_fzzC41Ff8_2;
	wire w_dff_B_SdaI9yDV7_2;
	wire w_dff_B_lVeuFj7i3_2;
	wire w_dff_B_l967Xkaa4_2;
	wire w_dff_B_PgL5sdK07_2;
	wire w_dff_B_F5KTOii04_2;
	wire w_dff_B_nRqDZMM19_2;
	wire w_dff_A_ETQstGiG0_0;
	wire w_dff_A_zZbIzLg79_0;
	wire w_dff_A_DbGLIGMI4_0;
	wire w_dff_A_pKRwmpZK3_0;
	wire w_dff_A_fhi3Q4gO4_0;
	wire w_dff_A_2dwXvW6g6_0;
	wire w_dff_A_E0sjAgrb3_0;
	wire w_dff_A_I1CYUHlT3_0;
	wire w_dff_A_KGSJOwy29_0;
	wire w_dff_A_Hp1puBtR0_0;
	wire w_dff_A_QlDhJh9o1_0;
	wire w_dff_A_15CWYWUg3_0;
	wire w_dff_A_U5XpNZBA8_0;
	wire w_dff_A_oTYYasxg4_0;
	wire w_dff_A_tLUHc9pw8_0;
	wire w_dff_A_Wispl0754_0;
	wire w_dff_A_BJdJbONd7_0;
	wire w_dff_A_vB8S38w90_0;
	wire w_dff_A_PjoCkbYc5_0;
	wire w_dff_A_nWrydaZy0_0;
	wire w_dff_A_i11qy3oI3_0;
	wire w_dff_B_9Ejn8SAM9_1;
	wire w_dff_B_b99rtdSG1_1;
	wire w_dff_B_O81W0fyS3_1;
	wire w_dff_B_0ibJyFA01_1;
	wire w_dff_B_ZT584fq39_1;
	wire w_dff_B_1YSV3hag4_1;
	wire w_dff_B_wxeByVvQ8_1;
	wire w_dff_B_JB9geFc13_1;
	wire w_dff_A_VbA1FYqv1_0;
	wire w_dff_A_3zMzafxQ0_0;
	wire w_dff_A_7chVJTYT4_0;
	wire w_dff_A_3lOcn6Ae6_0;
	wire w_dff_A_jRx41jlR4_0;
	wire w_dff_A_Iaa9LfoL2_0;
	wire w_dff_A_xlMAHoDw3_0;
	wire w_dff_A_WtCqoIhw8_0;
	wire w_dff_A_eMJEcvRX9_0;
	wire w_dff_A_6qyoy6ti4_0;
	wire w_dff_A_INV8YbR14_0;
	wire w_dff_A_QPC3tFcH5_0;
	wire w_dff_A_ulPa3Dcx5_0;
	wire w_dff_A_mdg1Qcp65_0;
	wire w_dff_A_XYS1mqVo8_0;
	wire w_dff_A_j6MGPAlk3_0;
	wire w_dff_A_f0KLnLm14_0;
	wire w_dff_A_8KnHbGtN8_0;
	wire w_dff_B_D3rm779A3_2;
	wire w_dff_B_VLsBj1Ob3_2;
	wire w_dff_B_a3N31SVR7_2;
	wire w_dff_B_wRLyrwcF8_2;
	wire w_dff_B_xxWt0xOr8_2;
	wire w_dff_B_0oOVepwL9_2;
	wire w_dff_B_LjiddWGy7_2;
	wire w_dff_A_75b5ul9A3_0;
	wire w_dff_A_Hc0Amted6_0;
	wire w_dff_A_JR78ul7R6_0;
	wire w_dff_A_Vkbw9zmX5_0;
	wire w_dff_A_vxywRz2Y0_0;
	wire w_dff_A_iXLtYgTW0_0;
	wire w_dff_A_HasXKJGy4_0;
	wire w_dff_A_8MlS1o3V7_0;
	wire w_dff_A_dNA4oHAQ7_0;
	wire w_dff_A_qFtG1D614_0;
	wire w_dff_A_ZZTgA83A1_0;
	wire w_dff_B_s9JpqwuC2_2;
	wire w_dff_B_zjrwG2rx1_2;
	wire w_dff_B_vo65AGxd4_2;
	wire w_dff_B_CDxLi0nf7_2;
	wire w_dff_B_TOOniKQo0_2;
	wire w_dff_B_sZxPAbMC2_2;
	wire w_dff_B_2383nTjN5_2;
	wire w_dff_B_UuWpBk8e4_1;
	wire w_dff_B_5jEXFLQw6_0;
	wire w_dff_A_wD8pm91g9_0;
	wire w_dff_A_B6bWZbTF0_0;
	wire w_dff_A_0MQiOCrZ5_0;
	wire w_dff_A_t26TpBhl1_0;
	wire w_dff_A_3FgFJ1Ds0_0;
	wire w_dff_A_dZUWnc8V7_0;
	wire w_dff_A_YYp97nOP6_0;
	wire w_dff_A_pHKS3yWJ1_0;
	wire w_dff_A_3bj74WQe9_0;
	wire w_dff_A_6ggCqFz20_0;
	wire w_dff_A_SlqBgjwD3_0;
	wire w_dff_B_6DwJa8ak8_2;
	wire w_dff_B_zpb7GV5u3_2;
	wire w_dff_B_co8Qk23n1_2;
	wire w_dff_B_q3JMA5Vy5_2;
	wire w_dff_B_iWkayhoz4_2;
	wire w_dff_B_cU3JyvQs4_2;
	wire w_dff_B_d94g1jne5_2;
	wire w_dff_A_Wd71qjV00_0;
	wire w_dff_A_vBHMAZOb3_0;
	wire w_dff_A_tf5nt8KM8_0;
	wire w_dff_A_wXORQXsF8_0;
	wire w_dff_A_7m7OL1VZ1_0;
	wire w_dff_A_HfQCzGGO4_0;
	wire w_dff_A_qdhEkhzh8_0;
	wire w_dff_A_h7uXJ1Za4_0;
	wire w_dff_A_HpukHOts3_0;
	wire w_dff_A_Df2fqTGy2_0;
	wire w_dff_A_iVbpCoSB7_0;
	wire w_dff_B_3NJJVuIR5_2;
	wire w_dff_B_xrr3inuy9_2;
	wire w_dff_B_lXatA0Gb7_2;
	wire w_dff_B_Q7cnN83r4_2;
	wire w_dff_B_T48b5iB48_2;
	wire w_dff_B_lYBSgovx5_2;
	wire w_dff_B_xZXqVwxy2_2;
	wire w_dff_B_0djgFnjH6_1;
	wire w_dff_B_2cWYEqb12_1;
	wire w_dff_B_fss9v9pb7_1;
	wire w_dff_B_tvSybPBs1_1;
	wire w_dff_B_Ylua8ZW21_1;
	wire w_dff_B_z4KKWFh40_1;
	wire w_dff_B_69IWdBfv7_1;
	wire w_dff_A_etusTHS08_0;
	wire w_dff_A_xSnmWATm5_0;
	wire w_dff_A_mtTomtmr4_0;
	wire w_dff_A_eC3ulkGY4_0;
	wire w_dff_A_O7ir2tha6_0;
	wire w_dff_A_zIBHdoei7_0;
	wire w_dff_A_5A7yxSpN6_0;
	wire w_dff_A_z9HeE6j80_0;
	wire w_dff_A_E2as1UsJ9_0;
	wire w_dff_A_w5h8NoPN9_0;
	wire w_dff_A_Vpuez0BJ8_0;
	wire w_dff_B_hvYkcC6P7_2;
	wire w_dff_B_bEFYQsCV1_2;
	wire w_dff_B_zPzNNgvb9_2;
	wire w_dff_B_jHY2UP930_2;
	wire w_dff_B_El9v8IRk6_2;
	wire w_dff_B_svnRpbIj0_2;
	wire w_dff_B_zXMf2XEi9_2;
	wire w_dff_A_yGXAjNQO9_1;
	wire w_dff_A_hD07DT974_1;
	wire w_dff_A_6y0FKlIA3_1;
	wire w_dff_A_lzWotW326_1;
	wire w_dff_A_U7C7JYPf9_1;
	wire w_dff_A_tsHqbiwq9_1;
	wire w_dff_A_0TP2qSA35_1;
	wire w_dff_A_Nhge5zT49_1;
	wire w_dff_A_btuvgOL03_1;
	wire w_dff_A_s10MHrKl5_1;
	wire w_dff_A_Y3y0ffj90_1;
	wire w_dff_A_eri90pHm3_1;
	wire w_dff_A_veiJWYq83_1;
	wire w_dff_A_93LQLPH25_1;
	wire w_dff_A_H0izGr0v9_1;
	wire w_dff_A_pWDz6cub2_0;
	wire w_dff_A_XgPVrpW43_0;
	wire w_dff_A_kqq7ADov6_0;
	wire w_dff_A_inpDNTQ21_0;
	wire w_dff_A_QSBh61bw9_0;
	wire w_dff_B_ByfiAHEG9_2;
	wire w_dff_B_yebf95lj0_2;
	wire w_dff_B_4P4Dj14L1_2;
	wire w_dff_B_2rPpI94R8_2;
	wire w_dff_B_3Ld2ROdY9_2;
	wire w_dff_B_MjrbvAuh6_2;
	wire w_dff_B_drRRZsue3_2;
	wire w_dff_B_MJhrWLMi7_2;
	wire w_dff_B_cObmXuED5_2;
	wire w_dff_B_8VuazdCD8_2;
	wire w_dff_B_k2SiN4JA2_2;
	wire w_dff_B_bqYDk4FS7_2;
	wire w_dff_B_X44NYGyM9_2;
	wire w_dff_B_zxrmMO796_2;
	wire w_dff_A_gaYOyXy37_0;
	wire w_dff_A_Mjlub2SV9_0;
	wire w_dff_A_8RjYcBBN2_0;
	wire w_dff_A_MkCc97db5_0;
	wire w_dff_A_hfzKUSQM4_0;
	wire w_dff_A_KUzs6dp26_0;
	wire w_dff_A_itPQSgbR6_0;
	wire w_dff_A_0XbUR4kT0_0;
	wire w_dff_A_ICPe4uHu8_0;
	wire w_dff_A_35SPAG2C1_0;
	wire w_dff_A_HXJgagCy8_0;
	wire w_dff_A_WHHALaDU3_0;
	wire w_dff_A_n57mvHM27_0;
	wire w_dff_A_EZ7PtoxU8_0;
	wire w_dff_A_4Hbif21O6_0;
	wire w_dff_A_vWsW9iQT5_0;
	wire w_dff_A_vEY9DlgU3_0;
	wire w_dff_A_zqEVtEAi9_0;
	wire w_dff_A_hDvUd3Kn1_0;
	wire w_dff_A_Y0v3swMy4_0;
	wire w_dff_A_sH5qWaTd4_0;
	wire w_dff_B_SDhLMKyS7_1;
	wire w_dff_B_xhPinsnU9_1;
	wire w_dff_A_bwF9LVaO1_0;
	wire w_dff_A_kQKLUrFv0_0;
	wire w_dff_A_i6lNTESq6_0;
	wire w_dff_A_90rAaKG98_0;
	wire w_dff_A_OlIjdwvL0_0;
	wire w_dff_A_8MfW7LCP6_0;
	wire w_dff_A_oQ31W50A7_0;
	wire w_dff_A_PNAk39HP3_0;
	wire w_dff_A_5EYzQs590_1;
	wire w_dff_A_ixdHPJ1C3_1;
	wire w_dff_A_UF9pdw1g6_1;
	wire w_dff_A_vNj5IGle3_1;
	wire w_dff_A_E1ZEBn9q1_1;
	wire w_dff_A_aEg1lPsR1_1;
	wire w_dff_A_Zf9CVxiy8_1;
	wire w_dff_A_xG03RLPb7_1;
	wire w_dff_A_rfXJqbez5_1;
	wire w_dff_A_n7eXfFcT5_1;
	wire w_dff_A_ET9R53Hk4_1;
	wire w_dff_A_tQ1hlDZD4_1;
	wire w_dff_A_wKWGJvJL1_1;
	wire w_dff_A_yfnhmTCl5_0;
	wire w_dff_A_g8narcgG7_0;
	wire w_dff_A_cEMPf0c93_0;
	wire w_dff_A_F5ALTxrE4_0;
	wire w_dff_A_9mhHPHMj0_0;
	wire w_dff_A_I1Wv4zCs2_0;
	wire w_dff_A_7gXa9zaa1_0;
	wire w_dff_A_jSH4mWPk3_0;
	wire w_dff_A_Cb8WFyt35_0;
	wire w_dff_A_Af1YuSND4_0;
	wire w_dff_A_7cD3xAYU8_0;
	wire w_dff_A_pgLAn1sp3_0;
	wire w_dff_A_uox7brt46_0;
	wire w_dff_A_s2qg08bX5_0;
	wire w_dff_A_CV8VZeWM0_0;
	wire w_dff_A_ejGkuxo42_0;
	wire w_dff_A_sHFDSFSc4_0;
	wire w_dff_A_b5MePVBU6_0;
	wire w_dff_A_22AEj7LU2_0;
	wire w_dff_A_vCaMbch46_1;
	wire w_dff_A_fbLuwnPe8_1;
	wire w_dff_A_r8IsYw6s7_1;
	wire w_dff_A_mbUctylG5_1;
	wire w_dff_A_ToATTP9q1_1;
	wire w_dff_A_6knYgbo40_1;
	wire w_dff_A_uKFuaD5e9_1;
	wire w_dff_A_jKSTLNsP8_1;
	wire w_dff_A_SvvGCQpD9_0;
	wire w_dff_A_DJpB76TI8_0;
	wire w_dff_A_ZTRatxce3_0;
	wire w_dff_A_R2fQV0xr7_0;
	wire w_dff_A_8x7MykNQ2_0;
	wire w_dff_A_RIKbZ0pK9_0;
	wire w_dff_A_Jndz8GqG8_0;
	wire w_dff_A_4knAMhm52_0;
	wire w_dff_A_PhVqGSUi3_0;
	wire w_dff_A_3KDphlJv9_0;
	wire w_dff_A_LFVeGlqI9_0;
	wire w_dff_A_QO8QSwik2_0;
	wire w_dff_A_qm0W7TaO1_0;
	wire w_dff_A_XUgkw1wy5_0;
	wire w_dff_A_eRpb26Ny0_0;
	wire w_dff_A_KSlA7fia0_0;
	wire w_dff_A_KuQL11Dh4_0;
	wire w_dff_A_hjmAjkzM8_0;
	wire w_dff_A_a8rZTlo97_0;
	wire w_dff_A_4jBlvItX0_1;
	wire w_dff_A_4lh03M5a6_1;
	wire w_dff_A_seaIE4A83_1;
	wire w_dff_A_rpIXkCx68_1;
	wire w_dff_A_g7R3sdOn7_1;
	wire w_dff_A_xIUS5okl1_1;
	wire w_dff_A_hMgvqrlX6_1;
	wire w_dff_A_e7w7KJmh4_1;
	wire w_dff_A_quDyM02J4_1;
	wire w_dff_A_bNchDfR86_1;
	wire w_dff_A_sx1E2CEi3_1;
	wire w_dff_A_Oe3fGkx99_1;
	wire w_dff_A_j5ZFPF3W7_1;
	wire w_dff_A_dJET2pmo5_1;
	wire w_dff_A_HsOYiziO0_1;
	wire w_dff_A_q34n06QX0_1;
	wire w_dff_A_Kjwjci5j6_0;
	wire w_dff_A_z9Sk57lB4_0;
	wire w_dff_A_z6wjh8qw1_0;
	wire w_dff_A_J19xxwDj7_0;
	wire w_dff_A_6OkFu1Y69_0;
	wire w_dff_B_FE8oe3zt8_2;
	wire w_dff_B_AuojKlfi3_2;
	wire w_dff_B_q2orjG034_2;
	wire w_dff_B_C6p35jO67_2;
	wire w_dff_B_yASvzsua5_2;
	wire w_dff_B_kr0qIfqT7_2;
	wire w_dff_B_6F2pPsVZ8_2;
	wire w_dff_A_DKireuJq5_0;
	wire w_dff_A_RDgVdBHK9_0;
	wire w_dff_A_luwGQRjV3_0;
	wire w_dff_A_M9DGxWoU6_0;
	wire w_dff_A_NU7gXzoF7_0;
	wire w_dff_A_jtd3syVZ6_0;
	wire w_dff_A_4lfgGwHj0_0;
	wire w_dff_A_6pkMR3F53_0;
	wire w_dff_A_VOCbAonh0_0;
	wire w_dff_A_XTmcFUYU3_0;
	wire w_dff_A_GTkSVVkd9_0;
	wire w_dff_A_WJS91CqH3_0;
	wire w_dff_A_YG8qQCjJ1_0;
	wire w_dff_B_L4jdTIV36_1;
	wire w_dff_B_LS2NnnOg9_0;
	wire w_dff_A_da2wEK4W8_0;
	wire w_dff_A_Go4Hd8746_0;
	wire w_dff_A_WBgjazlO6_0;
	wire w_dff_A_oVj8N9zX5_0;
	wire w_dff_A_SiTL53oB4_0;
	wire w_dff_A_0nTKHlM67_0;
	wire w_dff_B_mqLTv3ku5_1;
	wire w_dff_B_hlQwySnz8_1;
	wire w_dff_B_9ZGB8oOo6_1;
	wire w_dff_B_TkvD2zrK6_1;
	wire w_dff_B_MR1RBrVa4_1;
	wire w_dff_B_BOWiELq69_1;
	wire w_dff_A_RwybG6tX0_0;
	wire w_dff_A_LQDAvEqQ9_0;
	wire w_dff_A_XhwvFi4t7_0;
	wire w_dff_A_iQfPExlA8_0;
	wire w_dff_A_H04Op4pX0_0;
	wire w_dff_A_T5dfnjWx3_0;
	wire w_dff_A_P0Cvhqf03_0;
	wire w_dff_A_FgQvTQOT0_0;
	wire w_dff_A_ht2VrqHN6_0;
	wire w_dff_A_QjYuXeHI0_0;
	wire w_dff_A_ml1kpYNG4_0;
	wire w_dff_A_9c1ceGrW5_0;
	wire w_dff_A_Trkf7w596_0;
	wire w_dff_A_wDrIAQlP5_1;
	wire w_dff_A_ucYRhmgI0_1;
	wire w_dff_A_yco0T9be5_1;
	wire w_dff_A_LP808wx15_1;
	wire w_dff_A_3kyqLb242_1;
	wire w_dff_A_d9L3SHvs9_1;
	wire w_dff_A_KibjpU1d0_1;
	wire w_dff_A_vSKhQeS71_1;
	wire w_dff_A_qSALVIPY3_0;
	wire w_dff_A_VlKvZzBP8_0;
	wire w_dff_A_TN1YAt2a0_0;
	wire w_dff_A_l5XM0c368_0;
	wire w_dff_A_6KQD2n7m9_0;
	wire w_dff_A_xrX8NtgM4_0;
	wire w_dff_A_5JTPPUKV8_0;
	wire w_dff_A_WNeU2Jem0_0;
	wire w_dff_A_6ig9zHsH1_0;
	wire w_dff_A_uCFpV3yA3_0;
	wire w_dff_A_C5IXaVC89_0;
	wire w_dff_A_ogyN5u1A2_0;
	wire w_dff_A_NJKvVWLC5_0;
	wire w_dff_A_qxnsOABw3_0;
	wire w_dff_A_tWBVBbx02_0;
	wire w_dff_A_FKNzlUKt6_0;
	wire w_dff_A_RgASNUCH6_0;
	wire w_dff_A_neboB7sP3_0;
	wire w_dff_A_TtTMic2f7_0;
	wire w_dff_A_k1I87nsZ5_1;
	wire w_dff_A_rrmacSUs2_1;
	wire w_dff_A_fmBKZxip6_1;
	wire w_dff_A_zBfsPtvw5_1;
	wire w_dff_A_gx0pTNFj7_1;
	wire w_dff_A_YNJ6AOjQ2_1;
	wire w_dff_A_FmmN99Q40_1;
	wire w_dff_A_0qqjJV1q4_1;
	wire w_dff_A_MAuFFSEN3_0;
	wire w_dff_A_mjQk8Mm64_0;
	wire w_dff_A_978miXAZ9_0;
	wire w_dff_A_JEz8vuUG2_0;
	wire w_dff_A_3JMd7eMd4_0;
	wire w_dff_A_VGxBzT6Y2_0;
	wire w_dff_A_iUhGKo2b6_1;
	wire w_dff_A_S3391bGd9_1;
	wire w_dff_A_NK8WXUTU8_1;
	wire w_dff_A_CbNCsRrk0_1;
	wire w_dff_A_YnnGEYH09_1;
	wire w_dff_A_D620hIjN3_1;
	wire w_dff_A_EA4fEhLh9_0;
	wire w_dff_A_mZeqW5Xc3_0;
	wire w_dff_A_NioHEqBG4_0;
	wire w_dff_A_rHj2NQ2M1_0;
	wire w_dff_A_07mjf78m6_0;
	wire w_dff_A_JWi0SZFn6_0;
	wire w_dff_A_09M2gSEs1_0;
	wire w_dff_A_HWIp2MDX0_0;
	wire w_dff_A_zGPZz4L48_1;
	wire w_dff_A_vMZ8YF8h8_1;
	wire w_dff_A_g38jHedp6_1;
	wire w_dff_A_ePubq2rA8_1;
	wire w_dff_A_J7YzgHXy3_1;
	wire w_dff_A_K3HiBZhZ0_1;
	wire w_dff_A_9R5cDTOQ5_1;
	wire w_dff_A_rJxT69mx2_1;
	wire w_dff_A_pNZ02Kme4_1;
	wire w_dff_A_XPq9qGD88_1;
	wire w_dff_A_GiLn6BOZ3_1;
	wire w_dff_A_am0tLmpk8_1;
	wire w_dff_A_9Sv5mRmP8_1;
	wire w_dff_A_WCZ0mFjC7_0;
	wire w_dff_A_g9gBizeZ1_0;
	wire w_dff_A_loWXzfhA9_0;
	wire w_dff_A_0rNdRn0C5_0;
	wire w_dff_A_nUKewTiJ9_0;
	wire w_dff_A_DnJVo4kj9_0;
	wire w_dff_B_s0c1Tnw43_1;
	wire w_dff_B_rrynMJak1_1;
	wire w_dff_A_Fw0m2RSD9_0;
	wire w_dff_A_0iCzWIbG2_0;
	wire w_dff_A_yE7HAdrQ7_0;
	wire w_dff_A_xm6UIbV59_0;
	wire w_dff_A_7n9LOtu14_0;
	wire w_dff_A_hJNfhKKn3_0;
	wire w_dff_A_t59ejE1I7_0;
	wire w_dff_A_30qGjJbl3_0;
	wire w_dff_A_w5k1SJh39_0;
	wire w_dff_A_w2p70dmt4_0;
	wire w_dff_A_CpT96k2v0_0;
	wire w_dff_A_MTV7oEoe4_0;
	wire w_dff_A_gUjf7bgp9_0;
	wire w_dff_A_U3ECG0Ey4_0;
	wire w_dff_A_BXhbeJ6u9_0;
	wire w_dff_A_BRg9RaPD8_0;
	wire w_dff_A_sjZR4kzv5_0;
	wire w_dff_A_5LMN1alR9_0;
	wire w_dff_A_EghAq9VE0_0;
	wire w_dff_A_pnBdnbqj7_0;
	wire w_dff_A_5iR8ySs13_0;
	wire w_dff_A_TBOhhYWR0_0;
	wire w_dff_A_emfxJcVz0_0;
	wire w_dff_A_oqnyvqRT4_0;
	wire w_dff_A_m5XAkFSM9_0;
	wire w_dff_A_IpSgGjO59_0;
	wire w_dff_A_l45PGS1R4_0;
	wire w_dff_A_7RfAld141_0;
	wire w_dff_A_L2s6nSm88_0;
	wire w_dff_A_GW1TgdPw6_0;
	wire w_dff_A_UUIjfV6H9_0;
	wire w_dff_A_Fe8ugEQt2_0;
	wire w_dff_A_cYeha5vQ3_0;
	wire w_dff_A_zmuJEHr61_0;
	wire w_dff_A_jyBUWZxt2_0;
	wire w_dff_A_qxNhJFFj9_0;
	wire w_dff_A_eMw26Pmx1_0;
	wire w_dff_A_GFmMQHXB9_0;
	wire w_dff_A_oAujPlQh2_0;
	wire w_dff_A_hbs3gKxv1_0;
	wire w_dff_A_izcbH5rk2_0;
	wire w_dff_A_ZJZQzvDr9_0;
	wire w_dff_A_UE9Jyjob2_0;
	wire w_dff_A_sGjbF2kD1_0;
	wire w_dff_A_dHsrHFZ11_0;
	wire w_dff_A_axtwTHXH0_1;
	wire w_dff_A_REgmSQsm0_1;
	wire w_dff_A_LvvHirrd2_1;
	wire w_dff_A_kx8knwZf4_1;
	wire w_dff_A_eJFGdXfV6_1;
	wire w_dff_A_ajfTYSEm0_1;
	wire w_dff_A_A94sENI80_1;
	wire w_dff_A_gpuN8SLz2_1;
	wire w_dff_A_5bE7cs9u1_0;
	wire w_dff_A_7x6ncHxp5_0;
	wire w_dff_A_9JiKSFa46_0;
	wire w_dff_A_La0Lioxn3_0;
	wire w_dff_A_Up8MHMLe2_0;
	wire w_dff_B_egBKhqmp2_2;
	wire w_dff_B_kGUCirf42_2;
	wire w_dff_B_YcbZLqPw5_2;
	wire w_dff_B_iR8KAdii6_2;
	wire w_dff_B_yLq0bkSN3_2;
	wire w_dff_B_5YKmKlW35_2;
	wire w_dff_B_4eM6QmVo7_2;
	wire w_dff_A_ezEMIm566_0;
	wire w_dff_A_hTMZdTzv6_0;
	wire w_dff_A_e7yhCOKA5_0;
	wire w_dff_A_UIfke8RR2_0;
	wire w_dff_A_EY9DA8MV3_0;
	wire w_dff_A_BgwTVaKS1_0;
	wire w_dff_A_QZNzZTnj5_0;
	wire w_dff_A_1fdHG0aV6_0;
	wire w_dff_A_w6VFdMW76_0;
	wire w_dff_A_lk2s9mPd5_0;
	wire w_dff_A_XpQRtSzi7_0;
	wire w_dff_A_3CTgq0pL6_0;
	wire w_dff_A_oOw3wfMq8_0;
	wire w_dff_A_v4cc3wmn1_1;
	wire w_dff_A_U9Iwbpkv7_1;
	wire w_dff_A_1fzvDvob2_1;
	wire w_dff_A_4WvKJtRH4_1;
	wire w_dff_A_yHVOro008_1;
	wire w_dff_A_msO9EwR00_1;
	wire w_dff_A_kIzOScC21_1;
	wire w_dff_A_mkmU92eL9_1;
	wire w_dff_A_pUAz7cfj8_0;
	wire w_dff_A_d4L7to5l9_0;
	wire w_dff_A_lZeKiMiY3_0;
	wire w_dff_A_v6HKAFTI1_0;
	wire w_dff_A_CZqs8dwm3_0;
	wire w_dff_A_zxeppp4M2_0;
	wire w_dff_B_FXFeITBu7_1;
	wire w_dff_B_vtrJgknM1_1;
	wire w_dff_A_nTTTe9KR8_0;
	wire w_dff_A_zYlq5Etq3_0;
	wire w_dff_A_wGNpy5QZ2_0;
	wire w_dff_A_pctuj1dG3_0;
	wire w_dff_A_zSINf0dP3_0;
	wire w_dff_A_EhqGlHxz9_0;
	wire w_dff_A_Swk2Fr2z6_0;
	wire w_dff_A_sL3UCyQ09_0;
	wire w_dff_A_FOWyX1XP9_0;
	wire w_dff_A_FWkn7Djz2_0;
	wire w_dff_A_H92DG0GL3_0;
	wire w_dff_A_C9MKShi57_0;
	wire w_dff_A_8NwcASrU2_0;
	wire w_dff_A_QxQf8HVV3_2;
	wire w_dff_A_Lw6AVonP7_0;
	wire w_dff_A_sgLv7Sqh6_0;
	wire w_dff_A_qCEbS0iY1_0;
	wire w_dff_A_Xm31pBam3_0;
	wire w_dff_A_kzPWKD4u9_0;
	wire w_dff_A_m0axmQEX1_0;
	wire w_dff_A_SDsstCuO9_1;
	wire w_dff_A_8wKgaRna2_0;
	wire w_dff_A_uryQFvw91_0;
	wire w_dff_A_w8aiLEMO9_0;
	wire w_dff_A_mDfcpBla1_0;
	wire w_dff_A_ErQX5kCv7_0;
	wire w_dff_A_69aeXXNp3_0;
	wire w_dff_A_YfnHZVw77_0;
	wire w_dff_A_8zuRIUjp8_0;
	wire w_dff_A_SHlor39q6_0;
	wire w_dff_A_5XHH9LnT2_0;
	wire w_dff_A_DCEaacXu6_0;
	wire w_dff_A_zO9u0GcB2_0;
	wire w_dff_A_s6eqjM6c5_0;
	wire w_dff_A_EYXFSrfy1_2;
	wire w_dff_A_HMjUPUtq6_0;
	wire w_dff_A_Yp7kiGvO6_0;
	wire w_dff_A_F5QxENqL9_0;
	wire w_dff_A_SwLhpr7g5_0;
	wire w_dff_A_uyak5vtX8_0;
	wire w_dff_A_5c5qQ5998_0;
	wire w_dff_A_jsSRzS613_1;
	wire w_dff_A_Yle2qnlC2_0;
	wire w_dff_A_pM0DdqxR2_0;
	wire w_dff_A_uWU4UWII3_0;
	wire w_dff_A_SbPzlKR21_0;
	wire w_dff_A_hsy488Jo2_0;
	wire w_dff_A_jJ4botKv4_0;
	wire w_dff_A_MLFC6cQL6_0;
	wire w_dff_A_KdzitkGW9_0;
	wire w_dff_A_lGMJ01SH2_0;
	wire w_dff_A_f7UkhaFr8_0;
	wire w_dff_A_lZrKjVFF9_0;
	wire w_dff_A_Tlk1XYYi2_0;
	wire w_dff_A_dAcs90u54_0;
	wire w_dff_A_9TzEKDLb0_2;
	wire w_dff_A_nLswiUEQ4_0;
	wire w_dff_A_SgXvakfC7_0;
	wire w_dff_A_I04w0Ed15_0;
	wire w_dff_A_iyBw2BMF3_0;
	wire w_dff_A_6ErcL3651_0;
	wire w_dff_A_nuQVfrCK8_0;
	wire w_dff_A_bat33BQT1_1;
	wire w_dff_A_xBVxXj4H3_0;
	wire w_dff_A_Ibvd90Nt5_0;
	wire w_dff_A_BVNvk7AR9_0;
	wire w_dff_A_a03MK4F13_0;
	wire w_dff_A_2mHympoU3_0;
	wire w_dff_A_TFZNP5og8_0;
	wire w_dff_A_hzuSuDqq4_0;
	wire w_dff_A_k9oBrKtw7_0;
	wire w_dff_A_qb8llft07_0;
	wire w_dff_A_KVPLnuKV2_0;
	wire w_dff_A_wz1dhINR5_0;
	wire w_dff_A_ztoZ4Ik43_0;
	wire w_dff_A_AIYD32ue7_0;
	wire w_dff_A_3U8FYw7z2_0;
	wire w_dff_A_xchP7zrc5_0;
	wire w_dff_A_yQncFvPD4_0;
	wire w_dff_A_xa2axSfF4_0;
	wire w_dff_A_v8chX6U61_0;
	wire w_dff_A_840EB0C47_0;
	wire w_dff_A_wd53ojks9_0;
	wire w_dff_A_LO2AdWXo9_0;
	wire w_dff_A_6lDPQMiM6_0;
	wire w_dff_A_58rfLbq44_0;
	wire w_dff_A_GLScgb9d0_0;
	wire w_dff_A_PnGpoDEQ5_0;
	wire w_dff_A_putrv7vJ4_1;
	wire w_dff_A_17DCkZix0_1;
	wire w_dff_A_GGOXVVd55_1;
	wire w_dff_A_2G7GTXXA1_1;
	wire w_dff_A_WmTVgcOY8_1;
	wire w_dff_A_sf7ceMWh8_1;
	wire w_dff_A_uuRuBxWL8_1;
	wire w_dff_A_b7vCj8VR6_1;
	wire w_dff_A_YGd7f3wq6_1;
	wire w_dff_A_woP5CPUj6_1;
	wire w_dff_A_oAwbT1it9_1;
	wire w_dff_A_hFXxqUvB9_1;
	wire w_dff_A_ACcCLzje2_1;
	wire w_dff_A_aPtPo35h4_1;
	wire w_dff_A_3LW8RjDF0_1;
	wire w_dff_A_Zoh4t3ou5_1;
	wire w_dff_A_lv4hDV2y3_1;
	wire w_dff_A_cdXJ55VL2_1;
	wire w_dff_A_7ZANJyQm1_1;
	wire w_dff_A_BYVEcj0V7_1;
	wire w_dff_A_OAKd8djJ0_1;
	wire w_dff_A_uUhV7zC25_1;
	wire w_dff_A_JY1X5m9b9_1;
	wire w_dff_A_AX76BrwG9_2;
	wire w_dff_A_mORhmi6x1_2;
	wire w_dff_A_RIabsRvN7_2;
	wire w_dff_A_BkjMFss80_2;
	wire w_dff_A_fue3WWkf4_2;
	wire w_dff_A_7zXDXjEg5_2;
	wire w_dff_A_44uiDhtB2_2;
	wire w_dff_A_LSu6I9x51_0;
	wire w_dff_A_qpziZNcy2_0;
	wire w_dff_A_iw44Z7qf6_0;
	wire w_dff_A_uUu8MmDp4_0;
	wire w_dff_A_6GlWTpt34_0;
	wire w_dff_A_hWUgsm1k8_0;
	wire w_dff_A_xqQlZuPp8_0;
	wire w_dff_A_vCnhxTSl9_0;
	wire w_dff_A_BbHUDA3K2_0;
	wire w_dff_A_symnjcGt7_0;
	wire w_dff_A_enQQQfPp0_0;
	wire w_dff_A_GkBPbcJL9_0;
	wire w_dff_A_vhNZFhO60_0;
	wire w_dff_A_lHGipaW45_0;
	wire w_dff_A_40KTVuz15_2;
	wire w_dff_A_7i6jMMSp3_0;
	wire w_dff_A_pHMOnJ296_0;
	wire w_dff_A_Y3MK6xy55_0;
	wire w_dff_A_vuklsGmU3_0;
	wire w_dff_A_fRqyKCxj7_0;
	wire w_dff_A_FQ25SIfu6_0;
	wire w_dff_A_dvXEuoOL4_1;
	wire w_dff_A_WXFm6dcW9_0;
	wire w_dff_A_H1Oe7Lxx9_0;
	wire w_dff_A_lIQ7QlUT2_0;
	wire w_dff_A_TU3Lkj7o5_0;
	wire w_dff_A_RQEZTEaR6_0;
	wire w_dff_A_04nxMYQk2_0;
	wire w_dff_A_oSiZ7gDT6_0;
	wire w_dff_A_v169T4Al7_0;
	wire w_dff_A_DjWzpirg1_0;
	wire w_dff_A_Vcwr5R3U8_0;
	wire w_dff_A_RGLphzG85_0;
	wire w_dff_A_zCdpAzNl6_0;
	wire w_dff_A_JKbIRbPS4_0;
	wire w_dff_A_g7v9LeMl6_2;
	wire w_dff_A_rU0gyG9H0_0;
	wire w_dff_A_leS95rAp2_0;
	wire w_dff_A_14drUpLn5_0;
	wire w_dff_A_NCk2KTKr1_0;
	wire w_dff_A_32vJPTt17_0;
	wire w_dff_A_JFAWom510_0;
	wire w_dff_A_ZaaPI5mR8_1;
	wire w_dff_A_y4VQOozV3_0;
	wire w_dff_A_1HbrcX0L3_0;
	wire w_dff_A_18hYKMe90_0;
	wire w_dff_A_led2SLno8_0;
	wire w_dff_A_fnDq3uBZ4_0;
	wire w_dff_A_o9rGKiMQ7_0;
	wire w_dff_A_VJLj8OIH7_0;
	wire w_dff_A_O0q0vL7x6_0;
	wire w_dff_A_pm26wIVv4_0;
	wire w_dff_A_VrOYItL46_0;
	wire w_dff_A_7fkpechI8_0;
	wire w_dff_A_SPyXB4iA3_0;
	wire w_dff_A_FIg2GCjw0_0;
	wire w_dff_A_zygFzT2a9_2;
	wire w_dff_A_6UFmeu6I1_0;
	wire w_dff_A_aqlBCmgJ9_0;
	wire w_dff_A_6z0DgTKQ3_0;
	wire w_dff_A_wYaukfJb9_0;
	wire w_dff_A_A7eitZZH2_1;
	wire w_dff_B_xuLP8Eh94_1;
	wire w_dff_A_bgam7PBe5_0;
	wire w_dff_A_36kQpSaL0_0;
	wire w_dff_A_scUcDVEG6_0;
	wire w_dff_A_YuXhJ4Um4_0;
	wire w_dff_A_N5gcFe2e7_0;
	wire w_dff_A_geBB4Qix9_0;
	wire w_dff_A_Lejslc591_0;
	wire w_dff_A_zHlzfzZr8_0;
	wire w_dff_A_1NvjaUSz2_0;
	wire w_dff_A_qeepUeHI8_0;
	wire w_dff_A_gP9kfPVD8_0;
	wire w_dff_A_zX5oOBHJ6_0;
	wire w_dff_A_OUEB5VwY0_0;
	wire w_dff_A_JTuJefEr1_1;
	wire w_dff_A_Gwj2RSvC4_1;
	wire w_dff_A_j9sEVpXg1_1;
	wire w_dff_A_8CuQWF2Y1_1;
	wire w_dff_A_3klM5Thu5_1;
	wire w_dff_A_wGrMbDhJ8_1;
	wire w_dff_A_7iDJK7nM3_1;
	wire w_dff_A_hFEby3nc2_1;
	wire w_dff_A_rqEwo9jn8_2;
	wire w_dff_A_sZeNBXuB3_0;
	wire w_dff_A_K0G9mO477_0;
	wire w_dff_A_xdj6fnjM7_0;
	wire w_dff_A_B9arFAoA0_0;
	wire w_dff_A_xizCi96C2_0;
	wire w_dff_A_8Lux3dRq9_0;
	wire w_dff_A_1PGOAz6p4_0;
	wire w_dff_A_jfgelKNm7_0;
	wire w_dff_A_v1AH5uDF5_0;
	wire w_dff_A_Xnm3G1324_0;
	wire w_dff_A_hTDcbTfE3_0;
	wire w_dff_A_Vx6xWK0C8_0;
	wire w_dff_A_x36w9jM47_0;
	wire w_dff_A_UTPgT86y3_0;
	wire w_dff_A_7jISbaM68_0;
	wire w_dff_A_fIPF64IO4_0;
	wire w_dff_A_cev2CjdC9_0;
	wire w_dff_A_XGjrlVQB2_0;
	wire w_dff_A_UzbiHO6K5_0;
	wire w_dff_A_yhMk9iiA4_0;
	wire w_dff_A_P4Fkf42Z9_0;
	wire w_dff_A_xttPJG3s4_0;
	wire w_dff_A_xbIUcwZn2_1;
	wire w_dff_A_YfPI2v904_1;
	wire w_dff_A_njh5mEWr0_0;
	wire w_dff_A_oQwh5ee35_0;
	wire w_dff_A_ukaMzAcL2_0;
	wire w_dff_A_hatnZ07Q8_0;
	wire w_dff_A_nBB38dso0_0;
	wire w_dff_A_3DSdJ4Sk0_0;
	wire w_dff_A_HtasaU2e2_0;
	wire w_dff_A_7ldb0iwp0_0;
	wire w_dff_A_u5eVZI6s5_0;
	wire w_dff_A_lBlkwG4Y0_0;
	wire w_dff_A_Et6fxDxo6_0;
	wire w_dff_A_cQJbJjac7_0;
	wire w_dff_A_W91orP1H0_0;
	wire w_dff_A_0wake6Zx2_0;
	wire w_dff_A_WrNNn8z30_0;
	wire w_dff_A_jOKJLA681_0;
	wire w_dff_A_tGJMAIzP5_0;
	wire w_dff_A_T1BD899E4_0;
	wire w_dff_A_vEBV3Mnq0_0;
	wire w_dff_A_GdmBcFZY3_0;
	wire w_dff_A_zslZLxxx2_1;
	wire w_dff_A_fgKGFq3v6_0;
	wire w_dff_A_bCeJejtr7_0;
	wire w_dff_A_YvxgP7e18_0;
	wire w_dff_A_t7G4EAm29_0;
	wire w_dff_A_DsxUjxth7_0;
	wire w_dff_A_othRQFY30_0;
	wire w_dff_A_k0587dBx3_0;
	wire w_dff_A_fyuhdg9T0_0;
	wire w_dff_A_gOXwcJzZ9_0;
	wire w_dff_A_bJyxZgMB5_0;
	wire w_dff_A_iTSAjUzA0_0;
	wire w_dff_A_t8OamHmj4_0;
	wire w_dff_A_PlgHKSDr8_0;
	wire w_dff_A_pATUosgy8_2;
	wire w_dff_A_v8jZ1EzT4_0;
	wire w_dff_A_24bsNqOf1_0;
	wire w_dff_A_ZuZ75MTa6_0;
	wire w_dff_A_cnKnaLTX0_0;
	wire w_dff_A_YvfxF16g4_0;
	wire w_dff_A_Zx3vGH9S5_0;
	wire w_dff_A_U0JIoQ1W4_1;
	wire w_dff_A_ICoZLC8m9_0;
	jnot g000(.din(w_G102gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G108gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G43gat_0[1]),.dout(n45),.clk(gclk));
	jor g003(.dina(w_n45_0[1]),.dinb(w_dff_B_xuLP8Eh94_1),.dout(n46),.clk(gclk));
	jnot g004(.din(w_n46_0[2]),.dout(n47),.clk(gclk));
	jor g005(.dina(w_n47_0[1]),.dinb(w_n44_0[1]),.dout(n48),.clk(gclk));
	jnot g006(.din(w_G63gat_0[2]),.dout(n49),.clk(gclk));
	jand g007(.dina(w_G69gat_0[2]),.dinb(w_n49_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G11gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G17gat_0[2]),.dinb(w_n51_0[1]),.dout(n52),.clk(gclk));
	jor g010(.dina(n52),.dinb(n50),.dout(n53),.clk(gclk));
	jnot g011(.din(w_G24gat_0[2]),.dout(n54),.clk(gclk));
	jand g012(.dina(w_G30gat_0[2]),.dinb(w_n54_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G50gat_0[1]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G56gat_1[1]),.dinb(n56),.dout(n57),.clk(gclk));
	jor g015(.dina(w_n57_0[1]),.dinb(n55),.dout(n58),.clk(gclk));
	jor g016(.dina(n58),.dinb(n53),.dout(n59),.clk(gclk));
	jnot g017(.din(w_G1gat_0[2]),.dout(n60),.clk(gclk));
	jand g018(.dina(w_G4gat_0[2]),.dinb(w_n60_0[1]),.dout(n61),.clk(gclk));
	jnot g019(.din(w_G89gat_0[2]),.dout(n62),.clk(gclk));
	jand g020(.dina(w_G95gat_0[2]),.dinb(w_n62_0[1]),.dout(n63),.clk(gclk));
	jnot g021(.din(w_G76gat_0[2]),.dout(n64),.clk(gclk));
	jand g022(.dina(w_G82gat_0[2]),.dinb(w_n64_0[1]),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n63),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(w_dff_B_rrynMJak1_1),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(n59),.dout(n68),.clk(gclk));
	jor g026(.dina(n68),.dinb(w_dff_B_s0c1Tnw43_1),.dout(G223gat_fa_),.clk(gclk));
	jnot g027(.din(w_G21gat_0[2]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_n44_0[0]),.dout(n71),.clk(gclk));
	jand g029(.dina(w_n46_0[1]),.dinb(n71),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G69gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G63gat_0[1]),.dout(n74),.clk(gclk));
	jnot g032(.din(w_G17gat_0[1]),.dout(n75),.clk(gclk));
	jor g033(.dina(w_n75_0[1]),.dinb(w_G11gat_0[1]),.dout(n76),.clk(gclk));
	jand g034(.dina(n76),.dinb(n74),.dout(n77),.clk(gclk));
	jnot g035(.din(w_G30gat_0[1]),.dout(n78),.clk(gclk));
	jor g036(.dina(w_n78_0[1]),.dinb(w_G24gat_0[1]),.dout(n79),.clk(gclk));
	jnot g037(.din(w_G56gat_1[0]),.dout(n80),.clk(gclk));
	jor g038(.dina(w_n80_0[1]),.dinb(w_G50gat_0[0]),.dout(n81),.clk(gclk));
	jand g039(.dina(w_n81_0[1]),.dinb(n79),.dout(n82),.clk(gclk));
	jand g040(.dina(n82),.dinb(n77),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G4gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G1gat_0[1]),.dout(n85),.clk(gclk));
	jnot g043(.din(w_G95gat_0[1]),.dout(n86),.clk(gclk));
	jor g044(.dina(w_n86_0[1]),.dinb(w_G89gat_0[1]),.dout(n87),.clk(gclk));
	jnot g045(.din(w_G82gat_0[1]),.dout(n88),.clk(gclk));
	jor g046(.dina(w_n88_0[1]),.dinb(w_G76gat_0[1]),.dout(n89),.clk(gclk));
	jand g047(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(w_dff_B_vtrJgknM1_1),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n83),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(w_dff_B_FXFeITBu7_1),.dout(n93),.clk(gclk));
	jor g051(.dina(w_n93_3[2]),.dinb(w_n51_0[0]),.dout(n94),.clk(gclk));
	jand g052(.dina(n94),.dinb(w_G17gat_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(w_n95_0[1]),.dinb(w_n70_0[1]),.dout(n96),.clk(gclk));
	jnot g054(.din(w_G99gat_0[2]),.dout(n97),.clk(gclk));
	jor g055(.dina(w_n93_3[1]),.dinb(w_n62_0[0]),.dout(n98),.clk(gclk));
	jand g056(.dina(n98),.dinb(w_G95gat_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(w_dff_B_69IWdBfv7_1),.dout(n100),.clk(gclk));
	jor g058(.dina(n100),.dinb(n96),.dout(n101),.clk(gclk));
	jnot g059(.din(w_G73gat_0[2]),.dout(n102),.clk(gclk));
	jor g060(.dina(w_n93_3[0]),.dinb(w_n49_0[0]),.dout(n103),.clk(gclk));
	jand g061(.dina(n103),.dinb(w_G69gat_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(w_n104_0[1]),.dinb(w_n102_0[1]),.dout(n105),.clk(gclk));
	jnot g063(.din(w_G34gat_0[2]),.dout(n106),.clk(gclk));
	jor g064(.dina(w_n93_2[2]),.dinb(w_n54_0[0]),.dout(n107),.clk(gclk));
	jand g065(.dina(n107),.dinb(w_G30gat_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(w_n108_0[1]),.dinb(w_n106_0[1]),.dout(n109),.clk(gclk));
	jor g067(.dina(n109),.dinb(n105),.dout(n110),.clk(gclk));
	jnot g068(.din(w_G112gat_0[2]),.dout(n111),.clk(gclk));
	jor g069(.dina(w_n93_2[1]),.dinb(w_n43_0[0]),.dout(n112),.clk(gclk));
	jand g070(.dina(n112),.dinb(w_G108gat_0[1]),.dout(n113),.clk(gclk));
	jand g071(.dina(w_n113_0[1]),.dinb(w_n111_0[1]),.dout(n114),.clk(gclk));
	jor g072(.dina(w_dff_B_5jEXFLQw6_0),.dinb(n110),.dout(n115),.clk(gclk));
	jor g073(.dina(n115),.dinb(w_dff_B_UuWpBk8e4_1),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[1]),.dout(n117),.clk(gclk));
	jxor g075(.dina(w_n93_2[0]),.dinb(w_n57_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[2]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[2]),.dinb(w_n117_0[1]),.dout(n120),.clk(gclk));
	jnot g078(.din(w_G86gat_0[2]),.dout(n121),.clk(gclk));
	jor g079(.dina(w_n93_1[2]),.dinb(w_n64_0[0]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G82gat_0[0]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jnot g082(.din(w_G8gat_0[2]),.dout(n125),.clk(gclk));
	jor g083(.dina(w_n93_1[1]),.dinb(w_n60_0[0]),.dout(n126),.clk(gclk));
	jand g084(.dina(n126),.dinb(w_G4gat_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(w_n127_0[1]),.dinb(w_n125_0[1]),.dout(n128),.clk(gclk));
	jnot g086(.din(w_G47gat_0[2]),.dout(n129),.clk(gclk));
	jor g087(.dina(w_n93_1[0]),.dinb(w_n47_0[0]),.dout(n130),.clk(gclk));
	jand g088(.dina(n130),.dinb(w_G43gat_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(w_n131_0[2]),.dinb(w_dff_B_JB9geFc13_1),.dout(n132),.clk(gclk));
	jor g090(.dina(n132),.dinb(n128),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(w_dff_B_9Ejn8SAM9_1),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(w_n120_0[1]),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(n116),.dout(G329gat_fa_),.clk(gclk));
	jand g094(.dina(w_G223gat_4),.dinb(w_G89gat_0[0]),.dout(n137),.clk(gclk));
	jor g095(.dina(n137),.dinb(w_n86_0[0]),.dout(n138),.clk(gclk));
	jand g096(.dina(w_G329gat_4),.dinb(w_G99gat_0[1]),.dout(n139),.clk(gclk));
	jor g097(.dina(n139),.dinb(w_n138_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(w_n140_0[1]),.dinb(w_G105gat_0[1]),.dout(n141),.clk(gclk));
	jnot g099(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jand g100(.dina(w_G329gat_3[2]),.dinb(w_G47gat_0[1]),.dout(n143),.clk(gclk));
	jnot g101(.din(n143),.dout(n144),.clk(gclk));
	jnot g102(.din(w_G53gat_0[1]),.dout(n145),.clk(gclk));
	jand g103(.dina(w_n131_0[1]),.dinb(w_n145_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_dff_B_paiVXyJb5_0),.dinb(w_n144_0[1]),.dout(n147),.clk(gclk));
	jor g105(.dina(w_n147_0[1]),.dinb(n142),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G40gat_0[1]),.dout(n149),.clk(gclk));
	jand g107(.dina(w_G223gat_3[2]),.dinb(w_G11gat_0[0]),.dout(n150),.clk(gclk));
	jor g108(.dina(n150),.dinb(w_n75_0[0]),.dout(n151),.clk(gclk));
	jor g109(.dina(w_n151_0[1]),.dinb(w_G21gat_0[1]),.dout(n152),.clk(gclk));
	jor g110(.dina(w_n138_0[0]),.dinb(w_G99gat_0[0]),.dout(n153),.clk(gclk));
	jand g111(.dina(n153),.dinb(n152),.dout(n154),.clk(gclk));
	jand g112(.dina(w_G223gat_3[1]),.dinb(w_G63gat_0[0]),.dout(n155),.clk(gclk));
	jor g113(.dina(n155),.dinb(w_n73_0[0]),.dout(n156),.clk(gclk));
	jor g114(.dina(w_n156_0[1]),.dinb(w_G73gat_0[1]),.dout(n157),.clk(gclk));
	jand g115(.dina(w_G223gat_3[0]),.dinb(w_G24gat_0[0]),.dout(n158),.clk(gclk));
	jor g116(.dina(n158),.dinb(w_n78_0[0]),.dout(n159),.clk(gclk));
	jor g117(.dina(w_n159_0[1]),.dinb(w_G34gat_0[1]),.dout(n160),.clk(gclk));
	jand g118(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jnot g119(.din(w_G108gat_0[0]),.dout(n162),.clk(gclk));
	jand g120(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n163),.clk(gclk));
	jor g121(.dina(n163),.dinb(w_dff_B_BOWiELq69_1),.dout(n164),.clk(gclk));
	jor g122(.dina(w_n164_0[1]),.dinb(w_G112gat_0[1]),.dout(n165),.clk(gclk));
	jand g123(.dina(w_dff_B_LS2NnnOg9_0),.dinb(n161),.dout(n166),.clk(gclk));
	jand g124(.dina(n166),.dinb(w_dff_B_L4jdTIV36_1),.dout(n167),.clk(gclk));
	jnot g125(.din(w_n120_0[0]),.dout(n168),.clk(gclk));
	jand g126(.dina(w_G223gat_2[1]),.dinb(w_G76gat_0[0]),.dout(n169),.clk(gclk));
	jor g127(.dina(n169),.dinb(w_n88_0[0]),.dout(n170),.clk(gclk));
	jor g128(.dina(w_n170_0[1]),.dinb(w_G86gat_0[1]),.dout(n171),.clk(gclk));
	jand g129(.dina(w_G223gat_2[0]),.dinb(w_G1gat_0[0]),.dout(n172),.clk(gclk));
	jor g130(.dina(n172),.dinb(w_n84_0[0]),.dout(n173),.clk(gclk));
	jor g131(.dina(w_n173_0[1]),.dinb(w_G8gat_0[1]),.dout(n174),.clk(gclk));
	jand g132(.dina(w_G223gat_1[2]),.dinb(w_n46_0[0]),.dout(n175),.clk(gclk));
	jor g133(.dina(n175),.dinb(w_n45_0[0]),.dout(n176),.clk(gclk));
	jor g134(.dina(n176),.dinb(w_G47gat_0[0]),.dout(n177),.clk(gclk));
	jand g135(.dina(n177),.dinb(n174),.dout(n178),.clk(gclk));
	jand g136(.dina(n178),.dinb(w_dff_B_xhPinsnU9_1),.dout(n179),.clk(gclk));
	jand g137(.dina(n179),.dinb(w_dff_B_SDhLMKyS7_1),.dout(n180),.clk(gclk));
	jand g138(.dina(n180),.dinb(n167),.dout(n181),.clk(gclk));
	jor g139(.dina(w_n181_2[2]),.dinb(w_n106_0[0]),.dout(n182),.clk(gclk));
	jand g140(.dina(n182),.dinb(w_n108_0[0]),.dout(n183),.clk(gclk));
	jand g141(.dina(w_n183_0[1]),.dinb(w_n149_0[1]),.dout(n184),.clk(gclk));
	jnot g142(.din(w_G66gat_0[2]),.dout(n185),.clk(gclk));
	jor g143(.dina(w_n181_2[1]),.dinb(w_n117_0[0]),.dout(n186),.clk(gclk));
	jand g144(.dina(n186),.dinb(w_n119_0[1]),.dout(n187),.clk(gclk));
	jand g145(.dina(n187),.dinb(w_n185_0[1]),.dout(n188),.clk(gclk));
	jor g146(.dina(n188),.dinb(n184),.dout(n189),.clk(gclk));
	jnot g147(.din(w_G14gat_0[2]),.dout(n190),.clk(gclk));
	jor g148(.dina(w_n181_2[0]),.dinb(w_n125_0[0]),.dout(n191),.clk(gclk));
	jand g149(.dina(n191),.dinb(w_n127_0[0]),.dout(n192),.clk(gclk));
	jand g150(.dina(n192),.dinb(w_dff_B_1ab0SRD63_1),.dout(n193),.clk(gclk));
	jnot g151(.din(w_G92gat_0[2]),.dout(n194),.clk(gclk));
	jor g152(.dina(w_n181_1[2]),.dinb(w_n121_0[0]),.dout(n195),.clk(gclk));
	jand g153(.dina(n195),.dinb(w_n123_0[0]),.dout(n196),.clk(gclk));
	jand g154(.dina(n196),.dinb(w_dff_B_V6kzopNN6_1),.dout(n197),.clk(gclk));
	jor g155(.dina(n197),.dinb(n193),.dout(n198),.clk(gclk));
	jor g156(.dina(n198),.dinb(n189),.dout(n199),.clk(gclk));
	jnot g157(.din(w_G79gat_0[1]),.dout(n200),.clk(gclk));
	jor g158(.dina(w_n181_1[1]),.dinb(w_n102_0[0]),.dout(n201),.clk(gclk));
	jand g159(.dina(n201),.dinb(w_n104_0[0]),.dout(n202),.clk(gclk));
	jand g160(.dina(w_n202_0[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jnot g161(.din(w_G115gat_0[1]),.dout(n204),.clk(gclk));
	jor g162(.dina(w_n181_1[0]),.dinb(w_n111_0[0]),.dout(n205),.clk(gclk));
	jand g163(.dina(n205),.dinb(w_n113_0[0]),.dout(n206),.clk(gclk));
	jand g164(.dina(w_n206_0[1]),.dinb(w_n204_0[1]),.dout(n207),.clk(gclk));
	jor g165(.dina(n207),.dinb(n203),.dout(n208),.clk(gclk));
	jnot g166(.din(w_G27gat_0[1]),.dout(n209),.clk(gclk));
	jor g167(.dina(w_n181_0[2]),.dinb(w_n70_0[0]),.dout(n210),.clk(gclk));
	jand g168(.dina(n210),.dinb(w_n95_0[0]),.dout(n211),.clk(gclk));
	jand g169(.dina(w_n211_0[1]),.dinb(w_n209_0[1]),.dout(n212),.clk(gclk));
	jor g170(.dina(w_dff_B_qSKNWnMq2_0),.dinb(n208),.dout(n213),.clk(gclk));
	jor g171(.dina(n213),.dinb(n199),.dout(n214),.clk(gclk));
	jor g172(.dina(n214),.dinb(w_dff_B_YYPEZ8R58_1),.dout(G370gat_fa_),.clk(gclk));
	jnot g173(.din(w_n147_0[0]),.dout(n216),.clk(gclk));
	jand g174(.dina(n216),.dinb(w_n141_0[0]),.dout(n217),.clk(gclk));
	jand g175(.dina(w_G329gat_3[1]),.dinb(w_G34gat_0[0]),.dout(n218),.clk(gclk));
	jor g176(.dina(n218),.dinb(w_n159_0[0]),.dout(n219),.clk(gclk));
	jor g177(.dina(n219),.dinb(w_G40gat_0[0]),.dout(n220),.clk(gclk));
	jnot g178(.din(w_n119_0[0]),.dout(n221),.clk(gclk));
	jand g179(.dina(w_G329gat_3[0]),.dinb(w_G60gat_0[0]),.dout(n222),.clk(gclk));
	jor g180(.dina(w_n222_0[1]),.dinb(w_dff_B_0zhaWSMg6_1),.dout(n223),.clk(gclk));
	jor g181(.dina(n223),.dinb(w_G66gat_0[1]),.dout(n224),.clk(gclk));
	jand g182(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jand g183(.dina(w_G329gat_2[2]),.dinb(w_G8gat_0[0]),.dout(n226),.clk(gclk));
	jor g184(.dina(n226),.dinb(w_n173_0[0]),.dout(n227),.clk(gclk));
	jor g185(.dina(w_n227_0[1]),.dinb(w_G14gat_0[1]),.dout(n228),.clk(gclk));
	jand g186(.dina(w_G329gat_2[1]),.dinb(w_G86gat_0[0]),.dout(n229),.clk(gclk));
	jor g187(.dina(n229),.dinb(w_n170_0[0]),.dout(n230),.clk(gclk));
	jor g188(.dina(w_n230_0[1]),.dinb(w_G92gat_0[1]),.dout(n231),.clk(gclk));
	jand g189(.dina(n231),.dinb(n228),.dout(n232),.clk(gclk));
	jand g190(.dina(n232),.dinb(n225),.dout(n233),.clk(gclk));
	jand g191(.dina(w_G329gat_2[0]),.dinb(w_G73gat_0[0]),.dout(n234),.clk(gclk));
	jor g192(.dina(n234),.dinb(w_n156_0[0]),.dout(n235),.clk(gclk));
	jor g193(.dina(n235),.dinb(w_G79gat_0[0]),.dout(n236),.clk(gclk));
	jand g194(.dina(w_G329gat_1[2]),.dinb(w_G112gat_0[0]),.dout(n237),.clk(gclk));
	jor g195(.dina(n237),.dinb(w_n164_0[0]),.dout(n238),.clk(gclk));
	jor g196(.dina(n238),.dinb(w_G115gat_0[0]),.dout(n239),.clk(gclk));
	jand g197(.dina(n239),.dinb(n236),.dout(n240),.clk(gclk));
	jand g198(.dina(w_G329gat_1[1]),.dinb(w_G21gat_0[0]),.dout(n241),.clk(gclk));
	jor g199(.dina(n241),.dinb(w_n151_0[0]),.dout(n242),.clk(gclk));
	jor g200(.dina(n242),.dinb(w_G27gat_0[0]),.dout(n243),.clk(gclk));
	jand g201(.dina(w_dff_B_B7W15AHw3_0),.dinb(n240),.dout(n244),.clk(gclk));
	jand g202(.dina(n244),.dinb(n233),.dout(n245),.clk(gclk));
	jand g203(.dina(n245),.dinb(w_dff_B_LR9dAh5R7_1),.dout(n246),.clk(gclk));
	jor g204(.dina(w_n246_2[2]),.dinb(w_n209_0[0]),.dout(n247),.clk(gclk));
	jand g205(.dina(n247),.dinb(w_n211_0[0]),.dout(n248),.clk(gclk));
	jor g206(.dina(w_n246_2[1]),.dinb(w_n149_0[0]),.dout(n249),.clk(gclk));
	jand g207(.dina(n249),.dinb(w_n183_0[0]),.dout(n250),.clk(gclk));
	jor g208(.dina(w_n250_0[1]),.dinb(w_n248_0[1]),.dout(n251),.clk(gclk));
	jor g209(.dina(w_n246_2[0]),.dinb(w_n145_0[0]),.dout(n252),.clk(gclk));
	jand g210(.dina(w_n144_0[0]),.dinb(w_n131_0[0]),.dout(n253),.clk(gclk));
	jand g211(.dina(w_n253_0[1]),.dinb(n252),.dout(n254),.clk(gclk));
	jor g212(.dina(w_n246_1[2]),.dinb(w_n185_0[0]),.dout(n255),.clk(gclk));
	jand g213(.dina(w_G223gat_1[1]),.dinb(w_n81_0[0]),.dout(n256),.clk(gclk));
	jor g214(.dina(w_n222_0[0]),.dinb(w_dff_B_sm8nqeof3_1),.dout(n257),.clk(gclk));
	jnot g215(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g216(.dina(w_dff_B_haira9qa2_0),.dinb(n255),.dout(n259),.clk(gclk));
	jand g217(.dina(n259),.dinb(w_G56gat_0[1]),.dout(n260),.clk(gclk));
	jor g218(.dina(n260),.dinb(w_n254_0[1]),.dout(n261),.clk(gclk));
	jor g219(.dina(n261),.dinb(w_n251_0[1]),.dout(G430gat_fa_),.clk(gclk));
	jand g220(.dina(w_G370gat_1[1]),.dinb(w_G92gat_0[0]),.dout(n263),.clk(gclk));
	jor g221(.dina(n263),.dinb(w_n230_0[0]),.dout(n264),.clk(gclk));
	jnot g222(.din(w_n264_0[1]),.dout(n265),.clk(gclk));
	jnot g223(.din(w_n140_0[0]),.dout(n266),.clk(gclk));
	jnot g224(.din(w_G105gat_0[0]),.dout(n267),.clk(gclk));
	jor g225(.dina(w_n246_1[1]),.dinb(w_dff_B_sWI2zR2Z2_1),.dout(n268),.clk(gclk));
	jand g226(.dina(n268),.dinb(w_dff_B_4YKhSSsa8_1),.dout(n269),.clk(gclk));
	jor g227(.dina(w_n246_1[0]),.dinb(w_n200_0[0]),.dout(n270),.clk(gclk));
	jand g228(.dina(n270),.dinb(w_n202_0[0]),.dout(n271),.clk(gclk));
	jor g229(.dina(w_n246_0[2]),.dinb(w_n204_0[0]),.dout(n272),.clk(gclk));
	jand g230(.dina(n272),.dinb(w_n206_0[0]),.dout(n273),.clk(gclk));
	jor g231(.dina(n273),.dinb(w_n271_0[1]),.dout(n274),.clk(gclk));
	jor g232(.dina(n274),.dinb(w_n269_0[1]),.dout(n275),.clk(gclk));
	jor g233(.dina(n275),.dinb(w_n265_0[1]),.dout(n276),.clk(gclk));
	jor g234(.dina(n276),.dinb(w_G430gat_0),.dout(n277),.clk(gclk));
	jand g235(.dina(w_G370gat_1[0]),.dinb(w_G14gat_0[0]),.dout(n278),.clk(gclk));
	jor g236(.dina(n278),.dinb(w_n227_0[0]),.dout(n279),.clk(gclk));
	jand g237(.dina(w_dff_B_mm8gENSW7_0),.dinb(n277),.dout(G421gat),.clk(gclk));
	jnot g238(.din(w_n250_0[0]),.dout(n281),.clk(gclk));
	jand g239(.dina(w_G370gat_0[2]),.dinb(w_G53gat_0[0]),.dout(n282),.clk(gclk));
	jnot g240(.din(w_n253_0[0]),.dout(n283),.clk(gclk));
	jor g241(.dina(w_dff_B_Ia4EvD1F4_0),.dinb(n282),.dout(n284),.clk(gclk));
	jand g242(.dina(w_G370gat_0[1]),.dinb(w_G66gat_0[0]),.dout(n285),.clk(gclk));
	jor g243(.dina(w_n257_0[0]),.dinb(n285),.dout(n286),.clk(gclk));
	jor g244(.dina(n286),.dinb(w_n80_0[0]),.dout(n287),.clk(gclk));
	jand g245(.dina(n287),.dinb(w_dff_B_T4nIGQqQ2_1),.dout(n288),.clk(gclk));
	jand g246(.dina(w_n288_0[1]),.dinb(w_n281_0[1]),.dout(n289),.clk(gclk));
	jand g247(.dina(n289),.dinb(w_n271_0[0]),.dout(n290),.clk(gclk));
	jand g248(.dina(w_n265_0[0]),.dinb(w_n288_0[0]),.dout(n291),.clk(gclk));
	jor g249(.dina(n291),.dinb(w_n251_0[0]),.dout(n292),.clk(gclk));
	jor g250(.dina(n292),.dinb(w_n290_0[1]),.dout(G431gat),.clk(gclk));
	jand g251(.dina(w_n269_0[0]),.dinb(w_n264_0[0]),.dout(n294),.clk(gclk));
	jor g252(.dina(n294),.dinb(w_n254_0[0]),.dout(n295),.clk(gclk));
	jand g253(.dina(n295),.dinb(w_n281_0[0]),.dout(n296),.clk(gclk));
	jor g254(.dina(n296),.dinb(w_n248_0[0]),.dout(n297),.clk(gclk));
	jor g255(.dina(n297),.dinb(w_n290_0[0]),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_nuQVfrCK8_0),.doutb(w_dff_A_bat33BQT1_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_dAcs90u54_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_9TzEKDLb0_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_22AEj7LU2_0),.doutb(w_dff_A_jKSTLNsP8_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_dff_A_JFAWom510_0),.doutb(w_dff_A_ZaaPI5mR8_1),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_dff_A_B9LX9zz21_0),.doutb(w_dff_A_iA559QVq3_1),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_dff_A_JKbIRbPS4_0),.doutb(w_G17gat_0[1]),.doutc(w_dff_A_g7v9LeMl6_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_dff_A_dHsrHFZ11_0),.doutb(w_dff_A_gpuN8SLz2_1),.doutc(w_G21gat_0[2]),.din(G21gat));
	jspl3 jspl3_w_G24gat_0(.douta(w_dff_A_FQ25SIfu6_0),.doutb(w_dff_A_dvXEuoOL4_1),.doutc(w_G24gat_0[2]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_dff_A_t1lvHTWN3_0),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl3 jspl3_w_G30gat_0(.douta(w_dff_A_lHGipaW45_0),.doutb(w_G30gat_0[1]),.doutc(w_dff_A_40KTVuz15_2),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_TtTMic2f7_0),.doutb(w_dff_A_0qqjJV1q4_1),.doutc(w_G34gat_0[2]),.din(G34gat));
	jspl jspl_w_G40gat_0(.douta(w_dff_A_S9Y8jeJ59_0),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl jspl_w_G43gat_0(.douta(w_dff_A_OUEB5VwY0_0),.doutb(w_G43gat_0[1]),.din(G43gat));
	jspl3 jspl3_w_G47gat_0(.douta(w_dff_A_PNAk39HP3_0),.doutb(w_dff_A_wKWGJvJL1_1),.doutc(w_G47gat_0[2]),.din(G47gat));
	jspl jspl_w_G50gat_0(.douta(w_dff_A_LSu6I9x51_0),.doutb(w_G50gat_0[1]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_nWrydaZy0_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_G56gat_0[0]),.doutb(w_dff_A_JY1X5m9b9_1),.doutc(w_dff_A_44uiDhtB2_2),.din(G56gat));
	jspl jspl_w_G56gat_1(.douta(w_G56gat_1[0]),.doutb(w_dff_A_putrv7vJ4_1),.din(w_G56gat_0[0]));
	jspl jspl_w_G60gat_0(.douta(w_dff_A_YG8qQCjJ1_0),.doutb(w_G60gat_0[1]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_dff_A_xttPJG3s4_0),.doutb(w_dff_A_xbIUcwZn2_1),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl3 jspl3_w_G66gat_0(.douta(w_dff_A_40SG9CPg4_0),.doutb(w_dff_A_0ARvSZ8F9_1),.doutc(w_G66gat_0[2]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_FIg2GCjw0_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_zygFzT2a9_2),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_dff_A_oOw3wfMq8_0),.doutb(w_dff_A_mkmU92eL9_1),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl3 jspl3_w_G76gat_0(.douta(w_dff_A_m0axmQEX1_0),.doutb(w_dff_A_SDsstCuO9_1),.doutc(w_G76gat_0[2]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_dff_A_4Hbif21O6_0),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_dff_A_8NwcASrU2_0),.doutb(w_G82gat_0[1]),.doutc(w_dff_A_QxQf8HVV3_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_dff_A_a8rZTlo97_0),.doutb(w_dff_A_e7w7KJmh4_1),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_5c5qQ5998_0),.doutb(w_dff_A_jsSRzS613_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_sHVhMF8S9_0),.doutb(w_dff_A_YT8iWFLb1_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_s6eqjM6c5_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_EYXFSrfy1_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_HWIp2MDX0_0),.doutb(w_dff_A_9Sv5mRmP8_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl jspl_w_G102gat_0(.douta(w_dff_A_hTDcbTfE3_0),.doutb(w_G102gat_0[1]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_H0izGr0v9_1),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_G108gat_0[0]),.doutb(w_dff_A_hFEby3nc2_1),.doutc(w_dff_A_rqEwo9jn8_2),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_dff_A_Trkf7w596_0),.doutb(w_dff_A_vSKhQeS71_1),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_dff_A_BrB88TYv0_0),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_G223gat_3[2]),.din(w_G223gat_0[2]));
	jspl jspl_w_G223gat_4(.douta(w_G223gat_4),.doutb(w_dff_A_YfPI2v904_1),.din(w_G223gat_1[0]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl jspl_w_G329gat_4(.douta(w_G329gat_4),.doutb(w_dff_A_zslZLxxx2_1),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_dff_A_pATUosgy8_2),.din(w_G370gat_0[0]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_U0JIoQ1W4_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_dff_A_xizCi96C2_0),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_dff_A_JTuJefEr1_1),.din(n44));
	jspl jspl_w_n45_0(.douta(w_dff_A_geBB4Qix9_0),.doutb(w_n45_0[1]),.din(n45));
	jspl3 jspl3_w_n46_0(.douta(w_dff_A_wYaukfJb9_0),.doutb(w_dff_A_A7eitZZH2_1),.doutc(w_n46_0[2]),.din(n46));
	jspl jspl_w_n47_0(.douta(w_dff_A_Fe8ugEQt2_0),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n49_0(.douta(w_dff_A_fIPF64IO4_0),.doutb(w_n49_0[1]),.din(n49));
	jspl jspl_w_n51_0(.douta(w_dff_A_L2s6nSm88_0),.doutb(w_n51_0[1]),.din(n51));
	jspl jspl_w_n54_0(.douta(w_dff_A_oqnyvqRT4_0),.doutb(w_n54_0[1]),.din(n54));
	jspl jspl_w_n57_0(.douta(w_dff_A_EghAq9VE0_0),.doutb(w_n57_0[1]),.din(n57));
	jspl jspl_w_n60_0(.douta(w_dff_A_BXhbeJ6u9_0),.doutb(w_n60_0[1]),.din(n60));
	jspl jspl_w_n62_0(.douta(w_dff_A_w2p70dmt4_0),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n64_0(.douta(w_dff_A_7n9LOtu14_0),.doutb(w_n64_0[1]),.din(n64));
	jspl jspl_w_n70_0(.douta(w_dff_A_Vpuez0BJ8_0),.doutb(w_n70_0[1]),.din(w_dff_B_zXMf2XEi9_2));
	jspl jspl_w_n73_0(.douta(w_dff_A_o9rGKiMQ7_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n75_0(.douta(w_dff_A_04nxMYQk2_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n78_0(.douta(w_dff_A_xqQlZuPp8_0),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n80_0(.douta(w_dff_A_PnGpoDEQ5_0),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n81_0(.douta(w_dff_A_a03MK4F13_0),.doutb(w_n81_0[1]),.din(n81));
	jspl jspl_w_n84_0(.douta(w_dff_A_jJ4botKv4_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_69aeXXNp3_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_dff_A_EhqGlHxz9_0),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl3 jspl3_w_n93_1(.douta(w_n93_1[0]),.doutb(w_n93_1[1]),.doutc(w_n93_1[2]),.din(w_n93_0[0]));
	jspl3 jspl3_w_n93_2(.douta(w_n93_2[0]),.doutb(w_n93_2[1]),.doutc(w_n93_2[2]),.din(w_n93_0[1]));
	jspl3 jspl3_w_n93_3(.douta(w_n93_3[0]),.doutb(w_n93_3[1]),.doutc(w_n93_3[2]),.din(w_n93_0[2]));
	jspl jspl_w_n95_0(.douta(w_dff_A_zIBHdoei7_0),.doutb(w_n95_0[1]),.din(n95));
	jspl jspl_w_n102_0(.douta(w_dff_A_Up8MHMLe2_0),.doutb(w_n102_0[1]),.din(w_dff_B_4eM6QmVo7_2));
	jspl jspl_w_n104_0(.douta(w_dff_A_zxeppp4M2_0),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_dff_A_iVbpCoSB7_0),.doutb(w_n106_0[1]),.din(w_dff_B_xZXqVwxy2_2));
	jspl jspl_w_n108_0(.douta(w_dff_A_HfQCzGGO4_0),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n111_0(.douta(w_dff_A_SlqBgjwD3_0),.doutb(w_n111_0[1]),.din(w_dff_B_d94g1jne5_2));
	jspl jspl_w_n113_0(.douta(w_dff_A_dZUWnc8V7_0),.doutb(w_n113_0[1]),.din(n113));
	jspl jspl_w_n117_0(.douta(w_dff_A_6OkFu1Y69_0),.doutb(w_n117_0[1]),.din(w_dff_B_6F2pPsVZ8_2));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_dff_A_q34n06QX0_1),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_dff_A_bNchDfR86_1),.din(n120));
	jspl jspl_w_n121_0(.douta(w_dff_A_ZZTgA83A1_0),.doutb(w_n121_0[1]),.din(w_dff_B_2383nTjN5_2));
	jspl jspl_w_n123_0(.douta(w_dff_A_iXLtYgTW0_0),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_dff_A_8KnHbGtN8_0),.doutb(w_n125_0[1]),.din(w_dff_B_LjiddWGy7_2));
	jspl jspl_w_n127_0(.douta(w_dff_A_ulPa3Dcx5_0),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n131_0(.douta(w_dff_A_xlMAHoDw3_0),.doutb(w_n131_0[1]),.doutc(w_n131_0[2]),.din(n131));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_dff_A_D620hIjN3_1),.din(n138));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_i11qy3oI3_0),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(n144));
	jspl jspl_w_n145_0(.douta(w_dff_A_O0wQlBzA7_0),.doutb(w_n145_0[1]),.din(w_dff_B_nRqDZMM19_2));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_2nMf8lIr9_1),.din(n147));
	jspl jspl_w_n149_0(.douta(w_dff_A_xQpPy1Km9_0),.doutb(w_n149_0[1]),.din(w_dff_B_Ao6Eg4Y10_2));
	jspl jspl_w_n151_0(.douta(w_dff_A_DnJVo4kj9_0),.doutb(w_n151_0[1]),.din(n151));
	jspl jspl_w_n156_0(.douta(w_dff_A_VGxBzT6Y2_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_xrX8NtgM4_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_0nTKHlM67_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_RIKbZ0pK9_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_dff_A_I1Wv4zCs2_0),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n183_0(.douta(w_dff_A_npMJPdxG5_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n185_0(.douta(w_dff_A_KfpRo5LZ4_0),.doutb(w_n185_0[1]),.din(w_dff_B_8zFPGK4q8_2));
	jspl jspl_w_n200_0(.douta(w_dff_A_QSBh61bw9_0),.doutb(w_n200_0[1]),.din(w_dff_B_zxrmMO796_2));
	jspl jspl_w_n202_0(.douta(w_dff_A_sH5qWaTd4_0),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n204_0(.douta(w_dff_A_FkjMFXXK7_0),.doutb(w_n204_0[1]),.din(w_dff_B_11kHvXQO6_2));
	jspl jspl_w_n206_0(.douta(w_dff_A_xvjiRNkU4_0),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n209_0(.douta(w_dff_A_1IQXxtG49_0),.doutb(w_n209_0[1]),.din(w_dff_B_ZpqHa7210_2));
	jspl jspl_w_n211_0(.douta(w_dff_A_RLkBIp1p8_0),.doutb(w_n211_0[1]),.din(n211));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n227_0(.douta(w_dff_A_URiQhGSh9_0),.doutb(w_n227_0[1]),.din(n227));
	jspl jspl_w_n230_0(.douta(w_dff_A_MYdu8TrK4_0),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl3 jspl3_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.doutc(w_n246_1[2]),.din(w_n246_0[0]));
	jspl3 jspl3_w_n246_2(.douta(w_n246_2[0]),.doutb(w_n246_2[1]),.doutc(w_n246_2[2]),.din(w_n246_0[1]));
	jspl jspl_w_n248_0(.douta(w_dff_A_sQdHh1n37_0),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_dff_A_ecMX45fI9_0),.doutb(w_n251_0[1]),.din(w_dff_B_3lorr8c26_2));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_dff_A_clcYDvzU5_1),.din(n253));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_L6dqpViB0_2));
	jspl jspl_w_n257_0(.douta(w_dff_A_K4aNRt418_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(w_dff_B_Xk0lJJfU6_2));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_dff_A_5PGDgAJZ2_1),.din(n269));
	jspl jspl_w_n271_0(.douta(w_dff_A_re46KwVH6_0),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.din(w_dff_B_Dxuofd8Z2_2));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(n290));
	jdff dff_B_bPjHBH3h8_0(.din(n279),.dout(w_dff_B_bPjHBH3h8_0),.clk(gclk));
	jdff dff_B_yl2terfh9_0(.din(w_dff_B_bPjHBH3h8_0),.dout(w_dff_B_yl2terfh9_0),.clk(gclk));
	jdff dff_B_nMZ6D5Dx3_0(.din(w_dff_B_yl2terfh9_0),.dout(w_dff_B_nMZ6D5Dx3_0),.clk(gclk));
	jdff dff_B_mm8gENSW7_0(.din(w_dff_B_nMZ6D5Dx3_0),.dout(w_dff_B_mm8gENSW7_0),.clk(gclk));
	jdff dff_B_VtDiiVvS3_0(.din(n258),.dout(w_dff_B_VtDiiVvS3_0),.clk(gclk));
	jdff dff_B_QyI9FYcT2_0(.din(w_dff_B_VtDiiVvS3_0),.dout(w_dff_B_QyI9FYcT2_0),.clk(gclk));
	jdff dff_B_UDYFs09n4_0(.din(w_dff_B_QyI9FYcT2_0),.dout(w_dff_B_UDYFs09n4_0),.clk(gclk));
	jdff dff_B_6cLSZGCT2_0(.din(w_dff_B_UDYFs09n4_0),.dout(w_dff_B_6cLSZGCT2_0),.clk(gclk));
	jdff dff_B_haira9qa2_0(.din(w_dff_B_6cLSZGCT2_0),.dout(w_dff_B_haira9qa2_0),.clk(gclk));
	jdff dff_B_Xk0lJJfU6_2(.din(n265),.dout(w_dff_B_Xk0lJJfU6_2),.clk(gclk));
	jdff dff_A_ecMX45fI9_0(.dout(w_n251_0[0]),.din(w_dff_A_ecMX45fI9_0),.clk(gclk));
	jdff dff_B_3lorr8c26_2(.din(n251),.dout(w_dff_B_3lorr8c26_2),.clk(gclk));
	jdff dff_A_5PGDgAJZ2_1(.dout(w_n269_0[1]),.din(w_dff_A_5PGDgAJZ2_1),.clk(gclk));
	jdff dff_B_arOPje5Y0_1(.din(n266),.dout(w_dff_B_arOPje5Y0_1),.clk(gclk));
	jdff dff_B_wMWas1jf9_1(.din(w_dff_B_arOPje5Y0_1),.dout(w_dff_B_wMWas1jf9_1),.clk(gclk));
	jdff dff_B_gwwz2dgp4_1(.din(w_dff_B_wMWas1jf9_1),.dout(w_dff_B_gwwz2dgp4_1),.clk(gclk));
	jdff dff_B_UTeYUHQH9_1(.din(w_dff_B_gwwz2dgp4_1),.dout(w_dff_B_UTeYUHQH9_1),.clk(gclk));
	jdff dff_B_4YKhSSsa8_1(.din(w_dff_B_UTeYUHQH9_1),.dout(w_dff_B_4YKhSSsa8_1),.clk(gclk));
	jdff dff_B_KwnugGjf3_1(.din(n267),.dout(w_dff_B_KwnugGjf3_1),.clk(gclk));
	jdff dff_B_zFq2nHU27_1(.din(w_dff_B_KwnugGjf3_1),.dout(w_dff_B_zFq2nHU27_1),.clk(gclk));
	jdff dff_B_swwBgBw02_1(.din(w_dff_B_zFq2nHU27_1),.dout(w_dff_B_swwBgBw02_1),.clk(gclk));
	jdff dff_B_9WkdFLZQ5_1(.din(w_dff_B_swwBgBw02_1),.dout(w_dff_B_9WkdFLZQ5_1),.clk(gclk));
	jdff dff_B_WzV5yZLZ4_1(.din(w_dff_B_9WkdFLZQ5_1),.dout(w_dff_B_WzV5yZLZ4_1),.clk(gclk));
	jdff dff_B_pocnB0Ie0_1(.din(w_dff_B_WzV5yZLZ4_1),.dout(w_dff_B_pocnB0Ie0_1),.clk(gclk));
	jdff dff_B_gNmCbR4p6_1(.din(w_dff_B_pocnB0Ie0_1),.dout(w_dff_B_gNmCbR4p6_1),.clk(gclk));
	jdff dff_B_UVX5Q52q3_1(.din(w_dff_B_gNmCbR4p6_1),.dout(w_dff_B_UVX5Q52q3_1),.clk(gclk));
	jdff dff_B_mFrxlkXZ5_1(.din(w_dff_B_UVX5Q52q3_1),.dout(w_dff_B_mFrxlkXZ5_1),.clk(gclk));
	jdff dff_B_bhNwvLJR9_1(.din(w_dff_B_mFrxlkXZ5_1),.dout(w_dff_B_bhNwvLJR9_1),.clk(gclk));
	jdff dff_B_NwEF1kHj0_1(.din(w_dff_B_bhNwvLJR9_1),.dout(w_dff_B_NwEF1kHj0_1),.clk(gclk));
	jdff dff_B_hNun5WHj5_1(.din(w_dff_B_NwEF1kHj0_1),.dout(w_dff_B_hNun5WHj5_1),.clk(gclk));
	jdff dff_B_m3FlmHAJ4_1(.din(w_dff_B_hNun5WHj5_1),.dout(w_dff_B_m3FlmHAJ4_1),.clk(gclk));
	jdff dff_B_3rIGQKTy5_1(.din(w_dff_B_m3FlmHAJ4_1),.dout(w_dff_B_3rIGQKTy5_1),.clk(gclk));
	jdff dff_B_oZQrNMZb0_1(.din(w_dff_B_3rIGQKTy5_1),.dout(w_dff_B_oZQrNMZb0_1),.clk(gclk));
	jdff dff_B_YQ88Mjss7_1(.din(w_dff_B_oZQrNMZb0_1),.dout(w_dff_B_YQ88Mjss7_1),.clk(gclk));
	jdff dff_B_qmBZId8f7_1(.din(w_dff_B_YQ88Mjss7_1),.dout(w_dff_B_qmBZId8f7_1),.clk(gclk));
	jdff dff_B_MqXRGYB47_1(.din(w_dff_B_qmBZId8f7_1),.dout(w_dff_B_MqXRGYB47_1),.clk(gclk));
	jdff dff_B_sWI2zR2Z2_1(.din(w_dff_B_MqXRGYB47_1),.dout(w_dff_B_sWI2zR2Z2_1),.clk(gclk));
	jdff dff_B_L6dqpViB0_2(.din(n254),.dout(w_dff_B_L6dqpViB0_2),.clk(gclk));
	jdff dff_A_lk5oN2Px8_0(.dout(w_n248_0[0]),.din(w_dff_A_lk5oN2Px8_0),.clk(gclk));
	jdff dff_A_YmGPrnxB0_0(.dout(w_dff_A_lk5oN2Px8_0),.din(w_dff_A_YmGPrnxB0_0),.clk(gclk));
	jdff dff_A_sQdHh1n37_0(.dout(w_dff_A_YmGPrnxB0_0),.din(w_dff_A_sQdHh1n37_0),.clk(gclk));
	jdff dff_B_T4nIGQqQ2_1(.din(n284),.dout(w_dff_B_T4nIGQqQ2_1),.clk(gclk));
	jdff dff_A_pLGLSxkP3_0(.dout(w_n257_0[0]),.din(w_dff_A_pLGLSxkP3_0),.clk(gclk));
	jdff dff_A_6Feo5qj86_0(.dout(w_dff_A_pLGLSxkP3_0),.din(w_dff_A_6Feo5qj86_0),.clk(gclk));
	jdff dff_A_VufXFsyk5_0(.dout(w_dff_A_6Feo5qj86_0),.din(w_dff_A_VufXFsyk5_0),.clk(gclk));
	jdff dff_A_lDO0LMfw6_0(.dout(w_dff_A_VufXFsyk5_0),.din(w_dff_A_lDO0LMfw6_0),.clk(gclk));
	jdff dff_A_w6gnDch55_0(.dout(w_dff_A_lDO0LMfw6_0),.din(w_dff_A_w6gnDch55_0),.clk(gclk));
	jdff dff_A_K4aNRt418_0(.dout(w_dff_A_w6gnDch55_0),.din(w_dff_A_K4aNRt418_0),.clk(gclk));
	jdff dff_B_2uLaRsxG9_1(.din(n256),.dout(w_dff_B_2uLaRsxG9_1),.clk(gclk));
	jdff dff_B_1sNgVaS14_1(.din(w_dff_B_2uLaRsxG9_1),.dout(w_dff_B_1sNgVaS14_1),.clk(gclk));
	jdff dff_B_C2r8BW9j4_1(.din(w_dff_B_1sNgVaS14_1),.dout(w_dff_B_C2r8BW9j4_1),.clk(gclk));
	jdff dff_B_CyXqCiNp0_1(.din(w_dff_B_C2r8BW9j4_1),.dout(w_dff_B_CyXqCiNp0_1),.clk(gclk));
	jdff dff_B_ybIFUs8m1_1(.din(w_dff_B_CyXqCiNp0_1),.dout(w_dff_B_ybIFUs8m1_1),.clk(gclk));
	jdff dff_B_K7INepNu6_1(.din(w_dff_B_ybIFUs8m1_1),.dout(w_dff_B_K7INepNu6_1),.clk(gclk));
	jdff dff_B_sm8nqeof3_1(.din(w_dff_B_K7INepNu6_1),.dout(w_dff_B_sm8nqeof3_1),.clk(gclk));
	jdff dff_B_Gt05Sxcy8_0(.din(n283),.dout(w_dff_B_Gt05Sxcy8_0),.clk(gclk));
	jdff dff_B_F5NQ7doP6_0(.din(w_dff_B_Gt05Sxcy8_0),.dout(w_dff_B_F5NQ7doP6_0),.clk(gclk));
	jdff dff_B_1DnC2YYM8_0(.din(w_dff_B_F5NQ7doP6_0),.dout(w_dff_B_1DnC2YYM8_0),.clk(gclk));
	jdff dff_B_Ia4EvD1F4_0(.din(w_dff_B_1DnC2YYM8_0),.dout(w_dff_B_Ia4EvD1F4_0),.clk(gclk));
	jdff dff_A_y06fDyTX5_1(.dout(w_n253_0[1]),.din(w_dff_A_y06fDyTX5_1),.clk(gclk));
	jdff dff_A_00iMpKMO8_1(.dout(w_dff_A_y06fDyTX5_1),.din(w_dff_A_00iMpKMO8_1),.clk(gclk));
	jdff dff_A_kw7p7WYb9_1(.dout(w_dff_A_00iMpKMO8_1),.din(w_dff_A_kw7p7WYb9_1),.clk(gclk));
	jdff dff_A_n5gMisvx6_1(.dout(w_dff_A_kw7p7WYb9_1),.din(w_dff_A_n5gMisvx6_1),.clk(gclk));
	jdff dff_A_clcYDvzU5_1(.dout(w_dff_A_n5gMisvx6_1),.din(w_dff_A_clcYDvzU5_1),.clk(gclk));
	jdff dff_B_YYPEZ8R58_1(.din(n148),.dout(w_dff_B_YYPEZ8R58_1),.clk(gclk));
	jdff dff_B_qSKNWnMq2_0(.din(n212),.dout(w_dff_B_qSKNWnMq2_0),.clk(gclk));
	jdff dff_A_ZeHLK5Up7_0(.dout(w_n211_0[0]),.din(w_dff_A_ZeHLK5Up7_0),.clk(gclk));
	jdff dff_A_RLuC4rbH2_0(.dout(w_dff_A_ZeHLK5Up7_0),.din(w_dff_A_RLuC4rbH2_0),.clk(gclk));
	jdff dff_A_KjzGsVNx1_0(.dout(w_dff_A_RLuC4rbH2_0),.din(w_dff_A_KjzGsVNx1_0),.clk(gclk));
	jdff dff_A_45igkSop1_0(.dout(w_dff_A_KjzGsVNx1_0),.din(w_dff_A_45igkSop1_0),.clk(gclk));
	jdff dff_A_xBPB0U0t7_0(.dout(w_dff_A_45igkSop1_0),.din(w_dff_A_xBPB0U0t7_0),.clk(gclk));
	jdff dff_A_RLkBIp1p8_0(.dout(w_dff_A_xBPB0U0t7_0),.din(w_dff_A_RLkBIp1p8_0),.clk(gclk));
	jdff dff_A_RolMB63E2_0(.dout(w_n209_0[0]),.din(w_dff_A_RolMB63E2_0),.clk(gclk));
	jdff dff_A_e2DkesIj1_0(.dout(w_dff_A_RolMB63E2_0),.din(w_dff_A_e2DkesIj1_0),.clk(gclk));
	jdff dff_A_VLqdQm978_0(.dout(w_dff_A_e2DkesIj1_0),.din(w_dff_A_VLqdQm978_0),.clk(gclk));
	jdff dff_A_Cit0T6vd5_0(.dout(w_dff_A_VLqdQm978_0),.din(w_dff_A_Cit0T6vd5_0),.clk(gclk));
	jdff dff_A_1IQXxtG49_0(.dout(w_dff_A_Cit0T6vd5_0),.din(w_dff_A_1IQXxtG49_0),.clk(gclk));
	jdff dff_B_5QBn9vwG9_2(.din(n209),.dout(w_dff_B_5QBn9vwG9_2),.clk(gclk));
	jdff dff_B_UvZaV2l65_2(.din(w_dff_B_5QBn9vwG9_2),.dout(w_dff_B_UvZaV2l65_2),.clk(gclk));
	jdff dff_B_Jcb2xc3Y9_2(.din(w_dff_B_UvZaV2l65_2),.dout(w_dff_B_Jcb2xc3Y9_2),.clk(gclk));
	jdff dff_B_IPfJvSUz0_2(.din(w_dff_B_Jcb2xc3Y9_2),.dout(w_dff_B_IPfJvSUz0_2),.clk(gclk));
	jdff dff_B_lKj5Z0wb7_2(.din(w_dff_B_IPfJvSUz0_2),.dout(w_dff_B_lKj5Z0wb7_2),.clk(gclk));
	jdff dff_B_GsCLyO7a6_2(.din(w_dff_B_lKj5Z0wb7_2),.dout(w_dff_B_GsCLyO7a6_2),.clk(gclk));
	jdff dff_B_ckcbK40t4_2(.din(w_dff_B_GsCLyO7a6_2),.dout(w_dff_B_ckcbK40t4_2),.clk(gclk));
	jdff dff_B_zbMJB66E0_2(.din(w_dff_B_ckcbK40t4_2),.dout(w_dff_B_zbMJB66E0_2),.clk(gclk));
	jdff dff_B_pBv53cVB3_2(.din(w_dff_B_zbMJB66E0_2),.dout(w_dff_B_pBv53cVB3_2),.clk(gclk));
	jdff dff_B_u1gy6WZq5_2(.din(w_dff_B_pBv53cVB3_2),.dout(w_dff_B_u1gy6WZq5_2),.clk(gclk));
	jdff dff_B_JK1MxHSR1_2(.din(w_dff_B_u1gy6WZq5_2),.dout(w_dff_B_JK1MxHSR1_2),.clk(gclk));
	jdff dff_B_wxTuSRiP1_2(.din(w_dff_B_JK1MxHSR1_2),.dout(w_dff_B_wxTuSRiP1_2),.clk(gclk));
	jdff dff_B_Y5QRsITF6_2(.din(w_dff_B_wxTuSRiP1_2),.dout(w_dff_B_Y5QRsITF6_2),.clk(gclk));
	jdff dff_B_ZpqHa7210_2(.din(w_dff_B_Y5QRsITF6_2),.dout(w_dff_B_ZpqHa7210_2),.clk(gclk));
	jdff dff_A_Twl7KQTI4_0(.dout(w_n206_0[0]),.din(w_dff_A_Twl7KQTI4_0),.clk(gclk));
	jdff dff_A_2AwORB5l2_0(.dout(w_dff_A_Twl7KQTI4_0),.din(w_dff_A_2AwORB5l2_0),.clk(gclk));
	jdff dff_A_NRKkQU364_0(.dout(w_dff_A_2AwORB5l2_0),.din(w_dff_A_NRKkQU364_0),.clk(gclk));
	jdff dff_A_YW6uijQe5_0(.dout(w_dff_A_NRKkQU364_0),.din(w_dff_A_YW6uijQe5_0),.clk(gclk));
	jdff dff_A_keTKdMYW4_0(.dout(w_dff_A_YW6uijQe5_0),.din(w_dff_A_keTKdMYW4_0),.clk(gclk));
	jdff dff_A_xvjiRNkU4_0(.dout(w_dff_A_keTKdMYW4_0),.din(w_dff_A_xvjiRNkU4_0),.clk(gclk));
	jdff dff_A_zFeo3qiT8_0(.dout(w_n204_0[0]),.din(w_dff_A_zFeo3qiT8_0),.clk(gclk));
	jdff dff_A_KYaFkvxH3_0(.dout(w_dff_A_zFeo3qiT8_0),.din(w_dff_A_KYaFkvxH3_0),.clk(gclk));
	jdff dff_A_AQs67B543_0(.dout(w_dff_A_KYaFkvxH3_0),.din(w_dff_A_AQs67B543_0),.clk(gclk));
	jdff dff_A_GCx0MWnl7_0(.dout(w_dff_A_AQs67B543_0),.din(w_dff_A_GCx0MWnl7_0),.clk(gclk));
	jdff dff_A_FkjMFXXK7_0(.dout(w_dff_A_GCx0MWnl7_0),.din(w_dff_A_FkjMFXXK7_0),.clk(gclk));
	jdff dff_B_pyvjmihX0_2(.din(n204),.dout(w_dff_B_pyvjmihX0_2),.clk(gclk));
	jdff dff_B_Rqoa51le1_2(.din(w_dff_B_pyvjmihX0_2),.dout(w_dff_B_Rqoa51le1_2),.clk(gclk));
	jdff dff_B_FVRNWe4T3_2(.din(w_dff_B_Rqoa51le1_2),.dout(w_dff_B_FVRNWe4T3_2),.clk(gclk));
	jdff dff_B_2aIldgDc7_2(.din(w_dff_B_FVRNWe4T3_2),.dout(w_dff_B_2aIldgDc7_2),.clk(gclk));
	jdff dff_B_3MW6ahhJ6_2(.din(w_dff_B_2aIldgDc7_2),.dout(w_dff_B_3MW6ahhJ6_2),.clk(gclk));
	jdff dff_B_JN560gq67_2(.din(w_dff_B_3MW6ahhJ6_2),.dout(w_dff_B_JN560gq67_2),.clk(gclk));
	jdff dff_B_JiWso3Dt5_2(.din(w_dff_B_JN560gq67_2),.dout(w_dff_B_JiWso3Dt5_2),.clk(gclk));
	jdff dff_B_aoExucFl0_2(.din(w_dff_B_JiWso3Dt5_2),.dout(w_dff_B_aoExucFl0_2),.clk(gclk));
	jdff dff_B_aUO21Keg9_2(.din(w_dff_B_aoExucFl0_2),.dout(w_dff_B_aUO21Keg9_2),.clk(gclk));
	jdff dff_B_D9Qw4Dr58_2(.din(w_dff_B_aUO21Keg9_2),.dout(w_dff_B_D9Qw4Dr58_2),.clk(gclk));
	jdff dff_B_Ctc46mOx3_2(.din(w_dff_B_D9Qw4Dr58_2),.dout(w_dff_B_Ctc46mOx3_2),.clk(gclk));
	jdff dff_B_oPIgScKF0_2(.din(w_dff_B_Ctc46mOx3_2),.dout(w_dff_B_oPIgScKF0_2),.clk(gclk));
	jdff dff_B_x2nzTAyz6_2(.din(w_dff_B_oPIgScKF0_2),.dout(w_dff_B_x2nzTAyz6_2),.clk(gclk));
	jdff dff_B_11kHvXQO6_2(.din(w_dff_B_x2nzTAyz6_2),.dout(w_dff_B_11kHvXQO6_2),.clk(gclk));
	jdff dff_B_EWMUwY8D6_1(.din(n194),.dout(w_dff_B_EWMUwY8D6_1),.clk(gclk));
	jdff dff_B_NoK4utvG1_1(.din(w_dff_B_EWMUwY8D6_1),.dout(w_dff_B_NoK4utvG1_1),.clk(gclk));
	jdff dff_B_dWPghv9I9_1(.din(w_dff_B_NoK4utvG1_1),.dout(w_dff_B_dWPghv9I9_1),.clk(gclk));
	jdff dff_B_dt9IvtXm4_1(.din(w_dff_B_dWPghv9I9_1),.dout(w_dff_B_dt9IvtXm4_1),.clk(gclk));
	jdff dff_B_9lW2wGo79_1(.din(w_dff_B_dt9IvtXm4_1),.dout(w_dff_B_9lW2wGo79_1),.clk(gclk));
	jdff dff_B_NZTeA8Qx8_1(.din(w_dff_B_9lW2wGo79_1),.dout(w_dff_B_NZTeA8Qx8_1),.clk(gclk));
	jdff dff_B_YcQdMbcb1_1(.din(w_dff_B_NZTeA8Qx8_1),.dout(w_dff_B_YcQdMbcb1_1),.clk(gclk));
	jdff dff_B_REjk8CP10_1(.din(w_dff_B_YcQdMbcb1_1),.dout(w_dff_B_REjk8CP10_1),.clk(gclk));
	jdff dff_B_4qvRdGYB5_1(.din(w_dff_B_REjk8CP10_1),.dout(w_dff_B_4qvRdGYB5_1),.clk(gclk));
	jdff dff_B_3wJs1hff5_1(.din(w_dff_B_4qvRdGYB5_1),.dout(w_dff_B_3wJs1hff5_1),.clk(gclk));
	jdff dff_B_JsbSEA9S6_1(.din(w_dff_B_3wJs1hff5_1),.dout(w_dff_B_JsbSEA9S6_1),.clk(gclk));
	jdff dff_B_cHIierqT4_1(.din(w_dff_B_JsbSEA9S6_1),.dout(w_dff_B_cHIierqT4_1),.clk(gclk));
	jdff dff_B_fuA4Pupk1_1(.din(w_dff_B_cHIierqT4_1),.dout(w_dff_B_fuA4Pupk1_1),.clk(gclk));
	jdff dff_B_V6kzopNN6_1(.din(w_dff_B_fuA4Pupk1_1),.dout(w_dff_B_V6kzopNN6_1),.clk(gclk));
	jdff dff_B_q7cwNexr6_1(.din(n190),.dout(w_dff_B_q7cwNexr6_1),.clk(gclk));
	jdff dff_B_23izKn4C8_1(.din(w_dff_B_q7cwNexr6_1),.dout(w_dff_B_23izKn4C8_1),.clk(gclk));
	jdff dff_B_ASLHyAfW8_1(.din(w_dff_B_23izKn4C8_1),.dout(w_dff_B_ASLHyAfW8_1),.clk(gclk));
	jdff dff_B_idwTemFi1_1(.din(w_dff_B_ASLHyAfW8_1),.dout(w_dff_B_idwTemFi1_1),.clk(gclk));
	jdff dff_B_5Ugyj6ki2_1(.din(w_dff_B_idwTemFi1_1),.dout(w_dff_B_5Ugyj6ki2_1),.clk(gclk));
	jdff dff_B_ls6Ys0ht3_1(.din(w_dff_B_5Ugyj6ki2_1),.dout(w_dff_B_ls6Ys0ht3_1),.clk(gclk));
	jdff dff_B_rnRxmECU0_1(.din(w_dff_B_ls6Ys0ht3_1),.dout(w_dff_B_rnRxmECU0_1),.clk(gclk));
	jdff dff_B_8XewBiFj9_1(.din(w_dff_B_rnRxmECU0_1),.dout(w_dff_B_8XewBiFj9_1),.clk(gclk));
	jdff dff_B_Fk3MAnap5_1(.din(w_dff_B_8XewBiFj9_1),.dout(w_dff_B_Fk3MAnap5_1),.clk(gclk));
	jdff dff_B_w2tuWnAq2_1(.din(w_dff_B_Fk3MAnap5_1),.dout(w_dff_B_w2tuWnAq2_1),.clk(gclk));
	jdff dff_B_MQS63P3w3_1(.din(w_dff_B_w2tuWnAq2_1),.dout(w_dff_B_MQS63P3w3_1),.clk(gclk));
	jdff dff_B_2rjG9oEl4_1(.din(w_dff_B_MQS63P3w3_1),.dout(w_dff_B_2rjG9oEl4_1),.clk(gclk));
	jdff dff_B_M3IeiHw62_1(.din(w_dff_B_2rjG9oEl4_1),.dout(w_dff_B_M3IeiHw62_1),.clk(gclk));
	jdff dff_B_1ab0SRD63_1(.din(w_dff_B_M3IeiHw62_1),.dout(w_dff_B_1ab0SRD63_1),.clk(gclk));
	jdff dff_A_qEHxUWUw7_0(.dout(w_n185_0[0]),.din(w_dff_A_qEHxUWUw7_0),.clk(gclk));
	jdff dff_A_nmowiDWS1_0(.dout(w_dff_A_qEHxUWUw7_0),.din(w_dff_A_nmowiDWS1_0),.clk(gclk));
	jdff dff_A_wtAqk43u5_0(.dout(w_dff_A_nmowiDWS1_0),.din(w_dff_A_wtAqk43u5_0),.clk(gclk));
	jdff dff_A_o5aZb5hM7_0(.dout(w_dff_A_wtAqk43u5_0),.din(w_dff_A_o5aZb5hM7_0),.clk(gclk));
	jdff dff_A_KfpRo5LZ4_0(.dout(w_dff_A_o5aZb5hM7_0),.din(w_dff_A_KfpRo5LZ4_0),.clk(gclk));
	jdff dff_B_w3nCi8Ca7_2(.din(n185),.dout(w_dff_B_w3nCi8Ca7_2),.clk(gclk));
	jdff dff_B_X9S9FndA7_2(.din(w_dff_B_w3nCi8Ca7_2),.dout(w_dff_B_X9S9FndA7_2),.clk(gclk));
	jdff dff_B_Poaye4d59_2(.din(w_dff_B_X9S9FndA7_2),.dout(w_dff_B_Poaye4d59_2),.clk(gclk));
	jdff dff_B_aqUtM0TL6_2(.din(w_dff_B_Poaye4d59_2),.dout(w_dff_B_aqUtM0TL6_2),.clk(gclk));
	jdff dff_B_BrvhUVLZ7_2(.din(w_dff_B_aqUtM0TL6_2),.dout(w_dff_B_BrvhUVLZ7_2),.clk(gclk));
	jdff dff_B_pjjIQtIO9_2(.din(w_dff_B_BrvhUVLZ7_2),.dout(w_dff_B_pjjIQtIO9_2),.clk(gclk));
	jdff dff_B_cU2FmDGn3_2(.din(w_dff_B_pjjIQtIO9_2),.dout(w_dff_B_cU2FmDGn3_2),.clk(gclk));
	jdff dff_B_L2vDqohC6_2(.din(w_dff_B_cU2FmDGn3_2),.dout(w_dff_B_L2vDqohC6_2),.clk(gclk));
	jdff dff_B_Q7kbfaUg1_2(.din(w_dff_B_L2vDqohC6_2),.dout(w_dff_B_Q7kbfaUg1_2),.clk(gclk));
	jdff dff_B_63kkTZgB6_2(.din(w_dff_B_Q7kbfaUg1_2),.dout(w_dff_B_63kkTZgB6_2),.clk(gclk));
	jdff dff_B_ggr7m1UT8_2(.din(w_dff_B_63kkTZgB6_2),.dout(w_dff_B_ggr7m1UT8_2),.clk(gclk));
	jdff dff_B_SOcydkLC5_2(.din(w_dff_B_ggr7m1UT8_2),.dout(w_dff_B_SOcydkLC5_2),.clk(gclk));
	jdff dff_B_7yBeHPJ67_2(.din(w_dff_B_SOcydkLC5_2),.dout(w_dff_B_7yBeHPJ67_2),.clk(gclk));
	jdff dff_B_8zFPGK4q8_2(.din(w_dff_B_7yBeHPJ67_2),.dout(w_dff_B_8zFPGK4q8_2),.clk(gclk));
	jdff dff_B_Dxuofd8Z2_2(.din(n281),.dout(w_dff_B_Dxuofd8Z2_2),.clk(gclk));
	jdff dff_A_T9mV3NnG5_0(.dout(w_n149_0[0]),.din(w_dff_A_T9mV3NnG5_0),.clk(gclk));
	jdff dff_A_OZYfqWzk6_0(.dout(w_dff_A_T9mV3NnG5_0),.din(w_dff_A_OZYfqWzk6_0),.clk(gclk));
	jdff dff_A_aUFXydqr0_0(.dout(w_dff_A_OZYfqWzk6_0),.din(w_dff_A_aUFXydqr0_0),.clk(gclk));
	jdff dff_A_iyzUq9O70_0(.dout(w_dff_A_aUFXydqr0_0),.din(w_dff_A_iyzUq9O70_0),.clk(gclk));
	jdff dff_A_xQpPy1Km9_0(.dout(w_dff_A_iyzUq9O70_0),.din(w_dff_A_xQpPy1Km9_0),.clk(gclk));
	jdff dff_B_4HDTrH7R5_2(.din(n149),.dout(w_dff_B_4HDTrH7R5_2),.clk(gclk));
	jdff dff_B_u1Yo01bb8_2(.din(w_dff_B_4HDTrH7R5_2),.dout(w_dff_B_u1Yo01bb8_2),.clk(gclk));
	jdff dff_B_G8MiyEs00_2(.din(w_dff_B_u1Yo01bb8_2),.dout(w_dff_B_G8MiyEs00_2),.clk(gclk));
	jdff dff_B_H31XRr0r0_2(.din(w_dff_B_G8MiyEs00_2),.dout(w_dff_B_H31XRr0r0_2),.clk(gclk));
	jdff dff_B_G5dnU2xU5_2(.din(w_dff_B_H31XRr0r0_2),.dout(w_dff_B_G5dnU2xU5_2),.clk(gclk));
	jdff dff_B_sMGCvCnC6_2(.din(w_dff_B_G5dnU2xU5_2),.dout(w_dff_B_sMGCvCnC6_2),.clk(gclk));
	jdff dff_B_OEi3EvXT8_2(.din(w_dff_B_sMGCvCnC6_2),.dout(w_dff_B_OEi3EvXT8_2),.clk(gclk));
	jdff dff_B_hUJnCLyW7_2(.din(w_dff_B_OEi3EvXT8_2),.dout(w_dff_B_hUJnCLyW7_2),.clk(gclk));
	jdff dff_B_jxfeYicl8_2(.din(w_dff_B_hUJnCLyW7_2),.dout(w_dff_B_jxfeYicl8_2),.clk(gclk));
	jdff dff_B_htpEslNe9_2(.din(w_dff_B_jxfeYicl8_2),.dout(w_dff_B_htpEslNe9_2),.clk(gclk));
	jdff dff_B_8Hw6z0XB2_2(.din(w_dff_B_htpEslNe9_2),.dout(w_dff_B_8Hw6z0XB2_2),.clk(gclk));
	jdff dff_B_FNTAziHu9_2(.din(w_dff_B_8Hw6z0XB2_2),.dout(w_dff_B_FNTAziHu9_2),.clk(gclk));
	jdff dff_B_urenHQeE1_2(.din(w_dff_B_FNTAziHu9_2),.dout(w_dff_B_urenHQeE1_2),.clk(gclk));
	jdff dff_B_Ao6Eg4Y10_2(.din(w_dff_B_urenHQeE1_2),.dout(w_dff_B_Ao6Eg4Y10_2),.clk(gclk));
	jdff dff_A_PbtSaNKS8_0(.dout(w_n183_0[0]),.din(w_dff_A_PbtSaNKS8_0),.clk(gclk));
	jdff dff_A_u0WAQt203_0(.dout(w_dff_A_PbtSaNKS8_0),.din(w_dff_A_u0WAQt203_0),.clk(gclk));
	jdff dff_A_crKpqWTZ5_0(.dout(w_dff_A_u0WAQt203_0),.din(w_dff_A_crKpqWTZ5_0),.clk(gclk));
	jdff dff_A_ls0Xmgj72_0(.dout(w_dff_A_crKpqWTZ5_0),.din(w_dff_A_ls0Xmgj72_0),.clk(gclk));
	jdff dff_A_BHv2sUzV1_0(.dout(w_dff_A_ls0Xmgj72_0),.din(w_dff_A_BHv2sUzV1_0),.clk(gclk));
	jdff dff_A_npMJPdxG5_0(.dout(w_dff_A_BHv2sUzV1_0),.din(w_dff_A_npMJPdxG5_0),.clk(gclk));
	jdff dff_A_2cuzIc1f9_0(.dout(w_n271_0[0]),.din(w_dff_A_2cuzIc1f9_0),.clk(gclk));
	jdff dff_A_HkdP4Wa46_0(.dout(w_dff_A_2cuzIc1f9_0),.din(w_dff_A_HkdP4Wa46_0),.clk(gclk));
	jdff dff_A_re46KwVH6_0(.dout(w_dff_A_HkdP4Wa46_0),.din(w_dff_A_re46KwVH6_0),.clk(gclk));
	jdff dff_B_LR9dAh5R7_1(.din(n217),.dout(w_dff_B_LR9dAh5R7_1),.clk(gclk));
	jdff dff_B_B7W15AHw3_0(.din(n243),.dout(w_dff_B_B7W15AHw3_0),.clk(gclk));
	jdff dff_A_XrnIk4bn8_0(.dout(w_G27gat_0[0]),.din(w_dff_A_XrnIk4bn8_0),.clk(gclk));
	jdff dff_A_2ot3g6Jk2_0(.dout(w_dff_A_XrnIk4bn8_0),.din(w_dff_A_2ot3g6Jk2_0),.clk(gclk));
	jdff dff_A_X3C8Pmc37_0(.dout(w_dff_A_2ot3g6Jk2_0),.din(w_dff_A_X3C8Pmc37_0),.clk(gclk));
	jdff dff_A_xQdhGddt2_0(.dout(w_dff_A_X3C8Pmc37_0),.din(w_dff_A_xQdhGddt2_0),.clk(gclk));
	jdff dff_A_XWQsult97_0(.dout(w_dff_A_xQdhGddt2_0),.din(w_dff_A_XWQsult97_0),.clk(gclk));
	jdff dff_A_Q6oFFsFn8_0(.dout(w_dff_A_XWQsult97_0),.din(w_dff_A_Q6oFFsFn8_0),.clk(gclk));
	jdff dff_A_bW5LykPj5_0(.dout(w_dff_A_Q6oFFsFn8_0),.din(w_dff_A_bW5LykPj5_0),.clk(gclk));
	jdff dff_A_JXKToiTb4_0(.dout(w_dff_A_bW5LykPj5_0),.din(w_dff_A_JXKToiTb4_0),.clk(gclk));
	jdff dff_A_PXdvU1ov1_0(.dout(w_dff_A_JXKToiTb4_0),.din(w_dff_A_PXdvU1ov1_0),.clk(gclk));
	jdff dff_A_em0haHZN6_0(.dout(w_dff_A_PXdvU1ov1_0),.din(w_dff_A_em0haHZN6_0),.clk(gclk));
	jdff dff_A_2e6k5BFq9_0(.dout(w_dff_A_em0haHZN6_0),.din(w_dff_A_2e6k5BFq9_0),.clk(gclk));
	jdff dff_A_tdukIwAy8_0(.dout(w_dff_A_2e6k5BFq9_0),.din(w_dff_A_tdukIwAy8_0),.clk(gclk));
	jdff dff_A_M29Fgj9d8_0(.dout(w_dff_A_tdukIwAy8_0),.din(w_dff_A_M29Fgj9d8_0),.clk(gclk));
	jdff dff_A_xTlXDaKf3_0(.dout(w_dff_A_M29Fgj9d8_0),.din(w_dff_A_xTlXDaKf3_0),.clk(gclk));
	jdff dff_A_t1lvHTWN3_0(.dout(w_dff_A_xTlXDaKf3_0),.din(w_dff_A_t1lvHTWN3_0),.clk(gclk));
	jdff dff_A_gQ4GPX5n4_0(.dout(w_G115gat_0[0]),.din(w_dff_A_gQ4GPX5n4_0),.clk(gclk));
	jdff dff_A_bcu8cZWX0_0(.dout(w_dff_A_gQ4GPX5n4_0),.din(w_dff_A_bcu8cZWX0_0),.clk(gclk));
	jdff dff_A_HozFfQbX4_0(.dout(w_dff_A_bcu8cZWX0_0),.din(w_dff_A_HozFfQbX4_0),.clk(gclk));
	jdff dff_A_5Y8CGgZd9_0(.dout(w_dff_A_HozFfQbX4_0),.din(w_dff_A_5Y8CGgZd9_0),.clk(gclk));
	jdff dff_A_9dtdvi1f9_0(.dout(w_dff_A_5Y8CGgZd9_0),.din(w_dff_A_9dtdvi1f9_0),.clk(gclk));
	jdff dff_A_OPd7hUjC2_0(.dout(w_dff_A_9dtdvi1f9_0),.din(w_dff_A_OPd7hUjC2_0),.clk(gclk));
	jdff dff_A_fdKUXmEi0_0(.dout(w_dff_A_OPd7hUjC2_0),.din(w_dff_A_fdKUXmEi0_0),.clk(gclk));
	jdff dff_A_ZzhT5Luj8_0(.dout(w_dff_A_fdKUXmEi0_0),.din(w_dff_A_ZzhT5Luj8_0),.clk(gclk));
	jdff dff_A_FeSuzuR20_0(.dout(w_dff_A_ZzhT5Luj8_0),.din(w_dff_A_FeSuzuR20_0),.clk(gclk));
	jdff dff_A_Bk0xriSz6_0(.dout(w_dff_A_FeSuzuR20_0),.din(w_dff_A_Bk0xriSz6_0),.clk(gclk));
	jdff dff_A_pSUpvoc61_0(.dout(w_dff_A_Bk0xriSz6_0),.din(w_dff_A_pSUpvoc61_0),.clk(gclk));
	jdff dff_A_TeHHmgXQ8_0(.dout(w_dff_A_pSUpvoc61_0),.din(w_dff_A_TeHHmgXQ8_0),.clk(gclk));
	jdff dff_A_c897qPZX6_0(.dout(w_dff_A_TeHHmgXQ8_0),.din(w_dff_A_c897qPZX6_0),.clk(gclk));
	jdff dff_A_m2FxBFAN5_0(.dout(w_dff_A_c897qPZX6_0),.din(w_dff_A_m2FxBFAN5_0),.clk(gclk));
	jdff dff_A_BrB88TYv0_0(.dout(w_dff_A_m2FxBFAN5_0),.din(w_dff_A_BrB88TYv0_0),.clk(gclk));
	jdff dff_A_TE5ZFhsM0_0(.dout(w_n230_0[0]),.din(w_dff_A_TE5ZFhsM0_0),.clk(gclk));
	jdff dff_A_B8wPd7556_0(.dout(w_dff_A_TE5ZFhsM0_0),.din(w_dff_A_B8wPd7556_0),.clk(gclk));
	jdff dff_A_gxksOdZQ9_0(.dout(w_dff_A_B8wPd7556_0),.din(w_dff_A_gxksOdZQ9_0),.clk(gclk));
	jdff dff_A_SUSk2GZb9_0(.dout(w_dff_A_gxksOdZQ9_0),.din(w_dff_A_SUSk2GZb9_0),.clk(gclk));
	jdff dff_A_w9cGeVtq8_0(.dout(w_dff_A_SUSk2GZb9_0),.din(w_dff_A_w9cGeVtq8_0),.clk(gclk));
	jdff dff_A_MYdu8TrK4_0(.dout(w_dff_A_w9cGeVtq8_0),.din(w_dff_A_MYdu8TrK4_0),.clk(gclk));
	jdff dff_A_XPwPzKIp6_0(.dout(w_G92gat_0[0]),.din(w_dff_A_XPwPzKIp6_0),.clk(gclk));
	jdff dff_A_9IRuOFH21_0(.dout(w_dff_A_XPwPzKIp6_0),.din(w_dff_A_9IRuOFH21_0),.clk(gclk));
	jdff dff_A_IUafJYUi9_0(.dout(w_dff_A_9IRuOFH21_0),.din(w_dff_A_IUafJYUi9_0),.clk(gclk));
	jdff dff_A_k7Ha5SNK8_0(.dout(w_dff_A_IUafJYUi9_0),.din(w_dff_A_k7Ha5SNK8_0),.clk(gclk));
	jdff dff_A_EC2q37lL9_0(.dout(w_dff_A_k7Ha5SNK8_0),.din(w_dff_A_EC2q37lL9_0),.clk(gclk));
	jdff dff_A_77MK1I3v7_0(.dout(w_dff_A_EC2q37lL9_0),.din(w_dff_A_77MK1I3v7_0),.clk(gclk));
	jdff dff_A_mSy5WXBu8_0(.dout(w_dff_A_77MK1I3v7_0),.din(w_dff_A_mSy5WXBu8_0),.clk(gclk));
	jdff dff_A_EQPuw4Xx8_0(.dout(w_dff_A_mSy5WXBu8_0),.din(w_dff_A_EQPuw4Xx8_0),.clk(gclk));
	jdff dff_A_ZEM7Owvf2_0(.dout(w_dff_A_EQPuw4Xx8_0),.din(w_dff_A_ZEM7Owvf2_0),.clk(gclk));
	jdff dff_A_3jxfSrxU6_0(.dout(w_dff_A_ZEM7Owvf2_0),.din(w_dff_A_3jxfSrxU6_0),.clk(gclk));
	jdff dff_A_4vCTaY2l7_0(.dout(w_dff_A_3jxfSrxU6_0),.din(w_dff_A_4vCTaY2l7_0),.clk(gclk));
	jdff dff_A_ge7cvY329_0(.dout(w_dff_A_4vCTaY2l7_0),.din(w_dff_A_ge7cvY329_0),.clk(gclk));
	jdff dff_A_nKvyGjSi1_0(.dout(w_dff_A_ge7cvY329_0),.din(w_dff_A_nKvyGjSi1_0),.clk(gclk));
	jdff dff_A_s80YZnEh9_0(.dout(w_dff_A_nKvyGjSi1_0),.din(w_dff_A_s80YZnEh9_0),.clk(gclk));
	jdff dff_A_2tdWEtSC8_0(.dout(w_dff_A_s80YZnEh9_0),.din(w_dff_A_2tdWEtSC8_0),.clk(gclk));
	jdff dff_A_B20RmEEi8_0(.dout(w_dff_A_2tdWEtSC8_0),.din(w_dff_A_B20RmEEi8_0),.clk(gclk));
	jdff dff_A_ul9HRwnU4_0(.dout(w_dff_A_B20RmEEi8_0),.din(w_dff_A_ul9HRwnU4_0),.clk(gclk));
	jdff dff_A_A0eZaJkW1_0(.dout(w_dff_A_ul9HRwnU4_0),.din(w_dff_A_A0eZaJkW1_0),.clk(gclk));
	jdff dff_A_Htdhkaoi2_0(.dout(w_dff_A_A0eZaJkW1_0),.din(w_dff_A_Htdhkaoi2_0),.clk(gclk));
	jdff dff_A_sHVhMF8S9_0(.dout(w_dff_A_Htdhkaoi2_0),.din(w_dff_A_sHVhMF8S9_0),.clk(gclk));
	jdff dff_A_mnRhacPx5_1(.dout(w_G92gat_0[1]),.din(w_dff_A_mnRhacPx5_1),.clk(gclk));
	jdff dff_A_zP7Ve7Rj5_1(.dout(w_dff_A_mnRhacPx5_1),.din(w_dff_A_zP7Ve7Rj5_1),.clk(gclk));
	jdff dff_A_9WgDQZaW4_1(.dout(w_dff_A_zP7Ve7Rj5_1),.din(w_dff_A_9WgDQZaW4_1),.clk(gclk));
	jdff dff_A_rH22nS0W6_1(.dout(w_dff_A_9WgDQZaW4_1),.din(w_dff_A_rH22nS0W6_1),.clk(gclk));
	jdff dff_A_FVBT3PBs0_1(.dout(w_dff_A_rH22nS0W6_1),.din(w_dff_A_FVBT3PBs0_1),.clk(gclk));
	jdff dff_A_UcHNbOBb1_1(.dout(w_dff_A_FVBT3PBs0_1),.din(w_dff_A_UcHNbOBb1_1),.clk(gclk));
	jdff dff_A_a4uJBmZA5_1(.dout(w_dff_A_UcHNbOBb1_1),.din(w_dff_A_a4uJBmZA5_1),.clk(gclk));
	jdff dff_A_McnMWF4i8_1(.dout(w_dff_A_a4uJBmZA5_1),.din(w_dff_A_McnMWF4i8_1),.clk(gclk));
	jdff dff_A_kh3xpoMR7_1(.dout(w_dff_A_McnMWF4i8_1),.din(w_dff_A_kh3xpoMR7_1),.clk(gclk));
	jdff dff_A_FSe6SYPE6_1(.dout(w_dff_A_kh3xpoMR7_1),.din(w_dff_A_FSe6SYPE6_1),.clk(gclk));
	jdff dff_A_AHjkNldU9_1(.dout(w_dff_A_FSe6SYPE6_1),.din(w_dff_A_AHjkNldU9_1),.clk(gclk));
	jdff dff_A_DkAf5t1k3_1(.dout(w_dff_A_AHjkNldU9_1),.din(w_dff_A_DkAf5t1k3_1),.clk(gclk));
	jdff dff_A_6JHxCAyW2_1(.dout(w_dff_A_DkAf5t1k3_1),.din(w_dff_A_6JHxCAyW2_1),.clk(gclk));
	jdff dff_A_4LA2JJJp0_1(.dout(w_dff_A_6JHxCAyW2_1),.din(w_dff_A_4LA2JJJp0_1),.clk(gclk));
	jdff dff_A_YT8iWFLb1_1(.dout(w_dff_A_4LA2JJJp0_1),.din(w_dff_A_YT8iWFLb1_1),.clk(gclk));
	jdff dff_A_5YFQazP93_0(.dout(w_n227_0[0]),.din(w_dff_A_5YFQazP93_0),.clk(gclk));
	jdff dff_A_nPCNiFv90_0(.dout(w_dff_A_5YFQazP93_0),.din(w_dff_A_nPCNiFv90_0),.clk(gclk));
	jdff dff_A_fCmm0Yfz5_0(.dout(w_dff_A_nPCNiFv90_0),.din(w_dff_A_fCmm0Yfz5_0),.clk(gclk));
	jdff dff_A_R2rr5sTk3_0(.dout(w_dff_A_fCmm0Yfz5_0),.din(w_dff_A_R2rr5sTk3_0),.clk(gclk));
	jdff dff_A_iXbJSuJB2_0(.dout(w_dff_A_R2rr5sTk3_0),.din(w_dff_A_iXbJSuJB2_0),.clk(gclk));
	jdff dff_A_URiQhGSh9_0(.dout(w_dff_A_iXbJSuJB2_0),.din(w_dff_A_URiQhGSh9_0),.clk(gclk));
	jdff dff_A_omBVryHd6_0(.dout(w_G14gat_0[0]),.din(w_dff_A_omBVryHd6_0),.clk(gclk));
	jdff dff_A_rdeVdRNz3_0(.dout(w_dff_A_omBVryHd6_0),.din(w_dff_A_rdeVdRNz3_0),.clk(gclk));
	jdff dff_A_9oXFHW0V8_0(.dout(w_dff_A_rdeVdRNz3_0),.din(w_dff_A_9oXFHW0V8_0),.clk(gclk));
	jdff dff_A_b6jPoXU51_0(.dout(w_dff_A_9oXFHW0V8_0),.din(w_dff_A_b6jPoXU51_0),.clk(gclk));
	jdff dff_A_LsBEZ58d8_0(.dout(w_dff_A_b6jPoXU51_0),.din(w_dff_A_LsBEZ58d8_0),.clk(gclk));
	jdff dff_A_ggeOITuZ3_0(.dout(w_dff_A_LsBEZ58d8_0),.din(w_dff_A_ggeOITuZ3_0),.clk(gclk));
	jdff dff_A_6xg5YICe5_0(.dout(w_dff_A_ggeOITuZ3_0),.din(w_dff_A_6xg5YICe5_0),.clk(gclk));
	jdff dff_A_0fZNLKVp9_0(.dout(w_dff_A_6xg5YICe5_0),.din(w_dff_A_0fZNLKVp9_0),.clk(gclk));
	jdff dff_A_3rxHug5I6_0(.dout(w_dff_A_0fZNLKVp9_0),.din(w_dff_A_3rxHug5I6_0),.clk(gclk));
	jdff dff_A_SmMkBNte8_0(.dout(w_dff_A_3rxHug5I6_0),.din(w_dff_A_SmMkBNte8_0),.clk(gclk));
	jdff dff_A_7oKWTgbK1_0(.dout(w_dff_A_SmMkBNte8_0),.din(w_dff_A_7oKWTgbK1_0),.clk(gclk));
	jdff dff_A_8c7QOeGs8_0(.dout(w_dff_A_7oKWTgbK1_0),.din(w_dff_A_8c7QOeGs8_0),.clk(gclk));
	jdff dff_A_qNYUmA6T4_0(.dout(w_dff_A_8c7QOeGs8_0),.din(w_dff_A_qNYUmA6T4_0),.clk(gclk));
	jdff dff_A_oYrNu0tu8_0(.dout(w_dff_A_qNYUmA6T4_0),.din(w_dff_A_oYrNu0tu8_0),.clk(gclk));
	jdff dff_A_0uYgz50H6_0(.dout(w_dff_A_oYrNu0tu8_0),.din(w_dff_A_0uYgz50H6_0),.clk(gclk));
	jdff dff_A_t1Pd64y51_0(.dout(w_dff_A_0uYgz50H6_0),.din(w_dff_A_t1Pd64y51_0),.clk(gclk));
	jdff dff_A_uQBwZtPd6_0(.dout(w_dff_A_t1Pd64y51_0),.din(w_dff_A_uQBwZtPd6_0),.clk(gclk));
	jdff dff_A_Ffetb79U9_0(.dout(w_dff_A_uQBwZtPd6_0),.din(w_dff_A_Ffetb79U9_0),.clk(gclk));
	jdff dff_A_XLIG9Ewp3_0(.dout(w_dff_A_Ffetb79U9_0),.din(w_dff_A_XLIG9Ewp3_0),.clk(gclk));
	jdff dff_A_B9LX9zz21_0(.dout(w_dff_A_XLIG9Ewp3_0),.din(w_dff_A_B9LX9zz21_0),.clk(gclk));
	jdff dff_A_oWXfa6Cc4_1(.dout(w_G14gat_0[1]),.din(w_dff_A_oWXfa6Cc4_1),.clk(gclk));
	jdff dff_A_rdmP5a6T0_1(.dout(w_dff_A_oWXfa6Cc4_1),.din(w_dff_A_rdmP5a6T0_1),.clk(gclk));
	jdff dff_A_RzYyp0Ox5_1(.dout(w_dff_A_rdmP5a6T0_1),.din(w_dff_A_RzYyp0Ox5_1),.clk(gclk));
	jdff dff_A_ZMBjp6Q04_1(.dout(w_dff_A_RzYyp0Ox5_1),.din(w_dff_A_ZMBjp6Q04_1),.clk(gclk));
	jdff dff_A_nYGzuNUw7_1(.dout(w_dff_A_ZMBjp6Q04_1),.din(w_dff_A_nYGzuNUw7_1),.clk(gclk));
	jdff dff_A_u10Rjnzn5_1(.dout(w_dff_A_nYGzuNUw7_1),.din(w_dff_A_u10Rjnzn5_1),.clk(gclk));
	jdff dff_A_xDbOsd0l1_1(.dout(w_dff_A_u10Rjnzn5_1),.din(w_dff_A_xDbOsd0l1_1),.clk(gclk));
	jdff dff_A_fdyWZa240_1(.dout(w_dff_A_xDbOsd0l1_1),.din(w_dff_A_fdyWZa240_1),.clk(gclk));
	jdff dff_A_0Y0QXG8n4_1(.dout(w_dff_A_fdyWZa240_1),.din(w_dff_A_0Y0QXG8n4_1),.clk(gclk));
	jdff dff_A_AQjnpTW43_1(.dout(w_dff_A_0Y0QXG8n4_1),.din(w_dff_A_AQjnpTW43_1),.clk(gclk));
	jdff dff_A_pTR124rD5_1(.dout(w_dff_A_AQjnpTW43_1),.din(w_dff_A_pTR124rD5_1),.clk(gclk));
	jdff dff_A_RNUZXDNp4_1(.dout(w_dff_A_pTR124rD5_1),.din(w_dff_A_RNUZXDNp4_1),.clk(gclk));
	jdff dff_A_NKQ4mBEE9_1(.dout(w_dff_A_RNUZXDNp4_1),.din(w_dff_A_NKQ4mBEE9_1),.clk(gclk));
	jdff dff_A_RXeTVk6A3_1(.dout(w_dff_A_NKQ4mBEE9_1),.din(w_dff_A_RXeTVk6A3_1),.clk(gclk));
	jdff dff_A_iA559QVq3_1(.dout(w_dff_A_RXeTVk6A3_1),.din(w_dff_A_iA559QVq3_1),.clk(gclk));
	jdff dff_B_TSGJYjC88_1(.din(n221),.dout(w_dff_B_TSGJYjC88_1),.clk(gclk));
	jdff dff_B_Vor8q6b36_1(.din(w_dff_B_TSGJYjC88_1),.dout(w_dff_B_Vor8q6b36_1),.clk(gclk));
	jdff dff_B_t1m9d1w16_1(.din(w_dff_B_Vor8q6b36_1),.dout(w_dff_B_t1m9d1w16_1),.clk(gclk));
	jdff dff_B_h1iPyZE83_1(.din(w_dff_B_t1m9d1w16_1),.dout(w_dff_B_h1iPyZE83_1),.clk(gclk));
	jdff dff_B_0zhaWSMg6_1(.din(w_dff_B_h1iPyZE83_1),.dout(w_dff_B_0zhaWSMg6_1),.clk(gclk));
	jdff dff_A_YA4T75yo6_0(.dout(w_G66gat_0[0]),.din(w_dff_A_YA4T75yo6_0),.clk(gclk));
	jdff dff_A_hodyrOoN8_0(.dout(w_dff_A_YA4T75yo6_0),.din(w_dff_A_hodyrOoN8_0),.clk(gclk));
	jdff dff_A_7QvCauur8_0(.dout(w_dff_A_hodyrOoN8_0),.din(w_dff_A_7QvCauur8_0),.clk(gclk));
	jdff dff_A_D0tRt7ml1_0(.dout(w_dff_A_7QvCauur8_0),.din(w_dff_A_D0tRt7ml1_0),.clk(gclk));
	jdff dff_A_DGCf7jsN3_0(.dout(w_dff_A_D0tRt7ml1_0),.din(w_dff_A_DGCf7jsN3_0),.clk(gclk));
	jdff dff_A_L4RaDarK3_0(.dout(w_dff_A_DGCf7jsN3_0),.din(w_dff_A_L4RaDarK3_0),.clk(gclk));
	jdff dff_A_fMGEdRT69_0(.dout(w_dff_A_L4RaDarK3_0),.din(w_dff_A_fMGEdRT69_0),.clk(gclk));
	jdff dff_A_k5vx8KWr9_0(.dout(w_dff_A_fMGEdRT69_0),.din(w_dff_A_k5vx8KWr9_0),.clk(gclk));
	jdff dff_A_iKdmFnYb9_0(.dout(w_dff_A_k5vx8KWr9_0),.din(w_dff_A_iKdmFnYb9_0),.clk(gclk));
	jdff dff_A_HfdzV5iC9_0(.dout(w_dff_A_iKdmFnYb9_0),.din(w_dff_A_HfdzV5iC9_0),.clk(gclk));
	jdff dff_A_aLG49hB42_0(.dout(w_dff_A_HfdzV5iC9_0),.din(w_dff_A_aLG49hB42_0),.clk(gclk));
	jdff dff_A_ueuykuks7_0(.dout(w_dff_A_aLG49hB42_0),.din(w_dff_A_ueuykuks7_0),.clk(gclk));
	jdff dff_A_ZhVJwpZO3_0(.dout(w_dff_A_ueuykuks7_0),.din(w_dff_A_ZhVJwpZO3_0),.clk(gclk));
	jdff dff_A_YJBSrbur9_0(.dout(w_dff_A_ZhVJwpZO3_0),.din(w_dff_A_YJBSrbur9_0),.clk(gclk));
	jdff dff_A_iWhog36v9_0(.dout(w_dff_A_YJBSrbur9_0),.din(w_dff_A_iWhog36v9_0),.clk(gclk));
	jdff dff_A_M2OIffg29_0(.dout(w_dff_A_iWhog36v9_0),.din(w_dff_A_M2OIffg29_0),.clk(gclk));
	jdff dff_A_u07h95AP6_0(.dout(w_dff_A_M2OIffg29_0),.din(w_dff_A_u07h95AP6_0),.clk(gclk));
	jdff dff_A_4T3hAL9z2_0(.dout(w_dff_A_u07h95AP6_0),.din(w_dff_A_4T3hAL9z2_0),.clk(gclk));
	jdff dff_A_LoBPcUcI0_0(.dout(w_dff_A_4T3hAL9z2_0),.din(w_dff_A_LoBPcUcI0_0),.clk(gclk));
	jdff dff_A_40SG9CPg4_0(.dout(w_dff_A_LoBPcUcI0_0),.din(w_dff_A_40SG9CPg4_0),.clk(gclk));
	jdff dff_A_NMf0EbFR5_1(.dout(w_G66gat_0[1]),.din(w_dff_A_NMf0EbFR5_1),.clk(gclk));
	jdff dff_A_9XnP4ArK7_1(.dout(w_dff_A_NMf0EbFR5_1),.din(w_dff_A_9XnP4ArK7_1),.clk(gclk));
	jdff dff_A_tJAVIllD3_1(.dout(w_dff_A_9XnP4ArK7_1),.din(w_dff_A_tJAVIllD3_1),.clk(gclk));
	jdff dff_A_NMUZW6aA8_1(.dout(w_dff_A_tJAVIllD3_1),.din(w_dff_A_NMUZW6aA8_1),.clk(gclk));
	jdff dff_A_ajNIy8Tk0_1(.dout(w_dff_A_NMUZW6aA8_1),.din(w_dff_A_ajNIy8Tk0_1),.clk(gclk));
	jdff dff_A_4X8tPYDK9_1(.dout(w_dff_A_ajNIy8Tk0_1),.din(w_dff_A_4X8tPYDK9_1),.clk(gclk));
	jdff dff_A_kwZueTpZ6_1(.dout(w_dff_A_4X8tPYDK9_1),.din(w_dff_A_kwZueTpZ6_1),.clk(gclk));
	jdff dff_A_GYzVYy4W4_1(.dout(w_dff_A_kwZueTpZ6_1),.din(w_dff_A_GYzVYy4W4_1),.clk(gclk));
	jdff dff_A_ICeUlMas8_1(.dout(w_dff_A_GYzVYy4W4_1),.din(w_dff_A_ICeUlMas8_1),.clk(gclk));
	jdff dff_A_G1YXUitm2_1(.dout(w_dff_A_ICeUlMas8_1),.din(w_dff_A_G1YXUitm2_1),.clk(gclk));
	jdff dff_A_UbNZK9ix3_1(.dout(w_dff_A_G1YXUitm2_1),.din(w_dff_A_UbNZK9ix3_1),.clk(gclk));
	jdff dff_A_k1WU7RTL7_1(.dout(w_dff_A_UbNZK9ix3_1),.din(w_dff_A_k1WU7RTL7_1),.clk(gclk));
	jdff dff_A_K2oUXlZz3_1(.dout(w_dff_A_k1WU7RTL7_1),.din(w_dff_A_K2oUXlZz3_1),.clk(gclk));
	jdff dff_A_A1DlU1gM0_1(.dout(w_dff_A_K2oUXlZz3_1),.din(w_dff_A_A1DlU1gM0_1),.clk(gclk));
	jdff dff_A_0ARvSZ8F9_1(.dout(w_dff_A_A1DlU1gM0_1),.din(w_dff_A_0ARvSZ8F9_1),.clk(gclk));
	jdff dff_A_GqUV8JKA9_0(.dout(w_G40gat_0[0]),.din(w_dff_A_GqUV8JKA9_0),.clk(gclk));
	jdff dff_A_48eaq5Ir5_0(.dout(w_dff_A_GqUV8JKA9_0),.din(w_dff_A_48eaq5Ir5_0),.clk(gclk));
	jdff dff_A_NvyiPqS37_0(.dout(w_dff_A_48eaq5Ir5_0),.din(w_dff_A_NvyiPqS37_0),.clk(gclk));
	jdff dff_A_wuz6Fc069_0(.dout(w_dff_A_NvyiPqS37_0),.din(w_dff_A_wuz6Fc069_0),.clk(gclk));
	jdff dff_A_B9lTBLGU4_0(.dout(w_dff_A_wuz6Fc069_0),.din(w_dff_A_B9lTBLGU4_0),.clk(gclk));
	jdff dff_A_r0oD3pQw5_0(.dout(w_dff_A_B9lTBLGU4_0),.din(w_dff_A_r0oD3pQw5_0),.clk(gclk));
	jdff dff_A_TXKiECU73_0(.dout(w_dff_A_r0oD3pQw5_0),.din(w_dff_A_TXKiECU73_0),.clk(gclk));
	jdff dff_A_mp9hLhBg7_0(.dout(w_dff_A_TXKiECU73_0),.din(w_dff_A_mp9hLhBg7_0),.clk(gclk));
	jdff dff_A_RhnNqOOW1_0(.dout(w_dff_A_mp9hLhBg7_0),.din(w_dff_A_RhnNqOOW1_0),.clk(gclk));
	jdff dff_A_sottCIB02_0(.dout(w_dff_A_RhnNqOOW1_0),.din(w_dff_A_sottCIB02_0),.clk(gclk));
	jdff dff_A_rwc6q2dn2_0(.dout(w_dff_A_sottCIB02_0),.din(w_dff_A_rwc6q2dn2_0),.clk(gclk));
	jdff dff_A_gxtiFyyH8_0(.dout(w_dff_A_rwc6q2dn2_0),.din(w_dff_A_gxtiFyyH8_0),.clk(gclk));
	jdff dff_A_xbnXnNeJ5_0(.dout(w_dff_A_gxtiFyyH8_0),.din(w_dff_A_xbnXnNeJ5_0),.clk(gclk));
	jdff dff_A_3vOkVf0c5_0(.dout(w_dff_A_xbnXnNeJ5_0),.din(w_dff_A_3vOkVf0c5_0),.clk(gclk));
	jdff dff_A_S9Y8jeJ59_0(.dout(w_dff_A_3vOkVf0c5_0),.din(w_dff_A_S9Y8jeJ59_0),.clk(gclk));
	jdff dff_A_2nMf8lIr9_1(.dout(w_n147_0[1]),.din(w_dff_A_2nMf8lIr9_1),.clk(gclk));
	jdff dff_B_hgRNJLr90_0(.din(n146),.dout(w_dff_B_hgRNJLr90_0),.clk(gclk));
	jdff dff_B_8toNLRwD6_0(.din(w_dff_B_hgRNJLr90_0),.dout(w_dff_B_8toNLRwD6_0),.clk(gclk));
	jdff dff_B_YrCFl0P75_0(.din(w_dff_B_8toNLRwD6_0),.dout(w_dff_B_YrCFl0P75_0),.clk(gclk));
	jdff dff_B_TXJwmJs32_0(.din(w_dff_B_YrCFl0P75_0),.dout(w_dff_B_TXJwmJs32_0),.clk(gclk));
	jdff dff_B_T6Rc6Deo2_0(.din(w_dff_B_TXJwmJs32_0),.dout(w_dff_B_T6Rc6Deo2_0),.clk(gclk));
	jdff dff_B_paiVXyJb5_0(.din(w_dff_B_T6Rc6Deo2_0),.dout(w_dff_B_paiVXyJb5_0),.clk(gclk));
	jdff dff_A_VDhjwMVA7_0(.dout(w_n145_0[0]),.din(w_dff_A_VDhjwMVA7_0),.clk(gclk));
	jdff dff_A_HCaIh7oj7_0(.dout(w_dff_A_VDhjwMVA7_0),.din(w_dff_A_HCaIh7oj7_0),.clk(gclk));
	jdff dff_A_N8jagXYC1_0(.dout(w_dff_A_HCaIh7oj7_0),.din(w_dff_A_N8jagXYC1_0),.clk(gclk));
	jdff dff_A_GCm9gLmv1_0(.dout(w_dff_A_N8jagXYC1_0),.din(w_dff_A_GCm9gLmv1_0),.clk(gclk));
	jdff dff_A_H3at82mu6_0(.dout(w_dff_A_GCm9gLmv1_0),.din(w_dff_A_H3at82mu6_0),.clk(gclk));
	jdff dff_A_pPnQxv1e3_0(.dout(w_dff_A_H3at82mu6_0),.din(w_dff_A_pPnQxv1e3_0),.clk(gclk));
	jdff dff_A_WDJJMe4c4_0(.dout(w_dff_A_pPnQxv1e3_0),.din(w_dff_A_WDJJMe4c4_0),.clk(gclk));
	jdff dff_A_zEsNOJXv9_0(.dout(w_dff_A_WDJJMe4c4_0),.din(w_dff_A_zEsNOJXv9_0),.clk(gclk));
	jdff dff_A_iajL2Dnv6_0(.dout(w_dff_A_zEsNOJXv9_0),.din(w_dff_A_iajL2Dnv6_0),.clk(gclk));
	jdff dff_A_ti2L8lQ49_0(.dout(w_dff_A_iajL2Dnv6_0),.din(w_dff_A_ti2L8lQ49_0),.clk(gclk));
	jdff dff_A_fy2ss3vq8_0(.dout(w_dff_A_ti2L8lQ49_0),.din(w_dff_A_fy2ss3vq8_0),.clk(gclk));
	jdff dff_A_O0wQlBzA7_0(.dout(w_dff_A_fy2ss3vq8_0),.din(w_dff_A_O0wQlBzA7_0),.clk(gclk));
	jdff dff_B_fzzC41Ff8_2(.din(n145),.dout(w_dff_B_fzzC41Ff8_2),.clk(gclk));
	jdff dff_B_SdaI9yDV7_2(.din(w_dff_B_fzzC41Ff8_2),.dout(w_dff_B_SdaI9yDV7_2),.clk(gclk));
	jdff dff_B_lVeuFj7i3_2(.din(w_dff_B_SdaI9yDV7_2),.dout(w_dff_B_lVeuFj7i3_2),.clk(gclk));
	jdff dff_B_l967Xkaa4_2(.din(w_dff_B_lVeuFj7i3_2),.dout(w_dff_B_l967Xkaa4_2),.clk(gclk));
	jdff dff_B_PgL5sdK07_2(.din(w_dff_B_l967Xkaa4_2),.dout(w_dff_B_PgL5sdK07_2),.clk(gclk));
	jdff dff_B_F5KTOii04_2(.din(w_dff_B_PgL5sdK07_2),.dout(w_dff_B_F5KTOii04_2),.clk(gclk));
	jdff dff_B_nRqDZMM19_2(.din(w_dff_B_F5KTOii04_2),.dout(w_dff_B_nRqDZMM19_2),.clk(gclk));
	jdff dff_A_ETQstGiG0_0(.dout(w_G53gat_0[0]),.din(w_dff_A_ETQstGiG0_0),.clk(gclk));
	jdff dff_A_zZbIzLg79_0(.dout(w_dff_A_ETQstGiG0_0),.din(w_dff_A_zZbIzLg79_0),.clk(gclk));
	jdff dff_A_DbGLIGMI4_0(.dout(w_dff_A_zZbIzLg79_0),.din(w_dff_A_DbGLIGMI4_0),.clk(gclk));
	jdff dff_A_pKRwmpZK3_0(.dout(w_dff_A_DbGLIGMI4_0),.din(w_dff_A_pKRwmpZK3_0),.clk(gclk));
	jdff dff_A_fhi3Q4gO4_0(.dout(w_dff_A_pKRwmpZK3_0),.din(w_dff_A_fhi3Q4gO4_0),.clk(gclk));
	jdff dff_A_2dwXvW6g6_0(.dout(w_dff_A_fhi3Q4gO4_0),.din(w_dff_A_2dwXvW6g6_0),.clk(gclk));
	jdff dff_A_E0sjAgrb3_0(.dout(w_dff_A_2dwXvW6g6_0),.din(w_dff_A_E0sjAgrb3_0),.clk(gclk));
	jdff dff_A_I1CYUHlT3_0(.dout(w_dff_A_E0sjAgrb3_0),.din(w_dff_A_I1CYUHlT3_0),.clk(gclk));
	jdff dff_A_KGSJOwy29_0(.dout(w_dff_A_I1CYUHlT3_0),.din(w_dff_A_KGSJOwy29_0),.clk(gclk));
	jdff dff_A_Hp1puBtR0_0(.dout(w_dff_A_KGSJOwy29_0),.din(w_dff_A_Hp1puBtR0_0),.clk(gclk));
	jdff dff_A_QlDhJh9o1_0(.dout(w_dff_A_Hp1puBtR0_0),.din(w_dff_A_QlDhJh9o1_0),.clk(gclk));
	jdff dff_A_15CWYWUg3_0(.dout(w_dff_A_QlDhJh9o1_0),.din(w_dff_A_15CWYWUg3_0),.clk(gclk));
	jdff dff_A_U5XpNZBA8_0(.dout(w_dff_A_15CWYWUg3_0),.din(w_dff_A_U5XpNZBA8_0),.clk(gclk));
	jdff dff_A_oTYYasxg4_0(.dout(w_dff_A_U5XpNZBA8_0),.din(w_dff_A_oTYYasxg4_0),.clk(gclk));
	jdff dff_A_tLUHc9pw8_0(.dout(w_dff_A_oTYYasxg4_0),.din(w_dff_A_tLUHc9pw8_0),.clk(gclk));
	jdff dff_A_Wispl0754_0(.dout(w_dff_A_tLUHc9pw8_0),.din(w_dff_A_Wispl0754_0),.clk(gclk));
	jdff dff_A_BJdJbONd7_0(.dout(w_dff_A_Wispl0754_0),.din(w_dff_A_BJdJbONd7_0),.clk(gclk));
	jdff dff_A_vB8S38w90_0(.dout(w_dff_A_BJdJbONd7_0),.din(w_dff_A_vB8S38w90_0),.clk(gclk));
	jdff dff_A_PjoCkbYc5_0(.dout(w_dff_A_vB8S38w90_0),.din(w_dff_A_PjoCkbYc5_0),.clk(gclk));
	jdff dff_A_nWrydaZy0_0(.dout(w_dff_A_PjoCkbYc5_0),.din(w_dff_A_nWrydaZy0_0),.clk(gclk));
	jdff dff_A_i11qy3oI3_0(.dout(w_n141_0[0]),.din(w_dff_A_i11qy3oI3_0),.clk(gclk));
	jdff dff_B_9Ejn8SAM9_1(.din(n124),.dout(w_dff_B_9Ejn8SAM9_1),.clk(gclk));
	jdff dff_B_b99rtdSG1_1(.din(n129),.dout(w_dff_B_b99rtdSG1_1),.clk(gclk));
	jdff dff_B_O81W0fyS3_1(.din(w_dff_B_b99rtdSG1_1),.dout(w_dff_B_O81W0fyS3_1),.clk(gclk));
	jdff dff_B_0ibJyFA01_1(.din(w_dff_B_O81W0fyS3_1),.dout(w_dff_B_0ibJyFA01_1),.clk(gclk));
	jdff dff_B_ZT584fq39_1(.din(w_dff_B_0ibJyFA01_1),.dout(w_dff_B_ZT584fq39_1),.clk(gclk));
	jdff dff_B_1YSV3hag4_1(.din(w_dff_B_ZT584fq39_1),.dout(w_dff_B_1YSV3hag4_1),.clk(gclk));
	jdff dff_B_wxeByVvQ8_1(.din(w_dff_B_1YSV3hag4_1),.dout(w_dff_B_wxeByVvQ8_1),.clk(gclk));
	jdff dff_B_JB9geFc13_1(.din(w_dff_B_wxeByVvQ8_1),.dout(w_dff_B_JB9geFc13_1),.clk(gclk));
	jdff dff_A_VbA1FYqv1_0(.dout(w_n131_0[0]),.din(w_dff_A_VbA1FYqv1_0),.clk(gclk));
	jdff dff_A_3zMzafxQ0_0(.dout(w_dff_A_VbA1FYqv1_0),.din(w_dff_A_3zMzafxQ0_0),.clk(gclk));
	jdff dff_A_7chVJTYT4_0(.dout(w_dff_A_3zMzafxQ0_0),.din(w_dff_A_7chVJTYT4_0),.clk(gclk));
	jdff dff_A_3lOcn6Ae6_0(.dout(w_dff_A_7chVJTYT4_0),.din(w_dff_A_3lOcn6Ae6_0),.clk(gclk));
	jdff dff_A_jRx41jlR4_0(.dout(w_dff_A_3lOcn6Ae6_0),.din(w_dff_A_jRx41jlR4_0),.clk(gclk));
	jdff dff_A_Iaa9LfoL2_0(.dout(w_dff_A_jRx41jlR4_0),.din(w_dff_A_Iaa9LfoL2_0),.clk(gclk));
	jdff dff_A_xlMAHoDw3_0(.dout(w_dff_A_Iaa9LfoL2_0),.din(w_dff_A_xlMAHoDw3_0),.clk(gclk));
	jdff dff_A_WtCqoIhw8_0(.dout(w_n127_0[0]),.din(w_dff_A_WtCqoIhw8_0),.clk(gclk));
	jdff dff_A_eMJEcvRX9_0(.dout(w_dff_A_WtCqoIhw8_0),.din(w_dff_A_eMJEcvRX9_0),.clk(gclk));
	jdff dff_A_6qyoy6ti4_0(.dout(w_dff_A_eMJEcvRX9_0),.din(w_dff_A_6qyoy6ti4_0),.clk(gclk));
	jdff dff_A_INV8YbR14_0(.dout(w_dff_A_6qyoy6ti4_0),.din(w_dff_A_INV8YbR14_0),.clk(gclk));
	jdff dff_A_QPC3tFcH5_0(.dout(w_dff_A_INV8YbR14_0),.din(w_dff_A_QPC3tFcH5_0),.clk(gclk));
	jdff dff_A_ulPa3Dcx5_0(.dout(w_dff_A_QPC3tFcH5_0),.din(w_dff_A_ulPa3Dcx5_0),.clk(gclk));
	jdff dff_A_mdg1Qcp65_0(.dout(w_n125_0[0]),.din(w_dff_A_mdg1Qcp65_0),.clk(gclk));
	jdff dff_A_XYS1mqVo8_0(.dout(w_dff_A_mdg1Qcp65_0),.din(w_dff_A_XYS1mqVo8_0),.clk(gclk));
	jdff dff_A_j6MGPAlk3_0(.dout(w_dff_A_XYS1mqVo8_0),.din(w_dff_A_j6MGPAlk3_0),.clk(gclk));
	jdff dff_A_f0KLnLm14_0(.dout(w_dff_A_j6MGPAlk3_0),.din(w_dff_A_f0KLnLm14_0),.clk(gclk));
	jdff dff_A_8KnHbGtN8_0(.dout(w_dff_A_f0KLnLm14_0),.din(w_dff_A_8KnHbGtN8_0),.clk(gclk));
	jdff dff_B_D3rm779A3_2(.din(n125),.dout(w_dff_B_D3rm779A3_2),.clk(gclk));
	jdff dff_B_VLsBj1Ob3_2(.din(w_dff_B_D3rm779A3_2),.dout(w_dff_B_VLsBj1Ob3_2),.clk(gclk));
	jdff dff_B_a3N31SVR7_2(.din(w_dff_B_VLsBj1Ob3_2),.dout(w_dff_B_a3N31SVR7_2),.clk(gclk));
	jdff dff_B_wRLyrwcF8_2(.din(w_dff_B_a3N31SVR7_2),.dout(w_dff_B_wRLyrwcF8_2),.clk(gclk));
	jdff dff_B_xxWt0xOr8_2(.din(w_dff_B_wRLyrwcF8_2),.dout(w_dff_B_xxWt0xOr8_2),.clk(gclk));
	jdff dff_B_0oOVepwL9_2(.din(w_dff_B_xxWt0xOr8_2),.dout(w_dff_B_0oOVepwL9_2),.clk(gclk));
	jdff dff_B_LjiddWGy7_2(.din(w_dff_B_0oOVepwL9_2),.dout(w_dff_B_LjiddWGy7_2),.clk(gclk));
	jdff dff_A_75b5ul9A3_0(.dout(w_n123_0[0]),.din(w_dff_A_75b5ul9A3_0),.clk(gclk));
	jdff dff_A_Hc0Amted6_0(.dout(w_dff_A_75b5ul9A3_0),.din(w_dff_A_Hc0Amted6_0),.clk(gclk));
	jdff dff_A_JR78ul7R6_0(.dout(w_dff_A_Hc0Amted6_0),.din(w_dff_A_JR78ul7R6_0),.clk(gclk));
	jdff dff_A_Vkbw9zmX5_0(.dout(w_dff_A_JR78ul7R6_0),.din(w_dff_A_Vkbw9zmX5_0),.clk(gclk));
	jdff dff_A_vxywRz2Y0_0(.dout(w_dff_A_Vkbw9zmX5_0),.din(w_dff_A_vxywRz2Y0_0),.clk(gclk));
	jdff dff_A_iXLtYgTW0_0(.dout(w_dff_A_vxywRz2Y0_0),.din(w_dff_A_iXLtYgTW0_0),.clk(gclk));
	jdff dff_A_HasXKJGy4_0(.dout(w_n121_0[0]),.din(w_dff_A_HasXKJGy4_0),.clk(gclk));
	jdff dff_A_8MlS1o3V7_0(.dout(w_dff_A_HasXKJGy4_0),.din(w_dff_A_8MlS1o3V7_0),.clk(gclk));
	jdff dff_A_dNA4oHAQ7_0(.dout(w_dff_A_8MlS1o3V7_0),.din(w_dff_A_dNA4oHAQ7_0),.clk(gclk));
	jdff dff_A_qFtG1D614_0(.dout(w_dff_A_dNA4oHAQ7_0),.din(w_dff_A_qFtG1D614_0),.clk(gclk));
	jdff dff_A_ZZTgA83A1_0(.dout(w_dff_A_qFtG1D614_0),.din(w_dff_A_ZZTgA83A1_0),.clk(gclk));
	jdff dff_B_s9JpqwuC2_2(.din(n121),.dout(w_dff_B_s9JpqwuC2_2),.clk(gclk));
	jdff dff_B_zjrwG2rx1_2(.din(w_dff_B_s9JpqwuC2_2),.dout(w_dff_B_zjrwG2rx1_2),.clk(gclk));
	jdff dff_B_vo65AGxd4_2(.din(w_dff_B_zjrwG2rx1_2),.dout(w_dff_B_vo65AGxd4_2),.clk(gclk));
	jdff dff_B_CDxLi0nf7_2(.din(w_dff_B_vo65AGxd4_2),.dout(w_dff_B_CDxLi0nf7_2),.clk(gclk));
	jdff dff_B_TOOniKQo0_2(.din(w_dff_B_CDxLi0nf7_2),.dout(w_dff_B_TOOniKQo0_2),.clk(gclk));
	jdff dff_B_sZxPAbMC2_2(.din(w_dff_B_TOOniKQo0_2),.dout(w_dff_B_sZxPAbMC2_2),.clk(gclk));
	jdff dff_B_2383nTjN5_2(.din(w_dff_B_sZxPAbMC2_2),.dout(w_dff_B_2383nTjN5_2),.clk(gclk));
	jdff dff_B_UuWpBk8e4_1(.din(n101),.dout(w_dff_B_UuWpBk8e4_1),.clk(gclk));
	jdff dff_B_5jEXFLQw6_0(.din(n114),.dout(w_dff_B_5jEXFLQw6_0),.clk(gclk));
	jdff dff_A_wD8pm91g9_0(.dout(w_n113_0[0]),.din(w_dff_A_wD8pm91g9_0),.clk(gclk));
	jdff dff_A_B6bWZbTF0_0(.dout(w_dff_A_wD8pm91g9_0),.din(w_dff_A_B6bWZbTF0_0),.clk(gclk));
	jdff dff_A_0MQiOCrZ5_0(.dout(w_dff_A_B6bWZbTF0_0),.din(w_dff_A_0MQiOCrZ5_0),.clk(gclk));
	jdff dff_A_t26TpBhl1_0(.dout(w_dff_A_0MQiOCrZ5_0),.din(w_dff_A_t26TpBhl1_0),.clk(gclk));
	jdff dff_A_3FgFJ1Ds0_0(.dout(w_dff_A_t26TpBhl1_0),.din(w_dff_A_3FgFJ1Ds0_0),.clk(gclk));
	jdff dff_A_dZUWnc8V7_0(.dout(w_dff_A_3FgFJ1Ds0_0),.din(w_dff_A_dZUWnc8V7_0),.clk(gclk));
	jdff dff_A_YYp97nOP6_0(.dout(w_n111_0[0]),.din(w_dff_A_YYp97nOP6_0),.clk(gclk));
	jdff dff_A_pHKS3yWJ1_0(.dout(w_dff_A_YYp97nOP6_0),.din(w_dff_A_pHKS3yWJ1_0),.clk(gclk));
	jdff dff_A_3bj74WQe9_0(.dout(w_dff_A_pHKS3yWJ1_0),.din(w_dff_A_3bj74WQe9_0),.clk(gclk));
	jdff dff_A_6ggCqFz20_0(.dout(w_dff_A_3bj74WQe9_0),.din(w_dff_A_6ggCqFz20_0),.clk(gclk));
	jdff dff_A_SlqBgjwD3_0(.dout(w_dff_A_6ggCqFz20_0),.din(w_dff_A_SlqBgjwD3_0),.clk(gclk));
	jdff dff_B_6DwJa8ak8_2(.din(n111),.dout(w_dff_B_6DwJa8ak8_2),.clk(gclk));
	jdff dff_B_zpb7GV5u3_2(.din(w_dff_B_6DwJa8ak8_2),.dout(w_dff_B_zpb7GV5u3_2),.clk(gclk));
	jdff dff_B_co8Qk23n1_2(.din(w_dff_B_zpb7GV5u3_2),.dout(w_dff_B_co8Qk23n1_2),.clk(gclk));
	jdff dff_B_q3JMA5Vy5_2(.din(w_dff_B_co8Qk23n1_2),.dout(w_dff_B_q3JMA5Vy5_2),.clk(gclk));
	jdff dff_B_iWkayhoz4_2(.din(w_dff_B_q3JMA5Vy5_2),.dout(w_dff_B_iWkayhoz4_2),.clk(gclk));
	jdff dff_B_cU3JyvQs4_2(.din(w_dff_B_iWkayhoz4_2),.dout(w_dff_B_cU3JyvQs4_2),.clk(gclk));
	jdff dff_B_d94g1jne5_2(.din(w_dff_B_cU3JyvQs4_2),.dout(w_dff_B_d94g1jne5_2),.clk(gclk));
	jdff dff_A_Wd71qjV00_0(.dout(w_n108_0[0]),.din(w_dff_A_Wd71qjV00_0),.clk(gclk));
	jdff dff_A_vBHMAZOb3_0(.dout(w_dff_A_Wd71qjV00_0),.din(w_dff_A_vBHMAZOb3_0),.clk(gclk));
	jdff dff_A_tf5nt8KM8_0(.dout(w_dff_A_vBHMAZOb3_0),.din(w_dff_A_tf5nt8KM8_0),.clk(gclk));
	jdff dff_A_wXORQXsF8_0(.dout(w_dff_A_tf5nt8KM8_0),.din(w_dff_A_wXORQXsF8_0),.clk(gclk));
	jdff dff_A_7m7OL1VZ1_0(.dout(w_dff_A_wXORQXsF8_0),.din(w_dff_A_7m7OL1VZ1_0),.clk(gclk));
	jdff dff_A_HfQCzGGO4_0(.dout(w_dff_A_7m7OL1VZ1_0),.din(w_dff_A_HfQCzGGO4_0),.clk(gclk));
	jdff dff_A_qdhEkhzh8_0(.dout(w_n106_0[0]),.din(w_dff_A_qdhEkhzh8_0),.clk(gclk));
	jdff dff_A_h7uXJ1Za4_0(.dout(w_dff_A_qdhEkhzh8_0),.din(w_dff_A_h7uXJ1Za4_0),.clk(gclk));
	jdff dff_A_HpukHOts3_0(.dout(w_dff_A_h7uXJ1Za4_0),.din(w_dff_A_HpukHOts3_0),.clk(gclk));
	jdff dff_A_Df2fqTGy2_0(.dout(w_dff_A_HpukHOts3_0),.din(w_dff_A_Df2fqTGy2_0),.clk(gclk));
	jdff dff_A_iVbpCoSB7_0(.dout(w_dff_A_Df2fqTGy2_0),.din(w_dff_A_iVbpCoSB7_0),.clk(gclk));
	jdff dff_B_3NJJVuIR5_2(.din(n106),.dout(w_dff_B_3NJJVuIR5_2),.clk(gclk));
	jdff dff_B_xrr3inuy9_2(.din(w_dff_B_3NJJVuIR5_2),.dout(w_dff_B_xrr3inuy9_2),.clk(gclk));
	jdff dff_B_lXatA0Gb7_2(.din(w_dff_B_xrr3inuy9_2),.dout(w_dff_B_lXatA0Gb7_2),.clk(gclk));
	jdff dff_B_Q7cnN83r4_2(.din(w_dff_B_lXatA0Gb7_2),.dout(w_dff_B_Q7cnN83r4_2),.clk(gclk));
	jdff dff_B_T48b5iB48_2(.din(w_dff_B_Q7cnN83r4_2),.dout(w_dff_B_T48b5iB48_2),.clk(gclk));
	jdff dff_B_lYBSgovx5_2(.din(w_dff_B_T48b5iB48_2),.dout(w_dff_B_lYBSgovx5_2),.clk(gclk));
	jdff dff_B_xZXqVwxy2_2(.din(w_dff_B_lYBSgovx5_2),.dout(w_dff_B_xZXqVwxy2_2),.clk(gclk));
	jdff dff_B_0djgFnjH6_1(.din(n97),.dout(w_dff_B_0djgFnjH6_1),.clk(gclk));
	jdff dff_B_2cWYEqb12_1(.din(w_dff_B_0djgFnjH6_1),.dout(w_dff_B_2cWYEqb12_1),.clk(gclk));
	jdff dff_B_fss9v9pb7_1(.din(w_dff_B_2cWYEqb12_1),.dout(w_dff_B_fss9v9pb7_1),.clk(gclk));
	jdff dff_B_tvSybPBs1_1(.din(w_dff_B_fss9v9pb7_1),.dout(w_dff_B_tvSybPBs1_1),.clk(gclk));
	jdff dff_B_Ylua8ZW21_1(.din(w_dff_B_tvSybPBs1_1),.dout(w_dff_B_Ylua8ZW21_1),.clk(gclk));
	jdff dff_B_z4KKWFh40_1(.din(w_dff_B_Ylua8ZW21_1),.dout(w_dff_B_z4KKWFh40_1),.clk(gclk));
	jdff dff_B_69IWdBfv7_1(.din(w_dff_B_z4KKWFh40_1),.dout(w_dff_B_69IWdBfv7_1),.clk(gclk));
	jdff dff_A_etusTHS08_0(.dout(w_n95_0[0]),.din(w_dff_A_etusTHS08_0),.clk(gclk));
	jdff dff_A_xSnmWATm5_0(.dout(w_dff_A_etusTHS08_0),.din(w_dff_A_xSnmWATm5_0),.clk(gclk));
	jdff dff_A_mtTomtmr4_0(.dout(w_dff_A_xSnmWATm5_0),.din(w_dff_A_mtTomtmr4_0),.clk(gclk));
	jdff dff_A_eC3ulkGY4_0(.dout(w_dff_A_mtTomtmr4_0),.din(w_dff_A_eC3ulkGY4_0),.clk(gclk));
	jdff dff_A_O7ir2tha6_0(.dout(w_dff_A_eC3ulkGY4_0),.din(w_dff_A_O7ir2tha6_0),.clk(gclk));
	jdff dff_A_zIBHdoei7_0(.dout(w_dff_A_O7ir2tha6_0),.din(w_dff_A_zIBHdoei7_0),.clk(gclk));
	jdff dff_A_5A7yxSpN6_0(.dout(w_n70_0[0]),.din(w_dff_A_5A7yxSpN6_0),.clk(gclk));
	jdff dff_A_z9HeE6j80_0(.dout(w_dff_A_5A7yxSpN6_0),.din(w_dff_A_z9HeE6j80_0),.clk(gclk));
	jdff dff_A_E2as1UsJ9_0(.dout(w_dff_A_z9HeE6j80_0),.din(w_dff_A_E2as1UsJ9_0),.clk(gclk));
	jdff dff_A_w5h8NoPN9_0(.dout(w_dff_A_E2as1UsJ9_0),.din(w_dff_A_w5h8NoPN9_0),.clk(gclk));
	jdff dff_A_Vpuez0BJ8_0(.dout(w_dff_A_w5h8NoPN9_0),.din(w_dff_A_Vpuez0BJ8_0),.clk(gclk));
	jdff dff_B_hvYkcC6P7_2(.din(n70),.dout(w_dff_B_hvYkcC6P7_2),.clk(gclk));
	jdff dff_B_bEFYQsCV1_2(.din(w_dff_B_hvYkcC6P7_2),.dout(w_dff_B_bEFYQsCV1_2),.clk(gclk));
	jdff dff_B_zPzNNgvb9_2(.din(w_dff_B_bEFYQsCV1_2),.dout(w_dff_B_zPzNNgvb9_2),.clk(gclk));
	jdff dff_B_jHY2UP930_2(.din(w_dff_B_zPzNNgvb9_2),.dout(w_dff_B_jHY2UP930_2),.clk(gclk));
	jdff dff_B_El9v8IRk6_2(.din(w_dff_B_jHY2UP930_2),.dout(w_dff_B_El9v8IRk6_2),.clk(gclk));
	jdff dff_B_svnRpbIj0_2(.din(w_dff_B_El9v8IRk6_2),.dout(w_dff_B_svnRpbIj0_2),.clk(gclk));
	jdff dff_B_zXMf2XEi9_2(.din(w_dff_B_svnRpbIj0_2),.dout(w_dff_B_zXMf2XEi9_2),.clk(gclk));
	jdff dff_A_yGXAjNQO9_1(.dout(w_G105gat_0[1]),.din(w_dff_A_yGXAjNQO9_1),.clk(gclk));
	jdff dff_A_hD07DT974_1(.dout(w_dff_A_yGXAjNQO9_1),.din(w_dff_A_hD07DT974_1),.clk(gclk));
	jdff dff_A_6y0FKlIA3_1(.dout(w_dff_A_hD07DT974_1),.din(w_dff_A_6y0FKlIA3_1),.clk(gclk));
	jdff dff_A_lzWotW326_1(.dout(w_dff_A_6y0FKlIA3_1),.din(w_dff_A_lzWotW326_1),.clk(gclk));
	jdff dff_A_U7C7JYPf9_1(.dout(w_dff_A_lzWotW326_1),.din(w_dff_A_U7C7JYPf9_1),.clk(gclk));
	jdff dff_A_tsHqbiwq9_1(.dout(w_dff_A_U7C7JYPf9_1),.din(w_dff_A_tsHqbiwq9_1),.clk(gclk));
	jdff dff_A_0TP2qSA35_1(.dout(w_dff_A_tsHqbiwq9_1),.din(w_dff_A_0TP2qSA35_1),.clk(gclk));
	jdff dff_A_Nhge5zT49_1(.dout(w_dff_A_0TP2qSA35_1),.din(w_dff_A_Nhge5zT49_1),.clk(gclk));
	jdff dff_A_btuvgOL03_1(.dout(w_dff_A_Nhge5zT49_1),.din(w_dff_A_btuvgOL03_1),.clk(gclk));
	jdff dff_A_s10MHrKl5_1(.dout(w_dff_A_btuvgOL03_1),.din(w_dff_A_s10MHrKl5_1),.clk(gclk));
	jdff dff_A_Y3y0ffj90_1(.dout(w_dff_A_s10MHrKl5_1),.din(w_dff_A_Y3y0ffj90_1),.clk(gclk));
	jdff dff_A_eri90pHm3_1(.dout(w_dff_A_Y3y0ffj90_1),.din(w_dff_A_eri90pHm3_1),.clk(gclk));
	jdff dff_A_veiJWYq83_1(.dout(w_dff_A_eri90pHm3_1),.din(w_dff_A_veiJWYq83_1),.clk(gclk));
	jdff dff_A_93LQLPH25_1(.dout(w_dff_A_veiJWYq83_1),.din(w_dff_A_93LQLPH25_1),.clk(gclk));
	jdff dff_A_H0izGr0v9_1(.dout(w_dff_A_93LQLPH25_1),.din(w_dff_A_H0izGr0v9_1),.clk(gclk));
	jdff dff_A_pWDz6cub2_0(.dout(w_n200_0[0]),.din(w_dff_A_pWDz6cub2_0),.clk(gclk));
	jdff dff_A_XgPVrpW43_0(.dout(w_dff_A_pWDz6cub2_0),.din(w_dff_A_XgPVrpW43_0),.clk(gclk));
	jdff dff_A_kqq7ADov6_0(.dout(w_dff_A_XgPVrpW43_0),.din(w_dff_A_kqq7ADov6_0),.clk(gclk));
	jdff dff_A_inpDNTQ21_0(.dout(w_dff_A_kqq7ADov6_0),.din(w_dff_A_inpDNTQ21_0),.clk(gclk));
	jdff dff_A_QSBh61bw9_0(.dout(w_dff_A_inpDNTQ21_0),.din(w_dff_A_QSBh61bw9_0),.clk(gclk));
	jdff dff_B_ByfiAHEG9_2(.din(n200),.dout(w_dff_B_ByfiAHEG9_2),.clk(gclk));
	jdff dff_B_yebf95lj0_2(.din(w_dff_B_ByfiAHEG9_2),.dout(w_dff_B_yebf95lj0_2),.clk(gclk));
	jdff dff_B_4P4Dj14L1_2(.din(w_dff_B_yebf95lj0_2),.dout(w_dff_B_4P4Dj14L1_2),.clk(gclk));
	jdff dff_B_2rPpI94R8_2(.din(w_dff_B_4P4Dj14L1_2),.dout(w_dff_B_2rPpI94R8_2),.clk(gclk));
	jdff dff_B_3Ld2ROdY9_2(.din(w_dff_B_2rPpI94R8_2),.dout(w_dff_B_3Ld2ROdY9_2),.clk(gclk));
	jdff dff_B_MjrbvAuh6_2(.din(w_dff_B_3Ld2ROdY9_2),.dout(w_dff_B_MjrbvAuh6_2),.clk(gclk));
	jdff dff_B_drRRZsue3_2(.din(w_dff_B_MjrbvAuh6_2),.dout(w_dff_B_drRRZsue3_2),.clk(gclk));
	jdff dff_B_MJhrWLMi7_2(.din(w_dff_B_drRRZsue3_2),.dout(w_dff_B_MJhrWLMi7_2),.clk(gclk));
	jdff dff_B_cObmXuED5_2(.din(w_dff_B_MJhrWLMi7_2),.dout(w_dff_B_cObmXuED5_2),.clk(gclk));
	jdff dff_B_8VuazdCD8_2(.din(w_dff_B_cObmXuED5_2),.dout(w_dff_B_8VuazdCD8_2),.clk(gclk));
	jdff dff_B_k2SiN4JA2_2(.din(w_dff_B_8VuazdCD8_2),.dout(w_dff_B_k2SiN4JA2_2),.clk(gclk));
	jdff dff_B_bqYDk4FS7_2(.din(w_dff_B_k2SiN4JA2_2),.dout(w_dff_B_bqYDk4FS7_2),.clk(gclk));
	jdff dff_B_X44NYGyM9_2(.din(w_dff_B_bqYDk4FS7_2),.dout(w_dff_B_X44NYGyM9_2),.clk(gclk));
	jdff dff_B_zxrmMO796_2(.din(w_dff_B_X44NYGyM9_2),.dout(w_dff_B_zxrmMO796_2),.clk(gclk));
	jdff dff_A_gaYOyXy37_0(.dout(w_G79gat_0[0]),.din(w_dff_A_gaYOyXy37_0),.clk(gclk));
	jdff dff_A_Mjlub2SV9_0(.dout(w_dff_A_gaYOyXy37_0),.din(w_dff_A_Mjlub2SV9_0),.clk(gclk));
	jdff dff_A_8RjYcBBN2_0(.dout(w_dff_A_Mjlub2SV9_0),.din(w_dff_A_8RjYcBBN2_0),.clk(gclk));
	jdff dff_A_MkCc97db5_0(.dout(w_dff_A_8RjYcBBN2_0),.din(w_dff_A_MkCc97db5_0),.clk(gclk));
	jdff dff_A_hfzKUSQM4_0(.dout(w_dff_A_MkCc97db5_0),.din(w_dff_A_hfzKUSQM4_0),.clk(gclk));
	jdff dff_A_KUzs6dp26_0(.dout(w_dff_A_hfzKUSQM4_0),.din(w_dff_A_KUzs6dp26_0),.clk(gclk));
	jdff dff_A_itPQSgbR6_0(.dout(w_dff_A_KUzs6dp26_0),.din(w_dff_A_itPQSgbR6_0),.clk(gclk));
	jdff dff_A_0XbUR4kT0_0(.dout(w_dff_A_itPQSgbR6_0),.din(w_dff_A_0XbUR4kT0_0),.clk(gclk));
	jdff dff_A_ICPe4uHu8_0(.dout(w_dff_A_0XbUR4kT0_0),.din(w_dff_A_ICPe4uHu8_0),.clk(gclk));
	jdff dff_A_35SPAG2C1_0(.dout(w_dff_A_ICPe4uHu8_0),.din(w_dff_A_35SPAG2C1_0),.clk(gclk));
	jdff dff_A_HXJgagCy8_0(.dout(w_dff_A_35SPAG2C1_0),.din(w_dff_A_HXJgagCy8_0),.clk(gclk));
	jdff dff_A_WHHALaDU3_0(.dout(w_dff_A_HXJgagCy8_0),.din(w_dff_A_WHHALaDU3_0),.clk(gclk));
	jdff dff_A_n57mvHM27_0(.dout(w_dff_A_WHHALaDU3_0),.din(w_dff_A_n57mvHM27_0),.clk(gclk));
	jdff dff_A_EZ7PtoxU8_0(.dout(w_dff_A_n57mvHM27_0),.din(w_dff_A_EZ7PtoxU8_0),.clk(gclk));
	jdff dff_A_4Hbif21O6_0(.dout(w_dff_A_EZ7PtoxU8_0),.din(w_dff_A_4Hbif21O6_0),.clk(gclk));
	jdff dff_A_vWsW9iQT5_0(.dout(w_n202_0[0]),.din(w_dff_A_vWsW9iQT5_0),.clk(gclk));
	jdff dff_A_vEY9DlgU3_0(.dout(w_dff_A_vWsW9iQT5_0),.din(w_dff_A_vEY9DlgU3_0),.clk(gclk));
	jdff dff_A_zqEVtEAi9_0(.dout(w_dff_A_vEY9DlgU3_0),.din(w_dff_A_zqEVtEAi9_0),.clk(gclk));
	jdff dff_A_hDvUd3Kn1_0(.dout(w_dff_A_zqEVtEAi9_0),.din(w_dff_A_hDvUd3Kn1_0),.clk(gclk));
	jdff dff_A_Y0v3swMy4_0(.dout(w_dff_A_hDvUd3Kn1_0),.din(w_dff_A_Y0v3swMy4_0),.clk(gclk));
	jdff dff_A_sH5qWaTd4_0(.dout(w_dff_A_Y0v3swMy4_0),.din(w_dff_A_sH5qWaTd4_0),.clk(gclk));
	jdff dff_B_SDhLMKyS7_1(.din(n168),.dout(w_dff_B_SDhLMKyS7_1),.clk(gclk));
	jdff dff_B_xhPinsnU9_1(.din(n171),.dout(w_dff_B_xhPinsnU9_1),.clk(gclk));
	jdff dff_A_bwF9LVaO1_0(.dout(w_G47gat_0[0]),.din(w_dff_A_bwF9LVaO1_0),.clk(gclk));
	jdff dff_A_kQKLUrFv0_0(.dout(w_dff_A_bwF9LVaO1_0),.din(w_dff_A_kQKLUrFv0_0),.clk(gclk));
	jdff dff_A_i6lNTESq6_0(.dout(w_dff_A_kQKLUrFv0_0),.din(w_dff_A_i6lNTESq6_0),.clk(gclk));
	jdff dff_A_90rAaKG98_0(.dout(w_dff_A_i6lNTESq6_0),.din(w_dff_A_90rAaKG98_0),.clk(gclk));
	jdff dff_A_OlIjdwvL0_0(.dout(w_dff_A_90rAaKG98_0),.din(w_dff_A_OlIjdwvL0_0),.clk(gclk));
	jdff dff_A_8MfW7LCP6_0(.dout(w_dff_A_OlIjdwvL0_0),.din(w_dff_A_8MfW7LCP6_0),.clk(gclk));
	jdff dff_A_oQ31W50A7_0(.dout(w_dff_A_8MfW7LCP6_0),.din(w_dff_A_oQ31W50A7_0),.clk(gclk));
	jdff dff_A_PNAk39HP3_0(.dout(w_dff_A_oQ31W50A7_0),.din(w_dff_A_PNAk39HP3_0),.clk(gclk));
	jdff dff_A_5EYzQs590_1(.dout(w_G47gat_0[1]),.din(w_dff_A_5EYzQs590_1),.clk(gclk));
	jdff dff_A_ixdHPJ1C3_1(.dout(w_dff_A_5EYzQs590_1),.din(w_dff_A_ixdHPJ1C3_1),.clk(gclk));
	jdff dff_A_UF9pdw1g6_1(.dout(w_dff_A_ixdHPJ1C3_1),.din(w_dff_A_UF9pdw1g6_1),.clk(gclk));
	jdff dff_A_vNj5IGle3_1(.dout(w_dff_A_UF9pdw1g6_1),.din(w_dff_A_vNj5IGle3_1),.clk(gclk));
	jdff dff_A_E1ZEBn9q1_1(.dout(w_dff_A_vNj5IGle3_1),.din(w_dff_A_E1ZEBn9q1_1),.clk(gclk));
	jdff dff_A_aEg1lPsR1_1(.dout(w_dff_A_E1ZEBn9q1_1),.din(w_dff_A_aEg1lPsR1_1),.clk(gclk));
	jdff dff_A_Zf9CVxiy8_1(.dout(w_dff_A_aEg1lPsR1_1),.din(w_dff_A_Zf9CVxiy8_1),.clk(gclk));
	jdff dff_A_xG03RLPb7_1(.dout(w_dff_A_Zf9CVxiy8_1),.din(w_dff_A_xG03RLPb7_1),.clk(gclk));
	jdff dff_A_rfXJqbez5_1(.dout(w_dff_A_xG03RLPb7_1),.din(w_dff_A_rfXJqbez5_1),.clk(gclk));
	jdff dff_A_n7eXfFcT5_1(.dout(w_dff_A_rfXJqbez5_1),.din(w_dff_A_n7eXfFcT5_1),.clk(gclk));
	jdff dff_A_ET9R53Hk4_1(.dout(w_dff_A_n7eXfFcT5_1),.din(w_dff_A_ET9R53Hk4_1),.clk(gclk));
	jdff dff_A_tQ1hlDZD4_1(.dout(w_dff_A_ET9R53Hk4_1),.din(w_dff_A_tQ1hlDZD4_1),.clk(gclk));
	jdff dff_A_wKWGJvJL1_1(.dout(w_dff_A_tQ1hlDZD4_1),.din(w_dff_A_wKWGJvJL1_1),.clk(gclk));
	jdff dff_A_yfnhmTCl5_0(.dout(w_n173_0[0]),.din(w_dff_A_yfnhmTCl5_0),.clk(gclk));
	jdff dff_A_g8narcgG7_0(.dout(w_dff_A_yfnhmTCl5_0),.din(w_dff_A_g8narcgG7_0),.clk(gclk));
	jdff dff_A_cEMPf0c93_0(.dout(w_dff_A_g8narcgG7_0),.din(w_dff_A_cEMPf0c93_0),.clk(gclk));
	jdff dff_A_F5ALTxrE4_0(.dout(w_dff_A_cEMPf0c93_0),.din(w_dff_A_F5ALTxrE4_0),.clk(gclk));
	jdff dff_A_9mhHPHMj0_0(.dout(w_dff_A_F5ALTxrE4_0),.din(w_dff_A_9mhHPHMj0_0),.clk(gclk));
	jdff dff_A_I1Wv4zCs2_0(.dout(w_dff_A_9mhHPHMj0_0),.din(w_dff_A_I1Wv4zCs2_0),.clk(gclk));
	jdff dff_A_7gXa9zaa1_0(.dout(w_G8gat_0[0]),.din(w_dff_A_7gXa9zaa1_0),.clk(gclk));
	jdff dff_A_jSH4mWPk3_0(.dout(w_dff_A_7gXa9zaa1_0),.din(w_dff_A_jSH4mWPk3_0),.clk(gclk));
	jdff dff_A_Cb8WFyt35_0(.dout(w_dff_A_jSH4mWPk3_0),.din(w_dff_A_Cb8WFyt35_0),.clk(gclk));
	jdff dff_A_Af1YuSND4_0(.dout(w_dff_A_Cb8WFyt35_0),.din(w_dff_A_Af1YuSND4_0),.clk(gclk));
	jdff dff_A_7cD3xAYU8_0(.dout(w_dff_A_Af1YuSND4_0),.din(w_dff_A_7cD3xAYU8_0),.clk(gclk));
	jdff dff_A_pgLAn1sp3_0(.dout(w_dff_A_7cD3xAYU8_0),.din(w_dff_A_pgLAn1sp3_0),.clk(gclk));
	jdff dff_A_uox7brt46_0(.dout(w_dff_A_pgLAn1sp3_0),.din(w_dff_A_uox7brt46_0),.clk(gclk));
	jdff dff_A_s2qg08bX5_0(.dout(w_dff_A_uox7brt46_0),.din(w_dff_A_s2qg08bX5_0),.clk(gclk));
	jdff dff_A_CV8VZeWM0_0(.dout(w_dff_A_s2qg08bX5_0),.din(w_dff_A_CV8VZeWM0_0),.clk(gclk));
	jdff dff_A_ejGkuxo42_0(.dout(w_dff_A_CV8VZeWM0_0),.din(w_dff_A_ejGkuxo42_0),.clk(gclk));
	jdff dff_A_sHFDSFSc4_0(.dout(w_dff_A_ejGkuxo42_0),.din(w_dff_A_sHFDSFSc4_0),.clk(gclk));
	jdff dff_A_b5MePVBU6_0(.dout(w_dff_A_sHFDSFSc4_0),.din(w_dff_A_b5MePVBU6_0),.clk(gclk));
	jdff dff_A_22AEj7LU2_0(.dout(w_dff_A_b5MePVBU6_0),.din(w_dff_A_22AEj7LU2_0),.clk(gclk));
	jdff dff_A_vCaMbch46_1(.dout(w_G8gat_0[1]),.din(w_dff_A_vCaMbch46_1),.clk(gclk));
	jdff dff_A_fbLuwnPe8_1(.dout(w_dff_A_vCaMbch46_1),.din(w_dff_A_fbLuwnPe8_1),.clk(gclk));
	jdff dff_A_r8IsYw6s7_1(.dout(w_dff_A_fbLuwnPe8_1),.din(w_dff_A_r8IsYw6s7_1),.clk(gclk));
	jdff dff_A_mbUctylG5_1(.dout(w_dff_A_r8IsYw6s7_1),.din(w_dff_A_mbUctylG5_1),.clk(gclk));
	jdff dff_A_ToATTP9q1_1(.dout(w_dff_A_mbUctylG5_1),.din(w_dff_A_ToATTP9q1_1),.clk(gclk));
	jdff dff_A_6knYgbo40_1(.dout(w_dff_A_ToATTP9q1_1),.din(w_dff_A_6knYgbo40_1),.clk(gclk));
	jdff dff_A_uKFuaD5e9_1(.dout(w_dff_A_6knYgbo40_1),.din(w_dff_A_uKFuaD5e9_1),.clk(gclk));
	jdff dff_A_jKSTLNsP8_1(.dout(w_dff_A_uKFuaD5e9_1),.din(w_dff_A_jKSTLNsP8_1),.clk(gclk));
	jdff dff_A_SvvGCQpD9_0(.dout(w_n170_0[0]),.din(w_dff_A_SvvGCQpD9_0),.clk(gclk));
	jdff dff_A_DJpB76TI8_0(.dout(w_dff_A_SvvGCQpD9_0),.din(w_dff_A_DJpB76TI8_0),.clk(gclk));
	jdff dff_A_ZTRatxce3_0(.dout(w_dff_A_DJpB76TI8_0),.din(w_dff_A_ZTRatxce3_0),.clk(gclk));
	jdff dff_A_R2fQV0xr7_0(.dout(w_dff_A_ZTRatxce3_0),.din(w_dff_A_R2fQV0xr7_0),.clk(gclk));
	jdff dff_A_8x7MykNQ2_0(.dout(w_dff_A_R2fQV0xr7_0),.din(w_dff_A_8x7MykNQ2_0),.clk(gclk));
	jdff dff_A_RIKbZ0pK9_0(.dout(w_dff_A_8x7MykNQ2_0),.din(w_dff_A_RIKbZ0pK9_0),.clk(gclk));
	jdff dff_A_Jndz8GqG8_0(.dout(w_G86gat_0[0]),.din(w_dff_A_Jndz8GqG8_0),.clk(gclk));
	jdff dff_A_4knAMhm52_0(.dout(w_dff_A_Jndz8GqG8_0),.din(w_dff_A_4knAMhm52_0),.clk(gclk));
	jdff dff_A_PhVqGSUi3_0(.dout(w_dff_A_4knAMhm52_0),.din(w_dff_A_PhVqGSUi3_0),.clk(gclk));
	jdff dff_A_3KDphlJv9_0(.dout(w_dff_A_PhVqGSUi3_0),.din(w_dff_A_3KDphlJv9_0),.clk(gclk));
	jdff dff_A_LFVeGlqI9_0(.dout(w_dff_A_3KDphlJv9_0),.din(w_dff_A_LFVeGlqI9_0),.clk(gclk));
	jdff dff_A_QO8QSwik2_0(.dout(w_dff_A_LFVeGlqI9_0),.din(w_dff_A_QO8QSwik2_0),.clk(gclk));
	jdff dff_A_qm0W7TaO1_0(.dout(w_dff_A_QO8QSwik2_0),.din(w_dff_A_qm0W7TaO1_0),.clk(gclk));
	jdff dff_A_XUgkw1wy5_0(.dout(w_dff_A_qm0W7TaO1_0),.din(w_dff_A_XUgkw1wy5_0),.clk(gclk));
	jdff dff_A_eRpb26Ny0_0(.dout(w_dff_A_XUgkw1wy5_0),.din(w_dff_A_eRpb26Ny0_0),.clk(gclk));
	jdff dff_A_KSlA7fia0_0(.dout(w_dff_A_eRpb26Ny0_0),.din(w_dff_A_KSlA7fia0_0),.clk(gclk));
	jdff dff_A_KuQL11Dh4_0(.dout(w_dff_A_KSlA7fia0_0),.din(w_dff_A_KuQL11Dh4_0),.clk(gclk));
	jdff dff_A_hjmAjkzM8_0(.dout(w_dff_A_KuQL11Dh4_0),.din(w_dff_A_hjmAjkzM8_0),.clk(gclk));
	jdff dff_A_a8rZTlo97_0(.dout(w_dff_A_hjmAjkzM8_0),.din(w_dff_A_a8rZTlo97_0),.clk(gclk));
	jdff dff_A_4jBlvItX0_1(.dout(w_G86gat_0[1]),.din(w_dff_A_4jBlvItX0_1),.clk(gclk));
	jdff dff_A_4lh03M5a6_1(.dout(w_dff_A_4jBlvItX0_1),.din(w_dff_A_4lh03M5a6_1),.clk(gclk));
	jdff dff_A_seaIE4A83_1(.dout(w_dff_A_4lh03M5a6_1),.din(w_dff_A_seaIE4A83_1),.clk(gclk));
	jdff dff_A_rpIXkCx68_1(.dout(w_dff_A_seaIE4A83_1),.din(w_dff_A_rpIXkCx68_1),.clk(gclk));
	jdff dff_A_g7R3sdOn7_1(.dout(w_dff_A_rpIXkCx68_1),.din(w_dff_A_g7R3sdOn7_1),.clk(gclk));
	jdff dff_A_xIUS5okl1_1(.dout(w_dff_A_g7R3sdOn7_1),.din(w_dff_A_xIUS5okl1_1),.clk(gclk));
	jdff dff_A_hMgvqrlX6_1(.dout(w_dff_A_xIUS5okl1_1),.din(w_dff_A_hMgvqrlX6_1),.clk(gclk));
	jdff dff_A_e7w7KJmh4_1(.dout(w_dff_A_hMgvqrlX6_1),.din(w_dff_A_e7w7KJmh4_1),.clk(gclk));
	jdff dff_A_quDyM02J4_1(.dout(w_n120_0[1]),.din(w_dff_A_quDyM02J4_1),.clk(gclk));
	jdff dff_A_bNchDfR86_1(.dout(w_dff_A_quDyM02J4_1),.din(w_dff_A_bNchDfR86_1),.clk(gclk));
	jdff dff_A_sx1E2CEi3_1(.dout(w_n119_0[1]),.din(w_dff_A_sx1E2CEi3_1),.clk(gclk));
	jdff dff_A_Oe3fGkx99_1(.dout(w_dff_A_sx1E2CEi3_1),.din(w_dff_A_Oe3fGkx99_1),.clk(gclk));
	jdff dff_A_j5ZFPF3W7_1(.dout(w_dff_A_Oe3fGkx99_1),.din(w_dff_A_j5ZFPF3W7_1),.clk(gclk));
	jdff dff_A_dJET2pmo5_1(.dout(w_dff_A_j5ZFPF3W7_1),.din(w_dff_A_dJET2pmo5_1),.clk(gclk));
	jdff dff_A_HsOYiziO0_1(.dout(w_dff_A_dJET2pmo5_1),.din(w_dff_A_HsOYiziO0_1),.clk(gclk));
	jdff dff_A_q34n06QX0_1(.dout(w_dff_A_HsOYiziO0_1),.din(w_dff_A_q34n06QX0_1),.clk(gclk));
	jdff dff_A_Kjwjci5j6_0(.dout(w_n117_0[0]),.din(w_dff_A_Kjwjci5j6_0),.clk(gclk));
	jdff dff_A_z9Sk57lB4_0(.dout(w_dff_A_Kjwjci5j6_0),.din(w_dff_A_z9Sk57lB4_0),.clk(gclk));
	jdff dff_A_z6wjh8qw1_0(.dout(w_dff_A_z9Sk57lB4_0),.din(w_dff_A_z6wjh8qw1_0),.clk(gclk));
	jdff dff_A_J19xxwDj7_0(.dout(w_dff_A_z6wjh8qw1_0),.din(w_dff_A_J19xxwDj7_0),.clk(gclk));
	jdff dff_A_6OkFu1Y69_0(.dout(w_dff_A_J19xxwDj7_0),.din(w_dff_A_6OkFu1Y69_0),.clk(gclk));
	jdff dff_B_FE8oe3zt8_2(.din(n117),.dout(w_dff_B_FE8oe3zt8_2),.clk(gclk));
	jdff dff_B_AuojKlfi3_2(.din(w_dff_B_FE8oe3zt8_2),.dout(w_dff_B_AuojKlfi3_2),.clk(gclk));
	jdff dff_B_q2orjG034_2(.din(w_dff_B_AuojKlfi3_2),.dout(w_dff_B_q2orjG034_2),.clk(gclk));
	jdff dff_B_C6p35jO67_2(.din(w_dff_B_q2orjG034_2),.dout(w_dff_B_C6p35jO67_2),.clk(gclk));
	jdff dff_B_yASvzsua5_2(.din(w_dff_B_C6p35jO67_2),.dout(w_dff_B_yASvzsua5_2),.clk(gclk));
	jdff dff_B_kr0qIfqT7_2(.din(w_dff_B_yASvzsua5_2),.dout(w_dff_B_kr0qIfqT7_2),.clk(gclk));
	jdff dff_B_6F2pPsVZ8_2(.din(w_dff_B_kr0qIfqT7_2),.dout(w_dff_B_6F2pPsVZ8_2),.clk(gclk));
	jdff dff_A_DKireuJq5_0(.dout(w_G60gat_0[0]),.din(w_dff_A_DKireuJq5_0),.clk(gclk));
	jdff dff_A_RDgVdBHK9_0(.dout(w_dff_A_DKireuJq5_0),.din(w_dff_A_RDgVdBHK9_0),.clk(gclk));
	jdff dff_A_luwGQRjV3_0(.dout(w_dff_A_RDgVdBHK9_0),.din(w_dff_A_luwGQRjV3_0),.clk(gclk));
	jdff dff_A_M9DGxWoU6_0(.dout(w_dff_A_luwGQRjV3_0),.din(w_dff_A_M9DGxWoU6_0),.clk(gclk));
	jdff dff_A_NU7gXzoF7_0(.dout(w_dff_A_M9DGxWoU6_0),.din(w_dff_A_NU7gXzoF7_0),.clk(gclk));
	jdff dff_A_jtd3syVZ6_0(.dout(w_dff_A_NU7gXzoF7_0),.din(w_dff_A_jtd3syVZ6_0),.clk(gclk));
	jdff dff_A_4lfgGwHj0_0(.dout(w_dff_A_jtd3syVZ6_0),.din(w_dff_A_4lfgGwHj0_0),.clk(gclk));
	jdff dff_A_6pkMR3F53_0(.dout(w_dff_A_4lfgGwHj0_0),.din(w_dff_A_6pkMR3F53_0),.clk(gclk));
	jdff dff_A_VOCbAonh0_0(.dout(w_dff_A_6pkMR3F53_0),.din(w_dff_A_VOCbAonh0_0),.clk(gclk));
	jdff dff_A_XTmcFUYU3_0(.dout(w_dff_A_VOCbAonh0_0),.din(w_dff_A_XTmcFUYU3_0),.clk(gclk));
	jdff dff_A_GTkSVVkd9_0(.dout(w_dff_A_XTmcFUYU3_0),.din(w_dff_A_GTkSVVkd9_0),.clk(gclk));
	jdff dff_A_WJS91CqH3_0(.dout(w_dff_A_GTkSVVkd9_0),.din(w_dff_A_WJS91CqH3_0),.clk(gclk));
	jdff dff_A_YG8qQCjJ1_0(.dout(w_dff_A_WJS91CqH3_0),.din(w_dff_A_YG8qQCjJ1_0),.clk(gclk));
	jdff dff_B_L4jdTIV36_1(.din(n154),.dout(w_dff_B_L4jdTIV36_1),.clk(gclk));
	jdff dff_B_LS2NnnOg9_0(.din(n165),.dout(w_dff_B_LS2NnnOg9_0),.clk(gclk));
	jdff dff_A_da2wEK4W8_0(.dout(w_n164_0[0]),.din(w_dff_A_da2wEK4W8_0),.clk(gclk));
	jdff dff_A_Go4Hd8746_0(.dout(w_dff_A_da2wEK4W8_0),.din(w_dff_A_Go4Hd8746_0),.clk(gclk));
	jdff dff_A_WBgjazlO6_0(.dout(w_dff_A_Go4Hd8746_0),.din(w_dff_A_WBgjazlO6_0),.clk(gclk));
	jdff dff_A_oVj8N9zX5_0(.dout(w_dff_A_WBgjazlO6_0),.din(w_dff_A_oVj8N9zX5_0),.clk(gclk));
	jdff dff_A_SiTL53oB4_0(.dout(w_dff_A_oVj8N9zX5_0),.din(w_dff_A_SiTL53oB4_0),.clk(gclk));
	jdff dff_A_0nTKHlM67_0(.dout(w_dff_A_SiTL53oB4_0),.din(w_dff_A_0nTKHlM67_0),.clk(gclk));
	jdff dff_B_mqLTv3ku5_1(.din(n162),.dout(w_dff_B_mqLTv3ku5_1),.clk(gclk));
	jdff dff_B_hlQwySnz8_1(.din(w_dff_B_mqLTv3ku5_1),.dout(w_dff_B_hlQwySnz8_1),.clk(gclk));
	jdff dff_B_9ZGB8oOo6_1(.din(w_dff_B_hlQwySnz8_1),.dout(w_dff_B_9ZGB8oOo6_1),.clk(gclk));
	jdff dff_B_TkvD2zrK6_1(.din(w_dff_B_9ZGB8oOo6_1),.dout(w_dff_B_TkvD2zrK6_1),.clk(gclk));
	jdff dff_B_MR1RBrVa4_1(.din(w_dff_B_TkvD2zrK6_1),.dout(w_dff_B_MR1RBrVa4_1),.clk(gclk));
	jdff dff_B_BOWiELq69_1(.din(w_dff_B_MR1RBrVa4_1),.dout(w_dff_B_BOWiELq69_1),.clk(gclk));
	jdff dff_A_RwybG6tX0_0(.dout(w_G112gat_0[0]),.din(w_dff_A_RwybG6tX0_0),.clk(gclk));
	jdff dff_A_LQDAvEqQ9_0(.dout(w_dff_A_RwybG6tX0_0),.din(w_dff_A_LQDAvEqQ9_0),.clk(gclk));
	jdff dff_A_XhwvFi4t7_0(.dout(w_dff_A_LQDAvEqQ9_0),.din(w_dff_A_XhwvFi4t7_0),.clk(gclk));
	jdff dff_A_iQfPExlA8_0(.dout(w_dff_A_XhwvFi4t7_0),.din(w_dff_A_iQfPExlA8_0),.clk(gclk));
	jdff dff_A_H04Op4pX0_0(.dout(w_dff_A_iQfPExlA8_0),.din(w_dff_A_H04Op4pX0_0),.clk(gclk));
	jdff dff_A_T5dfnjWx3_0(.dout(w_dff_A_H04Op4pX0_0),.din(w_dff_A_T5dfnjWx3_0),.clk(gclk));
	jdff dff_A_P0Cvhqf03_0(.dout(w_dff_A_T5dfnjWx3_0),.din(w_dff_A_P0Cvhqf03_0),.clk(gclk));
	jdff dff_A_FgQvTQOT0_0(.dout(w_dff_A_P0Cvhqf03_0),.din(w_dff_A_FgQvTQOT0_0),.clk(gclk));
	jdff dff_A_ht2VrqHN6_0(.dout(w_dff_A_FgQvTQOT0_0),.din(w_dff_A_ht2VrqHN6_0),.clk(gclk));
	jdff dff_A_QjYuXeHI0_0(.dout(w_dff_A_ht2VrqHN6_0),.din(w_dff_A_QjYuXeHI0_0),.clk(gclk));
	jdff dff_A_ml1kpYNG4_0(.dout(w_dff_A_QjYuXeHI0_0),.din(w_dff_A_ml1kpYNG4_0),.clk(gclk));
	jdff dff_A_9c1ceGrW5_0(.dout(w_dff_A_ml1kpYNG4_0),.din(w_dff_A_9c1ceGrW5_0),.clk(gclk));
	jdff dff_A_Trkf7w596_0(.dout(w_dff_A_9c1ceGrW5_0),.din(w_dff_A_Trkf7w596_0),.clk(gclk));
	jdff dff_A_wDrIAQlP5_1(.dout(w_G112gat_0[1]),.din(w_dff_A_wDrIAQlP5_1),.clk(gclk));
	jdff dff_A_ucYRhmgI0_1(.dout(w_dff_A_wDrIAQlP5_1),.din(w_dff_A_ucYRhmgI0_1),.clk(gclk));
	jdff dff_A_yco0T9be5_1(.dout(w_dff_A_ucYRhmgI0_1),.din(w_dff_A_yco0T9be5_1),.clk(gclk));
	jdff dff_A_LP808wx15_1(.dout(w_dff_A_yco0T9be5_1),.din(w_dff_A_LP808wx15_1),.clk(gclk));
	jdff dff_A_3kyqLb242_1(.dout(w_dff_A_LP808wx15_1),.din(w_dff_A_3kyqLb242_1),.clk(gclk));
	jdff dff_A_d9L3SHvs9_1(.dout(w_dff_A_3kyqLb242_1),.din(w_dff_A_d9L3SHvs9_1),.clk(gclk));
	jdff dff_A_KibjpU1d0_1(.dout(w_dff_A_d9L3SHvs9_1),.din(w_dff_A_KibjpU1d0_1),.clk(gclk));
	jdff dff_A_vSKhQeS71_1(.dout(w_dff_A_KibjpU1d0_1),.din(w_dff_A_vSKhQeS71_1),.clk(gclk));
	jdff dff_A_qSALVIPY3_0(.dout(w_n159_0[0]),.din(w_dff_A_qSALVIPY3_0),.clk(gclk));
	jdff dff_A_VlKvZzBP8_0(.dout(w_dff_A_qSALVIPY3_0),.din(w_dff_A_VlKvZzBP8_0),.clk(gclk));
	jdff dff_A_TN1YAt2a0_0(.dout(w_dff_A_VlKvZzBP8_0),.din(w_dff_A_TN1YAt2a0_0),.clk(gclk));
	jdff dff_A_l5XM0c368_0(.dout(w_dff_A_TN1YAt2a0_0),.din(w_dff_A_l5XM0c368_0),.clk(gclk));
	jdff dff_A_6KQD2n7m9_0(.dout(w_dff_A_l5XM0c368_0),.din(w_dff_A_6KQD2n7m9_0),.clk(gclk));
	jdff dff_A_xrX8NtgM4_0(.dout(w_dff_A_6KQD2n7m9_0),.din(w_dff_A_xrX8NtgM4_0),.clk(gclk));
	jdff dff_A_5JTPPUKV8_0(.dout(w_G34gat_0[0]),.din(w_dff_A_5JTPPUKV8_0),.clk(gclk));
	jdff dff_A_WNeU2Jem0_0(.dout(w_dff_A_5JTPPUKV8_0),.din(w_dff_A_WNeU2Jem0_0),.clk(gclk));
	jdff dff_A_6ig9zHsH1_0(.dout(w_dff_A_WNeU2Jem0_0),.din(w_dff_A_6ig9zHsH1_0),.clk(gclk));
	jdff dff_A_uCFpV3yA3_0(.dout(w_dff_A_6ig9zHsH1_0),.din(w_dff_A_uCFpV3yA3_0),.clk(gclk));
	jdff dff_A_C5IXaVC89_0(.dout(w_dff_A_uCFpV3yA3_0),.din(w_dff_A_C5IXaVC89_0),.clk(gclk));
	jdff dff_A_ogyN5u1A2_0(.dout(w_dff_A_C5IXaVC89_0),.din(w_dff_A_ogyN5u1A2_0),.clk(gclk));
	jdff dff_A_NJKvVWLC5_0(.dout(w_dff_A_ogyN5u1A2_0),.din(w_dff_A_NJKvVWLC5_0),.clk(gclk));
	jdff dff_A_qxnsOABw3_0(.dout(w_dff_A_NJKvVWLC5_0),.din(w_dff_A_qxnsOABw3_0),.clk(gclk));
	jdff dff_A_tWBVBbx02_0(.dout(w_dff_A_qxnsOABw3_0),.din(w_dff_A_tWBVBbx02_0),.clk(gclk));
	jdff dff_A_FKNzlUKt6_0(.dout(w_dff_A_tWBVBbx02_0),.din(w_dff_A_FKNzlUKt6_0),.clk(gclk));
	jdff dff_A_RgASNUCH6_0(.dout(w_dff_A_FKNzlUKt6_0),.din(w_dff_A_RgASNUCH6_0),.clk(gclk));
	jdff dff_A_neboB7sP3_0(.dout(w_dff_A_RgASNUCH6_0),.din(w_dff_A_neboB7sP3_0),.clk(gclk));
	jdff dff_A_TtTMic2f7_0(.dout(w_dff_A_neboB7sP3_0),.din(w_dff_A_TtTMic2f7_0),.clk(gclk));
	jdff dff_A_k1I87nsZ5_1(.dout(w_G34gat_0[1]),.din(w_dff_A_k1I87nsZ5_1),.clk(gclk));
	jdff dff_A_rrmacSUs2_1(.dout(w_dff_A_k1I87nsZ5_1),.din(w_dff_A_rrmacSUs2_1),.clk(gclk));
	jdff dff_A_fmBKZxip6_1(.dout(w_dff_A_rrmacSUs2_1),.din(w_dff_A_fmBKZxip6_1),.clk(gclk));
	jdff dff_A_zBfsPtvw5_1(.dout(w_dff_A_fmBKZxip6_1),.din(w_dff_A_zBfsPtvw5_1),.clk(gclk));
	jdff dff_A_gx0pTNFj7_1(.dout(w_dff_A_zBfsPtvw5_1),.din(w_dff_A_gx0pTNFj7_1),.clk(gclk));
	jdff dff_A_YNJ6AOjQ2_1(.dout(w_dff_A_gx0pTNFj7_1),.din(w_dff_A_YNJ6AOjQ2_1),.clk(gclk));
	jdff dff_A_FmmN99Q40_1(.dout(w_dff_A_YNJ6AOjQ2_1),.din(w_dff_A_FmmN99Q40_1),.clk(gclk));
	jdff dff_A_0qqjJV1q4_1(.dout(w_dff_A_FmmN99Q40_1),.din(w_dff_A_0qqjJV1q4_1),.clk(gclk));
	jdff dff_A_MAuFFSEN3_0(.dout(w_n156_0[0]),.din(w_dff_A_MAuFFSEN3_0),.clk(gclk));
	jdff dff_A_mjQk8Mm64_0(.dout(w_dff_A_MAuFFSEN3_0),.din(w_dff_A_mjQk8Mm64_0),.clk(gclk));
	jdff dff_A_978miXAZ9_0(.dout(w_dff_A_mjQk8Mm64_0),.din(w_dff_A_978miXAZ9_0),.clk(gclk));
	jdff dff_A_JEz8vuUG2_0(.dout(w_dff_A_978miXAZ9_0),.din(w_dff_A_JEz8vuUG2_0),.clk(gclk));
	jdff dff_A_3JMd7eMd4_0(.dout(w_dff_A_JEz8vuUG2_0),.din(w_dff_A_3JMd7eMd4_0),.clk(gclk));
	jdff dff_A_VGxBzT6Y2_0(.dout(w_dff_A_3JMd7eMd4_0),.din(w_dff_A_VGxBzT6Y2_0),.clk(gclk));
	jdff dff_A_iUhGKo2b6_1(.dout(w_n138_0[1]),.din(w_dff_A_iUhGKo2b6_1),.clk(gclk));
	jdff dff_A_S3391bGd9_1(.dout(w_dff_A_iUhGKo2b6_1),.din(w_dff_A_S3391bGd9_1),.clk(gclk));
	jdff dff_A_NK8WXUTU8_1(.dout(w_dff_A_S3391bGd9_1),.din(w_dff_A_NK8WXUTU8_1),.clk(gclk));
	jdff dff_A_CbNCsRrk0_1(.dout(w_dff_A_NK8WXUTU8_1),.din(w_dff_A_CbNCsRrk0_1),.clk(gclk));
	jdff dff_A_YnnGEYH09_1(.dout(w_dff_A_CbNCsRrk0_1),.din(w_dff_A_YnnGEYH09_1),.clk(gclk));
	jdff dff_A_D620hIjN3_1(.dout(w_dff_A_YnnGEYH09_1),.din(w_dff_A_D620hIjN3_1),.clk(gclk));
	jdff dff_A_EA4fEhLh9_0(.dout(w_G99gat_0[0]),.din(w_dff_A_EA4fEhLh9_0),.clk(gclk));
	jdff dff_A_mZeqW5Xc3_0(.dout(w_dff_A_EA4fEhLh9_0),.din(w_dff_A_mZeqW5Xc3_0),.clk(gclk));
	jdff dff_A_NioHEqBG4_0(.dout(w_dff_A_mZeqW5Xc3_0),.din(w_dff_A_NioHEqBG4_0),.clk(gclk));
	jdff dff_A_rHj2NQ2M1_0(.dout(w_dff_A_NioHEqBG4_0),.din(w_dff_A_rHj2NQ2M1_0),.clk(gclk));
	jdff dff_A_07mjf78m6_0(.dout(w_dff_A_rHj2NQ2M1_0),.din(w_dff_A_07mjf78m6_0),.clk(gclk));
	jdff dff_A_JWi0SZFn6_0(.dout(w_dff_A_07mjf78m6_0),.din(w_dff_A_JWi0SZFn6_0),.clk(gclk));
	jdff dff_A_09M2gSEs1_0(.dout(w_dff_A_JWi0SZFn6_0),.din(w_dff_A_09M2gSEs1_0),.clk(gclk));
	jdff dff_A_HWIp2MDX0_0(.dout(w_dff_A_09M2gSEs1_0),.din(w_dff_A_HWIp2MDX0_0),.clk(gclk));
	jdff dff_A_zGPZz4L48_1(.dout(w_G99gat_0[1]),.din(w_dff_A_zGPZz4L48_1),.clk(gclk));
	jdff dff_A_vMZ8YF8h8_1(.dout(w_dff_A_zGPZz4L48_1),.din(w_dff_A_vMZ8YF8h8_1),.clk(gclk));
	jdff dff_A_g38jHedp6_1(.dout(w_dff_A_vMZ8YF8h8_1),.din(w_dff_A_g38jHedp6_1),.clk(gclk));
	jdff dff_A_ePubq2rA8_1(.dout(w_dff_A_g38jHedp6_1),.din(w_dff_A_ePubq2rA8_1),.clk(gclk));
	jdff dff_A_J7YzgHXy3_1(.dout(w_dff_A_ePubq2rA8_1),.din(w_dff_A_J7YzgHXy3_1),.clk(gclk));
	jdff dff_A_K3HiBZhZ0_1(.dout(w_dff_A_J7YzgHXy3_1),.din(w_dff_A_K3HiBZhZ0_1),.clk(gclk));
	jdff dff_A_9R5cDTOQ5_1(.dout(w_dff_A_K3HiBZhZ0_1),.din(w_dff_A_9R5cDTOQ5_1),.clk(gclk));
	jdff dff_A_rJxT69mx2_1(.dout(w_dff_A_9R5cDTOQ5_1),.din(w_dff_A_rJxT69mx2_1),.clk(gclk));
	jdff dff_A_pNZ02Kme4_1(.dout(w_dff_A_rJxT69mx2_1),.din(w_dff_A_pNZ02Kme4_1),.clk(gclk));
	jdff dff_A_XPq9qGD88_1(.dout(w_dff_A_pNZ02Kme4_1),.din(w_dff_A_XPq9qGD88_1),.clk(gclk));
	jdff dff_A_GiLn6BOZ3_1(.dout(w_dff_A_XPq9qGD88_1),.din(w_dff_A_GiLn6BOZ3_1),.clk(gclk));
	jdff dff_A_am0tLmpk8_1(.dout(w_dff_A_GiLn6BOZ3_1),.din(w_dff_A_am0tLmpk8_1),.clk(gclk));
	jdff dff_A_9Sv5mRmP8_1(.dout(w_dff_A_am0tLmpk8_1),.din(w_dff_A_9Sv5mRmP8_1),.clk(gclk));
	jdff dff_A_WCZ0mFjC7_0(.dout(w_n151_0[0]),.din(w_dff_A_WCZ0mFjC7_0),.clk(gclk));
	jdff dff_A_g9gBizeZ1_0(.dout(w_dff_A_WCZ0mFjC7_0),.din(w_dff_A_g9gBizeZ1_0),.clk(gclk));
	jdff dff_A_loWXzfhA9_0(.dout(w_dff_A_g9gBizeZ1_0),.din(w_dff_A_loWXzfhA9_0),.clk(gclk));
	jdff dff_A_0rNdRn0C5_0(.dout(w_dff_A_loWXzfhA9_0),.din(w_dff_A_0rNdRn0C5_0),.clk(gclk));
	jdff dff_A_nUKewTiJ9_0(.dout(w_dff_A_0rNdRn0C5_0),.din(w_dff_A_nUKewTiJ9_0),.clk(gclk));
	jdff dff_A_DnJVo4kj9_0(.dout(w_dff_A_nUKewTiJ9_0),.din(w_dff_A_DnJVo4kj9_0),.clk(gclk));
	jdff dff_B_s0c1Tnw43_1(.din(n48),.dout(w_dff_B_s0c1Tnw43_1),.clk(gclk));
	jdff dff_B_rrynMJak1_1(.din(n61),.dout(w_dff_B_rrynMJak1_1),.clk(gclk));
	jdff dff_A_Fw0m2RSD9_0(.dout(w_n64_0[0]),.din(w_dff_A_Fw0m2RSD9_0),.clk(gclk));
	jdff dff_A_0iCzWIbG2_0(.dout(w_dff_A_Fw0m2RSD9_0),.din(w_dff_A_0iCzWIbG2_0),.clk(gclk));
	jdff dff_A_yE7HAdrQ7_0(.dout(w_dff_A_0iCzWIbG2_0),.din(w_dff_A_yE7HAdrQ7_0),.clk(gclk));
	jdff dff_A_xm6UIbV59_0(.dout(w_dff_A_yE7HAdrQ7_0),.din(w_dff_A_xm6UIbV59_0),.clk(gclk));
	jdff dff_A_7n9LOtu14_0(.dout(w_dff_A_xm6UIbV59_0),.din(w_dff_A_7n9LOtu14_0),.clk(gclk));
	jdff dff_A_hJNfhKKn3_0(.dout(w_n62_0[0]),.din(w_dff_A_hJNfhKKn3_0),.clk(gclk));
	jdff dff_A_t59ejE1I7_0(.dout(w_dff_A_hJNfhKKn3_0),.din(w_dff_A_t59ejE1I7_0),.clk(gclk));
	jdff dff_A_30qGjJbl3_0(.dout(w_dff_A_t59ejE1I7_0),.din(w_dff_A_30qGjJbl3_0),.clk(gclk));
	jdff dff_A_w5k1SJh39_0(.dout(w_dff_A_30qGjJbl3_0),.din(w_dff_A_w5k1SJh39_0),.clk(gclk));
	jdff dff_A_w2p70dmt4_0(.dout(w_dff_A_w5k1SJh39_0),.din(w_dff_A_w2p70dmt4_0),.clk(gclk));
	jdff dff_A_CpT96k2v0_0(.dout(w_n60_0[0]),.din(w_dff_A_CpT96k2v0_0),.clk(gclk));
	jdff dff_A_MTV7oEoe4_0(.dout(w_dff_A_CpT96k2v0_0),.din(w_dff_A_MTV7oEoe4_0),.clk(gclk));
	jdff dff_A_gUjf7bgp9_0(.dout(w_dff_A_MTV7oEoe4_0),.din(w_dff_A_gUjf7bgp9_0),.clk(gclk));
	jdff dff_A_U3ECG0Ey4_0(.dout(w_dff_A_gUjf7bgp9_0),.din(w_dff_A_U3ECG0Ey4_0),.clk(gclk));
	jdff dff_A_BXhbeJ6u9_0(.dout(w_dff_A_U3ECG0Ey4_0),.din(w_dff_A_BXhbeJ6u9_0),.clk(gclk));
	jdff dff_A_BRg9RaPD8_0(.dout(w_n57_0[0]),.din(w_dff_A_BRg9RaPD8_0),.clk(gclk));
	jdff dff_A_sjZR4kzv5_0(.dout(w_dff_A_BRg9RaPD8_0),.din(w_dff_A_sjZR4kzv5_0),.clk(gclk));
	jdff dff_A_5LMN1alR9_0(.dout(w_dff_A_sjZR4kzv5_0),.din(w_dff_A_5LMN1alR9_0),.clk(gclk));
	jdff dff_A_EghAq9VE0_0(.dout(w_dff_A_5LMN1alR9_0),.din(w_dff_A_EghAq9VE0_0),.clk(gclk));
	jdff dff_A_pnBdnbqj7_0(.dout(w_n54_0[0]),.din(w_dff_A_pnBdnbqj7_0),.clk(gclk));
	jdff dff_A_5iR8ySs13_0(.dout(w_dff_A_pnBdnbqj7_0),.din(w_dff_A_5iR8ySs13_0),.clk(gclk));
	jdff dff_A_TBOhhYWR0_0(.dout(w_dff_A_5iR8ySs13_0),.din(w_dff_A_TBOhhYWR0_0),.clk(gclk));
	jdff dff_A_emfxJcVz0_0(.dout(w_dff_A_TBOhhYWR0_0),.din(w_dff_A_emfxJcVz0_0),.clk(gclk));
	jdff dff_A_oqnyvqRT4_0(.dout(w_dff_A_emfxJcVz0_0),.din(w_dff_A_oqnyvqRT4_0),.clk(gclk));
	jdff dff_A_m5XAkFSM9_0(.dout(w_n51_0[0]),.din(w_dff_A_m5XAkFSM9_0),.clk(gclk));
	jdff dff_A_IpSgGjO59_0(.dout(w_dff_A_m5XAkFSM9_0),.din(w_dff_A_IpSgGjO59_0),.clk(gclk));
	jdff dff_A_l45PGS1R4_0(.dout(w_dff_A_IpSgGjO59_0),.din(w_dff_A_l45PGS1R4_0),.clk(gclk));
	jdff dff_A_7RfAld141_0(.dout(w_dff_A_l45PGS1R4_0),.din(w_dff_A_7RfAld141_0),.clk(gclk));
	jdff dff_A_L2s6nSm88_0(.dout(w_dff_A_7RfAld141_0),.din(w_dff_A_L2s6nSm88_0),.clk(gclk));
	jdff dff_A_GW1TgdPw6_0(.dout(w_n47_0[0]),.din(w_dff_A_GW1TgdPw6_0),.clk(gclk));
	jdff dff_A_UUIjfV6H9_0(.dout(w_dff_A_GW1TgdPw6_0),.din(w_dff_A_UUIjfV6H9_0),.clk(gclk));
	jdff dff_A_Fe8ugEQt2_0(.dout(w_dff_A_UUIjfV6H9_0),.din(w_dff_A_Fe8ugEQt2_0),.clk(gclk));
	jdff dff_A_cYeha5vQ3_0(.dout(w_G21gat_0[0]),.din(w_dff_A_cYeha5vQ3_0),.clk(gclk));
	jdff dff_A_zmuJEHr61_0(.dout(w_dff_A_cYeha5vQ3_0),.din(w_dff_A_zmuJEHr61_0),.clk(gclk));
	jdff dff_A_jyBUWZxt2_0(.dout(w_dff_A_zmuJEHr61_0),.din(w_dff_A_jyBUWZxt2_0),.clk(gclk));
	jdff dff_A_qxNhJFFj9_0(.dout(w_dff_A_jyBUWZxt2_0),.din(w_dff_A_qxNhJFFj9_0),.clk(gclk));
	jdff dff_A_eMw26Pmx1_0(.dout(w_dff_A_qxNhJFFj9_0),.din(w_dff_A_eMw26Pmx1_0),.clk(gclk));
	jdff dff_A_GFmMQHXB9_0(.dout(w_dff_A_eMw26Pmx1_0),.din(w_dff_A_GFmMQHXB9_0),.clk(gclk));
	jdff dff_A_oAujPlQh2_0(.dout(w_dff_A_GFmMQHXB9_0),.din(w_dff_A_oAujPlQh2_0),.clk(gclk));
	jdff dff_A_hbs3gKxv1_0(.dout(w_dff_A_oAujPlQh2_0),.din(w_dff_A_hbs3gKxv1_0),.clk(gclk));
	jdff dff_A_izcbH5rk2_0(.dout(w_dff_A_hbs3gKxv1_0),.din(w_dff_A_izcbH5rk2_0),.clk(gclk));
	jdff dff_A_ZJZQzvDr9_0(.dout(w_dff_A_izcbH5rk2_0),.din(w_dff_A_ZJZQzvDr9_0),.clk(gclk));
	jdff dff_A_UE9Jyjob2_0(.dout(w_dff_A_ZJZQzvDr9_0),.din(w_dff_A_UE9Jyjob2_0),.clk(gclk));
	jdff dff_A_sGjbF2kD1_0(.dout(w_dff_A_UE9Jyjob2_0),.din(w_dff_A_sGjbF2kD1_0),.clk(gclk));
	jdff dff_A_dHsrHFZ11_0(.dout(w_dff_A_sGjbF2kD1_0),.din(w_dff_A_dHsrHFZ11_0),.clk(gclk));
	jdff dff_A_axtwTHXH0_1(.dout(w_G21gat_0[1]),.din(w_dff_A_axtwTHXH0_1),.clk(gclk));
	jdff dff_A_REgmSQsm0_1(.dout(w_dff_A_axtwTHXH0_1),.din(w_dff_A_REgmSQsm0_1),.clk(gclk));
	jdff dff_A_LvvHirrd2_1(.dout(w_dff_A_REgmSQsm0_1),.din(w_dff_A_LvvHirrd2_1),.clk(gclk));
	jdff dff_A_kx8knwZf4_1(.dout(w_dff_A_LvvHirrd2_1),.din(w_dff_A_kx8knwZf4_1),.clk(gclk));
	jdff dff_A_eJFGdXfV6_1(.dout(w_dff_A_kx8knwZf4_1),.din(w_dff_A_eJFGdXfV6_1),.clk(gclk));
	jdff dff_A_ajfTYSEm0_1(.dout(w_dff_A_eJFGdXfV6_1),.din(w_dff_A_ajfTYSEm0_1),.clk(gclk));
	jdff dff_A_A94sENI80_1(.dout(w_dff_A_ajfTYSEm0_1),.din(w_dff_A_A94sENI80_1),.clk(gclk));
	jdff dff_A_gpuN8SLz2_1(.dout(w_dff_A_A94sENI80_1),.din(w_dff_A_gpuN8SLz2_1),.clk(gclk));
	jdff dff_A_5bE7cs9u1_0(.dout(w_n102_0[0]),.din(w_dff_A_5bE7cs9u1_0),.clk(gclk));
	jdff dff_A_7x6ncHxp5_0(.dout(w_dff_A_5bE7cs9u1_0),.din(w_dff_A_7x6ncHxp5_0),.clk(gclk));
	jdff dff_A_9JiKSFa46_0(.dout(w_dff_A_7x6ncHxp5_0),.din(w_dff_A_9JiKSFa46_0),.clk(gclk));
	jdff dff_A_La0Lioxn3_0(.dout(w_dff_A_9JiKSFa46_0),.din(w_dff_A_La0Lioxn3_0),.clk(gclk));
	jdff dff_A_Up8MHMLe2_0(.dout(w_dff_A_La0Lioxn3_0),.din(w_dff_A_Up8MHMLe2_0),.clk(gclk));
	jdff dff_B_egBKhqmp2_2(.din(n102),.dout(w_dff_B_egBKhqmp2_2),.clk(gclk));
	jdff dff_B_kGUCirf42_2(.din(w_dff_B_egBKhqmp2_2),.dout(w_dff_B_kGUCirf42_2),.clk(gclk));
	jdff dff_B_YcbZLqPw5_2(.din(w_dff_B_kGUCirf42_2),.dout(w_dff_B_YcbZLqPw5_2),.clk(gclk));
	jdff dff_B_iR8KAdii6_2(.din(w_dff_B_YcbZLqPw5_2),.dout(w_dff_B_iR8KAdii6_2),.clk(gclk));
	jdff dff_B_yLq0bkSN3_2(.din(w_dff_B_iR8KAdii6_2),.dout(w_dff_B_yLq0bkSN3_2),.clk(gclk));
	jdff dff_B_5YKmKlW35_2(.din(w_dff_B_yLq0bkSN3_2),.dout(w_dff_B_5YKmKlW35_2),.clk(gclk));
	jdff dff_B_4eM6QmVo7_2(.din(w_dff_B_5YKmKlW35_2),.dout(w_dff_B_4eM6QmVo7_2),.clk(gclk));
	jdff dff_A_ezEMIm566_0(.dout(w_G73gat_0[0]),.din(w_dff_A_ezEMIm566_0),.clk(gclk));
	jdff dff_A_hTMZdTzv6_0(.dout(w_dff_A_ezEMIm566_0),.din(w_dff_A_hTMZdTzv6_0),.clk(gclk));
	jdff dff_A_e7yhCOKA5_0(.dout(w_dff_A_hTMZdTzv6_0),.din(w_dff_A_e7yhCOKA5_0),.clk(gclk));
	jdff dff_A_UIfke8RR2_0(.dout(w_dff_A_e7yhCOKA5_0),.din(w_dff_A_UIfke8RR2_0),.clk(gclk));
	jdff dff_A_EY9DA8MV3_0(.dout(w_dff_A_UIfke8RR2_0),.din(w_dff_A_EY9DA8MV3_0),.clk(gclk));
	jdff dff_A_BgwTVaKS1_0(.dout(w_dff_A_EY9DA8MV3_0),.din(w_dff_A_BgwTVaKS1_0),.clk(gclk));
	jdff dff_A_QZNzZTnj5_0(.dout(w_dff_A_BgwTVaKS1_0),.din(w_dff_A_QZNzZTnj5_0),.clk(gclk));
	jdff dff_A_1fdHG0aV6_0(.dout(w_dff_A_QZNzZTnj5_0),.din(w_dff_A_1fdHG0aV6_0),.clk(gclk));
	jdff dff_A_w6VFdMW76_0(.dout(w_dff_A_1fdHG0aV6_0),.din(w_dff_A_w6VFdMW76_0),.clk(gclk));
	jdff dff_A_lk2s9mPd5_0(.dout(w_dff_A_w6VFdMW76_0),.din(w_dff_A_lk2s9mPd5_0),.clk(gclk));
	jdff dff_A_XpQRtSzi7_0(.dout(w_dff_A_lk2s9mPd5_0),.din(w_dff_A_XpQRtSzi7_0),.clk(gclk));
	jdff dff_A_3CTgq0pL6_0(.dout(w_dff_A_XpQRtSzi7_0),.din(w_dff_A_3CTgq0pL6_0),.clk(gclk));
	jdff dff_A_oOw3wfMq8_0(.dout(w_dff_A_3CTgq0pL6_0),.din(w_dff_A_oOw3wfMq8_0),.clk(gclk));
	jdff dff_A_v4cc3wmn1_1(.dout(w_G73gat_0[1]),.din(w_dff_A_v4cc3wmn1_1),.clk(gclk));
	jdff dff_A_U9Iwbpkv7_1(.dout(w_dff_A_v4cc3wmn1_1),.din(w_dff_A_U9Iwbpkv7_1),.clk(gclk));
	jdff dff_A_1fzvDvob2_1(.dout(w_dff_A_U9Iwbpkv7_1),.din(w_dff_A_1fzvDvob2_1),.clk(gclk));
	jdff dff_A_4WvKJtRH4_1(.dout(w_dff_A_1fzvDvob2_1),.din(w_dff_A_4WvKJtRH4_1),.clk(gclk));
	jdff dff_A_yHVOro008_1(.dout(w_dff_A_4WvKJtRH4_1),.din(w_dff_A_yHVOro008_1),.clk(gclk));
	jdff dff_A_msO9EwR00_1(.dout(w_dff_A_yHVOro008_1),.din(w_dff_A_msO9EwR00_1),.clk(gclk));
	jdff dff_A_kIzOScC21_1(.dout(w_dff_A_msO9EwR00_1),.din(w_dff_A_kIzOScC21_1),.clk(gclk));
	jdff dff_A_mkmU92eL9_1(.dout(w_dff_A_kIzOScC21_1),.din(w_dff_A_mkmU92eL9_1),.clk(gclk));
	jdff dff_A_pUAz7cfj8_0(.dout(w_n104_0[0]),.din(w_dff_A_pUAz7cfj8_0),.clk(gclk));
	jdff dff_A_d4L7to5l9_0(.dout(w_dff_A_pUAz7cfj8_0),.din(w_dff_A_d4L7to5l9_0),.clk(gclk));
	jdff dff_A_lZeKiMiY3_0(.dout(w_dff_A_d4L7to5l9_0),.din(w_dff_A_lZeKiMiY3_0),.clk(gclk));
	jdff dff_A_v6HKAFTI1_0(.dout(w_dff_A_lZeKiMiY3_0),.din(w_dff_A_v6HKAFTI1_0),.clk(gclk));
	jdff dff_A_CZqs8dwm3_0(.dout(w_dff_A_v6HKAFTI1_0),.din(w_dff_A_CZqs8dwm3_0),.clk(gclk));
	jdff dff_A_zxeppp4M2_0(.dout(w_dff_A_CZqs8dwm3_0),.din(w_dff_A_zxeppp4M2_0),.clk(gclk));
	jdff dff_B_FXFeITBu7_1(.din(n72),.dout(w_dff_B_FXFeITBu7_1),.clk(gclk));
	jdff dff_B_vtrJgknM1_1(.din(n85),.dout(w_dff_B_vtrJgknM1_1),.clk(gclk));
	jdff dff_A_nTTTe9KR8_0(.dout(w_n88_0[0]),.din(w_dff_A_nTTTe9KR8_0),.clk(gclk));
	jdff dff_A_zYlq5Etq3_0(.dout(w_dff_A_nTTTe9KR8_0),.din(w_dff_A_zYlq5Etq3_0),.clk(gclk));
	jdff dff_A_wGNpy5QZ2_0(.dout(w_dff_A_zYlq5Etq3_0),.din(w_dff_A_wGNpy5QZ2_0),.clk(gclk));
	jdff dff_A_pctuj1dG3_0(.dout(w_dff_A_wGNpy5QZ2_0),.din(w_dff_A_pctuj1dG3_0),.clk(gclk));
	jdff dff_A_zSINf0dP3_0(.dout(w_dff_A_pctuj1dG3_0),.din(w_dff_A_zSINf0dP3_0),.clk(gclk));
	jdff dff_A_EhqGlHxz9_0(.dout(w_dff_A_zSINf0dP3_0),.din(w_dff_A_EhqGlHxz9_0),.clk(gclk));
	jdff dff_A_Swk2Fr2z6_0(.dout(w_G82gat_0[0]),.din(w_dff_A_Swk2Fr2z6_0),.clk(gclk));
	jdff dff_A_sL3UCyQ09_0(.dout(w_dff_A_Swk2Fr2z6_0),.din(w_dff_A_sL3UCyQ09_0),.clk(gclk));
	jdff dff_A_FOWyX1XP9_0(.dout(w_dff_A_sL3UCyQ09_0),.din(w_dff_A_FOWyX1XP9_0),.clk(gclk));
	jdff dff_A_FWkn7Djz2_0(.dout(w_dff_A_FOWyX1XP9_0),.din(w_dff_A_FWkn7Djz2_0),.clk(gclk));
	jdff dff_A_H92DG0GL3_0(.dout(w_dff_A_FWkn7Djz2_0),.din(w_dff_A_H92DG0GL3_0),.clk(gclk));
	jdff dff_A_C9MKShi57_0(.dout(w_dff_A_H92DG0GL3_0),.din(w_dff_A_C9MKShi57_0),.clk(gclk));
	jdff dff_A_8NwcASrU2_0(.dout(w_dff_A_C9MKShi57_0),.din(w_dff_A_8NwcASrU2_0),.clk(gclk));
	jdff dff_A_QxQf8HVV3_2(.dout(w_G82gat_0[2]),.din(w_dff_A_QxQf8HVV3_2),.clk(gclk));
	jdff dff_A_Lw6AVonP7_0(.dout(w_G76gat_0[0]),.din(w_dff_A_Lw6AVonP7_0),.clk(gclk));
	jdff dff_A_sgLv7Sqh6_0(.dout(w_dff_A_Lw6AVonP7_0),.din(w_dff_A_sgLv7Sqh6_0),.clk(gclk));
	jdff dff_A_qCEbS0iY1_0(.dout(w_dff_A_sgLv7Sqh6_0),.din(w_dff_A_qCEbS0iY1_0),.clk(gclk));
	jdff dff_A_Xm31pBam3_0(.dout(w_dff_A_qCEbS0iY1_0),.din(w_dff_A_Xm31pBam3_0),.clk(gclk));
	jdff dff_A_kzPWKD4u9_0(.dout(w_dff_A_Xm31pBam3_0),.din(w_dff_A_kzPWKD4u9_0),.clk(gclk));
	jdff dff_A_m0axmQEX1_0(.dout(w_dff_A_kzPWKD4u9_0),.din(w_dff_A_m0axmQEX1_0),.clk(gclk));
	jdff dff_A_SDsstCuO9_1(.dout(w_G76gat_0[1]),.din(w_dff_A_SDsstCuO9_1),.clk(gclk));
	jdff dff_A_8wKgaRna2_0(.dout(w_n86_0[0]),.din(w_dff_A_8wKgaRna2_0),.clk(gclk));
	jdff dff_A_uryQFvw91_0(.dout(w_dff_A_8wKgaRna2_0),.din(w_dff_A_uryQFvw91_0),.clk(gclk));
	jdff dff_A_w8aiLEMO9_0(.dout(w_dff_A_uryQFvw91_0),.din(w_dff_A_w8aiLEMO9_0),.clk(gclk));
	jdff dff_A_mDfcpBla1_0(.dout(w_dff_A_w8aiLEMO9_0),.din(w_dff_A_mDfcpBla1_0),.clk(gclk));
	jdff dff_A_ErQX5kCv7_0(.dout(w_dff_A_mDfcpBla1_0),.din(w_dff_A_ErQX5kCv7_0),.clk(gclk));
	jdff dff_A_69aeXXNp3_0(.dout(w_dff_A_ErQX5kCv7_0),.din(w_dff_A_69aeXXNp3_0),.clk(gclk));
	jdff dff_A_YfnHZVw77_0(.dout(w_G95gat_0[0]),.din(w_dff_A_YfnHZVw77_0),.clk(gclk));
	jdff dff_A_8zuRIUjp8_0(.dout(w_dff_A_YfnHZVw77_0),.din(w_dff_A_8zuRIUjp8_0),.clk(gclk));
	jdff dff_A_SHlor39q6_0(.dout(w_dff_A_8zuRIUjp8_0),.din(w_dff_A_SHlor39q6_0),.clk(gclk));
	jdff dff_A_5XHH9LnT2_0(.dout(w_dff_A_SHlor39q6_0),.din(w_dff_A_5XHH9LnT2_0),.clk(gclk));
	jdff dff_A_DCEaacXu6_0(.dout(w_dff_A_5XHH9LnT2_0),.din(w_dff_A_DCEaacXu6_0),.clk(gclk));
	jdff dff_A_zO9u0GcB2_0(.dout(w_dff_A_DCEaacXu6_0),.din(w_dff_A_zO9u0GcB2_0),.clk(gclk));
	jdff dff_A_s6eqjM6c5_0(.dout(w_dff_A_zO9u0GcB2_0),.din(w_dff_A_s6eqjM6c5_0),.clk(gclk));
	jdff dff_A_EYXFSrfy1_2(.dout(w_G95gat_0[2]),.din(w_dff_A_EYXFSrfy1_2),.clk(gclk));
	jdff dff_A_HMjUPUtq6_0(.dout(w_G89gat_0[0]),.din(w_dff_A_HMjUPUtq6_0),.clk(gclk));
	jdff dff_A_Yp7kiGvO6_0(.dout(w_dff_A_HMjUPUtq6_0),.din(w_dff_A_Yp7kiGvO6_0),.clk(gclk));
	jdff dff_A_F5QxENqL9_0(.dout(w_dff_A_Yp7kiGvO6_0),.din(w_dff_A_F5QxENqL9_0),.clk(gclk));
	jdff dff_A_SwLhpr7g5_0(.dout(w_dff_A_F5QxENqL9_0),.din(w_dff_A_SwLhpr7g5_0),.clk(gclk));
	jdff dff_A_uyak5vtX8_0(.dout(w_dff_A_SwLhpr7g5_0),.din(w_dff_A_uyak5vtX8_0),.clk(gclk));
	jdff dff_A_5c5qQ5998_0(.dout(w_dff_A_uyak5vtX8_0),.din(w_dff_A_5c5qQ5998_0),.clk(gclk));
	jdff dff_A_jsSRzS613_1(.dout(w_G89gat_0[1]),.din(w_dff_A_jsSRzS613_1),.clk(gclk));
	jdff dff_A_Yle2qnlC2_0(.dout(w_n84_0[0]),.din(w_dff_A_Yle2qnlC2_0),.clk(gclk));
	jdff dff_A_pM0DdqxR2_0(.dout(w_dff_A_Yle2qnlC2_0),.din(w_dff_A_pM0DdqxR2_0),.clk(gclk));
	jdff dff_A_uWU4UWII3_0(.dout(w_dff_A_pM0DdqxR2_0),.din(w_dff_A_uWU4UWII3_0),.clk(gclk));
	jdff dff_A_SbPzlKR21_0(.dout(w_dff_A_uWU4UWII3_0),.din(w_dff_A_SbPzlKR21_0),.clk(gclk));
	jdff dff_A_hsy488Jo2_0(.dout(w_dff_A_SbPzlKR21_0),.din(w_dff_A_hsy488Jo2_0),.clk(gclk));
	jdff dff_A_jJ4botKv4_0(.dout(w_dff_A_hsy488Jo2_0),.din(w_dff_A_jJ4botKv4_0),.clk(gclk));
	jdff dff_A_MLFC6cQL6_0(.dout(w_G4gat_0[0]),.din(w_dff_A_MLFC6cQL6_0),.clk(gclk));
	jdff dff_A_KdzitkGW9_0(.dout(w_dff_A_MLFC6cQL6_0),.din(w_dff_A_KdzitkGW9_0),.clk(gclk));
	jdff dff_A_lGMJ01SH2_0(.dout(w_dff_A_KdzitkGW9_0),.din(w_dff_A_lGMJ01SH2_0),.clk(gclk));
	jdff dff_A_f7UkhaFr8_0(.dout(w_dff_A_lGMJ01SH2_0),.din(w_dff_A_f7UkhaFr8_0),.clk(gclk));
	jdff dff_A_lZrKjVFF9_0(.dout(w_dff_A_f7UkhaFr8_0),.din(w_dff_A_lZrKjVFF9_0),.clk(gclk));
	jdff dff_A_Tlk1XYYi2_0(.dout(w_dff_A_lZrKjVFF9_0),.din(w_dff_A_Tlk1XYYi2_0),.clk(gclk));
	jdff dff_A_dAcs90u54_0(.dout(w_dff_A_Tlk1XYYi2_0),.din(w_dff_A_dAcs90u54_0),.clk(gclk));
	jdff dff_A_9TzEKDLb0_2(.dout(w_G4gat_0[2]),.din(w_dff_A_9TzEKDLb0_2),.clk(gclk));
	jdff dff_A_nLswiUEQ4_0(.dout(w_G1gat_0[0]),.din(w_dff_A_nLswiUEQ4_0),.clk(gclk));
	jdff dff_A_SgXvakfC7_0(.dout(w_dff_A_nLswiUEQ4_0),.din(w_dff_A_SgXvakfC7_0),.clk(gclk));
	jdff dff_A_I04w0Ed15_0(.dout(w_dff_A_SgXvakfC7_0),.din(w_dff_A_I04w0Ed15_0),.clk(gclk));
	jdff dff_A_iyBw2BMF3_0(.dout(w_dff_A_I04w0Ed15_0),.din(w_dff_A_iyBw2BMF3_0),.clk(gclk));
	jdff dff_A_6ErcL3651_0(.dout(w_dff_A_iyBw2BMF3_0),.din(w_dff_A_6ErcL3651_0),.clk(gclk));
	jdff dff_A_nuQVfrCK8_0(.dout(w_dff_A_6ErcL3651_0),.din(w_dff_A_nuQVfrCK8_0),.clk(gclk));
	jdff dff_A_bat33BQT1_1(.dout(w_G1gat_0[1]),.din(w_dff_A_bat33BQT1_1),.clk(gclk));
	jdff dff_A_xBVxXj4H3_0(.dout(w_n81_0[0]),.din(w_dff_A_xBVxXj4H3_0),.clk(gclk));
	jdff dff_A_Ibvd90Nt5_0(.dout(w_dff_A_xBVxXj4H3_0),.din(w_dff_A_Ibvd90Nt5_0),.clk(gclk));
	jdff dff_A_BVNvk7AR9_0(.dout(w_dff_A_Ibvd90Nt5_0),.din(w_dff_A_BVNvk7AR9_0),.clk(gclk));
	jdff dff_A_a03MK4F13_0(.dout(w_dff_A_BVNvk7AR9_0),.din(w_dff_A_a03MK4F13_0),.clk(gclk));
	jdff dff_A_2mHympoU3_0(.dout(w_n80_0[0]),.din(w_dff_A_2mHympoU3_0),.clk(gclk));
	jdff dff_A_TFZNP5og8_0(.dout(w_dff_A_2mHympoU3_0),.din(w_dff_A_TFZNP5og8_0),.clk(gclk));
	jdff dff_A_hzuSuDqq4_0(.dout(w_dff_A_TFZNP5og8_0),.din(w_dff_A_hzuSuDqq4_0),.clk(gclk));
	jdff dff_A_k9oBrKtw7_0(.dout(w_dff_A_hzuSuDqq4_0),.din(w_dff_A_k9oBrKtw7_0),.clk(gclk));
	jdff dff_A_qb8llft07_0(.dout(w_dff_A_k9oBrKtw7_0),.din(w_dff_A_qb8llft07_0),.clk(gclk));
	jdff dff_A_KVPLnuKV2_0(.dout(w_dff_A_qb8llft07_0),.din(w_dff_A_KVPLnuKV2_0),.clk(gclk));
	jdff dff_A_wz1dhINR5_0(.dout(w_dff_A_KVPLnuKV2_0),.din(w_dff_A_wz1dhINR5_0),.clk(gclk));
	jdff dff_A_ztoZ4Ik43_0(.dout(w_dff_A_wz1dhINR5_0),.din(w_dff_A_ztoZ4Ik43_0),.clk(gclk));
	jdff dff_A_AIYD32ue7_0(.dout(w_dff_A_ztoZ4Ik43_0),.din(w_dff_A_AIYD32ue7_0),.clk(gclk));
	jdff dff_A_3U8FYw7z2_0(.dout(w_dff_A_AIYD32ue7_0),.din(w_dff_A_3U8FYw7z2_0),.clk(gclk));
	jdff dff_A_xchP7zrc5_0(.dout(w_dff_A_3U8FYw7z2_0),.din(w_dff_A_xchP7zrc5_0),.clk(gclk));
	jdff dff_A_yQncFvPD4_0(.dout(w_dff_A_xchP7zrc5_0),.din(w_dff_A_yQncFvPD4_0),.clk(gclk));
	jdff dff_A_xa2axSfF4_0(.dout(w_dff_A_yQncFvPD4_0),.din(w_dff_A_xa2axSfF4_0),.clk(gclk));
	jdff dff_A_v8chX6U61_0(.dout(w_dff_A_xa2axSfF4_0),.din(w_dff_A_v8chX6U61_0),.clk(gclk));
	jdff dff_A_840EB0C47_0(.dout(w_dff_A_v8chX6U61_0),.din(w_dff_A_840EB0C47_0),.clk(gclk));
	jdff dff_A_wd53ojks9_0(.dout(w_dff_A_840EB0C47_0),.din(w_dff_A_wd53ojks9_0),.clk(gclk));
	jdff dff_A_LO2AdWXo9_0(.dout(w_dff_A_wd53ojks9_0),.din(w_dff_A_LO2AdWXo9_0),.clk(gclk));
	jdff dff_A_6lDPQMiM6_0(.dout(w_dff_A_LO2AdWXo9_0),.din(w_dff_A_6lDPQMiM6_0),.clk(gclk));
	jdff dff_A_58rfLbq44_0(.dout(w_dff_A_6lDPQMiM6_0),.din(w_dff_A_58rfLbq44_0),.clk(gclk));
	jdff dff_A_GLScgb9d0_0(.dout(w_dff_A_58rfLbq44_0),.din(w_dff_A_GLScgb9d0_0),.clk(gclk));
	jdff dff_A_PnGpoDEQ5_0(.dout(w_dff_A_GLScgb9d0_0),.din(w_dff_A_PnGpoDEQ5_0),.clk(gclk));
	jdff dff_A_putrv7vJ4_1(.dout(w_G56gat_1[1]),.din(w_dff_A_putrv7vJ4_1),.clk(gclk));
	jdff dff_A_17DCkZix0_1(.dout(w_G56gat_0[1]),.din(w_dff_A_17DCkZix0_1),.clk(gclk));
	jdff dff_A_GGOXVVd55_1(.dout(w_dff_A_17DCkZix0_1),.din(w_dff_A_GGOXVVd55_1),.clk(gclk));
	jdff dff_A_2G7GTXXA1_1(.dout(w_dff_A_GGOXVVd55_1),.din(w_dff_A_2G7GTXXA1_1),.clk(gclk));
	jdff dff_A_WmTVgcOY8_1(.dout(w_dff_A_2G7GTXXA1_1),.din(w_dff_A_WmTVgcOY8_1),.clk(gclk));
	jdff dff_A_sf7ceMWh8_1(.dout(w_dff_A_WmTVgcOY8_1),.din(w_dff_A_sf7ceMWh8_1),.clk(gclk));
	jdff dff_A_uuRuBxWL8_1(.dout(w_dff_A_sf7ceMWh8_1),.din(w_dff_A_uuRuBxWL8_1),.clk(gclk));
	jdff dff_A_b7vCj8VR6_1(.dout(w_dff_A_uuRuBxWL8_1),.din(w_dff_A_b7vCj8VR6_1),.clk(gclk));
	jdff dff_A_YGd7f3wq6_1(.dout(w_dff_A_b7vCj8VR6_1),.din(w_dff_A_YGd7f3wq6_1),.clk(gclk));
	jdff dff_A_woP5CPUj6_1(.dout(w_dff_A_YGd7f3wq6_1),.din(w_dff_A_woP5CPUj6_1),.clk(gclk));
	jdff dff_A_oAwbT1it9_1(.dout(w_dff_A_woP5CPUj6_1),.din(w_dff_A_oAwbT1it9_1),.clk(gclk));
	jdff dff_A_hFXxqUvB9_1(.dout(w_dff_A_oAwbT1it9_1),.din(w_dff_A_hFXxqUvB9_1),.clk(gclk));
	jdff dff_A_ACcCLzje2_1(.dout(w_dff_A_hFXxqUvB9_1),.din(w_dff_A_ACcCLzje2_1),.clk(gclk));
	jdff dff_A_aPtPo35h4_1(.dout(w_dff_A_ACcCLzje2_1),.din(w_dff_A_aPtPo35h4_1),.clk(gclk));
	jdff dff_A_3LW8RjDF0_1(.dout(w_dff_A_aPtPo35h4_1),.din(w_dff_A_3LW8RjDF0_1),.clk(gclk));
	jdff dff_A_Zoh4t3ou5_1(.dout(w_dff_A_3LW8RjDF0_1),.din(w_dff_A_Zoh4t3ou5_1),.clk(gclk));
	jdff dff_A_lv4hDV2y3_1(.dout(w_dff_A_Zoh4t3ou5_1),.din(w_dff_A_lv4hDV2y3_1),.clk(gclk));
	jdff dff_A_cdXJ55VL2_1(.dout(w_dff_A_lv4hDV2y3_1),.din(w_dff_A_cdXJ55VL2_1),.clk(gclk));
	jdff dff_A_7ZANJyQm1_1(.dout(w_dff_A_cdXJ55VL2_1),.din(w_dff_A_7ZANJyQm1_1),.clk(gclk));
	jdff dff_A_BYVEcj0V7_1(.dout(w_dff_A_7ZANJyQm1_1),.din(w_dff_A_BYVEcj0V7_1),.clk(gclk));
	jdff dff_A_OAKd8djJ0_1(.dout(w_dff_A_BYVEcj0V7_1),.din(w_dff_A_OAKd8djJ0_1),.clk(gclk));
	jdff dff_A_uUhV7zC25_1(.dout(w_dff_A_OAKd8djJ0_1),.din(w_dff_A_uUhV7zC25_1),.clk(gclk));
	jdff dff_A_JY1X5m9b9_1(.dout(w_dff_A_uUhV7zC25_1),.din(w_dff_A_JY1X5m9b9_1),.clk(gclk));
	jdff dff_A_AX76BrwG9_2(.dout(w_G56gat_0[2]),.din(w_dff_A_AX76BrwG9_2),.clk(gclk));
	jdff dff_A_mORhmi6x1_2(.dout(w_dff_A_AX76BrwG9_2),.din(w_dff_A_mORhmi6x1_2),.clk(gclk));
	jdff dff_A_RIabsRvN7_2(.dout(w_dff_A_mORhmi6x1_2),.din(w_dff_A_RIabsRvN7_2),.clk(gclk));
	jdff dff_A_BkjMFss80_2(.dout(w_dff_A_RIabsRvN7_2),.din(w_dff_A_BkjMFss80_2),.clk(gclk));
	jdff dff_A_fue3WWkf4_2(.dout(w_dff_A_BkjMFss80_2),.din(w_dff_A_fue3WWkf4_2),.clk(gclk));
	jdff dff_A_7zXDXjEg5_2(.dout(w_dff_A_fue3WWkf4_2),.din(w_dff_A_7zXDXjEg5_2),.clk(gclk));
	jdff dff_A_44uiDhtB2_2(.dout(w_dff_A_7zXDXjEg5_2),.din(w_dff_A_44uiDhtB2_2),.clk(gclk));
	jdff dff_A_LSu6I9x51_0(.dout(w_G50gat_0[0]),.din(w_dff_A_LSu6I9x51_0),.clk(gclk));
	jdff dff_A_qpziZNcy2_0(.dout(w_n78_0[0]),.din(w_dff_A_qpziZNcy2_0),.clk(gclk));
	jdff dff_A_iw44Z7qf6_0(.dout(w_dff_A_qpziZNcy2_0),.din(w_dff_A_iw44Z7qf6_0),.clk(gclk));
	jdff dff_A_uUu8MmDp4_0(.dout(w_dff_A_iw44Z7qf6_0),.din(w_dff_A_uUu8MmDp4_0),.clk(gclk));
	jdff dff_A_6GlWTpt34_0(.dout(w_dff_A_uUu8MmDp4_0),.din(w_dff_A_6GlWTpt34_0),.clk(gclk));
	jdff dff_A_hWUgsm1k8_0(.dout(w_dff_A_6GlWTpt34_0),.din(w_dff_A_hWUgsm1k8_0),.clk(gclk));
	jdff dff_A_xqQlZuPp8_0(.dout(w_dff_A_hWUgsm1k8_0),.din(w_dff_A_xqQlZuPp8_0),.clk(gclk));
	jdff dff_A_vCnhxTSl9_0(.dout(w_G30gat_0[0]),.din(w_dff_A_vCnhxTSl9_0),.clk(gclk));
	jdff dff_A_BbHUDA3K2_0(.dout(w_dff_A_vCnhxTSl9_0),.din(w_dff_A_BbHUDA3K2_0),.clk(gclk));
	jdff dff_A_symnjcGt7_0(.dout(w_dff_A_BbHUDA3K2_0),.din(w_dff_A_symnjcGt7_0),.clk(gclk));
	jdff dff_A_enQQQfPp0_0(.dout(w_dff_A_symnjcGt7_0),.din(w_dff_A_enQQQfPp0_0),.clk(gclk));
	jdff dff_A_GkBPbcJL9_0(.dout(w_dff_A_enQQQfPp0_0),.din(w_dff_A_GkBPbcJL9_0),.clk(gclk));
	jdff dff_A_vhNZFhO60_0(.dout(w_dff_A_GkBPbcJL9_0),.din(w_dff_A_vhNZFhO60_0),.clk(gclk));
	jdff dff_A_lHGipaW45_0(.dout(w_dff_A_vhNZFhO60_0),.din(w_dff_A_lHGipaW45_0),.clk(gclk));
	jdff dff_A_40KTVuz15_2(.dout(w_G30gat_0[2]),.din(w_dff_A_40KTVuz15_2),.clk(gclk));
	jdff dff_A_7i6jMMSp3_0(.dout(w_G24gat_0[0]),.din(w_dff_A_7i6jMMSp3_0),.clk(gclk));
	jdff dff_A_pHMOnJ296_0(.dout(w_dff_A_7i6jMMSp3_0),.din(w_dff_A_pHMOnJ296_0),.clk(gclk));
	jdff dff_A_Y3MK6xy55_0(.dout(w_dff_A_pHMOnJ296_0),.din(w_dff_A_Y3MK6xy55_0),.clk(gclk));
	jdff dff_A_vuklsGmU3_0(.dout(w_dff_A_Y3MK6xy55_0),.din(w_dff_A_vuklsGmU3_0),.clk(gclk));
	jdff dff_A_fRqyKCxj7_0(.dout(w_dff_A_vuklsGmU3_0),.din(w_dff_A_fRqyKCxj7_0),.clk(gclk));
	jdff dff_A_FQ25SIfu6_0(.dout(w_dff_A_fRqyKCxj7_0),.din(w_dff_A_FQ25SIfu6_0),.clk(gclk));
	jdff dff_A_dvXEuoOL4_1(.dout(w_G24gat_0[1]),.din(w_dff_A_dvXEuoOL4_1),.clk(gclk));
	jdff dff_A_WXFm6dcW9_0(.dout(w_n75_0[0]),.din(w_dff_A_WXFm6dcW9_0),.clk(gclk));
	jdff dff_A_H1Oe7Lxx9_0(.dout(w_dff_A_WXFm6dcW9_0),.din(w_dff_A_H1Oe7Lxx9_0),.clk(gclk));
	jdff dff_A_lIQ7QlUT2_0(.dout(w_dff_A_H1Oe7Lxx9_0),.din(w_dff_A_lIQ7QlUT2_0),.clk(gclk));
	jdff dff_A_TU3Lkj7o5_0(.dout(w_dff_A_lIQ7QlUT2_0),.din(w_dff_A_TU3Lkj7o5_0),.clk(gclk));
	jdff dff_A_RQEZTEaR6_0(.dout(w_dff_A_TU3Lkj7o5_0),.din(w_dff_A_RQEZTEaR6_0),.clk(gclk));
	jdff dff_A_04nxMYQk2_0(.dout(w_dff_A_RQEZTEaR6_0),.din(w_dff_A_04nxMYQk2_0),.clk(gclk));
	jdff dff_A_oSiZ7gDT6_0(.dout(w_G17gat_0[0]),.din(w_dff_A_oSiZ7gDT6_0),.clk(gclk));
	jdff dff_A_v169T4Al7_0(.dout(w_dff_A_oSiZ7gDT6_0),.din(w_dff_A_v169T4Al7_0),.clk(gclk));
	jdff dff_A_DjWzpirg1_0(.dout(w_dff_A_v169T4Al7_0),.din(w_dff_A_DjWzpirg1_0),.clk(gclk));
	jdff dff_A_Vcwr5R3U8_0(.dout(w_dff_A_DjWzpirg1_0),.din(w_dff_A_Vcwr5R3U8_0),.clk(gclk));
	jdff dff_A_RGLphzG85_0(.dout(w_dff_A_Vcwr5R3U8_0),.din(w_dff_A_RGLphzG85_0),.clk(gclk));
	jdff dff_A_zCdpAzNl6_0(.dout(w_dff_A_RGLphzG85_0),.din(w_dff_A_zCdpAzNl6_0),.clk(gclk));
	jdff dff_A_JKbIRbPS4_0(.dout(w_dff_A_zCdpAzNl6_0),.din(w_dff_A_JKbIRbPS4_0),.clk(gclk));
	jdff dff_A_g7v9LeMl6_2(.dout(w_G17gat_0[2]),.din(w_dff_A_g7v9LeMl6_2),.clk(gclk));
	jdff dff_A_rU0gyG9H0_0(.dout(w_G11gat_0[0]),.din(w_dff_A_rU0gyG9H0_0),.clk(gclk));
	jdff dff_A_leS95rAp2_0(.dout(w_dff_A_rU0gyG9H0_0),.din(w_dff_A_leS95rAp2_0),.clk(gclk));
	jdff dff_A_14drUpLn5_0(.dout(w_dff_A_leS95rAp2_0),.din(w_dff_A_14drUpLn5_0),.clk(gclk));
	jdff dff_A_NCk2KTKr1_0(.dout(w_dff_A_14drUpLn5_0),.din(w_dff_A_NCk2KTKr1_0),.clk(gclk));
	jdff dff_A_32vJPTt17_0(.dout(w_dff_A_NCk2KTKr1_0),.din(w_dff_A_32vJPTt17_0),.clk(gclk));
	jdff dff_A_JFAWom510_0(.dout(w_dff_A_32vJPTt17_0),.din(w_dff_A_JFAWom510_0),.clk(gclk));
	jdff dff_A_ZaaPI5mR8_1(.dout(w_G11gat_0[1]),.din(w_dff_A_ZaaPI5mR8_1),.clk(gclk));
	jdff dff_A_y4VQOozV3_0(.dout(w_n73_0[0]),.din(w_dff_A_y4VQOozV3_0),.clk(gclk));
	jdff dff_A_1HbrcX0L3_0(.dout(w_dff_A_y4VQOozV3_0),.din(w_dff_A_1HbrcX0L3_0),.clk(gclk));
	jdff dff_A_18hYKMe90_0(.dout(w_dff_A_1HbrcX0L3_0),.din(w_dff_A_18hYKMe90_0),.clk(gclk));
	jdff dff_A_led2SLno8_0(.dout(w_dff_A_18hYKMe90_0),.din(w_dff_A_led2SLno8_0),.clk(gclk));
	jdff dff_A_fnDq3uBZ4_0(.dout(w_dff_A_led2SLno8_0),.din(w_dff_A_fnDq3uBZ4_0),.clk(gclk));
	jdff dff_A_o9rGKiMQ7_0(.dout(w_dff_A_fnDq3uBZ4_0),.din(w_dff_A_o9rGKiMQ7_0),.clk(gclk));
	jdff dff_A_VJLj8OIH7_0(.dout(w_G69gat_0[0]),.din(w_dff_A_VJLj8OIH7_0),.clk(gclk));
	jdff dff_A_O0q0vL7x6_0(.dout(w_dff_A_VJLj8OIH7_0),.din(w_dff_A_O0q0vL7x6_0),.clk(gclk));
	jdff dff_A_pm26wIVv4_0(.dout(w_dff_A_O0q0vL7x6_0),.din(w_dff_A_pm26wIVv4_0),.clk(gclk));
	jdff dff_A_VrOYItL46_0(.dout(w_dff_A_pm26wIVv4_0),.din(w_dff_A_VrOYItL46_0),.clk(gclk));
	jdff dff_A_7fkpechI8_0(.dout(w_dff_A_VrOYItL46_0),.din(w_dff_A_7fkpechI8_0),.clk(gclk));
	jdff dff_A_SPyXB4iA3_0(.dout(w_dff_A_7fkpechI8_0),.din(w_dff_A_SPyXB4iA3_0),.clk(gclk));
	jdff dff_A_FIg2GCjw0_0(.dout(w_dff_A_SPyXB4iA3_0),.din(w_dff_A_FIg2GCjw0_0),.clk(gclk));
	jdff dff_A_zygFzT2a9_2(.dout(w_G69gat_0[2]),.din(w_dff_A_zygFzT2a9_2),.clk(gclk));
	jdff dff_A_6UFmeu6I1_0(.dout(w_n46_0[0]),.din(w_dff_A_6UFmeu6I1_0),.clk(gclk));
	jdff dff_A_aqlBCmgJ9_0(.dout(w_dff_A_6UFmeu6I1_0),.din(w_dff_A_aqlBCmgJ9_0),.clk(gclk));
	jdff dff_A_6z0DgTKQ3_0(.dout(w_dff_A_aqlBCmgJ9_0),.din(w_dff_A_6z0DgTKQ3_0),.clk(gclk));
	jdff dff_A_wYaukfJb9_0(.dout(w_dff_A_6z0DgTKQ3_0),.din(w_dff_A_wYaukfJb9_0),.clk(gclk));
	jdff dff_A_A7eitZZH2_1(.dout(w_n46_0[1]),.din(w_dff_A_A7eitZZH2_1),.clk(gclk));
	jdff dff_B_xuLP8Eh94_1(.din(G37gat),.dout(w_dff_B_xuLP8Eh94_1),.clk(gclk));
	jdff dff_A_bgam7PBe5_0(.dout(w_n45_0[0]),.din(w_dff_A_bgam7PBe5_0),.clk(gclk));
	jdff dff_A_36kQpSaL0_0(.dout(w_dff_A_bgam7PBe5_0),.din(w_dff_A_36kQpSaL0_0),.clk(gclk));
	jdff dff_A_scUcDVEG6_0(.dout(w_dff_A_36kQpSaL0_0),.din(w_dff_A_scUcDVEG6_0),.clk(gclk));
	jdff dff_A_YuXhJ4Um4_0(.dout(w_dff_A_scUcDVEG6_0),.din(w_dff_A_YuXhJ4Um4_0),.clk(gclk));
	jdff dff_A_N5gcFe2e7_0(.dout(w_dff_A_YuXhJ4Um4_0),.din(w_dff_A_N5gcFe2e7_0),.clk(gclk));
	jdff dff_A_geBB4Qix9_0(.dout(w_dff_A_N5gcFe2e7_0),.din(w_dff_A_geBB4Qix9_0),.clk(gclk));
	jdff dff_A_Lejslc591_0(.dout(w_G43gat_0[0]),.din(w_dff_A_Lejslc591_0),.clk(gclk));
	jdff dff_A_zHlzfzZr8_0(.dout(w_dff_A_Lejslc591_0),.din(w_dff_A_zHlzfzZr8_0),.clk(gclk));
	jdff dff_A_1NvjaUSz2_0(.dout(w_dff_A_zHlzfzZr8_0),.din(w_dff_A_1NvjaUSz2_0),.clk(gclk));
	jdff dff_A_qeepUeHI8_0(.dout(w_dff_A_1NvjaUSz2_0),.din(w_dff_A_qeepUeHI8_0),.clk(gclk));
	jdff dff_A_gP9kfPVD8_0(.dout(w_dff_A_qeepUeHI8_0),.din(w_dff_A_gP9kfPVD8_0),.clk(gclk));
	jdff dff_A_zX5oOBHJ6_0(.dout(w_dff_A_gP9kfPVD8_0),.din(w_dff_A_zX5oOBHJ6_0),.clk(gclk));
	jdff dff_A_OUEB5VwY0_0(.dout(w_dff_A_zX5oOBHJ6_0),.din(w_dff_A_OUEB5VwY0_0),.clk(gclk));
	jdff dff_A_JTuJefEr1_1(.dout(w_n44_0[1]),.din(w_dff_A_JTuJefEr1_1),.clk(gclk));
	jdff dff_A_Gwj2RSvC4_1(.dout(w_G108gat_0[1]),.din(w_dff_A_Gwj2RSvC4_1),.clk(gclk));
	jdff dff_A_j9sEVpXg1_1(.dout(w_dff_A_Gwj2RSvC4_1),.din(w_dff_A_j9sEVpXg1_1),.clk(gclk));
	jdff dff_A_8CuQWF2Y1_1(.dout(w_dff_A_j9sEVpXg1_1),.din(w_dff_A_8CuQWF2Y1_1),.clk(gclk));
	jdff dff_A_3klM5Thu5_1(.dout(w_dff_A_8CuQWF2Y1_1),.din(w_dff_A_3klM5Thu5_1),.clk(gclk));
	jdff dff_A_wGrMbDhJ8_1(.dout(w_dff_A_3klM5Thu5_1),.din(w_dff_A_wGrMbDhJ8_1),.clk(gclk));
	jdff dff_A_7iDJK7nM3_1(.dout(w_dff_A_wGrMbDhJ8_1),.din(w_dff_A_7iDJK7nM3_1),.clk(gclk));
	jdff dff_A_hFEby3nc2_1(.dout(w_dff_A_7iDJK7nM3_1),.din(w_dff_A_hFEby3nc2_1),.clk(gclk));
	jdff dff_A_rqEwo9jn8_2(.dout(w_G108gat_0[2]),.din(w_dff_A_rqEwo9jn8_2),.clk(gclk));
	jdff dff_A_sZeNBXuB3_0(.dout(w_n43_0[0]),.din(w_dff_A_sZeNBXuB3_0),.clk(gclk));
	jdff dff_A_K0G9mO477_0(.dout(w_dff_A_sZeNBXuB3_0),.din(w_dff_A_K0G9mO477_0),.clk(gclk));
	jdff dff_A_xdj6fnjM7_0(.dout(w_dff_A_K0G9mO477_0),.din(w_dff_A_xdj6fnjM7_0),.clk(gclk));
	jdff dff_A_B9arFAoA0_0(.dout(w_dff_A_xdj6fnjM7_0),.din(w_dff_A_B9arFAoA0_0),.clk(gclk));
	jdff dff_A_xizCi96C2_0(.dout(w_dff_A_B9arFAoA0_0),.din(w_dff_A_xizCi96C2_0),.clk(gclk));
	jdff dff_A_8Lux3dRq9_0(.dout(w_G102gat_0[0]),.din(w_dff_A_8Lux3dRq9_0),.clk(gclk));
	jdff dff_A_1PGOAz6p4_0(.dout(w_dff_A_8Lux3dRq9_0),.din(w_dff_A_1PGOAz6p4_0),.clk(gclk));
	jdff dff_A_jfgelKNm7_0(.dout(w_dff_A_1PGOAz6p4_0),.din(w_dff_A_jfgelKNm7_0),.clk(gclk));
	jdff dff_A_v1AH5uDF5_0(.dout(w_dff_A_jfgelKNm7_0),.din(w_dff_A_v1AH5uDF5_0),.clk(gclk));
	jdff dff_A_Xnm3G1324_0(.dout(w_dff_A_v1AH5uDF5_0),.din(w_dff_A_Xnm3G1324_0),.clk(gclk));
	jdff dff_A_hTDcbTfE3_0(.dout(w_dff_A_Xnm3G1324_0),.din(w_dff_A_hTDcbTfE3_0),.clk(gclk));
	jdff dff_A_Vx6xWK0C8_0(.dout(w_n49_0[0]),.din(w_dff_A_Vx6xWK0C8_0),.clk(gclk));
	jdff dff_A_x36w9jM47_0(.dout(w_dff_A_Vx6xWK0C8_0),.din(w_dff_A_x36w9jM47_0),.clk(gclk));
	jdff dff_A_UTPgT86y3_0(.dout(w_dff_A_x36w9jM47_0),.din(w_dff_A_UTPgT86y3_0),.clk(gclk));
	jdff dff_A_7jISbaM68_0(.dout(w_dff_A_UTPgT86y3_0),.din(w_dff_A_7jISbaM68_0),.clk(gclk));
	jdff dff_A_fIPF64IO4_0(.dout(w_dff_A_7jISbaM68_0),.din(w_dff_A_fIPF64IO4_0),.clk(gclk));
	jdff dff_A_cev2CjdC9_0(.dout(w_G63gat_0[0]),.din(w_dff_A_cev2CjdC9_0),.clk(gclk));
	jdff dff_A_XGjrlVQB2_0(.dout(w_dff_A_cev2CjdC9_0),.din(w_dff_A_XGjrlVQB2_0),.clk(gclk));
	jdff dff_A_UzbiHO6K5_0(.dout(w_dff_A_XGjrlVQB2_0),.din(w_dff_A_UzbiHO6K5_0),.clk(gclk));
	jdff dff_A_yhMk9iiA4_0(.dout(w_dff_A_UzbiHO6K5_0),.din(w_dff_A_yhMk9iiA4_0),.clk(gclk));
	jdff dff_A_P4Fkf42Z9_0(.dout(w_dff_A_yhMk9iiA4_0),.din(w_dff_A_P4Fkf42Z9_0),.clk(gclk));
	jdff dff_A_xttPJG3s4_0(.dout(w_dff_A_P4Fkf42Z9_0),.din(w_dff_A_xttPJG3s4_0),.clk(gclk));
	jdff dff_A_xbIUcwZn2_1(.dout(w_G63gat_0[1]),.din(w_dff_A_xbIUcwZn2_1),.clk(gclk));
	jdff dff_A_YfPI2v904_1(.dout(w_dff_A_njh5mEWr0_0),.din(w_dff_A_YfPI2v904_1),.clk(gclk));
	jdff dff_A_njh5mEWr0_0(.dout(w_dff_A_oQwh5ee35_0),.din(w_dff_A_njh5mEWr0_0),.clk(gclk));
	jdff dff_A_oQwh5ee35_0(.dout(w_dff_A_ukaMzAcL2_0),.din(w_dff_A_oQwh5ee35_0),.clk(gclk));
	jdff dff_A_ukaMzAcL2_0(.dout(w_dff_A_hatnZ07Q8_0),.din(w_dff_A_ukaMzAcL2_0),.clk(gclk));
	jdff dff_A_hatnZ07Q8_0(.dout(w_dff_A_nBB38dso0_0),.din(w_dff_A_hatnZ07Q8_0),.clk(gclk));
	jdff dff_A_nBB38dso0_0(.dout(w_dff_A_3DSdJ4Sk0_0),.din(w_dff_A_nBB38dso0_0),.clk(gclk));
	jdff dff_A_3DSdJ4Sk0_0(.dout(w_dff_A_HtasaU2e2_0),.din(w_dff_A_3DSdJ4Sk0_0),.clk(gclk));
	jdff dff_A_HtasaU2e2_0(.dout(w_dff_A_7ldb0iwp0_0),.din(w_dff_A_HtasaU2e2_0),.clk(gclk));
	jdff dff_A_7ldb0iwp0_0(.dout(w_dff_A_u5eVZI6s5_0),.din(w_dff_A_7ldb0iwp0_0),.clk(gclk));
	jdff dff_A_u5eVZI6s5_0(.dout(w_dff_A_lBlkwG4Y0_0),.din(w_dff_A_u5eVZI6s5_0),.clk(gclk));
	jdff dff_A_lBlkwG4Y0_0(.dout(w_dff_A_Et6fxDxo6_0),.din(w_dff_A_lBlkwG4Y0_0),.clk(gclk));
	jdff dff_A_Et6fxDxo6_0(.dout(w_dff_A_cQJbJjac7_0),.din(w_dff_A_Et6fxDxo6_0),.clk(gclk));
	jdff dff_A_cQJbJjac7_0(.dout(w_dff_A_W91orP1H0_0),.din(w_dff_A_cQJbJjac7_0),.clk(gclk));
	jdff dff_A_W91orP1H0_0(.dout(w_dff_A_0wake6Zx2_0),.din(w_dff_A_W91orP1H0_0),.clk(gclk));
	jdff dff_A_0wake6Zx2_0(.dout(w_dff_A_WrNNn8z30_0),.din(w_dff_A_0wake6Zx2_0),.clk(gclk));
	jdff dff_A_WrNNn8z30_0(.dout(w_dff_A_jOKJLA681_0),.din(w_dff_A_WrNNn8z30_0),.clk(gclk));
	jdff dff_A_jOKJLA681_0(.dout(w_dff_A_tGJMAIzP5_0),.din(w_dff_A_jOKJLA681_0),.clk(gclk));
	jdff dff_A_tGJMAIzP5_0(.dout(w_dff_A_T1BD899E4_0),.din(w_dff_A_tGJMAIzP5_0),.clk(gclk));
	jdff dff_A_T1BD899E4_0(.dout(w_dff_A_vEBV3Mnq0_0),.din(w_dff_A_T1BD899E4_0),.clk(gclk));
	jdff dff_A_vEBV3Mnq0_0(.dout(w_dff_A_GdmBcFZY3_0),.din(w_dff_A_vEBV3Mnq0_0),.clk(gclk));
	jdff dff_A_GdmBcFZY3_0(.dout(G223gat),.din(w_dff_A_GdmBcFZY3_0),.clk(gclk));
	jdff dff_A_zslZLxxx2_1(.dout(w_dff_A_fgKGFq3v6_0),.din(w_dff_A_zslZLxxx2_1),.clk(gclk));
	jdff dff_A_fgKGFq3v6_0(.dout(w_dff_A_bCeJejtr7_0),.din(w_dff_A_fgKGFq3v6_0),.clk(gclk));
	jdff dff_A_bCeJejtr7_0(.dout(w_dff_A_YvxgP7e18_0),.din(w_dff_A_bCeJejtr7_0),.clk(gclk));
	jdff dff_A_YvxgP7e18_0(.dout(w_dff_A_t7G4EAm29_0),.din(w_dff_A_YvxgP7e18_0),.clk(gclk));
	jdff dff_A_t7G4EAm29_0(.dout(w_dff_A_DsxUjxth7_0),.din(w_dff_A_t7G4EAm29_0),.clk(gclk));
	jdff dff_A_DsxUjxth7_0(.dout(w_dff_A_othRQFY30_0),.din(w_dff_A_DsxUjxth7_0),.clk(gclk));
	jdff dff_A_othRQFY30_0(.dout(w_dff_A_k0587dBx3_0),.din(w_dff_A_othRQFY30_0),.clk(gclk));
	jdff dff_A_k0587dBx3_0(.dout(w_dff_A_fyuhdg9T0_0),.din(w_dff_A_k0587dBx3_0),.clk(gclk));
	jdff dff_A_fyuhdg9T0_0(.dout(w_dff_A_gOXwcJzZ9_0),.din(w_dff_A_fyuhdg9T0_0),.clk(gclk));
	jdff dff_A_gOXwcJzZ9_0(.dout(w_dff_A_bJyxZgMB5_0),.din(w_dff_A_gOXwcJzZ9_0),.clk(gclk));
	jdff dff_A_bJyxZgMB5_0(.dout(w_dff_A_iTSAjUzA0_0),.din(w_dff_A_bJyxZgMB5_0),.clk(gclk));
	jdff dff_A_iTSAjUzA0_0(.dout(w_dff_A_t8OamHmj4_0),.din(w_dff_A_iTSAjUzA0_0),.clk(gclk));
	jdff dff_A_t8OamHmj4_0(.dout(w_dff_A_PlgHKSDr8_0),.din(w_dff_A_t8OamHmj4_0),.clk(gclk));
	jdff dff_A_PlgHKSDr8_0(.dout(G329gat),.din(w_dff_A_PlgHKSDr8_0),.clk(gclk));
	jdff dff_A_pATUosgy8_2(.dout(w_dff_A_v8jZ1EzT4_0),.din(w_dff_A_pATUosgy8_2),.clk(gclk));
	jdff dff_A_v8jZ1EzT4_0(.dout(w_dff_A_24bsNqOf1_0),.din(w_dff_A_v8jZ1EzT4_0),.clk(gclk));
	jdff dff_A_24bsNqOf1_0(.dout(w_dff_A_ZuZ75MTa6_0),.din(w_dff_A_24bsNqOf1_0),.clk(gclk));
	jdff dff_A_ZuZ75MTa6_0(.dout(w_dff_A_cnKnaLTX0_0),.din(w_dff_A_ZuZ75MTa6_0),.clk(gclk));
	jdff dff_A_cnKnaLTX0_0(.dout(w_dff_A_YvfxF16g4_0),.din(w_dff_A_cnKnaLTX0_0),.clk(gclk));
	jdff dff_A_YvfxF16g4_0(.dout(w_dff_A_Zx3vGH9S5_0),.din(w_dff_A_YvfxF16g4_0),.clk(gclk));
	jdff dff_A_Zx3vGH9S5_0(.dout(G370gat),.din(w_dff_A_Zx3vGH9S5_0),.clk(gclk));
	jdff dff_A_U0JIoQ1W4_1(.dout(w_dff_A_ICoZLC8m9_0),.din(w_dff_A_U0JIoQ1W4_1),.clk(gclk));
	jdff dff_A_ICoZLC8m9_0(.dout(G430gat),.din(w_dff_A_ICoZLC8m9_0),.clk(gclk));
endmodule

