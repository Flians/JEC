// Benchmark "top" written by ABC on Thu May 28 22:00:27 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] ;
  wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
    n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
    n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
    n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
    n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
    n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
    n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
    n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
    n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
    n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
    n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
    n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
    n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
    n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
    n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
    n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
    n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
    n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
    n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
    n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
    n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
    n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
    n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
    n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
    n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
    n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
    n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
    n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
    n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
    n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
    n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
    n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
    n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
    n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
    n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
    n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
    n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
    n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
    n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
    n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
    n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
    n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
    n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
    n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
    n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
    n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
    n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
    n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
    n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
    n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
    n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
    n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
    n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
    n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
    n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
    n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
    n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
    n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
    n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
    n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
    n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
    n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
    n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
    n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
    n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
    n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
    n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
    n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
    n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
    n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
    n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
    n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
    n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
    n6864, n6865, n6866, n6867, n6868, n6871, n6872, n6873, n6874, n6875,
    n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
    n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
    n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
    n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
    n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
    n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
    n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
    n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
    n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
    n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
    n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
    n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
    n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
    n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
    n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
    n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
    n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
    n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
    n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
    n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
    n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
    n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
    n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
    n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
    n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
    n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
    n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
    n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
    n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
    n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
    n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
    n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
    n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
    n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
    n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
    n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
    n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
    n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
    n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
    n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
    n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
    n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
    n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
    n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
    n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
    n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
    n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
    n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
    n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
    n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
    n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
    n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
    n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
    n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
    n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
    n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
    n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
    n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
    n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
    n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
    n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
    n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
    n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
    n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
    n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
    n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
    n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
    n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
    n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
    n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
    n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
    n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
    n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
    n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
    n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
    n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
    n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
    n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
    n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
    n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
    n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
    n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
    n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
    n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
    n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
    n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
    n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
    n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
    n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
    n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
    n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
    n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
    n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
    n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
    n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
    n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
    n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
    n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
    n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
    n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
    n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
    n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
    n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
    n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
    n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
    n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
    n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
    n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
    n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
    n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
    n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
    n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
    n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
    n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
    n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
    n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
    n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
    n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
    n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
    n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
    n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
    n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
    n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
    n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
    n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
    n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
    n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
    n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
    n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
    n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
    n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
    n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
    n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
    n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
    n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
    n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
    n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
    n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
    n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
    n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
    n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
    n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
    n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
    n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
    n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
    n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
    n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
    n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
    n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
    n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
    n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
    n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
    n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
    n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
    n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
    n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
    n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
    n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
    n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
    n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
    n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
    n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
    n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
    n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
    n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
    n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
    n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
    n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
    n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
    n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
    n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
    n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
    n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
    n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
    n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
    n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
    n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
    n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
    n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
    n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
    n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
    n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
    n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
    n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
    n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
    n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
    n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
    n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
    n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
    n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
    n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
    n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
    n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
    n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
    n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
    n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
    n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
    n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
    n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
    n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
    n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
    n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
    n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
    n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
    n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
    n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
    n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
    n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
    n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
    n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
    n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
    n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
    n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
    n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
    n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
    n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
    n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
    n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
    n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
    n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
    n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
    n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
    n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
    n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
    n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
    n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
    n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
    n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
    n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
    n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
    n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
    n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
    n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
    n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
    n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
    n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
    n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
    n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
    n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
    n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
    n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
    n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
    n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
    n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
    n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
    n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
    n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
    n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
    n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
    n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
    n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
    n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
    n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
    n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
    n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
    n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
    n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
    n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
    n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
    n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
    n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
    n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
    n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
    n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
    n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
    n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
    n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
    n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
    n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
    n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
    n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
    n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
    n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
    n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
    n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
    n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
    n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
    n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
    n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
    n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
    n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
    n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
    n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
    n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
    n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
    n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
    n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
    n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
    n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
    n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
    n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
    n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
    n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
    n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
    n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
    n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
    n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
    n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
    n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
    n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
    n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
    n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
    n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
    n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
    n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
    n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
    n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
    n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
    n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
    n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
    n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
    n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
    n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
    n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
    n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
    n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
    n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
    n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
    n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
    n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
    n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
    n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
    n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
    n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
    n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
    n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
    n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
    n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
    n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
    n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
    n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
    n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
    n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
    n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
    n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
    n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
    n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
    n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
    n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
    n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
    n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
    n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
    n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
    n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
    n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
    n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
    n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
    n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
    n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
    n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
    n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
    n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
    n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
    n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
    n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
    n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
    n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
    n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
    n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
    n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
    n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
    n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
    n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
    n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
    n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
    n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
    n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
    n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
    n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
    n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
    n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
    n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
    n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
    n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
    n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
    n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
    n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
    n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
    n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
    n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
    n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
    n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
    n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
    n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
    n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
    n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
    n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
    n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
    n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
    n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
    n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
    n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
    n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
    n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
    n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
    n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
    n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
    n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
    n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
    n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
    n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
    n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
    n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
    n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
    n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
    n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
    n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
    n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
    n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
    n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
    n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
    n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
    n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
    n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
    n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
    n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
    n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
    n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
    n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
    n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
    n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
    n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
    n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
    n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
    n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
    n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
    n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
    n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
    n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
    n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
    n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
    n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
    n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
    n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
    n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
    n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
    n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
    n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
    n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
    n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
    n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
    n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
    n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
    n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
    n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
    n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
    n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
    n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
    n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
    n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
    n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
    n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
    n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
    n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
    n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
    n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
    n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
    n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
    n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
    n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
    n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
    n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
    n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
    n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
    n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
    n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
    n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
    n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
    n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
    n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
    n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
    n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
    n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
    n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
    n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
    n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
    n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
    n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
    n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
    n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
    n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
    n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
    n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
    n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
    n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
    n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
    n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
    n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
    n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
    n14885, n14886, n14887, n14888, n14889, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14903, n14904,
    n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
    n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
    n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
    n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
    n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
    n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
    n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
    n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
    n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
    n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
    n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
    n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
    n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
    n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
    n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
    n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
    n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
    n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
    n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
    n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
    n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
    n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
    n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
    n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
    n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
    n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
    n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
    n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
    n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
    n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
    n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
    n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
    n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
    n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
    n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
    n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
    n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
    n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
    n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
    n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
    n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
    n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
    n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
    n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
    n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
    n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
    n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
    n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
    n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
    n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
    n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
    n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
    n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
    n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
    n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
    n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
    n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
    n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
    n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
    n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
    n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
    n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
    n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
    n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
    n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
    n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
    n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
    n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
    n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
    n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
    n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
    n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794, n15796, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
    n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
    n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
    n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
    n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
    n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
    n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
    n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
    n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
    n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
    n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
    n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
    n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
    n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
    n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
    n16070, n16071, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
    n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
    n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
    n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
    n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
    n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
    n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
    n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
    n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
    n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
    n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
    n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
    n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
    n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16339, n16342, n16343, n16344, n16345, n16346, n16347,
    n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
    n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
    n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
    n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
    n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
    n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
    n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
    n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
    n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
    n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
    n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
    n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
    n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
    n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
    n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
    n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
    n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
    n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
    n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
    n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
    n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
    n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16546,
    n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
    n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
    n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
    n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
    n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
    n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
    n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
    n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
    n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
    n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
    n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
    n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
    n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
    n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
    n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
    n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
    n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
    n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
    n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
    n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
    n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
    n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
    n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
    n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
    n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
    n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
    n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
    n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
    n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
    n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
    n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
    n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
    n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
    n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
    n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
    n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
    n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
    n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
    n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
    n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
    n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
    n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
    n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
    n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
    n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
    n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
    n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
    n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17291, n17292,
    n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
    n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
    n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
    n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
    n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
    n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
    n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
    n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
    n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
    n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
    n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
    n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
    n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
    n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
    n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
    n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
    n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
    n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
    n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
    n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
    n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
    n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
    n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
    n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
    n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
    n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
    n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
    n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
    n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
    n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
    n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
    n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
    n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
    n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
    n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
    n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
    n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
    n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
    n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
    n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
    n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
    n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
    n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
    n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
    n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
    n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
    n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
    n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17973, n17974,
    n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
    n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
    n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
    n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
    n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
    n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
    n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
    n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
    n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
    n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
    n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
    n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
    n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
    n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
    n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
    n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
    n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
    n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
    n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
    n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
    n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
    n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
    n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
    n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
    n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
    n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
    n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
    n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
    n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
    n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
    n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
    n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
    n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
    n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
    n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
    n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775, n18781, n18782, n18783,
    n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
    n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
    n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
    n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
    n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
    n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
    n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
    n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
    n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
    n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
    n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
    n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
    n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
    n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
    n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
    n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
    n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
    n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
    n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
    n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
    n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
    n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
    n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
    n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
    n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
    n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
    n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
    n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
    n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
    n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
    n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
    n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
    n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
    n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
    n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
    n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
    n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
    n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
    n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
    n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
    n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
    n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
    n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
    n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
    n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
    n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
    n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
    n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
    n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
    n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
    n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
    n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
    n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
    n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
    n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
    n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
    n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
    n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
    n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
    n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
    n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
    n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
    n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
    n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
    n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
    n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
    n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
    n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
    n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
    n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
    n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
    n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
    n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
    n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
    n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
    n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
    n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
    n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
    n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
    n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
    n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
    n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
    n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
    n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
    n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
    n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
    n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
    n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
    n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
    n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
    n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
    n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
    n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
    n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
    n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
    n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
    n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
    n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
    n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
    n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
    n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
    n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
    n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
    n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
    n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
    n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
    n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
    n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
    n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
    n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
    n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
    n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
    n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
    n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
    n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
    n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
    n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
    n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
    n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
    n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
    n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
    n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
    n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
    n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
    n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
    n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
    n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
    n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
    n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
    n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
    n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
    n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
    n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
    n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
    n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
    n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
    n20041, n20042, n20043, n20044, n20045, n20047, n20048, n20049, n20050,
    n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
    n20060, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
    n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
    n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
    n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
    n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
    n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
    n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
    n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
    n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
    n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
    n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
    n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
    n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
    n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
    n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
    n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
    n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
    n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
    n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
    n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
    n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
    n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
    n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
    n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
    n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
    n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
    n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
    n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
    n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
    n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
    n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
    n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
    n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
    n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
    n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
    n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
    n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
    n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
    n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
    n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
    n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
    n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
    n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
    n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
    n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
    n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
    n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
    n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
    n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
    n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
    n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
    n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
    n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
    n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
    n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
    n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
    n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
    n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
    n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
    n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
    n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
    n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
    n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
    n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
    n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
    n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
    n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
    n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
    n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
    n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
    n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
    n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
    n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
    n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
    n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
    n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
    n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
    n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
    n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
    n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
    n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
    n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
    n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
    n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
    n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
    n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
    n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
    n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
    n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
    n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
    n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
    n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
    n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
    n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
    n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
    n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
    n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
    n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
    n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
    n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
    n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
    n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
    n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
    n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
    n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
    n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
    n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
    n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
    n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
    n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
    n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
    n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
    n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
    n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
    n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
    n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
    n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
    n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
    n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
    n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22192,
    n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
    n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
    n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
    n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
    n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237,
    n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
    n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
    n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
    n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
    n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
    n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
    n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
    n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309,
    n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
    n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
    n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
    n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
    n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
    n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
    n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
    n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381,
    n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
    n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
    n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
    n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
    n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
    n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
    n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
    n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
    n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
    n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
    n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
    n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
    n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
    n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
    n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
    n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
    n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
    n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
    n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
    n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606,
    n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
    n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
    n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
    n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
    n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
    n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
    n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
    n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
    n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
    n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
    n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750,
    n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
    n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
    n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
    n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
    n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
    n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
    n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813,
    n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822,
    n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
    n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
    n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876,
    n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885,
    n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894,
    n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
    n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
    n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
    n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
    n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
    n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948,
    n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
    n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966,
    n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
    n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
    n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
    n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
    n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
    n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020,
    n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
    n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038,
    n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
    n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
    n23057, n23058, n23059, n23060, n23067, n23068, n23069, n23070, n23071,
    n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
    n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
    n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
    n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
    n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
    n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
    n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134,
    n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
    n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
    n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
    n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
    n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
    n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
    n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
    n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
    n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278,
    n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
    n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
    n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332,
    n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350,
    n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
    n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
    n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
    n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
    n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
    n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
    n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
    n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422,
    n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
    n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
    n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
    n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
    n23477, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23491, n23492, n23493, n23494, n23495, n23496,
    n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
    n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
    n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
    n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532,
    n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
    n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550,
    n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
    n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
    n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
    n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
    n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
    n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
    n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
    n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
    n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
    n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,
    n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
    n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
    n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
    n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676,
    n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
    n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
    n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
    n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,
    n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
    n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
    n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
    n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748,
    n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
    n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
    n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
    n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
    n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
    n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
    n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
    n23812, n23813, n23814, n23815, n23816, n23817, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
    n23831, n23832, n23833, n23842, n23843, n23844, n23845, n23846, n23847,
    n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
    n23857, n23858, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
    n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
    n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
    n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
    n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
    n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
    n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
    n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
    n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24089, n24090,
    n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
    n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108,
    n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117,
    n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126,
    n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135,
    n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,
    n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
    n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162,
    n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
    n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180,
    n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189,
    n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198,
    n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207,
    n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
    n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
    n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
    n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
    n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252,
    n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261,
    n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270,
    n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
    n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,
    n24289, n24290, n24291, n24293, n24294, n24295, n24296, n24297, n24298,
    n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
    n24308, n24309, n24310, n24311, n24312, n24313, n24315, n24316, n24317,
    n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
    n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
    n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
    n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
    n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
    n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
    n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
    n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
    n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
    n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494, n24496, n24497, n24498,
    n24499, n24500, n24501, n24503, n24504, n24505, n24506, n24507, n24508,
    n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
    n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
    n24527, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,
    n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
    n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
    n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
    n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572,
    n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581,
    n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590,
    n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
    n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,
    n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
    n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
    n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
    n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644,
    n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653,
    n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662,
    n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
    n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680,
    n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
    n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
    n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
    n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716,
    n24718, n24719, n24720, n24721, n24722, n24723, n24725, n24726, n24727,
    n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
    n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
    n24746, n24747, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
    n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764,
    n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773,
    n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782,
    n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
    n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,
    n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
    n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
    n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
    n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
    n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845,
    n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
    n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
    n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
    n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
    n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
    n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
    n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
    n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917,
    n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
    n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
    n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24945,
    n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
    n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
    n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972,
    n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981,
    n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990,
    n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
    n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
    n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
    n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
    n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
    n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
    n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053,
    n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062,
    n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071,
    n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
    n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
    n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
    n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
    n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116,
    n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125,
    n25126, n25127, n25128, n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
    n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
    n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180,
    n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
    n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
    n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
    n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
    n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
    n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
    n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
    n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252,
    n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
    n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270,
    n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
    n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
    n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
    n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
    n25307, n25308, n25309, n25310, n25311, n25312, n25314, n25315, n25316,
    n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
    n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334,
    n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
    n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
    n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
    n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
    n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
    n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
    n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
    n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
    n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
    n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
    n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
    n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
    n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
    n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
    n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
    n25488, n25489, n25490, n25491, n25492, n25493, n25495, n25496, n25497,
    n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
    n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
    n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524,
    n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533,
    n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542,
    n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551,
    n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
    n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
    n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
    n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
    n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
    n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605,
    n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614,
    n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623,
    n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
    n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
    n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
    n25651, n25652, n25653, n25654, n25655, n25656, n25658, n25659, n25660,
    n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678,
    n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
    n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
    n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
    n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
    n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
    n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
    n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
    n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25820, n25821, n25822, n25823,
    n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
    n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
    n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
    n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
    n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
    n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
    n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
    n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
    n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
    n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
    n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
    n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
    n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
    n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
    n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
    n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
    n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
    n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
    n25986, n25987, n25988, n25989, n25990, n25991, n25993, n25994, n25995,
    n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004,
    n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013,
    n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022,
    n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031,
    n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
    n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
    n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
    n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
    n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076,
    n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
    n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094,
    n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
    n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
    n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
    n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
    n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
    n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148,
    n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
    n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
    n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
    n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
    n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
    n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
    n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
    n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
    n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26302, n26303,
    n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
    n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
    n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
    n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
    n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348,
    n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357,
    n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366,
    n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
    n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
    n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
    n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
    n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
    n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420,
    n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429,
    n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438,
    n26439, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
    n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
    n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
    n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
    n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484,
    n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493,
    n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502,
    n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
    n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,
    n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
    n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
    n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
    n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556,
    n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565,
    n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574,
    n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26583, n26584,
    n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
    n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
    n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638,
    n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
    n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
    n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
    n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
    n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
    n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
    n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
    n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
    n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
    n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
    n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
    n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
    n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26846, n26847,
    n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
    n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
    n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
    n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
    n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
    n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
    n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910,
    n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
    n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,
    n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
    n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
    n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
    n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964,
    n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
    n26974, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
    n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
    n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
    n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046,
    n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
    n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
    n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
    n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101,
    n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110,
    n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119,
    n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
    n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
    n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
    n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
    n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
    n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
    n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182,
    n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191,
    n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,
    n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27209, n27210,
    n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
    n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228,
    n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237,
    n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246,
    n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255,
    n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264,
    n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
    n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
    n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
    n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
    n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309,
    n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318,
    n27319, n27320, n27322, n27323, n27324, n27325, n27326, n27327, n27328,
    n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
    n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
    n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
    n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
    n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373,
    n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382,
    n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
    n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
    n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
    n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
    n27419, n27420, n27421, n27423, n27424, n27425, n27426, n27427, n27428,
    n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
    n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
    n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
    n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
    n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
    n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
    n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509,
    n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518,
    n27519, n27520, n27521, n27522, n27523, n27525, n27526, n27527, n27528,
    n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
    n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
    n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
    n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
    n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
    n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582,
    n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591,
    n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600,
    n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
    n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
    n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646,
    n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
    n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
    n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
    n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27710,
    n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719,
    n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
    n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
    n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
    n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
    n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
    n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
    n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
    n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
    n27792, n27793, n27794, n27795, n27797, n27798, n27799, n27800, n27801,
    n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
    n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
    n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
    n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
    n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846,
    n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855,
    n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864,
    n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
    n27874, n27875, n27876, n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
    n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
    n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928,
    n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27946, n27947,
    n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
    n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965,
    n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974,
    n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983,
    n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992,
    n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
    n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
    n28011, n28012, n28013, n28014, n28016, n28017, n28018, n28019, n28020,
    n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029,
    n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038,
    n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047,
    n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056,
    n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
    n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
    n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
    n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
    n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116;
  jxor g00000(.dina(\a[27] ), .dinb(\a[26] ), .dout(n64));
  jnot g00001(.din(\a[23] ), .dout(n65));
  jxor g00002(.dina(\a[24] ), .dinb(n65), .dout(n66));
  jnot g00003(.din(n66), .dout(n67));
  jnot g00004(.din(\a[25] ), .dout(n68));
  jxor g00005(.dina(\a[26] ), .dinb(n68), .dout(n69));
  jnot g00006(.din(n69), .dout(n70));
  jand g00007(.dina(n70), .dinb(n67), .dout(n71));
  jnot g00008(.din(\a[27] ), .dout(n72));
  jand g00009(.dina(\a[28] ), .dinb(n72), .dout(n73));
  jnot g00010(.din(\a[30] ), .dout(n74));
  jand g00011(.dina(n74), .dinb(\a[29] ), .dout(n75));
  jand g00012(.dina(n75), .dinb(n73), .dout(n76));
  jnot g00013(.din(\a[26] ), .dout(n77));
  jand g00014(.dina(n77), .dinb(\a[23] ), .dout(n78));
  jand g00015(.dina(\a[25] ), .dinb(\a[24] ), .dout(n79));
  jand g00016(.dina(n79), .dinb(n78), .dout(n80));
  jand g00017(.dina(n80), .dinb(n76), .dout(n81));
  jnot g00018(.din(n81), .dout(n82));
  jnot g00019(.din(\a[24] ), .dout(n83));
  jand g00020(.dina(\a[25] ), .dinb(n83), .dout(n84));
  jand g00021(.dina(n77), .dinb(n65), .dout(n85));
  jand g00022(.dina(n85), .dinb(n84), .dout(n86));
  jnot g00023(.din(\a[28] ), .dout(n87));
  jand g00024(.dina(n87), .dinb(n72), .dout(n88));
  jand g00025(.dina(\a[30] ), .dinb(\a[29] ), .dout(n89));
  jand g00026(.dina(n89), .dinb(n88), .dout(n90));
  jand g00027(.dina(n90), .dinb(n86), .dout(n91));
  jnot g00028(.din(n91), .dout(n92));
  jnot g00029(.din(\a[29] ), .dout(n93));
  jand g00030(.dina(\a[30] ), .dinb(n93), .dout(n94));
  jand g00031(.dina(\a[28] ), .dinb(\a[27] ), .dout(n95));
  jand g00032(.dina(n95), .dinb(n94), .dout(n96));
  jand g00033(.dina(\a[26] ), .dinb(n65), .dout(n97));
  jand g00034(.dina(n97), .dinb(n79), .dout(n98));
  jand g00035(.dina(n98), .dinb(n96), .dout(n99));
  jnot g00036(.din(n99), .dout(n100));
  jand g00037(.dina(n100), .dinb(n92), .dout(n101));
  jor  g00038(.dina(n68), .dinb(n83), .dout(n102));
  jor  g00039(.dina(n77), .dinb(\a[23] ), .dout(n103));
  jor  g00040(.dina(n103), .dinb(n102), .dout(n104));
  jor  g00041(.dina(n87), .dinb(n72), .dout(n105));
  jor  g00042(.dina(\a[30] ), .dinb(\a[29] ), .dout(n106));
  jor  g00043(.dina(n106), .dinb(n105), .dout(n107));
  jor  g00044(.dina(n107), .dinb(n104), .dout(n108));
  jand g00045(.dina(n108), .dinb(n101), .dout(n109));
  jand g00046(.dina(n109), .dinb(n82), .dout(n110));
  jand g00047(.dina(n68), .dinb(\a[24] ), .dout(n111));
  jand g00048(.dina(n111), .dinb(n97), .dout(n112));
  jand g00049(.dina(n112), .dinb(n76), .dout(n113));
  jnot g00050(.din(n113), .dout(n114));
  jor  g00051(.dina(n87), .dinb(\a[27] ), .dout(n115));
  jor  g00052(.dina(\a[30] ), .dinb(n93), .dout(n116));
  jor  g00053(.dina(n116), .dinb(n115), .dout(n117));
  jor  g00054(.dina(\a[26] ), .dinb(n65), .dout(n118));
  jor  g00055(.dina(\a[25] ), .dinb(n83), .dout(n119));
  jor  g00056(.dina(n119), .dinb(n118), .dout(n120));
  jor  g00057(.dina(n120), .dinb(n117), .dout(n121));
  jand g00058(.dina(n121), .dinb(n114), .dout(n122));
  jand g00059(.dina(n122), .dinb(n110), .dout(n123));
  jnot g00060(.din(n123), .dout(n124));
  jand g00061(.dina(n87), .dinb(\a[27] ), .dout(n125));
  jand g00062(.dina(n125), .dinb(n89), .dout(n126));
  jand g00063(.dina(n68), .dinb(n83), .dout(n127));
  jand g00064(.dina(n127), .dinb(n85), .dout(n128));
  jand g00065(.dina(n128), .dinb(n126), .dout(n129));
  jnot g00066(.din(n129), .dout(n130));
  jand g00067(.dina(n96), .dinb(n80), .dout(n131));
  jnot g00068(.din(n131), .dout(n132));
  jand g00069(.dina(n111), .dinb(n85), .dout(n133));
  jand g00070(.dina(n133), .dinb(n76), .dout(n134));
  jnot g00071(.din(n134), .dout(n135));
  jand g00072(.dina(n135), .dinb(n132), .dout(n136));
  jand g00073(.dina(n136), .dinb(n130), .dout(n137));
  jnot g00074(.din(n137), .dout(n138));
  jand g00075(.dina(n85), .dinb(n79), .dout(n139));
  jand g00076(.dina(n125), .dinb(n94), .dout(n140));
  jand g00077(.dina(n140), .dinb(n139), .dout(n141));
  jand g00078(.dina(n74), .dinb(n93), .dout(n142));
  jand g00079(.dina(n125), .dinb(n142), .dout(n143));
  jand g00080(.dina(n97), .dinb(n84), .dout(n144));
  jand g00081(.dina(n144), .dinb(n143), .dout(n145));
  jand g00082(.dina(n142), .dinb(n73), .dout(n146));
  jand g00083(.dina(n146), .dinb(n139), .dout(n147));
  jor  g00084(.dina(n147), .dinb(n145), .dout(n148));
  jand g00085(.dina(n125), .dinb(n75), .dout(n149));
  jand g00086(.dina(n149), .dinb(n86), .dout(n150));
  jor  g00087(.dina(n150), .dinb(n148), .dout(n151));
  jand g00088(.dina(n139), .dinb(n76), .dout(n152));
  jand g00089(.dina(n142), .dinb(n88), .dout(n153));
  jand g00090(.dina(\a[26] ), .dinb(\a[23] ), .dout(n154));
  jand g00091(.dina(n154), .dinb(n127), .dout(n155));
  jand g00092(.dina(n155), .dinb(n153), .dout(n156));
  jor  g00093(.dina(n156), .dinb(n152), .dout(n157));
  jand g00094(.dina(n155), .dinb(n96), .dout(n158));
  jand g00095(.dina(n127), .dinb(n97), .dout(n159));
  jand g00096(.dina(n159), .dinb(n96), .dout(n160));
  jor  g00097(.dina(n160), .dinb(n158), .dout(n161));
  jor  g00098(.dina(n161), .dinb(n157), .dout(n162));
  jor  g00099(.dina(n162), .dinb(n151), .dout(n163));
  jor  g00100(.dina(n163), .dinb(n141), .dout(n164));
  jor  g00101(.dina(n164), .dinb(n138), .dout(n165));
  jand g00102(.dina(n89), .dinb(n73), .dout(n166));
  jand g00103(.dina(n166), .dinb(n80), .dout(n167));
  jnot g00104(.din(n167), .dout(n168));
  jand g00105(.dina(n95), .dinb(n75), .dout(n169));
  jand g00106(.dina(n169), .dinb(n159), .dout(n170));
  jnot g00107(.din(n170), .dout(n171));
  jand g00108(.dina(n171), .dinb(n168), .dout(n172));
  jnot g00109(.din(n172), .dout(n173));
  jand g00110(.dina(n169), .dinb(n128), .dout(n174));
  jnot g00111(.din(n174), .dout(n175));
  jand g00112(.dina(n111), .dinb(n78), .dout(n176));
  jand g00113(.dina(n153), .dinb(n176), .dout(n177));
  jnot g00114(.din(n177), .dout(n178));
  jand g00115(.dina(n178), .dinb(n175), .dout(n179));
  jnot g00116(.din(n179), .dout(n180));
  jand g00117(.dina(n154), .dinb(n111), .dout(n181));
  jand g00118(.dina(n181), .dinb(n90), .dout(n182));
  jand g00119(.dina(n127), .dinb(n78), .dout(n183));
  jand g00120(.dina(n183), .dinb(n96), .dout(n184));
  jor  g00121(.dina(n184), .dinb(n182), .dout(n185));
  jand g00122(.dina(n95), .dinb(n89), .dout(n186));
  jand g00123(.dina(n186), .dinb(n128), .dout(n187));
  jand g00124(.dina(n143), .dinb(n80), .dout(n188));
  jor  g00125(.dina(n188), .dinb(n187), .dout(n189));
  jor  g00126(.dina(n189), .dinb(n185), .dout(n190));
  jor  g00127(.dina(n190), .dinb(n180), .dout(n191));
  jor  g00128(.dina(n191), .dinb(n173), .dout(n192));
  jor  g00129(.dina(n192), .dinb(n165), .dout(n193));
  jand g00130(.dina(n155), .dinb(n143), .dout(n194));
  jand g00131(.dina(n154), .dinb(n84), .dout(n195));
  jand g00132(.dina(n195), .dinb(n153), .dout(n196));
  jand g00133(.dina(n94), .dinb(n73), .dout(n197));
  jand g00134(.dina(n197), .dinb(n139), .dout(n198));
  jand g00135(.dina(n159), .dinb(n149), .dout(n199));
  jor  g00136(.dina(n199), .dinb(n198), .dout(n200));
  jor  g00137(.dina(n200), .dinb(n196), .dout(n201));
  jand g00138(.dina(n149), .dinb(n176), .dout(n202));
  jor  g00139(.dina(n202), .dinb(n201), .dout(n203));
  jor  g00140(.dina(n203), .dinb(n194), .dout(n204));
  jand g00141(.dina(n146), .dinb(n144), .dout(n205));
  jand g00142(.dina(n159), .dinb(n126), .dout(n206));
  jor  g00143(.dina(n206), .dinb(n205), .dout(n207));
  jand g00144(.dina(n197), .dinb(n155), .dout(n208));
  jand g00145(.dina(n94), .dinb(n88), .dout(n209));
  jand g00146(.dina(n209), .dinb(n86), .dout(n210));
  jor  g00147(.dina(n210), .dinb(n208), .dout(n211));
  jand g00148(.dina(n84), .dinb(n78), .dout(n212));
  jand g00149(.dina(n212), .dinb(n90), .dout(n213));
  jor  g00150(.dina(n213), .dinb(n211), .dout(n214));
  jor  g00151(.dina(n214), .dinb(n207), .dout(n215));
  jand g00152(.dina(n183), .dinb(n90), .dout(n216));
  jand g00153(.dina(n143), .dinb(n133), .dout(n217));
  jor  g00154(.dina(n217), .dinb(n216), .dout(n218));
  jand g00155(.dina(n142), .dinb(n95), .dout(n219));
  jand g00156(.dina(n139), .dinb(n219), .dout(n220));
  jand g00157(.dina(n140), .dinb(n128), .dout(n221));
  jor  g00158(.dina(n221), .dinb(n220), .dout(n222));
  jor  g00159(.dina(n222), .dinb(n218), .dout(n223));
  jor  g00160(.dina(n223), .dinb(n215), .dout(n224));
  jor  g00161(.dina(n224), .dinb(n204), .dout(n225));
  jand g00162(.dina(n209), .dinb(n155), .dout(n226));
  jand g00163(.dina(n154), .dinb(n79), .dout(n227));
  jand g00164(.dina(n227), .dinb(n186), .dout(n228));
  jand g00165(.dina(n155), .dinb(n140), .dout(n229));
  jor  g00166(.dina(n229), .dinb(n228), .dout(n230));
  jand g00167(.dina(n169), .dinb(n80), .dout(n231));
  jor  g00168(.dina(n231), .dinb(n230), .dout(n232));
  jor  g00169(.dina(n232), .dinb(n226), .dout(n233));
  jand g00170(.dina(n195), .dinb(n149), .dout(n234));
  jor  g00171(.dina(n234), .dinb(n233), .dout(n235));
  jand g00172(.dina(n143), .dinb(n128), .dout(n236));
  jand g00173(.dina(n212), .dinb(n166), .dout(n237));
  jand g00174(.dina(n166), .dinb(n139), .dout(n238));
  jor  g00175(.dina(n238), .dinb(n237), .dout(n239));
  jor  g00176(.dina(n239), .dinb(n236), .dout(n240));
  jand g00177(.dina(n140), .dinb(n133), .dout(n241));
  jand g00178(.dina(n183), .dinb(n140), .dout(n242));
  jor  g00179(.dina(n242), .dinb(n241), .dout(n243));
  jand g00180(.dina(n209), .dinb(n176), .dout(n244));
  jand g00181(.dina(n227), .dinb(n90), .dout(n245));
  jor  g00182(.dina(n245), .dinb(n244), .dout(n246));
  jor  g00183(.dina(n246), .dinb(n243), .dout(n247));
  jor  g00184(.dina(n247), .dinb(n240), .dout(n248));
  jand g00185(.dina(n166), .dinb(n176), .dout(n249));
  jand g00186(.dina(n186), .dinb(n183), .dout(n250));
  jor  g00187(.dina(n250), .dinb(n249), .dout(n251));
  jand g00188(.dina(n88), .dinb(n75), .dout(n252));
  jand g00189(.dina(n252), .dinb(n159), .dout(n253));
  jand g00190(.dina(n181), .dinb(n76), .dout(n254));
  jor  g00191(.dina(n254), .dinb(n253), .dout(n255));
  jor  g00192(.dina(n255), .dinb(n251), .dout(n256));
  jor  g00193(.dina(n256), .dinb(n248), .dout(n257));
  jor  g00194(.dina(n257), .dinb(n235), .dout(n258));
  jor  g00195(.dina(n258), .dinb(n225), .dout(n259));
  jor  g00196(.dina(n259), .dinb(n193), .dout(n260));
  jor  g00197(.dina(n68), .dinb(\a[24] ), .dout(n261));
  jor  g00198(.dina(\a[26] ), .dinb(\a[23] ), .dout(n262));
  jor  g00199(.dina(n262), .dinb(n261), .dout(n263));
  jor  g00200(.dina(n74), .dinb(n93), .dout(n264));
  jor  g00201(.dina(n105), .dinb(n264), .dout(n265));
  jor  g00202(.dina(n265), .dinb(n263), .dout(n266));
  jor  g00203(.dina(n74), .dinb(\a[29] ), .dout(n267));
  jor  g00204(.dina(n105), .dinb(n267), .dout(n268));
  jor  g00205(.dina(n262), .dinb(n102), .dout(n269));
  jor  g00206(.dina(n269), .dinb(n268), .dout(n270));
  jand g00207(.dina(n270), .dinb(n266), .dout(n271));
  jnot g00208(.din(n271), .dout(n272));
  jand g00209(.dina(n181), .dinb(n219), .dout(n273));
  jand g00210(.dina(n186), .dinb(n159), .dout(n274));
  jand g00211(.dina(n252), .dinb(n139), .dout(n275));
  jor  g00212(.dina(n275), .dinb(n274), .dout(n276));
  jor  g00213(.dina(n276), .dinb(n273), .dout(n277));
  jor  g00214(.dina(n277), .dinb(n272), .dout(n278));
  jand g00215(.dina(n146), .dinb(n98), .dout(n279));
  jand g00216(.dina(n219), .dinb(n86), .dout(n280));
  jand g00217(.dina(n181), .dinb(n169), .dout(n281));
  jor  g00218(.dina(n281), .dinb(n280), .dout(n282));
  jor  g00219(.dina(n282), .dinb(n279), .dout(n283));
  jand g00220(.dina(n133), .dinb(n90), .dout(n284));
  jand g00221(.dina(n227), .dinb(n197), .dout(n285));
  jor  g00222(.dina(n285), .dinb(n284), .dout(n286));
  jand g00223(.dina(n153), .dinb(n144), .dout(n287));
  jand g00224(.dina(n143), .dinb(n139), .dout(n288));
  jor  g00225(.dina(n288), .dinb(n287), .dout(n289));
  jor  g00226(.dina(n289), .dinb(n286), .dout(n290));
  jor  g00227(.dina(n290), .dinb(n283), .dout(n291));
  jor  g00228(.dina(n291), .dinb(n278), .dout(n292));
  jand g00229(.dina(n155), .dinb(n126), .dout(n293));
  jand g00230(.dina(n186), .dinb(n139), .dout(n294));
  jand g00231(.dina(n176), .dinb(n96), .dout(n295));
  jor  g00232(.dina(n295), .dinb(n294), .dout(n296));
  jor  g00233(.dina(n296), .dinb(n293), .dout(n297));
  jand g00234(.dina(n126), .dinb(n86), .dout(n298));
  jand g00235(.dina(n197), .dinb(n86), .dout(n299));
  jor  g00236(.dina(n299), .dinb(n298), .dout(n300));
  jand g00237(.dina(n195), .dinb(n76), .dout(n301));
  jand g00238(.dina(n98), .dinb(n76), .dout(n302));
  jor  g00239(.dina(n302), .dinb(n301), .dout(n303));
  jor  g00240(.dina(n303), .dinb(n300), .dout(n304));
  jor  g00241(.dina(n304), .dinb(n297), .dout(n305));
  jand g00242(.dina(n155), .dinb(n146), .dout(n306));
  jand g00243(.dina(n186), .dinb(n155), .dout(n307));
  jor  g00244(.dina(n307), .dinb(n306), .dout(n308));
  jand g00245(.dina(n197), .dinb(n195), .dout(n309));
  jand g00246(.dina(n209), .dinb(n98), .dout(n310));
  jor  g00247(.dina(n310), .dinb(n309), .dout(n311));
  jand g00248(.dina(n186), .dinb(n144), .dout(n312));
  jand g00249(.dina(n140), .dinb(n98), .dout(n313));
  jor  g00250(.dina(n313), .dinb(n312), .dout(n314));
  jor  g00251(.dina(n314), .dinb(n311), .dout(n315));
  jor  g00252(.dina(n315), .dinb(n308), .dout(n316));
  jor  g00253(.dina(n316), .dinb(n305), .dout(n317));
  jor  g00254(.dina(n317), .dinb(n292), .dout(n318));
  jand g00255(.dina(n149), .dinb(n139), .dout(n319));
  jnot g00256(.din(n319), .dout(n320));
  jor  g00257(.dina(\a[28] ), .dinb(n72), .dout(n321));
  jor  g00258(.dina(n321), .dinb(n116), .dout(n322));
  jor  g00259(.dina(n77), .dinb(n65), .dout(n323));
  jor  g00260(.dina(n323), .dinb(n119), .dout(n324));
  jor  g00261(.dina(n324), .dinb(n322), .dout(n325));
  jand g00262(.dina(n325), .dinb(n320), .dout(n326));
  jand g00263(.dina(n181), .dinb(n166), .dout(n327));
  jnot g00264(.din(n327), .dout(n328));
  jand g00265(.dina(n328), .dinb(n326), .dout(n329));
  jnot g00266(.din(n329), .dout(n330));
  jand g00267(.dina(n252), .dinb(n212), .dout(n331));
  jand g00268(.dina(n252), .dinb(n80), .dout(n332));
  jor  g00269(.dina(n332), .dinb(n331), .dout(n333));
  jand g00270(.dina(n143), .dinb(n98), .dout(n334));
  jand g00271(.dina(n227), .dinb(n169), .dout(n335));
  jand g00272(.dina(n159), .dinb(n76), .dout(n336));
  jor  g00273(.dina(n336), .dinb(n335), .dout(n337));
  jor  g00274(.dina(n337), .dinb(n334), .dout(n338));
  jor  g00275(.dina(n338), .dinb(n333), .dout(n339));
  jand g00276(.dina(n140), .dinb(n112), .dout(n340));
  jand g00277(.dina(n159), .dinb(n219), .dout(n341));
  jand g00278(.dina(n126), .dinb(n176), .dout(n342));
  jor  g00279(.dina(n342), .dinb(n341), .dout(n343));
  jor  g00280(.dina(n343), .dinb(n340), .dout(n344));
  jor  g00281(.dina(n344), .dinb(n339), .dout(n345));
  jor  g00282(.dina(n345), .dinb(n330), .dout(n346));
  jor  g00283(.dina(n346), .dinb(n318), .dout(n347));
  jand g00284(.dina(n209), .dinb(n144), .dout(n348));
  jnot g00285(.din(n348), .dout(n349));
  jand g00286(.dina(n212), .dinb(n76), .dout(n350));
  jnot g00287(.din(n350), .dout(n351));
  jand g00288(.dina(n351), .dinb(n349), .dout(n352));
  jnot g00289(.din(n352), .dout(n353));
  jand g00290(.dina(n197), .dinb(n133), .dout(n354));
  jand g00291(.dina(n252), .dinb(n144), .dout(n355));
  jor  g00292(.dina(n355), .dinb(n354), .dout(n356));
  jand g00293(.dina(n227), .dinb(n76), .dout(n357));
  jor  g00294(.dina(n357), .dinb(n356), .dout(n358));
  jor  g00295(.dina(n358), .dinb(n353), .dout(n359));
  jand g00296(.dina(n197), .dinb(n144), .dout(n360));
  jand g00297(.dina(n181), .dinb(n146), .dout(n361));
  jand g00298(.dina(n181), .dinb(n96), .dout(n362));
  jor  g00299(.dina(n362), .dinb(n361), .dout(n363));
  jor  g00300(.dina(n363), .dinb(n360), .dout(n364));
  jand g00301(.dina(n252), .dinb(n181), .dout(n365));
  jand g00302(.dina(n159), .dinb(n90), .dout(n366));
  jor  g00303(.dina(n366), .dinb(n365), .dout(n367));
  jand g00304(.dina(n149), .dinb(n144), .dout(n368));
  jand g00305(.dina(n197), .dinb(n183), .dout(n369));
  jor  g00306(.dina(n369), .dinb(n368), .dout(n370));
  jor  g00307(.dina(n370), .dinb(n367), .dout(n371));
  jor  g00308(.dina(n371), .dinb(n364), .dout(n372));
  jand g00309(.dina(n146), .dinb(n176), .dout(n373));
  jand g00310(.dina(n169), .dinb(n176), .dout(n374));
  jand g00311(.dina(n96), .dinb(n86), .dout(n375));
  jor  g00312(.dina(n375), .dinb(n374), .dout(n376));
  jor  g00313(.dina(n376), .dinb(n373), .dout(n377));
  jor  g00314(.dina(n377), .dinb(n372), .dout(n378));
  jor  g00315(.dina(n378), .dinb(n359), .dout(n379));
  jand g00316(.dina(n166), .dinb(n112), .dout(n380));
  jand g00317(.dina(n212), .dinb(n126), .dout(n381));
  jor  g00318(.dina(n381), .dinb(n380), .dout(n382));
  jand g00319(.dina(n159), .dinb(n153), .dout(n383));
  jand g00320(.dina(n219), .dinb(n80), .dout(n384));
  jor  g00321(.dina(n384), .dinb(n383), .dout(n385));
  jor  g00322(.dina(n385), .dinb(n382), .dout(n386));
  jand g00323(.dina(n181), .dinb(n126), .dout(n387));
  jand g00324(.dina(n183), .dinb(n219), .dout(n388));
  jor  g00325(.dina(n388), .dinb(n387), .dout(n389));
  jand g00326(.dina(n212), .dinb(n149), .dout(n390));
  jand g00327(.dina(n227), .dinb(n96), .dout(n391));
  jor  g00328(.dina(n391), .dinb(n390), .dout(n392));
  jor  g00329(.dina(n392), .dinb(n389), .dout(n393));
  jor  g00330(.dina(n393), .dinb(n386), .dout(n394));
  jand g00331(.dina(n90), .dinb(n80), .dout(n395));
  jand g00332(.dina(n195), .dinb(n96), .dout(n396));
  jor  g00333(.dina(n396), .dinb(n395), .dout(n397));
  jand g00334(.dina(n227), .dinb(n143), .dout(n398));
  jand g00335(.dina(n209), .dinb(n112), .dout(n399));
  jor  g00336(.dina(n399), .dinb(n398), .dout(n400));
  jor  g00337(.dina(n400), .dinb(n397), .dout(n401));
  jand g00338(.dina(n195), .dinb(n219), .dout(n402));
  jand g00339(.dina(n159), .dinb(n143), .dout(n403));
  jor  g00340(.dina(n403), .dinb(n402), .dout(n404));
  jor  g00341(.dina(n404), .dinb(n401), .dout(n405));
  jor  g00342(.dina(n405), .dinb(n394), .dout(n406));
  jor  g00343(.dina(\a[25] ), .dinb(\a[24] ), .dout(n407));
  jor  g00344(.dina(n407), .dinb(n262), .dout(n408));
  jor  g00345(.dina(\a[28] ), .dinb(\a[27] ), .dout(n409));
  jor  g00346(.dina(n106), .dinb(n409), .dout(n410));
  jor  g00347(.dina(n410), .dinb(n408), .dout(n411));
  jnot g00348(.din(n411), .dout(n412));
  jand g00349(.dina(n252), .dinb(n227), .dout(n413));
  jor  g00350(.dina(n413), .dinb(n412), .dout(n414));
  jand g00351(.dina(n146), .dinb(n133), .dout(n415));
  jand g00352(.dina(n183), .dinb(n149), .dout(n416));
  jor  g00353(.dina(n416), .dinb(n415), .dout(n417));
  jor  g00354(.dina(n417), .dinb(n414), .dout(n418));
  jand g00355(.dina(n252), .dinb(n176), .dout(n419));
  jand g00356(.dina(n197), .dinb(n176), .dout(n420));
  jor  g00357(.dina(n420), .dinb(n419), .dout(n421));
  jand g00358(.dina(n166), .dinb(n128), .dout(n422));
  jand g00359(.dina(n227), .dinb(n149), .dout(n423));
  jor  g00360(.dina(n423), .dinb(n422), .dout(n424));
  jor  g00361(.dina(n424), .dinb(n421), .dout(n425));
  jor  g00362(.dina(n425), .dinb(n418), .dout(n426));
  jand g00363(.dina(n183), .dinb(n146), .dout(n427));
  jnot g00364(.din(n427), .dout(n428));
  jand g00365(.dina(n252), .dinb(n86), .dout(n429));
  jnot g00366(.din(n429), .dout(n430));
  jand g00367(.dina(n430), .dinb(n428), .dout(n431));
  jnot g00368(.din(n431), .dout(n432));
  jor  g00369(.dina(n432), .dinb(n426), .dout(n433));
  jor  g00370(.dina(n433), .dinb(n406), .dout(n434));
  jor  g00371(.dina(n434), .dinb(n379), .dout(n435));
  jor  g00372(.dina(n435), .dinb(n347), .dout(n436));
  jor  g00373(.dina(n436), .dinb(n260), .dout(n437));
  jor  g00374(.dina(n437), .dinb(n124), .dout(n438));
  jor  g00375(.dina(n103), .dinb(n261), .dout(n439));
  jor  g00376(.dina(n439), .dinb(n268), .dout(n440));
  jor  g00377(.dina(n409), .dinb(n116), .dout(n441));
  jor  g00378(.dina(n441), .dinb(n408), .dout(n442));
  jand g00379(.dina(n442), .dinb(n440), .dout(n443));
  jor  g00380(.dina(n261), .dinb(n118), .dout(n444));
  jor  g00381(.dina(n444), .dinb(n410), .dout(n445));
  jor  g00382(.dina(n323), .dinb(n261), .dout(n446));
  jor  g00383(.dina(n446), .dinb(n265), .dout(n447));
  jand g00384(.dina(n447), .dinb(n445), .dout(n448));
  jand g00385(.dina(n448), .dinb(n443), .dout(n449));
  jor  g00386(.dina(n444), .dinb(n322), .dout(n450));
  jor  g00387(.dina(n323), .dinb(n102), .dout(n451));
  jor  g00388(.dina(n451), .dinb(n268), .dout(n452));
  jand g00389(.dina(n452), .dinb(n450), .dout(n453));
  jor  g00390(.dina(n451), .dinb(n265), .dout(n454));
  jor  g00391(.dina(n102), .dinb(n118), .dout(n455));
  jor  g00392(.dina(n410), .dinb(n455), .dout(n456));
  jand g00393(.dina(n456), .dinb(n454), .dout(n457));
  jand g00394(.dina(n457), .dinb(n453), .dout(n458));
  jand g00395(.dina(n458), .dinb(n449), .dout(n459));
  jor  g00396(.dina(n321), .dinb(n264), .dout(n460));
  jor  g00397(.dina(n446), .dinb(n460), .dout(n461));
  jor  g00398(.dina(n407), .dinb(n118), .dout(n462));
  jor  g00399(.dina(n265), .dinb(n462), .dout(n463));
  jor  g00400(.dina(n105), .dinb(n116), .dout(n464));
  jor  g00401(.dina(n324), .dinb(n464), .dout(n465));
  jand g00402(.dina(n465), .dinb(n463), .dout(n466));
  jand g00403(.dina(n466), .dinb(n461), .dout(n467));
  jor  g00404(.dina(n407), .dinb(n103), .dout(n468));
  jor  g00405(.dina(n468), .dinb(n107), .dout(n469));
  jor  g00406(.dina(n446), .dinb(n117), .dout(n470));
  jor  g00407(.dina(n267), .dinb(n409), .dout(n471));
  jor  g00408(.dina(n451), .dinb(n471), .dout(n472));
  jand g00409(.dina(n472), .dinb(n470), .dout(n473));
  jand g00410(.dina(n473), .dinb(n469), .dout(n474));
  jand g00411(.dina(n474), .dinb(n467), .dout(n475));
  jand g00412(.dina(n475), .dinb(n459), .dout(n476));
  jand g00413(.dina(n144), .dinb(n140), .dout(n477));
  jor  g00414(.dina(n477), .dinb(n399), .dout(n478));
  jnot g00415(.din(n478), .dout(n479));
  jor  g00416(.dina(n451), .dinb(n464), .dout(n480));
  jor  g00417(.dina(n464), .dinb(n120), .dout(n481));
  jand g00418(.dina(n481), .dinb(n266), .dout(n482));
  jand g00419(.dina(n482), .dinb(n480), .dout(n483));
  jand g00420(.dina(n483), .dinb(n479), .dout(n484));
  jand g00421(.dina(n484), .dinb(n476), .dout(n485));
  jand g00422(.dina(n153), .dinb(n98), .dout(n486));
  jand g00423(.dina(n155), .dinb(n149), .dout(n487));
  jor  g00424(.dina(n487), .dinb(n174), .dout(n488));
  jor  g00425(.dina(n488), .dinb(n486), .dout(n489));
  jnot g00426(.din(n489), .dout(n490));
  jor  g00427(.dina(n267), .dinb(n115), .dout(n491));
  jor  g00428(.dina(n491), .dinb(n446), .dout(n492));
  jor  g00429(.dina(n269), .dinb(n117), .dout(n493));
  jor  g00430(.dina(n106), .dinb(n115), .dout(n494));
  jor  g00431(.dina(n494), .dinb(n408), .dout(n495));
  jand g00432(.dina(n495), .dinb(n493), .dout(n496));
  jand g00433(.dina(n496), .dinb(n492), .dout(n497));
  jand g00434(.dina(n149), .dinb(n112), .dout(n498));
  jnot g00435(.din(n498), .dout(n499));
  jor  g00436(.dina(n321), .dinb(n106), .dout(n500));
  jor  g00437(.dina(n439), .dinb(n500), .dout(n501));
  jor  g00438(.dina(n119), .dinb(n103), .dout(n502));
  jor  g00439(.dina(n500), .dinb(n502), .dout(n503));
  jand g00440(.dina(n503), .dinb(n501), .dout(n504));
  jand g00441(.dina(n504), .dinb(n499), .dout(n505));
  jand g00442(.dina(n505), .dinb(n497), .dout(n506));
  jand g00443(.dina(n506), .dinb(n490), .dout(n507));
  jand g00444(.dina(n507), .dinb(n485), .dout(n508));
  jor  g00445(.dina(n264), .dinb(n115), .dout(n509));
  jor  g00446(.dina(n509), .dinb(n502), .dout(n510));
  jor  g00447(.dina(n444), .dinb(n460), .dout(n511));
  jand g00448(.dina(n511), .dinb(n510), .dout(n512));
  jand g00449(.dina(n252), .dinb(n155), .dout(n513));
  jnot g00450(.din(n513), .dout(n514));
  jor  g00451(.dina(n264), .dinb(n409), .dout(n515));
  jor  g00452(.dina(n269), .dinb(n515), .dout(n516));
  jor  g00453(.dina(n446), .dinb(n322), .dout(n517));
  jand g00454(.dina(n325), .dinb(n517), .dout(n518));
  jand g00455(.dina(n518), .dinb(n516), .dout(n519));
  jand g00456(.dina(n186), .dinb(n112), .dout(n520));
  jnot g00457(.din(n520), .dout(n521));
  jand g00458(.dina(n521), .dinb(n519), .dout(n522));
  jand g00459(.dina(n522), .dinb(n514), .dout(n523));
  jor  g00460(.dina(n354), .dinb(n279), .dout(n524));
  jor  g00461(.dina(n220), .dinb(n91), .dout(n525));
  jor  g00462(.dina(n525), .dinb(n524), .dout(n526));
  jnot g00463(.din(n526), .dout(n527));
  jand g00464(.dina(n527), .dinb(n523), .dout(n528));
  jand g00465(.dina(n528), .dinb(n512), .dout(n529));
  jand g00466(.dina(n529), .dinb(n508), .dout(n530));
  jand g00467(.dina(n155), .dinb(n76), .dout(n531));
  jnot g00468(.din(n531), .dout(n532));
  jand g00469(.dina(n209), .dinb(n181), .dout(n533));
  jnot g00470(.din(n533), .dout(n534));
  jand g00471(.dina(n534), .dinb(n532), .dout(n535));
  jand g00472(.dina(n209), .dinb(n128), .dout(n536));
  jnot g00473(.din(n536), .dout(n537));
  jand g00474(.dina(n537), .dinb(n168), .dout(n538));
  jor  g00475(.dina(n119), .dinb(n262), .dout(n539));
  jor  g00476(.dina(n321), .dinb(n267), .dout(n540));
  jor  g00477(.dina(n540), .dinb(n539), .dout(n541));
  jor  g00478(.dina(n491), .dinb(n263), .dout(n542));
  jand g00479(.dina(n542), .dinb(n541), .dout(n543));
  jand g00480(.dina(n543), .dinb(n538), .dout(n544));
  jand g00481(.dina(n544), .dinb(n535), .dout(n545));
  jand g00482(.dina(n197), .dinb(n98), .dout(n546));
  jnot g00483(.din(n546), .dout(n547));
  jor  g00484(.dina(n269), .dinb(n460), .dout(n548));
  jand g00485(.dina(n548), .dinb(n547), .dout(n549));
  jand g00486(.dina(n549), .dinb(n545), .dout(n550));
  jor  g00487(.dina(n515), .dinb(n455), .dout(n551));
  jand g00488(.dina(n155), .dinb(n90), .dout(n552));
  jnot g00489(.din(n552), .dout(n553));
  jand g00490(.dina(n553), .dinb(n551), .dout(n554));
  jnot g00491(.din(n357), .dout(n555));
  jand g00492(.dina(n153), .dinb(n112), .dout(n556));
  jnot g00493(.din(n556), .dout(n557));
  jand g00494(.dina(n557), .dinb(n555), .dout(n558));
  jand g00495(.dina(n558), .dinb(n554), .dout(n559));
  jnot g00496(.din(n236), .dout(n560));
  jand g00497(.dina(n252), .dinb(n195), .dout(n561));
  jnot g00498(.din(n561), .dout(n562));
  jand g00499(.dina(n562), .dinb(n560), .dout(n563));
  jand g00500(.dina(n563), .dinb(n559), .dout(n564));
  jand g00501(.dina(n564), .dinb(n550), .dout(n565));
  jand g00502(.dina(n169), .dinb(n155), .dout(n566));
  jor  g00503(.dina(n566), .dinb(n129), .dout(n567));
  jor  g00504(.dina(n567), .dinb(n419), .dout(n568));
  jand g00505(.dina(n227), .dinb(n146), .dout(n569));
  jor  g00506(.dina(n569), .dinb(n158), .dout(n570));
  jor  g00507(.dina(n570), .dinb(n213), .dout(n571));
  jor  g00508(.dina(n571), .dinb(n568), .dout(n572));
  jand g00509(.dina(n166), .dinb(n98), .dout(n573));
  jand g00510(.dina(n186), .dinb(n98), .dout(n574));
  jor  g00511(.dina(n574), .dinb(n573), .dout(n575));
  jor  g00512(.dina(n575), .dinb(n205), .dout(n576));
  jand g00513(.dina(n197), .dinb(n159), .dout(n577));
  jor  g00514(.dina(n577), .dinb(n280), .dout(n578));
  jor  g00515(.dina(n578), .dinb(n295), .dout(n579));
  jor  g00516(.dina(n579), .dinb(n576), .dout(n580));
  jor  g00517(.dina(n580), .dinb(n572), .dout(n581));
  jnot g00518(.din(n231), .dout(n582));
  jnot g00519(.din(n402), .dout(n583));
  jand g00520(.dina(n583), .dinb(n582), .dout(n584));
  jand g00521(.dina(n144), .dinb(n76), .dout(n585));
  jnot g00522(.din(n585), .dout(n586));
  jand g00523(.dina(n195), .dinb(n166), .dout(n587));
  jnot g00524(.din(n587), .dout(n588));
  jand g00525(.dina(n588), .dinb(n586), .dout(n589));
  jand g00526(.dina(n589), .dinb(n584), .dout(n590));
  jnot g00527(.din(n590), .dout(n591));
  jor  g00528(.dina(n591), .dinb(n581), .dout(n592));
  jnot g00529(.din(n592), .dout(n593));
  jand g00530(.dina(n209), .dinb(n195), .dout(n594));
  jand g00531(.dina(n252), .dinb(n98), .dout(n595));
  jor  g00532(.dina(n595), .dinb(n334), .dout(n596));
  jor  g00533(.dina(n596), .dinb(n594), .dout(n597));
  jnot g00534(.din(n597), .dout(n598));
  jand g00535(.dina(n186), .dinb(n181), .dout(n599));
  jnot g00536(.din(n599), .dout(n600));
  jand g00537(.dina(n600), .dinb(n320), .dout(n601));
  jand g00538(.dina(n601), .dinb(n598), .dout(n602));
  jand g00539(.dina(n112), .dinb(n219), .dout(n603));
  jand g00540(.dina(n227), .dinb(n219), .dout(n604));
  jor  g00541(.dina(n604), .dinb(n603), .dout(n605));
  jand g00542(.dina(n128), .dinb(n76), .dout(n606));
  jor  g00543(.dina(n606), .dinb(n226), .dout(n607));
  jor  g00544(.dina(n607), .dinb(n605), .dout(n608));
  jand g00545(.dina(n227), .dinb(n126), .dout(n609));
  jor  g00546(.dina(n609), .dinb(n249), .dout(n610));
  jand g00547(.dina(n166), .dinb(n86), .dout(n611));
  jand g00548(.dina(n127), .dinb(n118), .dout(n612));
  jand g00549(.dina(n612), .dinb(n166), .dout(n613));
  jor  g00550(.dina(n613), .dinb(n611), .dout(n614));
  jor  g00551(.dina(n614), .dinb(n610), .dout(n615));
  jor  g00552(.dina(n615), .dinb(n608), .dout(n616));
  jnot g00553(.din(n616), .dout(n617));
  jand g00554(.dina(n617), .dinb(n602), .dout(n618));
  jor  g00555(.dina(n322), .dinb(n439), .dout(n619));
  jand g00556(.dina(n195), .dinb(n140), .dout(n620));
  jnot g00557(.din(n620), .dout(n621));
  jand g00558(.dina(n621), .dinb(n619), .dout(n622));
  jand g00559(.dina(n183), .dinb(n169), .dout(n623));
  jand g00560(.dina(n153), .dinb(n86), .dout(n624));
  jor  g00561(.dina(n624), .dinb(n623), .dout(n625));
  jor  g00562(.dina(n625), .dinb(n306), .dout(n626));
  jnot g00563(.din(n626), .dout(n627));
  jand g00564(.dina(n627), .dinb(n622), .dout(n628));
  jand g00565(.dina(n166), .dinb(n144), .dout(n629));
  jnot g00566(.din(n629), .dout(n630));
  jand g00567(.dina(n183), .dinb(n76), .dout(n631));
  jnot g00568(.din(n631), .dout(n632));
  jand g00569(.dina(n632), .dinb(n630), .dout(n633));
  jand g00570(.dina(n633), .dinb(n628), .dout(n634));
  jand g00571(.dina(n634), .dinb(n618), .dout(n635));
  jand g00572(.dina(n635), .dinb(n593), .dout(n636));
  jand g00573(.dina(n636), .dinb(n565), .dout(n637));
  jnot g00574(.din(n331), .dout(n638));
  jor  g00575(.dina(n265), .dinb(n468), .dout(n639));
  jand g00576(.dina(n140), .dinb(n86), .dout(n640));
  jnot g00577(.din(n640), .dout(n641));
  jand g00578(.dina(n641), .dinb(n639), .dout(n642));
  jand g00579(.dina(n642), .dinb(n349), .dout(n643));
  jand g00580(.dina(n183), .dinb(n126), .dout(n644));
  jnot g00581(.din(n644), .dout(n645));
  jand g00582(.dina(n176), .dinb(n90), .dout(n646));
  jnot g00583(.din(n646), .dout(n647));
  jand g00584(.dina(n647), .dinb(n645), .dout(n648));
  jand g00585(.dina(n143), .dinb(n86), .dout(n649));
  jnot g00586(.din(n649), .dout(n650));
  jand g00587(.dina(n650), .dinb(n108), .dout(n651));
  jor  g00588(.dina(n323), .dinb(n407), .dout(n652));
  jor  g00589(.dina(n652), .dinb(n410), .dout(n653));
  jor  g00590(.dina(n462), .dinb(n540), .dout(n654));
  jand g00591(.dina(n654), .dinb(n653), .dout(n655));
  jand g00592(.dina(n655), .dinb(n651), .dout(n656));
  jand g00593(.dina(n656), .dinb(n648), .dout(n657));
  jand g00594(.dina(n657), .dinb(n643), .dout(n658));
  jand g00595(.dina(n658), .dinb(n638), .dout(n659));
  jor  g00596(.dina(n540), .dinb(n455), .dout(n660));
  jand g00597(.dina(n660), .dinb(n411), .dout(n661));
  jnot g00598(.din(n196), .dout(n662));
  jand g00599(.dina(n212), .dinb(n96), .dout(n663));
  jnot g00600(.din(n663), .dout(n664));
  jand g00601(.dina(n664), .dinb(n662), .dout(n665));
  jand g00602(.dina(n665), .dinb(n661), .dout(n666));
  jand g00603(.dina(n140), .dinb(n176), .dout(n667));
  jnot g00604(.din(n667), .dout(n668));
  jand g00605(.dina(n169), .dinb(n98), .dout(n669));
  jnot g00606(.din(n669), .dout(n670));
  jand g00607(.dina(n212), .dinb(n186), .dout(n671));
  jnot g00608(.din(n671), .dout(n672));
  jand g00609(.dina(n672), .dinb(n670), .dout(n673));
  jand g00610(.dina(n673), .dinb(n668), .dout(n674));
  jand g00611(.dina(n674), .dinb(n666), .dout(n675));
  jnot g00612(.din(n206), .dout(n676));
  jand g00613(.dina(n144), .dinb(n126), .dout(n677));
  jnot g00614(.din(n677), .dout(n678));
  jand g00615(.dina(n183), .dinb(n166), .dout(n679));
  jnot g00616(.din(n679), .dout(n680));
  jand g00617(.dina(n680), .dinb(n678), .dout(n681));
  jand g00618(.dina(n681), .dinb(n676), .dout(n682));
  jnot g00619(.din(n253), .dout(n683));
  jand g00620(.dina(n149), .dinb(n133), .dout(n684));
  jnot g00621(.din(n684), .dout(n685));
  jand g00622(.dina(n685), .dinb(n683), .dout(n686));
  jand g00623(.dina(n686), .dinb(n100), .dout(n687));
  jand g00624(.dina(n687), .dinb(n682), .dout(n688));
  jand g00625(.dina(n688), .dinb(n675), .dout(n689));
  jand g00626(.dina(n209), .dinb(n183), .dout(n690));
  jnot g00627(.din(n690), .dout(n691));
  jand g00628(.dina(n209), .dinb(n139), .dout(n692));
  jnot g00629(.din(n692), .dout(n693));
  jand g00630(.dina(n693), .dinb(n691), .dout(n694));
  jnot g00631(.din(n375), .dout(n695));
  jor  g00632(.dina(n451), .dinb(n322), .dout(n696));
  jand g00633(.dina(n696), .dinb(n695), .dout(n697));
  jand g00634(.dina(n697), .dinb(n694), .dout(n698));
  jor  g00635(.dina(n468), .dinb(n117), .dout(n699));
  jor  g00636(.dina(n408), .dinb(n107), .dout(n700));
  jand g00637(.dina(n700), .dinb(n699), .dout(n701));
  jand g00638(.dina(n209), .dinb(n159), .dout(n702));
  jnot g00639(.din(n702), .dout(n703));
  jand g00640(.dina(n703), .dinb(n171), .dout(n704));
  jand g00641(.dina(n704), .dinb(n701), .dout(n705));
  jand g00642(.dina(n705), .dinb(n698), .dout(n706));
  jand g00643(.dina(n98), .dinb(n90), .dout(n707));
  jand g00644(.dina(n181), .dinb(n143), .dout(n708));
  jor  g00645(.dina(n708), .dinb(n361), .dout(n709));
  jor  g00646(.dina(n709), .dinb(n707), .dout(n710));
  jor  g00647(.dina(n710), .dinb(n150), .dout(n711));
  jnot g00648(.din(n711), .dout(n712));
  jnot g00649(.din(n355), .dout(n713));
  jor  g00650(.dina(n441), .dinb(n324), .dout(n714));
  jand g00651(.dina(n714), .dinb(n713), .dout(n715));
  jor  g00652(.dina(n494), .dinb(n539), .dout(n716));
  jand g00653(.dina(n146), .dinb(n86), .dout(n717));
  jnot g00654(.din(n717), .dout(n718));
  jand g00655(.dina(n718), .dinb(n716), .dout(n719));
  jand g00656(.dina(n719), .dinb(n715), .dout(n720));
  jand g00657(.dina(n720), .dinb(n712), .dout(n721));
  jand g00658(.dina(n721), .dinb(n706), .dout(n722));
  jand g00659(.dina(n722), .dinb(n689), .dout(n723));
  jand g00660(.dina(n723), .dinb(n659), .dout(n724));
  jand g00661(.dina(n724), .dinb(n637), .dout(n725));
  jand g00662(.dina(n725), .dinb(n530), .dout(n726));
  jxor g00663(.dina(n726), .dinb(n438), .dout(n727));
  jnot g00664(.din(n727), .dout(n728));
  jand g00665(.dina(n728), .dinb(n71), .dout(n729));
  jxor g00666(.dina(\a[25] ), .dinb(\a[24] ), .dout(n730));
  jand g00667(.dina(n730), .dinb(n66), .dout(n731));
  jand g00668(.dina(n731), .dinb(n438), .dout(n732));
  jand g00669(.dina(n144), .dinb(n96), .dout(n733));
  jand g00670(.dina(n252), .dinb(n128), .dout(n734));
  jor  g00671(.dina(n734), .dinb(n733), .dout(n735));
  jand g00672(.dina(n212), .dinb(n153), .dout(n736));
  jand g00673(.dina(n195), .dinb(n186), .dout(n737));
  jor  g00674(.dina(n737), .dinb(n736), .dout(n738));
  jor  g00675(.dina(n738), .dinb(n735), .dout(n739));
  jand g00676(.dina(n153), .dinb(n80), .dout(n740));
  jor  g00677(.dina(n740), .dinb(n228), .dout(n741));
  jor  g00678(.dina(n741), .dinb(n392), .dout(n742));
  jor  g00679(.dina(n742), .dinb(n739), .dout(n743));
  jand g00680(.dina(n195), .dinb(n126), .dout(n744));
  jor  g00681(.dina(n281), .dinb(n250), .dout(n745));
  jor  g00682(.dina(n745), .dinb(n744), .dout(n746));
  jand g00683(.dina(n227), .dinb(n209), .dout(n747));
  jor  g00684(.dina(n747), .dinb(n301), .dout(n748));
  jor  g00685(.dina(n748), .dinb(n341), .dout(n749));
  jor  g00686(.dina(n749), .dinb(n746), .dout(n750));
  jor  g00687(.dina(n750), .dinb(n743), .dout(n751));
  jand g00688(.dina(n186), .dinb(n86), .dout(n752));
  jor  g00689(.dina(n374), .dinb(n752), .dout(n753));
  jor  g00690(.dina(n753), .dinb(n335), .dout(n754));
  jor  g00691(.dina(n754), .dinb(n478), .dout(n755));
  jor  g00692(.dina(n755), .dinb(n751), .dout(n756));
  jand g00693(.dina(n146), .dinb(n128), .dout(n757));
  jor  g00694(.dina(n757), .dinb(n152), .dout(n758));
  jor  g00695(.dina(n758), .dinb(n309), .dout(n759));
  jand g00696(.dina(n143), .dinb(n112), .dout(n760));
  jor  g00697(.dina(n760), .dinb(n145), .dout(n761));
  jor  g00698(.dina(n761), .dinb(n498), .dout(n762));
  jor  g00699(.dina(n762), .dinb(n759), .dout(n763));
  jor  g00700(.dina(n763), .dinb(n489), .dout(n764));
  jor  g00701(.dina(n764), .dinb(n756), .dout(n765));
  jand g00702(.dina(n139), .dinb(n90), .dout(n766));
  jand g00703(.dina(n181), .dinb(n149), .dout(n767));
  jor  g00704(.dina(n767), .dinb(n234), .dout(n768));
  jor  g00705(.dina(n768), .dinb(n766), .dout(n769));
  jor  g00706(.dina(n520), .dinb(n769), .dout(n770));
  jor  g00707(.dina(n770), .dinb(n513), .dout(n771));
  jor  g00708(.dina(n526), .dinb(n771), .dout(n772));
  jor  g00709(.dina(n772), .dinb(n382), .dout(n773));
  jor  g00710(.dina(n773), .dinb(n765), .dout(n774));
  jnot g00711(.din(n565), .dout(n775));
  jnot g00712(.din(n601), .dout(n776));
  jor  g00713(.dina(n776), .dinb(n597), .dout(n777));
  jor  g00714(.dina(n616), .dinb(n777), .dout(n778));
  jnot g00715(.din(n622), .dout(n779));
  jor  g00716(.dina(n626), .dinb(n779), .dout(n780));
  jnot g00717(.din(n633), .dout(n781));
  jor  g00718(.dina(n781), .dinb(n780), .dout(n782));
  jor  g00719(.dina(n782), .dinb(n778), .dout(n783));
  jor  g00720(.dina(n783), .dinb(n592), .dout(n784));
  jor  g00721(.dina(n784), .dinb(n775), .dout(n785));
  jnot g00722(.din(n659), .dout(n786));
  jnot g00723(.din(n689), .dout(n787));
  jnot g00724(.din(n706), .dout(n788));
  jnot g00725(.din(n720), .dout(n789));
  jor  g00726(.dina(n789), .dinb(n711), .dout(n790));
  jor  g00727(.dina(n790), .dinb(n788), .dout(n791));
  jor  g00728(.dina(n791), .dinb(n787), .dout(n792));
  jor  g00729(.dina(n792), .dinb(n786), .dout(n793));
  jor  g00730(.dina(n793), .dinb(n785), .dout(n794));
  jor  g00731(.dina(n794), .dinb(n774), .dout(n795));
  jand g00732(.dina(n69), .dinb(n67), .dout(n796));
  jand g00733(.dina(n796), .dinb(n795), .dout(n797));
  jor  g00734(.dina(n797), .dinb(n732), .dout(n798));
  jor  g00735(.dina(n798), .dinb(n729), .dout(n799));
  jand g00736(.dina(n438), .dinb(n67), .dout(n800));
  jnot g00737(.din(n800), .dout(n801));
  jor  g00738(.dina(n801), .dinb(n77), .dout(n802));
  jxor g00739(.dina(n802), .dinb(n799), .dout(n803));
  jxor g00740(.dina(\a[21] ), .dinb(\a[20] ), .dout(n804));
  jxor g00741(.dina(\a[23] ), .dinb(\a[22] ), .dout(n805));
  jand g00742(.dina(n805), .dinb(n804), .dout(n806));
  jnot g00743(.din(n806), .dout(n807));
  jor  g00744(.dina(n265), .dinb(n439), .dout(n808));
  jand g00745(.dina(n521), .dinb(n808), .dout(n809));
  jand g00746(.dina(n809), .dinb(n619), .dout(n810));
  jnot g00747(.din(n194), .dout(n811));
  jand g00748(.dina(n456), .dinb(n542), .dout(n812));
  jand g00749(.dina(n812), .dinb(n811), .dout(n813));
  jand g00750(.dina(n813), .dinb(n810), .dout(n814));
  jand g00751(.dina(n814), .dinb(n704), .dout(n815));
  jand g00752(.dina(n547), .dinb(n499), .dout(n816));
  jand g00753(.dina(n816), .dinb(n562), .dout(n817));
  jor  g00754(.dina(n491), .dinb(n120), .dout(n818));
  jand g00755(.dina(n818), .dinb(n560), .dout(n819));
  jand g00756(.dina(n819), .dinb(n817), .dout(n820));
  jand g00757(.dina(n820), .dinb(n554), .dout(n821));
  jand g00758(.dina(n821), .dinb(n815), .dout(n822));
  jnot g00759(.din(n822), .dout(n823));
  jnot g00760(.din(n603), .dout(n824));
  jand g00761(.dina(n133), .dinb(n96), .dout(n825));
  jnot g00762(.din(n825), .dout(n826));
  jand g00763(.dina(n826), .dinb(n824), .dout(n827));
  jand g00764(.dina(n827), .dinb(n639), .dout(n828));
  jnot g00765(.din(n307), .dout(n829));
  jand g00766(.dina(n411), .dinb(n829), .dout(n830));
  jor  g00767(.dina(n451), .dinb(n491), .dout(n831));
  jand g00768(.dina(n197), .dinb(n112), .dout(n832));
  jnot g00769(.din(n832), .dout(n833));
  jand g00770(.dina(n833), .dinb(n831), .dout(n834));
  jand g00771(.dina(n834), .dinb(n830), .dout(n835));
  jand g00772(.dina(n835), .dinb(n828), .dout(n836));
  jnot g00773(.din(n836), .dout(n837));
  jor  g00774(.dina(n460), .dinb(n263), .dout(n838));
  jand g00775(.dina(n514), .dinb(n838), .dout(n839));
  jnot g00776(.din(n839), .dout(n840));
  jand g00777(.dina(n169), .dinb(n86), .dout(n841));
  jor  g00778(.dina(n841), .dinb(n574), .dout(n842));
  jor  g00779(.dina(n540), .dinb(n408), .dout(n843));
  jand g00780(.dina(n472), .dinb(n843), .dout(n844));
  jnot g00781(.din(n844), .dout(n845));
  jor  g00782(.dina(n845), .dinb(n842), .dout(n846));
  jand g00783(.dina(n126), .dinb(n80), .dout(n847));
  jnot g00784(.din(n847), .dout(n848));
  jand g00785(.dina(n848), .dinb(n442), .dout(n849));
  jnot g00786(.din(n849), .dout(n850));
  jor  g00787(.dina(n850), .dinb(n846), .dout(n851));
  jor  g00788(.dina(n851), .dinb(n840), .dout(n852));
  jor  g00789(.dina(n852), .dinb(n837), .dout(n853));
  jand g00790(.dina(n197), .dinb(n80), .dout(n854));
  jor  g00791(.dina(n854), .dinb(n717), .dout(n855));
  jor  g00792(.dina(n855), .dinb(n348), .dout(n856));
  jand g00793(.dina(n195), .dinb(n90), .dout(n857));
  jor  g00794(.dina(n857), .dinb(n198), .dout(n858));
  jand g00795(.dina(n700), .dinb(n481), .dout(n859));
  jnot g00796(.din(n859), .dout(n860));
  jor  g00797(.dina(n860), .dinb(n858), .dout(n861));
  jor  g00798(.dina(n861), .dinb(n856), .dout(n862));
  jand g00799(.dina(n219), .dinb(n98), .dout(n863));
  jand g00800(.dina(n197), .dinb(n181), .dout(n864));
  jor  g00801(.dina(n864), .dinb(n383), .dout(n865));
  jor  g00802(.dina(n865), .dinb(n310), .dout(n866));
  jor  g00803(.dina(n866), .dinb(n863), .dout(n867));
  jor  g00804(.dina(n867), .dinb(n862), .dout(n868));
  jnot g00805(.din(n606), .dout(n869));
  jand g00806(.dina(n632), .dinb(n869), .dout(n870));
  jor  g00807(.dina(n500), .dinb(n539), .dout(n871));
  jand g00808(.dina(n133), .dinb(n219), .dout(n872));
  jnot g00809(.din(n872), .dout(n873));
  jand g00810(.dina(n873), .dinb(n871), .dout(n874));
  jand g00811(.dina(n874), .dinb(n870), .dout(n875));
  jnot g00812(.din(n875), .dout(n876));
  jor  g00813(.dina(n876), .dinb(n868), .dout(n877));
  jor  g00814(.dina(n877), .dinb(n853), .dout(n878));
  jor  g00815(.dina(n878), .dinb(n823), .dout(n879));
  jnot g00816(.din(n150), .dout(n880));
  jnot g00817(.din(n577), .dout(n881));
  jand g00818(.dina(n881), .dinb(n880), .dout(n882));
  jnot g00819(.din(n882), .dout(n883));
  jnot g00820(.din(n486), .dout(n884));
  jand g00821(.dina(n144), .dinb(n219), .dout(n885));
  jnot g00822(.din(n885), .dout(n886));
  jand g00823(.dina(n886), .dinb(n884), .dout(n887));
  jnot g00824(.din(n887), .dout(n888));
  jor  g00825(.dina(n609), .dinb(n187), .dout(n889));
  jand g00826(.dina(n227), .dinb(n166), .dout(n890));
  jor  g00827(.dina(n890), .dinb(n361), .dout(n891));
  jor  g00828(.dina(n891), .dinb(n889), .dout(n892));
  jnot g00829(.din(n373), .dout(n893));
  jand g00830(.dina(n149), .dinb(n128), .dout(n894));
  jnot g00831(.din(n894), .dout(n895));
  jand g00832(.dina(n895), .dinb(n893), .dout(n896));
  jnot g00833(.din(n896), .dout(n897));
  jor  g00834(.dina(n897), .dinb(n892), .dout(n898));
  jand g00835(.dina(n638), .dinb(n517), .dout(n899));
  jor  g00836(.dina(n471), .dinb(n263), .dout(n900));
  jor  g00837(.dina(n471), .dinb(n120), .dout(n901));
  jand g00838(.dina(n901), .dinb(n900), .dout(n902));
  jand g00839(.dina(n902), .dinb(n445), .dout(n903));
  jand g00840(.dina(n903), .dinb(n899), .dout(n904));
  jnot g00841(.din(n904), .dout(n905));
  jor  g00842(.dina(n905), .dinb(n898), .dout(n906));
  jor  g00843(.dina(n509), .dinb(n269), .dout(n907));
  jnot g00844(.din(n707), .dout(n908));
  jand g00845(.dina(n908), .dinb(n465), .dout(n909));
  jand g00846(.dina(n909), .dinb(n907), .dout(n910));
  jnot g00847(.din(n910), .dout(n911));
  jor  g00848(.dina(n911), .dinb(n906), .dout(n912));
  jor  g00849(.dina(n912), .dinb(n888), .dout(n913));
  jor  g00850(.dina(n913), .dinb(n883), .dout(n914));
  jor  g00851(.dina(n914), .dinb(n879), .dout(n915));
  jnot g00852(.din(n332), .dout(n916));
  jor  g00853(.dina(n468), .dinb(n540), .dout(n917));
  jand g00854(.dina(n917), .dinb(n916), .dout(n918));
  jand g00855(.dina(n918), .dinb(n696), .dout(n919));
  jnot g00856(.din(n220), .dout(n920));
  jor  g00857(.dina(n322), .dinb(n455), .dout(n921));
  jand g00858(.dina(n921), .dinb(n480), .dout(n922));
  jand g00859(.dina(n922), .dinb(n920), .dout(n923));
  jand g00860(.dina(n923), .dinb(n919), .dout(n924));
  jor  g00861(.dina(n265), .dinb(n539), .dout(n925));
  jand g00862(.dina(n925), .dinb(n479), .dout(n926));
  jand g00863(.dina(n691), .dinb(n470), .dout(n927));
  jand g00864(.dina(n927), .dinb(n100), .dout(n928));
  jor  g00865(.dina(n539), .dinb(n515), .dout(n929));
  jand g00866(.dina(n112), .dinb(n90), .dout(n930));
  jnot g00867(.din(n930), .dout(n931));
  jand g00868(.dina(n931), .dinb(n929), .dout(n932));
  jnot g00869(.din(n249), .dout(n933));
  jand g00870(.dina(n503), .dinb(n933), .dout(n934));
  jand g00871(.dina(n934), .dinb(n932), .dout(n935));
  jand g00872(.dina(n935), .dinb(n928), .dout(n936));
  jand g00873(.dina(n936), .dinb(n926), .dout(n937));
  jand g00874(.dina(n937), .dinb(n924), .dout(n938));
  jnot g00875(.din(n938), .dout(n939));
  jand g00876(.dina(n159), .dinb(n146), .dout(n940));
  jand g00877(.dina(n212), .dinb(n143), .dout(n941));
  jor  g00878(.dina(n941), .dinb(n556), .dout(n942));
  jor  g00879(.dina(n942), .dinb(n288), .dout(n943));
  jor  g00880(.dina(n943), .dinb(n940), .dout(n944));
  jor  g00881(.dina(n944), .dinb(n536), .dout(n945));
  jor  g00882(.dina(n604), .dinb(n131), .dout(n946));
  jor  g00883(.dina(n946), .dinb(n566), .dout(n947));
  jor  g00884(.dina(n107), .dinb(n455), .dout(n948));
  jand g00885(.dina(n166), .dinb(n159), .dout(n949));
  jnot g00886(.din(n949), .dout(n950));
  jand g00887(.dina(n950), .dinb(n948), .dout(n951));
  jnot g00888(.din(n951), .dout(n952));
  jor  g00889(.dina(n952), .dinb(n947), .dout(n953));
  jor  g00890(.dina(n540), .dinb(n269), .dout(n954));
  jand g00891(.dina(n660), .dinb(n954), .dout(n955));
  jand g00892(.dina(n955), .dinb(n641), .dout(n956));
  jnot g00893(.din(n956), .dout(n957));
  jor  g00894(.dina(n957), .dinb(n953), .dout(n958));
  jor  g00895(.dina(n958), .dinb(n945), .dout(n959));
  jand g00896(.dina(n166), .dinb(n155), .dout(n960));
  jor  g00897(.dina(n960), .dinb(n573), .dout(n961));
  jor  g00898(.dina(n961), .dinb(n230), .dout(n962));
  jor  g00899(.dina(n962), .dinb(n113), .dout(n963));
  jor  g00900(.dina(n446), .dinb(n268), .dout(n964));
  jnot g00901(.din(n708), .dout(n965));
  jand g00902(.dina(n965), .dinb(n964), .dout(n966));
  jnot g00903(.din(n966), .dout(n967));
  jand g00904(.dina(n128), .dinb(n90), .dout(n968));
  jor  g00905(.dina(n968), .dinb(n294), .dout(n969));
  jor  g00906(.dina(n585), .dinb(n336), .dout(n970));
  jor  g00907(.dina(n970), .dinb(n969), .dout(n971));
  jor  g00908(.dina(n971), .dinb(n967), .dout(n972));
  jor  g00909(.dina(n972), .dinb(n963), .dout(n973));
  jor  g00910(.dina(n973), .dinb(n375), .dout(n974));
  jor  g00911(.dina(n974), .dinb(n959), .dout(n975));
  jor  g00912(.dina(n975), .dinb(n939), .dout(n976));
  jand g00913(.dina(n143), .dinb(n176), .dout(n977));
  jnot g00914(.din(n977), .dout(n978));
  jand g00915(.dina(n978), .dinb(n440), .dout(n979));
  jand g00916(.dina(n126), .dinb(n98), .dout(n980));
  jnot g00917(.din(n980), .dout(n981));
  jand g00918(.dina(n981), .dinb(n328), .dout(n982));
  jor  g00919(.dina(n441), .dinb(n539), .dout(n983));
  jand g00920(.dina(n983), .dinb(n461), .dout(n984));
  jand g00921(.dina(n984), .dinb(n982), .dout(n985));
  jand g00922(.dina(n985), .dinb(n979), .dout(n986));
  jnot g00923(.din(n986), .dout(n987));
  jor  g00924(.dina(n509), .dinb(n408), .dout(n988));
  jand g00925(.dina(n988), .dinb(n92), .dout(n989));
  jnot g00926(.din(n989), .dout(n990));
  jnot g00927(.din(n306), .dout(n991));
  jand g00928(.dina(n212), .dinb(n146), .dout(n992));
  jnot g00929(.din(n992), .dout(n993));
  jand g00930(.dina(n993), .dinb(n991), .dout(n994));
  jnot g00931(.din(n994), .dout(n995));
  jand g00932(.dina(n195), .dinb(n143), .dout(n996));
  jor  g00933(.dina(n996), .dinb(n279), .dout(n997));
  jand g00934(.dina(n195), .dinb(n169), .dout(n998));
  jor  g00935(.dina(n998), .dinb(n997), .dout(n999));
  jand g00936(.dina(n139), .dinb(n96), .dout(n1000));
  jor  g00937(.dina(n1000), .dinb(n188), .dout(n1001));
  jor  g00938(.dina(n1001), .dinb(n185), .dout(n1002));
  jor  g00939(.dina(n1002), .dinb(n999), .dout(n1003));
  jor  g00940(.dina(n1003), .dinb(n995), .dout(n1004));
  jnot g00941(.din(n594), .dout(n1005));
  jand g00942(.dina(n630), .dinb(n1005), .dout(n1006));
  jnot g00943(.din(n1006), .dout(n1007));
  jand g00944(.dina(n144), .dinb(n90), .dout(n1008));
  jor  g00945(.dina(n1008), .dinb(n362), .dout(n1009));
  jor  g00946(.dina(n1009), .dinb(n757), .dout(n1010));
  jor  g00947(.dina(n671), .dinb(n302), .dout(n1011));
  jor  g00948(.dina(n1011), .dinb(n1010), .dout(n1012));
  jor  g00949(.dina(n1012), .dinb(n1007), .dout(n1013));
  jor  g00950(.dina(n1013), .dinb(n1004), .dout(n1014));
  jand g00951(.dina(n146), .dinb(n80), .dout(n1015));
  jnot g00952(.din(n1015), .dout(n1016));
  jand g00953(.dina(n1016), .dinb(n493), .dout(n1017));
  jand g00954(.dina(n1017), .dinb(n492), .dout(n1018));
  jnot g00955(.din(n1018), .dout(n1019));
  jor  g00956(.dina(n1019), .dinb(n1014), .dout(n1020));
  jor  g00957(.dina(n1020), .dinb(n990), .dout(n1021));
  jor  g00958(.dina(n1021), .dinb(n987), .dout(n1022));
  jor  g00959(.dina(n1022), .dinb(n976), .dout(n1023));
  jor  g00960(.dina(n1023), .dinb(n915), .dout(n1024));
  jand g00961(.dina(n209), .dinb(n133), .dout(n1025));
  jor  g00962(.dina(n1025), .dinb(n872), .dout(n1026));
  jor  g00963(.dina(n244), .dinb(n202), .dout(n1027));
  jor  g00964(.dina(n1027), .dinb(n1026), .dout(n1028));
  jor  g00965(.dina(n1028), .dinb(n331), .dout(n1029));
  jor  g00966(.dina(n1029), .dinb(n960), .dout(n1030));
  jor  g00967(.dina(n603), .dinb(n287), .dout(n1031));
  jor  g00968(.dina(n1031), .dinb(n415), .dout(n1032));
  jor  g00969(.dina(n1032), .dinb(n667), .dout(n1033));
  jor  g00970(.dina(n1033), .dinb(n552), .dout(n1034));
  jor  g00971(.dina(n1034), .dinb(n1030), .dout(n1035));
  jor  g00972(.dina(n468), .dinb(n410), .dout(n1036));
  jnot g00973(.din(n968), .dout(n1037));
  jand g00974(.dina(n1037), .dinb(n1036), .dout(n1038));
  jnot g00975(.din(n1038), .dout(n1039));
  jnot g00976(.din(n205), .dout(n1040));
  jand g00977(.dina(n169), .dinb(n112), .dout(n1041));
  jnot g00978(.din(n1041), .dout(n1042));
  jand g00979(.dina(n1042), .dinb(n1040), .dout(n1043));
  jnot g00980(.din(n1043), .dout(n1044));
  jor  g00981(.dina(n1015), .dinb(n158), .dout(n1045));
  jor  g00982(.dina(n894), .dinb(n170), .dout(n1046));
  jor  g00983(.dina(n1046), .dinb(n1045), .dout(n1047));
  jor  g00984(.dina(n1047), .dinb(n1044), .dout(n1048));
  jor  g00985(.dina(n1048), .dinb(n113), .dout(n1049));
  jor  g00986(.dina(n1049), .dinb(n1039), .dout(n1050));
  jor  g00987(.dina(n1050), .dinb(n1035), .dout(n1051));
  jand g00988(.dina(n153), .dinb(n133), .dout(n1052));
  jnot g00989(.din(n1052), .dout(n1053));
  jand g00990(.dina(n1053), .dinb(n555), .dout(n1054));
  jand g00991(.dina(n1054), .dinb(n100), .dout(n1055));
  jnot g00992(.din(n1055), .dout(n1056));
  jand g00993(.dina(n212), .dinb(n140), .dout(n1057));
  jor  g00994(.dina(n629), .dinb(n236), .dout(n1058));
  jor  g00995(.dina(n1058), .dinb(n1057), .dout(n1059));
  jor  g00996(.dina(n1059), .dinb(n285), .dout(n1060));
  jor  g00997(.dina(n1060), .dinb(n1056), .dout(n1061));
  jnot g00998(.din(n697), .dout(n1062));
  jand g00999(.dina(n155), .dinb(n219), .dout(n1063));
  jand g01000(.dina(n212), .dinb(n219), .dout(n1064));
  jor  g01001(.dina(n1064), .dinb(n182), .dout(n1065));
  jand g01002(.dina(n126), .dinb(n112), .dout(n1066));
  jor  g01003(.dina(n1066), .dinb(n677), .dout(n1067));
  jor  g01004(.dina(n1067), .dinb(n1065), .dout(n1068));
  jor  g01005(.dina(n1068), .dinb(n1063), .dout(n1069));
  jor  g01006(.dina(n1069), .dinb(n1062), .dout(n1070));
  jor  g01007(.dina(n1070), .dinb(n1061), .dout(n1071));
  jand g01008(.dina(n159), .dinb(n140), .dout(n1072));
  jand g01009(.dina(n181), .dinb(n153), .dout(n1073));
  jor  g01010(.dina(n1073), .dinb(n1072), .dout(n1074));
  jor  g01011(.dina(n1074), .dinb(n254), .dout(n1075));
  jand g01012(.dina(n176), .dinb(n76), .dout(n1076));
  jor  g01013(.dina(n217), .dinb(n1076), .dout(n1077));
  jor  g01014(.dina(n1077), .dinb(n587), .dout(n1078));
  jor  g01015(.dina(n1078), .dinb(n1075), .dout(n1079));
  jand g01016(.dina(n128), .dinb(n96), .dout(n1080));
  jor  g01017(.dina(n1080), .dinb(n245), .dout(n1081));
  jand g01018(.dina(n195), .dinb(n146), .dout(n1082));
  jor  g01019(.dina(n1082), .dinb(n184), .dout(n1083));
  jor  g01020(.dina(n1083), .dinb(n1081), .dout(n1084));
  jor  g01021(.dina(n1084), .dinb(n1079), .dout(n1085));
  jor  g01022(.dina(n980), .dinb(n604), .dout(n1086));
  jor  g01023(.dina(n1086), .dinb(n280), .dout(n1087));
  jnot g01024(.din(n213), .dout(n1088));
  jand g01025(.dina(n166), .dinb(n133), .dout(n1089));
  jnot g01026(.din(n1089), .dout(n1090));
  jand g01027(.dina(n1090), .dinb(n1088), .dout(n1091));
  jnot g01028(.din(n1091), .dout(n1092));
  jor  g01029(.dina(n1092), .dinb(n1087), .dout(n1093));
  jor  g01030(.dina(n1093), .dinb(n1085), .dout(n1094));
  jand g01031(.dina(n181), .dinb(n140), .dout(n1095));
  jnot g01032(.din(n1095), .dout(n1096));
  jand g01033(.dina(n212), .dinb(n169), .dout(n1097));
  jnot g01034(.din(n1097), .dout(n1098));
  jand g01035(.dina(n1098), .dinb(n582), .dout(n1099));
  jand g01036(.dina(n1099), .dinb(n1096), .dout(n1100));
  jand g01037(.dina(n1100), .dinb(n352), .dout(n1101));
  jnot g01038(.din(n1101), .dout(n1102));
  jor  g01039(.dina(n1102), .dinb(n1094), .dout(n1103));
  jor  g01040(.dina(n1103), .dinb(n1071), .dout(n1104));
  jor  g01041(.dina(n1104), .dinb(n1051), .dout(n1105));
  jand g01042(.dina(n183), .dinb(n153), .dout(n1106));
  jnot g01043(.din(n1106), .dout(n1107));
  jand g01044(.dina(n1107), .dinb(n833), .dout(n1108));
  jnot g01045(.din(n1108), .dout(n1109));
  jand g01046(.dina(n140), .dinb(n80), .dout(n1110));
  jor  g01047(.dina(n1110), .dinb(n141), .dout(n1111));
  jor  g01048(.dina(n1111), .dinb(n275), .dout(n1112));
  jand g01049(.dina(n149), .dinb(n80), .dout(n1113));
  jor  g01050(.dina(n1113), .dinb(n208), .dout(n1114));
  jand g01051(.dina(n186), .dinb(n133), .dout(n1115));
  jand g01052(.dina(n227), .dinb(n153), .dout(n1116));
  jor  g01053(.dina(n1116), .dinb(n1115), .dout(n1117));
  jor  g01054(.dina(n1117), .dinb(n1114), .dout(n1118));
  jor  g01055(.dina(n1118), .dinb(n1112), .dout(n1119));
  jor  g01056(.dina(n1119), .dinb(n1109), .dout(n1120));
  jand g01057(.dina(n227), .dinb(n140), .dout(n1121));
  jand g01058(.dina(n128), .dinb(n219), .dout(n1122));
  jor  g01059(.dina(n1122), .dinb(n147), .dout(n1123));
  jor  g01060(.dina(n1123), .dinb(n396), .dout(n1124));
  jor  g01061(.dina(n1124), .dinb(n1121), .dout(n1125));
  jand g01062(.dina(n212), .dinb(n197), .dout(n1126));
  jor  g01063(.dina(n1126), .dinb(n360), .dout(n1127));
  jand g01064(.dina(n169), .dinb(n144), .dout(n1128));
  jor  g01065(.dina(n1128), .dinb(n998), .dout(n1129));
  jor  g01066(.dina(n1129), .dinb(n131), .dout(n1130));
  jor  g01067(.dina(n1130), .dinb(n1127), .dout(n1131));
  jor  g01068(.dina(n1131), .dinb(n1125), .dout(n1132));
  jor  g01069(.dina(n1132), .dinb(n1120), .dout(n1133));
  jand g01070(.dina(n186), .dinb(n80), .dout(n1134));
  jor  g01071(.dina(n1134), .dinb(n940), .dout(n1135));
  jor  g01072(.dina(n1135), .dinb(n160), .dout(n1136));
  jor  g01073(.dina(n1136), .dinb(n373), .dout(n1137));
  jor  g01074(.dina(n1137), .dinb(n229), .dout(n1138));
  jor  g01075(.dina(n1000), .dinb(n199), .dout(n1139));
  jor  g01076(.dina(n1139), .dinb(n307), .dout(n1140));
  jand g01077(.dina(n252), .dinb(n133), .dout(n1141));
  jor  g01078(.dina(n1141), .dinb(n221), .dout(n1142));
  jand g01079(.dina(n197), .dinb(n128), .dout(n1143));
  jor  g01080(.dina(n420), .dinb(n273), .dout(n1144));
  jor  g01081(.dina(n1144), .dinb(n1143), .dout(n1145));
  jor  g01082(.dina(n1145), .dinb(n1142), .dout(n1146));
  jor  g01083(.dina(n1146), .dinb(n1140), .dout(n1147));
  jor  g01084(.dina(n1147), .dinb(n1138), .dout(n1148));
  jor  g01085(.dina(n996), .dinb(n81), .dout(n1149));
  jand g01086(.dina(n252), .dinb(n183), .dout(n1150));
  jor  g01087(.dina(n1150), .dinb(n863), .dout(n1151));
  jor  g01088(.dina(n1151), .dinb(n302), .dout(n1152));
  jor  g01089(.dina(n1152), .dinb(n1149), .dout(n1153));
  jor  g01090(.dina(n1153), .dinb(n336), .dout(n1154));
  jor  g01091(.dina(n1154), .dinb(n1148), .dout(n1155));
  jor  g01092(.dina(n1155), .dinb(n1133), .dout(n1156));
  jor  g01093(.dina(n1156), .dinb(n774), .dout(n1157));
  jand g01094(.dina(n133), .dinb(n126), .dout(n1158));
  jnot g01095(.din(n1158), .dout(n1159));
  jnot g01096(.din(n189), .dout(n1160));
  jand g01097(.dina(n209), .dinb(n80), .dout(n1161));
  jnot g01098(.din(n1161), .dout(n1162));
  jand g01099(.dina(n1162), .dinb(n641), .dout(n1163));
  jand g01100(.dina(n1163), .dinb(n1160), .dout(n1164));
  jand g01101(.dina(n1164), .dinb(n1159), .dout(n1165));
  jand g01102(.dina(n252), .dinb(n112), .dout(n1166));
  jnot g01103(.din(n1166), .dout(n1167));
  jand g01104(.dina(n1167), .dinb(n993), .dout(n1168));
  jand g01105(.dina(n430), .dinb(n683), .dout(n1169));
  jand g01106(.dina(n1169), .dinb(n1168), .dout(n1170));
  jand g01107(.dina(n1170), .dinb(n1165), .dout(n1171));
  jand g01108(.dina(n1171), .dinb(n694), .dout(n1172));
  jnot g01109(.din(n1172), .dout(n1173));
  jor  g01110(.dina(n1173), .dinb(n1157), .dout(n1174));
  jor  g01111(.dina(n1174), .dinb(n1105), .dout(n1175));
  jand g01112(.dina(n1175), .dinb(n1024), .dout(n1176));
  jnot g01113(.din(n1176), .dout(n1177));
  jnot g01114(.din(n1035), .dout(n1178));
  jnot g01115(.din(n1047), .dout(n1179));
  jand g01116(.dina(n1179), .dinb(n1043), .dout(n1180));
  jand g01117(.dina(n1180), .dinb(n114), .dout(n1181));
  jand g01118(.dina(n1181), .dinb(n1038), .dout(n1182));
  jand g01119(.dina(n1182), .dinb(n1178), .dout(n1183));
  jnot g01120(.din(n1060), .dout(n1184));
  jand g01121(.dina(n1184), .dinb(n1055), .dout(n1185));
  jnot g01122(.din(n1070), .dout(n1186));
  jand g01123(.dina(n1186), .dinb(n1185), .dout(n1187));
  jnot g01124(.din(n254), .dout(n1188));
  jor  g01125(.dina(n324), .dinb(n410), .dout(n1189));
  jand g01126(.dina(n1189), .dinb(n917), .dout(n1190));
  jand g01127(.dina(n1190), .dinb(n1188), .dout(n1191));
  jand g01128(.dina(n871), .dinb(n121), .dout(n1192));
  jand g01129(.dina(n1192), .dinb(n588), .dout(n1193));
  jand g01130(.dina(n1193), .dinb(n1191), .dout(n1194));
  jnot g01131(.din(n1084), .dout(n1195));
  jand g01132(.dina(n1195), .dinb(n1194), .dout(n1196));
  jnot g01133(.din(n1087), .dout(n1197));
  jand g01134(.dina(n1091), .dinb(n1197), .dout(n1198));
  jand g01135(.dina(n1198), .dinb(n1196), .dout(n1199));
  jand g01136(.dina(n1101), .dinb(n1199), .dout(n1200));
  jand g01137(.dina(n1200), .dinb(n1187), .dout(n1201));
  jand g01138(.dina(n1201), .dinb(n1183), .dout(n1202));
  jor  g01139(.dina(n441), .dinb(n269), .dout(n1203));
  jand g01140(.dina(n955), .dinb(n1203), .dout(n1204));
  jor  g01141(.dina(n491), .dinb(n652), .dout(n1205));
  jand g01142(.dina(n921), .dinb(n1205), .dout(n1206));
  jor  g01143(.dina(n451), .dinb(n410), .dout(n1207));
  jand g01144(.dina(n1207), .dinb(n925), .dout(n1208));
  jand g01145(.dina(n1208), .dinb(n1206), .dout(n1209));
  jand g01146(.dina(n1209), .dinb(n1204), .dout(n1210));
  jand g01147(.dina(n1210), .dinb(n1108), .dout(n1211));
  jnot g01148(.din(n1121), .dout(n1212));
  jor  g01149(.dina(n494), .dinb(n269), .dout(n1213));
  jand g01150(.dina(n700), .dinb(n1213), .dout(n1214));
  jand g01151(.dina(n1214), .dinb(n964), .dout(n1215));
  jand g01152(.dina(n1215), .dinb(n1212), .dout(n1216));
  jnot g01153(.din(n1127), .dout(n1217));
  jor  g01154(.dina(n446), .dinb(n464), .dout(n1218));
  jor  g01155(.dina(n464), .dinb(n439), .dout(n1219));
  jand g01156(.dina(n1219), .dinb(n1218), .dout(n1220));
  jand g01157(.dina(n1220), .dinb(n132), .dout(n1221));
  jand g01158(.dina(n1221), .dinb(n1217), .dout(n1222));
  jand g01159(.dina(n1222), .dinb(n1216), .dout(n1223));
  jand g01160(.dina(n1223), .dinb(n1211), .dout(n1224));
  jor  g01161(.dina(n652), .dinb(n540), .dout(n1225));
  jor  g01162(.dina(n468), .dinb(n268), .dout(n1226));
  jor  g01163(.dina(n468), .dinb(n494), .dout(n1227));
  jor  g01164(.dina(n265), .dinb(n455), .dout(n1228));
  jand g01165(.dina(n1228), .dinb(n1227), .dout(n1229));
  jand g01166(.dina(n1229), .dinb(n1226), .dout(n1230));
  jand g01167(.dina(n1230), .dinb(n893), .dout(n1231));
  jand g01168(.dina(n1231), .dinb(n1225), .dout(n1232));
  jor  g01169(.dina(n468), .dinb(n322), .dout(n1233));
  jand g01170(.dina(n270), .dinb(n1233), .dout(n1234));
  jand g01171(.dina(n1234), .dinb(n829), .dout(n1235));
  jand g01172(.dina(n983), .dinb(n843), .dout(n1236));
  jor  g01173(.dina(n491), .dinb(n408), .dout(n1237));
  jor  g01174(.dina(n324), .dinb(n107), .dout(n1238));
  jand g01175(.dina(n818), .dinb(n1238), .dout(n1239));
  jand g01176(.dina(n1239), .dinb(n1237), .dout(n1240));
  jand g01177(.dina(n1240), .dinb(n1236), .dout(n1241));
  jand g01178(.dina(n1241), .dinb(n1235), .dout(n1242));
  jand g01179(.dina(n1242), .dinb(n1232), .dout(n1243));
  jnot g01180(.din(n1149), .dout(n1244));
  jor  g01181(.dina(n104), .dinb(n117), .dout(n1245));
  jor  g01182(.dina(n441), .dinb(n462), .dout(n1246));
  jand g01183(.dina(n1246), .dinb(n108), .dout(n1247));
  jand g01184(.dina(n1247), .dinb(n1245), .dout(n1248));
  jand g01185(.dina(n1248), .dinb(n1244), .dout(n1249));
  jand g01186(.dina(n1249), .dinb(n699), .dout(n1250));
  jand g01187(.dina(n1250), .dinb(n1243), .dout(n1251));
  jand g01188(.dina(n1251), .dinb(n1224), .dout(n1252));
  jand g01189(.dina(n1252), .dinb(n530), .dout(n1253));
  jand g01190(.dina(n1172), .dinb(n1253), .dout(n1254));
  jand g01191(.dina(n1254), .dinb(n1202), .dout(n1255));
  jxor g01192(.dina(n1255), .dinb(n1024), .dout(n1256));
  jand g01193(.dina(n1213), .dinb(n501), .dout(n1257));
  jand g01194(.dina(n880), .dinb(n1257), .dout(n1258));
  jand g01195(.dina(n653), .dinb(n493), .dout(n1259));
  jor  g01196(.dina(n652), .dinb(n268), .dout(n1260));
  jand g01197(.dina(n1226), .dinb(n1260), .dout(n1261));
  jand g01198(.dina(n1261), .dinb(n1259), .dout(n1262));
  jand g01199(.dina(n1262), .dinb(n1258), .dout(n1263));
  jand g01200(.dina(n1263), .dinb(n954), .dout(n1264));
  jand g01201(.dina(n1264), .dinb(n137), .dout(n1265));
  jnot g01202(.din(n190), .dout(n1266));
  jand g01203(.dina(n1266), .dinb(n179), .dout(n1267));
  jand g01204(.dina(n1267), .dinb(n172), .dout(n1268));
  jand g01205(.dina(n1268), .dinb(n1265), .dout(n1269));
  jor  g01206(.dina(n491), .dinb(n269), .dout(n1270));
  jand g01207(.dina(n1233), .dinb(n1270), .dout(n1271));
  jand g01208(.dina(n1271), .dinb(n662), .dout(n1272));
  jnot g01209(.din(n202), .dout(n1273));
  jand g01210(.dina(n1273), .dinb(n1272), .dout(n1274));
  jand g01211(.dina(n1274), .dinb(n811), .dout(n1275));
  jnot g01212(.din(n207), .dout(n1276));
  jand g01213(.dina(n900), .dinb(n1205), .dout(n1277));
  jand g01214(.dina(n1088), .dinb(n1277), .dout(n1278));
  jand g01215(.dina(n1278), .dinb(n1276), .dout(n1279));
  jnot g01216(.din(n223), .dout(n1280));
  jand g01217(.dina(n1280), .dinb(n1279), .dout(n1281));
  jand g01218(.dina(n1281), .dinb(n1275), .dout(n1282));
  jnot g01219(.din(n226), .dout(n1283));
  jand g01220(.dina(n1225), .dinb(n454), .dout(n1284));
  jand g01221(.dina(n582), .dinb(n1284), .dout(n1285));
  jand g01222(.dina(n1285), .dinb(n1283), .dout(n1286));
  jand g01223(.dina(n517), .dinb(n1286), .dout(n1287));
  jor  g01224(.dina(n444), .dinb(n509), .dout(n1288));
  jand g01225(.dina(n907), .dinb(n1288), .dout(n1289));
  jand g01226(.dina(n1289), .dinb(n560), .dout(n1290));
  jand g01227(.dina(n654), .dinb(n541), .dout(n1291));
  jor  g01228(.dina(n451), .dinb(n515), .dout(n1292));
  jand g01229(.dina(n1292), .dinb(n901), .dout(n1293));
  jand g01230(.dina(n1293), .dinb(n1291), .dout(n1294));
  jand g01231(.dina(n1294), .dinb(n1290), .dout(n1295));
  jnot g01232(.din(n256), .dout(n1296));
  jand g01233(.dina(n1296), .dinb(n1295), .dout(n1297));
  jand g01234(.dina(n1297), .dinb(n1287), .dout(n1298));
  jand g01235(.dina(n1298), .dinb(n1282), .dout(n1299));
  jand g01236(.dina(n1299), .dinb(n1269), .dout(n1300));
  jand g01237(.dina(n1203), .dinb(n639), .dout(n1301));
  jand g01238(.dina(n1301), .dinb(n1238), .dout(n1302));
  jand g01239(.dina(n1302), .dinb(n271), .dout(n1303));
  jor  g01240(.dina(n494), .dinb(n104), .dout(n1304));
  jor  g01241(.dina(n107), .dinb(n263), .dout(n1305));
  jand g01242(.dina(n465), .dinb(n1305), .dout(n1306));
  jand g01243(.dina(n1306), .dinb(n1304), .dout(n1307));
  jand g01244(.dina(n831), .dinb(n929), .dout(n1308));
  jor  g01245(.dina(n410), .dinb(n439), .dout(n1309));
  jor  g01246(.dina(n500), .dinb(n269), .dout(n1310));
  jand g01247(.dina(n1310), .dinb(n1309), .dout(n1311));
  jand g01248(.dina(n1311), .dinb(n1308), .dout(n1312));
  jand g01249(.dina(n1312), .dinb(n1307), .dout(n1313));
  jand g01250(.dina(n1313), .dinb(n1303), .dout(n1314));
  jnot g01251(.din(n293), .dout(n1315));
  jor  g01252(.dina(n265), .dinb(n269), .dout(n1316));
  jor  g01253(.dina(n120), .dinb(n268), .dout(n1317));
  jand g01254(.dina(n1317), .dinb(n1316), .dout(n1318));
  jand g01255(.dina(n1318), .dinb(n1315), .dout(n1319));
  jand g01256(.dina(n542), .dinb(n838), .dout(n1320));
  jand g01257(.dina(n1245), .dinb(n470), .dout(n1321));
  jand g01258(.dina(n1321), .dinb(n1320), .dout(n1322));
  jand g01259(.dina(n1322), .dinb(n1319), .dout(n1323));
  jnot g01260(.din(n308), .dout(n1324));
  jor  g01261(.dina(n471), .dinb(n104), .dout(n1325));
  jand g01262(.dina(n1325), .dinb(n492), .dout(n1326));
  jor  g01263(.dina(n540), .dinb(n104), .dout(n1327));
  jand g01264(.dina(n1327), .dinb(n808), .dout(n1328));
  jand g01265(.dina(n1328), .dinb(n1326), .dout(n1329));
  jand g01266(.dina(n1329), .dinb(n1324), .dout(n1330));
  jand g01267(.dina(n1330), .dinb(n1323), .dout(n1331));
  jand g01268(.dina(n1331), .dinb(n1314), .dout(n1332));
  jnot g01269(.din(n333), .dout(n1333));
  jnot g01270(.din(n334), .dout(n1334));
  jand g01271(.dina(n699), .dinb(n480), .dout(n1335));
  jand g01272(.dina(n1335), .dinb(n1334), .dout(n1336));
  jand g01273(.dina(n1336), .dinb(n1333), .dout(n1337));
  jnot g01274(.din(n344), .dout(n1338));
  jand g01275(.dina(n1338), .dinb(n1337), .dout(n1339));
  jand g01276(.dina(n1339), .dinb(n329), .dout(n1340));
  jand g01277(.dina(n1340), .dinb(n1332), .dout(n1341));
  jnot g01278(.din(n358), .dout(n1342));
  jand g01279(.dina(n1342), .dinb(n352), .dout(n1343));
  jnot g01280(.din(n360), .dout(n1344));
  jor  g01281(.dina(n324), .dinb(n494), .dout(n1345));
  jor  g01282(.dina(n324), .dinb(n268), .dout(n1346));
  jand g01283(.dina(n1346), .dinb(n1345), .dout(n1347));
  jand g01284(.dina(n1347), .dinb(n1344), .dout(n1348));
  jor  g01285(.dina(n468), .dinb(n515), .dout(n1349));
  jand g01286(.dina(n1349), .dinb(n714), .dout(n1350));
  jor  g01287(.dina(n491), .dinb(n462), .dout(n1351));
  jand g01288(.dina(n1351), .dinb(n619), .dout(n1352));
  jand g01289(.dina(n1352), .dinb(n1350), .dout(n1353));
  jand g01290(.dina(n1353), .dinb(n1348), .dout(n1354));
  jnot g01291(.din(n377), .dout(n1355));
  jand g01292(.dina(n1355), .dinb(n1354), .dout(n1356));
  jand g01293(.dina(n1356), .dinb(n1343), .dout(n1357));
  jand g01294(.dina(n948), .dinb(n1036), .dout(n1358));
  jand g01295(.dina(n1358), .dinb(n512), .dout(n1359));
  jor  g01296(.dina(n324), .dinb(n460), .dout(n1360));
  jor  g01297(.dina(n462), .dinb(n107), .dout(n1361));
  jand g01298(.dina(n1361), .dinb(n1360), .dout(n1362));
  jand g01299(.dina(n453), .dinb(n1362), .dout(n1363));
  jand g01300(.dina(n1363), .dinb(n1359), .dout(n1364));
  jand g01301(.dina(n964), .dinb(n551), .dout(n1365));
  jor  g01302(.dina(n451), .dinb(n500), .dout(n1366));
  jor  g01303(.dina(n471), .dinb(n502), .dout(n1367));
  jand g01304(.dina(n1367), .dinb(n1366), .dout(n1368));
  jand g01305(.dina(n1368), .dinb(n1365), .dout(n1369));
  jnot g01306(.din(n404), .dout(n1370));
  jand g01307(.dina(n1370), .dinb(n1369), .dout(n1371));
  jand g01308(.dina(n1371), .dinb(n1364), .dout(n1372));
  jor  g01309(.dina(n441), .dinb(n451), .dout(n1373));
  jand g01310(.dina(n1373), .dinb(n411), .dout(n1374));
  jor  g01311(.dina(n462), .dinb(n322), .dout(n1375));
  jand g01312(.dina(n1375), .dinb(n716), .dout(n1376));
  jand g01313(.dina(n1376), .dinb(n1374), .dout(n1377));
  jor  g01314(.dina(n441), .dinb(n120), .dout(n1378));
  jand g01315(.dina(n818), .dinb(n1378), .dout(n1379));
  jand g01316(.dina(n696), .dinb(n988), .dout(n1380));
  jand g01317(.dina(n1380), .dinb(n1379), .dout(n1381));
  jand g01318(.dina(n1381), .dinb(n1377), .dout(n1382));
  jand g01319(.dina(n431), .dinb(n1382), .dout(n1383));
  jand g01320(.dina(n1383), .dinb(n1372), .dout(n1384));
  jand g01321(.dina(n1384), .dinb(n1357), .dout(n1385));
  jand g01322(.dina(n1385), .dinb(n1341), .dout(n1386));
  jand g01323(.dina(n1386), .dinb(n1300), .dout(n1387));
  jand g01324(.dina(n1387), .dinb(n123), .dout(n1388));
  jand g01325(.dina(n1255), .dinb(n1388), .dout(n1389));
  jor  g01326(.dina(n1389), .dinb(n726), .dout(n1390));
  jor  g01327(.dina(n1390), .dinb(n1256), .dout(n1391));
  jand g01328(.dina(n1391), .dinb(n1177), .dout(n1392));
  jnot g01329(.din(n842), .dout(n1393));
  jand g01330(.dina(n844), .dinb(n1393), .dout(n1394));
  jand g01331(.dina(n849), .dinb(n1394), .dout(n1395));
  jand g01332(.dina(n1395), .dinb(n839), .dout(n1396));
  jand g01333(.dina(n1396), .dinb(n836), .dout(n1397));
  jnot g01334(.din(n856), .dout(n1398));
  jnot g01335(.din(n858), .dout(n1399));
  jand g01336(.dina(n859), .dinb(n1399), .dout(n1400));
  jand g01337(.dina(n1400), .dinb(n1398), .dout(n1401));
  jnot g01338(.din(n867), .dout(n1402));
  jand g01339(.dina(n1402), .dinb(n1401), .dout(n1403));
  jand g01340(.dina(n875), .dinb(n1403), .dout(n1404));
  jand g01341(.dina(n1404), .dinb(n1397), .dout(n1405));
  jand g01342(.dina(n1405), .dinb(n822), .dout(n1406));
  jnot g01343(.din(n892), .dout(n1407));
  jand g01344(.dina(n896), .dinb(n1407), .dout(n1408));
  jand g01345(.dina(n904), .dinb(n1408), .dout(n1409));
  jand g01346(.dina(n910), .dinb(n1409), .dout(n1410));
  jand g01347(.dina(n1410), .dinb(n887), .dout(n1411));
  jand g01348(.dina(n1411), .dinb(n882), .dout(n1412));
  jand g01349(.dina(n1412), .dinb(n1406), .dout(n1413));
  jnot g01350(.din(n945), .dout(n1414));
  jnot g01351(.din(n947), .dout(n1415));
  jand g01352(.dina(n951), .dinb(n1415), .dout(n1416));
  jand g01353(.dina(n956), .dinb(n1416), .dout(n1417));
  jand g01354(.dina(n1417), .dinb(n1414), .dout(n1418));
  jnot g01355(.din(n963), .dout(n1419));
  jnot g01356(.din(n971), .dout(n1420));
  jand g01357(.dina(n1420), .dinb(n966), .dout(n1421));
  jand g01358(.dina(n1421), .dinb(n1419), .dout(n1422));
  jand g01359(.dina(n1422), .dinb(n695), .dout(n1423));
  jand g01360(.dina(n1423), .dinb(n1418), .dout(n1424));
  jand g01361(.dina(n1424), .dinb(n938), .dout(n1425));
  jor  g01362(.dina(n446), .dinb(n500), .dout(n1426));
  jand g01363(.dina(n1426), .dinb(n1304), .dout(n1427));
  jand g01364(.dina(n1218), .dinb(n1427), .dout(n1428));
  jor  g01365(.dina(n324), .dinb(n515), .dout(n1429));
  jor  g01366(.dina(n462), .dinb(n268), .dout(n1430));
  jand g01367(.dina(n1430), .dinb(n1429), .dout(n1431));
  jor  g01368(.dina(n500), .dinb(n455), .dout(n1432));
  jand g01369(.dina(n270), .dinb(n1432), .dout(n1433));
  jand g01370(.dina(n1433), .dinb(n1431), .dout(n1434));
  jand g01371(.dina(n1434), .dinb(n1428), .dout(n1435));
  jand g01372(.dina(n1435), .dinb(n994), .dout(n1436));
  jor  g01373(.dina(n439), .dinb(n515), .dout(n1437));
  jand g01374(.dina(n1437), .dinb(n1346), .dout(n1438));
  jand g01375(.dina(n1438), .dinb(n495), .dout(n1439));
  jnot g01376(.din(n1011), .dout(n1440));
  jand g01377(.dina(n1440), .dinb(n1439), .dout(n1441));
  jand g01378(.dina(n1441), .dinb(n1006), .dout(n1442));
  jand g01379(.dina(n1442), .dinb(n1436), .dout(n1443));
  jand g01380(.dina(n1018), .dinb(n1443), .dout(n1444));
  jand g01381(.dina(n1444), .dinb(n989), .dout(n1445));
  jand g01382(.dina(n1445), .dinb(n986), .dout(n1446));
  jand g01383(.dina(n1446), .dinb(n1425), .dout(n1447));
  jand g01384(.dina(n1447), .dinb(n1413), .dout(n1448));
  jnot g01385(.din(n342), .dout(n1449));
  jand g01386(.dina(n112), .dinb(n96), .dout(n1450));
  jnot g01387(.din(n1450), .dout(n1451));
  jand g01388(.dina(n1451), .dinb(n1449), .dout(n1452));
  jnot g01389(.din(n864), .dout(n1453));
  jand g01390(.dina(n1453), .dinb(n901), .dout(n1454));
  jand g01391(.dina(n1454), .dinb(n1452), .dout(n1455));
  jand g01392(.dina(n1455), .dinb(n978), .dout(n1456));
  jand g01393(.dina(n1456), .dinb(n349), .dout(n1457));
  jand g01394(.dina(n1457), .dinb(n1304), .dout(n1458));
  jand g01395(.dina(n948), .dinb(n1213), .dout(n1459));
  jnot g01396(.din(n1082), .dout(n1460));
  jand g01397(.dina(n1460), .dinb(n445), .dout(n1461));
  jand g01398(.dina(n1005), .dinb(n1205), .dout(n1462));
  jand g01399(.dina(n1462), .dinb(n1461), .dout(n1463));
  jand g01400(.dina(n1463), .dinb(n1459), .dout(n1464));
  jnot g01401(.din(n573), .dout(n1465));
  jand g01402(.dina(n1465), .dinb(n320), .dout(n1466));
  jand g01403(.dina(n1466), .dinb(n518), .dout(n1467));
  jand g01404(.dina(n1467), .dinb(n1167), .dout(n1468));
  jand g01405(.dina(n176), .dinb(n219), .dout(n1469));
  jnot g01406(.din(n1469), .dout(n1470));
  jand g01407(.dina(n1470), .dinb(n921), .dout(n1471));
  jand g01408(.dina(n1471), .dinb(n481), .dout(n1472));
  jand g01409(.dina(n1207), .dinb(n650), .dout(n1473));
  jand g01410(.dina(n1473), .dinb(n676), .dout(n1474));
  jand g01411(.dina(n1474), .dinb(n1472), .dout(n1475));
  jnot g01412(.din(n487), .dout(n1476));
  jand g01413(.dina(n1476), .dinb(n1315), .dout(n1477));
  jand g01414(.dina(n1107), .dinb(n555), .dout(n1478));
  jand g01415(.dina(n1478), .dinb(n1477), .dout(n1479));
  jand g01416(.dina(n1479), .dinb(n848), .dout(n1480));
  jand g01417(.dina(n1480), .dinb(n1475), .dout(n1481));
  jand g01418(.dina(n1481), .dinb(n1468), .dout(n1482));
  jand g01419(.dina(n1482), .dinb(n1464), .dout(n1483));
  jand g01420(.dina(n1483), .dinb(n1458), .dout(n1484));
  jand g01421(.dina(n442), .dinb(n1349), .dout(n1485));
  jand g01422(.dina(n1016), .dinb(n411), .dout(n1486));
  jand g01423(.dina(n1486), .dinb(n600), .dout(n1487));
  jand g01424(.dina(n1487), .dinb(n1485), .dout(n1488));
  jand g01425(.dina(n871), .dinb(n132), .dout(n1489));
  jand g01426(.dina(n824), .dinb(n469), .dout(n1490));
  jand g01427(.dina(n1490), .dinb(n1316), .dout(n1491));
  jand g01428(.dina(n1491), .dinb(n1489), .dout(n1492));
  jand g01429(.dina(n1492), .dinb(n1488), .dout(n1493));
  jand g01430(.dina(n1493), .dinb(n547), .dout(n1494));
  jnot g01431(.din(n609), .dout(n1495));
  jand g01432(.dina(n680), .dinb(n178), .dout(n1496));
  jand g01433(.dina(n1496), .dinb(n1495), .dout(n1497));
  jand g01434(.dina(n538), .dinb(n541), .dout(n1498));
  jand g01435(.dina(n1498), .dinb(n1497), .dout(n1499));
  jand g01436(.dina(n1367), .dinb(n270), .dout(n1500));
  jand g01437(.dina(n1500), .dinb(n893), .dout(n1501));
  jand g01438(.dina(n1501), .dinb(n1439), .dout(n1502));
  jand g01439(.dina(n1502), .dinb(n1499), .dout(n1503));
  jand g01440(.dina(n619), .dinb(n1327), .dout(n1504));
  jand g01441(.dina(n1504), .dinb(n92), .dout(n1505));
  jnot g01442(.din(n1064), .dout(n1506));
  jand g01443(.dina(n1506), .dinb(n716), .dout(n1507));
  jand g01444(.dina(n1507), .dinb(n450), .dout(n1508));
  jand g01445(.dina(n1508), .dinb(n1505), .dout(n1509));
  jand g01446(.dina(n169), .dinb(n133), .dout(n1510));
  jnot g01447(.din(n1510), .dout(n1511));
  jand g01448(.dina(n1189), .dinb(n562), .dout(n1512));
  jand g01449(.dina(n1512), .dinb(n1511), .dout(n1513));
  jand g01450(.dina(n551), .dinb(n1292), .dout(n1514));
  jnot g01451(.din(n1126), .dout(n1515));
  jand g01452(.dina(n1515), .dinb(n1361), .dout(n1516));
  jand g01453(.dina(n1516), .dinb(n1514), .dout(n1517));
  jand g01454(.dina(n1517), .dinb(n1513), .dout(n1518));
  jand g01455(.dina(n1518), .dinb(n1509), .dout(n1519));
  jand g01456(.dina(n1519), .dinb(n1503), .dout(n1520));
  jand g01457(.dina(n1520), .dinb(n1494), .dout(n1521));
  jnot g01458(.din(n890), .dout(n1522));
  jand g01459(.dina(n1522), .dinb(n843), .dout(n1523));
  jnot g01460(.din(n1057), .dout(n1524));
  jand g01461(.dina(n1524), .dinb(n907), .dout(n1525));
  jand g01462(.dina(n1525), .dinb(n1523), .dout(n1526));
  jand g01463(.dina(n532), .dinb(n1366), .dout(n1527));
  jand g01464(.dina(n430), .dinb(n454), .dout(n1528));
  jand g01465(.dina(n1528), .dinb(n1527), .dout(n1529));
  jand g01466(.dina(n1529), .dinb(n1526), .dout(n1530));
  jand g01467(.dina(n703), .dinb(n664), .dout(n1531));
  jnot g01468(.din(n841), .dout(n1532));
  jand g01469(.dina(n1532), .dinb(n121), .dout(n1533));
  jnot g01470(.din(n611), .dout(n1534));
  jand g01471(.dina(n149), .dinb(n98), .dout(n1535));
  jnot g01472(.din(n1535), .dout(n1536));
  jand g01473(.dina(n1536), .dinb(n1534), .dout(n1537));
  jand g01474(.dina(n1537), .dinb(n1533), .dout(n1538));
  jand g01475(.dina(n1538), .dinb(n1531), .dout(n1539));
  jand g01476(.dina(n1539), .dinb(n1530), .dout(n1540));
  jnot g01477(.din(n1025), .dout(n1541));
  jand g01478(.dina(n1541), .dinb(n1218), .dout(n1542));
  jand g01479(.dina(n1163), .dinb(n534), .dout(n1543));
  jand g01480(.dina(n1543), .dinb(n1542), .dout(n1544));
  jand g01481(.dina(n351), .dinb(n470), .dout(n1545));
  jand g01482(.dina(n1545), .dinb(n1429), .dout(n1546));
  jand g01483(.dina(n920), .dinb(n1273), .dout(n1547));
  jand g01484(.dina(n548), .dinb(n521), .dout(n1548));
  jand g01485(.dina(n1548), .dinb(n1547), .dout(n1549));
  jand g01486(.dina(n1549), .dinb(n1546), .dout(n1550));
  jand g01487(.dina(n1550), .dinb(n1544), .dout(n1551));
  jand g01488(.dina(n511), .dinb(n1334), .dout(n1552));
  jand g01489(.dina(n560), .dinb(n662), .dout(n1553));
  jand g01490(.dina(n1553), .dinb(n621), .dout(n1554));
  jand g01491(.dina(n1554), .dinb(n929), .dout(n1555));
  jand g01492(.dina(n1555), .dinb(n1552), .dout(n1556));
  jand g01493(.dina(n1556), .dinb(n1551), .dout(n1557));
  jand g01494(.dina(n1557), .dinb(n1540), .dout(n1558));
  jnot g01495(.din(n595), .dout(n1559));
  jnot g01496(.din(n941), .dout(n1560));
  jand g01497(.dina(n1560), .dinb(n1559), .dout(n1561));
  jand g01498(.dina(n691), .dinb(n630), .dout(n1562));
  jand g01499(.dina(n1562), .dinb(n1561), .dout(n1563));
  jand g01500(.dina(n1344), .dinb(n175), .dout(n1564));
  jand g01501(.dina(n1098), .dinb(n831), .dout(n1565));
  jand g01502(.dina(n1565), .dinb(n1564), .dout(n1566));
  jand g01503(.dina(n1566), .dinb(n1563), .dout(n1567));
  jand g01504(.dina(n1228), .dinb(n718), .dout(n1568));
  jnot g01505(.din(n960), .dout(n1569));
  jand g01506(.dina(n1569), .dinb(n447), .dout(n1570));
  jand g01507(.dina(n1570), .dinb(n1568), .dout(n1571));
  jand g01508(.dina(n1037), .dinb(n933), .dout(n1572));
  jand g01509(.dina(n1572), .dinb(n1571), .dout(n1573));
  jand g01510(.dina(n1573), .dinb(n1567), .dout(n1574));
  jnot g01511(.din(n216), .dout(n1575));
  jand g01512(.dina(n153), .dinb(n139), .dout(n1576));
  jnot g01513(.din(n1576), .dout(n1577));
  jand g01514(.dina(n1577), .dinb(n1575), .dout(n1578));
  jand g01515(.dina(n1325), .dinb(n880), .dout(n1579));
  jand g01516(.dina(n1203), .dinb(n811), .dout(n1580));
  jand g01517(.dina(n1580), .dinb(n1579), .dout(n1581));
  jand g01518(.dina(n1426), .dinb(n983), .dout(n1582));
  jnot g01519(.din(n854), .dout(n1583));
  jand g01520(.dina(n1583), .dinb(n632), .dout(n1584));
  jand g01521(.dina(n1584), .dinb(n1582), .dout(n1585));
  jand g01522(.dina(n1585), .dinb(n1581), .dout(n1586));
  jand g01523(.dina(n1586), .dinb(n1578), .dout(n1587));
  jand g01524(.dina(n1587), .dinb(n1574), .dout(n1588));
  jand g01525(.dina(n917), .dinb(n1310), .dout(n1589));
  jand g01526(.dina(n1589), .dinb(n135), .dout(n1590));
  jnot g01527(.din(n604), .dout(n1591));
  jand g01528(.dina(n1591), .dinb(n964), .dout(n1592));
  jand g01529(.dina(n645), .dinb(n553), .dout(n1593));
  jand g01530(.dina(n1593), .dinb(n1592), .dout(n1594));
  jand g01531(.dina(n1594), .dinb(n1590), .dout(n1595));
  jnot g01532(.din(n570), .dout(n1596));
  jand g01533(.dina(n908), .dinb(n1596), .dout(n1597));
  jand g01534(.dina(n586), .dinb(n1373), .dout(n1598));
  jand g01535(.dina(n1598), .dinb(n1247), .dout(n1599));
  jand g01536(.dina(n1599), .dinb(n504), .dout(n1600));
  jand g01537(.dina(n1600), .dinb(n1597), .dout(n1601));
  jand g01538(.dina(n1601), .dinb(n1595), .dout(n1602));
  jand g01539(.dina(n1602), .dinb(n1588), .dout(n1603));
  jand g01540(.dina(n1603), .dinb(n1558), .dout(n1604));
  jand g01541(.dina(n1604), .dinb(n1521), .dout(n1605));
  jand g01542(.dina(n1605), .dinb(n1484), .dout(n1606));
  jxor g01543(.dina(n1606), .dinb(n1448), .dout(n1607));
  jxor g01544(.dina(n1607), .dinb(n1392), .dout(n1608));
  jor  g01545(.dina(n1608), .dinb(n807), .dout(n1609));
  jnot g01546(.din(n804), .dout(n1610));
  jxor g01547(.dina(\a[22] ), .dinb(\a[21] ), .dout(n1611));
  jand g01548(.dina(n1611), .dinb(n1610), .dout(n1612));
  jnot g01549(.din(n1612), .dout(n1613));
  jor  g01550(.dina(n1613), .dinb(n1448), .dout(n1614));
  jnot g01551(.din(n805), .dout(n1615));
  jor  g01552(.dina(n1611), .dinb(n804), .dout(n1616));
  jor  g01553(.dina(n1616), .dinb(n1615), .dout(n1617));
  jor  g01554(.dina(n1617), .dinb(n1255), .dout(n1618));
  jand g01555(.dina(n1618), .dinb(n1614), .dout(n1619));
  jand g01556(.dina(n1615), .dinb(n804), .dout(n1620));
  jnot g01557(.din(n1620), .dout(n1621));
  jor  g01558(.dina(n1621), .dinb(n1606), .dout(n1622));
  jand g01559(.dina(n1622), .dinb(n1619), .dout(n1623));
  jand g01560(.dina(n1623), .dinb(n1609), .dout(n1624));
  jxor g01561(.dina(n1624), .dinb(\a[23] ), .dout(n1625));
  jor  g01562(.dina(n1625), .dinb(n803), .dout(n1626));
  jand g01563(.dina(n806), .dinb(n728), .dout(n1627));
  jand g01564(.dina(n1612), .dinb(n438), .dout(n1628));
  jand g01565(.dina(n1620), .dinb(n795), .dout(n1629));
  jor  g01566(.dina(n1629), .dinb(n1628), .dout(n1630));
  jor  g01567(.dina(n1630), .dinb(n1627), .dout(n1631));
  jnot g01568(.din(n1631), .dout(n1632));
  jand g01569(.dina(n804), .dinb(n438), .dout(n1633));
  jnot g01570(.din(n1633), .dout(n1634));
  jand g01571(.dina(n1634), .dinb(\a[23] ), .dout(n1635));
  jand g01572(.dina(n1635), .dinb(n1632), .dout(n1636));
  jand g01573(.dina(n795), .dinb(n1388), .dout(n1637));
  jxor g01574(.dina(n1255), .dinb(n1637), .dout(n1638));
  jnot g01575(.din(n1638), .dout(n1639));
  jand g01576(.dina(n1639), .dinb(n806), .dout(n1640));
  jand g01577(.dina(n1612), .dinb(n795), .dout(n1641));
  jand g01578(.dina(n1620), .dinb(n1175), .dout(n1642));
  jor  g01579(.dina(n1642), .dinb(n1641), .dout(n1643));
  jnot g01580(.din(n1617), .dout(n1644));
  jand g01581(.dina(n1644), .dinb(n438), .dout(n1645));
  jor  g01582(.dina(n1645), .dinb(n1643), .dout(n1646));
  jor  g01583(.dina(n1646), .dinb(n1640), .dout(n1647));
  jnot g01584(.din(n1647), .dout(n1648));
  jand g01585(.dina(n1648), .dinb(n1636), .dout(n1649));
  jand g01586(.dina(n1649), .dinb(n800), .dout(n1650));
  jnot g01587(.din(n1650), .dout(n1651));
  jxor g01588(.dina(n1649), .dinb(n800), .dout(n1652));
  jnot g01589(.din(n1652), .dout(n1653));
  jor  g01590(.dina(n1175), .dinb(n438), .dout(n1654));
  jand g01591(.dina(n1654), .dinb(n795), .dout(n1655));
  jxor g01592(.dina(n1655), .dinb(n1256), .dout(n1656));
  jor  g01593(.dina(n1656), .dinb(n807), .dout(n1657));
  jor  g01594(.dina(n1621), .dinb(n1448), .dout(n1658));
  jor  g01595(.dina(n1613), .dinb(n1255), .dout(n1659));
  jand g01596(.dina(n1659), .dinb(n1658), .dout(n1660));
  jor  g01597(.dina(n1617), .dinb(n726), .dout(n1661));
  jand g01598(.dina(n1661), .dinb(n1660), .dout(n1662));
  jand g01599(.dina(n1662), .dinb(n1657), .dout(n1663));
  jxor g01600(.dina(n1663), .dinb(\a[23] ), .dout(n1664));
  jor  g01601(.dina(n1664), .dinb(n1653), .dout(n1665));
  jand g01602(.dina(n1665), .dinb(n1651), .dout(n1666));
  jnot g01603(.din(n1666), .dout(n1667));
  jxor g01604(.dina(n1625), .dinb(n803), .dout(n1668));
  jand g01605(.dina(n1668), .dinb(n1667), .dout(n1669));
  jnot g01606(.din(n1669), .dout(n1670));
  jand g01607(.dina(n1670), .dinb(n1626), .dout(n1671));
  jnot g01608(.din(n1671), .dout(n1672));
  jnot g01609(.din(n1606), .dout(n1673));
  jand g01610(.dina(n1673), .dinb(n1024), .dout(n1674));
  jnot g01611(.din(n1674), .dout(n1675));
  jnot g01612(.din(n1607), .dout(n1676));
  jor  g01613(.dina(n1676), .dinb(n1392), .dout(n1677));
  jand g01614(.dina(n1677), .dinb(n1675), .dout(n1678));
  jand g01615(.dina(n873), .dinb(n1532), .dout(n1679));
  jand g01616(.dina(n1577), .dinb(n933), .dout(n1680));
  jand g01617(.dina(n1680), .dinb(n1679), .dout(n1681));
  jnot g01618(.din(n403), .dout(n1682));
  jand g01619(.dina(n534), .dinb(n1682), .dout(n1683));
  jand g01620(.dina(n1683), .dinb(n465), .dout(n1684));
  jand g01621(.dina(n1684), .dinb(n1681), .dout(n1685));
  jand g01622(.dina(n447), .dinb(n818), .dout(n1686));
  jand g01623(.dina(n826), .dinb(n900), .dout(n1687));
  jand g01624(.dina(n1036), .dinb(n1288), .dout(n1688));
  jand g01625(.dina(n1688), .dinb(n1687), .dout(n1689));
  jand g01626(.dina(n1689), .dinb(n1686), .dout(n1690));
  jand g01627(.dina(n1690), .dinb(n1685), .dout(n1691));
  jand g01628(.dina(n1691), .dinb(n1275), .dout(n1692));
  jand g01629(.dina(n557), .dinb(n831), .dout(n1693));
  jand g01630(.dina(n1693), .dinb(n521), .dout(n1694));
  jand g01631(.dina(n1694), .dinb(n921), .dout(n1695));
  jand g01632(.dina(n1460), .dinb(n650), .dout(n1696));
  jnot g01633(.din(n569), .dout(n1697));
  jand g01634(.dina(n978), .dinb(n1697), .dout(n1698));
  jand g01635(.dina(n1698), .dinb(n1696), .dout(n1699));
  jand g01636(.dina(n1212), .dinb(n931), .dout(n1700));
  jnot g01637(.din(n187), .dout(n1701));
  jand g01638(.dina(n1451), .dinb(n1701), .dout(n1702));
  jand g01639(.dina(n1702), .dinb(n1700), .dout(n1703));
  jand g01640(.dina(n1703), .dinb(n1699), .dout(n1704));
  jand g01641(.dina(n1159), .dinb(n1315), .dout(n1705));
  jand g01642(.dina(n1705), .dinb(n668), .dout(n1706));
  jand g01643(.dina(n670), .dinb(n560), .dout(n1707));
  jnot g01644(.din(n477), .dout(n1708));
  jand g01645(.dina(n1708), .dinb(n517), .dout(n1709));
  jand g01646(.dina(n1709), .dinb(n1707), .dout(n1710));
  jand g01647(.dina(n1710), .dinb(n1706), .dout(n1711));
  jand g01648(.dina(n1711), .dinb(n1704), .dout(n1712));
  jnot g01649(.din(n1080), .dout(n1713));
  jand g01650(.dina(n1713), .dinb(n1378), .dout(n1714));
  jand g01651(.dina(n1714), .dinb(n630), .dout(n1715));
  jand g01652(.dina(n638), .dinb(n542), .dout(n1716));
  jand g01653(.dina(n983), .dinb(n493), .dout(n1717));
  jand g01654(.dina(n1717), .dinb(n1716), .dout(n1718));
  jand g01655(.dina(n1718), .dinb(n1715), .dout(n1719));
  jand g01656(.dina(n186), .dinb(n176), .dout(n1720));
  jnot g01657(.din(n1720), .dout(n1721));
  jand g01658(.dina(n583), .dinb(n100), .dout(n1722));
  jand g01659(.dina(n621), .dinb(n1304), .dout(n1723));
  jand g01660(.dina(n1723), .dinb(n1722), .dout(n1724));
  jand g01661(.dina(n1724), .dinb(n1721), .dout(n1725));
  jand g01662(.dina(n1725), .dinb(n1719), .dout(n1726));
  jand g01663(.dina(n1726), .dinb(n1712), .dout(n1727));
  jand g01664(.dina(n1727), .dinb(n1695), .dout(n1728));
  jand g01665(.dina(n1728), .dinb(n1692), .dout(n1729));
  jand g01666(.dina(n183), .dinb(n143), .dout(n1730));
  jnot g01667(.din(n1730), .dout(n1731));
  jand g01668(.dina(n1731), .dinb(n672), .dout(n1732));
  jand g01669(.dina(n1732), .dinb(n1042), .dout(n1733));
  jand g01670(.dina(n1733), .dinb(n1521), .dout(n1734));
  jand g01671(.dina(n1470), .dinb(n1305), .dout(n1735));
  jand g01672(.dina(n440), .dinb(n654), .dout(n1736));
  jand g01673(.dina(n1736), .dinb(n1735), .dout(n1737));
  jnot g01674(.din(n354), .dout(n1738));
  jand g01675(.dina(n1375), .dinb(n320), .dout(n1739));
  jand g01676(.dina(n1739), .dinb(n1738), .dout(n1740));
  jand g01677(.dina(n1740), .dinb(n1737), .dout(n1741));
  jand g01678(.dina(n86), .dinb(n76), .dout(n1742));
  jnot g01679(.din(n1742), .dout(n1743));
  jand g01680(.dina(n1743), .dinb(n703), .dout(n1744));
  jand g01681(.dina(n1744), .dinb(n701), .dout(n1745));
  jand g01682(.dina(n1053), .dinb(n1088), .dout(n1746));
  jand g01683(.dina(n929), .dinb(n1188), .dout(n1747));
  jand g01684(.dina(n1747), .dinb(n1746), .dout(n1748));
  jand g01685(.dina(n1748), .dinb(n1745), .dout(n1749));
  jand g01686(.dina(n1749), .dinb(n1741), .dout(n1750));
  jand g01687(.dina(n514), .dinb(n829), .dout(n1751));
  jand g01688(.dina(n1090), .dinb(n693), .dout(n1752));
  jand g01689(.dina(n349), .dinb(n1283), .dout(n1753));
  jand g01690(.dina(n1753), .dinb(n1752), .dout(n1754));
  jand g01691(.dina(n1754), .dinb(n1751), .dout(n1755));
  jnot g01692(.din(n574), .dout(n1756));
  jand g01693(.dina(n1756), .dinb(n1225), .dout(n1757));
  jand g01694(.dina(n1757), .dinb(n848), .dout(n1758));
  jand g01695(.dina(n1758), .dinb(n887), .dout(n1759));
  jand g01696(.dina(n1759), .dinb(n1755), .dout(n1760));
  jand g01697(.dina(n1760), .dinb(n1750), .dout(n1761));
  jand g01698(.dina(n993), .dinb(n696), .dout(n1762));
  jand g01699(.dina(n1476), .dinb(n456), .dout(n1763));
  jand g01700(.dina(n1763), .dinb(n1762), .dout(n1764));
  jand g01701(.dina(n1107), .dinb(n653), .dout(n1765));
  jand g01702(.dina(n1765), .dinb(n981), .dout(n1766));
  jand g01703(.dina(n1522), .dinb(n1430), .dout(n1767));
  jand g01704(.dina(n718), .dinb(n1213), .dout(n1768));
  jand g01705(.dina(n1768), .dinb(n1767), .dout(n1769));
  jand g01706(.dina(n1769), .dinb(n1766), .dout(n1770));
  jand g01707(.dina(n169), .dinb(n139), .dout(n1771));
  jnot g01708(.din(n1771), .dout(n1772));
  jand g01709(.dina(n1772), .dinb(n683), .dout(n1773));
  jand g01710(.dina(n645), .dinb(n1345), .dout(n1774));
  jand g01711(.dina(n1774), .dinb(n1773), .dout(n1775));
  jand g01712(.dina(n1775), .dinb(n950), .dout(n1776));
  jand g01713(.dina(n1776), .dinb(n1770), .dout(n1777));
  jnot g01714(.din(n623), .dout(n1778));
  jand g01715(.dina(n1778), .dinb(n428), .dout(n1779));
  jand g01716(.dina(n1541), .dinb(n916), .dout(n1780));
  jand g01717(.dina(n1780), .dinb(n1779), .dout(n1781));
  jnot g01718(.din(n1067), .dout(n1782));
  jand g01719(.dina(n1536), .dinb(n114), .dout(n1783));
  jand g01720(.dina(n1783), .dinb(n1782), .dout(n1784));
  jand g01721(.dina(n1784), .dinb(n1781), .dout(n1785));
  jand g01722(.dina(n1785), .dinb(n1777), .dout(n1786));
  jand g01723(.dina(n1786), .dinb(n1764), .dout(n1787));
  jand g01724(.dina(n1787), .dinb(n1761), .dout(n1788));
  jand g01725(.dina(n1788), .dinb(n1734), .dout(n1789));
  jand g01726(.dina(n1789), .dinb(n1729), .dout(n1790));
  jxor g01727(.dina(n1790), .dinb(n1606), .dout(n1791));
  jxor g01728(.dina(n1791), .dinb(n1678), .dout(n1792));
  jor  g01729(.dina(n1792), .dinb(n807), .dout(n1793));
  jor  g01730(.dina(n1790), .dinb(n1621), .dout(n1794));
  jor  g01731(.dina(n1617), .dinb(n1448), .dout(n1795));
  jor  g01732(.dina(n1613), .dinb(n1606), .dout(n1796));
  jand g01733(.dina(n1796), .dinb(n1795), .dout(n1797));
  jand g01734(.dina(n1797), .dinb(n1794), .dout(n1798));
  jand g01735(.dina(n1798), .dinb(n1793), .dout(n1799));
  jxor g01736(.dina(n1799), .dinb(n65), .dout(n1800));
  jand g01737(.dina(n1639), .dinb(n71), .dout(n1801));
  jand g01738(.dina(n731), .dinb(n795), .dout(n1802));
  jand g01739(.dina(n1175), .dinb(n796), .dout(n1803));
  jor  g01740(.dina(n1803), .dinb(n1802), .dout(n1804));
  jand g01741(.dina(n468), .dinb(n455), .dout(n1805));
  jnot g01742(.din(n1805), .dout(n1806));
  jand g01743(.dina(n1806), .dinb(n438), .dout(n1807));
  jor  g01744(.dina(n1807), .dinb(n1804), .dout(n1808));
  jor  g01745(.dina(n1808), .dinb(n1801), .dout(n1809));
  jor  g01746(.dina(n800), .dinb(n77), .dout(n1810));
  jor  g01747(.dina(n1810), .dinb(n799), .dout(n1811));
  jand g01748(.dina(n1811), .dinb(\a[26] ), .dout(n1812));
  jxor g01749(.dina(n1812), .dinb(n1809), .dout(n1813));
  jxor g01750(.dina(n1813), .dinb(n1800), .dout(n1814));
  jxor g01751(.dina(n1814), .dinb(n1672), .dout(n1815));
  jnot g01752(.din(n1815), .dout(n1816));
  jxor g01753(.dina(\a[18] ), .dinb(\a[17] ), .dout(n1817));
  jxor g01754(.dina(\a[20] ), .dinb(\a[19] ), .dout(n1818));
  jand g01755(.dina(n1818), .dinb(n1817), .dout(n1819));
  jnot g01756(.din(n1819), .dout(n1820));
  jand g01757(.dina(n537), .dinb(n988), .dout(n1821));
  jnot g01758(.din(n340), .dout(n1822));
  jand g01759(.dina(n1822), .dinb(n480), .dout(n1823));
  jand g01760(.dina(n445), .dinb(n1238), .dout(n1824));
  jand g01761(.dina(n1824), .dinb(n1823), .dout(n1825));
  jand g01762(.dina(n1825), .dinb(n1821), .dout(n1826));
  jand g01763(.dina(n650), .dinb(n1349), .dout(n1827));
  jand g01764(.dina(n1162), .dinb(n978), .dout(n1828));
  jand g01765(.dina(n1828), .dinb(n1827), .dout(n1829));
  jand g01766(.dina(n1829), .dinb(n925), .dout(n1830));
  jand g01767(.dina(n1830), .dinb(n1826), .dout(n1831));
  jand g01768(.dina(n1756), .dinb(n948), .dout(n1832));
  jand g01769(.dina(n1832), .dinb(n678), .dout(n1833));
  jand g01770(.dina(n654), .dinb(n1205), .dout(n1834));
  jand g01771(.dina(n1042), .dinb(n908), .dout(n1835));
  jand g01772(.dina(n1835), .dinb(n1834), .dout(n1836));
  jand g01773(.dina(n1836), .dinb(n1833), .dout(n1837));
  jand g01774(.dina(n1370), .dinb(n829), .dout(n1838));
  jand g01775(.dina(n1838), .dinb(n900), .dout(n1839));
  jand g01776(.dina(n1839), .dinb(n1837), .dout(n1840));
  jand g01777(.dina(n1840), .dinb(n1831), .dout(n1841));
  jand g01778(.dina(n1841), .dinb(n1283), .dout(n1842));
  jand g01779(.dina(n270), .dinb(n920), .dout(n1843));
  jand g01780(.dina(n1843), .dinb(n1426), .dout(n1844));
  jand g01781(.dina(n146), .dinb(n112), .dout(n1845));
  jnot g01782(.din(n1845), .dout(n1846));
  jand g01783(.dina(n1846), .dinb(n1053), .dout(n1847));
  jand g01784(.dina(n1847), .dinb(n1559), .dout(n1848));
  jand g01785(.dina(n1848), .dinb(n1844), .dout(n1849));
  jand g01786(.dina(n1849), .dinb(n1005), .dout(n1850));
  jand g01787(.dina(n695), .dinb(n901), .dout(n1851));
  jand g01788(.dina(n1373), .dinb(n916), .dout(n1852));
  jand g01789(.dina(n1591), .dinb(n442), .dout(n1853));
  jand g01790(.dina(n1853), .dinb(n638), .dout(n1854));
  jand g01791(.dina(n514), .dinb(n1378), .dout(n1855));
  jand g01792(.dina(n1855), .dinb(n1247), .dout(n1856));
  jand g01793(.dina(n1856), .dinb(n1854), .dout(n1857));
  jand g01794(.dina(n1857), .dinb(n1852), .dout(n1858));
  jand g01795(.dina(n1858), .dinb(n1851), .dout(n1859));
  jand g01796(.dina(n1859), .dinb(n1850), .dout(n1860));
  jand g01797(.dina(n1344), .dinb(n1088), .dout(n1861));
  jand g01798(.dina(n1861), .dinb(n101), .dout(n1862));
  jand g01799(.dina(n873), .dinb(n700), .dout(n1863));
  jand g01800(.dina(n1863), .dinb(n1862), .dout(n1864));
  jand g01801(.dina(n993), .dinb(n1351), .dout(n1865));
  jand g01802(.dina(n1865), .dinb(n1037), .dout(n1866));
  jnot g01803(.din(n1066), .dout(n1867));
  jand g01804(.dina(n1212), .dinb(n1867), .dout(n1868));
  jand g01805(.dina(n647), .dinb(n472), .dout(n1869));
  jand g01806(.dina(n1869), .dinb(n1868), .dout(n1870));
  jand g01807(.dina(n1870), .dinb(n1866), .dout(n1871));
  jand g01808(.dina(n1237), .dinb(n1361), .dout(n1872));
  jand g01809(.dina(n826), .dinb(n510), .dout(n1873));
  jand g01810(.dina(n1873), .dinb(n1872), .dout(n1874));
  jand g01811(.dina(n1874), .dinb(n1871), .dout(n1875));
  jand g01812(.dina(n1875), .dinb(n1864), .dout(n1876));
  jand g01813(.dina(n542), .dinb(n933), .dout(n1877));
  jand g01814(.dina(n1877), .dinb(n1565), .dout(n1878));
  jand g01815(.dina(n1878), .dinb(n691), .dout(n1879));
  jand g01816(.dina(n1879), .dinb(n1876), .dout(n1880));
  jand g01817(.dina(n1880), .dinb(n1860), .dout(n1881));
  jand g01818(.dina(n1881), .dinb(n1842), .dout(n1882));
  jand g01819(.dina(n1545), .dinb(n326), .dout(n1883));
  jand g01820(.dina(n880), .dinb(n121), .dout(n1884));
  jand g01821(.dina(n1884), .dinb(n1783), .dout(n1885));
  jand g01822(.dina(n1885), .dinb(n1883), .dout(n1886));
  jand g01823(.dina(n1886), .dinb(n870), .dout(n1887));
  jand g01824(.dina(n1233), .dinb(n493), .dout(n1888));
  jand g01825(.dina(n1888), .dinb(n696), .dout(n1889));
  jand g01826(.dina(n1743), .dinb(n1245), .dout(n1890));
  jand g01827(.dina(n1375), .dinb(n555), .dout(n1891));
  jand g01828(.dina(n1891), .dinb(n499), .dout(n1892));
  jand g01829(.dina(n1892), .dinb(n1890), .dout(n1893));
  jand g01830(.dina(n1893), .dinb(n1889), .dout(n1894));
  jand g01831(.dina(n1894), .dinb(n1887), .dout(n1895));
  jand g01832(.dina(n1895), .dinb(n1167), .dout(n1896));
  jand g01833(.dina(n1896), .dinb(n895), .dout(n1897));
  jand g01834(.dina(n1228), .dinb(n1399), .dout(n1898));
  jand g01835(.dina(n621), .dinb(n929), .dout(n1899));
  jand g01836(.dina(n428), .dinb(n893), .dout(n1900));
  jand g01837(.dina(n1900), .dinb(n1899), .dout(n1901));
  jand g01838(.dina(n1901), .dinb(n1898), .dout(n1902));
  jnot g01839(.din(n624), .dout(n1903));
  jand g01840(.dina(n1903), .dinb(n1040), .dout(n1904));
  jand g01841(.dina(n1904), .dinb(n549), .dout(n1905));
  jand g01842(.dina(n1905), .dinb(n440), .dout(n1906));
  jand g01843(.dina(n1906), .dinb(n1902), .dout(n1907));
  jand g01844(.dina(n1453), .dinb(n848), .dout(n1908));
  jand g01845(.dina(n1908), .dinb(n917), .dout(n1909));
  jand g01846(.dina(n1909), .dinb(n653), .dout(n1910));
  jand g01847(.dina(n1910), .dinb(n1495), .dout(n1911));
  jand g01848(.dina(n461), .dinb(n1334), .dout(n1912));
  jand g01849(.dina(n1912), .dinb(n982), .dout(n1913));
  jand g01850(.dina(n1913), .dinb(n1328), .dout(n1914));
  jand g01851(.dina(n1583), .dinb(n668), .dout(n1915));
  jand g01852(.dina(n630), .dinb(n1316), .dout(n1916));
  jand g01853(.dina(n1916), .dinb(n818), .dout(n1917));
  jand g01854(.dina(n1917), .dinb(n1915), .dout(n1918));
  jand g01855(.dina(n1918), .dinb(n1914), .dout(n1919));
  jand g01856(.dina(n1919), .dinb(n1911), .dout(n1920));
  jand g01857(.dina(n1920), .dinb(n1907), .dout(n1921));
  jand g01858(.dina(n551), .dinb(n1317), .dout(n1922));
  jand g01859(.dina(n1922), .dinb(n1532), .dout(n1923));
  jand g01860(.dina(n1430), .dinb(n130), .dout(n1924));
  jand g01861(.dina(n582), .dinb(n501), .dout(n1925));
  jand g01862(.dina(n1925), .dinb(n1924), .dout(n1926));
  jand g01863(.dina(n1926), .dinb(n1923), .dout(n1927));
  jand g01864(.dina(n1731), .dinb(n1360), .dout(n1928));
  jnot g01865(.din(n1065), .dout(n1929));
  jand g01866(.dina(n660), .dinb(n349), .dout(n1930));
  jand g01867(.dina(n1930), .dinb(n1929), .dout(n1931));
  jand g01868(.dina(n1931), .dinb(n1928), .dout(n1932));
  jand g01869(.dina(n1449), .dinb(n1309), .dout(n1933));
  jand g01870(.dina(n456), .dinb(n1292), .dout(n1934));
  jand g01871(.dina(n1934), .dinb(n1933), .dout(n1935));
  jand g01872(.dina(n1345), .dinb(n168), .dout(n1936));
  jand g01873(.dina(n1936), .dinb(n1935), .dout(n1937));
  jand g01874(.dina(n1937), .dinb(n1932), .dout(n1938));
  jand g01875(.dina(n1938), .dinb(n1927), .dout(n1939));
  jnot g01876(.din(n944), .dout(n1940));
  jand g01877(.dina(n1735), .dinb(n1325), .dout(n1941));
  jand g01878(.dina(n1941), .dinb(n1515), .dout(n1942));
  jand g01879(.dina(n1090), .dinb(n964), .dout(n1943));
  jand g01880(.dina(n1697), .dinb(n1432), .dout(n1944));
  jand g01881(.dina(n1944), .dinb(n1943), .dout(n1945));
  jand g01882(.dina(n645), .dinb(n676), .dout(n1946));
  jand g01883(.dina(n1946), .dinb(n1541), .dout(n1947));
  jand g01884(.dina(n1947), .dinb(n1945), .dout(n1948));
  jand g01885(.dina(n1948), .dinb(n1942), .dout(n1949));
  jand g01886(.dina(n1949), .dinb(n1940), .dout(n1950));
  jand g01887(.dina(n1950), .dinb(n1939), .dout(n1951));
  jand g01888(.dina(n1951), .dinb(n1921), .dout(n1952));
  jand g01889(.dina(n1952), .dinb(n1897), .dout(n1953));
  jand g01890(.dina(n1953), .dinb(n1882), .dout(n1954));
  jnot g01891(.din(n1954), .dout(n1955));
  jand g01892(.dina(n925), .dinb(n450), .dout(n1956));
  jand g01893(.dina(n1449), .dinb(n920), .dout(n1957));
  jand g01894(.dina(n1957), .dinb(n1956), .dout(n1958));
  jand g01895(.dina(n1958), .dinb(n1053), .dout(n1959));
  jand g01896(.dina(n672), .dinb(n1347), .dout(n1960));
  jand g01897(.dina(n1506), .dinb(n521), .dout(n1961));
  jand g01898(.dina(n1961), .dinb(n1960), .dout(n1962));
  jand g01899(.dina(n1962), .dinb(n1959), .dout(n1963));
  jand g01900(.dina(n1569), .dinb(n1310), .dout(n1964));
  jand g01901(.dina(n1964), .dinb(n555), .dout(n1965));
  jand g01902(.dina(n718), .dinb(n1226), .dout(n1966));
  jand g01903(.dina(n1966), .dinb(n1965), .dout(n1967));
  jand g01904(.dina(n1237), .dinb(n1098), .dout(n1968));
  jand g01905(.dina(n1968), .dinb(n685), .dout(n1969));
  jand g01906(.dina(n1969), .dinb(n1967), .dout(n1970));
  jand g01907(.dina(n1772), .dinb(n1515), .dout(n1971));
  jand g01908(.dina(n1852), .dinb(n978), .dout(n1972));
  jand g01909(.dina(n1972), .dinb(n1971), .dout(n1973));
  jand g01910(.dina(n1973), .dinb(n545), .dout(n1974));
  jand g01911(.dina(n1974), .dinb(n1970), .dout(n1975));
  jnot g01912(.din(n970), .dout(n1976));
  jand g01913(.dina(n548), .dinb(n1360), .dout(n1977));
  jand g01914(.dina(n1977), .dinb(n1976), .dout(n1978));
  jand g01915(.dina(n1713), .dinb(n848), .dout(n1979));
  jand g01916(.dina(n1979), .dinb(n1708), .dout(n1980));
  jand g01917(.dina(n1980), .dinb(n1978), .dout(n1981));
  jand g01918(.dina(n1868), .dinb(n1756), .dout(n1982));
  jand g01919(.dina(n1982), .dinb(n928), .dout(n1983));
  jand g01920(.dina(n1983), .dinb(n1981), .dout(n1984));
  jand g01921(.dina(n1984), .dinb(n1975), .dout(n1985));
  jand g01922(.dina(n1985), .dinb(n1963), .dout(n1986));
  jand g01923(.dina(n553), .dinb(n493), .dout(n1987));
  jand g01924(.dina(n1987), .dinb(n1219), .dout(n1988));
  jand g01925(.dina(n1534), .dinb(n1270), .dout(n1989));
  jand g01926(.dina(n829), .dinb(n1273), .dout(n1990));
  jand g01927(.dina(n1990), .dinb(n1989), .dout(n1991));
  jand g01928(.dina(n1991), .dinb(n1988), .dout(n1992));
  jand g01929(.dina(n1992), .dinb(n271), .dout(n1993));
  jand g01930(.dina(n1993), .dinb(n658), .dout(n1994));
  jand g01931(.dina(n1366), .dinb(n501), .dout(n1995));
  jand g01932(.dina(n1995), .dinb(n517), .dout(n1996));
  jand g01933(.dina(n1532), .dinb(n452), .dout(n1997));
  jand g01934(.dina(n1997), .dinb(n583), .dout(n1998));
  jand g01935(.dina(n693), .dinb(n964), .dout(n1999));
  jand g01936(.dina(n1437), .dinb(n1188), .dout(n2000));
  jand g01937(.dina(n2000), .dinb(n1999), .dout(n2001));
  jand g01938(.dina(n2001), .dinb(n1998), .dout(n2002));
  jand g01939(.dina(n2002), .dinb(n1996), .dout(n2003));
  jand g01940(.dina(n1823), .dinb(n1580), .dout(n2004));
  jand g01941(.dina(n2004), .dinb(n816), .dout(n2005));
  jand g01942(.dina(n2005), .dinb(n2003), .dout(n2006));
  jand g01943(.dina(n2006), .dinb(n1994), .dout(n2007));
  jand g01944(.dina(n869), .dinb(n991), .dout(n2008));
  jand g01945(.dina(n2008), .dinb(n1315), .dout(n2009));
  jand g01946(.dina(n2009), .dinb(n463), .dout(n2010));
  jand g01947(.dina(n1451), .dinb(n1378), .dout(n2011));
  jand g01948(.dina(n351), .dinb(n1309), .dout(n2012));
  jand g01949(.dina(n2012), .dinb(n2011), .dout(n2013));
  jand g01950(.dina(n2013), .dinb(n2010), .dout(n2014));
  jand g01951(.dina(n1779), .dinb(n1038), .dout(n2015));
  jand g01952(.dina(n2015), .dinb(n1218), .dout(n2016));
  jand g01953(.dina(n2016), .dinb(n2014), .dout(n2017));
  jand g01954(.dina(n2017), .dinb(n2007), .dout(n2018));
  jnot g01955(.din(n1045), .dout(n2019));
  jand g01956(.dina(n908), .dinb(n824), .dout(n2020));
  jand g01957(.dina(n2020), .dinb(n1461), .dout(n2021));
  jand g01958(.dina(n2021), .dinb(n2019), .dout(n2022));
  jnot g01959(.din(n1063), .dout(n2023));
  jand g01960(.dina(n2023), .dinb(n1334), .dout(n2024));
  jand g01961(.dina(n2024), .dinb(n588), .dout(n2025));
  jand g01962(.dina(n2025), .dinb(n1327), .dout(n2026));
  jand g01963(.dina(n2026), .dinb(n2022), .dout(n2027));
  jnot g01964(.din(n578), .dout(n2028));
  jand g01965(.dina(n461), .dinb(n683), .dout(n2029));
  jand g01966(.dina(n2029), .dinb(n2028), .dout(n2030));
  jand g01967(.dina(n1522), .dinb(n716), .dout(n2031));
  jand g01968(.dina(n1743), .dinb(n503), .dout(n2032));
  jand g01969(.dina(n2032), .dinb(n2031), .dout(n2033));
  jand g01970(.dina(n2033), .dinb(n1429), .dout(n2034));
  jand g01971(.dina(n2034), .dinb(n2030), .dout(n2035));
  jand g01972(.dina(n2035), .dinb(n2027), .dout(n2036));
  jand g01973(.dina(n514), .dinb(n582), .dout(n2037));
  jand g01974(.dina(n2037), .dinb(n1213), .dout(n2038));
  jand g01975(.dina(n1162), .dinb(n662), .dout(n2039));
  jand g01976(.dina(n2039), .dinb(n1349), .dout(n2040));
  jand g01977(.dina(n2040), .dinb(n2038), .dout(n2041));
  jand g01978(.dina(n808), .dinb(n114), .dout(n2042));
  jand g01979(.dina(n1701), .dinb(n132), .dout(n2043));
  jand g01980(.dina(n2043), .dinb(n1189), .dout(n2044));
  jand g01981(.dina(n2044), .dinb(n2042), .dout(n2045));
  jand g01982(.dina(n2045), .dinb(n2041), .dout(n2046));
  jand g01983(.dina(n826), .dinb(n1325), .dout(n2047));
  jand g01984(.dina(n2047), .dinb(n563), .dout(n2048));
  jand g01985(.dina(n2048), .dinb(n1236), .dout(n2049));
  jand g01986(.dina(n2049), .dinb(n2046), .dout(n2050));
  jand g01987(.dina(n2050), .dinb(n2036), .dout(n2051));
  jand g01988(.dina(n1591), .dinb(n1245), .dout(n2052));
  jand g01989(.dina(n993), .dinb(n430), .dout(n2053));
  jand g01990(.dina(n2053), .dinb(n2052), .dout(n2054));
  jand g01991(.dina(n2054), .dinb(n2051), .dout(n2055));
  jand g01992(.dina(n2055), .dinb(n2018), .dout(n2056));
  jand g01993(.dina(n2056), .dinb(n1986), .dout(n2057));
  jnot g01994(.din(n2057), .dout(n2058));
  jand g01995(.dina(n2058), .dinb(n1955), .dout(n2059));
  jnot g01996(.din(n2059), .dout(n2060));
  jnot g01997(.din(n1790), .dout(n2061));
  jand g01998(.dina(n2058), .dinb(n2061), .dout(n2062));
  jnot g01999(.din(n2062), .dout(n2063));
  jand g02000(.dina(n2061), .dinb(n1673), .dout(n2064));
  jnot g02001(.din(n2064), .dout(n2065));
  jnot g02002(.din(n1791), .dout(n2066));
  jor  g02003(.dina(n2066), .dinb(n1678), .dout(n2067));
  jand g02004(.dina(n2067), .dinb(n2065), .dout(n2068));
  jxor g02005(.dina(n2057), .dinb(n1790), .dout(n2069));
  jnot g02006(.din(n2069), .dout(n2070));
  jor  g02007(.dina(n2070), .dinb(n2068), .dout(n2071));
  jand g02008(.dina(n2071), .dinb(n2063), .dout(n2072));
  jxor g02009(.dina(n2057), .dinb(n1954), .dout(n2073));
  jnot g02010(.din(n2073), .dout(n2074));
  jor  g02011(.dina(n2074), .dinb(n2072), .dout(n2075));
  jand g02012(.dina(n2075), .dinb(n2060), .dout(n2076));
  jand g02013(.dina(n1903), .dinb(n884), .dout(n2077));
  jand g02014(.dina(n1470), .dinb(n1042), .dout(n2078));
  jand g02015(.dina(n2078), .dinb(n1352), .dout(n2079));
  jand g02016(.dina(n1246), .dinb(n501), .dout(n2080));
  jand g02017(.dina(n1334), .dinb(n991), .dout(n2081));
  jand g02018(.dina(n2081), .dinb(n2080), .dout(n2082));
  jand g02019(.dina(n1159), .dinb(n266), .dout(n2083));
  jand g02020(.dina(n2083), .dinb(n1218), .dout(n2084));
  jand g02021(.dina(n2084), .dinb(n2082), .dout(n2085));
  jand g02022(.dina(n886), .dinb(n1465), .dout(n2086));
  jand g02023(.dina(n516), .dinb(n639), .dout(n2087));
  jand g02024(.dina(n2087), .dinb(n2086), .dout(n2088));
  jand g02025(.dina(n630), .dinb(n175), .dout(n2089));
  jand g02026(.dina(n2089), .dinb(n2088), .dout(n2090));
  jand g02027(.dina(n2090), .dinb(n2085), .dout(n2091));
  jand g02028(.dina(n2091), .dinb(n2079), .dout(n2092));
  jand g02029(.dina(n1721), .dinb(n1316), .dout(n2093));
  jand g02030(.dina(n2093), .dinb(n988), .dout(n2094));
  jand g02031(.dina(n2094), .dinb(n638), .dout(n2095));
  jand g02032(.dina(n1212), .dinb(n1708), .dout(n2096));
  jand g02033(.dina(n2096), .dinb(n917), .dout(n2097));
  jand g02034(.dina(n1768), .dinb(n1580), .dout(n2098));
  jand g02035(.dina(n212), .dinb(n209), .dout(n2099));
  jnot g02036(.din(n2099), .dout(n2100));
  jand g02037(.dina(n2100), .dinb(n680), .dout(n2101));
  jand g02038(.dina(n2101), .dinb(n1713), .dout(n2102));
  jand g02039(.dina(n2102), .dinb(n2098), .dout(n2103));
  jand g02040(.dina(n2103), .dinb(n2097), .dout(n2104));
  jand g02041(.dina(n2104), .dinb(n2095), .dout(n2105));
  jand g02042(.dina(n1506), .dinb(n645), .dout(n2106));
  jand g02043(.dina(n1976), .dinb(n1326), .dout(n2107));
  jand g02044(.dina(n2107), .dinb(n1923), .dout(n2108));
  jand g02045(.dina(n2108), .dinb(n2106), .dout(n2109));
  jand g02046(.dina(n925), .dinb(n700), .dout(n2110));
  jand g02047(.dina(n2110), .dinb(n929), .dout(n2111));
  jand g02048(.dina(n2111), .dinb(n2109), .dout(n2112));
  jand g02049(.dina(n2112), .dinb(n2105), .dout(n2113));
  jand g02050(.dina(n2113), .dinb(n2092), .dout(n2114));
  jand g02051(.dina(n2114), .dinb(n600), .dout(n2115));
  jand g02052(.dina(n2115), .dinb(n2077), .dout(n2116));
  jnot g02053(.din(n255), .dout(n2117));
  jand g02054(.dina(n882), .dinb(n2117), .dout(n2118));
  jand g02055(.dina(n993), .dinb(n450), .dout(n2119));
  jand g02056(.dina(n1772), .dinb(n1273), .dout(n2120));
  jand g02057(.dina(n2120), .dinb(n1489), .dout(n2121));
  jand g02058(.dina(n2121), .dinb(n2119), .dout(n2122));
  jand g02059(.dina(n2122), .dinb(n2118), .dout(n2123));
  jnot g02060(.din(n857), .dout(n2124));
  jand g02061(.dina(n2124), .dinb(n472), .dout(n2125));
  jand g02062(.dina(n1309), .dinb(n933), .dout(n2126));
  jand g02063(.dina(n2126), .dinb(n2125), .dout(n2127));
  jand g02064(.dina(n1107), .dinb(n1756), .dout(n2128));
  jand g02065(.dina(n2128), .dinb(n714), .dout(n2129));
  jand g02066(.dina(n2129), .dinb(n2127), .dout(n2130));
  jand g02067(.dina(n1534), .dinb(n121), .dout(n2131));
  jand g02068(.dina(n2131), .dinb(n442), .dout(n2132));
  jand g02069(.dina(n2132), .dinb(n2130), .dout(n2133));
  jand g02070(.dina(n2133), .dinb(n2123), .dout(n2134));
  jand g02071(.dina(n660), .dinb(n818), .dout(n2135));
  jand g02072(.dina(n553), .dinb(n829), .dout(n2136));
  jand g02073(.dina(n2136), .dinb(n2135), .dout(n2137));
  jand g02074(.dina(n2137), .dinb(n1862), .dout(n2138));
  jand g02075(.dina(n2138), .dinb(n1260), .dout(n2139));
  jand g02076(.dina(n2139), .dinb(n1189), .dout(n2140));
  jand g02077(.dina(n2140), .dinb(n2134), .dout(n2141));
  jand g02078(.dina(n1473), .dinb(n499), .dout(n2142));
  jand g02079(.dina(n2142), .dinb(n447), .dout(n2143));
  jand g02080(.dina(n2143), .dinb(n869), .dout(n2144));
  jand g02081(.dina(n1516), .dinb(n920), .dout(n2145));
  jand g02082(.dina(n2145), .dinb(n1702), .dout(n2146));
  jand g02083(.dina(n2146), .dinb(n2144), .dout(n2147));
  jnot g02084(.din(n566), .dout(n2148));
  jand g02085(.dina(n1536), .dinb(n2148), .dout(n2149));
  jand g02086(.dina(n2149), .dinb(n809), .dout(n2150));
  jand g02087(.dina(n2150), .dinb(n827), .dout(n2151));
  jand g02088(.dina(n557), .dinb(n1360), .dout(n2152));
  jand g02089(.dina(n2152), .dinb(n2151), .dout(n2153));
  jand g02090(.dina(n647), .dinb(n907), .dout(n2154));
  jand g02091(.dina(n2154), .dinb(n1965), .dout(n2155));
  jand g02092(.dina(n2155), .dinb(n2153), .dout(n2156));
  jand g02093(.dina(n2156), .dinb(n2147), .dout(n2157));
  jand g02094(.dina(n1753), .dinb(n548), .dout(n2158));
  jand g02095(.dina(n2158), .dinb(n1427), .dout(n2159));
  jand g02096(.dina(n2159), .dinb(n1541), .dout(n2160));
  jand g02097(.dina(n1162), .dinb(n503), .dout(n2161));
  jand g02098(.dina(n452), .dinb(n916), .dout(n2162));
  jand g02099(.dina(n2162), .dinb(n135), .dout(n2163));
  jand g02100(.dina(n2163), .dinb(n2161), .dout(n2164));
  jand g02101(.dina(n1577), .dinb(n1453), .dout(n2165));
  jand g02102(.dina(n672), .dinb(n325), .dout(n2166));
  jand g02103(.dina(n2166), .dinb(n2165), .dout(n2167));
  jand g02104(.dina(n2167), .dinb(n1438), .dout(n2168));
  jand g02105(.dina(n2168), .dinb(n588), .dout(n2169));
  jand g02106(.dina(n2169), .dinb(n2164), .dout(n2170));
  jand g02107(.dina(n2170), .dinb(n2160), .dout(n2171));
  jand g02108(.dina(n2171), .dinb(n2157), .dout(n2172));
  jand g02109(.dina(n2172), .dinb(n2141), .dout(n2173));
  jand g02110(.dina(n2173), .dinb(n2116), .dout(n2174));
  jxor g02111(.dina(n2174), .dinb(n1954), .dout(n2175));
  jxor g02112(.dina(n2175), .dinb(n2076), .dout(n2176));
  jor  g02113(.dina(n2176), .dinb(n1820), .dout(n2177));
  jnot g02114(.din(n1817), .dout(n2178));
  jxor g02115(.dina(\a[19] ), .dinb(\a[18] ), .dout(n2179));
  jand g02116(.dina(n2179), .dinb(n2178), .dout(n2180));
  jnot g02117(.din(n2180), .dout(n2181));
  jor  g02118(.dina(n2181), .dinb(n1954), .dout(n2182));
  jor  g02119(.dina(n2179), .dinb(n1817), .dout(n2183));
  jnot g02120(.din(n2183), .dout(n2184));
  jand g02121(.dina(n2184), .dinb(n1818), .dout(n2185));
  jnot g02122(.din(n2185), .dout(n2186));
  jor  g02123(.dina(n2186), .dinb(n2057), .dout(n2187));
  jand g02124(.dina(n2187), .dinb(n2182), .dout(n2188));
  jor  g02125(.dina(n1818), .dinb(n2178), .dout(n2189));
  jor  g02126(.dina(n2189), .dinb(n2174), .dout(n2190));
  jand g02127(.dina(n2190), .dinb(n2188), .dout(n2191));
  jand g02128(.dina(n2191), .dinb(n2177), .dout(n2192));
  jxor g02129(.dina(n2192), .dinb(\a[20] ), .dout(n2193));
  jor  g02130(.dina(n2193), .dinb(n1816), .dout(n2194));
  jxor g02131(.dina(n1668), .dinb(n1667), .dout(n2195));
  jnot g02132(.din(\a[20] ), .dout(n2196));
  jxor g02133(.dina(n2073), .dinb(n2072), .dout(n2197));
  jor  g02134(.dina(n2197), .dinb(n1820), .dout(n2198));
  jor  g02135(.dina(n2186), .dinb(n1790), .dout(n2199));
  jor  g02136(.dina(n2189), .dinb(n1954), .dout(n2200));
  jor  g02137(.dina(n2181), .dinb(n2057), .dout(n2201));
  jand g02138(.dina(n2201), .dinb(n2200), .dout(n2202));
  jand g02139(.dina(n2202), .dinb(n2199), .dout(n2203));
  jand g02140(.dina(n2203), .dinb(n2198), .dout(n2204));
  jxor g02141(.dina(n2204), .dinb(n2196), .dout(n2205));
  jand g02142(.dina(n2205), .dinb(n2195), .dout(n2206));
  jxor g02143(.dina(n1664), .dinb(n1653), .dout(n2207));
  jxor g02144(.dina(n2069), .dinb(n2068), .dout(n2208));
  jor  g02145(.dina(n2208), .dinb(n1820), .dout(n2209));
  jor  g02146(.dina(n2181), .dinb(n1790), .dout(n2210));
  jor  g02147(.dina(n2186), .dinb(n1606), .dout(n2211));
  jor  g02148(.dina(n2189), .dinb(n2057), .dout(n2212));
  jand g02149(.dina(n2212), .dinb(n2211), .dout(n2213));
  jand g02150(.dina(n2213), .dinb(n2210), .dout(n2214));
  jand g02151(.dina(n2214), .dinb(n2209), .dout(n2215));
  jxor g02152(.dina(n2215), .dinb(n2196), .dout(n2216));
  jand g02153(.dina(n2216), .dinb(n2207), .dout(n2217));
  jor  g02154(.dina(n1820), .dinb(n1792), .dout(n2218));
  jor  g02155(.dina(n2189), .dinb(n1790), .dout(n2219));
  jor  g02156(.dina(n2186), .dinb(n1448), .dout(n2220));
  jor  g02157(.dina(n2181), .dinb(n1606), .dout(n2221));
  jand g02158(.dina(n2221), .dinb(n2220), .dout(n2222));
  jand g02159(.dina(n2222), .dinb(n2219), .dout(n2223));
  jand g02160(.dina(n2223), .dinb(n2218), .dout(n2224));
  jxor g02161(.dina(n2224), .dinb(n2196), .dout(n2225));
  jor  g02162(.dina(n1636), .dinb(n65), .dout(n2226));
  jxor g02163(.dina(n2226), .dinb(n1648), .dout(n2227));
  jand g02164(.dina(n2227), .dinb(n2225), .dout(n2228));
  jand g02165(.dina(n1633), .dinb(\a[23] ), .dout(n2229));
  jxor g02166(.dina(n2229), .dinb(n1631), .dout(n2230));
  jnot g02167(.din(n2230), .dout(n2231));
  jor  g02168(.dina(n1820), .dinb(n1608), .dout(n2232));
  jor  g02169(.dina(n2181), .dinb(n1448), .dout(n2233));
  jor  g02170(.dina(n2186), .dinb(n1255), .dout(n2234));
  jand g02171(.dina(n2234), .dinb(n2233), .dout(n2235));
  jor  g02172(.dina(n2189), .dinb(n1606), .dout(n2236));
  jand g02173(.dina(n2236), .dinb(n2235), .dout(n2237));
  jand g02174(.dina(n2237), .dinb(n2232), .dout(n2238));
  jxor g02175(.dina(n2238), .dinb(\a[20] ), .dout(n2239));
  jor  g02176(.dina(n2239), .dinb(n2231), .dout(n2240));
  jand g02177(.dina(n1819), .dinb(n728), .dout(n2241));
  jand g02178(.dina(n2180), .dinb(n438), .dout(n2242));
  jnot g02179(.din(n2189), .dout(n2243));
  jand g02180(.dina(n2243), .dinb(n795), .dout(n2244));
  jor  g02181(.dina(n2244), .dinb(n2242), .dout(n2245));
  jor  g02182(.dina(n2245), .dinb(n2241), .dout(n2246));
  jnot g02183(.din(n2246), .dout(n2247));
  jand g02184(.dina(n1817), .dinb(n438), .dout(n2248));
  jnot g02185(.din(n2248), .dout(n2249));
  jand g02186(.dina(n2249), .dinb(\a[20] ), .dout(n2250));
  jand g02187(.dina(n2250), .dinb(n2247), .dout(n2251));
  jand g02188(.dina(n1819), .dinb(n1639), .dout(n2252));
  jand g02189(.dina(n2180), .dinb(n795), .dout(n2253));
  jand g02190(.dina(n2243), .dinb(n1175), .dout(n2254));
  jor  g02191(.dina(n2254), .dinb(n2253), .dout(n2255));
  jand g02192(.dina(n2185), .dinb(n438), .dout(n2256));
  jor  g02193(.dina(n2256), .dinb(n2255), .dout(n2257));
  jor  g02194(.dina(n2257), .dinb(n2252), .dout(n2258));
  jnot g02195(.din(n2258), .dout(n2259));
  jand g02196(.dina(n2259), .dinb(n2251), .dout(n2260));
  jand g02197(.dina(n2260), .dinb(n1633), .dout(n2261));
  jnot g02198(.din(n2261), .dout(n2262));
  jxor g02199(.dina(n2260), .dinb(n1633), .dout(n2263));
  jnot g02200(.din(n2263), .dout(n2264));
  jor  g02201(.dina(n1820), .dinb(n1656), .dout(n2265));
  jor  g02202(.dina(n2186), .dinb(n726), .dout(n2266));
  jor  g02203(.dina(n2181), .dinb(n1255), .dout(n2267));
  jand g02204(.dina(n2267), .dinb(n2266), .dout(n2268));
  jor  g02205(.dina(n2189), .dinb(n1448), .dout(n2269));
  jand g02206(.dina(n2269), .dinb(n2268), .dout(n2270));
  jand g02207(.dina(n2270), .dinb(n2265), .dout(n2271));
  jxor g02208(.dina(n2271), .dinb(\a[20] ), .dout(n2272));
  jor  g02209(.dina(n2272), .dinb(n2264), .dout(n2273));
  jand g02210(.dina(n2273), .dinb(n2262), .dout(n2274));
  jnot g02211(.din(n2274), .dout(n2275));
  jxor g02212(.dina(n2239), .dinb(n2231), .dout(n2276));
  jand g02213(.dina(n2276), .dinb(n2275), .dout(n2277));
  jnot g02214(.din(n2277), .dout(n2278));
  jand g02215(.dina(n2278), .dinb(n2240), .dout(n2279));
  jnot g02216(.din(n2279), .dout(n2280));
  jxor g02217(.dina(n2227), .dinb(n2225), .dout(n2281));
  jand g02218(.dina(n2281), .dinb(n2280), .dout(n2282));
  jor  g02219(.dina(n2282), .dinb(n2228), .dout(n2283));
  jxor g02220(.dina(n2216), .dinb(n2207), .dout(n2284));
  jand g02221(.dina(n2284), .dinb(n2283), .dout(n2285));
  jor  g02222(.dina(n2285), .dinb(n2217), .dout(n2286));
  jxor g02223(.dina(n2205), .dinb(n2195), .dout(n2287));
  jand g02224(.dina(n2287), .dinb(n2286), .dout(n2288));
  jor  g02225(.dina(n2288), .dinb(n2206), .dout(n2289));
  jxor g02226(.dina(n2193), .dinb(n1816), .dout(n2290));
  jand g02227(.dina(n2290), .dinb(n2289), .dout(n2291));
  jnot g02228(.din(n2291), .dout(n2292));
  jand g02229(.dina(n2292), .dinb(n2194), .dout(n2293));
  jnot g02230(.din(n2293), .dout(n2294));
  jand g02231(.dina(n1813), .dinb(n1800), .dout(n2295));
  jand g02232(.dina(n1814), .dinb(n1672), .dout(n2296));
  jor  g02233(.dina(n2296), .dinb(n2295), .dout(n2297));
  jand g02234(.dina(n438), .dinb(n64), .dout(n2298));
  jnot g02235(.din(n2298), .dout(n2299));
  jor  g02236(.dina(n1811), .dinb(n1809), .dout(n2300));
  jxor g02237(.dina(n2300), .dinb(n2299), .dout(n2301));
  jnot g02238(.din(n2301), .dout(n2302));
  jnot g02239(.din(n71), .dout(n2303));
  jor  g02240(.dina(n1656), .dinb(n2303), .dout(n2304));
  jor  g02241(.dina(n1805), .dinb(n726), .dout(n2305));
  jnot g02242(.din(n731), .dout(n2306));
  jor  g02243(.dina(n1255), .dinb(n2306), .dout(n2307));
  jand g02244(.dina(n2307), .dinb(n2305), .dout(n2308));
  jnot g02245(.din(n796), .dout(n2309));
  jor  g02246(.dina(n1448), .dinb(n2309), .dout(n2310));
  jand g02247(.dina(n2310), .dinb(n2308), .dout(n2311));
  jand g02248(.dina(n2311), .dinb(n2304), .dout(n2312));
  jxor g02249(.dina(n2312), .dinb(\a[26] ), .dout(n2313));
  jxor g02250(.dina(n2313), .dinb(n2302), .dout(n2314));
  jor  g02251(.dina(n2208), .dinb(n807), .dout(n2315));
  jor  g02252(.dina(n1790), .dinb(n1613), .dout(n2316));
  jor  g02253(.dina(n1617), .dinb(n1606), .dout(n2317));
  jor  g02254(.dina(n2057), .dinb(n1621), .dout(n2318));
  jand g02255(.dina(n2318), .dinb(n2317), .dout(n2319));
  jand g02256(.dina(n2319), .dinb(n2316), .dout(n2320));
  jand g02257(.dina(n2320), .dinb(n2315), .dout(n2321));
  jxor g02258(.dina(n2321), .dinb(n65), .dout(n2322));
  jxor g02259(.dina(n2322), .dinb(n2314), .dout(n2323));
  jxor g02260(.dina(n2323), .dinb(n2297), .dout(n2324));
  jnot g02261(.din(n2174), .dout(n2325));
  jand g02262(.dina(n2325), .dinb(n1955), .dout(n2326));
  jnot g02263(.din(n2326), .dout(n2327));
  jnot g02264(.din(n2175), .dout(n2328));
  jor  g02265(.dina(n2328), .dinb(n2076), .dout(n2329));
  jand g02266(.dina(n2329), .dinb(n2327), .dout(n2330));
  jand g02267(.dina(n1346), .dinb(n1575), .dout(n2331));
  jand g02268(.dina(n2331), .dinb(n1327), .dout(n2332));
  jand g02269(.dina(n510), .dinb(n1203), .dout(n2333));
  jand g02270(.dina(n2333), .dinb(n2052), .dout(n2334));
  jand g02271(.dina(n2100), .dinb(n1005), .dout(n2335));
  jand g02272(.dina(n2335), .dinb(n1090), .dout(n2336));
  jand g02273(.dina(n2336), .dinb(n2334), .dout(n2337));
  jand g02274(.dina(n1961), .dinb(n537), .dout(n2338));
  jand g02275(.dina(n2338), .dinb(n583), .dout(n2339));
  jand g02276(.dina(n2339), .dinb(n2337), .dout(n2340));
  jand g02277(.dina(n1495), .dinb(n101), .dout(n2341));
  jand g02278(.dina(n2341), .dinb(n685), .dout(n2342));
  jand g02279(.dina(n660), .dinb(n1305), .dout(n2343));
  jand g02280(.dina(n1524), .dinb(n175), .dout(n2344));
  jand g02281(.dina(n2344), .dinb(n270), .dout(n2345));
  jand g02282(.dina(n2345), .dinb(n2343), .dout(n2346));
  jand g02283(.dina(n2346), .dinb(n2342), .dout(n2347));
  jand g02284(.dina(n2347), .dinb(n2340), .dout(n2348));
  jand g02285(.dina(n2348), .dinb(n2332), .dout(n2349));
  jand g02286(.dina(n1324), .dinb(n676), .dout(n2350));
  jand g02287(.dina(n2350), .dinb(n932), .dout(n2351));
  jand g02288(.dina(n1361), .dinb(n880), .dout(n2352));
  jand g02289(.dina(n2352), .dinb(n2351), .dout(n2353));
  jand g02290(.dina(n2353), .dinb(n1691), .dout(n2354));
  jand g02291(.dina(n2354), .dinb(n551), .dout(n2355));
  jand g02292(.dina(n2355), .dinb(n2349), .dout(n2356));
  jand g02293(.dina(n461), .dinb(n266), .dout(n2357));
  jand g02294(.dina(n965), .dinb(n452), .dout(n2358));
  jand g02295(.dina(n668), .dinb(n1822), .dout(n2359));
  jand g02296(.dina(n2359), .dinb(n2358), .dout(n2360));
  jand g02297(.dina(n1846), .dinb(n1212), .dout(n2361));
  jand g02298(.dina(n907), .dinb(n1226), .dout(n2362));
  jand g02299(.dina(n2362), .dinb(n2361), .dout(n2363));
  jand g02300(.dina(n2363), .dinb(n2360), .dout(n2364));
  jand g02301(.dina(n2364), .dinb(n2357), .dout(n2365));
  jand g02302(.dina(n511), .dinb(n695), .dout(n2366));
  jand g02303(.dina(n470), .dinb(n130), .dout(n2367));
  jand g02304(.dina(n2367), .dinb(n2366), .dout(n2368));
  jand g02305(.dina(n2368), .dinb(n887), .dout(n2369));
  jand g02306(.dina(n2369), .dinb(n1698), .dout(n2370));
  jand g02307(.dina(n2370), .dinb(n2365), .dout(n2371));
  jand g02308(.dina(n1541), .dinb(n1569), .dout(n2372));
  jand g02309(.dina(n672), .dinb(n328), .dout(n2373));
  jand g02310(.dina(n2373), .dinb(n2087), .dout(n2374));
  jand g02311(.dina(n2374), .dinb(n2372), .dout(n2375));
  jand g02312(.dina(n1360), .dinb(n1344), .dout(n2376));
  jand g02313(.dina(n2376), .dinb(n2117), .dout(n2377));
  jand g02314(.dina(n833), .dinb(n1534), .dout(n2378));
  jand g02315(.dina(n1345), .dinb(n1233), .dout(n2379));
  jand g02316(.dina(n2379), .dinb(n2378), .dout(n2380));
  jand g02317(.dina(n2380), .dinb(n1429), .dout(n2381));
  jand g02318(.dina(n2381), .dinb(n2377), .dout(n2382));
  jand g02319(.dina(n2382), .dinb(n2375), .dout(n2383));
  jand g02320(.dina(n2383), .dinb(n2371), .dout(n2384));
  jand g02321(.dina(n808), .dinb(n1270), .dout(n2385));
  jand g02322(.dina(n1246), .dinb(n650), .dout(n2386));
  jand g02323(.dina(n2386), .dinb(n2385), .dout(n2387));
  jand g02324(.dina(n2387), .dinb(n2023), .dout(n2388));
  jand g02325(.dina(n2388), .dinb(n681), .dout(n2389));
  jand g02326(.dina(n1317), .dinb(n121), .dout(n2390));
  jand g02327(.dina(n2390), .dinb(n2389), .dout(n2391));
  jand g02328(.dina(n2391), .dinb(n2384), .dout(n2392));
  jand g02329(.dina(n1971), .dinb(n831), .dout(n2393));
  jand g02330(.dina(n168), .dinb(n501), .dout(n2394));
  jand g02331(.dina(n411), .dinb(n108), .dout(n2395));
  jand g02332(.dina(n2395), .dinb(n2394), .dout(n2396));
  jand g02333(.dina(n2396), .dinb(n2393), .dout(n2397));
  jand g02334(.dina(n2397), .dinb(n703), .dout(n2398));
  jand g02335(.dina(n1968), .dinb(n1190), .dout(n2399));
  jand g02336(.dina(n2124), .dinb(n555), .dout(n2400));
  jand g02337(.dina(n1708), .dinb(n1304), .dout(n2401));
  jand g02338(.dina(n2401), .dinb(n2400), .dout(n2402));
  jand g02339(.dina(n2402), .dinb(n2399), .dout(n2403));
  jand g02340(.dina(n2403), .dinb(n1934), .dout(n2404));
  jand g02341(.dina(n2404), .dinb(n2398), .dout(n2405));
  jand g02342(.dina(n1743), .dinb(n1219), .dout(n2406));
  jand g02343(.dina(n553), .dinb(n481), .dout(n2407));
  jand g02344(.dina(n2407), .dinb(n2406), .dout(n2408));
  jand g02345(.dina(n562), .dinb(n1088), .dout(n2409));
  jand g02346(.dina(n2409), .dinb(n1753), .dout(n2410));
  jand g02347(.dina(n2410), .dinb(n983), .dout(n2411));
  jand g02348(.dina(n2411), .dinb(n2408), .dout(n2412));
  jand g02349(.dina(n981), .dinb(n454), .dout(n2413));
  jand g02350(.dina(n893), .dinb(n178), .dout(n2414));
  jand g02351(.dina(n2414), .dinb(n2413), .dout(n2415));
  jand g02352(.dina(n1437), .dinb(n541), .dout(n2416));
  jand g02353(.dina(n2416), .dinb(n132), .dout(n2417));
  jand g02354(.dina(n2417), .dinb(n2415), .dout(n2418));
  jand g02355(.dina(n492), .dinb(n653), .dout(n2419));
  jand g02356(.dina(n1536), .dinb(n696), .dout(n2420));
  jand g02357(.dina(n1159), .dinb(n1309), .dout(n2421));
  jand g02358(.dina(n2421), .dinb(n2420), .dout(n2422));
  jand g02359(.dina(n2422), .dinb(n2419), .dout(n2423));
  jand g02360(.dina(n2423), .dinb(n2418), .dout(n2424));
  jand g02361(.dina(n2424), .dinb(n2412), .dout(n2425));
  jand g02362(.dina(n2425), .dinb(n2405), .dout(n2426));
  jand g02363(.dina(n2426), .dinb(n2392), .dout(n2427));
  jand g02364(.dina(n2427), .dinb(n2356), .dout(n2428));
  jxor g02365(.dina(n2428), .dinb(n2174), .dout(n2429));
  jxor g02366(.dina(n2429), .dinb(n2330), .dout(n2430));
  jor  g02367(.dina(n2430), .dinb(n1820), .dout(n2431));
  jor  g02368(.dina(n2181), .dinb(n2174), .dout(n2432));
  jor  g02369(.dina(n2428), .dinb(n2189), .dout(n2433));
  jor  g02370(.dina(n2186), .dinb(n1954), .dout(n2434));
  jand g02371(.dina(n2434), .dinb(n2433), .dout(n2435));
  jand g02372(.dina(n2435), .dinb(n2432), .dout(n2436));
  jand g02373(.dina(n2436), .dinb(n2431), .dout(n2437));
  jxor g02374(.dina(n2437), .dinb(n2196), .dout(n2438));
  jxor g02375(.dina(n2438), .dinb(n2324), .dout(n2439));
  jxor g02376(.dina(n2439), .dinb(n2294), .dout(n2440));
  jnot g02377(.din(\a[17] ), .dout(n2441));
  jand g02378(.dina(n351), .dinb(n100), .dout(n2442));
  jand g02379(.dina(n2442), .dinb(n1096), .dout(n2443));
  jand g02380(.dina(n1846), .dinb(n654), .dout(n2444));
  jand g02381(.dina(n886), .dinb(n501), .dout(n2445));
  jand g02382(.dina(n2445), .dinb(n2444), .dout(n2446));
  jand g02383(.dina(n2446), .dinb(n2443), .dout(n2447));
  jand g02384(.dina(n588), .dinb(n516), .dout(n2448));
  jand g02385(.dina(n2448), .dinb(n700), .dout(n2449));
  jand g02386(.dina(n1697), .dinb(n108), .dout(n2450));
  jand g02387(.dina(n2450), .dinb(n2449), .dout(n2451));
  jand g02388(.dina(n2451), .dinb(n2447), .dout(n2452));
  jand g02389(.dina(n2452), .dinb(n1438), .dout(n2453));
  jand g02390(.dina(n328), .dinb(n900), .dout(n2454));
  jand g02391(.dina(n931), .dinb(n873), .dout(n2455));
  jand g02392(.dina(n1349), .dinb(n469), .dout(n2456));
  jand g02393(.dina(n2456), .dinb(n2455), .dout(n2457));
  jand g02394(.dina(n1360), .dinb(n541), .dout(n2458));
  jand g02395(.dina(n2458), .dinb(n326), .dout(n2459));
  jand g02396(.dina(n2459), .dinb(n2457), .dout(n2460));
  jand g02397(.dina(n2460), .dinb(n2454), .dout(n2461));
  jand g02398(.dina(n826), .dinb(n818), .dout(n2462));
  jand g02399(.dina(n1219), .dinb(n621), .dout(n2463));
  jand g02400(.dina(n2463), .dinb(n1473), .dout(n2464));
  jand g02401(.dina(n2464), .dinb(n2462), .dout(n2465));
  jand g02402(.dina(n1961), .dinb(n1708), .dout(n2466));
  jand g02403(.dina(n2466), .dinb(n1168), .dout(n2467));
  jand g02404(.dina(n2467), .dinb(n2465), .dout(n2468));
  jand g02405(.dina(n2468), .dinb(n1189), .dout(n2469));
  jand g02406(.dina(n2469), .dinb(n2461), .dout(n2470));
  jand g02407(.dina(n2470), .dinb(n2453), .dout(n2471));
  jand g02408(.dina(n1037), .dinb(n1213), .dout(n2472));
  jand g02409(.dina(n2472), .dinb(n2471), .dout(n2473));
  jand g02410(.dina(n981), .dinb(n411), .dout(n2474));
  jand g02411(.dina(n2474), .dinb(n1843), .dout(n2475));
  jand g02412(.dina(n2475), .dinb(n1822), .dout(n2476));
  jand g02413(.dina(n1451), .dinb(n442), .dout(n2477));
  jand g02414(.dina(n2477), .dinb(n917), .dout(n2478));
  jand g02415(.dina(n1534), .dinb(n430), .dout(n2479));
  jand g02416(.dina(n2479), .dinb(n82), .dout(n2480));
  jand g02417(.dina(n2480), .dinb(n2478), .dout(n2481));
  jand g02418(.dina(n1352), .dinb(n1345), .dout(n2482));
  jand g02419(.dina(n547), .dinb(n1375), .dout(n2483));
  jand g02420(.dina(n2483), .dinb(n1569), .dout(n2484));
  jand g02421(.dina(n2484), .dinb(n2482), .dout(n2485));
  jand g02422(.dina(n2485), .dinb(n2481), .dout(n2486));
  jand g02423(.dina(n2486), .dinb(n2476), .dout(n2487));
  jand g02424(.dina(n1017), .dinb(n716), .dout(n2488));
  jand g02425(.dina(n2488), .dinb(n1898), .dout(n2489));
  jand g02426(.dina(n893), .dinb(n1575), .dout(n2490));
  jand g02427(.dina(n2490), .dinb(n685), .dout(n2491));
  jand g02428(.dina(n824), .dinb(n171), .dout(n2492));
  jand g02429(.dina(n2492), .dinb(n1107), .dout(n2493));
  jand g02430(.dina(n2493), .dinb(n1043), .dout(n2494));
  jand g02431(.dina(n2494), .dinb(n2491), .dout(n2495));
  jand g02432(.dina(n2495), .dinb(n2489), .dout(n2496));
  jand g02433(.dina(n2023), .dinb(n440), .dout(n2497));
  jand g02434(.dina(n534), .dinb(n1327), .dout(n2498));
  jand g02435(.dina(n2498), .dinb(n2497), .dout(n2499));
  jand g02436(.dina(n1053), .dinb(n178), .dout(n2500));
  jand g02437(.dina(n670), .dinb(n632), .dout(n2501));
  jand g02438(.dina(n2501), .dinb(n2500), .dout(n2502));
  jand g02439(.dina(n2502), .dinb(n2499), .dout(n2503));
  jand g02440(.dina(n1088), .dinb(n662), .dout(n2504));
  jand g02441(.dina(n2504), .dinb(n2503), .dout(n2505));
  jand g02442(.dina(n2505), .dinb(n2496), .dout(n2506));
  jand g02443(.dina(n2506), .dinb(n2487), .dout(n2507));
  jand g02444(.dina(n1495), .dinb(n1225), .dout(n2508));
  jand g02445(.dina(n2508), .dinb(n554), .dout(n2509));
  jand g02446(.dina(n2509), .dinb(n514), .dout(n2510));
  jnot g02447(.din(n488), .dout(n2511));
  jand g02448(.dina(n1515), .dinb(n600), .dout(n2512));
  jand g02449(.dina(n2512), .dinb(n562), .dout(n2513));
  jand g02450(.dina(n2513), .dinb(n2511), .dout(n2514));
  jand g02451(.dina(n2514), .dinb(n2510), .dout(n2515));
  jand g02452(.dina(n1721), .dinb(n1449), .dout(n2516));
  jand g02453(.dina(n2516), .dinb(n1205), .dout(n2517));
  jand g02454(.dina(n2517), .dinb(n1580), .dout(n2518));
  jand g02455(.dina(n2518), .dinb(n555), .dout(n2519));
  jand g02456(.dina(n2519), .dinb(n2515), .dout(n2520));
  jand g02457(.dina(n664), .dinb(n463), .dout(n2521));
  jand g02458(.dina(n1367), .dinb(n114), .dout(n2522));
  jand g02459(.dina(n2522), .dinb(n1324), .dout(n2523));
  jand g02460(.dina(n2523), .dinb(n1579), .dout(n2524));
  jand g02461(.dina(n2524), .dinb(n2521), .dout(n2525));
  jand g02462(.dina(n1090), .dinb(n510), .dout(n2526));
  jand g02463(.dina(n2526), .dinb(n1308), .dout(n2527));
  jand g02464(.dina(n2527), .dinb(n638), .dout(n2528));
  jand g02465(.dina(n1159), .dinb(n908), .dout(n2529));
  jand g02466(.dina(n2529), .dinb(n1373), .dout(n2530));
  jand g02467(.dina(n1237), .dinb(n1432), .dout(n2531));
  jand g02468(.dina(n2148), .dinb(n1305), .dout(n2532));
  jand g02469(.dina(n2532), .dinb(n2531), .dout(n2533));
  jand g02470(.dina(n2533), .dinb(n2530), .dout(n2534));
  jand g02471(.dina(n2534), .dinb(n2528), .dout(n2535));
  jand g02472(.dina(n2535), .dinb(n1380), .dout(n2536));
  jand g02473(.dina(n2536), .dinb(n2525), .dout(n2537));
  jand g02474(.dina(n884), .dinb(n1273), .dout(n2538));
  jand g02475(.dina(n2538), .dinb(n642), .dout(n2539));
  jand g02476(.dina(n1541), .dinb(n1344), .dout(n2540));
  jand g02477(.dina(n703), .dinb(n808), .dout(n2541));
  jand g02478(.dina(n978), .dinb(n933), .dout(n2542));
  jand g02479(.dina(n2542), .dinb(n2541), .dout(n2543));
  jand g02480(.dina(n869), .dinb(n428), .dout(n2544));
  jand g02481(.dina(n2544), .dinb(n517), .dout(n2545));
  jand g02482(.dina(n2545), .dinb(n2543), .dout(n2546));
  jand g02483(.dina(n2546), .dinb(n2540), .dout(n2547));
  jand g02484(.dina(n2547), .dinb(n1560), .dout(n2548));
  jand g02485(.dina(n2548), .dinb(n2539), .dout(n2549));
  jand g02486(.dina(n2549), .dinb(n2537), .dout(n2550));
  jand g02487(.dina(n2550), .dinb(n2520), .dout(n2551));
  jand g02488(.dina(n2551), .dinb(n2507), .dout(n2552));
  jand g02489(.dina(n2552), .dinb(n2473), .dout(n2553));
  jnot g02490(.din(n2553), .dout(n2554));
  jand g02491(.dina(n1237), .dinb(n480), .dout(n2555));
  jand g02492(.dina(n2555), .dinb(n1305), .dout(n2556));
  jand g02493(.dina(n2556), .dinb(n266), .dout(n2557));
  jand g02494(.dina(n2557), .dinb(n328), .dout(n2558));
  jand g02495(.dina(n694), .dinb(n411), .dout(n2559));
  jand g02496(.dina(n2559), .dinb(n1525), .dout(n2560));
  jand g02497(.dina(n1090), .dinb(n1569), .dout(n2561));
  jand g02498(.dina(n2561), .dinb(n1247), .dout(n2562));
  jand g02499(.dina(n2562), .dinb(n2560), .dout(n2563));
  jand g02500(.dina(n2563), .dinb(n554), .dout(n2564));
  jand g02501(.dina(n2564), .dinb(n2558), .dout(n2565));
  jand g02502(.dina(n950), .dinb(n534), .dout(n2566));
  jand g02503(.dina(n2566), .dinb(n1218), .dout(n2567));
  jand g02504(.dina(n1559), .dinb(n1205), .dout(n2568));
  jand g02505(.dina(n2568), .dinb(n2567), .dout(n2569));
  jnot g02506(.din(n1026), .dout(n2570));
  jand g02507(.dina(n900), .dinb(n1432), .dout(n2571));
  jand g02508(.dina(n2571), .dinb(n2570), .dout(n2572));
  jand g02509(.dina(n647), .dinb(n1376), .dout(n2573));
  jand g02510(.dina(n2573), .dinb(n2572), .dout(n2574));
  jand g02511(.dina(n2574), .dinb(n490), .dout(n2575));
  jand g02512(.dina(n2575), .dinb(n2569), .dout(n2576));
  jand g02513(.dina(n1361), .dinb(n325), .dout(n2577));
  jand g02514(.dina(n2577), .dinb(n1591), .dout(n2578));
  jand g02515(.dina(n2578), .dinb(n672), .dout(n2579));
  jand g02516(.dina(n1778), .dinb(n481), .dout(n2580));
  jand g02517(.dina(n917), .dinb(n954), .dout(n2581));
  jand g02518(.dina(n2581), .dinb(n2580), .dout(n2582));
  jand g02519(.dina(n2409), .dinb(n654), .dout(n2583));
  jand g02520(.dina(n2583), .dinb(n2582), .dout(n2584));
  jand g02521(.dina(n2584), .dinb(n2579), .dout(n2585));
  jand g02522(.dina(n1189), .dinb(n1238), .dout(n2586));
  jand g02523(.dina(n988), .dinb(n469), .dout(n2587));
  jand g02524(.dina(n600), .dinb(n1273), .dout(n2588));
  jand g02525(.dina(n2588), .dinb(n2587), .dout(n2589));
  jand g02526(.dina(n2589), .dinb(n2586), .dout(n2590));
  jand g02527(.dina(n2590), .dinb(n2079), .dout(n2591));
  jand g02528(.dina(n2591), .dinb(n1438), .dout(n2592));
  jand g02529(.dina(n2592), .dinb(n2585), .dout(n2593));
  jand g02530(.dina(n2593), .dinb(n2576), .dout(n2594));
  jand g02531(.dina(n886), .dinb(n824), .dout(n2595));
  jand g02532(.dina(n2595), .dinb(n2390), .dout(n2596));
  jand g02533(.dina(n685), .dinb(n135), .dout(n2597));
  jand g02534(.dina(n2597), .dinb(n1903), .dout(n2598));
  jand g02535(.dina(n2598), .dinb(n2596), .dout(n2599));
  jand g02536(.dina(n1053), .dinb(n1310), .dout(n2600));
  jand g02537(.dina(n548), .dinb(n893), .dout(n2601));
  jand g02538(.dina(n2601), .dinb(n452), .dout(n2602));
  jand g02539(.dina(n2602), .dinb(n2600), .dout(n2603));
  jand g02540(.dina(n2603), .dinb(n2599), .dout(n2604));
  jand g02541(.dina(n695), .dinb(n1245), .dout(n2605));
  jand g02542(.dina(n2605), .dinb(n1349), .dout(n2606));
  jand g02543(.dina(n2606), .dinb(n1283), .dout(n2607));
  jand g02544(.dina(n1367), .dinb(n450), .dout(n2608));
  jand g02545(.dina(n2608), .dinb(n848), .dout(n2609));
  jand g02546(.dina(n2609), .dinb(n2607), .dout(n2610));
  jand g02547(.dina(n2610), .dinb(n2604), .dout(n2611));
  jand g02548(.dina(n1188), .dinb(n582), .dout(n2612));
  jand g02549(.dina(n2612), .dinb(n2333), .dout(n2613));
  jand g02550(.dina(n1096), .dinb(n492), .dout(n2614));
  jand g02551(.dina(n2614), .dinb(n1016), .dout(n2615));
  jand g02552(.dina(n2615), .dinb(n1207), .dout(n2616));
  jand g02553(.dina(n2616), .dinb(n2613), .dout(n2617));
  jand g02554(.dina(n1167), .dinb(n1225), .dout(n2618));
  jand g02555(.dina(n2618), .dinb(n1373), .dout(n2619));
  jand g02556(.dina(n1560), .dinb(n586), .dout(n2620));
  jand g02557(.dina(n2620), .dinb(n2619), .dout(n2621));
  jand g02558(.dina(n2012), .dinb(n1328), .dout(n2622));
  jand g02559(.dina(n2622), .dinb(n1506), .dout(n2623));
  jand g02560(.dina(n2623), .dinb(n2621), .dout(n2624));
  jand g02561(.dina(n2624), .dinb(n2617), .dout(n2625));
  jand g02562(.dina(n2625), .dinb(n2611), .dout(n2626));
  jand g02563(.dina(n2626), .dinb(n1728), .dout(n2627));
  jand g02564(.dina(n2627), .dinb(n2594), .dout(n2628));
  jand g02565(.dina(n2628), .dinb(n2565), .dout(n2629));
  jnot g02566(.din(n2629), .dout(n2630));
  jand g02567(.dina(n2630), .dinb(n2554), .dout(n2631));
  jnot g02568(.din(n2631), .dout(n2632));
  jnot g02569(.din(n2428), .dout(n2633));
  jand g02570(.dina(n2630), .dinb(n2633), .dout(n2634));
  jnot g02571(.din(n2634), .dout(n2635));
  jand g02572(.dina(n2633), .dinb(n2325), .dout(n2636));
  jnot g02573(.din(n2636), .dout(n2637));
  jnot g02574(.din(n2429), .dout(n2638));
  jor  g02575(.dina(n2638), .dinb(n2330), .dout(n2639));
  jand g02576(.dina(n2639), .dinb(n2637), .dout(n2640));
  jxor g02577(.dina(n2629), .dinb(n2428), .dout(n2641));
  jnot g02578(.din(n2641), .dout(n2642));
  jor  g02579(.dina(n2642), .dinb(n2640), .dout(n2643));
  jand g02580(.dina(n2643), .dinb(n2635), .dout(n2644));
  jxor g02581(.dina(n2629), .dinb(n2553), .dout(n2645));
  jnot g02582(.din(n2645), .dout(n2646));
  jor  g02583(.dina(n2646), .dinb(n2644), .dout(n2647));
  jand g02584(.dina(n2647), .dinb(n2632), .dout(n2648));
  jand g02585(.dina(n1721), .dinb(n1903), .dout(n2649));
  jand g02586(.dina(n2649), .dinb(n1470), .dout(n2650));
  jand g02587(.dina(n2650), .dinb(n848), .dout(n2651));
  jand g02588(.dina(n881), .dinb(n1366), .dout(n2652));
  jand g02589(.dina(n2652), .dinb(n2148), .dout(n2653));
  jand g02590(.dina(n2653), .dinb(n630), .dout(n2654));
  jand g02591(.dina(n2654), .dinb(n2651), .dout(n2655));
  jand g02592(.dina(n2655), .dinb(n908), .dout(n2656));
  jand g02593(.dina(n1534), .dinb(n1360), .dout(n2657));
  jand g02594(.dina(n2657), .dinb(n1310), .dout(n2658));
  jand g02595(.dina(n869), .dinb(n1238), .dout(n2659));
  jand g02596(.dina(n1532), .dinb(n664), .dout(n2660));
  jand g02597(.dina(n2660), .dinb(n2659), .dout(n2661));
  jand g02598(.dina(n2661), .dinb(n2658), .dout(n2662));
  jand g02599(.dina(n1476), .dinb(n1276), .dout(n2663));
  jand g02600(.dina(n2663), .dinb(n2106), .dout(n2664));
  jand g02601(.dina(n2664), .dinb(n2662), .dout(n2665));
  jand g02602(.dina(n1714), .dinb(n499), .dout(n2666));
  jand g02603(.dina(n1162), .dinb(n668), .dout(n2667));
  jand g02604(.dina(n2667), .dinb(n542), .dout(n2668));
  jand g02605(.dina(n2668), .dinb(n2666), .dout(n2669));
  jand g02606(.dina(n1700), .dinb(n511), .dout(n2670));
  jand g02607(.dina(n2670), .dinb(n2587), .dout(n2671));
  jand g02608(.dina(n2671), .dinb(n2669), .dout(n2672));
  jand g02609(.dina(n2672), .dinb(n2665), .dout(n2673));
  jand g02610(.dina(n351), .dinb(n1575), .dout(n2674));
  jand g02611(.dina(n2674), .dinb(n320), .dout(n2675));
  jand g02612(.dina(n2675), .dinb(n2122), .dout(n2676));
  jand g02613(.dina(n2676), .dinb(n1524), .dout(n2677));
  jand g02614(.dina(n2677), .dinb(n2673), .dout(n2678));
  jand g02615(.dina(n2678), .dinb(n2656), .dout(n2679));
  jand g02616(.dina(n632), .dinb(n893), .dout(n2680));
  jand g02617(.dina(n696), .dinb(n1317), .dout(n2681));
  jand g02618(.dina(n2681), .dinb(n2680), .dout(n2682));
  jand g02619(.dina(n2682), .dinb(n495), .dout(n2683));
  jand g02620(.dina(n833), .dinb(n553), .dout(n2684));
  jand g02621(.dina(n2684), .dinb(n699), .dout(n2685));
  jand g02622(.dina(n2685), .dinb(n2367), .dout(n2686));
  jand g02623(.dina(n2686), .dinb(n2683), .dout(n2687));
  jand g02624(.dina(n950), .dinb(n1778), .dout(n2688));
  jand g02625(.dina(n2688), .dinb(n447), .dout(n2689));
  jand g02626(.dina(n2689), .dinb(n2047), .dout(n2690));
  jand g02627(.dina(n2690), .dinb(n1709), .dout(n2691));
  jand g02628(.dina(n2691), .dinb(n2687), .dout(n2692));
  jand g02629(.dina(n1189), .dinb(n557), .dout(n2693));
  jand g02630(.dina(n1738), .dinb(n1822), .dout(n2694));
  jand g02631(.dina(n2694), .dinb(n2693), .dout(n2695));
  jand g02632(.dina(n2695), .dinb(n639), .dout(n2696));
  jand g02633(.dina(n2696), .dinb(n1246), .dout(n2697));
  jand g02634(.dina(n1867), .dinb(n838), .dout(n2698));
  jand g02635(.dina(n2698), .dinb(n1227), .dout(n2699));
  jand g02636(.dina(n873), .dinb(n503), .dout(n2700));
  jand g02637(.dina(n2700), .dinb(n660), .dout(n2701));
  jand g02638(.dina(n2701), .dinb(n2699), .dout(n2702));
  jand g02639(.dina(n2702), .dinb(n1347), .dout(n2703));
  jand g02640(.dina(n2703), .dinb(n2697), .dout(n2704));
  jand g02641(.dina(n1843), .dinb(n809), .dout(n2705));
  jand g02642(.dina(n2705), .dinb(n2704), .dout(n2706));
  jand g02643(.dina(n2706), .dinb(n2692), .dout(n2707));
  jand g02644(.dina(n1233), .dinb(n1430), .dout(n2708));
  jand g02645(.dina(n2708), .dinb(n456), .dout(n2709));
  jand g02646(.dina(n2101), .dinb(n887), .dout(n2710));
  jand g02647(.dina(n2710), .dinb(n2709), .dout(n2711));
  jand g02648(.dina(n2711), .dinb(n1516), .dout(n2712));
  jand g02649(.dina(n641), .dinb(n452), .dout(n2713));
  jand g02650(.dina(n2713), .dinb(n1834), .dout(n2714));
  jand g02651(.dina(n2714), .dinb(n1349), .dout(n2715));
  jand g02652(.dina(n547), .dinb(n516), .dout(n2716));
  jand g02653(.dina(n2716), .dinb(n551), .dout(n2717));
  jand g02654(.dina(n2717), .dinb(n2715), .dout(n2718));
  jand g02655(.dina(n2718), .dinb(n2712), .dout(n2719));
  jand g02656(.dina(n1098), .dinb(n178), .dout(n2720));
  jand g02657(.dina(n2720), .dinb(n1437), .dout(n2721));
  jand g02658(.dina(n463), .dinb(n1429), .dout(n2722));
  jand g02659(.dina(n2722), .dinb(n2721), .dout(n2723));
  jand g02660(.dina(n1504), .dinb(n535), .dout(n2724));
  jand g02661(.dina(n2724), .dinb(n2167), .dout(n2725));
  jand g02662(.dina(n2725), .dinb(n2723), .dout(n2726));
  jand g02663(.dina(n2619), .dinb(n2130), .dout(n2727));
  jand g02664(.dina(n2727), .dinb(n2726), .dout(n2728));
  jand g02665(.dina(n1159), .dinb(n582), .dout(n2729));
  jand g02666(.dina(n2729), .dinb(n121), .dout(n2730));
  jand g02667(.dina(n2730), .dinb(n2031), .dout(n2731));
  jand g02668(.dina(n1582), .dinb(n430), .dout(n2732));
  jand g02669(.dina(n2732), .dinb(n925), .dout(n2733));
  jand g02670(.dina(n2733), .dinb(n2731), .dout(n2734));
  jand g02671(.dina(n2734), .dinb(n2728), .dout(n2735));
  jand g02672(.dina(n2735), .dinb(n2719), .dout(n2736));
  jand g02673(.dina(n2736), .dinb(n2707), .dout(n2737));
  jand g02674(.dina(n2737), .dinb(n2679), .dout(n2738));
  jxor g02675(.dina(n2738), .dinb(n2553), .dout(n2739));
  jxor g02676(.dina(n2739), .dinb(n2648), .dout(n2740));
  jxor g02677(.dina(\a[15] ), .dinb(\a[14] ), .dout(n2741));
  jxor g02678(.dina(\a[17] ), .dinb(\a[16] ), .dout(n2742));
  jand g02679(.dina(n2742), .dinb(n2741), .dout(n2743));
  jnot g02680(.din(n2743), .dout(n2744));
  jor  g02681(.dina(n2744), .dinb(n2740), .dout(n2745));
  jnot g02682(.din(n2741), .dout(n2746));
  jxor g02683(.dina(\a[16] ), .dinb(\a[15] ), .dout(n2747));
  jand g02684(.dina(n2747), .dinb(n2746), .dout(n2748));
  jnot g02685(.din(n2748), .dout(n2749));
  jor  g02686(.dina(n2749), .dinb(n2553), .dout(n2750));
  jnot g02687(.din(n2742), .dout(n2751));
  jand g02688(.dina(n2751), .dinb(n2741), .dout(n2752));
  jnot g02689(.din(n2752), .dout(n2753));
  jor  g02690(.dina(n2753), .dinb(n2738), .dout(n2754));
  jor  g02691(.dina(n2747), .dinb(n2741), .dout(n2755));
  jnot g02692(.din(n2755), .dout(n2756));
  jand g02693(.dina(n2756), .dinb(n2742), .dout(n2757));
  jnot g02694(.din(n2757), .dout(n2758));
  jor  g02695(.dina(n2758), .dinb(n2629), .dout(n2759));
  jand g02696(.dina(n2759), .dinb(n2754), .dout(n2760));
  jand g02697(.dina(n2760), .dinb(n2750), .dout(n2761));
  jand g02698(.dina(n2761), .dinb(n2745), .dout(n2762));
  jxor g02699(.dina(n2762), .dinb(n2441), .dout(n2763));
  jand g02700(.dina(n2763), .dinb(n2440), .dout(n2764));
  jxor g02701(.dina(n2290), .dinb(n2289), .dout(n2765));
  jnot g02702(.din(n2765), .dout(n2766));
  jor  g02703(.dina(n2753), .dinb(n2553), .dout(n2767));
  jxor g02704(.dina(n2645), .dinb(n2644), .dout(n2768));
  jor  g02705(.dina(n2768), .dinb(n2744), .dout(n2769));
  jor  g02706(.dina(n2758), .dinb(n2428), .dout(n2770));
  jor  g02707(.dina(n2749), .dinb(n2629), .dout(n2771));
  jand g02708(.dina(n2771), .dinb(n2770), .dout(n2772));
  jand g02709(.dina(n2772), .dinb(n2769), .dout(n2773));
  jand g02710(.dina(n2773), .dinb(n2767), .dout(n2774));
  jxor g02711(.dina(n2774), .dinb(\a[17] ), .dout(n2775));
  jor  g02712(.dina(n2775), .dinb(n2766), .dout(n2776));
  jxor g02713(.dina(n2287), .dinb(n2286), .dout(n2777));
  jnot g02714(.din(n2777), .dout(n2778));
  jxor g02715(.dina(n2641), .dinb(n2640), .dout(n2779));
  jor  g02716(.dina(n2779), .dinb(n2744), .dout(n2780));
  jor  g02717(.dina(n2749), .dinb(n2428), .dout(n2781));
  jor  g02718(.dina(n2753), .dinb(n2629), .dout(n2782));
  jand g02719(.dina(n2782), .dinb(n2781), .dout(n2783));
  jor  g02720(.dina(n2758), .dinb(n2174), .dout(n2784));
  jand g02721(.dina(n2784), .dinb(n2783), .dout(n2785));
  jand g02722(.dina(n2785), .dinb(n2780), .dout(n2786));
  jxor g02723(.dina(n2786), .dinb(\a[17] ), .dout(n2787));
  jor  g02724(.dina(n2787), .dinb(n2778), .dout(n2788));
  jxor g02725(.dina(n2284), .dinb(n2283), .dout(n2789));
  jor  g02726(.dina(n2744), .dinb(n2430), .dout(n2790));
  jor  g02727(.dina(n2749), .dinb(n2174), .dout(n2791));
  jor  g02728(.dina(n2753), .dinb(n2428), .dout(n2792));
  jor  g02729(.dina(n2758), .dinb(n1954), .dout(n2793));
  jand g02730(.dina(n2793), .dinb(n2792), .dout(n2794));
  jand g02731(.dina(n2794), .dinb(n2791), .dout(n2795));
  jand g02732(.dina(n2795), .dinb(n2790), .dout(n2796));
  jxor g02733(.dina(n2796), .dinb(n2441), .dout(n2797));
  jand g02734(.dina(n2797), .dinb(n2789), .dout(n2798));
  jxor g02735(.dina(n2281), .dinb(n2280), .dout(n2799));
  jnot g02736(.din(n2799), .dout(n2800));
  jor  g02737(.dina(n2744), .dinb(n2176), .dout(n2801));
  jor  g02738(.dina(n2749), .dinb(n1954), .dout(n2802));
  jor  g02739(.dina(n2758), .dinb(n2057), .dout(n2803));
  jand g02740(.dina(n2803), .dinb(n2802), .dout(n2804));
  jor  g02741(.dina(n2753), .dinb(n2174), .dout(n2805));
  jand g02742(.dina(n2805), .dinb(n2804), .dout(n2806));
  jand g02743(.dina(n2806), .dinb(n2801), .dout(n2807));
  jxor g02744(.dina(n2807), .dinb(\a[17] ), .dout(n2808));
  jor  g02745(.dina(n2808), .dinb(n2800), .dout(n2809));
  jxor g02746(.dina(n2276), .dinb(n2275), .dout(n2810));
  jor  g02747(.dina(n2744), .dinb(n2197), .dout(n2811));
  jor  g02748(.dina(n2758), .dinb(n1790), .dout(n2812));
  jor  g02749(.dina(n2753), .dinb(n1954), .dout(n2813));
  jor  g02750(.dina(n2749), .dinb(n2057), .dout(n2814));
  jand g02751(.dina(n2814), .dinb(n2813), .dout(n2815));
  jand g02752(.dina(n2815), .dinb(n2812), .dout(n2816));
  jand g02753(.dina(n2816), .dinb(n2811), .dout(n2817));
  jxor g02754(.dina(n2817), .dinb(n2441), .dout(n2818));
  jand g02755(.dina(n2818), .dinb(n2810), .dout(n2819));
  jxor g02756(.dina(n2272), .dinb(n2264), .dout(n2820));
  jor  g02757(.dina(n2744), .dinb(n2208), .dout(n2821));
  jor  g02758(.dina(n2749), .dinb(n1790), .dout(n2822));
  jor  g02759(.dina(n2758), .dinb(n1606), .dout(n2823));
  jor  g02760(.dina(n2753), .dinb(n2057), .dout(n2824));
  jand g02761(.dina(n2824), .dinb(n2823), .dout(n2825));
  jand g02762(.dina(n2825), .dinb(n2822), .dout(n2826));
  jand g02763(.dina(n2826), .dinb(n2821), .dout(n2827));
  jxor g02764(.dina(n2827), .dinb(n2441), .dout(n2828));
  jand g02765(.dina(n2828), .dinb(n2820), .dout(n2829));
  jor  g02766(.dina(n2753), .dinb(n1790), .dout(n2830));
  jor  g02767(.dina(n2744), .dinb(n1792), .dout(n2831));
  jor  g02768(.dina(n2758), .dinb(n1448), .dout(n2832));
  jor  g02769(.dina(n2749), .dinb(n1606), .dout(n2833));
  jand g02770(.dina(n2833), .dinb(n2832), .dout(n2834));
  jand g02771(.dina(n2834), .dinb(n2831), .dout(n2835));
  jand g02772(.dina(n2835), .dinb(n2830), .dout(n2836));
  jxor g02773(.dina(n2836), .dinb(\a[17] ), .dout(n2837));
  jnot g02774(.din(n2837), .dout(n2838));
  jor  g02775(.dina(n2251), .dinb(n2196), .dout(n2839));
  jxor g02776(.dina(n2839), .dinb(n2259), .dout(n2840));
  jand g02777(.dina(n2840), .dinb(n2838), .dout(n2841));
  jand g02778(.dina(n2248), .dinb(\a[20] ), .dout(n2842));
  jxor g02779(.dina(n2842), .dinb(n2246), .dout(n2843));
  jnot g02780(.din(n2843), .dout(n2844));
  jor  g02781(.dina(n2744), .dinb(n1608), .dout(n2845));
  jor  g02782(.dina(n2749), .dinb(n1448), .dout(n2846));
  jor  g02783(.dina(n2758), .dinb(n1255), .dout(n2847));
  jand g02784(.dina(n2847), .dinb(n2846), .dout(n2848));
  jor  g02785(.dina(n2753), .dinb(n1606), .dout(n2849));
  jand g02786(.dina(n2849), .dinb(n2848), .dout(n2850));
  jand g02787(.dina(n2850), .dinb(n2845), .dout(n2851));
  jxor g02788(.dina(n2851), .dinb(\a[17] ), .dout(n2852));
  jor  g02789(.dina(n2852), .dinb(n2844), .dout(n2853));
  jand g02790(.dina(n2743), .dinb(n728), .dout(n2854));
  jand g02791(.dina(n2748), .dinb(n438), .dout(n2855));
  jand g02792(.dina(n2752), .dinb(n795), .dout(n2856));
  jor  g02793(.dina(n2856), .dinb(n2855), .dout(n2857));
  jor  g02794(.dina(n2857), .dinb(n2854), .dout(n2858));
  jnot g02795(.din(n2858), .dout(n2859));
  jand g02796(.dina(n2741), .dinb(n438), .dout(n2860));
  jnot g02797(.din(n2860), .dout(n2861));
  jand g02798(.dina(n2861), .dinb(\a[17] ), .dout(n2862));
  jand g02799(.dina(n2862), .dinb(n2859), .dout(n2863));
  jand g02800(.dina(n2743), .dinb(n1639), .dout(n2864));
  jand g02801(.dina(n2748), .dinb(n795), .dout(n2865));
  jand g02802(.dina(n2752), .dinb(n1175), .dout(n2866));
  jor  g02803(.dina(n2866), .dinb(n2865), .dout(n2867));
  jand g02804(.dina(n2757), .dinb(n438), .dout(n2868));
  jor  g02805(.dina(n2868), .dinb(n2867), .dout(n2869));
  jor  g02806(.dina(n2869), .dinb(n2864), .dout(n2870));
  jnot g02807(.din(n2870), .dout(n2871));
  jand g02808(.dina(n2871), .dinb(n2863), .dout(n2872));
  jand g02809(.dina(n2872), .dinb(n2248), .dout(n2873));
  jnot g02810(.din(n2873), .dout(n2874));
  jxor g02811(.dina(n2872), .dinb(n2248), .dout(n2875));
  jnot g02812(.din(n2875), .dout(n2876));
  jor  g02813(.dina(n2744), .dinb(n1656), .dout(n2877));
  jor  g02814(.dina(n2753), .dinb(n1448), .dout(n2878));
  jor  g02815(.dina(n2749), .dinb(n1255), .dout(n2879));
  jand g02816(.dina(n2879), .dinb(n2878), .dout(n2880));
  jor  g02817(.dina(n2758), .dinb(n726), .dout(n2881));
  jand g02818(.dina(n2881), .dinb(n2880), .dout(n2882));
  jand g02819(.dina(n2882), .dinb(n2877), .dout(n2883));
  jxor g02820(.dina(n2883), .dinb(\a[17] ), .dout(n2884));
  jor  g02821(.dina(n2884), .dinb(n2876), .dout(n2885));
  jand g02822(.dina(n2885), .dinb(n2874), .dout(n2886));
  jnot g02823(.din(n2886), .dout(n2887));
  jxor g02824(.dina(n2852), .dinb(n2844), .dout(n2888));
  jand g02825(.dina(n2888), .dinb(n2887), .dout(n2889));
  jnot g02826(.din(n2889), .dout(n2890));
  jand g02827(.dina(n2890), .dinb(n2853), .dout(n2891));
  jnot g02828(.din(n2891), .dout(n2892));
  jxor g02829(.dina(n2840), .dinb(n2838), .dout(n2893));
  jand g02830(.dina(n2893), .dinb(n2892), .dout(n2894));
  jor  g02831(.dina(n2894), .dinb(n2841), .dout(n2895));
  jxor g02832(.dina(n2828), .dinb(n2820), .dout(n2896));
  jand g02833(.dina(n2896), .dinb(n2895), .dout(n2897));
  jor  g02834(.dina(n2897), .dinb(n2829), .dout(n2898));
  jxor g02835(.dina(n2818), .dinb(n2810), .dout(n2899));
  jand g02836(.dina(n2899), .dinb(n2898), .dout(n2900));
  jor  g02837(.dina(n2900), .dinb(n2819), .dout(n2901));
  jxor g02838(.dina(n2808), .dinb(n2800), .dout(n2902));
  jand g02839(.dina(n2902), .dinb(n2901), .dout(n2903));
  jnot g02840(.din(n2903), .dout(n2904));
  jand g02841(.dina(n2904), .dinb(n2809), .dout(n2905));
  jnot g02842(.din(n2905), .dout(n2906));
  jxor g02843(.dina(n2797), .dinb(n2789), .dout(n2907));
  jand g02844(.dina(n2907), .dinb(n2906), .dout(n2908));
  jor  g02845(.dina(n2908), .dinb(n2798), .dout(n2909));
  jxor g02846(.dina(n2787), .dinb(n2778), .dout(n2910));
  jand g02847(.dina(n2910), .dinb(n2909), .dout(n2911));
  jnot g02848(.din(n2911), .dout(n2912));
  jand g02849(.dina(n2912), .dinb(n2788), .dout(n2913));
  jnot g02850(.din(n2913), .dout(n2914));
  jxor g02851(.dina(n2775), .dinb(n2766), .dout(n2915));
  jand g02852(.dina(n2915), .dinb(n2914), .dout(n2916));
  jnot g02853(.din(n2916), .dout(n2917));
  jand g02854(.dina(n2917), .dinb(n2776), .dout(n2918));
  jnot g02855(.din(n2918), .dout(n2919));
  jxor g02856(.dina(n2763), .dinb(n2440), .dout(n2920));
  jand g02857(.dina(n2920), .dinb(n2919), .dout(n2921));
  jor  g02858(.dina(n2921), .dinb(n2764), .dout(n2922));
  jand g02859(.dina(n2438), .dinb(n2324), .dout(n2923));
  jand g02860(.dina(n2439), .dinb(n2294), .dout(n2924));
  jor  g02861(.dina(n2924), .dinb(n2923), .dout(n2925));
  jand g02862(.dina(n2322), .dinb(n2314), .dout(n2926));
  jand g02863(.dina(n2323), .dinb(n2297), .dout(n2927));
  jor  g02864(.dina(n2927), .dinb(n2926), .dout(n2928));
  jnot g02865(.din(n2300), .dout(n2929));
  jand g02866(.dina(n2929), .dinb(n2298), .dout(n2930));
  jnot g02867(.din(n2930), .dout(n2931));
  jor  g02868(.dina(n2313), .dinb(n2302), .dout(n2932));
  jand g02869(.dina(n2932), .dinb(n2931), .dout(n2933));
  jnot g02870(.din(n2933), .dout(n2934));
  jxor g02871(.dina(\a[29] ), .dinb(\a[28] ), .dout(n2935));
  jand g02872(.dina(n2935), .dinb(n64), .dout(n2936));
  jand g02873(.dina(n2936), .dinb(n728), .dout(n2937));
  jnot g02874(.din(n64), .dout(n2938));
  jxor g02875(.dina(\a[28] ), .dinb(\a[27] ), .dout(n2939));
  jand g02876(.dina(n2939), .dinb(n2938), .dout(n2940));
  jand g02877(.dina(n2940), .dinb(n438), .dout(n2941));
  jnot g02878(.din(n2935), .dout(n2942));
  jand g02879(.dina(n2942), .dinb(n64), .dout(n2943));
  jand g02880(.dina(n2943), .dinb(n795), .dout(n2944));
  jor  g02881(.dina(n2944), .dinb(n2941), .dout(n2945));
  jor  g02882(.dina(n2945), .dinb(n2937), .dout(n2946));
  jor  g02883(.dina(n2299), .dinb(n93), .dout(n2947));
  jxor g02884(.dina(n2947), .dinb(n2946), .dout(n2948));
  jor  g02885(.dina(n1608), .dinb(n2303), .dout(n2949));
  jor  g02886(.dina(n1448), .dinb(n2306), .dout(n2950));
  jor  g02887(.dina(n1805), .dinb(n1255), .dout(n2951));
  jand g02888(.dina(n2951), .dinb(n2950), .dout(n2952));
  jor  g02889(.dina(n1606), .dinb(n2309), .dout(n2953));
  jand g02890(.dina(n2953), .dinb(n2952), .dout(n2954));
  jand g02891(.dina(n2954), .dinb(n2949), .dout(n2955));
  jxor g02892(.dina(n2955), .dinb(\a[26] ), .dout(n2956));
  jxor g02893(.dina(n2956), .dinb(n2948), .dout(n2957));
  jxor g02894(.dina(n2957), .dinb(n2934), .dout(n2958));
  jor  g02895(.dina(n2197), .dinb(n807), .dout(n2959));
  jor  g02896(.dina(n2057), .dinb(n1613), .dout(n2960));
  jor  g02897(.dina(n1954), .dinb(n1621), .dout(n2961));
  jor  g02898(.dina(n1790), .dinb(n1617), .dout(n2962));
  jand g02899(.dina(n2962), .dinb(n2961), .dout(n2963));
  jand g02900(.dina(n2963), .dinb(n2960), .dout(n2964));
  jand g02901(.dina(n2964), .dinb(n2959), .dout(n2965));
  jxor g02902(.dina(n2965), .dinb(n65), .dout(n2966));
  jxor g02903(.dina(n2966), .dinb(n2958), .dout(n2967));
  jxor g02904(.dina(n2967), .dinb(n2928), .dout(n2968));
  jnot g02905(.din(n2968), .dout(n2969));
  jor  g02906(.dina(n2779), .dinb(n1820), .dout(n2970));
  jor  g02907(.dina(n2428), .dinb(n2181), .dout(n2971));
  jor  g02908(.dina(n2629), .dinb(n2189), .dout(n2972));
  jand g02909(.dina(n2972), .dinb(n2971), .dout(n2973));
  jor  g02910(.dina(n2186), .dinb(n2174), .dout(n2974));
  jand g02911(.dina(n2974), .dinb(n2973), .dout(n2975));
  jand g02912(.dina(n2975), .dinb(n2970), .dout(n2976));
  jxor g02913(.dina(n2976), .dinb(\a[20] ), .dout(n2977));
  jxor g02914(.dina(n2977), .dinb(n2969), .dout(n2978));
  jxor g02915(.dina(n2978), .dinb(n2925), .dout(n2979));
  jnot g02916(.din(n2979), .dout(n2980));
  jand g02917(.dina(n512), .dinb(n880), .dout(n2981));
  jand g02918(.dina(n2981), .dinb(n1779), .dout(n2982));
  jand g02919(.dina(n2982), .dinb(n1245), .dout(n2983));
  jand g02920(.dina(n1686), .dinb(n1432), .dout(n2984));
  jand g02921(.dina(n848), .dinb(n680), .dout(n2985));
  jand g02922(.dina(n2985), .dinb(n1832), .dout(n2986));
  jand g02923(.dina(n2986), .dinb(n2984), .dout(n2987));
  jand g02924(.dina(n983), .dinb(n1532), .dout(n2988));
  jand g02925(.dina(n2988), .dinb(n2987), .dout(n2989));
  jand g02926(.dina(n2989), .dinb(n2983), .dout(n2990));
  jand g02927(.dina(n1868), .dinb(n703), .dout(n2991));
  jand g02928(.dina(n2586), .dinb(n136), .dout(n2992));
  jand g02929(.dina(n1218), .dinb(n1591), .dout(n2993));
  jand g02930(.dina(n1713), .dinb(n320), .dout(n2994));
  jand g02931(.dina(n2994), .dinb(n2993), .dout(n2995));
  jand g02932(.dina(n2995), .dinb(n2992), .dout(n2996));
  jand g02933(.dina(n660), .dinb(n1465), .dout(n2997));
  jand g02934(.dina(n2997), .dinb(n988), .dout(n2998));
  jand g02935(.dina(n2998), .dinb(n2996), .dout(n2999));
  jand g02936(.dina(n2999), .dinb(n2991), .dout(n3000));
  jand g02937(.dina(n1038), .dinb(n718), .dout(n3001));
  jand g02938(.dina(n3001), .dinb(n1283), .dout(n3002));
  jand g02939(.dina(n445), .dinb(n492), .dout(n3003));
  jand g02940(.dina(n1708), .dinb(n551), .dout(n3004));
  jand g02941(.dina(n3004), .dinb(n3003), .dout(n3005));
  jand g02942(.dina(n3005), .dinb(n3002), .dout(n3006));
  jand g02943(.dina(n1167), .dinb(n713), .dout(n3007));
  jand g02944(.dina(n3007), .dinb(n966), .dout(n3008));
  jand g02945(.dina(n3008), .dinb(n3006), .dout(n3009));
  jand g02946(.dina(n3009), .dinb(n3000), .dout(n3010));
  jand g02947(.dina(n3010), .dinb(n2990), .dout(n3011));
  jand g02948(.dina(n3011), .dinb(n600), .dout(n3012));
  jand g02949(.dina(n3012), .dinb(n1310), .dout(n3013));
  jand g02950(.dina(n1697), .dinb(n716), .dout(n3014));
  jand g02951(.dina(n1159), .dinb(n168), .dout(n3015));
  jand g02952(.dina(n3015), .dinb(n1366), .dout(n3016));
  jand g02953(.dina(n3016), .dinb(n2332), .dout(n3017));
  jand g02954(.dina(n3017), .dinb(n3014), .dout(n3018));
  jand g02955(.dina(n1470), .dinb(n548), .dout(n3019));
  jand g02956(.dina(n950), .dinb(n440), .dout(n3020));
  jand g02957(.dina(n1580), .dinb(n622), .dout(n3021));
  jand g02958(.dina(n3021), .dinb(n3020), .dout(n3022));
  jand g02959(.dina(n3022), .dinb(n3019), .dout(n3023));
  jand g02960(.dina(n3023), .dinb(n3018), .dout(n3024));
  jand g02961(.dina(n1767), .dinb(n844), .dout(n3025));
  jand g02962(.dina(n869), .dinb(n537), .dout(n3026));
  jand g02963(.dina(n3026), .dinb(n1163), .dout(n3027));
  jand g02964(.dina(n3027), .dinb(n672), .dout(n3028));
  jand g02965(.dina(n3028), .dinb(n3025), .dout(n3029));
  jand g02966(.dina(n1743), .dinb(n1226), .dout(n3030));
  jand g02967(.dina(n3030), .dinb(n1449), .dout(n3031));
  jand g02968(.dina(n1246), .dinb(n900), .dout(n3032));
  jand g02969(.dina(n3032), .dinb(n3031), .dout(n3033));
  jand g02970(.dina(n3033), .dinb(n908), .dout(n3034));
  jand g02971(.dina(n3034), .dinb(n3029), .dout(n3035));
  jand g02972(.dina(n3035), .dinb(n3024), .dout(n3036));
  jand g02973(.dina(n1473), .dinb(n1257), .dout(n3037));
  jand g02974(.dina(n3037), .dinb(n1324), .dout(n3038));
  jand g02975(.dina(n1098), .dinb(n678), .dout(n3039));
  jand g02976(.dina(n3039), .dinb(n1292), .dout(n3040));
  jand g02977(.dina(n3040), .dinb(n2561), .dout(n3041));
  jand g02978(.dina(n3041), .dinb(n3038), .dout(n3042));
  jand g02979(.dina(n3042), .dinb(n2687), .dout(n3043));
  jand g02980(.dina(n461), .dinb(n463), .dout(n3044));
  jand g02981(.dina(n1560), .dinb(n411), .dout(n3045));
  jand g02982(.dina(n1378), .dinb(n654), .dout(n3046));
  jand g02983(.dina(n3046), .dinb(n3045), .dout(n3047));
  jnot g02984(.din(n1059), .dout(n3048));
  jand g02985(.dina(n1453), .dinb(n1361), .dout(n3049));
  jand g02986(.dina(n1219), .dinb(n929), .dout(n3050));
  jand g02987(.dina(n3050), .dinb(n3049), .dout(n3051));
  jand g02988(.dina(n3051), .dinb(n3048), .dout(n3052));
  jand g02989(.dina(n3052), .dinb(n3047), .dout(n3053));
  jand g02990(.dina(n3053), .dinb(n3044), .dout(n3054));
  jand g02991(.dina(n3054), .dinb(n3043), .dout(n3055));
  jand g02992(.dina(n442), .dinb(n582), .dout(n3056));
  jand g02993(.dina(n3056), .dinb(n328), .dout(n3057));
  jand g02994(.dina(n1515), .dinb(n917), .dout(n3058));
  jand g02995(.dina(n3058), .dinb(n1315), .dout(n3059));
  jand g02996(.dina(n3059), .dinb(n3057), .dout(n3060));
  jand g02997(.dina(n3060), .dinb(n122), .dout(n3061));
  jand g02998(.dina(n2154), .dinb(n2077), .dout(n3062));
  jand g02999(.dina(n685), .dinb(n1334), .dout(n3063));
  jand g03000(.dina(n3063), .dinb(n638), .dout(n3064));
  jand g03001(.dina(n3064), .dinb(n3062), .dout(n3065));
  jand g03002(.dina(n481), .dinb(n1316), .dout(n3066));
  jand g03003(.dina(n3066), .dinb(n1852), .dout(n3067));
  jand g03004(.dina(n3067), .dinb(n3065), .dout(n3068));
  jand g03005(.dina(n3068), .dinb(n3061), .dout(n3069));
  jand g03006(.dina(n3069), .dinb(n3055), .dout(n3070));
  jand g03007(.dina(n3070), .dinb(n3036), .dout(n3071));
  jand g03008(.dina(n3071), .dinb(n3013), .dout(n3072));
  jor  g03009(.dina(n3072), .dinb(n2753), .dout(n3073));
  jnot g03010(.din(n2738), .dout(n3074));
  jand g03011(.dina(n3074), .dinb(n2554), .dout(n3075));
  jnot g03012(.din(n3075), .dout(n3076));
  jnot g03013(.din(n2739), .dout(n3077));
  jor  g03014(.dina(n3077), .dinb(n2648), .dout(n3078));
  jand g03015(.dina(n3078), .dinb(n3076), .dout(n3079));
  jxor g03016(.dina(n3072), .dinb(n2738), .dout(n3080));
  jxor g03017(.dina(n3080), .dinb(n3079), .dout(n3081));
  jor  g03018(.dina(n3081), .dinb(n2744), .dout(n3082));
  jor  g03019(.dina(n2749), .dinb(n2738), .dout(n3083));
  jor  g03020(.dina(n2758), .dinb(n2553), .dout(n3084));
  jand g03021(.dina(n3084), .dinb(n3083), .dout(n3085));
  jand g03022(.dina(n3085), .dinb(n3082), .dout(n3086));
  jand g03023(.dina(n3086), .dinb(n3073), .dout(n3087));
  jxor g03024(.dina(n3087), .dinb(\a[17] ), .dout(n3088));
  jxor g03025(.dina(n3088), .dinb(n2980), .dout(n3089));
  jxor g03026(.dina(n3089), .dinb(n2922), .dout(n3090));
  jnot g03027(.din(n3090), .dout(n3091));
  jand g03028(.dina(n1108), .dinb(n871), .dout(n3092));
  jand g03029(.dina(n1559), .dinb(n1213), .dout(n3093));
  jand g03030(.dina(n3093), .dinb(n1772), .dout(n3094));
  jand g03031(.dina(n3094), .dinb(n811), .dout(n3095));
  jand g03032(.dina(n3095), .dinb(n3092), .dout(n3096));
  jand g03033(.dina(n3096), .dinb(n978), .dout(n3097));
  jand g03034(.dina(n1218), .dinb(n496), .dout(n3098));
  jand g03035(.dina(n1016), .dinb(n1583), .dout(n3099));
  jand g03036(.dina(n3099), .dinb(n1702), .dout(n3100));
  jand g03037(.dina(n3100), .dinb(n3098), .dout(n3101));
  jnot g03038(.din(n1081), .dout(n3102));
  jand g03039(.dina(n1237), .dinb(n3102), .dout(n3103));
  jand g03040(.dina(n3103), .dinb(n880), .dout(n3104));
  jand g03041(.dina(n3104), .dinb(n3101), .dout(n3105));
  jand g03042(.dina(n3105), .dinb(n3097), .dout(n3106));
  jand g03043(.dina(n3106), .dinb(n1779), .dout(n3107));
  jand g03044(.dina(n1453), .dinb(n1575), .dout(n3108));
  jand g03045(.dina(n3108), .dinb(n1495), .dout(n3109));
  jand g03046(.dina(n3109), .dinb(n1743), .dout(n3110));
  jand g03047(.dina(n3110), .dinb(n1096), .dout(n3111));
  jand g03048(.dina(n672), .dinb(n411), .dout(n3112));
  jand g03049(.dina(n3112), .dinb(n2721), .dout(n3113));
  jand g03050(.dina(n3113), .dinb(n121), .dout(n3114));
  jand g03051(.dina(n3114), .dinb(n3111), .dout(n3115));
  jand g03052(.dina(n1042), .dinb(n132), .dout(n3116));
  jand g03053(.dina(n685), .dinb(n1238), .dout(n3117));
  jand g03054(.dina(n3117), .dinb(n465), .dout(n3118));
  jand g03055(.dina(n3118), .dinb(n1782), .dout(n3119));
  jand g03056(.dina(n848), .dinb(n1429), .dout(n3120));
  jand g03057(.dina(n3120), .dinb(n2385), .dout(n3121));
  jand g03058(.dina(n553), .dinb(n831), .dout(n3122));
  jand g03059(.dina(n3122), .dinb(n3121), .dout(n3123));
  jand g03060(.dina(n3123), .dinb(n3119), .dout(n3124));
  jand g03061(.dina(n1725), .dinb(n1393), .dout(n3125));
  jand g03062(.dina(n3125), .dinb(n3124), .dout(n3126));
  jand g03063(.dina(n3126), .dinb(n3116), .dout(n3127));
  jand g03064(.dina(n3127), .dinb(n3115), .dout(n3128));
  jand g03065(.dina(n3128), .dinb(n3107), .dout(n3129));
  jand g03066(.dina(n1360), .dinb(n1036), .dout(n3130));
  jand g03067(.dina(n3130), .dinb(n948), .dout(n3131));
  jand g03068(.dina(n3131), .dinb(n1167), .dout(n3132));
  jand g03069(.dina(n2100), .dinb(n1309), .dout(n3133));
  jand g03070(.dina(n3133), .dinb(n1700), .dout(n3134));
  jand g03071(.dina(n3134), .dinb(n3132), .dout(n3135));
  jand g03072(.dina(n1207), .dinb(n1460), .dout(n3136));
  jand g03073(.dina(n3136), .dinb(n463), .dout(n3137));
  jand g03074(.dina(n3137), .dinb(n900), .dout(n3138));
  jand g03075(.dina(n3138), .dinb(n521), .dout(n3139));
  jand g03076(.dina(n3139), .dinb(n3135), .dout(n3140));
  jand g03077(.dina(n3140), .dinb(n3129), .dout(n3141));
  jand g03078(.dina(n1227), .dinb(n600), .dout(n3142));
  jand g03079(.dina(n3142), .dinb(n1345), .dout(n3143));
  jand g03080(.dina(n3143), .dinb(n1260), .dout(n3144));
  jand g03081(.dina(n884), .dinb(n135), .dout(n3145));
  jand g03082(.dina(n3145), .dinb(n320), .dout(n3146));
  jand g03083(.dina(n1738), .dinb(n1283), .dout(n3147));
  jand g03084(.dina(n3147), .dinb(n3146), .dout(n3148));
  jand g03085(.dina(n3148), .dinb(n3144), .dout(n3149));
  jand g03086(.dina(n1219), .dinb(n670), .dout(n3150));
  jand g03087(.dina(n3150), .dinb(n1942), .dout(n3151));
  jand g03088(.dina(n3151), .dinb(n3149), .dout(n3152));
  jand g03089(.dina(n430), .dinb(n582), .dout(n3153));
  jand g03090(.dina(n1591), .dinb(n130), .dout(n3154));
  jand g03091(.dina(n901), .dinb(n108), .dout(n3155));
  jand g03092(.dina(n3155), .dinb(n3154), .dout(n3156));
  jand g03093(.dina(n3156), .dinb(n3153), .dout(n3157));
  jand g03094(.dina(n3157), .dinb(n839), .dout(n3158));
  jand g03095(.dina(n3158), .dinb(n3152), .dout(n3159));
  jand g03096(.dina(n1697), .dinb(n492), .dout(n3160));
  jand g03097(.dina(n693), .dinb(n1344), .dout(n3161));
  jand g03098(.dina(n3161), .dinb(n3160), .dout(n3162));
  jand g03099(.dina(n3162), .dinb(n1511), .dout(n3163));
  jand g03100(.dina(n664), .dinb(n655), .dout(n3164));
  jand g03101(.dina(n3164), .dinb(n1822), .dout(n3165));
  jand g03102(.dina(n3165), .dinb(n3163), .dout(n3166));
  jand g03103(.dina(n1361), .dinb(n1203), .dout(n3167));
  jand g03104(.dina(n503), .dinb(n818), .dout(n3168));
  jand g03105(.dina(n3168), .dinb(n3167), .dout(n3169));
  jand g03106(.dina(n3169), .dinb(n1333), .dout(n3170));
  jand g03107(.dina(n3170), .dinb(n2029), .dout(n3171));
  jand g03108(.dina(n3171), .dinb(n3166), .dout(n3172));
  jand g03109(.dina(n826), .dinb(n641), .dout(n3173));
  jand g03110(.dina(n3173), .dinb(n447), .dout(n3174));
  jand g03111(.dina(n3174), .dinb(n1246), .dout(n3175));
  jand g03112(.dina(n925), .dinb(n588), .dout(n3176));
  jand g03113(.dina(n3176), .dinb(n516), .dout(n3177));
  jand g03114(.dina(n895), .dinb(n511), .dout(n3178));
  jand g03115(.dina(n1465), .dinb(n562), .dout(n3179));
  jand g03116(.dina(n3179), .dinb(n3178), .dout(n3180));
  jand g03117(.dina(n3180), .dinb(n3177), .dout(n3181));
  jand g03118(.dina(n965), .dinb(n1233), .dout(n3182));
  jand g03119(.dina(n1315), .dinb(n168), .dout(n3183));
  jand g03120(.dina(n3183), .dinb(n3182), .dout(n3184));
  jnot g03121(.din(n525), .dout(n3185));
  jand g03122(.dina(n3185), .dinb(n510), .dout(n3186));
  jand g03123(.dina(n3186), .dinb(n3184), .dout(n3187));
  jand g03124(.dina(n3187), .dinb(n3181), .dout(n3188));
  jand g03125(.dina(n3188), .dinb(n3175), .dout(n3189));
  jand g03126(.dina(n3189), .dinb(n3172), .dout(n3190));
  jand g03127(.dina(n3020), .dinb(n481), .dout(n3191));
  jand g03128(.dina(n873), .dinb(n470), .dout(n3192));
  jand g03129(.dina(n3192), .dinb(n662), .dout(n3193));
  jand g03130(.dina(n3193), .dinb(n3191), .dout(n3194));
  jand g03131(.dina(n534), .dinb(n472), .dout(n3195));
  jand g03132(.dina(n3195), .dinb(n1334), .dout(n3196));
  jand g03133(.dina(n3196), .dinb(n3194), .dout(n3197));
  jand g03134(.dina(n469), .dinb(n954), .dout(n3198));
  jand g03135(.dina(n3198), .dinb(n704), .dout(n3199));
  jand g03136(.dina(n3199), .dinb(n3197), .dout(n3200));
  jand g03137(.dina(n3200), .dinb(n3190), .dout(n3201));
  jand g03138(.dina(n3201), .dinb(n3159), .dout(n3202));
  jand g03139(.dina(n3202), .dinb(n3141), .dout(n3203));
  jxor g03140(.dina(\a[14] ), .dinb(\a[13] ), .dout(n3204));
  jxor g03141(.dina(\a[12] ), .dinb(\a[11] ), .dout(n3205));
  jnot g03142(.din(n3205), .dout(n3206));
  jxor g03143(.dina(\a[13] ), .dinb(\a[12] ), .dout(n3207));
  jnot g03144(.din(n3207), .dout(n3208));
  jand g03145(.dina(n3208), .dinb(n3206), .dout(n3209));
  jand g03146(.dina(n3209), .dinb(n3204), .dout(n3210));
  jnot g03147(.din(n3210), .dout(n3211));
  jor  g03148(.dina(n3211), .dinb(n3203), .dout(n3212));
  jnot g03149(.din(n3203), .dout(n3213));
  jand g03150(.dina(n718), .dinb(n1317), .dout(n3214));
  jand g03151(.dina(n965), .dinb(n1682), .dout(n3215));
  jand g03152(.dina(n3215), .dinb(n3214), .dout(n3216));
  jand g03153(.dina(n1373), .dinb(n266), .dout(n3217));
  jand g03154(.dina(n645), .dinb(n130), .dout(n3218));
  jand g03155(.dina(n3218), .dinb(n3217), .dout(n3219));
  jand g03156(.dina(n3219), .dinb(n3173), .dout(n3220));
  jand g03157(.dina(n3220), .dinb(n3216), .dout(n3221));
  jand g03158(.dina(n1460), .dinb(n1270), .dout(n3222));
  jand g03159(.dina(n3222), .dinb(n1301), .dout(n3223));
  jand g03160(.dina(n3223), .dinb(n696), .dout(n3224));
  jand g03161(.dina(n1426), .dinb(n691), .dout(n3225));
  jand g03162(.dina(n1511), .dinb(n1532), .dout(n3226));
  jand g03163(.dina(n3226), .dinb(n703), .dout(n3227));
  jand g03164(.dina(n3227), .dinb(n3225), .dout(n3228));
  jand g03165(.dina(n3228), .dinb(n3224), .dout(n3229));
  jand g03166(.dina(n3229), .dinb(n3221), .dout(n3230));
  jand g03167(.dina(n352), .dinb(n1701), .dout(n3231));
  jand g03168(.dina(n981), .dinb(n178), .dout(n3232));
  jand g03169(.dina(n1237), .dinb(n82), .dout(n3233));
  jand g03170(.dina(n3233), .dinb(n3232), .dout(n3234));
  jand g03171(.dina(n3234), .dinb(n3231), .dout(n3235));
  jand g03172(.dina(n1583), .dinb(n470), .dout(n3236));
  jand g03173(.dina(n3236), .dinb(n583), .dout(n3237));
  jand g03174(.dina(n632), .dinb(n1310), .dout(n3238));
  jand g03175(.dina(n3238), .dinb(n560), .dout(n3239));
  jand g03176(.dina(n1522), .dinb(n92), .dout(n3240));
  jand g03177(.dina(n3240), .dinb(n1260), .dout(n3241));
  jand g03178(.dina(n3241), .dinb(n3239), .dout(n3242));
  jand g03179(.dina(n3242), .dinb(n3237), .dout(n3243));
  jand g03180(.dina(n3243), .dinb(n3235), .dout(n3244));
  jand g03181(.dina(n3244), .dinb(n2576), .dout(n3245));
  jand g03182(.dina(n3245), .dinb(n3230), .dout(n3246));
  jand g03183(.dina(n1495), .dinb(n270), .dout(n3247));
  jand g03184(.dina(n638), .dinb(n1040), .dout(n3248));
  jand g03185(.dina(n3248), .dinb(n3247), .dout(n3249));
  jand g03186(.dina(n1098), .dinb(n1315), .dout(n3250));
  jand g03187(.dina(n2100), .dinb(n1903), .dout(n3251));
  jand g03188(.dina(n3251), .dinb(n3250), .dout(n3252));
  jand g03189(.dina(n3252), .dinb(n3249), .dout(n3253));
  jand g03190(.dina(n1167), .dinb(n135), .dout(n3254));
  jand g03191(.dina(n3254), .dinb(n700), .dout(n3255));
  jand g03192(.dina(n1890), .dinb(n1688), .dout(n3256));
  jand g03193(.dina(n3256), .dinb(n3255), .dout(n3257));
  jand g03194(.dina(n3257), .dinb(n3253), .dout(n3258));
  jand g03195(.dina(n871), .dinb(n653), .dout(n3259));
  jand g03196(.dina(n3259), .dinb(n2522), .dout(n3260));
  jand g03197(.dina(n925), .dinb(n1756), .dout(n3261));
  jand g03198(.dina(n3261), .dinb(n685), .dout(n3262));
  jand g03199(.dina(n3262), .dinb(n3260), .dout(n3263));
  jand g03200(.dina(n1005), .dinb(n480), .dout(n3264));
  jand g03201(.dina(n1366), .dinb(n1292), .dout(n3265));
  jand g03202(.dina(n3265), .dinb(n3264), .dout(n3266));
  jand g03203(.dina(n442), .dinb(n541), .dout(n3267));
  jand g03204(.dina(n3267), .dinb(n2716), .dout(n3268));
  jand g03205(.dina(n3268), .dinb(n3266), .dout(n3269));
  jand g03206(.dina(n3269), .dinb(n3263), .dout(n3270));
  jand g03207(.dina(n630), .dinb(n2028), .dout(n3271));
  jand g03208(.dina(n1246), .dinb(n1228), .dout(n3272));
  jand g03209(.dina(n3272), .dinb(n472), .dout(n3273));
  jand g03210(.dina(n3273), .dinb(n3271), .dout(n3274));
  jand g03211(.dina(n3274), .dinb(n2152), .dout(n3275));
  jand g03212(.dina(n1846), .dinb(n843), .dout(n3276));
  jand g03213(.dina(n3276), .dinb(n1751), .dout(n3277));
  jand g03214(.dina(n3277), .dinb(n2380), .dout(n3278));
  jand g03215(.dina(n1731), .dinb(n454), .dout(n3279));
  jand g03216(.dina(n3279), .dinb(n2526), .dout(n3280));
  jand g03217(.dina(n3280), .dinb(n3278), .dout(n3281));
  jand g03218(.dina(n3281), .dinb(n3275), .dout(n3282));
  jand g03219(.dina(n3282), .dinb(n3270), .dout(n3283));
  jand g03220(.dina(n3283), .dinb(n2593), .dout(n3284));
  jand g03221(.dina(n3284), .dinb(n3258), .dout(n3285));
  jand g03222(.dina(n3285), .dinb(n3246), .dout(n3286));
  jnot g03223(.din(n3286), .dout(n3287));
  jand g03224(.dina(n3287), .dinb(n3213), .dout(n3288));
  jnot g03225(.din(n3288), .dout(n3289));
  jnot g03226(.din(n3072), .dout(n3290));
  jand g03227(.dina(n3213), .dinb(n3290), .dout(n3291));
  jnot g03228(.din(n3291), .dout(n3292));
  jand g03229(.dina(n3290), .dinb(n3074), .dout(n3293));
  jnot g03230(.din(n3293), .dout(n3294));
  jnot g03231(.din(n3080), .dout(n3295));
  jor  g03232(.dina(n3295), .dinb(n3079), .dout(n3296));
  jand g03233(.dina(n3296), .dinb(n3294), .dout(n3297));
  jxor g03234(.dina(n3203), .dinb(n3072), .dout(n3298));
  jnot g03235(.din(n3298), .dout(n3299));
  jor  g03236(.dina(n3299), .dinb(n3297), .dout(n3300));
  jand g03237(.dina(n3300), .dinb(n3292), .dout(n3301));
  jxor g03238(.dina(n3286), .dinb(n3203), .dout(n3302));
  jnot g03239(.din(n3302), .dout(n3303));
  jor  g03240(.dina(n3303), .dinb(n3301), .dout(n3304));
  jand g03241(.dina(n3304), .dinb(n3289), .dout(n3305));
  jand g03242(.dina(n695), .dinb(n171), .dout(n3306));
  jand g03243(.dina(n3306), .dinb(n583), .dout(n3307));
  jand g03244(.dina(n826), .dinb(n465), .dout(n3308));
  jand g03245(.dina(n3308), .dinb(n3307), .dout(n3309));
  jand g03246(.dina(n3309), .dinb(n3143), .dout(n3310));
  jand g03247(.dina(n713), .dinb(n493), .dout(n3311));
  jand g03248(.dina(n1207), .dinb(n981), .dout(n3312));
  jand g03249(.dina(n3312), .dinb(n3311), .dout(n3313));
  jand g03250(.dina(n3313), .dinb(n1751), .dout(n3314));
  jand g03251(.dina(n3314), .dinb(n1688), .dout(n3315));
  jand g03252(.dina(n3315), .dinb(n3310), .dout(n3316));
  jand g03253(.dina(n1203), .dinb(n501), .dout(n3317));
  jand g03254(.dina(n1465), .dinb(n1360), .dout(n3318));
  jand g03255(.dina(n3318), .dinb(n3317), .dout(n3319));
  jand g03256(.dina(n3319), .dinb(n718), .dout(n3320));
  jand g03257(.dina(n3320), .dinb(n1973), .dout(n3321));
  jand g03258(.dina(n1577), .dinb(n931), .dout(n3322));
  jand g03259(.dina(n3322), .dinb(n2597), .dout(n3323));
  jand g03260(.dina(n548), .dinb(n1349), .dout(n3324));
  jand g03261(.dina(n1534), .dinb(n555), .dout(n3325));
  jand g03262(.dina(n3325), .dinb(n3324), .dout(n3326));
  jand g03263(.dina(n3326), .dinb(n3323), .dout(n3327));
  jand g03264(.dina(n1245), .dinb(n560), .dout(n3328));
  jand g03265(.dina(n480), .dinb(n1292), .dout(n3329));
  jand g03266(.dina(n3329), .dinb(n1352), .dout(n3330));
  jand g03267(.dina(n3330), .dinb(n3328), .dout(n3331));
  jand g03268(.dina(n3331), .dinb(n3327), .dout(n3332));
  jand g03269(.dina(n3332), .dinb(n3321), .dout(n3333));
  jand g03270(.dina(n2666), .dinb(n1432), .dout(n3334));
  jand g03271(.dina(n3334), .dinb(n3150), .dout(n3335));
  jand g03272(.dina(n693), .dinb(n454), .dout(n3336));
  jand g03273(.dina(n1511), .dinb(n676), .dout(n3337));
  jand g03274(.dina(n3337), .dinb(n3336), .dout(n3338));
  jand g03275(.dina(n3338), .dinb(n2008), .dout(n3339));
  jand g03276(.dina(n3339), .dinb(n3335), .dout(n3340));
  jand g03277(.dina(n3340), .dinb(n3333), .dout(n3341));
  jand g03278(.dina(n3341), .dinb(n3316), .dout(n3342));
  jand g03279(.dina(n1732), .dinb(n882), .dout(n3343));
  jand g03280(.dina(n3343), .dinb(n3092), .dout(n3344));
  jand g03281(.dina(n921), .dinb(n893), .dout(n3345));
  jand g03282(.dina(n3345), .dinb(n535), .dout(n3346));
  jand g03283(.dina(n3346), .dinb(n2477), .dout(n3347));
  jand g03284(.dina(n3347), .dinb(n3344), .dout(n3348));
  jand g03285(.dina(n1524), .dinb(n1708), .dout(n3349));
  jand g03286(.dina(n1559), .dinb(n114), .dout(n3350));
  jand g03287(.dina(n3350), .dinb(n3349), .dout(n3351));
  jand g03288(.dina(n1495), .dinb(n696), .dout(n3352));
  jand g03289(.dina(n3352), .dinb(n900), .dout(n3353));
  jand g03290(.dina(n3353), .dinb(n3351), .dout(n3354));
  jand g03291(.dina(n3354), .dinb(n3155), .dout(n3355));
  jand g03292(.dina(n1042), .dinb(n1305), .dout(n3356));
  jand g03293(.dina(n1506), .dinb(n1053), .dout(n3357));
  jand g03294(.dina(n3357), .dinb(n351), .dout(n3358));
  jand g03295(.dina(n3358), .dinb(n3356), .dout(n3359));
  jand g03296(.dina(n3359), .dinb(n3355), .dout(n3360));
  jand g03297(.dina(n3360), .dinb(n3348), .dout(n3361));
  jand g03298(.dina(n3361), .dinb(n3342), .dout(n3362));
  jand g03299(.dina(n1437), .dinb(n933), .dout(n3363));
  jand g03300(.dina(n1560), .dinb(n349), .dout(n3364));
  jand g03301(.dina(n1016), .dinb(n1226), .dout(n3365));
  jand g03302(.dina(n3365), .dinb(n3364), .dout(n3366));
  jand g03303(.dina(n3366), .dinb(n1744), .dout(n3367));
  jand g03304(.dina(n463), .dinb(n1040), .dout(n3368));
  jand g03305(.dina(n3368), .dinb(n2608), .dout(n3369));
  jand g03306(.dina(n3369), .dinb(n428), .dout(n3370));
  jand g03307(.dina(n1246), .dinb(n517), .dout(n3371));
  jand g03308(.dina(n3371), .dinb(n632), .dout(n3372));
  jand g03309(.dina(n3372), .dinb(n1167), .dout(n3373));
  jand g03310(.dina(n3373), .dinb(n3370), .dout(n3374));
  jand g03311(.dina(n3374), .dinb(n3367), .dout(n3375));
  jand g03312(.dina(n3375), .dinb(n3363), .dout(n3376));
  jand g03313(.dina(n993), .dinb(n586), .dout(n3377));
  jand g03314(.dina(n3377), .dinb(n2124), .dout(n3378));
  jand g03315(.dina(n461), .dinb(n1317), .dout(n3379));
  jand g03316(.dina(n3379), .dinb(n1846), .dout(n3380));
  jand g03317(.dina(n553), .dinb(n714), .dout(n3381));
  jand g03318(.dina(n3381), .dinb(n1366), .dout(n3382));
  jand g03319(.dina(n3382), .dinb(n3380), .dout(n3383));
  jand g03320(.dina(n3383), .dinb(n3378), .dout(n3384));
  jand g03321(.dina(n983), .dinb(n700), .dout(n3385));
  jand g03322(.dina(n907), .dinb(n1273), .dout(n3386));
  jand g03323(.dina(n3386), .dinb(n3385), .dout(n3387));
  jand g03324(.dina(n678), .dinb(n811), .dout(n3388));
  jand g03325(.dina(n3388), .dinb(n440), .dout(n3389));
  jand g03326(.dina(n1806), .dinb(n186), .dout(n3390));
  jor  g03327(.dina(n3390), .dinb(n1720), .dout(n3391));
  jnot g03328(.din(n3391), .dout(n3392));
  jand g03329(.dina(n3392), .dinb(n3389), .dout(n3393));
  jand g03330(.dina(n3393), .dinb(n3387), .dout(n3394));
  jand g03331(.dina(n3394), .dinb(n3384), .dout(n3395));
  jand g03332(.dina(n1212), .dinb(n1778), .dout(n3396));
  jand g03333(.dina(n1682), .dinb(n542), .dout(n3397));
  jand g03334(.dina(n2148), .dinb(n481), .dout(n3398));
  jand g03335(.dina(n3398), .dinb(n3397), .dout(n3399));
  jand g03336(.dina(n3399), .dinb(n3396), .dout(n3400));
  jand g03337(.dina(n3400), .dinb(n3395), .dout(n3401));
  jand g03338(.dina(n3401), .dinb(n3376), .dout(n3402));
  jand g03339(.dina(n824), .dinb(n516), .dout(n3403));
  jand g03340(.dina(n3403), .dinb(n1738), .dout(n3404));
  jand g03341(.dina(n1583), .dinb(n954), .dout(n3405));
  jand g03342(.dina(n3405), .dinb(n175), .dout(n3406));
  jand g03343(.dina(n3406), .dinb(n3404), .dout(n3407));
  jand g03344(.dina(n1541), .dinb(n1522), .dout(n3408));
  jand g03345(.dina(n647), .dinb(n1316), .dout(n3409));
  jand g03346(.dina(n1375), .dinb(n831), .dout(n3410));
  jand g03347(.dina(n3410), .dinb(n3409), .dout(n3411));
  jand g03348(.dina(n3411), .dinb(n3408), .dout(n3412));
  jand g03349(.dina(n3412), .dinb(n3407), .dout(n3413));
  jand g03350(.dina(n1872), .dinb(n1903), .dout(n3414));
  jand g03351(.dina(n1163), .dinb(n326), .dout(n3415));
  jand g03352(.dina(n3415), .dinb(n1244), .dout(n3416));
  jand g03353(.dina(n3416), .dinb(n3414), .dout(n3417));
  jand g03354(.dina(n3417), .dinb(n3413), .dout(n3418));
  jand g03355(.dina(n3418), .dinb(n3402), .dout(n3419));
  jand g03356(.dina(n3419), .dinb(n3362), .dout(n3420));
  jxor g03357(.dina(n3420), .dinb(n3286), .dout(n3421));
  jxor g03358(.dina(n3421), .dinb(n3305), .dout(n3422));
  jand g03359(.dina(n3205), .dinb(n3204), .dout(n3423));
  jnot g03360(.din(n3423), .dout(n3424));
  jor  g03361(.dina(n3424), .dinb(n3422), .dout(n3425));
  jor  g03362(.dina(n3206), .dinb(n3204), .dout(n3426));
  jor  g03363(.dina(n3426), .dinb(n3420), .dout(n3427));
  jand g03364(.dina(n3207), .dinb(n3206), .dout(n3428));
  jnot g03365(.din(n3428), .dout(n3429));
  jor  g03366(.dina(n3429), .dinb(n3286), .dout(n3430));
  jand g03367(.dina(n3430), .dinb(n3427), .dout(n3431));
  jand g03368(.dina(n3431), .dinb(n3425), .dout(n3432));
  jand g03369(.dina(n3432), .dinb(n3212), .dout(n3433));
  jxor g03370(.dina(n3433), .dinb(\a[14] ), .dout(n3434));
  jor  g03371(.dina(n3434), .dinb(n3091), .dout(n3435));
  jnot g03372(.din(n3435), .dout(n3436));
  jxor g03373(.dina(n2920), .dinb(n2919), .dout(n3437));
  jnot g03374(.din(n3437), .dout(n3438));
  jor  g03375(.dina(n3211), .dinb(n3072), .dout(n3439));
  jxor g03376(.dina(n3302), .dinb(n3301), .dout(n3440));
  jor  g03377(.dina(n3440), .dinb(n3424), .dout(n3441));
  jor  g03378(.dina(n3426), .dinb(n3286), .dout(n3442));
  jor  g03379(.dina(n3429), .dinb(n3203), .dout(n3443));
  jand g03380(.dina(n3443), .dinb(n3442), .dout(n3444));
  jand g03381(.dina(n3444), .dinb(n3441), .dout(n3445));
  jand g03382(.dina(n3445), .dinb(n3439), .dout(n3446));
  jxor g03383(.dina(n3446), .dinb(\a[14] ), .dout(n3447));
  jor  g03384(.dina(n3447), .dinb(n3438), .dout(n3448));
  jxor g03385(.dina(n2915), .dinb(n2914), .dout(n3449));
  jnot g03386(.din(n3449), .dout(n3450));
  jxor g03387(.dina(n3298), .dinb(n3297), .dout(n3451));
  jor  g03388(.dina(n3451), .dinb(n3424), .dout(n3452));
  jor  g03389(.dina(n3429), .dinb(n3072), .dout(n3453));
  jor  g03390(.dina(n3211), .dinb(n2738), .dout(n3454));
  jand g03391(.dina(n3454), .dinb(n3453), .dout(n3455));
  jor  g03392(.dina(n3426), .dinb(n3203), .dout(n3456));
  jand g03393(.dina(n3456), .dinb(n3455), .dout(n3457));
  jand g03394(.dina(n3457), .dinb(n3452), .dout(n3458));
  jxor g03395(.dina(n3458), .dinb(\a[14] ), .dout(n3459));
  jor  g03396(.dina(n3459), .dinb(n3450), .dout(n3460));
  jxor g03397(.dina(n2910), .dinb(n2909), .dout(n3461));
  jnot g03398(.din(n3461), .dout(n3462));
  jor  g03399(.dina(n3426), .dinb(n3072), .dout(n3463));
  jor  g03400(.dina(n3424), .dinb(n3081), .dout(n3464));
  jor  g03401(.dina(n3429), .dinb(n2738), .dout(n3465));
  jor  g03402(.dina(n3211), .dinb(n2553), .dout(n3466));
  jand g03403(.dina(n3466), .dinb(n3465), .dout(n3467));
  jand g03404(.dina(n3467), .dinb(n3464), .dout(n3468));
  jand g03405(.dina(n3468), .dinb(n3463), .dout(n3469));
  jxor g03406(.dina(n3469), .dinb(\a[14] ), .dout(n3470));
  jor  g03407(.dina(n3470), .dinb(n3462), .dout(n3471));
  jxor g03408(.dina(n2907), .dinb(n2906), .dout(n3472));
  jnot g03409(.din(\a[14] ), .dout(n3473));
  jor  g03410(.dina(n3424), .dinb(n2740), .dout(n3474));
  jor  g03411(.dina(n3429), .dinb(n2553), .dout(n3475));
  jor  g03412(.dina(n3211), .dinb(n2629), .dout(n3476));
  jor  g03413(.dina(n3426), .dinb(n2738), .dout(n3477));
  jand g03414(.dina(n3477), .dinb(n3476), .dout(n3478));
  jand g03415(.dina(n3478), .dinb(n3475), .dout(n3479));
  jand g03416(.dina(n3479), .dinb(n3474), .dout(n3480));
  jxor g03417(.dina(n3480), .dinb(n3473), .dout(n3481));
  jand g03418(.dina(n3481), .dinb(n3472), .dout(n3482));
  jxor g03419(.dina(n2902), .dinb(n2901), .dout(n3483));
  jor  g03420(.dina(n3424), .dinb(n2768), .dout(n3484));
  jor  g03421(.dina(n3426), .dinb(n2553), .dout(n3485));
  jor  g03422(.dina(n3211), .dinb(n2428), .dout(n3486));
  jor  g03423(.dina(n3429), .dinb(n2629), .dout(n3487));
  jand g03424(.dina(n3487), .dinb(n3486), .dout(n3488));
  jand g03425(.dina(n3488), .dinb(n3485), .dout(n3489));
  jand g03426(.dina(n3489), .dinb(n3484), .dout(n3490));
  jxor g03427(.dina(n3490), .dinb(n3473), .dout(n3491));
  jand g03428(.dina(n3491), .dinb(n3483), .dout(n3492));
  jxor g03429(.dina(n2899), .dinb(n2898), .dout(n3493));
  jnot g03430(.din(n3493), .dout(n3494));
  jor  g03431(.dina(n3424), .dinb(n2779), .dout(n3495));
  jor  g03432(.dina(n3429), .dinb(n2428), .dout(n3496));
  jor  g03433(.dina(n3426), .dinb(n2629), .dout(n3497));
  jand g03434(.dina(n3497), .dinb(n3496), .dout(n3498));
  jor  g03435(.dina(n3211), .dinb(n2174), .dout(n3499));
  jand g03436(.dina(n3499), .dinb(n3498), .dout(n3500));
  jand g03437(.dina(n3500), .dinb(n3495), .dout(n3501));
  jxor g03438(.dina(n3501), .dinb(\a[14] ), .dout(n3502));
  jor  g03439(.dina(n3502), .dinb(n3494), .dout(n3503));
  jxor g03440(.dina(n2896), .dinb(n2895), .dout(n3504));
  jor  g03441(.dina(n3424), .dinb(n2430), .dout(n3505));
  jor  g03442(.dina(n3429), .dinb(n2174), .dout(n3506));
  jor  g03443(.dina(n3426), .dinb(n2428), .dout(n3507));
  jor  g03444(.dina(n3211), .dinb(n1954), .dout(n3508));
  jand g03445(.dina(n3508), .dinb(n3507), .dout(n3509));
  jand g03446(.dina(n3509), .dinb(n3506), .dout(n3510));
  jand g03447(.dina(n3510), .dinb(n3505), .dout(n3511));
  jxor g03448(.dina(n3511), .dinb(n3473), .dout(n3512));
  jand g03449(.dina(n3512), .dinb(n3504), .dout(n3513));
  jxor g03450(.dina(n2893), .dinb(n2892), .dout(n3514));
  jor  g03451(.dina(n3424), .dinb(n2176), .dout(n3515));
  jor  g03452(.dina(n3426), .dinb(n2174), .dout(n3516));
  jor  g03453(.dina(n3211), .dinb(n2057), .dout(n3517));
  jor  g03454(.dina(n3429), .dinb(n1954), .dout(n3518));
  jand g03455(.dina(n3518), .dinb(n3517), .dout(n3519));
  jand g03456(.dina(n3519), .dinb(n3516), .dout(n3520));
  jand g03457(.dina(n3520), .dinb(n3515), .dout(n3521));
  jxor g03458(.dina(n3521), .dinb(n3473), .dout(n3522));
  jand g03459(.dina(n3522), .dinb(n3514), .dout(n3523));
  jxor g03460(.dina(n2888), .dinb(n2887), .dout(n3524));
  jor  g03461(.dina(n3424), .dinb(n2197), .dout(n3525));
  jor  g03462(.dina(n3429), .dinb(n2057), .dout(n3526));
  jor  g03463(.dina(n3426), .dinb(n1954), .dout(n3527));
  jor  g03464(.dina(n3211), .dinb(n1790), .dout(n3528));
  jand g03465(.dina(n3528), .dinb(n3527), .dout(n3529));
  jand g03466(.dina(n3529), .dinb(n3526), .dout(n3530));
  jand g03467(.dina(n3530), .dinb(n3525), .dout(n3531));
  jxor g03468(.dina(n3531), .dinb(n3473), .dout(n3532));
  jand g03469(.dina(n3532), .dinb(n3524), .dout(n3533));
  jxor g03470(.dina(n2884), .dinb(n2876), .dout(n3534));
  jor  g03471(.dina(n3424), .dinb(n2208), .dout(n3535));
  jor  g03472(.dina(n3429), .dinb(n1790), .dout(n3536));
  jor  g03473(.dina(n3211), .dinb(n1606), .dout(n3537));
  jor  g03474(.dina(n3426), .dinb(n2057), .dout(n3538));
  jand g03475(.dina(n3538), .dinb(n3537), .dout(n3539));
  jand g03476(.dina(n3539), .dinb(n3536), .dout(n3540));
  jand g03477(.dina(n3540), .dinb(n3535), .dout(n3541));
  jxor g03478(.dina(n3541), .dinb(n3473), .dout(n3542));
  jand g03479(.dina(n3542), .dinb(n3534), .dout(n3543));
  jor  g03480(.dina(n3424), .dinb(n1792), .dout(n3544));
  jor  g03481(.dina(n3426), .dinb(n1790), .dout(n3545));
  jor  g03482(.dina(n3211), .dinb(n1448), .dout(n3546));
  jor  g03483(.dina(n3429), .dinb(n1606), .dout(n3547));
  jand g03484(.dina(n3547), .dinb(n3546), .dout(n3548));
  jand g03485(.dina(n3548), .dinb(n3545), .dout(n3549));
  jand g03486(.dina(n3549), .dinb(n3544), .dout(n3550));
  jxor g03487(.dina(n3550), .dinb(n3473), .dout(n3551));
  jor  g03488(.dina(n2863), .dinb(n2441), .dout(n3552));
  jxor g03489(.dina(n3552), .dinb(n2871), .dout(n3553));
  jand g03490(.dina(n3553), .dinb(n3551), .dout(n3554));
  jand g03491(.dina(n2860), .dinb(\a[17] ), .dout(n3555));
  jxor g03492(.dina(n3555), .dinb(n2858), .dout(n3556));
  jnot g03493(.din(n3556), .dout(n3557));
  jor  g03494(.dina(n3424), .dinb(n1608), .dout(n3558));
  jor  g03495(.dina(n3429), .dinb(n1448), .dout(n3559));
  jor  g03496(.dina(n3211), .dinb(n1255), .dout(n3560));
  jand g03497(.dina(n3560), .dinb(n3559), .dout(n3561));
  jor  g03498(.dina(n3426), .dinb(n1606), .dout(n3562));
  jand g03499(.dina(n3562), .dinb(n3561), .dout(n3563));
  jand g03500(.dina(n3563), .dinb(n3558), .dout(n3564));
  jxor g03501(.dina(n3564), .dinb(\a[14] ), .dout(n3565));
  jor  g03502(.dina(n3565), .dinb(n3557), .dout(n3566));
  jand g03503(.dina(n3423), .dinb(n728), .dout(n3567));
  jand g03504(.dina(n3428), .dinb(n438), .dout(n3568));
  jnot g03505(.din(n3426), .dout(n3569));
  jand g03506(.dina(n3569), .dinb(n795), .dout(n3570));
  jor  g03507(.dina(n3570), .dinb(n3568), .dout(n3571));
  jor  g03508(.dina(n3571), .dinb(n3567), .dout(n3572));
  jnot g03509(.din(n3572), .dout(n3573));
  jand g03510(.dina(n3205), .dinb(n438), .dout(n3574));
  jnot g03511(.din(n3574), .dout(n3575));
  jand g03512(.dina(n3575), .dinb(\a[14] ), .dout(n3576));
  jand g03513(.dina(n3576), .dinb(n3573), .dout(n3577));
  jand g03514(.dina(n3423), .dinb(n1639), .dout(n3578));
  jand g03515(.dina(n3428), .dinb(n795), .dout(n3579));
  jand g03516(.dina(n3569), .dinb(n1175), .dout(n3580));
  jor  g03517(.dina(n3580), .dinb(n3579), .dout(n3581));
  jand g03518(.dina(n3210), .dinb(n438), .dout(n3582));
  jor  g03519(.dina(n3582), .dinb(n3581), .dout(n3583));
  jor  g03520(.dina(n3583), .dinb(n3578), .dout(n3584));
  jnot g03521(.din(n3584), .dout(n3585));
  jand g03522(.dina(n3585), .dinb(n3577), .dout(n3586));
  jand g03523(.dina(n3586), .dinb(n2860), .dout(n3587));
  jnot g03524(.din(n3587), .dout(n3588));
  jxor g03525(.dina(n3586), .dinb(n2860), .dout(n3589));
  jnot g03526(.din(n3589), .dout(n3590));
  jor  g03527(.dina(n3424), .dinb(n1656), .dout(n3591));
  jor  g03528(.dina(n3426), .dinb(n1448), .dout(n3592));
  jor  g03529(.dina(n3429), .dinb(n1255), .dout(n3593));
  jand g03530(.dina(n3593), .dinb(n3592), .dout(n3594));
  jor  g03531(.dina(n3211), .dinb(n726), .dout(n3595));
  jand g03532(.dina(n3595), .dinb(n3594), .dout(n3596));
  jand g03533(.dina(n3596), .dinb(n3591), .dout(n3597));
  jxor g03534(.dina(n3597), .dinb(\a[14] ), .dout(n3598));
  jor  g03535(.dina(n3598), .dinb(n3590), .dout(n3599));
  jand g03536(.dina(n3599), .dinb(n3588), .dout(n3600));
  jnot g03537(.din(n3600), .dout(n3601));
  jxor g03538(.dina(n3565), .dinb(n3557), .dout(n3602));
  jand g03539(.dina(n3602), .dinb(n3601), .dout(n3603));
  jnot g03540(.din(n3603), .dout(n3604));
  jand g03541(.dina(n3604), .dinb(n3566), .dout(n3605));
  jnot g03542(.din(n3605), .dout(n3606));
  jxor g03543(.dina(n3553), .dinb(n3551), .dout(n3607));
  jand g03544(.dina(n3607), .dinb(n3606), .dout(n3608));
  jor  g03545(.dina(n3608), .dinb(n3554), .dout(n3609));
  jxor g03546(.dina(n3542), .dinb(n3534), .dout(n3610));
  jand g03547(.dina(n3610), .dinb(n3609), .dout(n3611));
  jor  g03548(.dina(n3611), .dinb(n3543), .dout(n3612));
  jxor g03549(.dina(n3532), .dinb(n3524), .dout(n3613));
  jand g03550(.dina(n3613), .dinb(n3612), .dout(n3614));
  jor  g03551(.dina(n3614), .dinb(n3533), .dout(n3615));
  jxor g03552(.dina(n3522), .dinb(n3514), .dout(n3616));
  jand g03553(.dina(n3616), .dinb(n3615), .dout(n3617));
  jor  g03554(.dina(n3617), .dinb(n3523), .dout(n3618));
  jxor g03555(.dina(n3512), .dinb(n3504), .dout(n3619));
  jand g03556(.dina(n3619), .dinb(n3618), .dout(n3620));
  jor  g03557(.dina(n3620), .dinb(n3513), .dout(n3621));
  jxor g03558(.dina(n3502), .dinb(n3494), .dout(n3622));
  jand g03559(.dina(n3622), .dinb(n3621), .dout(n3623));
  jnot g03560(.din(n3623), .dout(n3624));
  jand g03561(.dina(n3624), .dinb(n3503), .dout(n3625));
  jnot g03562(.din(n3625), .dout(n3626));
  jxor g03563(.dina(n3491), .dinb(n3483), .dout(n3627));
  jand g03564(.dina(n3627), .dinb(n3626), .dout(n3628));
  jor  g03565(.dina(n3628), .dinb(n3492), .dout(n3629));
  jxor g03566(.dina(n3481), .dinb(n3472), .dout(n3630));
  jand g03567(.dina(n3630), .dinb(n3629), .dout(n3631));
  jor  g03568(.dina(n3631), .dinb(n3482), .dout(n3632));
  jxor g03569(.dina(n3470), .dinb(n3462), .dout(n3633));
  jand g03570(.dina(n3633), .dinb(n3632), .dout(n3634));
  jnot g03571(.din(n3634), .dout(n3635));
  jand g03572(.dina(n3635), .dinb(n3471), .dout(n3636));
  jnot g03573(.din(n3636), .dout(n3637));
  jxor g03574(.dina(n3459), .dinb(n3450), .dout(n3638));
  jand g03575(.dina(n3638), .dinb(n3637), .dout(n3639));
  jnot g03576(.din(n3639), .dout(n3640));
  jand g03577(.dina(n3640), .dinb(n3460), .dout(n3641));
  jnot g03578(.din(n3641), .dout(n3642));
  jxor g03579(.dina(n3447), .dinb(n3438), .dout(n3643));
  jand g03580(.dina(n3643), .dinb(n3642), .dout(n3644));
  jnot g03581(.din(n3644), .dout(n3645));
  jand g03582(.dina(n3645), .dinb(n3448), .dout(n3646));
  jnot g03583(.din(n3646), .dout(n3647));
  jxor g03584(.dina(n3434), .dinb(n3091), .dout(n3648));
  jand g03585(.dina(n3648), .dinb(n3647), .dout(n3649));
  jor  g03586(.dina(n3649), .dinb(n3436), .dout(n3650));
  jor  g03587(.dina(n3088), .dinb(n2980), .dout(n3651));
  jand g03588(.dina(n3089), .dinb(n2922), .dout(n3652));
  jnot g03589(.din(n3652), .dout(n3653));
  jand g03590(.dina(n3653), .dinb(n3651), .dout(n3654));
  jnot g03591(.din(n3654), .dout(n3655));
  jor  g03592(.dina(n2977), .dinb(n2969), .dout(n3656));
  jand g03593(.dina(n2978), .dinb(n2925), .dout(n3657));
  jnot g03594(.din(n3657), .dout(n3658));
  jand g03595(.dina(n3658), .dinb(n3656), .dout(n3659));
  jnot g03596(.din(n3659), .dout(n3660));
  jand g03597(.dina(n2966), .dinb(n2958), .dout(n3661));
  jand g03598(.dina(n2967), .dinb(n2928), .dout(n3662));
  jor  g03599(.dina(n3662), .dinb(n3661), .dout(n3663));
  jor  g03600(.dina(n2956), .dinb(n2948), .dout(n3664));
  jand g03601(.dina(n2957), .dinb(n2934), .dout(n3665));
  jnot g03602(.din(n3665), .dout(n3666));
  jand g03603(.dina(n3666), .dinb(n3664), .dout(n3667));
  jnot g03604(.din(n3667), .dout(n3668));
  jor  g03605(.dina(n1790), .dinb(n2309), .dout(n3669));
  jor  g03606(.dina(n1792), .dinb(n2303), .dout(n3670));
  jor  g03607(.dina(n1805), .dinb(n1448), .dout(n3671));
  jor  g03608(.dina(n1606), .dinb(n2306), .dout(n3672));
  jand g03609(.dina(n3672), .dinb(n3671), .dout(n3673));
  jand g03610(.dina(n3673), .dinb(n3670), .dout(n3674));
  jand g03611(.dina(n3674), .dinb(n3669), .dout(n3675));
  jxor g03612(.dina(n3675), .dinb(\a[26] ), .dout(n3676));
  jnot g03613(.din(n3676), .dout(n3677));
  jand g03614(.dina(n2936), .dinb(n1639), .dout(n3678));
  jand g03615(.dina(n2940), .dinb(n795), .dout(n3679));
  jand g03616(.dina(n2943), .dinb(n1175), .dout(n3680));
  jor  g03617(.dina(n3680), .dinb(n3679), .dout(n3681));
  jor  g03618(.dina(n2939), .dinb(n64), .dout(n3682));
  jor  g03619(.dina(n3682), .dinb(n2942), .dout(n3683));
  jnot g03620(.din(n3683), .dout(n3684));
  jand g03621(.dina(n3684), .dinb(n438), .dout(n3685));
  jor  g03622(.dina(n3685), .dinb(n3681), .dout(n3686));
  jor  g03623(.dina(n3686), .dinb(n3678), .dout(n3687));
  jnot g03624(.din(n2946), .dout(n3688));
  jand g03625(.dina(n2299), .dinb(\a[29] ), .dout(n3689));
  jand g03626(.dina(n3689), .dinb(n3688), .dout(n3690));
  jnot g03627(.din(n3690), .dout(n3691));
  jand g03628(.dina(n3691), .dinb(\a[29] ), .dout(n3692));
  jxor g03629(.dina(n3692), .dinb(n3687), .dout(n3693));
  jxor g03630(.dina(n3693), .dinb(n3677), .dout(n3694));
  jxor g03631(.dina(n3694), .dinb(n3668), .dout(n3695));
  jnot g03632(.din(n3695), .dout(n3696));
  jor  g03633(.dina(n2174), .dinb(n1621), .dout(n3697));
  jor  g03634(.dina(n2176), .dinb(n807), .dout(n3698));
  jor  g03635(.dina(n2057), .dinb(n1617), .dout(n3699));
  jor  g03636(.dina(n1954), .dinb(n1613), .dout(n3700));
  jand g03637(.dina(n3700), .dinb(n3699), .dout(n3701));
  jand g03638(.dina(n3701), .dinb(n3698), .dout(n3702));
  jand g03639(.dina(n3702), .dinb(n3697), .dout(n3703));
  jxor g03640(.dina(n3703), .dinb(\a[23] ), .dout(n3704));
  jxor g03641(.dina(n3704), .dinb(n3696), .dout(n3705));
  jxor g03642(.dina(n3705), .dinb(n3663), .dout(n3706));
  jor  g03643(.dina(n2768), .dinb(n1820), .dout(n3707));
  jor  g03644(.dina(n2553), .dinb(n2189), .dout(n3708));
  jor  g03645(.dina(n2428), .dinb(n2186), .dout(n3709));
  jor  g03646(.dina(n2629), .dinb(n2181), .dout(n3710));
  jand g03647(.dina(n3710), .dinb(n3709), .dout(n3711));
  jand g03648(.dina(n3711), .dinb(n3708), .dout(n3712));
  jand g03649(.dina(n3712), .dinb(n3707), .dout(n3713));
  jxor g03650(.dina(n3713), .dinb(n2196), .dout(n3714));
  jxor g03651(.dina(n3714), .dinb(n3706), .dout(n3715));
  jxor g03652(.dina(n3715), .dinb(n3660), .dout(n3716));
  jnot g03653(.din(n3716), .dout(n3717));
  jor  g03654(.dina(n3451), .dinb(n2744), .dout(n3718));
  jor  g03655(.dina(n3072), .dinb(n2749), .dout(n3719));
  jor  g03656(.dina(n2758), .dinb(n2738), .dout(n3720));
  jand g03657(.dina(n3720), .dinb(n3719), .dout(n3721));
  jor  g03658(.dina(n3203), .dinb(n2753), .dout(n3722));
  jand g03659(.dina(n3722), .dinb(n3721), .dout(n3723));
  jand g03660(.dina(n3723), .dinb(n3718), .dout(n3724));
  jxor g03661(.dina(n3724), .dinb(\a[17] ), .dout(n3725));
  jxor g03662(.dina(n3725), .dinb(n3717), .dout(n3726));
  jxor g03663(.dina(n3726), .dinb(n3655), .dout(n3727));
  jnot g03664(.din(n3727), .dout(n3728));
  jnot g03665(.din(n3420), .dout(n3729));
  jand g03666(.dina(n3729), .dinb(n3287), .dout(n3730));
  jnot g03667(.din(n3730), .dout(n3731));
  jnot g03668(.din(n3421), .dout(n3732));
  jor  g03669(.dina(n3732), .dinb(n3305), .dout(n3733));
  jand g03670(.dina(n3733), .dinb(n3731), .dout(n3734));
  jand g03671(.dina(n2116), .dinb(n695), .dout(n3735));
  jand g03672(.dina(n982), .dinb(n135), .dout(n3736));
  jand g03673(.dina(n3736), .dinb(n691), .dout(n3737));
  jand g03674(.dina(n3737), .dinb(n666), .dout(n3738));
  jand g03675(.dina(n1867), .dinb(n1327), .dout(n3739));
  jand g03676(.dina(n3739), .dinb(n320), .dout(n3740));
  jand g03677(.dina(n3740), .dinb(n534), .dout(n3741));
  jand g03678(.dina(n3741), .dinb(n3367), .dout(n3742));
  jand g03679(.dina(n696), .dinb(n1292), .dout(n3743));
  jand g03680(.dina(n3743), .dinb(n2118), .dout(n3744));
  jand g03681(.dina(n3744), .dinb(n1451), .dout(n3745));
  jand g03682(.dina(n3745), .dinb(n3742), .dout(n3746));
  jnot g03683(.din(n356), .dout(n3747));
  jand g03684(.dina(n2409), .dinb(n3747), .dout(n3748));
  jand g03685(.dina(n3748), .dinb(n621), .dout(n3749));
  jnot g03686(.din(n1027), .dout(n3750));
  jand g03687(.dina(n1227), .dinb(n647), .dout(n3751));
  jand g03688(.dina(n495), .dinb(n1366), .dout(n3752));
  jand g03689(.dina(n3752), .dinb(n3751), .dout(n3753));
  jand g03690(.dina(n3753), .dinb(n3750), .dout(n3754));
  jand g03691(.dina(n3754), .dinb(n3749), .dout(n3755));
  jand g03692(.dina(n3755), .dinb(n3746), .dout(n3756));
  jand g03693(.dina(n3756), .dinb(n3738), .dout(n3757));
  jand g03694(.dina(n895), .dinb(n583), .dout(n3758));
  jand g03695(.dina(n3758), .dinb(n3757), .dout(n3759));
  jand g03696(.dina(n931), .dinb(n838), .dout(n3760));
  jand g03697(.dina(n3760), .dinb(n1756), .dout(n3761));
  jand g03698(.dina(n1511), .dinb(n833), .dout(n3762));
  jand g03699(.dina(n3762), .dinb(n3761), .dout(n3763));
  jand g03700(.dina(n3763), .dinb(n3759), .dout(n3764));
  jand g03701(.dina(n351), .dinb(n900), .dout(n3765));
  jand g03702(.dina(n3765), .dinb(n653), .dout(n3766));
  jand g03703(.dina(n1559), .dinb(n1682), .dout(n3767));
  jand g03704(.dina(n2023), .dinb(n1449), .dout(n3768));
  jand g03705(.dina(n3768), .dinb(n3767), .dout(n3769));
  jand g03706(.dina(n3769), .dinb(n3766), .dout(n3770));
  jand g03707(.dina(n1701), .dinb(n108), .dout(n3771));
  jand g03708(.dina(n3771), .dinb(n428), .dout(n3772));
  jand g03709(.dina(n3772), .dinb(n1237), .dout(n3773));
  jand g03710(.dina(n3773), .dinb(n3770), .dout(n3774));
  jand g03711(.dina(n3774), .dinb(n476), .dout(n3775));
  jand g03712(.dina(n1207), .dinb(n1375), .dout(n3776));
  jand g03713(.dina(n3776), .dinb(n1090), .dout(n3777));
  jand g03714(.dina(n3777), .dinb(n3184), .dout(n3778));
  jand g03715(.dina(n1583), .dinb(n1349), .dout(n3779));
  jand g03716(.dina(n2124), .dinb(n808), .dout(n3780));
  jand g03717(.dina(n3780), .dinb(n3779), .dout(n3781));
  jand g03718(.dina(n1846), .dinb(n1345), .dout(n3782));
  jand g03719(.dina(n3782), .dinb(n3781), .dout(n3783));
  jand g03720(.dina(n3783), .dinb(n3778), .dout(n3784));
  jand g03721(.dina(n3784), .dinb(n3775), .dout(n3785));
  jand g03722(.dina(n3785), .dinb(n3764), .dout(n3786));
  jand g03723(.dina(n3786), .dinb(n3735), .dout(n3787));
  jxor g03724(.dina(n3787), .dinb(n3420), .dout(n3788));
  jxor g03725(.dina(n3788), .dinb(n3734), .dout(n3789));
  jor  g03726(.dina(n3789), .dinb(n3424), .dout(n3790));
  jor  g03727(.dina(n3429), .dinb(n3420), .dout(n3791));
  jor  g03728(.dina(n3286), .dinb(n3211), .dout(n3792));
  jand g03729(.dina(n3792), .dinb(n3791), .dout(n3793));
  jor  g03730(.dina(n3787), .dinb(n3426), .dout(n3794));
  jand g03731(.dina(n3794), .dinb(n3793), .dout(n3795));
  jand g03732(.dina(n3795), .dinb(n3790), .dout(n3796));
  jxor g03733(.dina(n3796), .dinb(\a[14] ), .dout(n3797));
  jxor g03734(.dina(n3797), .dinb(n3728), .dout(n3798));
  jxor g03735(.dina(n3798), .dinb(n3650), .dout(n3799));
  jnot g03736(.din(n3799), .dout(n3800));
  jand g03737(.dina(n3316), .dinb(n1421), .dout(n3801));
  jand g03738(.dina(n1460), .dinb(n921), .dout(n3802));
  jand g03739(.dina(n3802), .dinb(n3801), .dout(n3803));
  jand g03740(.dina(n1228), .dinb(n1708), .dout(n3804));
  jand g03741(.dina(n1315), .dinb(n929), .dout(n3805));
  jand g03742(.dina(n3805), .dinb(n3804), .dout(n3806));
  jand g03743(.dina(n3806), .dinb(n3150), .dout(n3807));
  jand g03744(.dina(n838), .dinb(n82), .dout(n3808));
  jand g03745(.dina(n1682), .dinb(n1305), .dout(n3809));
  jand g03746(.dina(n3809), .dinb(n3808), .dout(n3810));
  jand g03747(.dina(n3810), .dinb(n3807), .dout(n3811));
  jand g03748(.dina(n349), .dinb(n1088), .dout(n3812));
  jand g03749(.dina(n3812), .dinb(n3811), .dout(n3813));
  jand g03750(.dina(n1449), .dinb(n130), .dout(n3814));
  jand g03751(.dina(n818), .dinb(n880), .dout(n3815));
  jand g03752(.dina(n3815), .dinb(n3814), .dout(n3816));
  jand g03753(.dina(n588), .dinb(n557), .dout(n3817));
  jand g03754(.dina(n3817), .dinb(n843), .dout(n3818));
  jand g03755(.dina(n1237), .dinb(n660), .dout(n3819));
  jand g03756(.dina(n3819), .dinb(n563), .dout(n3820));
  jand g03757(.dina(n1326), .dinb(n92), .dout(n3821));
  jand g03758(.dina(n3821), .dinb(n3820), .dout(n3822));
  jand g03759(.dina(n3822), .dinb(n3818), .dout(n3823));
  jand g03760(.dina(n3823), .dinb(n3816), .dout(n3824));
  jand g03761(.dina(n3824), .dinb(n3813), .dout(n3825));
  jand g03762(.dina(n3825), .dinb(n3803), .dout(n3826));
  jand g03763(.dina(n1107), .dinb(n1367), .dout(n3827));
  jand g03764(.dina(n3827), .dinb(n983), .dout(n3828));
  jand g03765(.dina(n1569), .dinb(n1346), .dout(n3829));
  jand g03766(.dina(n3829), .dinb(n1260), .dout(n3830));
  jand g03767(.dina(n3830), .dinb(n495), .dout(n3831));
  jand g03768(.dina(n3831), .dinb(n3828), .dout(n3832));
  jand g03769(.dina(n1205), .dinb(n122), .dout(n3833));
  jand g03770(.dina(n3833), .dinb(n1430), .dout(n3834));
  jand g03771(.dina(n672), .dinb(n621), .dout(n3835));
  jand g03772(.dina(n3835), .dinb(n1822), .dout(n3836));
  jand g03773(.dina(n3836), .dinb(n3834), .dout(n3837));
  jand g03774(.dina(n3837), .dinb(n3832), .dout(n3838));
  jand g03775(.dina(n2526), .dinb(n1516), .dout(n3839));
  jand g03776(.dina(n1511), .dinb(n2124), .dout(n3840));
  jand g03777(.dina(n833), .dinb(n703), .dout(n3841));
  jand g03778(.dina(n3841), .dinb(n3840), .dout(n3842));
  jand g03779(.dina(n2567), .dinb(n548), .dout(n3843));
  jand g03780(.dina(n3843), .dinb(n3842), .dout(n3844));
  jand g03781(.dina(n3844), .dinb(n3839), .dout(n3845));
  jand g03782(.dina(n3845), .dinb(n3838), .dout(n3846));
  jand g03783(.dina(n1778), .dinb(n456), .dout(n3847));
  jand g03784(.dina(n3847), .dinb(n179), .dout(n3848));
  jand g03785(.dina(n3848), .dinb(n919), .dout(n3849));
  jand g03786(.dina(n3255), .dinb(n653), .dout(n3850));
  jand g03787(.dina(n3850), .dinb(n3849), .dout(n3851));
  jand g03788(.dina(n1560), .dinb(n1465), .dout(n3852));
  jand g03789(.dina(n3264), .dinb(n2052), .dout(n3853));
  jand g03790(.dina(n3853), .dinb(n445), .dout(n3854));
  jand g03791(.dina(n3854), .dinb(n3852), .dout(n3855));
  jand g03792(.dina(n3855), .dinb(n3851), .dout(n3856));
  jand g03793(.dina(n948), .dinb(n1327), .dout(n3857));
  jand g03794(.dina(n3857), .dinb(n2388), .dout(n3858));
  jand g03795(.dina(n3858), .dinb(n1849), .dout(n3859));
  jand g03796(.dina(n3859), .dinb(n3856), .dout(n3860));
  jand g03797(.dina(n3860), .dinb(n3846), .dout(n3861));
  jand g03798(.dina(n3861), .dinb(n2679), .dout(n3862));
  jand g03799(.dina(n3862), .dinb(n3826), .dout(n3863));
  jxor g03800(.dina(\a[11] ), .dinb(\a[10] ), .dout(n3864));
  jxor g03801(.dina(\a[9] ), .dinb(\a[8] ), .dout(n3865));
  jnot g03802(.din(n3865), .dout(n3866));
  jxor g03803(.dina(\a[10] ), .dinb(\a[9] ), .dout(n3867));
  jnot g03804(.din(n3867), .dout(n3868));
  jand g03805(.dina(n3868), .dinb(n3866), .dout(n3869));
  jand g03806(.dina(n3869), .dinb(n3864), .dout(n3870));
  jnot g03807(.din(n3870), .dout(n3871));
  jor  g03808(.dina(n3871), .dinb(n3863), .dout(n3872));
  jnot g03809(.din(n3863), .dout(n3873));
  jand g03810(.dina(n2077), .dinb(n1189), .dout(n3874));
  jand g03811(.dina(n3874), .dinb(n3098), .dout(n3875));
  jand g03812(.dina(n3875), .dinb(n2566), .dout(n3876));
  jand g03813(.dina(n3876), .dinb(n1498), .dout(n3877));
  jand g03814(.dina(n2149), .dinb(n1697), .dout(n3878));
  jand g03815(.dina(n3878), .dinb(n647), .dout(n3879));
  jand g03816(.dina(n2106), .dinb(n699), .dout(n3880));
  jand g03817(.dina(n3747), .dinb(n1449), .dout(n3881));
  jand g03818(.dina(n3881), .dinb(n3880), .dout(n3882));
  jand g03819(.dina(n1037), .dinb(n447), .dout(n3883));
  jand g03820(.dina(n1351), .dinb(n916), .dout(n3884));
  jand g03821(.dina(n3884), .dinb(n3883), .dout(n3885));
  jand g03822(.dina(n2023), .dinb(n1822), .dout(n3886));
  jand g03823(.dina(n1575), .dinb(n1040), .dout(n3887));
  jand g03824(.dina(n3887), .dinb(n3886), .dout(n3888));
  jand g03825(.dina(n3888), .dinb(n3885), .dout(n3889));
  jand g03826(.dina(n3889), .dinb(n3882), .dout(n3890));
  jand g03827(.dina(n3890), .dinb(n3879), .dout(n3891));
  jand g03828(.dina(n2117), .dinb(n92), .dout(n3892));
  jand g03829(.dina(n3892), .dinb(n2343), .dout(n3893));
  jand g03830(.dina(n3893), .dinb(n1971), .dout(n3894));
  jand g03831(.dina(n3894), .dinb(n3891), .dout(n3895));
  jand g03832(.dina(n3895), .dinb(n3877), .dout(n3896));
  jand g03833(.dina(n588), .dinb(n555), .dout(n3897));
  jand g03834(.dina(n3897), .dinb(n3337), .dout(n3898));
  jand g03835(.dina(n3093), .dinb(n2012), .dout(n3899));
  jand g03836(.dina(n1096), .dinb(n662), .dout(n3900));
  jand g03837(.dina(n3900), .dinb(n1782), .dout(n3901));
  jand g03838(.dina(n3901), .dinb(n3899), .dout(n3902));
  jand g03839(.dina(n516), .dinb(n82), .dout(n3903));
  jand g03840(.dina(n3903), .dinb(n453), .dout(n3904));
  jand g03841(.dina(n3904), .dinb(n3902), .dout(n3905));
  jand g03842(.dina(n3905), .dinb(n3898), .dout(n3906));
  jand g03843(.dina(n1731), .dinb(n328), .dout(n3907));
  jand g03844(.dina(n3907), .dinb(n921), .dout(n3908));
  jand g03845(.dina(n2571), .dinb(n1228), .dout(n3909));
  jand g03846(.dina(n3909), .dinb(n3908), .dout(n3910));
  jand g03847(.dina(n1346), .dinb(n130), .dout(n3911));
  jand g03848(.dina(n3911), .dinb(n954), .dout(n3912));
  jand g03849(.dina(n1016), .dinb(n1366), .dout(n3913));
  jand g03850(.dina(n3913), .dinb(n266), .dout(n3914));
  jand g03851(.dina(n3914), .dinb(n3912), .dout(n3915));
  jand g03852(.dina(n3915), .dinb(n583), .dout(n3916));
  jand g03853(.dina(n3916), .dinb(n3910), .dout(n3917));
  jand g03854(.dina(n3917), .dinb(n3906), .dout(n3918));
  jand g03855(.dina(n670), .dinb(n1288), .dout(n3919));
  jand g03856(.dina(n3919), .dinb(n557), .dout(n3920));
  jand g03857(.dina(n320), .dinb(n132), .dout(n3921));
  jand g03858(.dina(n3921), .dinb(n3750), .dout(n3922));
  jand g03859(.dina(n3922), .dinb(n2082), .dout(n3923));
  jand g03860(.dina(n3923), .dinb(n586), .dout(n3924));
  jand g03861(.dina(n3924), .dinb(n3920), .dout(n3925));
  jand g03862(.dina(n3925), .dinb(n2734), .dout(n3926));
  jand g03863(.dina(n3926), .dinb(n3918), .dout(n3927));
  jand g03864(.dina(n3927), .dinb(n1406), .dout(n3928));
  jand g03865(.dina(n3928), .dinb(n3896), .dout(n3929));
  jnot g03866(.din(n3929), .dout(n3930));
  jand g03867(.dina(n3930), .dinb(n3873), .dout(n3931));
  jnot g03868(.din(n3931), .dout(n3932));
  jnot g03869(.din(n3787), .dout(n3933));
  jand g03870(.dina(n3873), .dinb(n3933), .dout(n3934));
  jnot g03871(.din(n3934), .dout(n3935));
  jand g03872(.dina(n3933), .dinb(n3729), .dout(n3936));
  jnot g03873(.din(n3936), .dout(n3937));
  jnot g03874(.din(n3788), .dout(n3938));
  jor  g03875(.dina(n3938), .dinb(n3734), .dout(n3939));
  jand g03876(.dina(n3939), .dinb(n3937), .dout(n3940));
  jxor g03877(.dina(n3863), .dinb(n3787), .dout(n3941));
  jnot g03878(.din(n3941), .dout(n3942));
  jor  g03879(.dina(n3942), .dinb(n3940), .dout(n3943));
  jand g03880(.dina(n3943), .dinb(n3935), .dout(n3944));
  jxor g03881(.dina(n3929), .dinb(n3863), .dout(n3945));
  jnot g03882(.din(n3945), .dout(n3946));
  jor  g03883(.dina(n3946), .dinb(n3944), .dout(n3947));
  jand g03884(.dina(n3947), .dinb(n3932), .dout(n3948));
  jand g03885(.dina(n1736), .dinb(n1233), .dout(n3949));
  jand g03886(.dina(n1721), .dinb(n492), .dout(n3950));
  jand g03887(.dina(n3950), .dinb(n1713), .dout(n3951));
  jand g03888(.dina(n3951), .dinb(n3949), .dout(n3952));
  jand g03889(.dina(n2597), .dinb(n175), .dout(n3953));
  jand g03890(.dina(n3953), .dinb(n718), .dout(n3954));
  jand g03891(.dina(n3857), .dinb(n3381), .dout(n3955));
  jand g03892(.dina(n1453), .dinb(n510), .dout(n3956));
  jand g03893(.dina(n3956), .dinb(n1451), .dout(n3957));
  jand g03894(.dina(n3957), .dinb(n3955), .dout(n3958));
  jand g03895(.dina(n3958), .dinb(n3954), .dout(n3959));
  jand g03896(.dina(n3959), .dinb(n3952), .dout(n3960));
  jnot g03897(.din(n710), .dout(n3961));
  jand g03898(.dina(n532), .dinb(n325), .dout(n3962));
  jand g03899(.dina(n3962), .dinb(n838), .dout(n3963));
  jand g03900(.dina(n978), .dinb(n873), .dout(n3964));
  jand g03901(.dina(n3964), .dinb(n3963), .dout(n3965));
  jand g03902(.dina(n3965), .dinb(n3961), .dout(n3966));
  jand g03903(.dina(n428), .dinb(n481), .dout(n3967));
  jand g03904(.dina(n3967), .dinb(n694), .dout(n3968));
  jand g03905(.dina(n3968), .dinb(n827), .dout(n3969));
  jand g03906(.dina(n3969), .dinb(n1580), .dout(n3970));
  jand g03907(.dina(n3970), .dinb(n3966), .dout(n3971));
  jand g03908(.dina(n3971), .dinb(n3960), .dout(n3972));
  jand g03909(.dina(n3972), .dinb(n3896), .dout(n3973));
  jnot g03910(.din(n942), .dout(n3974));
  jand g03911(.dina(n1053), .dinb(n1476), .dout(n3975));
  jand g03912(.dina(n3975), .dinb(n3974), .dout(n3976));
  jand g03913(.dina(n3976), .dinb(n621), .dout(n3977));
  jand g03914(.dina(n983), .dinb(n871), .dout(n3978));
  jand g03915(.dina(n3978), .dinb(n1245), .dout(n3979));
  jand g03916(.dina(n1005), .dinb(n954), .dout(n3980));
  jand g03917(.dina(n3980), .dinb(n2087), .dout(n3981));
  jand g03918(.dina(n3981), .dinb(n3979), .dout(n3982));
  jand g03919(.dina(n3982), .dinb(n3977), .dout(n3983));
  jand g03920(.dina(n2352), .dinb(n442), .dout(n3984));
  jand g03921(.dina(n1577), .dinb(n680), .dout(n3985));
  jand g03922(.dina(n3985), .dinb(n3984), .dout(n3986));
  jand g03923(.dina(n3986), .dinb(n1927), .dout(n3987));
  jand g03924(.dina(n3987), .dinb(n3983), .dout(n3988));
  jand g03925(.dina(n695), .dinb(n517), .dout(n3989));
  jand g03926(.dina(n700), .dinb(n461), .dout(n3990));
  jand g03927(.dina(n3990), .dinb(n3989), .dout(n3991));
  jand g03928(.dina(n917), .dinb(n1270), .dout(n3992));
  jand g03929(.dina(n3992), .dinb(n931), .dout(n3993));
  jand g03930(.dina(n3993), .dinb(n3991), .dout(n3994));
  jand g03931(.dina(n886), .dinb(n499), .dout(n3995));
  jand g03932(.dina(n1437), .dinb(n1344), .dout(n3996));
  jand g03933(.dina(n3996), .dinb(n3995), .dout(n3997));
  jand g03934(.dina(n3997), .dinb(n3994), .dout(n3998));
  jand g03935(.dina(n1016), .dinb(n121), .dout(n3999));
  jand g03936(.dina(n3999), .dinb(n1168), .dout(n4000));
  jand g03937(.dina(n4000), .dinb(n668), .dout(n4001));
  jand g03938(.dina(n4001), .dinb(n921), .dout(n4002));
  jand g03939(.dina(n4002), .dinb(n3998), .dout(n4003));
  jand g03940(.dina(n4003), .dinb(n3988), .dout(n4004));
  jand g03941(.dina(n1765), .dinb(n563), .dout(n4005));
  jand g03942(.dina(n870), .dinb(n1465), .dout(n4006));
  jand g03943(.dina(n1373), .dinb(n1315), .dout(n4007));
  jand g03944(.dina(n4007), .dinb(n456), .dout(n4008));
  jand g03945(.dina(n4008), .dinb(n548), .dout(n4009));
  jand g03946(.dina(n4009), .dinb(n4006), .dout(n4010));
  jand g03947(.dina(n3136), .dinb(n1162), .dout(n4011));
  jand g03948(.dina(n4011), .dinb(n1238), .dout(n4012));
  jand g03949(.dina(n844), .dinb(n480), .dout(n4013));
  jand g03950(.dina(n4013), .dinb(n1205), .dout(n4014));
  jand g03951(.dina(n4014), .dinb(n4012), .dout(n4015));
  jand g03952(.dina(n4015), .dinb(n4010), .dout(n4016));
  jand g03953(.dina(n4016), .dinb(n4005), .dout(n4017));
  jand g03954(.dina(n4017), .dinb(n4004), .dout(n4018));
  jand g03955(.dina(n4018), .dinb(n3973), .dout(n4019));
  jxor g03956(.dina(n4019), .dinb(n3929), .dout(n4020));
  jxor g03957(.dina(n4020), .dinb(n3948), .dout(n4021));
  jand g03958(.dina(n3865), .dinb(n3864), .dout(n4022));
  jnot g03959(.din(n4022), .dout(n4023));
  jor  g03960(.dina(n4023), .dinb(n4021), .dout(n4024));
  jor  g03961(.dina(n3866), .dinb(n3864), .dout(n4025));
  jor  g03962(.dina(n4025), .dinb(n4019), .dout(n4026));
  jand g03963(.dina(n3867), .dinb(n3866), .dout(n4027));
  jnot g03964(.din(n4027), .dout(n4028));
  jor  g03965(.dina(n4028), .dinb(n3929), .dout(n4029));
  jand g03966(.dina(n4029), .dinb(n4026), .dout(n4030));
  jand g03967(.dina(n4030), .dinb(n4024), .dout(n4031));
  jand g03968(.dina(n4031), .dinb(n3872), .dout(n4032));
  jxor g03969(.dina(n4032), .dinb(\a[11] ), .dout(n4033));
  jor  g03970(.dina(n4033), .dinb(n3800), .dout(n4034));
  jnot g03971(.din(n4034), .dout(n4035));
  jxor g03972(.dina(n3648), .dinb(n3647), .dout(n4036));
  jnot g03973(.din(n4036), .dout(n4037));
  jxor g03974(.dina(n3945), .dinb(n3944), .dout(n4038));
  jor  g03975(.dina(n4038), .dinb(n4023), .dout(n4039));
  jor  g03976(.dina(n4028), .dinb(n3863), .dout(n4040));
  jor  g03977(.dina(n4025), .dinb(n3929), .dout(n4041));
  jand g03978(.dina(n4041), .dinb(n4040), .dout(n4042));
  jor  g03979(.dina(n3871), .dinb(n3787), .dout(n4043));
  jand g03980(.dina(n4043), .dinb(n4042), .dout(n4044));
  jand g03981(.dina(n4044), .dinb(n4039), .dout(n4045));
  jxor g03982(.dina(n4045), .dinb(\a[11] ), .dout(n4046));
  jor  g03983(.dina(n4046), .dinb(n4037), .dout(n4047));
  jnot g03984(.din(n4047), .dout(n4048));
  jxor g03985(.dina(n3643), .dinb(n3642), .dout(n4049));
  jnot g03986(.din(\a[11] ), .dout(n4050));
  jxor g03987(.dina(n3941), .dinb(n3940), .dout(n4051));
  jor  g03988(.dina(n4051), .dinb(n4023), .dout(n4052));
  jor  g03989(.dina(n4028), .dinb(n3787), .dout(n4053));
  jor  g03990(.dina(n4025), .dinb(n3863), .dout(n4054));
  jor  g03991(.dina(n3871), .dinb(n3420), .dout(n4055));
  jand g03992(.dina(n4055), .dinb(n4054), .dout(n4056));
  jand g03993(.dina(n4056), .dinb(n4053), .dout(n4057));
  jand g03994(.dina(n4057), .dinb(n4052), .dout(n4058));
  jxor g03995(.dina(n4058), .dinb(n4050), .dout(n4059));
  jand g03996(.dina(n4059), .dinb(n4049), .dout(n4060));
  jxor g03997(.dina(n3638), .dinb(n3637), .dout(n4061));
  jnot g03998(.din(n4061), .dout(n4062));
  jor  g03999(.dina(n4023), .dinb(n3789), .dout(n4063));
  jor  g04000(.dina(n4028), .dinb(n3420), .dout(n4064));
  jor  g04001(.dina(n3871), .dinb(n3286), .dout(n4065));
  jand g04002(.dina(n4065), .dinb(n4064), .dout(n4066));
  jor  g04003(.dina(n4025), .dinb(n3787), .dout(n4067));
  jand g04004(.dina(n4067), .dinb(n4066), .dout(n4068));
  jand g04005(.dina(n4068), .dinb(n4063), .dout(n4069));
  jxor g04006(.dina(n4069), .dinb(\a[11] ), .dout(n4070));
  jor  g04007(.dina(n4070), .dinb(n4062), .dout(n4071));
  jnot g04008(.din(n4071), .dout(n4072));
  jxor g04009(.dina(n3633), .dinb(n3632), .dout(n4073));
  jnot g04010(.din(n4073), .dout(n4074));
  jor  g04011(.dina(n3871), .dinb(n3203), .dout(n4075));
  jor  g04012(.dina(n4023), .dinb(n3422), .dout(n4076));
  jor  g04013(.dina(n4025), .dinb(n3420), .dout(n4077));
  jor  g04014(.dina(n4028), .dinb(n3286), .dout(n4078));
  jand g04015(.dina(n4078), .dinb(n4077), .dout(n4079));
  jand g04016(.dina(n4079), .dinb(n4076), .dout(n4080));
  jand g04017(.dina(n4080), .dinb(n4075), .dout(n4081));
  jxor g04018(.dina(n4081), .dinb(\a[11] ), .dout(n4082));
  jor  g04019(.dina(n4082), .dinb(n4074), .dout(n4083));
  jnot g04020(.din(n4083), .dout(n4084));
  jxor g04021(.dina(n3630), .dinb(n3629), .dout(n4085));
  jor  g04022(.dina(n4023), .dinb(n3440), .dout(n4086));
  jor  g04023(.dina(n4028), .dinb(n3203), .dout(n4087));
  jor  g04024(.dina(n4025), .dinb(n3286), .dout(n4088));
  jor  g04025(.dina(n3871), .dinb(n3072), .dout(n4089));
  jand g04026(.dina(n4089), .dinb(n4088), .dout(n4090));
  jand g04027(.dina(n4090), .dinb(n4087), .dout(n4091));
  jand g04028(.dina(n4091), .dinb(n4086), .dout(n4092));
  jxor g04029(.dina(n4092), .dinb(n4050), .dout(n4093));
  jand g04030(.dina(n4093), .dinb(n4085), .dout(n4094));
  jxor g04031(.dina(n3627), .dinb(n3626), .dout(n4095));
  jnot g04032(.din(n4095), .dout(n4096));
  jor  g04033(.dina(n4023), .dinb(n3451), .dout(n4097));
  jor  g04034(.dina(n4028), .dinb(n3072), .dout(n4098));
  jor  g04035(.dina(n3871), .dinb(n2738), .dout(n4099));
  jand g04036(.dina(n4099), .dinb(n4098), .dout(n4100));
  jor  g04037(.dina(n4025), .dinb(n3203), .dout(n4101));
  jand g04038(.dina(n4101), .dinb(n4100), .dout(n4102));
  jand g04039(.dina(n4102), .dinb(n4097), .dout(n4103));
  jxor g04040(.dina(n4103), .dinb(\a[11] ), .dout(n4104));
  jor  g04041(.dina(n4104), .dinb(n4096), .dout(n4105));
  jnot g04042(.din(n4105), .dout(n4106));
  jxor g04043(.dina(n3622), .dinb(n3621), .dout(n4107));
  jnot g04044(.din(n4107), .dout(n4108));
  jor  g04045(.dina(n4023), .dinb(n3081), .dout(n4109));
  jor  g04046(.dina(n3871), .dinb(n2553), .dout(n4110));
  jor  g04047(.dina(n4028), .dinb(n2738), .dout(n4111));
  jand g04048(.dina(n4111), .dinb(n4110), .dout(n4112));
  jor  g04049(.dina(n4025), .dinb(n3072), .dout(n4113));
  jand g04050(.dina(n4113), .dinb(n4112), .dout(n4114));
  jand g04051(.dina(n4114), .dinb(n4109), .dout(n4115));
  jxor g04052(.dina(n4115), .dinb(\a[11] ), .dout(n4116));
  jor  g04053(.dina(n4116), .dinb(n4108), .dout(n4117));
  jxor g04054(.dina(n3619), .dinb(n3618), .dout(n4118));
  jnot g04055(.din(n4118), .dout(n4119));
  jor  g04056(.dina(n4023), .dinb(n2740), .dout(n4120));
  jor  g04057(.dina(n4028), .dinb(n2553), .dout(n4121));
  jor  g04058(.dina(n3871), .dinb(n2629), .dout(n4122));
  jand g04059(.dina(n4122), .dinb(n4121), .dout(n4123));
  jor  g04060(.dina(n4025), .dinb(n2738), .dout(n4124));
  jand g04061(.dina(n4124), .dinb(n4123), .dout(n4125));
  jand g04062(.dina(n4125), .dinb(n4120), .dout(n4126));
  jxor g04063(.dina(n4126), .dinb(\a[11] ), .dout(n4127));
  jor  g04064(.dina(n4127), .dinb(n4119), .dout(n4128));
  jxor g04065(.dina(n3616), .dinb(n3615), .dout(n4129));
  jor  g04066(.dina(n4023), .dinb(n2768), .dout(n4130));
  jor  g04067(.dina(n4025), .dinb(n2553), .dout(n4131));
  jor  g04068(.dina(n3871), .dinb(n2428), .dout(n4132));
  jor  g04069(.dina(n4028), .dinb(n2629), .dout(n4133));
  jand g04070(.dina(n4133), .dinb(n4132), .dout(n4134));
  jand g04071(.dina(n4134), .dinb(n4131), .dout(n4135));
  jand g04072(.dina(n4135), .dinb(n4130), .dout(n4136));
  jxor g04073(.dina(n4136), .dinb(n4050), .dout(n4137));
  jand g04074(.dina(n4137), .dinb(n4129), .dout(n4138));
  jnot g04075(.din(n4138), .dout(n4139));
  jxor g04076(.dina(n3613), .dinb(n3612), .dout(n4140));
  jor  g04077(.dina(n4023), .dinb(n2779), .dout(n4141));
  jor  g04078(.dina(n3871), .dinb(n2174), .dout(n4142));
  jor  g04079(.dina(n4025), .dinb(n2629), .dout(n4143));
  jor  g04080(.dina(n4028), .dinb(n2428), .dout(n4144));
  jand g04081(.dina(n4144), .dinb(n4143), .dout(n4145));
  jand g04082(.dina(n4145), .dinb(n4142), .dout(n4146));
  jand g04083(.dina(n4146), .dinb(n4141), .dout(n4147));
  jxor g04084(.dina(n4147), .dinb(n4050), .dout(n4148));
  jand g04085(.dina(n4148), .dinb(n4140), .dout(n4149));
  jnot g04086(.din(n4149), .dout(n4150));
  jxor g04087(.dina(n3610), .dinb(n3609), .dout(n4151));
  jor  g04088(.dina(n4023), .dinb(n2430), .dout(n4152));
  jor  g04089(.dina(n4028), .dinb(n2174), .dout(n4153));
  jor  g04090(.dina(n4025), .dinb(n2428), .dout(n4154));
  jor  g04091(.dina(n3871), .dinb(n1954), .dout(n4155));
  jand g04092(.dina(n4155), .dinb(n4154), .dout(n4156));
  jand g04093(.dina(n4156), .dinb(n4153), .dout(n4157));
  jand g04094(.dina(n4157), .dinb(n4152), .dout(n4158));
  jxor g04095(.dina(n4158), .dinb(n4050), .dout(n4159));
  jand g04096(.dina(n4159), .dinb(n4151), .dout(n4160));
  jnot g04097(.din(n4160), .dout(n4161));
  jxor g04098(.dina(n3607), .dinb(n3606), .dout(n4162));
  jnot g04099(.din(n4162), .dout(n4163));
  jor  g04100(.dina(n4023), .dinb(n2176), .dout(n4164));
  jor  g04101(.dina(n4028), .dinb(n1954), .dout(n4165));
  jor  g04102(.dina(n3871), .dinb(n2057), .dout(n4166));
  jand g04103(.dina(n4166), .dinb(n4165), .dout(n4167));
  jor  g04104(.dina(n4025), .dinb(n2174), .dout(n4168));
  jand g04105(.dina(n4168), .dinb(n4167), .dout(n4169));
  jand g04106(.dina(n4169), .dinb(n4164), .dout(n4170));
  jxor g04107(.dina(n4170), .dinb(\a[11] ), .dout(n4171));
  jor  g04108(.dina(n4171), .dinb(n4163), .dout(n4172));
  jxor g04109(.dina(n3602), .dinb(n3601), .dout(n4173));
  jnot g04110(.din(n4173), .dout(n4174));
  jor  g04111(.dina(n3871), .dinb(n1790), .dout(n4175));
  jor  g04112(.dina(n4023), .dinb(n2197), .dout(n4176));
  jor  g04113(.dina(n4025), .dinb(n1954), .dout(n4177));
  jor  g04114(.dina(n4028), .dinb(n2057), .dout(n4178));
  jand g04115(.dina(n4178), .dinb(n4177), .dout(n4179));
  jand g04116(.dina(n4179), .dinb(n4176), .dout(n4180));
  jand g04117(.dina(n4180), .dinb(n4175), .dout(n4181));
  jxor g04118(.dina(n4181), .dinb(\a[11] ), .dout(n4182));
  jor  g04119(.dina(n4182), .dinb(n4174), .dout(n4183));
  jxor g04120(.dina(n3598), .dinb(n3590), .dout(n4184));
  jor  g04121(.dina(n4023), .dinb(n2208), .dout(n4185));
  jor  g04122(.dina(n4028), .dinb(n1790), .dout(n4186));
  jor  g04123(.dina(n3871), .dinb(n1606), .dout(n4187));
  jor  g04124(.dina(n4025), .dinb(n2057), .dout(n4188));
  jand g04125(.dina(n4188), .dinb(n4187), .dout(n4189));
  jand g04126(.dina(n4189), .dinb(n4186), .dout(n4190));
  jand g04127(.dina(n4190), .dinb(n4185), .dout(n4191));
  jxor g04128(.dina(n4191), .dinb(n4050), .dout(n4192));
  jand g04129(.dina(n4192), .dinb(n4184), .dout(n4193));
  jor  g04130(.dina(n4025), .dinb(n1790), .dout(n4194));
  jor  g04131(.dina(n4023), .dinb(n1792), .dout(n4195));
  jor  g04132(.dina(n3871), .dinb(n1448), .dout(n4196));
  jor  g04133(.dina(n4028), .dinb(n1606), .dout(n4197));
  jand g04134(.dina(n4197), .dinb(n4196), .dout(n4198));
  jand g04135(.dina(n4198), .dinb(n4195), .dout(n4199));
  jand g04136(.dina(n4199), .dinb(n4194), .dout(n4200));
  jxor g04137(.dina(n4200), .dinb(\a[11] ), .dout(n4201));
  jnot g04138(.din(n4201), .dout(n4202));
  jor  g04139(.dina(n3577), .dinb(n3473), .dout(n4203));
  jxor g04140(.dina(n4203), .dinb(n3585), .dout(n4204));
  jand g04141(.dina(n4204), .dinb(n4202), .dout(n4205));
  jand g04142(.dina(n3574), .dinb(\a[14] ), .dout(n4206));
  jxor g04143(.dina(n4206), .dinb(n3572), .dout(n4207));
  jnot g04144(.din(n4207), .dout(n4208));
  jor  g04145(.dina(n4023), .dinb(n1608), .dout(n4209));
  jor  g04146(.dina(n4028), .dinb(n1448), .dout(n4210));
  jor  g04147(.dina(n3871), .dinb(n1255), .dout(n4211));
  jand g04148(.dina(n4211), .dinb(n4210), .dout(n4212));
  jor  g04149(.dina(n4025), .dinb(n1606), .dout(n4213));
  jand g04150(.dina(n4213), .dinb(n4212), .dout(n4214));
  jand g04151(.dina(n4214), .dinb(n4209), .dout(n4215));
  jxor g04152(.dina(n4215), .dinb(\a[11] ), .dout(n4216));
  jor  g04153(.dina(n4216), .dinb(n4208), .dout(n4217));
  jand g04154(.dina(n4022), .dinb(n728), .dout(n4218));
  jand g04155(.dina(n4027), .dinb(n438), .dout(n4219));
  jnot g04156(.din(n4025), .dout(n4220));
  jand g04157(.dina(n4220), .dinb(n795), .dout(n4221));
  jor  g04158(.dina(n4221), .dinb(n4219), .dout(n4222));
  jor  g04159(.dina(n4222), .dinb(n4218), .dout(n4223));
  jnot g04160(.din(n4223), .dout(n4224));
  jand g04161(.dina(n3865), .dinb(n438), .dout(n4225));
  jnot g04162(.din(n4225), .dout(n4226));
  jand g04163(.dina(n4226), .dinb(\a[11] ), .dout(n4227));
  jand g04164(.dina(n4227), .dinb(n4224), .dout(n4228));
  jand g04165(.dina(n4022), .dinb(n1639), .dout(n4229));
  jand g04166(.dina(n4027), .dinb(n795), .dout(n4230));
  jand g04167(.dina(n4220), .dinb(n1175), .dout(n4231));
  jor  g04168(.dina(n4231), .dinb(n4230), .dout(n4232));
  jand g04169(.dina(n3870), .dinb(n438), .dout(n4233));
  jor  g04170(.dina(n4233), .dinb(n4232), .dout(n4234));
  jor  g04171(.dina(n4234), .dinb(n4229), .dout(n4235));
  jnot g04172(.din(n4235), .dout(n4236));
  jand g04173(.dina(n4236), .dinb(n4228), .dout(n4237));
  jand g04174(.dina(n4237), .dinb(n3574), .dout(n4238));
  jnot g04175(.din(n4238), .dout(n4239));
  jxor g04176(.dina(n4237), .dinb(n3574), .dout(n4240));
  jnot g04177(.din(n4240), .dout(n4241));
  jor  g04178(.dina(n4023), .dinb(n1656), .dout(n4242));
  jor  g04179(.dina(n3871), .dinb(n726), .dout(n4243));
  jor  g04180(.dina(n4028), .dinb(n1255), .dout(n4244));
  jand g04181(.dina(n4244), .dinb(n4243), .dout(n4245));
  jor  g04182(.dina(n4025), .dinb(n1448), .dout(n4246));
  jand g04183(.dina(n4246), .dinb(n4245), .dout(n4247));
  jand g04184(.dina(n4247), .dinb(n4242), .dout(n4248));
  jxor g04185(.dina(n4248), .dinb(\a[11] ), .dout(n4249));
  jor  g04186(.dina(n4249), .dinb(n4241), .dout(n4250));
  jand g04187(.dina(n4250), .dinb(n4239), .dout(n4251));
  jnot g04188(.din(n4251), .dout(n4252));
  jxor g04189(.dina(n4216), .dinb(n4208), .dout(n4253));
  jand g04190(.dina(n4253), .dinb(n4252), .dout(n4254));
  jnot g04191(.din(n4254), .dout(n4255));
  jand g04192(.dina(n4255), .dinb(n4217), .dout(n4256));
  jnot g04193(.din(n4256), .dout(n4257));
  jxor g04194(.dina(n4204), .dinb(n4202), .dout(n4258));
  jand g04195(.dina(n4258), .dinb(n4257), .dout(n4259));
  jor  g04196(.dina(n4259), .dinb(n4205), .dout(n4260));
  jxor g04197(.dina(n4192), .dinb(n4184), .dout(n4261));
  jand g04198(.dina(n4261), .dinb(n4260), .dout(n4262));
  jor  g04199(.dina(n4262), .dinb(n4193), .dout(n4263));
  jxor g04200(.dina(n4182), .dinb(n4174), .dout(n4264));
  jand g04201(.dina(n4264), .dinb(n4263), .dout(n4265));
  jnot g04202(.din(n4265), .dout(n4266));
  jand g04203(.dina(n4266), .dinb(n4183), .dout(n4267));
  jnot g04204(.din(n4267), .dout(n4268));
  jxor g04205(.dina(n4171), .dinb(n4163), .dout(n4269));
  jand g04206(.dina(n4269), .dinb(n4268), .dout(n4270));
  jnot g04207(.din(n4270), .dout(n4271));
  jand g04208(.dina(n4271), .dinb(n4172), .dout(n4272));
  jxor g04209(.dina(n4159), .dinb(n4151), .dout(n4273));
  jnot g04210(.din(n4273), .dout(n4274));
  jor  g04211(.dina(n4274), .dinb(n4272), .dout(n4275));
  jand g04212(.dina(n4275), .dinb(n4161), .dout(n4276));
  jxor g04213(.dina(n4148), .dinb(n4140), .dout(n4277));
  jnot g04214(.din(n4277), .dout(n4278));
  jor  g04215(.dina(n4278), .dinb(n4276), .dout(n4279));
  jand g04216(.dina(n4279), .dinb(n4150), .dout(n4280));
  jxor g04217(.dina(n4137), .dinb(n4129), .dout(n4281));
  jnot g04218(.din(n4281), .dout(n4282));
  jor  g04219(.dina(n4282), .dinb(n4280), .dout(n4283));
  jand g04220(.dina(n4283), .dinb(n4139), .dout(n4284));
  jxor g04221(.dina(n4127), .dinb(n4119), .dout(n4285));
  jnot g04222(.din(n4285), .dout(n4286));
  jor  g04223(.dina(n4286), .dinb(n4284), .dout(n4287));
  jand g04224(.dina(n4287), .dinb(n4128), .dout(n4288));
  jxor g04225(.dina(n4116), .dinb(n4108), .dout(n4289));
  jnot g04226(.din(n4289), .dout(n4290));
  jor  g04227(.dina(n4290), .dinb(n4288), .dout(n4291));
  jand g04228(.dina(n4291), .dinb(n4117), .dout(n4292));
  jnot g04229(.din(n4292), .dout(n4293));
  jxor g04230(.dina(n4104), .dinb(n4096), .dout(n4294));
  jand g04231(.dina(n4294), .dinb(n4293), .dout(n4295));
  jor  g04232(.dina(n4295), .dinb(n4106), .dout(n4296));
  jxor g04233(.dina(n4093), .dinb(n4085), .dout(n4297));
  jand g04234(.dina(n4297), .dinb(n4296), .dout(n4298));
  jor  g04235(.dina(n4298), .dinb(n4094), .dout(n4299));
  jxor g04236(.dina(n4082), .dinb(n4074), .dout(n4300));
  jand g04237(.dina(n4300), .dinb(n4299), .dout(n4301));
  jor  g04238(.dina(n4301), .dinb(n4084), .dout(n4302));
  jxor g04239(.dina(n4070), .dinb(n4062), .dout(n4303));
  jand g04240(.dina(n4303), .dinb(n4302), .dout(n4304));
  jor  g04241(.dina(n4304), .dinb(n4072), .dout(n4305));
  jxor g04242(.dina(n4059), .dinb(n4049), .dout(n4306));
  jand g04243(.dina(n4306), .dinb(n4305), .dout(n4307));
  jor  g04244(.dina(n4307), .dinb(n4060), .dout(n4308));
  jxor g04245(.dina(n4046), .dinb(n4036), .dout(n4309));
  jnot g04246(.din(n4309), .dout(n4310));
  jand g04247(.dina(n4310), .dinb(n4308), .dout(n4311));
  jor  g04248(.dina(n4311), .dinb(n4048), .dout(n4312));
  jxor g04249(.dina(n4033), .dinb(n3799), .dout(n4313));
  jnot g04250(.din(n4313), .dout(n4314));
  jand g04251(.dina(n4314), .dinb(n4312), .dout(n4315));
  jor  g04252(.dina(n4315), .dinb(n4035), .dout(n4316));
  jor  g04253(.dina(n3797), .dinb(n3728), .dout(n4317));
  jnot g04254(.din(n4317), .dout(n4318));
  jand g04255(.dina(n3798), .dinb(n3650), .dout(n4319));
  jor  g04256(.dina(n4319), .dinb(n4318), .dout(n4320));
  jor  g04257(.dina(n3725), .dinb(n3717), .dout(n4321));
  jand g04258(.dina(n3726), .dinb(n3655), .dout(n4322));
  jnot g04259(.din(n4322), .dout(n4323));
  jand g04260(.dina(n4323), .dinb(n4321), .dout(n4324));
  jnot g04261(.din(n4324), .dout(n4325));
  jand g04262(.dina(n3714), .dinb(n3706), .dout(n4326));
  jand g04263(.dina(n3715), .dinb(n3660), .dout(n4327));
  jor  g04264(.dina(n4327), .dinb(n4326), .dout(n4328));
  jor  g04265(.dina(n3704), .dinb(n3696), .dout(n4329));
  jand g04266(.dina(n3705), .dinb(n3663), .dout(n4330));
  jnot g04267(.din(n4330), .dout(n4331));
  jand g04268(.dina(n4331), .dinb(n4329), .dout(n4332));
  jnot g04269(.din(n4332), .dout(n4333));
  jand g04270(.dina(n3693), .dinb(n3677), .dout(n4334));
  jand g04271(.dina(n3694), .dinb(n3668), .dout(n4335));
  jor  g04272(.dina(n4335), .dinb(n4334), .dout(n4336));
  jxor g04273(.dina(\a[30] ), .dinb(n93), .dout(n4337));
  jnot g04274(.din(n4337), .dout(n4338));
  jand g04275(.dina(n4338), .dinb(n438), .dout(n4339));
  jor  g04276(.dina(n3691), .dinb(n3687), .dout(n4340));
  jnot g04277(.din(n4340), .dout(n4341));
  jxor g04278(.dina(n4341), .dinb(n4339), .dout(n4342));
  jnot g04279(.din(n2936), .dout(n4343));
  jor  g04280(.dina(n4343), .dinb(n1656), .dout(n4344));
  jor  g04281(.dina(n3683), .dinb(n726), .dout(n4345));
  jnot g04282(.din(n2940), .dout(n4346));
  jor  g04283(.dina(n4346), .dinb(n1255), .dout(n4347));
  jnot g04284(.din(n2943), .dout(n4348));
  jor  g04285(.dina(n4348), .dinb(n1448), .dout(n4349));
  jand g04286(.dina(n4349), .dinb(n4347), .dout(n4350));
  jand g04287(.dina(n4350), .dinb(n4345), .dout(n4351));
  jand g04288(.dina(n4351), .dinb(n4344), .dout(n4352));
  jxor g04289(.dina(n4352), .dinb(n93), .dout(n4353));
  jxor g04290(.dina(n4353), .dinb(n4342), .dout(n4354));
  jor  g04291(.dina(n2208), .dinb(n2303), .dout(n4355));
  jor  g04292(.dina(n1790), .dinb(n2306), .dout(n4356));
  jor  g04293(.dina(n1805), .dinb(n1606), .dout(n4357));
  jor  g04294(.dina(n2057), .dinb(n2309), .dout(n4358));
  jand g04295(.dina(n4358), .dinb(n4357), .dout(n4359));
  jand g04296(.dina(n4359), .dinb(n4356), .dout(n4360));
  jand g04297(.dina(n4360), .dinb(n4355), .dout(n4361));
  jxor g04298(.dina(n4361), .dinb(n77), .dout(n4362));
  jxor g04299(.dina(n4362), .dinb(n4354), .dout(n4363));
  jxor g04300(.dina(n4363), .dinb(n4336), .dout(n4364));
  jor  g04301(.dina(n2430), .dinb(n807), .dout(n4365));
  jor  g04302(.dina(n2174), .dinb(n1613), .dout(n4366));
  jor  g04303(.dina(n2428), .dinb(n1621), .dout(n4367));
  jor  g04304(.dina(n1954), .dinb(n1617), .dout(n4368));
  jand g04305(.dina(n4368), .dinb(n4367), .dout(n4369));
  jand g04306(.dina(n4369), .dinb(n4366), .dout(n4370));
  jand g04307(.dina(n4370), .dinb(n4365), .dout(n4371));
  jxor g04308(.dina(n4371), .dinb(n65), .dout(n4372));
  jxor g04309(.dina(n4372), .dinb(n4364), .dout(n4373));
  jxor g04310(.dina(n4373), .dinb(n4333), .dout(n4374));
  jor  g04311(.dina(n2740), .dinb(n1820), .dout(n4375));
  jor  g04312(.dina(n2553), .dinb(n2181), .dout(n4376));
  jor  g04313(.dina(n2629), .dinb(n2186), .dout(n4377));
  jor  g04314(.dina(n2738), .dinb(n2189), .dout(n4378));
  jand g04315(.dina(n4378), .dinb(n4377), .dout(n4379));
  jand g04316(.dina(n4379), .dinb(n4376), .dout(n4380));
  jand g04317(.dina(n4380), .dinb(n4375), .dout(n4381));
  jxor g04318(.dina(n4381), .dinb(n2196), .dout(n4382));
  jxor g04319(.dina(n4382), .dinb(n4374), .dout(n4383));
  jxor g04320(.dina(n4383), .dinb(n4328), .dout(n4384));
  jnot g04321(.din(n4384), .dout(n4385));
  jor  g04322(.dina(n3440), .dinb(n2744), .dout(n4386));
  jor  g04323(.dina(n3203), .dinb(n2749), .dout(n4387));
  jor  g04324(.dina(n3286), .dinb(n2753), .dout(n4388));
  jand g04325(.dina(n4388), .dinb(n4387), .dout(n4389));
  jor  g04326(.dina(n3072), .dinb(n2758), .dout(n4390));
  jand g04327(.dina(n4390), .dinb(n4389), .dout(n4391));
  jand g04328(.dina(n4391), .dinb(n4386), .dout(n4392));
  jxor g04329(.dina(n4392), .dinb(\a[17] ), .dout(n4393));
  jxor g04330(.dina(n4393), .dinb(n4385), .dout(n4394));
  jxor g04331(.dina(n4394), .dinb(n4325), .dout(n4395));
  jor  g04332(.dina(n4051), .dinb(n3424), .dout(n4396));
  jor  g04333(.dina(n3787), .dinb(n3429), .dout(n4397));
  jor  g04334(.dina(n3863), .dinb(n3426), .dout(n4398));
  jor  g04335(.dina(n3420), .dinb(n3211), .dout(n4399));
  jand g04336(.dina(n4399), .dinb(n4398), .dout(n4400));
  jand g04337(.dina(n4400), .dinb(n4397), .dout(n4401));
  jand g04338(.dina(n4401), .dinb(n4396), .dout(n4402));
  jxor g04339(.dina(n4402), .dinb(n3473), .dout(n4403));
  jxor g04340(.dina(n4403), .dinb(n4395), .dout(n4404));
  jxor g04341(.dina(n4404), .dinb(n4320), .dout(n4405));
  jnot g04342(.din(n4019), .dout(n4406));
  jand g04343(.dina(n4406), .dinb(n3930), .dout(n4407));
  jnot g04344(.din(n4407), .dout(n4408));
  jnot g04345(.din(n4020), .dout(n4409));
  jor  g04346(.dina(n4409), .dinb(n3948), .dout(n4410));
  jand g04347(.dina(n4410), .dinb(n4408), .dout(n4411));
  jand g04348(.dina(n1203), .dinb(n1575), .dout(n4412));
  jand g04349(.dina(n4412), .dinb(n678), .dout(n4413));
  jand g04350(.dina(n886), .dinb(n662), .dout(n4414));
  jand g04351(.dina(n4414), .dinb(n880), .dout(n4415));
  jand g04352(.dina(n4415), .dinb(n4413), .dout(n4416));
  jand g04353(.dina(n1532), .dinb(n171), .dout(n4417));
  jand g04354(.dina(n1351), .dinb(n683), .dout(n4418));
  jand g04355(.dina(n4418), .dinb(n4417), .dout(n4419));
  jand g04356(.dina(n4419), .dinb(n4416), .dout(n4420));
  jand g04357(.dina(n4420), .dinb(n1561), .dout(n4421));
  jand g04358(.dina(n600), .dinb(n454), .dout(n4422));
  jand g04359(.dina(n4422), .dinb(n3178), .dout(n4423));
  jand g04360(.dina(n1536), .dinb(n1470), .dout(n4424));
  jand g04361(.dina(n516), .dinb(n108), .dout(n4425));
  jand g04362(.dina(n4425), .dinb(n4424), .dout(n4426));
  jand g04363(.dina(n4426), .dinb(n816), .dout(n4427));
  jand g04364(.dina(n1316), .dinb(n1205), .dout(n4428));
  jand g04365(.dina(n4428), .dinb(n931), .dout(n4429));
  jand g04366(.dina(n1017), .dinb(n694), .dout(n4430));
  jand g04367(.dina(n4430), .dinb(n4429), .dout(n4431));
  jand g04368(.dina(n4431), .dinb(n4427), .dout(n4432));
  jand g04369(.dina(n4432), .dinb(n4423), .dout(n4433));
  jand g04370(.dina(n3908), .dinb(n1324), .dout(n4434));
  jand g04371(.dina(n700), .dinb(n650), .dout(n4435));
  jand g04372(.dina(n1534), .dinb(n1088), .dout(n4436));
  jand g04373(.dina(n4436), .dinb(n1426), .dout(n4437));
  jand g04374(.dina(n4437), .dinb(n4435), .dout(n4438));
  jand g04375(.dina(n4438), .dinb(n4434), .dout(n4439));
  jand g04376(.dina(n645), .dinb(n1373), .dout(n4440));
  jand g04377(.dina(n713), .dinb(n542), .dout(n4441));
  jand g04378(.dina(n4441), .dinb(n1459), .dout(n4442));
  jand g04379(.dina(n4442), .dinb(n4440), .dout(n4443));
  jand g04380(.dina(n1851), .dinb(n1308), .dout(n4444));
  jand g04381(.dina(n4444), .dinb(n4443), .dout(n4445));
  jand g04382(.dina(n4445), .dinb(n4439), .dout(n4446));
  jand g04383(.dina(n4446), .dinb(n4433), .dout(n4447));
  jand g04384(.dina(n965), .dinb(n501), .dout(n4448));
  jand g04385(.dina(n4448), .dinb(n1697), .dout(n4449));
  jand g04386(.dina(n4449), .dinb(n1212), .dout(n4450));
  jand g04387(.dina(n1163), .dinb(n1453), .dout(n4451));
  jand g04388(.dina(n811), .dinb(n168), .dout(n4452));
  jand g04389(.dina(n4452), .dinb(n993), .dout(n4453));
  jand g04390(.dina(n4453), .dinb(n4451), .dout(n4454));
  jand g04391(.dina(n4454), .dinb(n4450), .dout(n4455));
  jand g04392(.dina(n3003), .dinb(n2124), .dout(n4456));
  jand g04393(.dina(n4456), .dinb(n266), .dout(n4457));
  jand g04394(.dina(n1090), .dinb(n824), .dout(n4458));
  jand g04395(.dina(n4458), .dinb(n3405), .dout(n4459));
  jand g04396(.dina(n4459), .dinb(n4457), .dout(n4460));
  jand g04397(.dina(n3026), .dinb(n654), .dout(n4461));
  jand g04398(.dina(n1713), .dinb(n900), .dout(n4462));
  jand g04399(.dina(n4462), .dinb(n3978), .dout(n4463));
  jand g04400(.dina(n4463), .dinb(n4461), .dout(n4464));
  jand g04401(.dina(n3897), .dinb(n1043), .dout(n4465));
  jand g04402(.dina(n4465), .dinb(n4464), .dout(n4466));
  jand g04403(.dina(n4466), .dinb(n4460), .dout(n4467));
  jand g04404(.dina(n4467), .dinb(n4455), .dout(n4468));
  jand g04405(.dina(n4468), .dinb(n4447), .dout(n4469));
  jand g04406(.dina(n4469), .dinb(n2707), .dout(n4470));
  jand g04407(.dina(n4470), .dinb(n4421), .dout(n4471));
  jxor g04408(.dina(n4471), .dinb(n4019), .dout(n4472));
  jxor g04409(.dina(n4472), .dinb(n4411), .dout(n4473));
  jor  g04410(.dina(n4473), .dinb(n4023), .dout(n4474));
  jor  g04411(.dina(n4028), .dinb(n4019), .dout(n4475));
  jor  g04412(.dina(n3929), .dinb(n3871), .dout(n4476));
  jor  g04413(.dina(n4471), .dinb(n4025), .dout(n4477));
  jand g04414(.dina(n4477), .dinb(n4476), .dout(n4478));
  jand g04415(.dina(n4478), .dinb(n4475), .dout(n4479));
  jand g04416(.dina(n4479), .dinb(n4474), .dout(n4480));
  jxor g04417(.dina(n4480), .dinb(n4050), .dout(n4481));
  jxor g04418(.dina(n4481), .dinb(n4405), .dout(n4482));
  jxor g04419(.dina(n4482), .dinb(n4316), .dout(n4483));
  jnot g04420(.din(n4483), .dout(n4484));
  jand g04421(.dina(n2144), .dinb(n1456), .dout(n4485));
  jand g04422(.dina(n4485), .dinb(n814), .dout(n4486));
  jand g04423(.dina(n1515), .dinb(n1437), .dout(n4487));
  jand g04424(.dina(n4487), .dinb(n1228), .dout(n4488));
  jand g04425(.dina(n4488), .dinb(n653), .dout(n4489));
  jand g04426(.dina(n1536), .dinb(n1304), .dout(n4490));
  jand g04427(.dina(n4490), .dinb(n3324), .dout(n4491));
  jand g04428(.dina(n1928), .dinb(n1283), .dout(n4492));
  jand g04429(.dina(n4492), .dinb(n4491), .dout(n4493));
  jand g04430(.dina(n4493), .dinb(n4489), .dout(n4494));
  jand g04431(.dina(n1346), .dinb(n1334), .dout(n4495));
  jand g04432(.dina(n4495), .dinb(n440), .dout(n4496));
  jand g04433(.dina(n4496), .dinb(n2587), .dout(n4497));
  jand g04434(.dina(n1247), .dinb(n1042), .dout(n4498));
  jand g04435(.dina(n4498), .dinb(n4497), .dout(n4499));
  jand g04436(.dina(n4499), .dinb(n4494), .dout(n4500));
  jand g04437(.dina(n3178), .dinb(n328), .dout(n4501));
  jand g04438(.dina(n886), .dinb(n1238), .dout(n4502));
  jand g04439(.dina(n4502), .dinb(n463), .dout(n4503));
  jand g04440(.dina(n4503), .dinb(n4501), .dout(n4504));
  jand g04441(.dina(n4504), .dinb(n3258), .dout(n4505));
  jand g04442(.dina(n4505), .dinb(n4500), .dout(n4506));
  jand g04443(.dina(n4506), .dinb(n4486), .dout(n4507));
  jand g04444(.dina(n1397), .dinb(n1233), .dout(n4508));
  jand g04445(.dina(n4508), .dinb(n3749), .dout(n4509));
  jand g04446(.dina(n4509), .dinb(n4507), .dout(n4510));
  jand g04447(.dina(n1219), .dinb(n541), .dout(n4511));
  jand g04448(.dina(n1460), .dinb(n1682), .dout(n4512));
  jand g04449(.dina(n4512), .dinb(n4511), .dout(n4513));
  jand g04450(.dina(n1189), .dinb(n1541), .dout(n4514));
  jand g04451(.dina(n4514), .dinb(n1575), .dout(n4515));
  jand g04452(.dina(n4515), .dinb(n4513), .dout(n4516));
  jand g04453(.dina(n1203), .dinb(n175), .dout(n4517));
  jand g04454(.dina(n4517), .dinb(n600), .dout(n4518));
  jand g04455(.dina(n4518), .dinb(n1476), .dout(n4519));
  jand g04456(.dina(n4519), .dinb(n4516), .dout(n4520));
  jand g04457(.dina(n3103), .dinb(n693), .dout(n4521));
  jand g04458(.dina(n4521), .dinb(n1205), .dout(n4522));
  jand g04459(.dina(n4522), .dinb(n3906), .dout(n4523));
  jand g04460(.dina(n4523), .dinb(n4520), .dout(n4524));
  jand g04461(.dina(n4524), .dinb(n1425), .dout(n4525));
  jand g04462(.dina(n4525), .dinb(n4510), .dout(n4526));
  jnot g04463(.din(n4526), .dout(n4527));
  jand g04464(.dina(n2500), .dinb(n1036), .dout(n4528));
  jand g04465(.dina(n4528), .dinb(n1916), .dout(n4529));
  jand g04466(.dina(n454), .dinb(n92), .dout(n4530));
  jand g04467(.dina(n4530), .dinb(n1682), .dout(n4531));
  jand g04468(.dina(n1042), .dinb(n1378), .dout(n4532));
  jand g04469(.dina(n4532), .dinb(n4531), .dout(n4533));
  jand g04470(.dina(n929), .dinb(n1429), .dout(n4534));
  jand g04471(.dina(n4534), .dinb(n551), .dout(n4535));
  jand g04472(.dina(n4535), .dinb(n1823), .dout(n4536));
  jand g04473(.dina(n4536), .dinb(n4533), .dout(n4537));
  jand g04474(.dina(n3978), .dinb(n988), .dout(n4538));
  jand g04475(.dina(n4538), .dinb(n4537), .dout(n4539));
  jand g04476(.dina(n4539), .dinb(n4529), .dout(n4540));
  jand g04477(.dina(n1536), .dinb(n833), .dout(n4541));
  jand g04478(.dina(n4522), .dinb(n2124), .dout(n4542));
  jand g04479(.dina(n4542), .dinb(n4541), .dout(n4543));
  jand g04480(.dina(n1767), .dinb(n1561), .dout(n4544));
  jand g04481(.dina(n715), .dinb(n172), .dout(n4545));
  jand g04482(.dina(n4545), .dinb(n1366), .dout(n4546));
  jand g04483(.dina(n4546), .dinb(n4544), .dout(n4547));
  jand g04484(.dina(n1580), .dinb(n1226), .dout(n4548));
  jand g04485(.dina(n4548), .dinb(n1773), .dout(n4549));
  jand g04486(.dina(n4549), .dinb(n4547), .dout(n4550));
  jand g04487(.dina(n4550), .dinb(n1458), .dout(n4551));
  jand g04488(.dina(n4551), .dinb(n4543), .dout(n4552));
  jand g04489(.dina(n4552), .dinb(n4540), .dout(n4553));
  jand g04490(.dina(n818), .dinb(n893), .dout(n4554));
  jand g04491(.dina(n1016), .dinb(n465), .dout(n4555));
  jand g04492(.dina(n4555), .dinb(n4554), .dout(n4556));
  jand g04493(.dina(n1005), .dinb(n469), .dout(n4557));
  jand g04494(.dina(n4557), .dinb(n4556), .dout(n4558));
  jand g04495(.dina(n2449), .dinb(n2345), .dout(n4559));
  jand g04496(.dina(n4559), .dinb(n4558), .dout(n4560));
  jand g04497(.dina(n1721), .dinb(n1246), .dout(n4561));
  jand g04498(.dina(n981), .dinb(n621), .dout(n4562));
  jand g04499(.dina(n4562), .dinb(n843), .dout(n4563));
  jand g04500(.dina(n4563), .dinb(n933), .dout(n4564));
  jand g04501(.dina(n4564), .dinb(n4561), .dout(n4565));
  jand g04502(.dina(n4565), .dinb(n4560), .dout(n4566));
  jand g04503(.dina(n1090), .dinb(n696), .dout(n4567));
  jand g04504(.dina(n4567), .dinb(n563), .dout(n4568));
  jand g04505(.dina(n4568), .dinb(n1162), .dout(n4569));
  jand g04506(.dina(n4569), .dinb(n4566), .dout(n4570));
  jand g04507(.dina(n4570), .dinb(n2152), .dout(n4571));
  jand g04508(.dina(n1167), .dinb(n542), .dout(n4572));
  jand g04509(.dina(n4572), .dinb(n2570), .dout(n4573));
  jand g04510(.dina(n869), .dinb(n1756), .dout(n4574));
  jand g04511(.dina(n1437), .dinb(n954), .dout(n4575));
  jand g04512(.dina(n4575), .dinb(n4574), .dout(n4576));
  jand g04513(.dina(n4576), .dinb(n2483), .dout(n4577));
  jand g04514(.dina(n2406), .dinb(n1283), .dout(n4578));
  jand g04515(.dina(n4578), .dinb(n1228), .dout(n4579));
  jand g04516(.dina(n4579), .dinb(n4577), .dout(n4580));
  jand g04517(.dina(n4580), .dinb(n3876), .dout(n4581));
  jand g04518(.dina(n4581), .dinb(n4573), .dout(n4582));
  jand g04519(.dina(n3153), .dinb(n1212), .dout(n4583));
  jand g04520(.dina(n4583), .dinb(n1506), .dout(n4584));
  jand g04521(.dina(n678), .dinb(n1270), .dout(n4585));
  jand g04522(.dina(n4585), .dinb(n2521), .dout(n4586));
  jand g04523(.dina(n4586), .dinb(n4584), .dout(n4587));
  jand g04524(.dina(n1325), .dinb(n920), .dout(n4588));
  jand g04525(.dina(n4588), .dinb(n130), .dout(n4589));
  jand g04526(.dina(n586), .dinb(n1349), .dout(n4590));
  jand g04527(.dina(n4590), .dinb(n1310), .dout(n4591));
  jand g04528(.dina(n4591), .dinb(n4589), .dout(n4592));
  jand g04529(.dina(n4592), .dinb(n4587), .dout(n4593));
  jand g04530(.dina(n4593), .dinb(n4582), .dout(n4594));
  jand g04531(.dina(n4594), .dinb(n4571), .dout(n4595));
  jand g04532(.dina(n4595), .dinb(n4553), .dout(n4596));
  jnot g04533(.din(n4596), .dout(n4597));
  jand g04534(.dina(n4597), .dinb(n4527), .dout(n4598));
  jnot g04535(.din(n4598), .dout(n4599));
  jnot g04536(.din(n4471), .dout(n4600));
  jand g04537(.dina(n4597), .dinb(n4600), .dout(n4601));
  jnot g04538(.din(n4601), .dout(n4602));
  jand g04539(.dina(n4600), .dinb(n4406), .dout(n4603));
  jnot g04540(.din(n4603), .dout(n4604));
  jnot g04541(.din(n4472), .dout(n4605));
  jor  g04542(.dina(n4605), .dinb(n4411), .dout(n4606));
  jand g04543(.dina(n4606), .dinb(n4604), .dout(n4607));
  jxor g04544(.dina(n4596), .dinb(n4471), .dout(n4608));
  jnot g04545(.din(n4608), .dout(n4609));
  jor  g04546(.dina(n4609), .dinb(n4607), .dout(n4610));
  jand g04547(.dina(n4610), .dinb(n4602), .dout(n4611));
  jxor g04548(.dina(n4596), .dinb(n4526), .dout(n4612));
  jnot g04549(.din(n4612), .dout(n4613));
  jor  g04550(.dina(n4613), .dinb(n4611), .dout(n4614));
  jand g04551(.dina(n4614), .dinb(n4599), .dout(n4615));
  jand g04552(.dina(n3355), .dinb(n1834), .dout(n4616));
  jand g04553(.dina(n600), .dinb(n1432), .dout(n4617));
  jand g04554(.dina(n3911), .dinb(n1306), .dout(n4618));
  jand g04555(.dina(n4618), .dinb(n3897), .dout(n4619));
  jand g04556(.dina(n4619), .dinb(n4617), .dout(n4620));
  jand g04557(.dina(n4620), .dinb(n931), .dout(n4621));
  jand g04558(.dina(n4621), .dinb(n4616), .dout(n4622));
  jand g04559(.dina(n989), .dinb(n271), .dout(n4623));
  jand g04560(.dina(n1589), .dinb(n1430), .dout(n4624));
  jand g04561(.dina(n4624), .dinb(n1562), .dout(n4625));
  jand g04562(.dina(n4625), .dinb(n1292), .dout(n4626));
  jand g04563(.dina(n4626), .dinb(n4623), .dout(n4627));
  jand g04564(.dina(n4627), .dinb(n4622), .dout(n4628));
  jand g04565(.dina(n833), .dinb(n693), .dout(n4629));
  jand g04566(.dina(n1822), .dinb(n1288), .dout(n4630));
  jand g04567(.dina(n4630), .dinb(n4629), .dout(n4631));
  jand g04568(.dina(n645), .dinb(n481), .dout(n4632));
  jand g04569(.dina(n4632), .dinb(n2538), .dout(n4633));
  jand g04570(.dina(n4633), .dinb(n4631), .dout(n4634));
  jand g04571(.dina(n874), .dinb(n480), .dout(n4635));
  jand g04572(.dina(n4635), .dinb(n557), .dout(n4636));
  jand g04573(.dina(n4636), .dinb(n4634), .dout(n4637));
  jand g04574(.dina(n4637), .dinb(n664), .dout(n4638));
  jand g04575(.dina(n1511), .dinb(n442), .dout(n4639));
  jand g04576(.dina(n4639), .dinb(n1765), .dout(n4640));
  jand g04577(.dina(n2023), .dinb(n470), .dout(n4641));
  jand g04578(.dina(n4641), .dinb(n4640), .dout(n4642));
  jand g04579(.dina(n4642), .dinb(n2164), .dout(n4643));
  jand g04580(.dina(n1846), .dinb(n551), .dout(n4644));
  jand g04581(.dina(n1159), .dinb(n981), .dout(n4645));
  jand g04582(.dina(n4645), .dinb(n4644), .dout(n4646));
  jand g04583(.dina(n4646), .dinb(n3747), .dout(n4647));
  jand g04584(.dina(n4647), .dinb(n4643), .dout(n4648));
  jand g04585(.dina(n4648), .dinb(n4638), .dout(n4649));
  jand g04586(.dina(n583), .dinb(n920), .dout(n4650));
  jand g04587(.dina(n4650), .dinb(n1751), .dout(n4651));
  jand g04588(.dina(n450), .dinb(n1304), .dout(n4652));
  jand g04589(.dina(n4652), .dinb(n1575), .dout(n4653));
  jand g04590(.dina(n4653), .dinb(n4651), .dout(n4654));
  jand g04591(.dina(n461), .dinb(n121), .dout(n4655));
  jand g04592(.dina(n1212), .dinb(n1375), .dout(n4656));
  jand g04593(.dina(n4656), .dinb(n4655), .dout(n4657));
  jand g04594(.dina(n4657), .dinb(n1768), .dout(n4658));
  jand g04595(.dina(n4658), .dinb(n4654), .dout(n4659));
  jand g04596(.dina(n1460), .dinb(n964), .dout(n4660));
  jand g04597(.dina(n4660), .dinb(n1036), .dout(n4661));
  jand g04598(.dina(n4661), .dinb(n1569), .dout(n4662));
  jand g04599(.dina(n4662), .dinb(n1230), .dout(n4663));
  jand g04600(.dina(n4663), .dinb(n4659), .dout(n4664));
  jand g04601(.dina(n1016), .dinb(n454), .dout(n4665));
  jand g04602(.dina(n4665), .dinb(n4664), .dout(n4666));
  jand g04603(.dina(n4666), .dinb(n4649), .dout(n4667));
  jand g04604(.dina(n1522), .dinb(n541), .dout(n4668));
  jand g04605(.dina(n925), .dinb(n619), .dout(n4669));
  jand g04606(.dina(n1453), .dinb(n516), .dout(n4670));
  jand g04607(.dina(n4670), .dinb(n1040), .dout(n4671));
  jand g04608(.dina(n1929), .dinb(n562), .dout(n4672));
  jand g04609(.dina(n4672), .dinb(n4671), .dout(n4673));
  jand g04610(.dina(n4673), .dinb(n4669), .dout(n4674));
  jand g04611(.dina(n1470), .dinb(n826), .dout(n4675));
  jand g04612(.dina(n4675), .dinb(n4674), .dout(n4676));
  jand g04613(.dina(n4676), .dinb(n4668), .dout(n4677));
  jand g04614(.dina(n703), .dinb(n1534), .dout(n4678));
  jand g04615(.dina(n4678), .dinb(n1527), .dout(n4679));
  jand g04616(.dina(n3150), .dinb(n326), .dout(n4680));
  jand g04617(.dina(n4680), .dinb(n3198), .dout(n4681));
  jand g04618(.dina(n4681), .dinb(n4679), .dout(n4682));
  jand g04619(.dina(n4682), .dinb(n1686), .dout(n4683));
  jand g04620(.dina(n4683), .dinb(n4677), .dout(n4684));
  jand g04621(.dina(n4684), .dinb(n4667), .dout(n4685));
  jand g04622(.dina(n4685), .dinb(n4628), .dout(n4686));
  jxor g04623(.dina(n4686), .dinb(n4526), .dout(n4687));
  jxor g04624(.dina(n4687), .dinb(n4615), .dout(n4688));
  jxor g04625(.dina(\a[6] ), .dinb(\a[5] ), .dout(n4689));
  jxor g04626(.dina(\a[8] ), .dinb(\a[7] ), .dout(n4690));
  jand g04627(.dina(n4690), .dinb(n4689), .dout(n4691));
  jnot g04628(.din(n4691), .dout(n4692));
  jor  g04629(.dina(n4692), .dinb(n4688), .dout(n4693));
  jnot g04630(.din(n4689), .dout(n4694));
  jxor g04631(.dina(\a[7] ), .dinb(\a[6] ), .dout(n4695));
  jand g04632(.dina(n4695), .dinb(n4694), .dout(n4696));
  jnot g04633(.din(n4696), .dout(n4697));
  jor  g04634(.dina(n4697), .dinb(n4526), .dout(n4698));
  jor  g04635(.dina(n4695), .dinb(n4689), .dout(n4699));
  jnot g04636(.din(n4699), .dout(n4700));
  jand g04637(.dina(n4700), .dinb(n4690), .dout(n4701));
  jnot g04638(.din(n4701), .dout(n4702));
  jor  g04639(.dina(n4702), .dinb(n4596), .dout(n4703));
  jand g04640(.dina(n4703), .dinb(n4698), .dout(n4704));
  jor  g04641(.dina(n4690), .dinb(n4694), .dout(n4705));
  jor  g04642(.dina(n4705), .dinb(n4686), .dout(n4706));
  jand g04643(.dina(n4706), .dinb(n4704), .dout(n4707));
  jand g04644(.dina(n4707), .dinb(n4693), .dout(n4708));
  jxor g04645(.dina(n4708), .dinb(\a[8] ), .dout(n4709));
  jor  g04646(.dina(n4709), .dinb(n4484), .dout(n4710));
  jnot g04647(.din(n4710), .dout(n4711));
  jxor g04648(.dina(n4314), .dinb(n4312), .dout(n4712));
  jnot g04649(.din(\a[8] ), .dout(n4713));
  jxor g04650(.dina(n4612), .dinb(n4611), .dout(n4714));
  jor  g04651(.dina(n4714), .dinb(n4692), .dout(n4715));
  jor  g04652(.dina(n4697), .dinb(n4596), .dout(n4716));
  jor  g04653(.dina(n4702), .dinb(n4471), .dout(n4717));
  jor  g04654(.dina(n4705), .dinb(n4526), .dout(n4718));
  jand g04655(.dina(n4718), .dinb(n4717), .dout(n4719));
  jand g04656(.dina(n4719), .dinb(n4716), .dout(n4720));
  jand g04657(.dina(n4720), .dinb(n4715), .dout(n4721));
  jxor g04658(.dina(n4721), .dinb(n4713), .dout(n4722));
  jand g04659(.dina(n4722), .dinb(n4712), .dout(n4723));
  jxor g04660(.dina(n4309), .dinb(n4308), .dout(n4724));
  jnot g04661(.din(n4724), .dout(n4725));
  jxor g04662(.dina(n4608), .dinb(n4607), .dout(n4726));
  jor  g04663(.dina(n4726), .dinb(n4692), .dout(n4727));
  jor  g04664(.dina(n4697), .dinb(n4471), .dout(n4728));
  jor  g04665(.dina(n4702), .dinb(n4019), .dout(n4729));
  jor  g04666(.dina(n4705), .dinb(n4596), .dout(n4730));
  jand g04667(.dina(n4730), .dinb(n4729), .dout(n4731));
  jand g04668(.dina(n4731), .dinb(n4728), .dout(n4732));
  jand g04669(.dina(n4732), .dinb(n4727), .dout(n4733));
  jxor g04670(.dina(n4733), .dinb(n4713), .dout(n4734));
  jand g04671(.dina(n4734), .dinb(n4725), .dout(n4735));
  jxor g04672(.dina(n4306), .dinb(n4305), .dout(n4736));
  jnot g04673(.din(n4736), .dout(n4737));
  jor  g04674(.dina(n4692), .dinb(n4473), .dout(n4738));
  jor  g04675(.dina(n4697), .dinb(n4019), .dout(n4739));
  jor  g04676(.dina(n4702), .dinb(n3929), .dout(n4740));
  jand g04677(.dina(n4740), .dinb(n4739), .dout(n4741));
  jor  g04678(.dina(n4705), .dinb(n4471), .dout(n4742));
  jand g04679(.dina(n4742), .dinb(n4741), .dout(n4743));
  jand g04680(.dina(n4743), .dinb(n4738), .dout(n4744));
  jxor g04681(.dina(n4744), .dinb(\a[8] ), .dout(n4745));
  jor  g04682(.dina(n4745), .dinb(n4737), .dout(n4746));
  jnot g04683(.din(n4746), .dout(n4747));
  jxor g04684(.dina(n4303), .dinb(n4302), .dout(n4748));
  jor  g04685(.dina(n4692), .dinb(n4021), .dout(n4749));
  jor  g04686(.dina(n4697), .dinb(n3929), .dout(n4750));
  jor  g04687(.dina(n4705), .dinb(n4019), .dout(n4751));
  jor  g04688(.dina(n4702), .dinb(n3863), .dout(n4752));
  jand g04689(.dina(n4752), .dinb(n4751), .dout(n4753));
  jand g04690(.dina(n4753), .dinb(n4750), .dout(n4754));
  jand g04691(.dina(n4754), .dinb(n4749), .dout(n4755));
  jxor g04692(.dina(n4755), .dinb(n4713), .dout(n4756));
  jand g04693(.dina(n4756), .dinb(n4748), .dout(n4757));
  jxor g04694(.dina(n4300), .dinb(n4299), .dout(n4758));
  jnot g04695(.din(n4758), .dout(n4759));
  jor  g04696(.dina(n4692), .dinb(n4038), .dout(n4760));
  jor  g04697(.dina(n4697), .dinb(n3863), .dout(n4761));
  jor  g04698(.dina(n4705), .dinb(n3929), .dout(n4762));
  jand g04699(.dina(n4762), .dinb(n4761), .dout(n4763));
  jor  g04700(.dina(n4702), .dinb(n3787), .dout(n4764));
  jand g04701(.dina(n4764), .dinb(n4763), .dout(n4765));
  jand g04702(.dina(n4765), .dinb(n4760), .dout(n4766));
  jxor g04703(.dina(n4766), .dinb(\a[8] ), .dout(n4767));
  jor  g04704(.dina(n4767), .dinb(n4759), .dout(n4768));
  jnot g04705(.din(n4768), .dout(n4769));
  jxor g04706(.dina(n4297), .dinb(n4296), .dout(n4770));
  jor  g04707(.dina(n4692), .dinb(n4051), .dout(n4771));
  jor  g04708(.dina(n4697), .dinb(n3787), .dout(n4772));
  jor  g04709(.dina(n4705), .dinb(n3863), .dout(n4773));
  jor  g04710(.dina(n4702), .dinb(n3420), .dout(n4774));
  jand g04711(.dina(n4774), .dinb(n4773), .dout(n4775));
  jand g04712(.dina(n4775), .dinb(n4772), .dout(n4776));
  jand g04713(.dina(n4776), .dinb(n4771), .dout(n4777));
  jxor g04714(.dina(n4777), .dinb(n4713), .dout(n4778));
  jand g04715(.dina(n4778), .dinb(n4770), .dout(n4779));
  jxor g04716(.dina(n4294), .dinb(n4292), .dout(n4780));
  jor  g04717(.dina(n4692), .dinb(n3789), .dout(n4781));
  jor  g04718(.dina(n4697), .dinb(n3420), .dout(n4782));
  jor  g04719(.dina(n4702), .dinb(n3286), .dout(n4783));
  jand g04720(.dina(n4783), .dinb(n4782), .dout(n4784));
  jor  g04721(.dina(n4705), .dinb(n3787), .dout(n4785));
  jand g04722(.dina(n4785), .dinb(n4784), .dout(n4786));
  jand g04723(.dina(n4786), .dinb(n4781), .dout(n4787));
  jxor g04724(.dina(n4787), .dinb(\a[8] ), .dout(n4788));
  jor  g04725(.dina(n4788), .dinb(n4780), .dout(n4789));
  jnot g04726(.din(n4789), .dout(n4790));
  jxor g04727(.dina(n4290), .dinb(n4288), .dout(n4791));
  jnot g04728(.din(n4791), .dout(n4792));
  jor  g04729(.dina(n4702), .dinb(n3203), .dout(n4793));
  jor  g04730(.dina(n4692), .dinb(n3422), .dout(n4794));
  jor  g04731(.dina(n4705), .dinb(n3420), .dout(n4795));
  jor  g04732(.dina(n4697), .dinb(n3286), .dout(n4796));
  jand g04733(.dina(n4796), .dinb(n4795), .dout(n4797));
  jand g04734(.dina(n4797), .dinb(n4794), .dout(n4798));
  jand g04735(.dina(n4798), .dinb(n4793), .dout(n4799));
  jxor g04736(.dina(n4799), .dinb(\a[8] ), .dout(n4800));
  jor  g04737(.dina(n4800), .dinb(n4792), .dout(n4801));
  jnot g04738(.din(n4801), .dout(n4802));
  jxor g04739(.dina(n4286), .dinb(n4284), .dout(n4803));
  jnot g04740(.din(n4803), .dout(n4804));
  jor  g04741(.dina(n4692), .dinb(n3440), .dout(n4805));
  jor  g04742(.dina(n4697), .dinb(n3203), .dout(n4806));
  jor  g04743(.dina(n4705), .dinb(n3286), .dout(n4807));
  jand g04744(.dina(n4807), .dinb(n4806), .dout(n4808));
  jor  g04745(.dina(n4702), .dinb(n3072), .dout(n4809));
  jand g04746(.dina(n4809), .dinb(n4808), .dout(n4810));
  jand g04747(.dina(n4810), .dinb(n4805), .dout(n4811));
  jxor g04748(.dina(n4811), .dinb(\a[8] ), .dout(n4812));
  jor  g04749(.dina(n4812), .dinb(n4804), .dout(n4813));
  jnot g04750(.din(n4813), .dout(n4814));
  jxor g04751(.dina(n4282), .dinb(n4280), .dout(n4815));
  jnot g04752(.din(n4815), .dout(n4816));
  jor  g04753(.dina(n4692), .dinb(n3451), .dout(n4817));
  jor  g04754(.dina(n4697), .dinb(n3072), .dout(n4818));
  jor  g04755(.dina(n4705), .dinb(n3203), .dout(n4819));
  jand g04756(.dina(n4819), .dinb(n4818), .dout(n4820));
  jor  g04757(.dina(n4702), .dinb(n2738), .dout(n4821));
  jand g04758(.dina(n4821), .dinb(n4820), .dout(n4822));
  jand g04759(.dina(n4822), .dinb(n4817), .dout(n4823));
  jxor g04760(.dina(n4823), .dinb(\a[8] ), .dout(n4824));
  jor  g04761(.dina(n4824), .dinb(n4816), .dout(n4825));
  jnot g04762(.din(n4825), .dout(n4826));
  jxor g04763(.dina(n4278), .dinb(n4276), .dout(n4827));
  jnot g04764(.din(n4827), .dout(n4828));
  jor  g04765(.dina(n4692), .dinb(n3081), .dout(n4829));
  jor  g04766(.dina(n4702), .dinb(n2553), .dout(n4830));
  jor  g04767(.dina(n4697), .dinb(n2738), .dout(n4831));
  jand g04768(.dina(n4831), .dinb(n4830), .dout(n4832));
  jor  g04769(.dina(n4705), .dinb(n3072), .dout(n4833));
  jand g04770(.dina(n4833), .dinb(n4832), .dout(n4834));
  jand g04771(.dina(n4834), .dinb(n4829), .dout(n4835));
  jxor g04772(.dina(n4835), .dinb(\a[8] ), .dout(n4836));
  jor  g04773(.dina(n4836), .dinb(n4828), .dout(n4837));
  jnot g04774(.din(n4837), .dout(n4838));
  jxor g04775(.dina(n4274), .dinb(n4272), .dout(n4839));
  jor  g04776(.dina(n4692), .dinb(n2740), .dout(n4840));
  jor  g04777(.dina(n4697), .dinb(n2553), .dout(n4841));
  jor  g04778(.dina(n4702), .dinb(n2629), .dout(n4842));
  jor  g04779(.dina(n4705), .dinb(n2738), .dout(n4843));
  jand g04780(.dina(n4843), .dinb(n4842), .dout(n4844));
  jand g04781(.dina(n4844), .dinb(n4841), .dout(n4845));
  jand g04782(.dina(n4845), .dinb(n4840), .dout(n4846));
  jxor g04783(.dina(n4846), .dinb(n4713), .dout(n4847));
  jand g04784(.dina(n4847), .dinb(n4839), .dout(n4848));
  jxor g04785(.dina(n4269), .dinb(n4268), .dout(n4849));
  jor  g04786(.dina(n4692), .dinb(n2768), .dout(n4850));
  jor  g04787(.dina(n4705), .dinb(n2553), .dout(n4851));
  jor  g04788(.dina(n4702), .dinb(n2428), .dout(n4852));
  jor  g04789(.dina(n4697), .dinb(n2629), .dout(n4853));
  jand g04790(.dina(n4853), .dinb(n4852), .dout(n4854));
  jand g04791(.dina(n4854), .dinb(n4851), .dout(n4855));
  jand g04792(.dina(n4855), .dinb(n4850), .dout(n4856));
  jxor g04793(.dina(n4856), .dinb(n4713), .dout(n4857));
  jand g04794(.dina(n4857), .dinb(n4849), .dout(n4858));
  jnot g04795(.din(n4858), .dout(n4859));
  jxor g04796(.dina(n4264), .dinb(n4263), .dout(n4860));
  jnot g04797(.din(n4860), .dout(n4861));
  jor  g04798(.dina(n4692), .dinb(n2779), .dout(n4862));
  jor  g04799(.dina(n4697), .dinb(n2428), .dout(n4863));
  jor  g04800(.dina(n4705), .dinb(n2629), .dout(n4864));
  jand g04801(.dina(n4864), .dinb(n4863), .dout(n4865));
  jor  g04802(.dina(n4702), .dinb(n2174), .dout(n4866));
  jand g04803(.dina(n4866), .dinb(n4865), .dout(n4867));
  jand g04804(.dina(n4867), .dinb(n4862), .dout(n4868));
  jxor g04805(.dina(n4868), .dinb(\a[8] ), .dout(n4869));
  jor  g04806(.dina(n4869), .dinb(n4861), .dout(n4870));
  jxor g04807(.dina(n4261), .dinb(n4260), .dout(n4871));
  jor  g04808(.dina(n4692), .dinb(n2430), .dout(n4872));
  jor  g04809(.dina(n4697), .dinb(n2174), .dout(n4873));
  jor  g04810(.dina(n4705), .dinb(n2428), .dout(n4874));
  jor  g04811(.dina(n4702), .dinb(n1954), .dout(n4875));
  jand g04812(.dina(n4875), .dinb(n4874), .dout(n4876));
  jand g04813(.dina(n4876), .dinb(n4873), .dout(n4877));
  jand g04814(.dina(n4877), .dinb(n4872), .dout(n4878));
  jxor g04815(.dina(n4878), .dinb(n4713), .dout(n4879));
  jand g04816(.dina(n4879), .dinb(n4871), .dout(n4880));
  jnot g04817(.din(n4880), .dout(n4881));
  jxor g04818(.dina(n4258), .dinb(n4257), .dout(n4882));
  jor  g04819(.dina(n4692), .dinb(n2176), .dout(n4883));
  jor  g04820(.dina(n4705), .dinb(n2174), .dout(n4884));
  jor  g04821(.dina(n4702), .dinb(n2057), .dout(n4885));
  jor  g04822(.dina(n4697), .dinb(n1954), .dout(n4886));
  jand g04823(.dina(n4886), .dinb(n4885), .dout(n4887));
  jand g04824(.dina(n4887), .dinb(n4884), .dout(n4888));
  jand g04825(.dina(n4888), .dinb(n4883), .dout(n4889));
  jxor g04826(.dina(n4889), .dinb(n4713), .dout(n4890));
  jand g04827(.dina(n4890), .dinb(n4882), .dout(n4891));
  jnot g04828(.din(n4891), .dout(n4892));
  jxor g04829(.dina(n4253), .dinb(n4252), .dout(n4893));
  jnot g04830(.din(n4893), .dout(n4894));
  jor  g04831(.dina(n4702), .dinb(n1790), .dout(n4895));
  jor  g04832(.dina(n4692), .dinb(n2197), .dout(n4896));
  jor  g04833(.dina(n4705), .dinb(n1954), .dout(n4897));
  jor  g04834(.dina(n4697), .dinb(n2057), .dout(n4898));
  jand g04835(.dina(n4898), .dinb(n4897), .dout(n4899));
  jand g04836(.dina(n4899), .dinb(n4896), .dout(n4900));
  jand g04837(.dina(n4900), .dinb(n4895), .dout(n4901));
  jxor g04838(.dina(n4901), .dinb(\a[8] ), .dout(n4902));
  jor  g04839(.dina(n4902), .dinb(n4894), .dout(n4903));
  jxor g04840(.dina(n4249), .dinb(n4241), .dout(n4904));
  jor  g04841(.dina(n4692), .dinb(n2208), .dout(n4905));
  jor  g04842(.dina(n4697), .dinb(n1790), .dout(n4906));
  jor  g04843(.dina(n4702), .dinb(n1606), .dout(n4907));
  jor  g04844(.dina(n4705), .dinb(n2057), .dout(n4908));
  jand g04845(.dina(n4908), .dinb(n4907), .dout(n4909));
  jand g04846(.dina(n4909), .dinb(n4906), .dout(n4910));
  jand g04847(.dina(n4910), .dinb(n4905), .dout(n4911));
  jxor g04848(.dina(n4911), .dinb(n4713), .dout(n4912));
  jand g04849(.dina(n4912), .dinb(n4904), .dout(n4913));
  jnot g04850(.din(n4913), .dout(n4914));
  jor  g04851(.dina(n4705), .dinb(n1790), .dout(n4915));
  jor  g04852(.dina(n4692), .dinb(n1792), .dout(n4916));
  jor  g04853(.dina(n4702), .dinb(n1448), .dout(n4917));
  jor  g04854(.dina(n4697), .dinb(n1606), .dout(n4918));
  jand g04855(.dina(n4918), .dinb(n4917), .dout(n4919));
  jand g04856(.dina(n4919), .dinb(n4916), .dout(n4920));
  jand g04857(.dina(n4920), .dinb(n4915), .dout(n4921));
  jxor g04858(.dina(n4921), .dinb(\a[8] ), .dout(n4922));
  jnot g04859(.din(n4922), .dout(n4923));
  jor  g04860(.dina(n4228), .dinb(n4050), .dout(n4924));
  jxor g04861(.dina(n4924), .dinb(n4236), .dout(n4925));
  jand g04862(.dina(n4925), .dinb(n4923), .dout(n4926));
  jnot g04863(.din(n4926), .dout(n4927));
  jand g04864(.dina(n4225), .dinb(\a[11] ), .dout(n4928));
  jxor g04865(.dina(n4928), .dinb(n4223), .dout(n4929));
  jnot g04866(.din(n4929), .dout(n4930));
  jor  g04867(.dina(n4692), .dinb(n1608), .dout(n4931));
  jor  g04868(.dina(n4697), .dinb(n1448), .dout(n4932));
  jor  g04869(.dina(n4702), .dinb(n1255), .dout(n4933));
  jand g04870(.dina(n4933), .dinb(n4932), .dout(n4934));
  jor  g04871(.dina(n4705), .dinb(n1606), .dout(n4935));
  jand g04872(.dina(n4935), .dinb(n4934), .dout(n4936));
  jand g04873(.dina(n4936), .dinb(n4931), .dout(n4937));
  jxor g04874(.dina(n4937), .dinb(\a[8] ), .dout(n4938));
  jor  g04875(.dina(n4938), .dinb(n4930), .dout(n4939));
  jand g04876(.dina(n4691), .dinb(n728), .dout(n4940));
  jnot g04877(.din(n4705), .dout(n4941));
  jand g04878(.dina(n4941), .dinb(n795), .dout(n4942));
  jand g04879(.dina(n4696), .dinb(n438), .dout(n4943));
  jor  g04880(.dina(n4943), .dinb(n4942), .dout(n4944));
  jor  g04881(.dina(n4944), .dinb(n4940), .dout(n4945));
  jnot g04882(.din(n4945), .dout(n4946));
  jand g04883(.dina(n4689), .dinb(n438), .dout(n4947));
  jnot g04884(.din(n4947), .dout(n4948));
  jand g04885(.dina(n4948), .dinb(\a[8] ), .dout(n4949));
  jand g04886(.dina(n4949), .dinb(n4946), .dout(n4950));
  jand g04887(.dina(n4691), .dinb(n1639), .dout(n4951));
  jand g04888(.dina(n4696), .dinb(n795), .dout(n4952));
  jand g04889(.dina(n4941), .dinb(n1175), .dout(n4953));
  jor  g04890(.dina(n4953), .dinb(n4952), .dout(n4954));
  jand g04891(.dina(n4701), .dinb(n438), .dout(n4955));
  jor  g04892(.dina(n4955), .dinb(n4954), .dout(n4956));
  jor  g04893(.dina(n4956), .dinb(n4951), .dout(n4957));
  jnot g04894(.din(n4957), .dout(n4958));
  jand g04895(.dina(n4958), .dinb(n4950), .dout(n4959));
  jand g04896(.dina(n4959), .dinb(n4225), .dout(n4960));
  jnot g04897(.din(n4960), .dout(n4961));
  jxor g04898(.dina(n4959), .dinb(n4225), .dout(n4962));
  jnot g04899(.din(n4962), .dout(n4963));
  jor  g04900(.dina(n4692), .dinb(n1656), .dout(n4964));
  jor  g04901(.dina(n4702), .dinb(n726), .dout(n4965));
  jor  g04902(.dina(n4697), .dinb(n1255), .dout(n4966));
  jand g04903(.dina(n4966), .dinb(n4965), .dout(n4967));
  jor  g04904(.dina(n4705), .dinb(n1448), .dout(n4968));
  jand g04905(.dina(n4968), .dinb(n4967), .dout(n4969));
  jand g04906(.dina(n4969), .dinb(n4964), .dout(n4970));
  jxor g04907(.dina(n4970), .dinb(\a[8] ), .dout(n4971));
  jor  g04908(.dina(n4971), .dinb(n4963), .dout(n4972));
  jand g04909(.dina(n4972), .dinb(n4961), .dout(n4973));
  jnot g04910(.din(n4973), .dout(n4974));
  jxor g04911(.dina(n4938), .dinb(n4930), .dout(n4975));
  jand g04912(.dina(n4975), .dinb(n4974), .dout(n4976));
  jnot g04913(.din(n4976), .dout(n4977));
  jand g04914(.dina(n4977), .dinb(n4939), .dout(n4978));
  jxor g04915(.dina(n4925), .dinb(n4923), .dout(n4979));
  jnot g04916(.din(n4979), .dout(n4980));
  jor  g04917(.dina(n4980), .dinb(n4978), .dout(n4981));
  jand g04918(.dina(n4981), .dinb(n4927), .dout(n4982));
  jxor g04919(.dina(n4912), .dinb(n4904), .dout(n4983));
  jnot g04920(.din(n4983), .dout(n4984));
  jor  g04921(.dina(n4984), .dinb(n4982), .dout(n4985));
  jand g04922(.dina(n4985), .dinb(n4914), .dout(n4986));
  jxor g04923(.dina(n4902), .dinb(n4894), .dout(n4987));
  jnot g04924(.din(n4987), .dout(n4988));
  jor  g04925(.dina(n4988), .dinb(n4986), .dout(n4989));
  jand g04926(.dina(n4989), .dinb(n4903), .dout(n4990));
  jxor g04927(.dina(n4890), .dinb(n4882), .dout(n4991));
  jnot g04928(.din(n4991), .dout(n4992));
  jor  g04929(.dina(n4992), .dinb(n4990), .dout(n4993));
  jand g04930(.dina(n4993), .dinb(n4892), .dout(n4994));
  jxor g04931(.dina(n4879), .dinb(n4871), .dout(n4995));
  jnot g04932(.din(n4995), .dout(n4996));
  jor  g04933(.dina(n4996), .dinb(n4994), .dout(n4997));
  jand g04934(.dina(n4997), .dinb(n4881), .dout(n4998));
  jxor g04935(.dina(n4869), .dinb(n4861), .dout(n4999));
  jnot g04936(.din(n4999), .dout(n5000));
  jor  g04937(.dina(n5000), .dinb(n4998), .dout(n5001));
  jand g04938(.dina(n5001), .dinb(n4870), .dout(n5002));
  jxor g04939(.dina(n4857), .dinb(n4849), .dout(n5003));
  jnot g04940(.din(n5003), .dout(n5004));
  jor  g04941(.dina(n5004), .dinb(n5002), .dout(n5005));
  jand g04942(.dina(n5005), .dinb(n4859), .dout(n5006));
  jnot g04943(.din(n5006), .dout(n5007));
  jxor g04944(.dina(n4847), .dinb(n4839), .dout(n5008));
  jand g04945(.dina(n5008), .dinb(n5007), .dout(n5009));
  jor  g04946(.dina(n5009), .dinb(n4848), .dout(n5010));
  jxor g04947(.dina(n4836), .dinb(n4827), .dout(n5011));
  jnot g04948(.din(n5011), .dout(n5012));
  jand g04949(.dina(n5012), .dinb(n5010), .dout(n5013));
  jor  g04950(.dina(n5013), .dinb(n4838), .dout(n5014));
  jxor g04951(.dina(n4824), .dinb(n4815), .dout(n5015));
  jnot g04952(.din(n5015), .dout(n5016));
  jand g04953(.dina(n5016), .dinb(n5014), .dout(n5017));
  jor  g04954(.dina(n5017), .dinb(n4826), .dout(n5018));
  jxor g04955(.dina(n4812), .dinb(n4803), .dout(n5019));
  jnot g04956(.din(n5019), .dout(n5020));
  jand g04957(.dina(n5020), .dinb(n5018), .dout(n5021));
  jor  g04958(.dina(n5021), .dinb(n4814), .dout(n5022));
  jxor g04959(.dina(n4800), .dinb(n4792), .dout(n5023));
  jand g04960(.dina(n5023), .dinb(n5022), .dout(n5024));
  jor  g04961(.dina(n5024), .dinb(n4802), .dout(n5025));
  jxor g04962(.dina(n4788), .dinb(n4780), .dout(n5026));
  jand g04963(.dina(n5026), .dinb(n5025), .dout(n5027));
  jor  g04964(.dina(n5027), .dinb(n4790), .dout(n5028));
  jxor g04965(.dina(n4778), .dinb(n4770), .dout(n5029));
  jand g04966(.dina(n5029), .dinb(n5028), .dout(n5030));
  jor  g04967(.dina(n5030), .dinb(n4779), .dout(n5031));
  jxor g04968(.dina(n4767), .dinb(n4758), .dout(n5032));
  jnot g04969(.din(n5032), .dout(n5033));
  jand g04970(.dina(n5033), .dinb(n5031), .dout(n5034));
  jor  g04971(.dina(n5034), .dinb(n4769), .dout(n5035));
  jxor g04972(.dina(n4756), .dinb(n4748), .dout(n5036));
  jand g04973(.dina(n5036), .dinb(n5035), .dout(n5037));
  jor  g04974(.dina(n5037), .dinb(n4757), .dout(n5038));
  jxor g04975(.dina(n4745), .dinb(n4736), .dout(n5039));
  jnot g04976(.din(n5039), .dout(n5040));
  jand g04977(.dina(n5040), .dinb(n5038), .dout(n5041));
  jor  g04978(.dina(n5041), .dinb(n4747), .dout(n5042));
  jxor g04979(.dina(n4734), .dinb(n4724), .dout(n5043));
  jnot g04980(.din(n5043), .dout(n5044));
  jand g04981(.dina(n5044), .dinb(n5042), .dout(n5045));
  jor  g04982(.dina(n5045), .dinb(n4735), .dout(n5046));
  jxor g04983(.dina(n4722), .dinb(n4712), .dout(n5047));
  jand g04984(.dina(n5047), .dinb(n5046), .dout(n5048));
  jor  g04985(.dina(n5048), .dinb(n4723), .dout(n5049));
  jxor g04986(.dina(n4709), .dinb(n4484), .dout(n5050));
  jand g04987(.dina(n5050), .dinb(n5049), .dout(n5051));
  jor  g04988(.dina(n5051), .dinb(n4711), .dout(n5052));
  jand g04989(.dina(n4481), .dinb(n4405), .dout(n5053));
  jand g04990(.dina(n4482), .dinb(n4316), .dout(n5054));
  jor  g04991(.dina(n5054), .dinb(n5053), .dout(n5055));
  jand g04992(.dina(n4403), .dinb(n4395), .dout(n5056));
  jand g04993(.dina(n4404), .dinb(n4320), .dout(n5057));
  jor  g04994(.dina(n5057), .dinb(n5056), .dout(n5058));
  jor  g04995(.dina(n4393), .dinb(n4385), .dout(n5059));
  jand g04996(.dina(n4394), .dinb(n4325), .dout(n5060));
  jnot g04997(.din(n5060), .dout(n5061));
  jand g04998(.dina(n5061), .dinb(n5059), .dout(n5062));
  jnot g04999(.din(n5062), .dout(n5063));
  jand g05000(.dina(n4382), .dinb(n4374), .dout(n5064));
  jand g05001(.dina(n4383), .dinb(n4328), .dout(n5065));
  jor  g05002(.dina(n5065), .dinb(n5064), .dout(n5066));
  jand g05003(.dina(n4372), .dinb(n4364), .dout(n5067));
  jand g05004(.dina(n4373), .dinb(n4333), .dout(n5068));
  jor  g05005(.dina(n5068), .dinb(n5067), .dout(n5069));
  jand g05006(.dina(n4362), .dinb(n4354), .dout(n5070));
  jand g05007(.dina(n4363), .dinb(n4336), .dout(n5071));
  jor  g05008(.dina(n5071), .dinb(n5070), .dout(n5072));
  jand g05009(.dina(n4341), .dinb(n4339), .dout(n5073));
  jand g05010(.dina(n4353), .dinb(n4342), .dout(n5074));
  jor  g05011(.dina(n5074), .dinb(n5073), .dout(n5075));
  jand g05012(.dina(n4338), .dinb(\a[31] ), .dout(n5076));
  jand g05013(.dina(n5076), .dinb(n728), .dout(n5077));
  jnot g05014(.din(\a[31] ), .dout(n5078));
  jand g05015(.dina(n264), .dinb(n5078), .dout(n5079));
  jand g05016(.dina(n106), .dinb(\a[31] ), .dout(n5080));
  jor  g05017(.dina(n5080), .dinb(n5079), .dout(n5081));
  jnot g05018(.din(n5081), .dout(n5082));
  jand g05019(.dina(n5082), .dinb(n438), .dout(n5083));
  jand g05020(.dina(n4338), .dinb(n5078), .dout(n5084));
  jand g05021(.dina(n5084), .dinb(n795), .dout(n5085));
  jor  g05022(.dina(n5085), .dinb(n5083), .dout(n5086));
  jor  g05023(.dina(n5086), .dinb(n5077), .dout(n5087));
  jnot g05024(.din(n5087), .dout(n5088));
  jor  g05025(.dina(n4343), .dinb(n1608), .dout(n5089));
  jor  g05026(.dina(n4346), .dinb(n1448), .dout(n5090));
  jor  g05027(.dina(n3683), .dinb(n1255), .dout(n5091));
  jand g05028(.dina(n5091), .dinb(n5090), .dout(n5092));
  jor  g05029(.dina(n4348), .dinb(n1606), .dout(n5093));
  jand g05030(.dina(n5093), .dinb(n5092), .dout(n5094));
  jand g05031(.dina(n5094), .dinb(n5089), .dout(n5095));
  jxor g05032(.dina(n5095), .dinb(\a[29] ), .dout(n5096));
  jxor g05033(.dina(n5096), .dinb(n5088), .dout(n5097));
  jxor g05034(.dina(n5097), .dinb(n5075), .dout(n5098));
  jnot g05035(.din(n5098), .dout(n5099));
  jor  g05036(.dina(n1805), .dinb(n1790), .dout(n5100));
  jor  g05037(.dina(n2197), .dinb(n2303), .dout(n5101));
  jor  g05038(.dina(n1954), .dinb(n2309), .dout(n5102));
  jor  g05039(.dina(n2057), .dinb(n2306), .dout(n5103));
  jand g05040(.dina(n5103), .dinb(n5102), .dout(n5104));
  jand g05041(.dina(n5104), .dinb(n5101), .dout(n5105));
  jand g05042(.dina(n5105), .dinb(n5100), .dout(n5106));
  jxor g05043(.dina(n5106), .dinb(\a[26] ), .dout(n5107));
  jxor g05044(.dina(n5107), .dinb(n5099), .dout(n5108));
  jxor g05045(.dina(n5108), .dinb(n5072), .dout(n5109));
  jnot g05046(.din(n5109), .dout(n5110));
  jor  g05047(.dina(n2779), .dinb(n807), .dout(n5111));
  jor  g05048(.dina(n2428), .dinb(n1613), .dout(n5112));
  jor  g05049(.dina(n2629), .dinb(n1621), .dout(n5113));
  jand g05050(.dina(n5113), .dinb(n5112), .dout(n5114));
  jor  g05051(.dina(n2174), .dinb(n1617), .dout(n5115));
  jand g05052(.dina(n5115), .dinb(n5114), .dout(n5116));
  jand g05053(.dina(n5116), .dinb(n5111), .dout(n5117));
  jxor g05054(.dina(n5117), .dinb(\a[23] ), .dout(n5118));
  jxor g05055(.dina(n5118), .dinb(n5110), .dout(n5119));
  jxor g05056(.dina(n5119), .dinb(n5069), .dout(n5120));
  jor  g05057(.dina(n3081), .dinb(n1820), .dout(n5121));
  jor  g05058(.dina(n2553), .dinb(n2186), .dout(n5122));
  jor  g05059(.dina(n2738), .dinb(n2181), .dout(n5123));
  jor  g05060(.dina(n3072), .dinb(n2189), .dout(n5124));
  jand g05061(.dina(n5124), .dinb(n5123), .dout(n5125));
  jand g05062(.dina(n5125), .dinb(n5122), .dout(n5126));
  jand g05063(.dina(n5126), .dinb(n5121), .dout(n5127));
  jxor g05064(.dina(n5127), .dinb(n2196), .dout(n5128));
  jxor g05065(.dina(n5128), .dinb(n5120), .dout(n5129));
  jxor g05066(.dina(n5129), .dinb(n5066), .dout(n5130));
  jnot g05067(.din(n5130), .dout(n5131));
  jor  g05068(.dina(n3203), .dinb(n2758), .dout(n5132));
  jor  g05069(.dina(n3422), .dinb(n2744), .dout(n5133));
  jor  g05070(.dina(n3420), .dinb(n2753), .dout(n5134));
  jor  g05071(.dina(n3286), .dinb(n2749), .dout(n5135));
  jand g05072(.dina(n5135), .dinb(n5134), .dout(n5136));
  jand g05073(.dina(n5136), .dinb(n5133), .dout(n5137));
  jand g05074(.dina(n5137), .dinb(n5132), .dout(n5138));
  jxor g05075(.dina(n5138), .dinb(\a[17] ), .dout(n5139));
  jxor g05076(.dina(n5139), .dinb(n5131), .dout(n5140));
  jxor g05077(.dina(n5140), .dinb(n5063), .dout(n5141));
  jor  g05078(.dina(n4038), .dinb(n3424), .dout(n5142));
  jor  g05079(.dina(n3863), .dinb(n3429), .dout(n5143));
  jor  g05080(.dina(n3929), .dinb(n3426), .dout(n5144));
  jand g05081(.dina(n5144), .dinb(n5143), .dout(n5145));
  jor  g05082(.dina(n3787), .dinb(n3211), .dout(n5146));
  jand g05083(.dina(n5146), .dinb(n5145), .dout(n5147));
  jand g05084(.dina(n5147), .dinb(n5142), .dout(n5148));
  jxor g05085(.dina(n5148), .dinb(\a[14] ), .dout(n5149));
  jxor g05086(.dina(n5149), .dinb(n5141), .dout(n5150));
  jxor g05087(.dina(n5150), .dinb(n5058), .dout(n5151));
  jor  g05088(.dina(n4726), .dinb(n4023), .dout(n5152));
  jor  g05089(.dina(n4471), .dinb(n4028), .dout(n5153));
  jor  g05090(.dina(n4596), .dinb(n4025), .dout(n5154));
  jor  g05091(.dina(n4019), .dinb(n3871), .dout(n5155));
  jand g05092(.dina(n5155), .dinb(n5154), .dout(n5156));
  jand g05093(.dina(n5156), .dinb(n5153), .dout(n5157));
  jand g05094(.dina(n5157), .dinb(n5152), .dout(n5158));
  jxor g05095(.dina(n5158), .dinb(n4050), .dout(n5159));
  jxor g05096(.dina(n5159), .dinb(n5151), .dout(n5160));
  jnot g05097(.din(n5160), .dout(n5161));
  jxor g05098(.dina(n5161), .dinb(n5055), .dout(n5162));
  jnot g05099(.din(n4686), .dout(n5163));
  jand g05100(.dina(n5163), .dinb(n4527), .dout(n5164));
  jnot g05101(.din(n5164), .dout(n5165));
  jnot g05102(.din(n4687), .dout(n5166));
  jor  g05103(.dina(n5166), .dinb(n4615), .dout(n5167));
  jand g05104(.dina(n5167), .dinb(n5165), .dout(n5168));
  jand g05105(.dina(n4528), .dinb(n1577), .dout(n5169));
  jand g05106(.dina(n5169), .dinb(n514), .dout(n5170));
  jand g05107(.dina(n714), .dinb(n1292), .dout(n5171));
  jand g05108(.dina(n1349), .dinb(n266), .dout(n5172));
  jand g05109(.dina(n5172), .dinb(n5171), .dout(n5173));
  jand g05110(.dina(n5173), .dinb(n1851), .dout(n5174));
  jand g05111(.dina(n1591), .dinb(n1432), .dout(n5175));
  jand g05112(.dina(n5175), .dinb(n1706), .dout(n5176));
  jand g05113(.dina(n5176), .dinb(n5174), .dout(n5177));
  jand g05114(.dina(n5177), .dinb(n5170), .dout(n5178));
  jand g05115(.dina(n172), .dinb(n100), .dout(n5179));
  jand g05116(.dina(n461), .dinb(n1309), .dout(n5180));
  jand g05117(.dina(n5180), .dinb(n2508), .dout(n5181));
  jand g05118(.dina(n5181), .dinb(n5179), .dout(n5182));
  jand g05119(.dina(n1891), .dinb(n1885), .dout(n5183));
  jand g05120(.dina(n5183), .dinb(n5182), .dout(n5184));
  jand g05121(.dina(n5184), .dinb(n5178), .dout(n5185));
  jand g05122(.dina(n351), .dinb(n1324), .dout(n5186));
  jand g05123(.dina(n5186), .dinb(n532), .dout(n5187));
  jand g05124(.dina(n678), .dinb(n1361), .dout(n5188));
  jand g05125(.dina(n5188), .dinb(n1569), .dout(n5189));
  jand g05126(.dina(n5189), .dinb(n136), .dout(n5190));
  jand g05127(.dina(n5190), .dinb(n5187), .dout(n5191));
  jand g05128(.dina(n5191), .dinb(n2154), .dout(n5192));
  jand g05129(.dina(n5192), .dinb(n5185), .dout(n5193));
  jand g05130(.dina(n1042), .dinb(n325), .dout(n5194));
  jand g05131(.dina(n5194), .dinb(n2700), .dout(n5195));
  jand g05132(.dina(n5195), .dinb(n1772), .dout(n5196));
  jand g05133(.dina(n833), .dinb(n1449), .dout(n5197));
  jand g05134(.dina(n818), .dinb(n811), .dout(n5198));
  jand g05135(.dina(n5198), .dinb(n1987), .dout(n5199));
  jand g05136(.dina(n5199), .dinb(n5197), .dout(n5200));
  jand g05137(.dina(n3328), .dinb(n1305), .dout(n5201));
  jand g05138(.dina(n641), .dinb(n1822), .dout(n5202));
  jand g05139(.dina(n5202), .dinb(n5201), .dout(n5203));
  jand g05140(.dina(n5203), .dinb(n5200), .dout(n5204));
  jand g05141(.dina(n5204), .dinb(n5196), .dout(n5205));
  jand g05142(.dina(n1731), .dinb(n645), .dout(n5206));
  jand g05143(.dina(n5206), .dinb(n1476), .dout(n5207));
  jand g05144(.dina(n2100), .dinb(n895), .dout(n5208));
  jand g05145(.dina(n5208), .dinb(n2077), .dout(n5209));
  jand g05146(.dina(n5209), .dinb(n5207), .dout(n5210));
  jand g05147(.dina(n4639), .dinb(n1168), .dout(n5211));
  jand g05148(.dina(n5211), .dinb(n5210), .dout(n5212));
  jand g05149(.dina(n5212), .dinb(n1365), .dout(n5213));
  jand g05150(.dina(n5213), .dinb(n5205), .dout(n5214));
  jand g05151(.dina(n2152), .dinb(n951), .dout(n5215));
  jand g05152(.dina(n2406), .dinb(n1308), .dout(n5216));
  jand g05153(.dina(n5216), .dinb(n5215), .dout(n5217));
  jand g05154(.dina(n1451), .dinb(n1107), .dout(n5218));
  jand g05155(.dina(n981), .dinb(n548), .dout(n5219));
  jand g05156(.dina(n5219), .dinb(n5218), .dout(n5220));
  jand g05157(.dina(n5220), .dinb(n1532), .dout(n5221));
  jand g05158(.dina(n1515), .dinb(n450), .dout(n5222));
  jand g05159(.dina(n5222), .dinb(n3802), .dout(n5223));
  jand g05160(.dina(n639), .dinb(n954), .dout(n5224));
  jand g05161(.dina(n5224), .dinb(n5223), .dout(n5225));
  jand g05162(.dina(n5225), .dinb(n5221), .dout(n5226));
  jand g05163(.dina(n5226), .dinb(n5217), .dout(n5227));
  jand g05164(.dina(n5227), .dinb(n5214), .dout(n5228));
  jand g05165(.dina(n1575), .dinb(n676), .dout(n5229));
  jand g05166(.dina(n5229), .dinb(n516), .dout(n5230));
  jand g05167(.dina(n1524), .dinb(n130), .dout(n5231));
  jand g05168(.dina(n1227), .dinb(n1583), .dout(n5232));
  jand g05169(.dina(n5232), .dinb(n5231), .dout(n5233));
  jand g05170(.dina(n5233), .dinb(n5230), .dout(n5234));
  jand g05171(.dina(n430), .dinb(n1373), .dout(n5235));
  jand g05172(.dina(n5235), .dinb(n3950), .dout(n5236));
  jand g05173(.dina(n2698), .dinb(n1767), .dout(n5237));
  jand g05174(.dina(n5237), .dinb(n5236), .dout(n5238));
  jand g05175(.dina(n5238), .dinb(n5234), .dout(n5239));
  jand g05176(.dina(n3233), .dinb(n511), .dout(n5240));
  jand g05177(.dina(n5240), .dinb(n537), .dout(n5241));
  jand g05178(.dina(n1778), .dinb(n900), .dout(n5242));
  jand g05179(.dina(n5242), .dinb(n5241), .dout(n5243));
  jand g05180(.dina(n5243), .dinb(n5239), .dout(n5244));
  jand g05181(.dina(n1473), .dinb(n1304), .dout(n5245));
  jand g05182(.dina(n5245), .dinb(n5244), .dout(n5246));
  jand g05183(.dina(n4538), .dinb(n653), .dout(n5247));
  jand g05184(.dina(n447), .dinb(n1203), .dout(n5248));
  jand g05185(.dina(n920), .dinb(n1040), .dout(n5249));
  jand g05186(.dina(n5249), .dinb(n5248), .dout(n5250));
  jand g05187(.dina(n5250), .dinb(n5247), .dout(n5251));
  jand g05188(.dina(n1310), .dinb(n1257), .dout(n5252));
  jand g05189(.dina(n1465), .dinb(n1682), .dout(n5253));
  jand g05190(.dina(n848), .dinb(n621), .dout(n5254));
  jand g05191(.dina(n1218), .dinb(n270), .dout(n5255));
  jand g05192(.dina(n5255), .dinb(n5254), .dout(n5256));
  jand g05193(.dina(n5256), .dinb(n5253), .dout(n5257));
  jand g05194(.dina(n5257), .dinb(n5252), .dout(n5258));
  jand g05195(.dina(n1336), .dinb(n808), .dout(n5259));
  jand g05196(.dina(n5259), .dinb(n5258), .dout(n5260));
  jand g05197(.dina(n5260), .dinb(n5251), .dout(n5261));
  jand g05198(.dina(n5261), .dinb(n5246), .dout(n5262));
  jand g05199(.dina(n5262), .dinb(n5228), .dout(n5263));
  jand g05200(.dina(n5263), .dinb(n5193), .dout(n5264));
  jxor g05201(.dina(n5264), .dinb(n4686), .dout(n5265));
  jxor g05202(.dina(n5265), .dinb(n5168), .dout(n5266));
  jor  g05203(.dina(n5266), .dinb(n4692), .dout(n5267));
  jor  g05204(.dina(n4697), .dinb(n4686), .dout(n5268));
  jor  g05205(.dina(n4702), .dinb(n4526), .dout(n5269));
  jor  g05206(.dina(n5264), .dinb(n4705), .dout(n5270));
  jand g05207(.dina(n5270), .dinb(n5269), .dout(n5271));
  jand g05208(.dina(n5271), .dinb(n5268), .dout(n5272));
  jand g05209(.dina(n5272), .dinb(n5267), .dout(n5273));
  jxor g05210(.dina(n5273), .dinb(n4713), .dout(n5274));
  jxor g05211(.dina(n5274), .dinb(n5162), .dout(n5275));
  jxor g05212(.dina(n5275), .dinb(n5052), .dout(n5276));
  jnot g05213(.din(\a[5] ), .dout(n5277));
  jxor g05214(.dina(\a[5] ), .dinb(\a[4] ), .dout(n5278));
  jxor g05215(.dina(\a[3] ), .dinb(\a[2] ), .dout(n5279));
  jand g05216(.dina(n5279), .dinb(n5278), .dout(n5280));
  jnot g05217(.din(n5280), .dout(n5281));
  jand g05218(.dina(n1315), .dinb(n266), .dout(n5282));
  jand g05219(.dina(n654), .dinb(n135), .dout(n5283));
  jand g05220(.dina(n5283), .dinb(n5282), .dout(n5284));
  jand g05221(.dina(n1107), .dinb(n411), .dout(n5285));
  jand g05222(.dina(n632), .dinb(n1366), .dout(n5286));
  jand g05223(.dina(n5286), .dinb(n5285), .dout(n5287));
  jand g05224(.dina(n5287), .dinb(n1775), .dout(n5288));
  jand g05225(.dina(n5288), .dinb(n5284), .dout(n5289));
  jand g05226(.dina(n5289), .dinb(n982), .dout(n5290));
  jand g05227(.dina(n5290), .dinb(n2366), .dout(n5291));
  jand g05228(.dina(n2100), .dinb(n880), .dout(n5292));
  jand g05229(.dina(n5292), .dinb(n1306), .dout(n5293));
  jand g05230(.dina(n5293), .dinb(n1709), .dout(n5294));
  jand g05231(.dina(n3150), .dinb(n3065), .dout(n5295));
  jand g05232(.dina(n5295), .dinb(n5294), .dout(n5296));
  jand g05233(.dina(n5296), .dinb(n5291), .dout(n5297));
  jand g05234(.dina(n931), .dinb(n456), .dout(n5298));
  jand g05235(.dina(n3345), .dinb(n871), .dout(n5299));
  jand g05236(.dina(n5299), .dinb(n5298), .dout(n5300));
  jand g05237(.dina(n430), .dinb(n1283), .dout(n5301));
  jand g05238(.dina(n5301), .dinb(n3750), .dout(n5302));
  jand g05239(.dina(n5302), .dinb(n5300), .dout(n5303));
  jand g05240(.dina(n521), .dinb(n481), .dout(n5304));
  jand g05241(.dina(n5304), .dinb(n1522), .dout(n5305));
  jand g05242(.dina(n5305), .dinb(n1460), .dout(n5306));
  jand g05243(.dina(n1564), .dinb(n470), .dout(n5307));
  jand g05244(.dina(n5307), .dinb(n92), .dout(n5308));
  jand g05245(.dina(n5308), .dinb(n5306), .dout(n5309));
  jand g05246(.dina(n1532), .dinb(n537), .dout(n5310));
  jand g05247(.dina(n1190), .dinb(n991), .dout(n5311));
  jand g05248(.dina(n5311), .dinb(n1822), .dout(n5312));
  jand g05249(.dina(n5312), .dinb(n5310), .dout(n5313));
  jand g05250(.dina(n5313), .dinb(n5309), .dout(n5314));
  jand g05251(.dina(n1524), .dinb(n1361), .dout(n5315));
  jand g05252(.dina(n824), .dinb(n1270), .dout(n5316));
  jand g05253(.dina(n5316), .dinb(n5315), .dout(n5317));
  jand g05254(.dina(n5317), .dinb(n1917), .dout(n5318));
  jand g05255(.dina(n600), .dinb(n1351), .dout(n5319));
  jand g05256(.dina(n1238), .dinb(n82), .dout(n5320));
  jand g05257(.dina(n5320), .dinb(n1459), .dout(n5321));
  jand g05258(.dina(n5321), .dinb(n5319), .dout(n5322));
  jand g05259(.dina(n5322), .dinb(n5318), .dout(n5323));
  jand g05260(.dina(n5323), .dinb(n3044), .dout(n5324));
  jand g05261(.dina(n5324), .dinb(n5314), .dout(n5325));
  jand g05262(.dina(n5325), .dinb(n5303), .dout(n5326));
  jand g05263(.dina(n1451), .dinb(n1426), .dout(n5327));
  jand g05264(.dina(n5327), .dinb(n1259), .dout(n5328));
  jand g05265(.dina(n5328), .dinb(n1877), .dout(n5329));
  jand g05266(.dina(n1462), .dinb(n549), .dout(n5330));
  jand g05267(.dina(n5330), .dinb(n5329), .dout(n5331));
  jand g05268(.dina(n1732), .dinb(n122), .dout(n5332));
  jand g05269(.dina(n450), .dinb(n916), .dout(n5333));
  jand g05270(.dina(n5333), .dinb(n1868), .dout(n5334));
  jand g05271(.dina(n5334), .dinb(n5332), .dout(n5335));
  jand g05272(.dina(n3771), .dinb(n2529), .dout(n5336));
  jand g05273(.dina(n5336), .dinb(n5335), .dout(n5337));
  jand g05274(.dina(n5337), .dinb(n5331), .dout(n5338));
  jand g05275(.dina(n1162), .dinb(n1541), .dout(n5339));
  jand g05276(.dina(n5339), .dinb(n3195), .dout(n5340));
  jand g05277(.dina(n1698), .dinb(n1429), .dout(n5341));
  jand g05278(.dina(n5341), .dinb(n1415), .dout(n5342));
  jand g05279(.dina(n619), .dinb(n1203), .dout(n5343));
  jand g05280(.dina(n5343), .dinb(n1778), .dout(n5344));
  jand g05281(.dina(n5344), .dinb(n5342), .dout(n5345));
  jand g05282(.dina(n5345), .dinb(n5340), .dout(n5346));
  jand g05283(.dina(n5346), .dinb(n5338), .dout(n5347));
  jand g05284(.dina(n1536), .dinb(n1090), .dout(n5348));
  jand g05285(.dina(n5348), .dinb(n1365), .dout(n5349));
  jand g05286(.dina(n5349), .dinb(n716), .dout(n5350));
  jand g05287(.dina(n1037), .dinb(n516), .dout(n5351));
  jand g05288(.dina(n5351), .dinb(n1430), .dout(n5352));
  jand g05289(.dina(n5352), .dinb(n668), .dout(n5353));
  jand g05290(.dina(n454), .dinb(n168), .dout(n5354));
  jand g05291(.dina(n320), .dinb(n1245), .dout(n5355));
  jand g05292(.dina(n1453), .dinb(n829), .dout(n5356));
  jand g05293(.dina(n5356), .dinb(n5355), .dout(n5357));
  jand g05294(.dina(n5357), .dinb(n5354), .dout(n5358));
  jand g05295(.dina(n5358), .dinb(n5353), .dout(n5359));
  jand g05296(.dina(n5359), .dinb(n5350), .dout(n5360));
  jand g05297(.dina(n5360), .dinb(n1843), .dout(n5361));
  jand g05298(.dina(n5361), .dinb(n5347), .dout(n5362));
  jand g05299(.dina(n5362), .dinb(n5326), .dout(n5363));
  jand g05300(.dina(n5363), .dinb(n5297), .dout(n5364));
  jnot g05301(.din(n5364), .dout(n5365));
  jand g05302(.dina(n1449), .dinb(n178), .dout(n5366));
  jand g05303(.dina(n5366), .dinb(n921), .dout(n5367));
  jand g05304(.dina(n670), .dinb(n1325), .dout(n5368));
  jand g05305(.dina(n5368), .dinb(n2567), .dout(n5369));
  jand g05306(.dina(n3371), .dinb(n3178), .dout(n5370));
  jand g05307(.dina(n3980), .dinb(n816), .dout(n5371));
  jand g05308(.dina(n5371), .dinb(n5370), .dout(n5372));
  jand g05309(.dina(n5372), .dinb(n5369), .dout(n5373));
  jand g05310(.dina(n1843), .dinb(n1292), .dout(n5374));
  jand g05311(.dina(n1778), .dinb(n1495), .dout(n5375));
  jand g05312(.dina(n5375), .dinb(n2020), .dout(n5376));
  jand g05313(.dina(n5376), .dinb(n5374), .dout(n5377));
  jand g05314(.dina(n965), .dinb(n1309), .dout(n5378));
  jand g05315(.dina(n925), .dinb(n1226), .dout(n5379));
  jand g05316(.dina(n5379), .dinb(n5378), .dout(n5380));
  jand g05317(.dina(n5380), .dinb(n5377), .dout(n5381));
  jand g05318(.dina(n5381), .dinb(n5373), .dout(n5382));
  jand g05319(.dina(n5382), .dinb(n5367), .dout(n5383));
  jand g05320(.dina(n2620), .dinb(n1732), .dout(n5384));
  jand g05321(.dina(n2148), .dinb(n1375), .dout(n5385));
  jand g05322(.dina(n5385), .dinb(n5384), .dout(n5386));
  jand g05323(.dina(n4440), .dinb(n1163), .dout(n5387));
  jand g05324(.dina(n5387), .dinb(n5386), .dout(n5388));
  jand g05325(.dina(n647), .dinb(n1345), .dout(n5389));
  jand g05326(.dina(n1361), .dinb(n1351), .dout(n5390));
  jand g05327(.dina(n5390), .dinb(n2009), .dout(n5391));
  jand g05328(.dina(n5391), .dinb(n5389), .dout(n5392));
  jand g05329(.dina(n5392), .dinb(n5388), .dout(n5393));
  jand g05330(.dina(n1578), .dinb(n442), .dout(n5394));
  jand g05331(.dina(n472), .dinb(n82), .dout(n5395));
  jand g05332(.dina(n2100), .dinb(n848), .dout(n5396));
  jand g05333(.dina(n5396), .dinb(n5395), .dout(n5397));
  jand g05334(.dina(n5397), .dinb(n2385), .dout(n5398));
  jand g05335(.dina(n5398), .dinb(n5394), .dout(n5399));
  jand g05336(.dina(n5399), .dinb(n3827), .dout(n5400));
  jand g05337(.dina(n5400), .dinb(n5393), .dout(n5401));
  jand g05338(.dina(n5401), .dinb(n5383), .dout(n5402));
  jand g05339(.dina(n1037), .dinb(n715), .dout(n5403));
  jand g05340(.dina(n1454), .dinb(n1738), .dout(n5404));
  jand g05341(.dina(n5404), .dinb(n1900), .dout(n5405));
  jand g05342(.dina(n5405), .dinb(n5403), .dout(n5406));
  jand g05343(.dina(n5406), .dinb(n1540), .dout(n5407));
  jand g05344(.dina(n411), .dinb(n1245), .dout(n5408));
  jand g05345(.dina(n5408), .dinb(n1565), .dout(n5409));
  jand g05346(.dina(n5409), .dinb(n2409), .dout(n5410));
  jand g05347(.dina(n1701), .dinb(n171), .dout(n5411));
  jand g05348(.dina(n5411), .dinb(n1915), .dout(n5412));
  jand g05349(.dina(n5412), .dinb(n1559), .dout(n5413));
  jand g05350(.dina(n5413), .dinb(n5410), .dout(n5414));
  jand g05351(.dina(n456), .dinb(n638), .dout(n5415));
  jand g05352(.dina(n2357), .dinb(n1229), .dout(n5416));
  jand g05353(.dina(n5416), .dinb(n5415), .dout(n5417));
  jand g05354(.dina(n5417), .dinb(n1755), .dout(n5418));
  jand g05355(.dina(n5418), .dinb(n5414), .dout(n5419));
  jand g05356(.dina(n5419), .dinb(n5407), .dout(n5420));
  jand g05357(.dina(n5420), .dinb(n2471), .dout(n5421));
  jand g05358(.dina(n5421), .dinb(n5402), .dout(n5422));
  jnot g05359(.din(n5422), .dout(n5423));
  jand g05360(.dina(n5423), .dinb(n5365), .dout(n5424));
  jnot g05361(.din(n5424), .dout(n5425));
  jnot g05362(.din(n5264), .dout(n5426));
  jand g05363(.dina(n5423), .dinb(n5426), .dout(n5427));
  jnot g05364(.din(n5427), .dout(n5428));
  jand g05365(.dina(n5426), .dinb(n5163), .dout(n5429));
  jnot g05366(.din(n5429), .dout(n5430));
  jnot g05367(.din(n5265), .dout(n5431));
  jor  g05368(.dina(n5431), .dinb(n5168), .dout(n5432));
  jand g05369(.dina(n5432), .dinb(n5430), .dout(n5433));
  jxor g05370(.dina(n5422), .dinb(n5264), .dout(n5434));
  jnot g05371(.din(n5434), .dout(n5435));
  jor  g05372(.dina(n5435), .dinb(n5433), .dout(n5436));
  jand g05373(.dina(n5436), .dinb(n5428), .dout(n5437));
  jxor g05374(.dina(n5422), .dinb(n5364), .dout(n5438));
  jnot g05375(.din(n5438), .dout(n5439));
  jor  g05376(.dina(n5439), .dinb(n5437), .dout(n5440));
  jand g05377(.dina(n5440), .dinb(n5425), .dout(n5441));
  jand g05378(.dina(n3762), .dinb(n551), .dout(n5442));
  jand g05379(.dina(n2600), .dinb(n1206), .dout(n5443));
  jand g05380(.dina(n5443), .dinb(n5442), .dout(n5444));
  jand g05381(.dina(n5444), .dinb(n1698), .dout(n5445));
  jand g05382(.dina(n5445), .dinb(n4659), .dout(n5446));
  jand g05383(.dina(n521), .dinb(n499), .dout(n5447));
  jand g05384(.dina(n5447), .dinb(n5231), .dout(n5448));
  jand g05385(.dina(n5448), .dinb(n1852), .dout(n5449));
  jand g05386(.dina(n1756), .dinb(n1283), .dout(n5450));
  jand g05387(.dina(n5450), .dinb(n2366), .dout(n5451));
  jand g05388(.dina(n5451), .dinb(n1367), .dout(n5452));
  jand g05389(.dina(n5452), .dinb(n5449), .dout(n5453));
  jand g05390(.dina(n3847), .dinb(n1325), .dout(n5454));
  jand g05391(.dina(n5454), .dinb(n4590), .dout(n5455));
  jand g05392(.dina(n993), .dinb(n988), .dout(n5456));
  jand g05393(.dina(n5456), .dinb(n1936), .dout(n5457));
  jand g05394(.dina(n5457), .dinb(n5396), .dout(n5458));
  jand g05395(.dina(n5458), .dinb(n5455), .dout(n5459));
  jand g05396(.dina(n5459), .dinb(n5453), .dout(n5460));
  jand g05397(.dina(n5460), .dinb(n5446), .dout(n5461));
  jand g05398(.dina(n4417), .dinb(n811), .dout(n5462));
  jand g05399(.dina(n5462), .dinb(n680), .dout(n5463));
  jand g05400(.dina(n2444), .dinb(n445), .dout(n5464));
  jand g05401(.dina(n1822), .dinb(n463), .dout(n5465));
  jand g05402(.dina(n5465), .dinb(n1495), .dout(n5466));
  jand g05403(.dina(n5466), .dinb(n5464), .dout(n5467));
  jand g05404(.dina(n5467), .dinb(n5463), .dout(n5468));
  jand g05405(.dina(n1716), .dinb(n1713), .dout(n5469));
  jand g05406(.dina(n5469), .dinb(n1309), .dout(n5470));
  jand g05407(.dina(n5470), .dinb(n5468), .dout(n5471));
  jand g05408(.dina(n5471), .dinb(n5461), .dout(n5472));
  jand g05409(.dina(n1426), .dinb(n1560), .dout(n5473));
  jand g05410(.dina(n5473), .dinb(n555), .dout(n5474));
  jand g05411(.dina(n696), .dinb(n510), .dout(n5475));
  jand g05412(.dina(n5475), .dinb(n1968), .dout(n5476));
  jand g05413(.dina(n5476), .dinb(n3900), .dout(n5477));
  jand g05414(.dina(n5477), .dinb(n5474), .dout(n5478));
  jand g05415(.dina(n664), .dinb(n808), .dout(n5479));
  jand g05416(.dina(n5479), .dinb(n909), .dout(n5480));
  jand g05417(.dina(n4669), .dinb(n108), .dout(n5481));
  jand g05418(.dina(n5481), .dinb(n5480), .dout(n5482));
  jand g05419(.dina(n4448), .dinb(n3978), .dout(n5483));
  jand g05420(.dina(n5483), .dinb(n2586), .dout(n5484));
  jand g05421(.dina(n5484), .dinb(n5482), .dout(n5485));
  jand g05422(.dina(n5485), .dinb(n5478), .dout(n5486));
  jand g05423(.dina(n1721), .dinb(n950), .dout(n5487));
  jand g05424(.dina(n2716), .dinb(n1987), .dout(n5488));
  jand g05425(.dina(n5488), .dinb(n4668), .dout(n5489));
  jand g05426(.dina(n5489), .dinb(n5487), .dout(n5490));
  jand g05427(.dina(n2372), .dinb(n1366), .dout(n5491));
  jand g05428(.dina(n5491), .dinb(n1903), .dout(n5492));
  jand g05429(.dina(n1743), .dinb(n1515), .dout(n5493));
  jand g05430(.dina(n5493), .dinb(n1308), .dout(n5494));
  jand g05431(.dina(n5494), .dinb(n4496), .dout(n5495));
  jand g05432(.dina(n5495), .dinb(n5492), .dout(n5496));
  jand g05433(.dina(n5496), .dinb(n5490), .dout(n5497));
  jand g05434(.dina(n5497), .dinb(n5486), .dout(n5498));
  jand g05435(.dina(n632), .dinb(n1233), .dout(n5499));
  jand g05436(.dina(n5499), .dinb(n954), .dout(n5500));
  jand g05437(.dina(n562), .dinb(n442), .dout(n5501));
  jand g05438(.dina(n1682), .dinb(n1036), .dout(n5502));
  jand g05439(.dina(n5502), .dinb(n5501), .dout(n5503));
  jand g05440(.dina(n5503), .dinb(n5500), .dout(n5504));
  jand g05441(.dina(n1506), .dinb(n670), .dout(n5505));
  jand g05442(.dina(n5505), .dinb(n1160), .dout(n5506));
  jand g05443(.dina(n5171), .dinb(n1245), .dout(n5507));
  jand g05444(.dina(n5507), .dinb(n5506), .dout(n5508));
  jand g05445(.dina(n5508), .dinb(n5504), .dout(n5509));
  jand g05446(.dina(n5220), .dinb(n2701), .dout(n5510));
  jand g05447(.dina(n1037), .dinb(n469), .dout(n5511));
  jand g05448(.dina(n5511), .dinb(n1536), .dout(n5512));
  jand g05449(.dina(n5512), .dinb(n1686), .dout(n5513));
  jand g05450(.dina(n5513), .dinb(n5510), .dout(n5514));
  jand g05451(.dina(n1731), .dinb(n532), .dout(n5515));
  jand g05452(.dina(n5515), .dinb(n650), .dout(n5516));
  jand g05453(.dina(n5516), .dinb(n3264), .dout(n5517));
  jand g05454(.dina(n693), .dinb(n676), .dout(n5518));
  jand g05455(.dina(n2588), .dinb(n907), .dout(n5519));
  jand g05456(.dina(n5519), .dinb(n5518), .dout(n5520));
  jand g05457(.dina(n5520), .dinb(n5517), .dout(n5521));
  jand g05458(.dina(n5521), .dinb(n5514), .dout(n5522));
  jand g05459(.dina(n5522), .dinb(n5509), .dout(n5523));
  jand g05460(.dina(n5523), .dinb(n5498), .dout(n5524));
  jand g05461(.dina(n5524), .dinb(n5472), .dout(n5525));
  jxor g05462(.dina(n5525), .dinb(n5364), .dout(n5526));
  jxor g05463(.dina(n5526), .dinb(n5441), .dout(n5527));
  jor  g05464(.dina(n5527), .dinb(n5281), .dout(n5528));
  jnot g05465(.din(n5279), .dout(n5529));
  jxor g05466(.dina(\a[4] ), .dinb(\a[3] ), .dout(n5530));
  jand g05467(.dina(n5530), .dinb(n5529), .dout(n5531));
  jnot g05468(.din(n5531), .dout(n5532));
  jor  g05469(.dina(n5532), .dinb(n5364), .dout(n5533));
  jor  g05470(.dina(n5530), .dinb(n5279), .dout(n5534));
  jnot g05471(.din(n5534), .dout(n5535));
  jand g05472(.dina(n5535), .dinb(n5278), .dout(n5536));
  jnot g05473(.din(n5536), .dout(n5537));
  jor  g05474(.dina(n5537), .dinb(n5422), .dout(n5538));
  jor  g05475(.dina(n5529), .dinb(n5278), .dout(n5539));
  jor  g05476(.dina(n5539), .dinb(n5525), .dout(n5540));
  jand g05477(.dina(n5540), .dinb(n5538), .dout(n5541));
  jand g05478(.dina(n5541), .dinb(n5533), .dout(n5542));
  jand g05479(.dina(n5542), .dinb(n5528), .dout(n5543));
  jxor g05480(.dina(n5543), .dinb(n5277), .dout(n5544));
  jand g05481(.dina(n5544), .dinb(n5276), .dout(n5545));
  jnot g05482(.din(n5545), .dout(n5546));
  jxor g05483(.dina(n5050), .dinb(n5049), .dout(n5547));
  jnot g05484(.din(n5547), .dout(n5548));
  jxor g05485(.dina(n5438), .dinb(n5437), .dout(n5549));
  jor  g05486(.dina(n5549), .dinb(n5281), .dout(n5550));
  jor  g05487(.dina(n5532), .dinb(n5422), .dout(n5551));
  jor  g05488(.dina(n5537), .dinb(n5264), .dout(n5552));
  jand g05489(.dina(n5552), .dinb(n5551), .dout(n5553));
  jor  g05490(.dina(n5539), .dinb(n5364), .dout(n5554));
  jand g05491(.dina(n5554), .dinb(n5553), .dout(n5555));
  jand g05492(.dina(n5555), .dinb(n5550), .dout(n5556));
  jxor g05493(.dina(n5556), .dinb(\a[5] ), .dout(n5557));
  jor  g05494(.dina(n5557), .dinb(n5548), .dout(n5558));
  jxor g05495(.dina(n5047), .dinb(n5046), .dout(n5559));
  jxor g05496(.dina(n5434), .dinb(n5433), .dout(n5560));
  jor  g05497(.dina(n5560), .dinb(n5281), .dout(n5561));
  jor  g05498(.dina(n5532), .dinb(n5264), .dout(n5562));
  jor  g05499(.dina(n5539), .dinb(n5422), .dout(n5563));
  jor  g05500(.dina(n5537), .dinb(n4686), .dout(n5564));
  jand g05501(.dina(n5564), .dinb(n5563), .dout(n5565));
  jand g05502(.dina(n5565), .dinb(n5562), .dout(n5566));
  jand g05503(.dina(n5566), .dinb(n5561), .dout(n5567));
  jxor g05504(.dina(n5567), .dinb(n5277), .dout(n5568));
  jand g05505(.dina(n5568), .dinb(n5559), .dout(n5569));
  jxor g05506(.dina(n5044), .dinb(n5042), .dout(n5570));
  jor  g05507(.dina(n5281), .dinb(n5266), .dout(n5571));
  jor  g05508(.dina(n5532), .dinb(n4686), .dout(n5572));
  jor  g05509(.dina(n5537), .dinb(n4526), .dout(n5573));
  jor  g05510(.dina(n5539), .dinb(n5264), .dout(n5574));
  jand g05511(.dina(n5574), .dinb(n5573), .dout(n5575));
  jand g05512(.dina(n5575), .dinb(n5572), .dout(n5576));
  jand g05513(.dina(n5576), .dinb(n5571), .dout(n5577));
  jxor g05514(.dina(n5577), .dinb(n5277), .dout(n5578));
  jand g05515(.dina(n5578), .dinb(n5570), .dout(n5579));
  jxor g05516(.dina(n5040), .dinb(n5038), .dout(n5580));
  jnot g05517(.din(n5580), .dout(n5581));
  jor  g05518(.dina(n5281), .dinb(n4688), .dout(n5582));
  jor  g05519(.dina(n5532), .dinb(n4526), .dout(n5583));
  jor  g05520(.dina(n5539), .dinb(n4686), .dout(n5584));
  jand g05521(.dina(n5584), .dinb(n5583), .dout(n5585));
  jor  g05522(.dina(n5537), .dinb(n4596), .dout(n5586));
  jand g05523(.dina(n5586), .dinb(n5585), .dout(n5587));
  jand g05524(.dina(n5587), .dinb(n5582), .dout(n5588));
  jxor g05525(.dina(n5588), .dinb(\a[5] ), .dout(n5589));
  jor  g05526(.dina(n5589), .dinb(n5581), .dout(n5590));
  jnot g05527(.din(n5590), .dout(n5591));
  jxor g05528(.dina(n5036), .dinb(n5035), .dout(n5592));
  jor  g05529(.dina(n5281), .dinb(n4714), .dout(n5593));
  jor  g05530(.dina(n5532), .dinb(n4596), .dout(n5594));
  jor  g05531(.dina(n5537), .dinb(n4471), .dout(n5595));
  jor  g05532(.dina(n5539), .dinb(n4526), .dout(n5596));
  jand g05533(.dina(n5596), .dinb(n5595), .dout(n5597));
  jand g05534(.dina(n5597), .dinb(n5594), .dout(n5598));
  jand g05535(.dina(n5598), .dinb(n5593), .dout(n5599));
  jxor g05536(.dina(n5599), .dinb(n5277), .dout(n5600));
  jand g05537(.dina(n5600), .dinb(n5592), .dout(n5601));
  jxor g05538(.dina(n5032), .dinb(n5031), .dout(n5602));
  jnot g05539(.din(n5602), .dout(n5603));
  jor  g05540(.dina(n5281), .dinb(n4726), .dout(n5604));
  jor  g05541(.dina(n5532), .dinb(n4471), .dout(n5605));
  jor  g05542(.dina(n5537), .dinb(n4019), .dout(n5606));
  jor  g05543(.dina(n5539), .dinb(n4596), .dout(n5607));
  jand g05544(.dina(n5607), .dinb(n5606), .dout(n5608));
  jand g05545(.dina(n5608), .dinb(n5605), .dout(n5609));
  jand g05546(.dina(n5609), .dinb(n5604), .dout(n5610));
  jxor g05547(.dina(n5610), .dinb(n5277), .dout(n5611));
  jand g05548(.dina(n5611), .dinb(n5603), .dout(n5612));
  jxor g05549(.dina(n5029), .dinb(n5028), .dout(n5613));
  jor  g05550(.dina(n5281), .dinb(n4473), .dout(n5614));
  jor  g05551(.dina(n5532), .dinb(n4019), .dout(n5615));
  jor  g05552(.dina(n5537), .dinb(n3929), .dout(n5616));
  jor  g05553(.dina(n5539), .dinb(n4471), .dout(n5617));
  jand g05554(.dina(n5617), .dinb(n5616), .dout(n5618));
  jand g05555(.dina(n5618), .dinb(n5615), .dout(n5619));
  jand g05556(.dina(n5619), .dinb(n5614), .dout(n5620));
  jxor g05557(.dina(n5620), .dinb(n5277), .dout(n5621));
  jand g05558(.dina(n5621), .dinb(n5613), .dout(n5622));
  jxor g05559(.dina(n5026), .dinb(n5025), .dout(n5623));
  jor  g05560(.dina(n5281), .dinb(n4021), .dout(n5624));
  jor  g05561(.dina(n5532), .dinb(n3929), .dout(n5625));
  jor  g05562(.dina(n5539), .dinb(n4019), .dout(n5626));
  jor  g05563(.dina(n5537), .dinb(n3863), .dout(n5627));
  jand g05564(.dina(n5627), .dinb(n5626), .dout(n5628));
  jand g05565(.dina(n5628), .dinb(n5625), .dout(n5629));
  jand g05566(.dina(n5629), .dinb(n5624), .dout(n5630));
  jxor g05567(.dina(n5630), .dinb(n5277), .dout(n5631));
  jand g05568(.dina(n5631), .dinb(n5623), .dout(n5632));
  jxor g05569(.dina(n5023), .dinb(n5022), .dout(n5633));
  jnot g05570(.din(n5633), .dout(n5634));
  jor  g05571(.dina(n5281), .dinb(n4038), .dout(n5635));
  jor  g05572(.dina(n5532), .dinb(n3863), .dout(n5636));
  jor  g05573(.dina(n5539), .dinb(n3929), .dout(n5637));
  jand g05574(.dina(n5637), .dinb(n5636), .dout(n5638));
  jor  g05575(.dina(n5537), .dinb(n3787), .dout(n5639));
  jand g05576(.dina(n5639), .dinb(n5638), .dout(n5640));
  jand g05577(.dina(n5640), .dinb(n5635), .dout(n5641));
  jxor g05578(.dina(n5641), .dinb(\a[5] ), .dout(n5642));
  jor  g05579(.dina(n5642), .dinb(n5634), .dout(n5643));
  jnot g05580(.din(n5643), .dout(n5644));
  jxor g05581(.dina(n5020), .dinb(n5018), .dout(n5645));
  jor  g05582(.dina(n5281), .dinb(n4051), .dout(n5646));
  jor  g05583(.dina(n5532), .dinb(n3787), .dout(n5647));
  jor  g05584(.dina(n5539), .dinb(n3863), .dout(n5648));
  jor  g05585(.dina(n5537), .dinb(n3420), .dout(n5649));
  jand g05586(.dina(n5649), .dinb(n5648), .dout(n5650));
  jand g05587(.dina(n5650), .dinb(n5647), .dout(n5651));
  jand g05588(.dina(n5651), .dinb(n5646), .dout(n5652));
  jxor g05589(.dina(n5652), .dinb(n5277), .dout(n5653));
  jand g05590(.dina(n5653), .dinb(n5645), .dout(n5654));
  jxor g05591(.dina(n5016), .dinb(n5014), .dout(n5655));
  jnot g05592(.din(n5655), .dout(n5656));
  jor  g05593(.dina(n5281), .dinb(n3789), .dout(n5657));
  jor  g05594(.dina(n5532), .dinb(n3420), .dout(n5658));
  jor  g05595(.dina(n5537), .dinb(n3286), .dout(n5659));
  jand g05596(.dina(n5659), .dinb(n5658), .dout(n5660));
  jor  g05597(.dina(n5539), .dinb(n3787), .dout(n5661));
  jand g05598(.dina(n5661), .dinb(n5660), .dout(n5662));
  jand g05599(.dina(n5662), .dinb(n5657), .dout(n5663));
  jxor g05600(.dina(n5663), .dinb(\a[5] ), .dout(n5664));
  jor  g05601(.dina(n5664), .dinb(n5656), .dout(n5665));
  jnot g05602(.din(n5665), .dout(n5666));
  jxor g05603(.dina(n5012), .dinb(n5010), .dout(n5667));
  jnot g05604(.din(n5667), .dout(n5668));
  jor  g05605(.dina(n5537), .dinb(n3203), .dout(n5669));
  jor  g05606(.dina(n5281), .dinb(n3422), .dout(n5670));
  jor  g05607(.dina(n5539), .dinb(n3420), .dout(n5671));
  jor  g05608(.dina(n5532), .dinb(n3286), .dout(n5672));
  jand g05609(.dina(n5672), .dinb(n5671), .dout(n5673));
  jand g05610(.dina(n5673), .dinb(n5670), .dout(n5674));
  jand g05611(.dina(n5674), .dinb(n5669), .dout(n5675));
  jxor g05612(.dina(n5675), .dinb(\a[5] ), .dout(n5676));
  jor  g05613(.dina(n5676), .dinb(n5668), .dout(n5677));
  jnot g05614(.din(n5677), .dout(n5678));
  jxor g05615(.dina(n5008), .dinb(n5006), .dout(n5679));
  jor  g05616(.dina(n5281), .dinb(n3440), .dout(n5680));
  jor  g05617(.dina(n5532), .dinb(n3203), .dout(n5681));
  jor  g05618(.dina(n5539), .dinb(n3286), .dout(n5682));
  jand g05619(.dina(n5682), .dinb(n5681), .dout(n5683));
  jor  g05620(.dina(n5537), .dinb(n3072), .dout(n5684));
  jand g05621(.dina(n5684), .dinb(n5683), .dout(n5685));
  jand g05622(.dina(n5685), .dinb(n5680), .dout(n5686));
  jxor g05623(.dina(n5686), .dinb(\a[5] ), .dout(n5687));
  jor  g05624(.dina(n5687), .dinb(n5679), .dout(n5688));
  jxor g05625(.dina(n5004), .dinb(n5002), .dout(n5689));
  jnot g05626(.din(n5689), .dout(n5690));
  jor  g05627(.dina(n5281), .dinb(n3451), .dout(n5691));
  jor  g05628(.dina(n5532), .dinb(n3072), .dout(n5692));
  jor  g05629(.dina(n5537), .dinb(n2738), .dout(n5693));
  jand g05630(.dina(n5693), .dinb(n5692), .dout(n5694));
  jor  g05631(.dina(n5539), .dinb(n3203), .dout(n5695));
  jand g05632(.dina(n5695), .dinb(n5694), .dout(n5696));
  jand g05633(.dina(n5696), .dinb(n5691), .dout(n5697));
  jxor g05634(.dina(n5697), .dinb(\a[5] ), .dout(n5698));
  jor  g05635(.dina(n5698), .dinb(n5690), .dout(n5699));
  jxor g05636(.dina(n5000), .dinb(n4998), .dout(n5700));
  jor  g05637(.dina(n5281), .dinb(n3081), .dout(n5701));
  jor  g05638(.dina(n5537), .dinb(n2553), .dout(n5702));
  jor  g05639(.dina(n5532), .dinb(n2738), .dout(n5703));
  jor  g05640(.dina(n5539), .dinb(n3072), .dout(n5704));
  jand g05641(.dina(n5704), .dinb(n5703), .dout(n5705));
  jand g05642(.dina(n5705), .dinb(n5702), .dout(n5706));
  jand g05643(.dina(n5706), .dinb(n5701), .dout(n5707));
  jxor g05644(.dina(n5707), .dinb(n5277), .dout(n5708));
  jand g05645(.dina(n5708), .dinb(n5700), .dout(n5709));
  jnot g05646(.din(n5709), .dout(n5710));
  jxor g05647(.dina(n4996), .dinb(n4994), .dout(n5711));
  jor  g05648(.dina(n5281), .dinb(n2740), .dout(n5712));
  jor  g05649(.dina(n5532), .dinb(n2553), .dout(n5713));
  jor  g05650(.dina(n5537), .dinb(n2629), .dout(n5714));
  jor  g05651(.dina(n5539), .dinb(n2738), .dout(n5715));
  jand g05652(.dina(n5715), .dinb(n5714), .dout(n5716));
  jand g05653(.dina(n5716), .dinb(n5713), .dout(n5717));
  jand g05654(.dina(n5717), .dinb(n5712), .dout(n5718));
  jxor g05655(.dina(n5718), .dinb(n5277), .dout(n5719));
  jand g05656(.dina(n5719), .dinb(n5711), .dout(n5720));
  jnot g05657(.din(n5720), .dout(n5721));
  jxor g05658(.dina(n4992), .dinb(n4990), .dout(n5722));
  jor  g05659(.dina(n5281), .dinb(n2768), .dout(n5723));
  jor  g05660(.dina(n5539), .dinb(n2553), .dout(n5724));
  jor  g05661(.dina(n5537), .dinb(n2428), .dout(n5725));
  jor  g05662(.dina(n5532), .dinb(n2629), .dout(n5726));
  jand g05663(.dina(n5726), .dinb(n5725), .dout(n5727));
  jand g05664(.dina(n5727), .dinb(n5724), .dout(n5728));
  jand g05665(.dina(n5728), .dinb(n5723), .dout(n5729));
  jxor g05666(.dina(n5729), .dinb(n5277), .dout(n5730));
  jand g05667(.dina(n5730), .dinb(n5722), .dout(n5731));
  jnot g05668(.din(n5731), .dout(n5732));
  jxor g05669(.dina(n4988), .dinb(n4986), .dout(n5733));
  jnot g05670(.din(n5733), .dout(n5734));
  jor  g05671(.dina(n5537), .dinb(n2174), .dout(n5735));
  jor  g05672(.dina(n5281), .dinb(n2779), .dout(n5736));
  jor  g05673(.dina(n5539), .dinb(n2629), .dout(n5737));
  jor  g05674(.dina(n5532), .dinb(n2428), .dout(n5738));
  jand g05675(.dina(n5738), .dinb(n5737), .dout(n5739));
  jand g05676(.dina(n5739), .dinb(n5736), .dout(n5740));
  jand g05677(.dina(n5740), .dinb(n5735), .dout(n5741));
  jxor g05678(.dina(n5741), .dinb(\a[5] ), .dout(n5742));
  jor  g05679(.dina(n5742), .dinb(n5734), .dout(n5743));
  jxor g05680(.dina(n4984), .dinb(n4982), .dout(n5744));
  jor  g05681(.dina(n5281), .dinb(n2430), .dout(n5745));
  jor  g05682(.dina(n5532), .dinb(n2174), .dout(n5746));
  jor  g05683(.dina(n5539), .dinb(n2428), .dout(n5747));
  jor  g05684(.dina(n5537), .dinb(n1954), .dout(n5748));
  jand g05685(.dina(n5748), .dinb(n5747), .dout(n5749));
  jand g05686(.dina(n5749), .dinb(n5746), .dout(n5750));
  jand g05687(.dina(n5750), .dinb(n5745), .dout(n5751));
  jxor g05688(.dina(n5751), .dinb(n5277), .dout(n5752));
  jand g05689(.dina(n5752), .dinb(n5744), .dout(n5753));
  jnot g05690(.din(n5753), .dout(n5754));
  jxor g05691(.dina(n4980), .dinb(n4978), .dout(n5755));
  jnot g05692(.din(n5755), .dout(n5756));
  jor  g05693(.dina(n5281), .dinb(n2176), .dout(n5757));
  jor  g05694(.dina(n5532), .dinb(n1954), .dout(n5758));
  jor  g05695(.dina(n5537), .dinb(n2057), .dout(n5759));
  jand g05696(.dina(n5759), .dinb(n5758), .dout(n5760));
  jor  g05697(.dina(n5539), .dinb(n2174), .dout(n5761));
  jand g05698(.dina(n5761), .dinb(n5760), .dout(n5762));
  jand g05699(.dina(n5762), .dinb(n5757), .dout(n5763));
  jxor g05700(.dina(n5763), .dinb(\a[5] ), .dout(n5764));
  jor  g05701(.dina(n5764), .dinb(n5756), .dout(n5765));
  jxor g05702(.dina(n4975), .dinb(n4974), .dout(n5766));
  jor  g05703(.dina(n5281), .dinb(n2197), .dout(n5767));
  jor  g05704(.dina(n5537), .dinb(n1790), .dout(n5768));
  jor  g05705(.dina(n5539), .dinb(n1954), .dout(n5769));
  jor  g05706(.dina(n5532), .dinb(n2057), .dout(n5770));
  jand g05707(.dina(n5770), .dinb(n5769), .dout(n5771));
  jand g05708(.dina(n5771), .dinb(n5768), .dout(n5772));
  jand g05709(.dina(n5772), .dinb(n5767), .dout(n5773));
  jxor g05710(.dina(n5773), .dinb(n5277), .dout(n5774));
  jand g05711(.dina(n5774), .dinb(n5766), .dout(n5775));
  jnot g05712(.din(n5775), .dout(n5776));
  jxor g05713(.dina(n4971), .dinb(n4963), .dout(n5777));
  jnot g05714(.din(n5777), .dout(n5778));
  jor  g05715(.dina(n5281), .dinb(n2208), .dout(n5779));
  jor  g05716(.dina(n5532), .dinb(n1790), .dout(n5780));
  jor  g05717(.dina(n5539), .dinb(n2057), .dout(n5781));
  jand g05718(.dina(n5781), .dinb(n5780), .dout(n5782));
  jor  g05719(.dina(n5537), .dinb(n1606), .dout(n5783));
  jand g05720(.dina(n5783), .dinb(n5782), .dout(n5784));
  jand g05721(.dina(n5784), .dinb(n5779), .dout(n5785));
  jxor g05722(.dina(n5785), .dinb(\a[5] ), .dout(n5786));
  jor  g05723(.dina(n5786), .dinb(n5778), .dout(n5787));
  jor  g05724(.dina(n5281), .dinb(n1792), .dout(n5788));
  jor  g05725(.dina(n5539), .dinb(n1790), .dout(n5789));
  jor  g05726(.dina(n5537), .dinb(n1448), .dout(n5790));
  jor  g05727(.dina(n5532), .dinb(n1606), .dout(n5791));
  jand g05728(.dina(n5791), .dinb(n5790), .dout(n5792));
  jand g05729(.dina(n5792), .dinb(n5789), .dout(n5793));
  jand g05730(.dina(n5793), .dinb(n5788), .dout(n5794));
  jxor g05731(.dina(n5794), .dinb(n5277), .dout(n5795));
  jor  g05732(.dina(n4950), .dinb(n4713), .dout(n5796));
  jxor g05733(.dina(n5796), .dinb(n4958), .dout(n5797));
  jand g05734(.dina(n5797), .dinb(n5795), .dout(n5798));
  jnot g05735(.din(n5798), .dout(n5799));
  jand g05736(.dina(n4947), .dinb(\a[8] ), .dout(n5800));
  jxor g05737(.dina(n5800), .dinb(n4945), .dout(n5801));
  jnot g05738(.din(n5801), .dout(n5802));
  jor  g05739(.dina(n5281), .dinb(n1608), .dout(n5803));
  jor  g05740(.dina(n5532), .dinb(n1448), .dout(n5804));
  jor  g05741(.dina(n5537), .dinb(n1255), .dout(n5805));
  jand g05742(.dina(n5805), .dinb(n5804), .dout(n5806));
  jor  g05743(.dina(n5539), .dinb(n1606), .dout(n5807));
  jand g05744(.dina(n5807), .dinb(n5806), .dout(n5808));
  jand g05745(.dina(n5808), .dinb(n5803), .dout(n5809));
  jxor g05746(.dina(n5809), .dinb(\a[5] ), .dout(n5810));
  jor  g05747(.dina(n5810), .dinb(n5802), .dout(n5811));
  jor  g05748(.dina(n5281), .dinb(n727), .dout(n5812));
  jand g05749(.dina(n5531), .dinb(n438), .dout(n5813));
  jnot g05750(.din(n5539), .dout(n5814));
  jand g05751(.dina(n5814), .dinb(n795), .dout(n5815));
  jor  g05752(.dina(n5815), .dinb(n5813), .dout(n5816));
  jnot g05753(.din(n5816), .dout(n5817));
  jand g05754(.dina(n5817), .dinb(n5812), .dout(n5818));
  jand g05755(.dina(n5279), .dinb(n438), .dout(n5819));
  jnot g05756(.din(n5819), .dout(n5820));
  jand g05757(.dina(n5820), .dinb(\a[5] ), .dout(n5821));
  jand g05758(.dina(n5821), .dinb(n5818), .dout(n5822));
  jand g05759(.dina(n5280), .dinb(n1639), .dout(n5823));
  jand g05760(.dina(n5531), .dinb(n795), .dout(n5824));
  jand g05761(.dina(n5814), .dinb(n1175), .dout(n5825));
  jor  g05762(.dina(n5825), .dinb(n5824), .dout(n5826));
  jand g05763(.dina(n5536), .dinb(n438), .dout(n5827));
  jor  g05764(.dina(n5827), .dinb(n5826), .dout(n5828));
  jor  g05765(.dina(n5828), .dinb(n5823), .dout(n5829));
  jnot g05766(.din(n5829), .dout(n5830));
  jand g05767(.dina(n5830), .dinb(n5822), .dout(n5831));
  jand g05768(.dina(n5831), .dinb(n4947), .dout(n5832));
  jnot g05769(.din(n5832), .dout(n5833));
  jxor g05770(.dina(n5831), .dinb(n4947), .dout(n5834));
  jnot g05771(.din(n5834), .dout(n5835));
  jor  g05772(.dina(n5281), .dinb(n1656), .dout(n5836));
  jor  g05773(.dina(n5539), .dinb(n1448), .dout(n5837));
  jor  g05774(.dina(n5532), .dinb(n1255), .dout(n5838));
  jand g05775(.dina(n5838), .dinb(n5837), .dout(n5839));
  jor  g05776(.dina(n5537), .dinb(n726), .dout(n5840));
  jand g05777(.dina(n5840), .dinb(n5839), .dout(n5841));
  jand g05778(.dina(n5841), .dinb(n5836), .dout(n5842));
  jxor g05779(.dina(n5842), .dinb(\a[5] ), .dout(n5843));
  jor  g05780(.dina(n5843), .dinb(n5835), .dout(n5844));
  jand g05781(.dina(n5844), .dinb(n5833), .dout(n5845));
  jxor g05782(.dina(n5810), .dinb(n5802), .dout(n5846));
  jnot g05783(.din(n5846), .dout(n5847));
  jor  g05784(.dina(n5847), .dinb(n5845), .dout(n5848));
  jand g05785(.dina(n5848), .dinb(n5811), .dout(n5849));
  jxor g05786(.dina(n5797), .dinb(n5795), .dout(n5850));
  jnot g05787(.din(n5850), .dout(n5851));
  jor  g05788(.dina(n5851), .dinb(n5849), .dout(n5852));
  jand g05789(.dina(n5852), .dinb(n5799), .dout(n5853));
  jxor g05790(.dina(n5786), .dinb(n5778), .dout(n5854));
  jnot g05791(.din(n5854), .dout(n5855));
  jor  g05792(.dina(n5855), .dinb(n5853), .dout(n5856));
  jand g05793(.dina(n5856), .dinb(n5787), .dout(n5857));
  jxor g05794(.dina(n5774), .dinb(n5766), .dout(n5858));
  jnot g05795(.din(n5858), .dout(n5859));
  jor  g05796(.dina(n5859), .dinb(n5857), .dout(n5860));
  jand g05797(.dina(n5860), .dinb(n5776), .dout(n5861));
  jxor g05798(.dina(n5764), .dinb(n5756), .dout(n5862));
  jnot g05799(.din(n5862), .dout(n5863));
  jor  g05800(.dina(n5863), .dinb(n5861), .dout(n5864));
  jand g05801(.dina(n5864), .dinb(n5765), .dout(n5865));
  jxor g05802(.dina(n5752), .dinb(n5744), .dout(n5866));
  jnot g05803(.din(n5866), .dout(n5867));
  jor  g05804(.dina(n5867), .dinb(n5865), .dout(n5868));
  jand g05805(.dina(n5868), .dinb(n5754), .dout(n5869));
  jxor g05806(.dina(n5742), .dinb(n5734), .dout(n5870));
  jnot g05807(.din(n5870), .dout(n5871));
  jor  g05808(.dina(n5871), .dinb(n5869), .dout(n5872));
  jand g05809(.dina(n5872), .dinb(n5743), .dout(n5873));
  jxor g05810(.dina(n5730), .dinb(n5722), .dout(n5874));
  jnot g05811(.din(n5874), .dout(n5875));
  jor  g05812(.dina(n5875), .dinb(n5873), .dout(n5876));
  jand g05813(.dina(n5876), .dinb(n5732), .dout(n5877));
  jxor g05814(.dina(n5719), .dinb(n5711), .dout(n5878));
  jnot g05815(.din(n5878), .dout(n5879));
  jor  g05816(.dina(n5879), .dinb(n5877), .dout(n5880));
  jand g05817(.dina(n5880), .dinb(n5721), .dout(n5881));
  jxor g05818(.dina(n5708), .dinb(n5700), .dout(n5882));
  jnot g05819(.din(n5882), .dout(n5883));
  jor  g05820(.dina(n5883), .dinb(n5881), .dout(n5884));
  jand g05821(.dina(n5884), .dinb(n5710), .dout(n5885));
  jxor g05822(.dina(n5698), .dinb(n5690), .dout(n5886));
  jnot g05823(.din(n5886), .dout(n5887));
  jor  g05824(.dina(n5887), .dinb(n5885), .dout(n5888));
  jand g05825(.dina(n5888), .dinb(n5699), .dout(n5889));
  jxor g05826(.dina(n5687), .dinb(n5679), .dout(n5890));
  jnot g05827(.din(n5890), .dout(n5891));
  jor  g05828(.dina(n5891), .dinb(n5889), .dout(n5892));
  jand g05829(.dina(n5892), .dinb(n5688), .dout(n5893));
  jnot g05830(.din(n5893), .dout(n5894));
  jxor g05831(.dina(n5676), .dinb(n5668), .dout(n5895));
  jand g05832(.dina(n5895), .dinb(n5894), .dout(n5896));
  jor  g05833(.dina(n5896), .dinb(n5678), .dout(n5897));
  jxor g05834(.dina(n5664), .dinb(n5656), .dout(n5898));
  jand g05835(.dina(n5898), .dinb(n5897), .dout(n5899));
  jor  g05836(.dina(n5899), .dinb(n5666), .dout(n5900));
  jxor g05837(.dina(n5653), .dinb(n5645), .dout(n5901));
  jand g05838(.dina(n5901), .dinb(n5900), .dout(n5902));
  jor  g05839(.dina(n5902), .dinb(n5654), .dout(n5903));
  jxor g05840(.dina(n5642), .dinb(n5634), .dout(n5904));
  jand g05841(.dina(n5904), .dinb(n5903), .dout(n5905));
  jor  g05842(.dina(n5905), .dinb(n5644), .dout(n5906));
  jxor g05843(.dina(n5631), .dinb(n5623), .dout(n5907));
  jand g05844(.dina(n5907), .dinb(n5906), .dout(n5908));
  jor  g05845(.dina(n5908), .dinb(n5632), .dout(n5909));
  jxor g05846(.dina(n5621), .dinb(n5613), .dout(n5910));
  jand g05847(.dina(n5910), .dinb(n5909), .dout(n5911));
  jor  g05848(.dina(n5911), .dinb(n5622), .dout(n5912));
  jxor g05849(.dina(n5611), .dinb(n5602), .dout(n5913));
  jnot g05850(.din(n5913), .dout(n5914));
  jand g05851(.dina(n5914), .dinb(n5912), .dout(n5915));
  jor  g05852(.dina(n5915), .dinb(n5612), .dout(n5916));
  jxor g05853(.dina(n5600), .dinb(n5592), .dout(n5917));
  jand g05854(.dina(n5917), .dinb(n5916), .dout(n5918));
  jor  g05855(.dina(n5918), .dinb(n5601), .dout(n5919));
  jxor g05856(.dina(n5589), .dinb(n5581), .dout(n5920));
  jand g05857(.dina(n5920), .dinb(n5919), .dout(n5921));
  jor  g05858(.dina(n5921), .dinb(n5591), .dout(n5922));
  jxor g05859(.dina(n5578), .dinb(n5570), .dout(n5923));
  jand g05860(.dina(n5923), .dinb(n5922), .dout(n5924));
  jor  g05861(.dina(n5924), .dinb(n5579), .dout(n5925));
  jxor g05862(.dina(n5568), .dinb(n5559), .dout(n5926));
  jand g05863(.dina(n5926), .dinb(n5925), .dout(n5927));
  jor  g05864(.dina(n5927), .dinb(n5569), .dout(n5928));
  jnot g05865(.din(n5928), .dout(n5929));
  jxor g05866(.dina(n5557), .dinb(n5547), .dout(n5930));
  jor  g05867(.dina(n5930), .dinb(n5929), .dout(n5931));
  jand g05868(.dina(n5931), .dinb(n5558), .dout(n5932));
  jxor g05869(.dina(n5544), .dinb(n5276), .dout(n5933));
  jnot g05870(.din(n5933), .dout(n5934));
  jor  g05871(.dina(n5934), .dinb(n5932), .dout(n5935));
  jand g05872(.dina(n5935), .dinb(n5546), .dout(n5936));
  jand g05873(.dina(n5274), .dinb(n5162), .dout(n5937));
  jand g05874(.dina(n5275), .dinb(n5052), .dout(n5938));
  jor  g05875(.dina(n5938), .dinb(n5937), .dout(n5939));
  jnot g05876(.din(n5151), .dout(n5940));
  jand g05877(.dina(n5159), .dinb(n5940), .dout(n5941));
  jand g05878(.dina(n5161), .dinb(n5055), .dout(n5942));
  jor  g05879(.dina(n5942), .dinb(n5941), .dout(n5943));
  jnot g05880(.din(n5141), .dout(n5944));
  jor  g05881(.dina(n5149), .dinb(n5944), .dout(n5945));
  jnot g05882(.din(n5945), .dout(n5946));
  jnot g05883(.din(n5150), .dout(n5947));
  jand g05884(.dina(n5947), .dinb(n5058), .dout(n5948));
  jor  g05885(.dina(n5948), .dinb(n5946), .dout(n5949));
  jor  g05886(.dina(n5139), .dinb(n5131), .dout(n5950));
  jnot g05887(.din(n5950), .dout(n5951));
  jand g05888(.dina(n5140), .dinb(n5063), .dout(n5952));
  jor  g05889(.dina(n5952), .dinb(n5951), .dout(n5953));
  jand g05890(.dina(n5128), .dinb(n5120), .dout(n5954));
  jand g05891(.dina(n5129), .dinb(n5066), .dout(n5955));
  jor  g05892(.dina(n5955), .dinb(n5954), .dout(n5956));
  jor  g05893(.dina(n5118), .dinb(n5110), .dout(n5957));
  jand g05894(.dina(n5119), .dinb(n5069), .dout(n5958));
  jnot g05895(.din(n5958), .dout(n5959));
  jand g05896(.dina(n5959), .dinb(n5957), .dout(n5960));
  jnot g05897(.din(n5960), .dout(n5961));
  jor  g05898(.dina(n5107), .dinb(n5099), .dout(n5962));
  jand g05899(.dina(n5108), .dinb(n5072), .dout(n5963));
  jnot g05900(.din(n5963), .dout(n5964));
  jand g05901(.dina(n5964), .dinb(n5962), .dout(n5965));
  jnot g05902(.din(n5965), .dout(n5966));
  jor  g05903(.dina(n5096), .dinb(n5088), .dout(n5967));
  jand g05904(.dina(n5097), .dinb(n5075), .dout(n5968));
  jnot g05905(.din(n5968), .dout(n5969));
  jand g05906(.dina(n5969), .dinb(n5967), .dout(n5970));
  jnot g05907(.din(n5970), .dout(n5971));
  jand g05908(.dina(n480), .dinb(n270), .dout(n5972));
  jand g05909(.dina(n5972), .dinb(n3066), .dout(n5973));
  jand g05910(.dina(n5973), .dinb(n2106), .dout(n5974));
  jand g05911(.dina(n5974), .dinb(n2149), .dout(n5975));
  jand g05912(.dina(n5975), .dinb(n2388), .dout(n5976));
  jand g05913(.dina(n2571), .dinb(n639), .dout(n5977));
  jand g05914(.dina(n5977), .dinb(n838), .dout(n5978));
  jand g05915(.dina(n1470), .dinb(n320), .dout(n5979));
  jand g05916(.dina(n5979), .dinb(n1738), .dout(n5980));
  jand g05917(.dina(n5980), .dinb(n685), .dout(n5981));
  jand g05918(.dina(n5981), .dinb(n5978), .dout(n5982));
  jand g05919(.dina(n510), .dinb(n907), .dout(n5983));
  jand g05920(.dina(n1159), .dinb(n1429), .dout(n5984));
  jand g05921(.dina(n5984), .dinb(n4451), .dout(n5985));
  jand g05922(.dina(n5985), .dinb(n5983), .dout(n5986));
  jand g05923(.dina(n5986), .dinb(n5982), .dout(n5987));
  jand g05924(.dina(n3116), .dinb(n932), .dout(n5988));
  jand g05925(.dina(n1721), .dinb(n1426), .dout(n5989));
  jand g05926(.dina(n886), .dinb(n495), .dout(n5990));
  jand g05927(.dina(n5990), .dinb(n5989), .dout(n5991));
  jand g05928(.dina(n1227), .dinb(n1559), .dout(n5992));
  jand g05929(.dina(n5992), .dinb(n3996), .dout(n5993));
  jand g05930(.dina(n5993), .dinb(n5991), .dout(n5994));
  jand g05931(.dina(n5994), .dinb(n5988), .dout(n5995));
  jand g05932(.dina(n5995), .dinb(n5248), .dout(n5996));
  jand g05933(.dina(n5996), .dinb(n5987), .dout(n5997));
  jand g05934(.dina(n5997), .dinb(n5976), .dout(n5998));
  jand g05935(.dina(n1583), .dinb(n1245), .dout(n5999));
  jand g05936(.dina(n5999), .dinb(n584), .dout(n6000));
  jand g05937(.dina(n6000), .dinb(n1578), .dout(n6001));
  jand g05938(.dina(n881), .dinb(n1334), .dout(n6002));
  jand g05939(.dina(n6002), .dinb(n1228), .dout(n6003));
  jand g05940(.dina(n6003), .dinb(n1366), .dout(n6004));
  jand g05941(.dina(n6004), .dinb(n6001), .dout(n6005));
  jand g05942(.dina(n6005), .dinb(n328), .dout(n6006));
  jand g05943(.dina(n6006), .dinb(n2405), .dout(n6007));
  jand g05944(.dina(n6007), .dinb(n5998), .dout(n6008));
  jand g05945(.dina(n2603), .dinb(n683), .dout(n6009));
  jand g05946(.dina(n1511), .dinb(n588), .dout(n6010));
  jand g05947(.dina(n1212), .dinb(n541), .dout(n6011));
  jand g05948(.dina(n6011), .dinb(n621), .dout(n6012));
  jand g05949(.dina(n6012), .dinb(n1904), .dout(n6013));
  jand g05950(.dina(n6013), .dinb(n6010), .dout(n6014));
  jand g05951(.dina(n3007), .dinb(n101), .dout(n6015));
  jand g05952(.dina(n6015), .dinb(n2570), .dout(n6016));
  jand g05953(.dina(n6016), .dinb(n557), .dout(n6017));
  jand g05954(.dina(n6017), .dinb(n6014), .dout(n6018));
  jand g05955(.dina(n670), .dinb(n351), .dout(n6019));
  jand g05956(.dina(n6019), .dinb(n869), .dout(n6020));
  jand g05957(.dina(n6020), .dinb(n880), .dout(n6021));
  jand g05958(.dina(n844), .dinb(n1261), .dout(n6022));
  jand g05959(.dina(n978), .dinb(n718), .dout(n6023));
  jand g05960(.dina(n6023), .dinb(n951), .dout(n6024));
  jand g05961(.dina(n6024), .dinb(n6022), .dout(n6025));
  jand g05962(.dina(n6025), .dinb(n6021), .dout(n6026));
  jand g05963(.dina(n6026), .dinb(n6018), .dout(n6027));
  jand g05964(.dina(n6027), .dinb(n6009), .dout(n6028));
  jand g05965(.dina(n2100), .dinb(n954), .dout(n6029));
  jand g05966(.dina(n6029), .dinb(n1449), .dout(n6030));
  jand g05967(.dina(n1852), .dinb(n630), .dout(n6031));
  jand g05968(.dina(n6031), .dinb(n465), .dout(n6032));
  jand g05969(.dina(n6032), .dinb(n1188), .dout(n6033));
  jand g05970(.dina(n6033), .dinb(n6030), .dout(n6034));
  jand g05971(.dina(n934), .dinb(n965), .dout(n6035));
  jand g05972(.dina(n6035), .dinb(n1702), .dout(n6036));
  jand g05973(.dina(n2588), .dinb(n1851), .dout(n6037));
  jand g05974(.dina(n6037), .dinb(n4588), .dout(n6038));
  jand g05975(.dina(n6038), .dinb(n6036), .dout(n6039));
  jand g05976(.dina(n1757), .dinb(n1688), .dout(n6040));
  jand g05977(.dina(n6040), .dinb(n547), .dout(n6041));
  jand g05978(.dina(n1732), .dinb(n1462), .dout(n6042));
  jand g05979(.dina(n6042), .dinb(n6041), .dout(n6043));
  jand g05980(.dina(n6043), .dinb(n6039), .dout(n6044));
  jand g05981(.dina(n6044), .dinb(n6034), .dout(n6045));
  jand g05982(.dina(n6045), .dinb(n6028), .dout(n6046));
  jand g05983(.dina(n6046), .dinb(n6008), .dout(n6047));
  jnot g05984(.din(n6047), .dout(n6048));
  jand g05985(.dina(n5076), .dinb(n1639), .dout(n6049));
  jand g05986(.dina(n89), .dinb(\a[31] ), .dout(n6050));
  jand g05987(.dina(n6050), .dinb(n438), .dout(n6051));
  jor  g05988(.dina(n6051), .dinb(n6049), .dout(n6052));
  jand g05989(.dina(n5084), .dinb(n1175), .dout(n6053));
  jand g05990(.dina(n5082), .dinb(n795), .dout(n6054));
  jor  g05991(.dina(n6054), .dinb(n6053), .dout(n6055));
  jor  g05992(.dina(n6055), .dinb(n6052), .dout(n6056));
  jxor g05993(.dina(n6056), .dinb(n6048), .dout(n6057));
  jor  g05994(.dina(n4343), .dinb(n1792), .dout(n6058));
  jor  g05995(.dina(n4348), .dinb(n1790), .dout(n6059));
  jor  g05996(.dina(n3683), .dinb(n1448), .dout(n6060));
  jor  g05997(.dina(n4346), .dinb(n1606), .dout(n6061));
  jand g05998(.dina(n6061), .dinb(n6060), .dout(n6062));
  jand g05999(.dina(n6062), .dinb(n6059), .dout(n6063));
  jand g06000(.dina(n6063), .dinb(n6058), .dout(n6064));
  jxor g06001(.dina(n6064), .dinb(n93), .dout(n6065));
  jxor g06002(.dina(n6065), .dinb(n6057), .dout(n6066));
  jxor g06003(.dina(n6066), .dinb(n5971), .dout(n6067));
  jor  g06004(.dina(n2176), .dinb(n2303), .dout(n6068));
  jor  g06005(.dina(n2174), .dinb(n2309), .dout(n6069));
  jor  g06006(.dina(n2057), .dinb(n1805), .dout(n6070));
  jor  g06007(.dina(n1954), .dinb(n2306), .dout(n6071));
  jand g06008(.dina(n6071), .dinb(n6070), .dout(n6072));
  jand g06009(.dina(n6072), .dinb(n6069), .dout(n6073));
  jand g06010(.dina(n6073), .dinb(n6068), .dout(n6074));
  jxor g06011(.dina(n6074), .dinb(n77), .dout(n6075));
  jxor g06012(.dina(n6075), .dinb(n6067), .dout(n6076));
  jxor g06013(.dina(n6076), .dinb(n5966), .dout(n6077));
  jor  g06014(.dina(n2768), .dinb(n807), .dout(n6078));
  jor  g06015(.dina(n2553), .dinb(n1621), .dout(n6079));
  jor  g06016(.dina(n2428), .dinb(n1617), .dout(n6080));
  jor  g06017(.dina(n2629), .dinb(n1613), .dout(n6081));
  jand g06018(.dina(n6081), .dinb(n6080), .dout(n6082));
  jand g06019(.dina(n6082), .dinb(n6079), .dout(n6083));
  jand g06020(.dina(n6083), .dinb(n6078), .dout(n6084));
  jxor g06021(.dina(n6084), .dinb(n65), .dout(n6085));
  jxor g06022(.dina(n6085), .dinb(n6077), .dout(n6086));
  jxor g06023(.dina(n6086), .dinb(n5961), .dout(n6087));
  jnot g06024(.din(n6087), .dout(n6088));
  jor  g06025(.dina(n3451), .dinb(n1820), .dout(n6089));
  jor  g06026(.dina(n3072), .dinb(n2181), .dout(n6090));
  jor  g06027(.dina(n3203), .dinb(n2189), .dout(n6091));
  jand g06028(.dina(n6091), .dinb(n6090), .dout(n6092));
  jor  g06029(.dina(n2738), .dinb(n2186), .dout(n6093));
  jand g06030(.dina(n6093), .dinb(n6092), .dout(n6094));
  jand g06031(.dina(n6094), .dinb(n6089), .dout(n6095));
  jxor g06032(.dina(n6095), .dinb(\a[20] ), .dout(n6096));
  jxor g06033(.dina(n6096), .dinb(n6088), .dout(n6097));
  jxor g06034(.dina(n6097), .dinb(n5956), .dout(n6098));
  jnot g06035(.din(n6098), .dout(n6099));
  jor  g06036(.dina(n3789), .dinb(n2744), .dout(n6100));
  jor  g06037(.dina(n3420), .dinb(n2749), .dout(n6101));
  jor  g06038(.dina(n3286), .dinb(n2758), .dout(n6102));
  jand g06039(.dina(n6102), .dinb(n6101), .dout(n6103));
  jor  g06040(.dina(n3787), .dinb(n2753), .dout(n6104));
  jand g06041(.dina(n6104), .dinb(n6103), .dout(n6105));
  jand g06042(.dina(n6105), .dinb(n6100), .dout(n6106));
  jxor g06043(.dina(n6106), .dinb(\a[17] ), .dout(n6107));
  jxor g06044(.dina(n6107), .dinb(n6099), .dout(n6108));
  jxor g06045(.dina(n6108), .dinb(n5953), .dout(n6109));
  jor  g06046(.dina(n4021), .dinb(n3424), .dout(n6110));
  jor  g06047(.dina(n3863), .dinb(n3211), .dout(n6111));
  jor  g06048(.dina(n4019), .dinb(n3426), .dout(n6112));
  jor  g06049(.dina(n3929), .dinb(n3429), .dout(n6113));
  jand g06050(.dina(n6113), .dinb(n6112), .dout(n6114));
  jand g06051(.dina(n6114), .dinb(n6111), .dout(n6115));
  jand g06052(.dina(n6115), .dinb(n6110), .dout(n6116));
  jxor g06053(.dina(n6116), .dinb(n3473), .dout(n6117));
  jxor g06054(.dina(n6117), .dinb(n6109), .dout(n6118));
  jxor g06055(.dina(n6118), .dinb(n5949), .dout(n6119));
  jor  g06056(.dina(n4714), .dinb(n4023), .dout(n6120));
  jor  g06057(.dina(n4596), .dinb(n4028), .dout(n6121));
  jor  g06058(.dina(n4471), .dinb(n3871), .dout(n6122));
  jor  g06059(.dina(n4526), .dinb(n4025), .dout(n6123));
  jand g06060(.dina(n6123), .dinb(n6122), .dout(n6124));
  jand g06061(.dina(n6124), .dinb(n6121), .dout(n6125));
  jand g06062(.dina(n6125), .dinb(n6120), .dout(n6126));
  jxor g06063(.dina(n6126), .dinb(n4050), .dout(n6127));
  jxor g06064(.dina(n6127), .dinb(n6119), .dout(n6128));
  jxor g06065(.dina(n6128), .dinb(n5943), .dout(n6129));
  jor  g06066(.dina(n5560), .dinb(n4692), .dout(n6130));
  jor  g06067(.dina(n5264), .dinb(n4697), .dout(n6131));
  jor  g06068(.dina(n4702), .dinb(n4686), .dout(n6132));
  jor  g06069(.dina(n5422), .dinb(n4705), .dout(n6133));
  jand g06070(.dina(n6133), .dinb(n6132), .dout(n6134));
  jand g06071(.dina(n6134), .dinb(n6131), .dout(n6135));
  jand g06072(.dina(n6135), .dinb(n6130), .dout(n6136));
  jxor g06073(.dina(n6136), .dinb(n4713), .dout(n6137));
  jxor g06074(.dina(n6137), .dinb(n6129), .dout(n6138));
  jxor g06075(.dina(n6138), .dinb(n5939), .dout(n6139));
  jnot g06076(.din(n5525), .dout(n6140));
  jand g06077(.dina(n6140), .dinb(n5365), .dout(n6141));
  jnot g06078(.din(n6141), .dout(n6142));
  jnot g06079(.din(n5526), .dout(n6143));
  jor  g06080(.dina(n6143), .dinb(n5441), .dout(n6144));
  jand g06081(.dina(n6144), .dinb(n6142), .dout(n6145));
  jand g06082(.dina(n1227), .dinb(n532), .dout(n6146));
  jand g06083(.dina(n1541), .dinb(n983), .dout(n6147));
  jand g06084(.dina(n6147), .dinb(n662), .dout(n6148));
  jand g06085(.dina(n6148), .dinb(n6146), .dout(n6149));
  jand g06086(.dina(n6149), .dinb(n2603), .dout(n6150));
  jand g06087(.dina(n950), .dinb(n2124), .dout(n6151));
  jand g06088(.dina(n696), .dinb(n1365), .dout(n6152));
  jand g06089(.dina(n6152), .dinb(n6151), .dout(n6153));
  jand g06090(.dina(n6153), .dinb(n6150), .dout(n6154));
  jand g06091(.dina(n3397), .dinb(n2522), .dout(n6155));
  jand g06092(.dina(n349), .dinb(n907), .dout(n6156));
  jand g06093(.dina(n6156), .dinb(n2513), .dout(n6157));
  jand g06094(.dina(n511), .dinb(n1188), .dout(n6158));
  jand g06095(.dina(n6158), .dinb(n6157), .dout(n6159));
  jand g06096(.dina(n6159), .dinb(n6155), .dout(n6160));
  jand g06097(.dina(n6160), .dinb(n6154), .dout(n6161));
  jand g06098(.dina(n1915), .dinb(n557), .dout(n6162));
  jand g06099(.dina(n6162), .dinb(n503), .dout(n6163));
  jand g06100(.dina(n881), .dinb(n871), .dout(n6164));
  jand g06101(.dina(n6164), .dinb(n5354), .dout(n6165));
  jand g06102(.dina(n6165), .dinb(n6163), .dout(n6166));
  jand g06103(.dina(n6166), .dinb(n3124), .dout(n6167));
  jand g06104(.dina(n6167), .dinb(n6161), .dout(n6168));
  jand g06105(.dina(n1772), .dinb(n1099), .dout(n6169));
  jand g06106(.dina(n6169), .dinb(n428), .dout(n6170));
  jand g06107(.dina(n6170), .dinb(n1451), .dout(n6171));
  jnot g06108(.din(n575), .dout(n6172));
  jand g06109(.dina(n630), .dinb(n447), .dout(n6173));
  jand g06110(.dina(n6173), .dinb(n829), .dout(n6174));
  jand g06111(.dina(n6174), .dinb(n6172), .dout(n6175));
  jand g06112(.dina(n6175), .dinb(n1893), .dout(n6176));
  jand g06113(.dina(n6176), .dinb(n6171), .dout(n6177));
  jand g06114(.dina(n1532), .dinb(n1334), .dout(n6178));
  jand g06115(.dina(n1536), .dinb(n1036), .dout(n6179));
  jand g06116(.dina(n6179), .dinb(n6178), .dout(n6180));
  jand g06117(.dina(n6180), .dinb(n1461), .dout(n6181));
  jand g06118(.dina(n6181), .dinb(n2390), .dout(n6182));
  jand g06119(.dina(n6182), .dinb(n6177), .dout(n6183));
  jand g06120(.dina(n1822), .dinb(n1283), .dout(n6184));
  jand g06121(.dina(n6184), .dinb(n676), .dout(n6185));
  jand g06122(.dina(n6185), .dinb(n450), .dout(n6186));
  jand g06123(.dina(n6186), .dinb(n641), .dout(n6187));
  jand g06124(.dina(n6187), .dinb(n6183), .dout(n6188));
  jand g06125(.dina(n6188), .dinb(n6168), .dout(n6189));
  jand g06126(.dina(n4517), .dinb(n1470), .dout(n6190));
  jand g06127(.dina(n6190), .dinb(n1315), .dout(n6191));
  jand g06128(.dina(n547), .dinb(n510), .dout(n6192));
  jand g06129(.dina(n6192), .dinb(n2499), .dout(n6193));
  jand g06130(.dina(n6193), .dinb(n6191), .dout(n6194));
  jand g06131(.dina(n2993), .dinb(n1714), .dout(n6195));
  jand g06132(.dina(n638), .dinb(n1430), .dout(n6196));
  jand g06133(.dina(n6196), .dinb(n514), .dout(n6197));
  jand g06134(.dina(n6197), .dinb(n6195), .dout(n6198));
  jand g06135(.dina(n869), .dinb(n901), .dout(n6199));
  jand g06136(.dina(n6199), .dinb(n1559), .dout(n6200));
  jand g06137(.dina(n6200), .dinb(n1569), .dout(n6201));
  jand g06138(.dina(n6201), .dinb(n6198), .dout(n6202));
  jand g06139(.dina(n6202), .dinb(n6194), .dout(n6203));
  jand g06140(.dina(n6203), .dinb(n2471), .dout(n6204));
  jand g06141(.dina(n6204), .dinb(n6189), .dout(n6205));
  jxor g06142(.dina(n6205), .dinb(n5525), .dout(n6206));
  jxor g06143(.dina(n6206), .dinb(n6145), .dout(n6207));
  jor  g06144(.dina(n6207), .dinb(n5281), .dout(n6208));
  jor  g06145(.dina(n5532), .dinb(n5525), .dout(n6209));
  jor  g06146(.dina(n6205), .dinb(n5539), .dout(n6210));
  jand g06147(.dina(n6210), .dinb(n6209), .dout(n6211));
  jor  g06148(.dina(n5537), .dinb(n5364), .dout(n6212));
  jand g06149(.dina(n6212), .dinb(n6211), .dout(n6213));
  jand g06150(.dina(n6213), .dinb(n6208), .dout(n6214));
  jxor g06151(.dina(n6214), .dinb(\a[5] ), .dout(n6215));
  jxor g06152(.dina(n6215), .dinb(n6139), .dout(n6216));
  jnot g06153(.din(n6216), .dout(n6217));
  jxor g06154(.dina(n6217), .dinb(n5936), .dout(n6218));
  jnot g06155(.din(\a[2] ), .dout(n6219));
  jand g06156(.dina(n440), .dinb(n452), .dout(n6220));
  jand g06157(.dina(n1038), .dinb(n537), .dout(n6221));
  jand g06158(.dina(n3743), .dinb(n1237), .dout(n6222));
  jand g06159(.dina(n6222), .dinb(n6221), .dout(n6223));
  jand g06160(.dina(n6223), .dinb(n6220), .dout(n6224));
  jand g06161(.dina(n6224), .dinb(n1324), .dout(n6225));
  jand g06162(.dina(n641), .dinb(n621), .dout(n6226));
  jand g06163(.dina(n6226), .dinb(n668), .dout(n6227));
  jand g06164(.dina(n653), .dinb(n100), .dout(n6228));
  jand g06165(.dina(n931), .dinb(n447), .dout(n6229));
  jand g06166(.dina(n6229), .dinb(n6228), .dout(n6230));
  jand g06167(.dina(n6230), .dinb(n6227), .dout(n6231));
  jand g06168(.dina(n6231), .dinb(n2149), .dout(n6232));
  jand g06169(.dina(n3782), .dinb(n909), .dout(n6233));
  jand g06170(.dina(n6233), .dinb(n6232), .dout(n6234));
  jand g06171(.dina(n6234), .dinb(n6225), .dout(n6235));
  jand g06172(.dina(n1218), .dinb(n1738), .dout(n6236));
  jand g06173(.dina(n6236), .dinb(n4617), .dout(n6237));
  jand g06174(.dina(n6237), .dinb(n1708), .dout(n6238));
  jand g06175(.dina(n6238), .dinb(n4537), .dout(n6239));
  jand g06176(.dina(n1247), .dinb(n660), .dout(n6240));
  jand g06177(.dina(n1349), .dinb(n1225), .dout(n6241));
  jand g06178(.dina(n516), .dinb(n811), .dout(n6242));
  jand g06179(.dina(n6242), .dinb(n6241), .dout(n6243));
  jand g06180(.dina(n6243), .dinb(n6240), .dout(n6244));
  jand g06181(.dina(n5231), .dinb(n1099), .dout(n6245));
  jand g06182(.dina(n6245), .dinb(n6244), .dout(n6246));
  jand g06183(.dina(n6246), .dinb(n6239), .dout(n6247));
  jand g06184(.dina(n6247), .dinb(n6235), .dout(n6248));
  jand g06185(.dina(n1595), .dinb(n2124), .dout(n6249));
  jand g06186(.dina(n442), .dinb(n1040), .dout(n6250));
  jand g06187(.dina(n6250), .dinb(n4576), .dout(n6251));
  jand g06188(.dina(n6251), .dinb(n1351), .dout(n6252));
  jand g06189(.dina(n6252), .dinb(n6249), .dout(n6253));
  jand g06190(.dina(n4417), .dinb(n1096), .dout(n6254));
  jand g06191(.dina(n6254), .dinb(n3150), .dout(n6255));
  jand g06192(.dina(n1159), .dinb(n1088), .dout(n6256));
  jand g06193(.dina(n6256), .dinb(n3751), .dout(n6257));
  jand g06194(.dina(n6257), .dinb(n6255), .dout(n6258));
  jand g06195(.dina(n6258), .dinb(n2332), .dout(n6259));
  jand g06196(.dina(n983), .dinb(n557), .dout(n6260));
  jand g06197(.dina(n6260), .dinb(n632), .dout(n6261));
  jand g06198(.dina(n6261), .dinb(n809), .dout(n6262));
  jand g06199(.dina(n1212), .dinb(n430), .dout(n6263));
  jand g06200(.dina(n6263), .dinb(n6262), .dout(n6264));
  jand g06201(.dina(n6264), .dinb(n1772), .dout(n6265));
  jand g06202(.dina(n6265), .dinb(n6259), .dout(n6266));
  jand g06203(.dina(n6266), .dinb(n6253), .dout(n6267));
  jand g06204(.dina(n6267), .dinb(n6248), .dout(n6268));
  jand g06205(.dina(n1731), .dinb(n1903), .dout(n6269));
  jand g06206(.dina(n1559), .dinb(n1273), .dout(n6270));
  jand g06207(.dina(n3752), .dinb(n880), .dout(n6271));
  jand g06208(.dina(n6271), .dinb(n6270), .dout(n6272));
  jand g06209(.dina(n895), .dinb(n428), .dout(n6273));
  jand g06210(.dina(n6273), .dinb(n1376), .dout(n6274));
  jand g06211(.dina(n6274), .dinb(n3063), .dout(n6275));
  jand g06212(.dina(n6275), .dinb(n6272), .dout(n6276));
  jand g06213(.dina(n6276), .dinb(n563), .dout(n6277));
  jand g06214(.dina(n6277), .dinb(n6269), .dout(n6278));
  jand g06215(.dina(n873), .dinb(n948), .dout(n6279));
  jand g06216(.dina(n6279), .dinb(n1207), .dout(n6280));
  jand g06217(.dina(n6280), .dinb(n3808), .dout(n6281));
  jand g06218(.dina(n6281), .dinb(n6278), .dout(n6282));
  jand g06219(.dina(n1506), .dinb(n493), .dout(n6283));
  jand g06220(.dina(n6283), .dinb(n699), .dout(n6284));
  jand g06221(.dina(n1743), .dinb(n691), .dout(n6285));
  jand g06222(.dina(n351), .dinb(n121), .dout(n6286));
  jand g06223(.dina(n6286), .dinb(n6285), .dout(n6287));
  jand g06224(.dina(n6287), .dinb(n1957), .dout(n6288));
  jand g06225(.dina(n6288), .dinb(n6284), .dout(n6289));
  jand g06226(.dina(n2500), .dinb(n1735), .dout(n6290));
  jand g06227(.dina(n6290), .dinb(n6289), .dout(n6291));
  jand g06228(.dina(n1451), .dinb(n541), .dout(n6292));
  jand g06229(.dina(n1373), .dinb(n654), .dout(n6293));
  jand g06230(.dina(n6293), .dinb(n6292), .dout(n6294));
  jand g06231(.dina(n6294), .dinb(n6291), .dout(n6295));
  jand g06232(.dina(n6295), .dinb(n6282), .dout(n6296));
  jand g06233(.dina(n6296), .dinb(n6268), .dout(n6297));
  jnot g06234(.din(n6297), .dout(n6298));
  jand g06235(.dina(n3130), .dinb(n1772), .dout(n6299));
  jand g06236(.dina(n6299), .dinb(n981), .dout(n6300));
  jand g06237(.dina(n1225), .dinb(n1270), .dout(n6301));
  jand g06238(.dina(n6301), .dinb(n1334), .dout(n6302));
  jand g06239(.dina(n6302), .dinb(n5979), .dout(n6303));
  jand g06240(.dina(n6303), .dinb(n6300), .dout(n6304));
  jand g06241(.dina(n6304), .dinb(n3751), .dout(n6305));
  jand g06242(.dina(n917), .dinb(n563), .dout(n6306));
  jand g06243(.dina(n6306), .dinb(n2571), .dout(n6307));
  jand g06244(.dina(n6307), .dinb(n1476), .dout(n6308));
  jand g06245(.dina(n1532), .dinb(n901), .dout(n6309));
  jand g06246(.dina(n6309), .dinb(n548), .dout(n6310));
  jand g06247(.dina(n833), .dinb(n411), .dout(n6311));
  jand g06248(.dina(n6311), .dinb(n532), .dout(n6312));
  jand g06249(.dina(n6312), .dinb(n6310), .dout(n6313));
  jand g06250(.dina(n6313), .dinb(n6308), .dout(n6314));
  jand g06251(.dina(n881), .dinb(n929), .dout(n6315));
  jand g06252(.dina(n6315), .dinb(n1592), .dout(n6316));
  jand g06253(.dina(n6316), .dinb(n1346), .dout(n6317));
  jand g06254(.dina(n2029), .dinb(n582), .dout(n6318));
  jand g06255(.dina(n6318), .dinb(n1205), .dout(n6319));
  jand g06256(.dina(n6319), .dinb(n6317), .dout(n6320));
  jand g06257(.dina(n6320), .dinb(n5396), .dout(n6321));
  jand g06258(.dina(n6321), .dinb(n6314), .dout(n6322));
  jand g06259(.dina(n6322), .dinb(n6305), .dout(n6323));
  jand g06260(.dina(n1088), .dinb(n101), .dout(n6324));
  jand g06261(.dina(n6324), .dinb(n6220), .dout(n6325));
  jand g06262(.dina(n1247), .dinb(n704), .dout(n6326));
  jand g06263(.dina(n6326), .dinb(n5518), .dout(n6327));
  jand g06264(.dina(n6327), .dinb(n6325), .dout(n6328));
  jand g06265(.dina(n1037), .dinb(n1310), .dout(n6329));
  jand g06266(.dina(n6329), .dinb(n3752), .dout(n6330));
  jand g06267(.dina(n6330), .dinb(n2570), .dout(n6331));
  jand g06268(.dina(n6331), .dinb(n2343), .dout(n6332));
  jand g06269(.dina(n6332), .dinb(n6328), .dout(n6333));
  jand g06270(.dina(n1915), .dinb(n1324), .dout(n6334));
  jand g06271(.dina(n921), .dinb(n450), .dout(n6335));
  jand g06272(.dina(n1098), .dinb(n442), .dout(n6336));
  jand g06273(.dina(n6336), .dinb(n6335), .dout(n6337));
  jand g06274(.dina(n6337), .dinb(n6334), .dout(n6338));
  jand g06275(.dina(n511), .dinb(n1315), .dout(n6339));
  jand g06276(.dina(n6339), .dinb(n4451), .dout(n6340));
  jand g06277(.dina(n6340), .dinb(n6338), .dout(n6341));
  jand g06278(.dina(n1867), .dinb(n521), .dout(n6342));
  jand g06279(.dina(n1524), .dinb(n954), .dout(n6343));
  jand g06280(.dina(n6343), .dinb(n1233), .dout(n6344));
  jand g06281(.dina(n6344), .dinb(n678), .dout(n6345));
  jand g06282(.dina(n1207), .dinb(n1344), .dout(n6346));
  jand g06283(.dina(n3003), .dinb(n1578), .dout(n6347));
  jand g06284(.dina(n6347), .dinb(n6346), .dout(n6348));
  jand g06285(.dina(n6348), .dinb(n6345), .dout(n6349));
  jand g06286(.dina(n6349), .dinb(n6342), .dout(n6350));
  jand g06287(.dina(n6350), .dinb(n6341), .dout(n6351));
  jand g06288(.dina(n6351), .dinb(n6333), .dout(n6352));
  jand g06289(.dina(n6352), .dinb(n6323), .dout(n6353));
  jand g06290(.dina(n1852), .dinb(n893), .dout(n6354));
  jand g06291(.dina(n6354), .dinb(n1460), .dout(n6355));
  jand g06292(.dina(n1042), .dinb(n638), .dout(n6356));
  jand g06293(.dina(n6356), .dinb(n1188), .dout(n6357));
  jand g06294(.dina(n6357), .dinb(n4641), .dout(n6358));
  jand g06295(.dina(n6358), .dinb(n6355), .dout(n6359));
  jand g06296(.dina(n978), .dinb(n871), .dout(n6360));
  jand g06297(.dina(n6360), .dinb(n1189), .dout(n6361));
  jand g06298(.dina(n4422), .dinb(n895), .dout(n6362));
  jand g06299(.dina(n6362), .dinb(n6361), .dout(n6363));
  jand g06300(.dina(n1053), .dinb(n718), .dout(n6364));
  jand g06301(.dina(n6364), .dinb(n2148), .dout(n6365));
  jand g06302(.dina(n6365), .dinb(n5348), .dout(n6366));
  jand g06303(.dina(n6366), .dinb(n6363), .dout(n6367));
  jand g06304(.dina(n824), .dinb(n1559), .dout(n6368));
  jand g06305(.dina(n6368), .dinb(n586), .dout(n6369));
  jand g06306(.dina(n6369), .dinb(n4574), .dout(n6370));
  jand g06307(.dina(n6370), .dinb(n6367), .dout(n6371));
  jand g06308(.dina(n1304), .dinb(n653), .dout(n6372));
  jand g06309(.dina(n6372), .dinb(n2042), .dout(n6373));
  jand g06310(.dina(n1534), .dinb(n469), .dout(n6374));
  jand g06311(.dina(n818), .dinb(n542), .dout(n6375));
  jand g06312(.dina(n6375), .dinb(n6374), .dout(n6376));
  jand g06313(.dina(n6376), .dinb(n6373), .dout(n6377));
  jand g06314(.dina(n1515), .dinb(n1288), .dout(n6378));
  jand g06315(.dina(n6378), .dinb(n632), .dout(n6379));
  jand g06316(.dina(n6379), .dinb(n1497), .dout(n6380));
  jand g06317(.dina(n6380), .dinb(n6377), .dout(n6381));
  jand g06318(.dina(n5378), .dinb(n934), .dout(n6382));
  jand g06319(.dina(n5283), .dinb(n1380), .dout(n6383));
  jand g06320(.dina(n6383), .dinb(n5248), .dout(n6384));
  jand g06321(.dina(n6384), .dinb(n6382), .dout(n6385));
  jand g06322(.dina(n6385), .dinb(n6292), .dout(n6386));
  jand g06323(.dina(n6386), .dinb(n6381), .dout(n6387));
  jand g06324(.dina(n6387), .dinb(n6371), .dout(n6388));
  jand g06325(.dina(n6388), .dinb(n6359), .dout(n6389));
  jand g06326(.dina(n6389), .dinb(n6353), .dout(n6390));
  jnot g06327(.din(n6390), .dout(n6391));
  jand g06328(.dina(n6391), .dinb(n6298), .dout(n6392));
  jnot g06329(.din(n6392), .dout(n6393));
  jnot g06330(.din(n6205), .dout(n6394));
  jand g06331(.dina(n6391), .dinb(n6394), .dout(n6395));
  jnot g06332(.din(n6395), .dout(n6396));
  jand g06333(.dina(n6394), .dinb(n6140), .dout(n6397));
  jnot g06334(.din(n6397), .dout(n6398));
  jnot g06335(.din(n6206), .dout(n6399));
  jor  g06336(.dina(n6399), .dinb(n6145), .dout(n6400));
  jand g06337(.dina(n6400), .dinb(n6398), .dout(n6401));
  jxor g06338(.dina(n6390), .dinb(n6205), .dout(n6402));
  jnot g06339(.din(n6402), .dout(n6403));
  jor  g06340(.dina(n6403), .dinb(n6401), .dout(n6404));
  jand g06341(.dina(n6404), .dinb(n6396), .dout(n6405));
  jxor g06342(.dina(n6390), .dinb(n6297), .dout(n6406));
  jnot g06343(.din(n6406), .dout(n6407));
  jor  g06344(.dina(n6407), .dinb(n6405), .dout(n6408));
  jand g06345(.dina(n6408), .dinb(n6393), .dout(n6409));
  jand g06346(.dina(n447), .dinb(n811), .dout(n6410));
  jand g06347(.dina(n6410), .dinb(n1378), .dout(n6411));
  jand g06348(.dina(n983), .dinb(n114), .dout(n6412));
  jand g06349(.dina(n6412), .dinb(n1890), .dout(n6413));
  jand g06350(.dina(n6413), .dinb(n1460), .dout(n6414));
  jand g06351(.dina(n6414), .dinb(n6411), .dout(n6415));
  jand g06352(.dina(n683), .dinb(n1432), .dout(n6416));
  jand g06353(.dina(n6416), .dinb(n1040), .dout(n6417));
  jand g06354(.dina(n6417), .dinb(n5232), .dout(n6418));
  jand g06355(.dina(n6418), .dinb(n3170), .dout(n6419));
  jand g06356(.dina(n6419), .dinb(n6415), .dout(n6420));
  jand g06357(.dina(n881), .dinb(n492), .dout(n6421));
  jand g06358(.dina(n6421), .dinb(n1430), .dout(n6422));
  jand g06359(.dina(n1515), .dinb(n547), .dout(n6423));
  jand g06360(.dina(n1453), .dinb(n1270), .dout(n6424));
  jand g06361(.dina(n6424), .dinb(n6423), .dout(n6425));
  jand g06362(.dina(n6425), .dinb(n6422), .dout(n6426));
  jand g06363(.dina(n6426), .dinb(n834), .dout(n6427));
  jand g06364(.dina(n6427), .dinb(n1344), .dout(n6428));
  jand g06365(.dina(n6428), .dinb(n5187), .dout(n6429));
  jand g06366(.dina(n701), .dinb(n514), .dout(n6430));
  jand g06367(.dina(n6430), .dinb(n1846), .dout(n6431));
  jand g06368(.dina(n493), .dinb(n121), .dout(n6432));
  jand g06369(.dina(n1697), .dinb(n1310), .dout(n6433));
  jand g06370(.dina(n6433), .dinb(n6432), .dout(n6434));
  jand g06371(.dina(n1713), .dinb(n826), .dout(n6435));
  jand g06372(.dina(n6435), .dinb(n1756), .dout(n6436));
  jand g06373(.dina(n6436), .dinb(n6434), .dout(n6437));
  jand g06374(.dina(n6437), .dinb(n6431), .dout(n6438));
  jand g06375(.dina(n714), .dinb(n82), .dout(n6439));
  jand g06376(.dina(n6439), .dinb(n3007), .dout(n6440));
  jnot g06377(.din(n524), .dout(n6441));
  jand g06378(.dina(n6441), .dinb(n470), .dout(n6442));
  jand g06379(.dina(n430), .dinb(n1188), .dout(n6443));
  jand g06380(.dina(n6443), .dinb(n3397), .dout(n6444));
  jand g06381(.dina(n6444), .dinb(n6442), .dout(n6445));
  jand g06382(.dina(n6445), .dinb(n6440), .dout(n6446));
  jand g06383(.dina(n6446), .dinb(n6438), .dout(n6447));
  jand g06384(.dina(n586), .dinb(n1205), .dout(n6448));
  jand g06385(.dina(n4422), .dinb(n809), .dout(n6449));
  jand g06386(.dina(n6449), .dinb(n1345), .dout(n6450));
  jand g06387(.dina(n6450), .dinb(n6448), .dout(n6451));
  jand g06388(.dina(n6451), .dinb(n6447), .dout(n6452));
  jand g06389(.dina(n6452), .dinb(n6429), .dout(n6453));
  jand g06390(.dina(n6453), .dinb(n6420), .dout(n6454));
  jand g06391(.dina(n3819), .dinb(n1327), .dout(n6455));
  jand g06392(.dina(n6455), .dinb(n6227), .dout(n6456));
  jand g06393(.dina(n6456), .dinb(n6343), .dout(n6457));
  jand g06394(.dina(n1096), .dinb(n1822), .dout(n6458));
  jand g06395(.dina(n1351), .dinb(n1225), .dout(n6459));
  jand g06396(.dina(n6459), .dinb(n2097), .dout(n6460));
  jand g06397(.dina(n6460), .dinb(n6458), .dout(n6461));
  jand g06398(.dina(n6461), .dinb(n6457), .dout(n6462));
  jand g06399(.dina(n270), .dinb(n1261), .dout(n6463));
  jand g06400(.dina(n6463), .dinb(n664), .dout(n6464));
  jand g06401(.dina(n558), .dinb(n175), .dout(n6465));
  jand g06402(.dina(n6465), .dinb(n1309), .dout(n6466));
  jand g06403(.dina(n6466), .dinb(n6464), .dout(n6467));
  jand g06404(.dina(n1189), .dinb(n662), .dout(n6468));
  jand g06405(.dina(n6468), .dinb(n1853), .dout(n6469));
  jand g06406(.dina(n6469), .dinb(n653), .dout(n6470));
  jand g06407(.dina(n6470), .dinb(n6467), .dout(n6471));
  jand g06408(.dina(n2580), .dinb(n1511), .dout(n6472));
  jand g06409(.dina(n6472), .dinb(n411), .dout(n6473));
  jand g06410(.dina(n1107), .dinb(n884), .dout(n6474));
  jand g06411(.dina(n6474), .dinb(n1036), .dout(n6475));
  jand g06412(.dina(n6475), .dinb(n1426), .dout(n6476));
  jand g06413(.dina(n6476), .dinb(n6473), .dout(n6477));
  jand g06414(.dina(n965), .dinb(n1317), .dout(n6478));
  jand g06415(.dina(n6478), .dinb(n136), .dout(n6479));
  jand g06416(.dina(n1247), .dinb(n697), .dout(n6480));
  jand g06417(.dina(n6480), .dinb(n1536), .dout(n6481));
  jand g06418(.dina(n6481), .dinb(n6479), .dout(n6482));
  jand g06419(.dina(n870), .dinb(n501), .dout(n6483));
  jand g06420(.dina(n6483), .dinb(n1291), .dout(n6484));
  jand g06421(.dina(n6484), .dinb(n6482), .dout(n6485));
  jand g06422(.dina(n6485), .dinb(n6477), .dout(n6486));
  jand g06423(.dina(n6486), .dinb(n6471), .dout(n6487));
  jand g06424(.dina(n6487), .dinb(n6462), .dout(n6488));
  jand g06425(.dina(n6488), .dinb(n6454), .dout(n6489));
  jxor g06426(.dina(n6489), .dinb(n6297), .dout(n6490));
  jxor g06427(.dina(n6490), .dinb(n6409), .dout(n6491));
  jnot g06428(.din(\a[1] ), .dout(n6492));
  jxor g06429(.dina(\a[2] ), .dinb(n6492), .dout(n6493));
  jnot g06430(.din(n6493), .dout(n6494));
  jand g06431(.dina(n6494), .dinb(\a[0] ), .dout(n6495));
  jnot g06432(.din(n6495), .dout(n6496));
  jor  g06433(.dina(n6496), .dinb(n6491), .dout(n6497));
  jnot g06434(.din(\a[0] ), .dout(n6498));
  jand g06435(.dina(n6492), .dinb(n6498), .dout(n6499));
  jand g06436(.dina(n6499), .dinb(\a[2] ), .dout(n6500));
  jnot g06437(.din(n6500), .dout(n6501));
  jor  g06438(.dina(n6501), .dinb(n6390), .dout(n6502));
  jand g06439(.dina(n6493), .dinb(\a[0] ), .dout(n6503));
  jnot g06440(.din(n6503), .dout(n6504));
  jor  g06441(.dina(n6504), .dinb(n6489), .dout(n6505));
  jand g06442(.dina(\a[1] ), .dinb(n6498), .dout(n6506));
  jnot g06443(.din(n6506), .dout(n6507));
  jor  g06444(.dina(n6507), .dinb(n6297), .dout(n6508));
  jand g06445(.dina(n6508), .dinb(n6505), .dout(n6509));
  jand g06446(.dina(n6509), .dinb(n6502), .dout(n6510));
  jand g06447(.dina(n6510), .dinb(n6497), .dout(n6511));
  jxor g06448(.dina(n6511), .dinb(n6219), .dout(n6512));
  jxor g06449(.dina(n6512), .dinb(n6218), .dout(n6513));
  jxor g06450(.dina(n5930), .dinb(n5928), .dout(n6514));
  jnot g06451(.din(n6514), .dout(n6515));
  jxor g06452(.dina(n6402), .dinb(n6401), .dout(n6516));
  jor  g06453(.dina(n6516), .dinb(n6496), .dout(n6517));
  jor  g06454(.dina(n6507), .dinb(n6205), .dout(n6518));
  jor  g06455(.dina(n6504), .dinb(n6390), .dout(n6519));
  jand g06456(.dina(n6519), .dinb(n6518), .dout(n6520));
  jor  g06457(.dina(n6501), .dinb(n5525), .dout(n6521));
  jand g06458(.dina(n6521), .dinb(n6520), .dout(n6522));
  jand g06459(.dina(n6522), .dinb(n6517), .dout(n6523));
  jxor g06460(.dina(n6523), .dinb(n6219), .dout(n6524));
  jand g06461(.dina(n6524), .dinb(n6515), .dout(n6525));
  jnot g06462(.din(n6525), .dout(n6526));
  jxor g06463(.dina(n6523), .dinb(\a[2] ), .dout(n6527));
  jand g06464(.dina(n6527), .dinb(n6514), .dout(n6528));
  jxor g06465(.dina(n5926), .dinb(n5925), .dout(n6529));
  jor  g06466(.dina(n6496), .dinb(n6207), .dout(n6530));
  jor  g06467(.dina(n6507), .dinb(n5525), .dout(n6531));
  jor  g06468(.dina(n6504), .dinb(n6205), .dout(n6532));
  jand g06469(.dina(n6532), .dinb(n6531), .dout(n6533));
  jor  g06470(.dina(n6501), .dinb(n5364), .dout(n6534));
  jand g06471(.dina(n6534), .dinb(n6533), .dout(n6535));
  jand g06472(.dina(n6535), .dinb(n6530), .dout(n6536));
  jxor g06473(.dina(n6536), .dinb(n6219), .dout(n6537));
  jand g06474(.dina(n6537), .dinb(n6529), .dout(n6538));
  jnot g06475(.din(n6538), .dout(n6539));
  jnot g06476(.din(n6529), .dout(n6540));
  jxor g06477(.dina(n6536), .dinb(\a[2] ), .dout(n6541));
  jand g06478(.dina(n6541), .dinb(n6540), .dout(n6542));
  jxor g06479(.dina(n5923), .dinb(n5922), .dout(n6543));
  jor  g06480(.dina(n6496), .dinb(n5527), .dout(n6544));
  jor  g06481(.dina(n6507), .dinb(n5364), .dout(n6545));
  jor  g06482(.dina(n6504), .dinb(n5525), .dout(n6546));
  jand g06483(.dina(n6546), .dinb(n6545), .dout(n6547));
  jor  g06484(.dina(n6501), .dinb(n5422), .dout(n6548));
  jand g06485(.dina(n6548), .dinb(n6547), .dout(n6549));
  jand g06486(.dina(n6549), .dinb(n6544), .dout(n6550));
  jxor g06487(.dina(n6550), .dinb(n6219), .dout(n6551));
  jand g06488(.dina(n6551), .dinb(n6543), .dout(n6552));
  jnot g06489(.din(n6552), .dout(n6553));
  jnot g06490(.din(n6543), .dout(n6554));
  jxor g06491(.dina(n6550), .dinb(\a[2] ), .dout(n6555));
  jand g06492(.dina(n6555), .dinb(n6554), .dout(n6556));
  jxor g06493(.dina(n5920), .dinb(n5919), .dout(n6557));
  jor  g06494(.dina(n6496), .dinb(n5549), .dout(n6558));
  jor  g06495(.dina(n6507), .dinb(n5422), .dout(n6559));
  jor  g06496(.dina(n6504), .dinb(n5364), .dout(n6560));
  jand g06497(.dina(n6560), .dinb(n6559), .dout(n6561));
  jor  g06498(.dina(n6501), .dinb(n5264), .dout(n6562));
  jand g06499(.dina(n6562), .dinb(n6561), .dout(n6563));
  jand g06500(.dina(n6563), .dinb(n6558), .dout(n6564));
  jxor g06501(.dina(n6564), .dinb(n6219), .dout(n6565));
  jand g06502(.dina(n6565), .dinb(n6557), .dout(n6566));
  jnot g06503(.din(n6566), .dout(n6567));
  jnot g06504(.din(n6557), .dout(n6568));
  jxor g06505(.dina(n6564), .dinb(\a[2] ), .dout(n6569));
  jand g06506(.dina(n6569), .dinb(n6568), .dout(n6570));
  jxor g06507(.dina(n5917), .dinb(n5916), .dout(n6571));
  jor  g06508(.dina(n6496), .dinb(n5560), .dout(n6572));
  jor  g06509(.dina(n6507), .dinb(n5264), .dout(n6573));
  jor  g06510(.dina(n6504), .dinb(n5422), .dout(n6574));
  jand g06511(.dina(n6574), .dinb(n6573), .dout(n6575));
  jor  g06512(.dina(n6501), .dinb(n4686), .dout(n6576));
  jand g06513(.dina(n6576), .dinb(n6575), .dout(n6577));
  jand g06514(.dina(n6577), .dinb(n6572), .dout(n6578));
  jxor g06515(.dina(n6578), .dinb(n6219), .dout(n6579));
  jand g06516(.dina(n6579), .dinb(n6571), .dout(n6580));
  jnot g06517(.din(n6580), .dout(n6581));
  jnot g06518(.din(n6571), .dout(n6582));
  jxor g06519(.dina(n6578), .dinb(\a[2] ), .dout(n6583));
  jand g06520(.dina(n6583), .dinb(n6582), .dout(n6584));
  jxor g06521(.dina(n5914), .dinb(n5912), .dout(n6585));
  jor  g06522(.dina(n6496), .dinb(n5266), .dout(n6586));
  jor  g06523(.dina(n6507), .dinb(n4686), .dout(n6587));
  jor  g06524(.dina(n6504), .dinb(n5264), .dout(n6588));
  jand g06525(.dina(n6588), .dinb(n6587), .dout(n6589));
  jor  g06526(.dina(n6501), .dinb(n4526), .dout(n6590));
  jand g06527(.dina(n6590), .dinb(n6589), .dout(n6591));
  jand g06528(.dina(n6591), .dinb(n6586), .dout(n6592));
  jxor g06529(.dina(n6592), .dinb(n6219), .dout(n6593));
  jand g06530(.dina(n6593), .dinb(n6585), .dout(n6594));
  jnot g06531(.din(n6594), .dout(n6595));
  jnot g06532(.din(n6585), .dout(n6596));
  jxor g06533(.dina(n6592), .dinb(\a[2] ), .dout(n6597));
  jand g06534(.dina(n6597), .dinb(n6596), .dout(n6598));
  jxor g06535(.dina(n5910), .dinb(n5909), .dout(n6599));
  jor  g06536(.dina(n6496), .dinb(n4688), .dout(n6600));
  jor  g06537(.dina(n6507), .dinb(n4526), .dout(n6601));
  jor  g06538(.dina(n6504), .dinb(n4686), .dout(n6602));
  jand g06539(.dina(n6602), .dinb(n6601), .dout(n6603));
  jor  g06540(.dina(n6501), .dinb(n4596), .dout(n6604));
  jand g06541(.dina(n6604), .dinb(n6603), .dout(n6605));
  jand g06542(.dina(n6605), .dinb(n6600), .dout(n6606));
  jxor g06543(.dina(n6606), .dinb(n6219), .dout(n6607));
  jand g06544(.dina(n6607), .dinb(n6599), .dout(n6608));
  jnot g06545(.din(n6608), .dout(n6609));
  jnot g06546(.din(n6599), .dout(n6610));
  jxor g06547(.dina(n6606), .dinb(\a[2] ), .dout(n6611));
  jand g06548(.dina(n6611), .dinb(n6610), .dout(n6612));
  jnot g06549(.din(n5907), .dout(n6613));
  jxor g06550(.dina(n6613), .dinb(n5906), .dout(n6614));
  jor  g06551(.dina(n6496), .dinb(n4714), .dout(n6615));
  jor  g06552(.dina(n6507), .dinb(n4596), .dout(n6616));
  jor  g06553(.dina(n6504), .dinb(n4526), .dout(n6617));
  jand g06554(.dina(n6617), .dinb(n6616), .dout(n6618));
  jor  g06555(.dina(n6501), .dinb(n4471), .dout(n6619));
  jand g06556(.dina(n6619), .dinb(n6618), .dout(n6620));
  jand g06557(.dina(n6620), .dinb(n6615), .dout(n6621));
  jxor g06558(.dina(n6621), .dinb(\a[2] ), .dout(n6622));
  jand g06559(.dina(n6622), .dinb(n6614), .dout(n6623));
  jxor g06560(.dina(n5898), .dinb(n5897), .dout(n6624));
  jnot g06561(.din(n6624), .dout(n6625));
  jxor g06562(.dina(n5895), .dinb(n5894), .dout(n6626));
  jor  g06563(.dina(n6496), .dinb(n4038), .dout(n6627));
  jor  g06564(.dina(n6507), .dinb(n3863), .dout(n6628));
  jor  g06565(.dina(n6504), .dinb(n3929), .dout(n6629));
  jand g06566(.dina(n6629), .dinb(n6628), .dout(n6630));
  jor  g06567(.dina(n6501), .dinb(n3787), .dout(n6631));
  jand g06568(.dina(n6631), .dinb(n6630), .dout(n6632));
  jand g06569(.dina(n6632), .dinb(n6627), .dout(n6633));
  jxor g06570(.dina(n6633), .dinb(n6219), .dout(n6634));
  jand g06571(.dina(n6634), .dinb(n6626), .dout(n6635));
  jnot g06572(.din(n6635), .dout(n6636));
  jnot g06573(.din(n6626), .dout(n6637));
  jxor g06574(.dina(n6633), .dinb(\a[2] ), .dout(n6638));
  jand g06575(.dina(n6638), .dinb(n6637), .dout(n6639));
  jxor g06576(.dina(n5891), .dinb(n5889), .dout(n6640));
  jor  g06577(.dina(n6496), .dinb(n4051), .dout(n6641));
  jor  g06578(.dina(n6501), .dinb(n3420), .dout(n6642));
  jor  g06579(.dina(n6504), .dinb(n3863), .dout(n6643));
  jand g06580(.dina(n6643), .dinb(n6642), .dout(n6644));
  jor  g06581(.dina(n6507), .dinb(n3787), .dout(n6645));
  jand g06582(.dina(n6645), .dinb(n6644), .dout(n6646));
  jand g06583(.dina(n6646), .dinb(n6641), .dout(n6647));
  jxor g06584(.dina(n6647), .dinb(n6219), .dout(n6648));
  jand g06585(.dina(n6648), .dinb(n6640), .dout(n6649));
  jnot g06586(.din(n6649), .dout(n6650));
  jnot g06587(.din(n6640), .dout(n6651));
  jxor g06588(.dina(n6647), .dinb(\a[2] ), .dout(n6652));
  jand g06589(.dina(n6652), .dinb(n6651), .dout(n6653));
  jxor g06590(.dina(n5887), .dinb(n5885), .dout(n6654));
  jor  g06591(.dina(n6496), .dinb(n3789), .dout(n6655));
  jor  g06592(.dina(n6507), .dinb(n3420), .dout(n6656));
  jor  g06593(.dina(n6501), .dinb(n3286), .dout(n6657));
  jand g06594(.dina(n6657), .dinb(n6656), .dout(n6658));
  jor  g06595(.dina(n6504), .dinb(n3787), .dout(n6659));
  jand g06596(.dina(n6659), .dinb(n6658), .dout(n6660));
  jand g06597(.dina(n6660), .dinb(n6655), .dout(n6661));
  jxor g06598(.dina(n6661), .dinb(n6219), .dout(n6662));
  jand g06599(.dina(n6662), .dinb(n6654), .dout(n6663));
  jnot g06600(.din(n6663), .dout(n6664));
  jnot g06601(.din(n6654), .dout(n6665));
  jxor g06602(.dina(n6661), .dinb(\a[2] ), .dout(n6666));
  jand g06603(.dina(n6666), .dinb(n6665), .dout(n6667));
  jxor g06604(.dina(n5883), .dinb(n5881), .dout(n6668));
  jnot g06605(.din(n6668), .dout(n6669));
  jor  g06606(.dina(n6496), .dinb(n3422), .dout(n6670));
  jand g06607(.dina(n6503), .dinb(n3729), .dout(n6671));
  jand g06608(.dina(n6506), .dinb(n3287), .dout(n6672));
  jor  g06609(.dina(n6672), .dinb(n6671), .dout(n6673));
  jnot g06610(.din(n6673), .dout(n6674));
  jand g06611(.dina(n6674), .dinb(n6670), .dout(n6675));
  jor  g06612(.dina(n6675), .dinb(\a[2] ), .dout(n6676));
  jxor g06613(.dina(n1255), .dinb(n1448), .dout(n6677));
  jand g06614(.dina(n1655), .dinb(n6677), .dout(n6678));
  jor  g06615(.dina(n6678), .dinb(n1176), .dout(n6679));
  jand g06616(.dina(n1607), .dinb(n6679), .dout(n6680));
  jor  g06617(.dina(n6680), .dinb(n1674), .dout(n6681));
  jand g06618(.dina(n1791), .dinb(n6681), .dout(n6682));
  jor  g06619(.dina(n6682), .dinb(n2064), .dout(n6683));
  jand g06620(.dina(n2069), .dinb(n6683), .dout(n6684));
  jor  g06621(.dina(n6684), .dinb(n2062), .dout(n6685));
  jand g06622(.dina(n2073), .dinb(n6685), .dout(n6686));
  jor  g06623(.dina(n6686), .dinb(n2059), .dout(n6687));
  jand g06624(.dina(n2175), .dinb(n6687), .dout(n6688));
  jor  g06625(.dina(n6688), .dinb(n2326), .dout(n6689));
  jand g06626(.dina(n2429), .dinb(n6689), .dout(n6690));
  jor  g06627(.dina(n6690), .dinb(n2636), .dout(n6691));
  jand g06628(.dina(n2641), .dinb(n6691), .dout(n6692));
  jor  g06629(.dina(n6692), .dinb(n2634), .dout(n6693));
  jand g06630(.dina(n2645), .dinb(n6693), .dout(n6694));
  jor  g06631(.dina(n6694), .dinb(n2631), .dout(n6695));
  jand g06632(.dina(n2739), .dinb(n6695), .dout(n6696));
  jor  g06633(.dina(n6696), .dinb(n3075), .dout(n6697));
  jand g06634(.dina(n3080), .dinb(n6697), .dout(n6698));
  jor  g06635(.dina(n6698), .dinb(n3293), .dout(n6699));
  jand g06636(.dina(n3298), .dinb(n6699), .dout(n6700));
  jor  g06637(.dina(n6700), .dinb(n3291), .dout(n6701));
  jand g06638(.dina(n3302), .dinb(n6701), .dout(n6702));
  jor  g06639(.dina(n6702), .dinb(n3288), .dout(n6703));
  jxor g06640(.dina(n3421), .dinb(n6703), .dout(n6704));
  jand g06641(.dina(n6495), .dinb(n6704), .dout(n6705));
  jor  g06642(.dina(n6673), .dinb(n6705), .dout(n6706));
  jand g06643(.dina(n6500), .dinb(n3213), .dout(n6707));
  jor  g06644(.dina(n6707), .dinb(n6219), .dout(n6708));
  jor  g06645(.dina(n6708), .dinb(n6706), .dout(n6709));
  jand g06646(.dina(n6709), .dinb(n6676), .dout(n6710));
  jor  g06647(.dina(n6710), .dinb(n6669), .dout(n6711));
  jand g06648(.dina(n6710), .dinb(n6669), .dout(n6712));
  jxor g06649(.dina(n5879), .dinb(n5877), .dout(n6713));
  jnot g06650(.din(n6713), .dout(n6714));
  jor  g06651(.dina(n6507), .dinb(n3203), .dout(n6715));
  jor  g06652(.dina(n6496), .dinb(n3440), .dout(n6716));
  jor  g06653(.dina(n6504), .dinb(n3286), .dout(n6717));
  jor  g06654(.dina(n6501), .dinb(n3072), .dout(n6718));
  jand g06655(.dina(n6718), .dinb(n6717), .dout(n6719));
  jand g06656(.dina(n6719), .dinb(n6716), .dout(n6720));
  jand g06657(.dina(n6720), .dinb(n6715), .dout(n6721));
  jxor g06658(.dina(n6721), .dinb(\a[2] ), .dout(n6722));
  jor  g06659(.dina(n6722), .dinb(n6714), .dout(n6723));
  jand g06660(.dina(n6722), .dinb(n6714), .dout(n6724));
  jxor g06661(.dina(n5875), .dinb(n5873), .dout(n6725));
  jnot g06662(.din(n6725), .dout(n6726));
  jor  g06663(.dina(n6496), .dinb(n3451), .dout(n6727));
  jor  g06664(.dina(n6507), .dinb(n3072), .dout(n6728));
  jor  g06665(.dina(n6504), .dinb(n3203), .dout(n6729));
  jand g06666(.dina(n6729), .dinb(n6728), .dout(n6730));
  jor  g06667(.dina(n6501), .dinb(n2738), .dout(n6731));
  jand g06668(.dina(n6731), .dinb(n6730), .dout(n6732));
  jand g06669(.dina(n6732), .dinb(n6727), .dout(n6733));
  jxor g06670(.dina(n6733), .dinb(\a[2] ), .dout(n6734));
  jand g06671(.dina(n6734), .dinb(n6726), .dout(n6735));
  jor  g06672(.dina(n6734), .dinb(n6726), .dout(n6736));
  jxor g06673(.dina(n5871), .dinb(n5869), .dout(n6737));
  jor  g06674(.dina(n6496), .dinb(n3081), .dout(n6738));
  jor  g06675(.dina(n6501), .dinb(n2553), .dout(n6739));
  jor  g06676(.dina(n6507), .dinb(n2738), .dout(n6740));
  jand g06677(.dina(n6740), .dinb(n6739), .dout(n6741));
  jor  g06678(.dina(n6504), .dinb(n3072), .dout(n6742));
  jand g06679(.dina(n6742), .dinb(n6741), .dout(n6743));
  jand g06680(.dina(n6743), .dinb(n6738), .dout(n6744));
  jxor g06681(.dina(n6744), .dinb(n6219), .dout(n6745));
  jand g06682(.dina(n6745), .dinb(n6737), .dout(n6746));
  jnot g06683(.din(n6746), .dout(n6747));
  jnot g06684(.din(n6737), .dout(n6748));
  jxor g06685(.dina(n6744), .dinb(\a[2] ), .dout(n6749));
  jand g06686(.dina(n6749), .dinb(n6748), .dout(n6750));
  jxor g06687(.dina(n5867), .dinb(n5865), .dout(n6751));
  jor  g06688(.dina(n6496), .dinb(n2740), .dout(n6752));
  jor  g06689(.dina(n6507), .dinb(n2553), .dout(n6753));
  jor  g06690(.dina(n6504), .dinb(n2738), .dout(n6754));
  jor  g06691(.dina(n6501), .dinb(n2629), .dout(n6755));
  jand g06692(.dina(n6755), .dinb(n6754), .dout(n6756));
  jand g06693(.dina(n6756), .dinb(n6753), .dout(n6757));
  jand g06694(.dina(n6757), .dinb(n6752), .dout(n6758));
  jxor g06695(.dina(n6758), .dinb(n6219), .dout(n6759));
  jand g06696(.dina(n6759), .dinb(n6751), .dout(n6760));
  jnot g06697(.din(n6760), .dout(n6761));
  jnot g06698(.din(n6751), .dout(n6762));
  jxor g06699(.dina(n6758), .dinb(\a[2] ), .dout(n6763));
  jand g06700(.dina(n6763), .dinb(n6762), .dout(n6764));
  jxor g06701(.dina(n5863), .dinb(n5861), .dout(n6765));
  jor  g06702(.dina(n6496), .dinb(n2768), .dout(n6766));
  jor  g06703(.dina(n6504), .dinb(n2553), .dout(n6767));
  jor  g06704(.dina(n6501), .dinb(n2428), .dout(n6768));
  jand g06705(.dina(n6768), .dinb(n6767), .dout(n6769));
  jor  g06706(.dina(n6507), .dinb(n2629), .dout(n6770));
  jand g06707(.dina(n6770), .dinb(n6769), .dout(n6771));
  jand g06708(.dina(n6771), .dinb(n6766), .dout(n6772));
  jxor g06709(.dina(n6772), .dinb(n6219), .dout(n6773));
  jand g06710(.dina(n6773), .dinb(n6765), .dout(n6774));
  jnot g06711(.din(n6774), .dout(n6775));
  jnot g06712(.din(n6765), .dout(n6776));
  jxor g06713(.dina(n6772), .dinb(\a[2] ), .dout(n6777));
  jand g06714(.dina(n6777), .dinb(n6776), .dout(n6778));
  jxor g06715(.dina(n5859), .dinb(n5857), .dout(n6779));
  jor  g06716(.dina(n6496), .dinb(n2779), .dout(n6780));
  jor  g06717(.dina(n6507), .dinb(n2428), .dout(n6781));
  jor  g06718(.dina(n6504), .dinb(n2629), .dout(n6782));
  jand g06719(.dina(n6782), .dinb(n6781), .dout(n6783));
  jor  g06720(.dina(n6501), .dinb(n2174), .dout(n6784));
  jand g06721(.dina(n6784), .dinb(n6783), .dout(n6785));
  jand g06722(.dina(n6785), .dinb(n6780), .dout(n6786));
  jxor g06723(.dina(n6786), .dinb(n6219), .dout(n6787));
  jand g06724(.dina(n6787), .dinb(n6779), .dout(n6788));
  jnot g06725(.din(n6788), .dout(n6789));
  jnot g06726(.din(n6779), .dout(n6790));
  jxor g06727(.dina(n6786), .dinb(\a[2] ), .dout(n6791));
  jand g06728(.dina(n6791), .dinb(n6790), .dout(n6792));
  jor  g06729(.dina(n6496), .dinb(n2430), .dout(n6793));
  jor  g06730(.dina(n6507), .dinb(n2174), .dout(n6794));
  jor  g06731(.dina(n6504), .dinb(n2428), .dout(n6795));
  jor  g06732(.dina(n6501), .dinb(n1954), .dout(n6796));
  jand g06733(.dina(n6796), .dinb(n6795), .dout(n6797));
  jand g06734(.dina(n6797), .dinb(n6794), .dout(n6798));
  jand g06735(.dina(n6798), .dinb(n6793), .dout(n6799));
  jxor g06736(.dina(n6799), .dinb(n6219), .dout(n6800));
  jxor g06737(.dina(n5855), .dinb(n5853), .dout(n6801));
  jand g06738(.dina(n6801), .dinb(n6800), .dout(n6802));
  jnot g06739(.din(n6802), .dout(n6803));
  jxor g06740(.dina(n6799), .dinb(\a[2] ), .dout(n6804));
  jnot g06741(.din(n6801), .dout(n6805));
  jand g06742(.dina(n6805), .dinb(n6804), .dout(n6806));
  jor  g06743(.dina(n6496), .dinb(n2176), .dout(n6807));
  jor  g06744(.dina(n6504), .dinb(n2174), .dout(n6808));
  jor  g06745(.dina(n6501), .dinb(n2057), .dout(n6809));
  jor  g06746(.dina(n6507), .dinb(n1954), .dout(n6810));
  jand g06747(.dina(n6810), .dinb(n6809), .dout(n6811));
  jand g06748(.dina(n6811), .dinb(n6808), .dout(n6812));
  jand g06749(.dina(n6812), .dinb(n6807), .dout(n6813));
  jxor g06750(.dina(n6813), .dinb(n6219), .dout(n6814));
  jxor g06751(.dina(n5851), .dinb(n5849), .dout(n6815));
  jand g06752(.dina(n6815), .dinb(n6814), .dout(n6816));
  jnot g06753(.din(n6816), .dout(n6817));
  jxor g06754(.dina(n6813), .dinb(\a[2] ), .dout(n6818));
  jnot g06755(.din(n6815), .dout(n6819));
  jand g06756(.dina(n6819), .dinb(n6818), .dout(n6820));
  jxor g06757(.dina(n5847), .dinb(n5845), .dout(n6821));
  jor  g06758(.dina(n6496), .dinb(n2197), .dout(n6822));
  jor  g06759(.dina(n6501), .dinb(n1790), .dout(n6823));
  jor  g06760(.dina(n6504), .dinb(n1954), .dout(n6824));
  jor  g06761(.dina(n6507), .dinb(n2057), .dout(n6825));
  jand g06762(.dina(n6825), .dinb(n6824), .dout(n6826));
  jand g06763(.dina(n6826), .dinb(n6823), .dout(n6827));
  jand g06764(.dina(n6827), .dinb(n6822), .dout(n6828));
  jxor g06765(.dina(n6828), .dinb(n6219), .dout(n6829));
  jand g06766(.dina(n6829), .dinb(n6821), .dout(n6830));
  jnot g06767(.din(n6830), .dout(n6831));
  jnot g06768(.din(n6821), .dout(n6832));
  jxor g06769(.dina(n6828), .dinb(\a[2] ), .dout(n6833));
  jand g06770(.dina(n6833), .dinb(n6832), .dout(n6834));
  jxor g06771(.dina(n5843), .dinb(n5835), .dout(n6835));
  jnot g06772(.din(n6835), .dout(n6836));
  jor  g06773(.dina(n6507), .dinb(n1790), .dout(n6837));
  jor  g06774(.dina(n6496), .dinb(n2208), .dout(n6838));
  jor  g06775(.dina(n6504), .dinb(n2057), .dout(n6839));
  jor  g06776(.dina(n6501), .dinb(n1606), .dout(n6840));
  jand g06777(.dina(n6840), .dinb(n6839), .dout(n6841));
  jand g06778(.dina(n6841), .dinb(n6838), .dout(n6842));
  jand g06779(.dina(n6842), .dinb(n6837), .dout(n6843));
  jxor g06780(.dina(n6843), .dinb(\a[2] ), .dout(n6844));
  jor  g06781(.dina(n6844), .dinb(n6836), .dout(n6845));
  jor  g06782(.dina(n6496), .dinb(n1792), .dout(n6846));
  jor  g06783(.dina(n6504), .dinb(n1790), .dout(n6847));
  jor  g06784(.dina(n6501), .dinb(n1448), .dout(n6848));
  jand g06785(.dina(n6848), .dinb(n6847), .dout(n6849));
  jor  g06786(.dina(n6507), .dinb(n1606), .dout(n6850));
  jand g06787(.dina(n6850), .dinb(n6849), .dout(n6851));
  jand g06788(.dina(n6851), .dinb(n6846), .dout(n6852));
  jxor g06789(.dina(n6852), .dinb(n6219), .dout(n6853));
  jnot g06790(.din(n6853), .dout(n6854));
  jand g06791(.dina(\a[2] ), .dinb(\a[1] ), .dout(n6855));
  jor  g06792(.dina(n6855), .dinb(n6506), .dout(n6856));
  jand g06793(.dina(n6856), .dinb(n795), .dout(n6857));
  jnot g06794(.din(n6857), .dout(n6858));
  jand g06795(.dina(\a[2] ), .dinb(n6492), .dout(n6859));
  jand g06796(.dina(n6859), .dinb(\a[0] ), .dout(n6860));
  jnot g06797(.din(n6860), .dout(n6861));
  jand g06798(.dina(n6861), .dinb(n6504), .dout(n6862));
  jor  g06799(.dina(n6862), .dinb(n1255), .dout(n6863));
  jand g06800(.dina(n6863), .dinb(n6858), .dout(n6864));
  jor  g06801(.dina(n6861), .dinb(n726), .dout(n6865));
  jand g06802(.dina(n6865), .dinb(n1388), .dout(n6866));
  jand g06803(.dina(n6866), .dinb(\a[2] ), .dout(n6867));
  jand g06804(.dina(n6867), .dinb(n6864), .dout(n6868));
  jnot g06805(.din(n6863), .dout(n6871));
  jor  g06806(.dina(n6871), .dinb(n6857), .dout(n6872));
  jand g06807(.dina(n6860), .dinb(n795), .dout(n6873));
  jor  g06808(.dina(n6873), .dinb(n438), .dout(n6874));
  jor  g06809(.dina(n6874), .dinb(n6219), .dout(n6875));
  jor  g06810(.dina(n6875), .dinb(n6872), .dout(n6876));
  jand g06811(.dina(n6876), .dinb(n5820), .dout(n6877));
  jor  g06812(.dina(n6496), .dinb(n1656), .dout(n6878));
  jor  g06813(.dina(n6501), .dinb(n726), .dout(n6879));
  jor  g06814(.dina(n6507), .dinb(n1255), .dout(n6880));
  jand g06815(.dina(n6880), .dinb(n6879), .dout(n6881));
  jor  g06816(.dina(n6504), .dinb(n1448), .dout(n6882));
  jand g06817(.dina(n6882), .dinb(n6881), .dout(n6883));
  jand g06818(.dina(n6883), .dinb(n6878), .dout(n6884));
  jxor g06819(.dina(n6884), .dinb(\a[2] ), .dout(n6885));
  jor  g06820(.dina(n6885), .dinb(n6877), .dout(n6886));
  jand g06821(.dina(n5819), .dinb(\a[5] ), .dout(n6888));
  jxor g06822(.dina(n6888), .dinb(n5818), .dout(n6889));
  jor  g06823(.dina(n6889), .dinb(n6886), .dout(n6890));
  jand g06824(.dina(n6889), .dinb(n6886), .dout(n6891));
  jor  g06825(.dina(n6496), .dinb(n1608), .dout(n6892));
  jor  g06826(.dina(n6501), .dinb(n1255), .dout(n6893));
  jor  g06827(.dina(n6507), .dinb(n1448), .dout(n6894));
  jor  g06828(.dina(n6504), .dinb(n1606), .dout(n6895));
  jand g06829(.dina(n6895), .dinb(n6894), .dout(n6896));
  jand g06830(.dina(n6896), .dinb(n6893), .dout(n6897));
  jand g06831(.dina(n6897), .dinb(n6892), .dout(n6898));
  jxor g06832(.dina(n6898), .dinb(\a[2] ), .dout(n6899));
  jor  g06833(.dina(n6899), .dinb(n6891), .dout(n6900));
  jand g06834(.dina(n6900), .dinb(n6890), .dout(n6901));
  jnot g06835(.din(n5822), .dout(n6902));
  jand g06836(.dina(n6902), .dinb(\a[5] ), .dout(n6903));
  jxor g06837(.dina(n6903), .dinb(n5829), .dout(n6904));
  jnot g06838(.din(n6904), .dout(n6905));
  jor  g06839(.dina(n6905), .dinb(n6901), .dout(n6906));
  jand g06840(.dina(n6906), .dinb(n6854), .dout(n6907));
  jand g06841(.dina(n6905), .dinb(n6901), .dout(n6908));
  jor  g06842(.dina(n6908), .dinb(n6907), .dout(n6909));
  jand g06843(.dina(n6844), .dinb(n6836), .dout(n6910));
  jor  g06844(.dina(n6910), .dinb(n6909), .dout(n6911));
  jand g06845(.dina(n6911), .dinb(n6845), .dout(n6912));
  jor  g06846(.dina(n6912), .dinb(n6834), .dout(n6913));
  jand g06847(.dina(n6913), .dinb(n6831), .dout(n6914));
  jor  g06848(.dina(n6914), .dinb(n6820), .dout(n6915));
  jand g06849(.dina(n6915), .dinb(n6817), .dout(n6916));
  jor  g06850(.dina(n6916), .dinb(n6806), .dout(n6917));
  jand g06851(.dina(n6917), .dinb(n6803), .dout(n6918));
  jor  g06852(.dina(n6918), .dinb(n6792), .dout(n6919));
  jand g06853(.dina(n6919), .dinb(n6789), .dout(n6920));
  jor  g06854(.dina(n6920), .dinb(n6778), .dout(n6921));
  jand g06855(.dina(n6921), .dinb(n6775), .dout(n6922));
  jor  g06856(.dina(n6922), .dinb(n6764), .dout(n6923));
  jand g06857(.dina(n6923), .dinb(n6761), .dout(n6924));
  jor  g06858(.dina(n6924), .dinb(n6750), .dout(n6925));
  jand g06859(.dina(n6925), .dinb(n6747), .dout(n6926));
  jand g06860(.dina(n6926), .dinb(n6736), .dout(n6927));
  jor  g06861(.dina(n6927), .dinb(n6735), .dout(n6928));
  jor  g06862(.dina(n6928), .dinb(n6724), .dout(n6929));
  jand g06863(.dina(n6929), .dinb(n6723), .dout(n6930));
  jor  g06864(.dina(n6930), .dinb(n6712), .dout(n6931));
  jand g06865(.dina(n6931), .dinb(n6711), .dout(n6932));
  jor  g06866(.dina(n6932), .dinb(n6667), .dout(n6933));
  jand g06867(.dina(n6933), .dinb(n6664), .dout(n6934));
  jor  g06868(.dina(n6934), .dinb(n6653), .dout(n6935));
  jand g06869(.dina(n6935), .dinb(n6650), .dout(n6936));
  jor  g06870(.dina(n6936), .dinb(n6639), .dout(n6937));
  jand g06871(.dina(n6937), .dinb(n6636), .dout(n6938));
  jand g06872(.dina(n6938), .dinb(n6625), .dout(n6939));
  jor  g06873(.dina(n6938), .dinb(n6625), .dout(n6940));
  jor  g06874(.dina(n6496), .dinb(n4021), .dout(n6941));
  jor  g06875(.dina(n6501), .dinb(n3863), .dout(n6942));
  jor  g06876(.dina(n6504), .dinb(n4019), .dout(n6943));
  jand g06877(.dina(n6943), .dinb(n6942), .dout(n6944));
  jor  g06878(.dina(n6507), .dinb(n3929), .dout(n6945));
  jand g06879(.dina(n6945), .dinb(n6944), .dout(n6946));
  jand g06880(.dina(n6946), .dinb(n6941), .dout(n6947));
  jxor g06881(.dina(n6947), .dinb(\a[2] ), .dout(n6948));
  jand g06882(.dina(n6948), .dinb(n6940), .dout(n6949));
  jor  g06883(.dina(n6949), .dinb(n6939), .dout(n6950));
  jxor g06884(.dina(n5901), .dinb(n5900), .dout(n6951));
  jor  g06885(.dina(n6496), .dinb(n4473), .dout(n6952));
  jor  g06886(.dina(n6507), .dinb(n4019), .dout(n6953));
  jor  g06887(.dina(n6504), .dinb(n4471), .dout(n6954));
  jand g06888(.dina(n6954), .dinb(n6953), .dout(n6955));
  jor  g06889(.dina(n6501), .dinb(n3929), .dout(n6956));
  jand g06890(.dina(n6956), .dinb(n6955), .dout(n6957));
  jand g06891(.dina(n6957), .dinb(n6952), .dout(n6958));
  jxor g06892(.dina(n6958), .dinb(n6219), .dout(n6959));
  jand g06893(.dina(n6959), .dinb(n6951), .dout(n6960));
  jnot g06894(.din(n6960), .dout(n6961));
  jand g06895(.dina(n6961), .dinb(n6950), .dout(n6962));
  jor  g06896(.dina(n6959), .dinb(n6951), .dout(n6963));
  jnot g06897(.din(n6963), .dout(n6964));
  jor  g06898(.dina(n6964), .dinb(n6962), .dout(n6965));
  jxor g06899(.dina(n5904), .dinb(n5903), .dout(n6966));
  jor  g06900(.dina(n6496), .dinb(n4726), .dout(n6967));
  jor  g06901(.dina(n6507), .dinb(n4471), .dout(n6968));
  jor  g06902(.dina(n6504), .dinb(n4596), .dout(n6969));
  jand g06903(.dina(n6969), .dinb(n6968), .dout(n6970));
  jor  g06904(.dina(n6501), .dinb(n4019), .dout(n6971));
  jand g06905(.dina(n6971), .dinb(n6970), .dout(n6972));
  jand g06906(.dina(n6972), .dinb(n6967), .dout(n6973));
  jxor g06907(.dina(n6973), .dinb(n6219), .dout(n6974));
  jor  g06908(.dina(n6974), .dinb(n6966), .dout(n6975));
  jnot g06909(.din(n6975), .dout(n6976));
  jor  g06910(.dina(n6976), .dinb(n6965), .dout(n6977));
  jor  g06911(.dina(n6622), .dinb(n6614), .dout(n6978));
  jand g06912(.dina(n6974), .dinb(n6966), .dout(n6979));
  jnot g06913(.din(n6979), .dout(n6980));
  jand g06914(.dina(n6980), .dinb(n6978), .dout(n6981));
  jand g06915(.dina(n6981), .dinb(n6977), .dout(n6982));
  jor  g06916(.dina(n6982), .dinb(n6623), .dout(n6983));
  jor  g06917(.dina(n6983), .dinb(n6612), .dout(n6984));
  jand g06918(.dina(n6984), .dinb(n6609), .dout(n6985));
  jor  g06919(.dina(n6985), .dinb(n6598), .dout(n6986));
  jand g06920(.dina(n6986), .dinb(n6595), .dout(n6987));
  jor  g06921(.dina(n6987), .dinb(n6584), .dout(n6988));
  jand g06922(.dina(n6988), .dinb(n6581), .dout(n6989));
  jor  g06923(.dina(n6989), .dinb(n6570), .dout(n6990));
  jand g06924(.dina(n6990), .dinb(n6567), .dout(n6991));
  jor  g06925(.dina(n6991), .dinb(n6556), .dout(n6992));
  jand g06926(.dina(n6992), .dinb(n6553), .dout(n6993));
  jor  g06927(.dina(n6993), .dinb(n6542), .dout(n6994));
  jand g06928(.dina(n6994), .dinb(n6539), .dout(n6995));
  jor  g06929(.dina(n6995), .dinb(n6528), .dout(n6996));
  jand g06930(.dina(n6996), .dinb(n6526), .dout(n6997));
  jxor g06931(.dina(n5933), .dinb(n5932), .dout(n6998));
  jxor g06932(.dina(n6406), .dinb(n6405), .dout(n6999));
  jor  g06933(.dina(n6999), .dinb(n6496), .dout(n7000));
  jor  g06934(.dina(n6501), .dinb(n6205), .dout(n7001));
  jor  g06935(.dina(n6504), .dinb(n6297), .dout(n7002));
  jor  g06936(.dina(n6507), .dinb(n6390), .dout(n7003));
  jand g06937(.dina(n7003), .dinb(n7002), .dout(n7004));
  jand g06938(.dina(n7004), .dinb(n7001), .dout(n7005));
  jand g06939(.dina(n7005), .dinb(n7000), .dout(n7006));
  jxor g06940(.dina(n7006), .dinb(\a[2] ), .dout(n7007));
  jand g06941(.dina(n7007), .dinb(n6998), .dout(n7008));
  jor  g06942(.dina(n7008), .dinb(n6997), .dout(n7009));
  jnot g06943(.din(n5558), .dout(n7010));
  jnot g06944(.din(n5930), .dout(n7011));
  jand g06945(.dina(n7011), .dinb(n5928), .dout(n7012));
  jor  g06946(.dina(n7012), .dinb(n7010), .dout(n7013));
  jxor g06947(.dina(n5933), .dinb(n7013), .dout(n7014));
  jxor g06948(.dina(n7006), .dinb(n6219), .dout(n7015));
  jand g06949(.dina(n7015), .dinb(n7014), .dout(n7016));
  jnot g06950(.din(n7016), .dout(n7017));
  jand g06951(.dina(n7017), .dinb(n7009), .dout(n7018));
  jxor g06952(.dina(n7018), .dinb(n6513), .dout(n7019));
  jand g06953(.dina(n7019), .dinb(n67), .dout(n7020));
  jnot g06954(.din(n7019), .dout(n7021));
  jand g06955(.dina(n5933), .dinb(n7013), .dout(n7022));
  jor  g06956(.dina(n7022), .dinb(n5545), .dout(n7023));
  jxor g06957(.dina(n6217), .dinb(n7023), .dout(n7024));
  jand g06958(.dina(n6512), .dinb(n7024), .dout(n7025));
  jnot g06959(.din(n7025), .dout(n7026));
  jor  g06960(.dina(n7018), .dinb(n6513), .dout(n7027));
  jand g06961(.dina(n7027), .dinb(n7026), .dout(n7028));
  jnot g06962(.din(n6139), .dout(n7029));
  jor  g06963(.dina(n6215), .dinb(n7029), .dout(n7030));
  jnot g06964(.din(n7030), .dout(n7031));
  jand g06965(.dina(n6217), .dinb(n7023), .dout(n7032));
  jor  g06966(.dina(n7032), .dinb(n7031), .dout(n7033));
  jand g06967(.dina(n6137), .dinb(n6129), .dout(n7034));
  jand g06968(.dina(n6138), .dinb(n5939), .dout(n7035));
  jor  g06969(.dina(n7035), .dinb(n7034), .dout(n7036));
  jand g06970(.dina(n6127), .dinb(n6119), .dout(n7037));
  jand g06971(.dina(n6128), .dinb(n5943), .dout(n7038));
  jor  g06972(.dina(n7038), .dinb(n7037), .dout(n7039));
  jand g06973(.dina(n6117), .dinb(n6109), .dout(n7040));
  jand g06974(.dina(n6118), .dinb(n5949), .dout(n7041));
  jor  g06975(.dina(n7041), .dinb(n7040), .dout(n7042));
  jor  g06976(.dina(n6107), .dinb(n6099), .dout(n7043));
  jnot g06977(.din(n7043), .dout(n7044));
  jand g06978(.dina(n6108), .dinb(n5953), .dout(n7045));
  jor  g06979(.dina(n7045), .dinb(n7044), .dout(n7046));
  jor  g06980(.dina(n6096), .dinb(n6088), .dout(n7047));
  jand g06981(.dina(n6097), .dinb(n5956), .dout(n7048));
  jnot g06982(.din(n7048), .dout(n7049));
  jand g06983(.dina(n7049), .dinb(n7047), .dout(n7050));
  jnot g06984(.din(n7050), .dout(n7051));
  jand g06985(.dina(n6085), .dinb(n6077), .dout(n7052));
  jand g06986(.dina(n6086), .dinb(n5961), .dout(n7053));
  jor  g06987(.dina(n7053), .dinb(n7052), .dout(n7054));
  jand g06988(.dina(n6075), .dinb(n6067), .dout(n7055));
  jand g06989(.dina(n6076), .dinb(n5966), .dout(n7056));
  jor  g06990(.dina(n7056), .dinb(n7055), .dout(n7057));
  jand g06991(.dina(n6065), .dinb(n6057), .dout(n7058));
  jand g06992(.dina(n6066), .dinb(n5971), .dout(n7059));
  jor  g06993(.dina(n7059), .dinb(n7058), .dout(n7060));
  jnot g06994(.din(n5076), .dout(n7061));
  jor  g06995(.dina(n7061), .dinb(n1656), .dout(n7062));
  jand g06996(.dina(n6050), .dinb(n795), .dout(n7063));
  jnot g06997(.din(n7063), .dout(n7064));
  jand g06998(.dina(n7064), .dinb(n7062), .dout(n7065));
  jand g06999(.dina(n5082), .dinb(n1175), .dout(n7066));
  jand g07000(.dina(n5084), .dinb(n1024), .dout(n7067));
  jor  g07001(.dina(n7067), .dinb(n7066), .dout(n7068));
  jnot g07002(.din(n7068), .dout(n7069));
  jand g07003(.dina(n7069), .dinb(n7065), .dout(n7070));
  jnot g07004(.din(n7070), .dout(n7071));
  jand g07005(.dina(n6056), .dinb(n6048), .dout(n7072));
  jnot g07006(.din(n7072), .dout(n7073));
  jand g07007(.dina(n466), .dinb(n411), .dout(n7074));
  jand g07008(.dina(n6439), .dinb(n5518), .dout(n7075));
  jand g07009(.dina(n7075), .dinb(n7074), .dout(n7076));
  jand g07010(.dina(n921), .dinb(n6441), .dout(n7077));
  jand g07011(.dina(n7077), .dinb(n3237), .dout(n7078));
  jand g07012(.dina(n7078), .dinb(n7076), .dout(n7079));
  jand g07013(.dina(n7079), .dinb(n535), .dout(n7080));
  jand g07014(.dina(n650), .dinb(n495), .dout(n7081));
  jand g07015(.dina(n1107), .dinb(n916), .dout(n7082));
  jand g07016(.dina(n7082), .dinb(n7081), .dout(n7083));
  jand g07017(.dina(n6184), .dinb(n325), .dout(n7084));
  jand g07018(.dina(n7084), .dinb(n428), .dout(n7085));
  jand g07019(.dina(n833), .dinb(n132), .dout(n7086));
  jand g07020(.dina(n7086), .dinb(n1783), .dout(n7087));
  jand g07021(.dina(n1373), .dinb(n653), .dout(n7088));
  jand g07022(.dina(n1743), .dinb(n510), .dout(n7089));
  jand g07023(.dina(n7089), .dinb(n7088), .dout(n7090));
  jand g07024(.dina(n7090), .dinb(n7087), .dout(n7091));
  jand g07025(.dina(n7091), .dinb(n7085), .dout(n7092));
  jand g07026(.dina(n7092), .dinb(n7083), .dout(n7093));
  jand g07027(.dina(n3178), .dinb(n966), .dout(n7094));
  jand g07028(.dina(n7094), .dinb(n1512), .dout(n7095));
  jand g07029(.dina(n2393), .dinb(n537), .dout(n7096));
  jand g07030(.dina(n7096), .dinb(n7095), .dout(n7097));
  jand g07031(.dina(n7097), .dinb(n7093), .dout(n7098));
  jand g07032(.dina(n7098), .dinb(n7080), .dout(n7099));
  jand g07033(.dina(n7099), .dinb(n685), .dout(n7100));
  jand g07034(.dina(n3920), .dinb(n1243), .dout(n7101));
  jand g07035(.dina(n1561), .dinb(n873), .dout(n7102));
  jand g07036(.dina(n7102), .dinb(n950), .dout(n7103));
  jand g07037(.dina(n469), .dinb(n108), .dout(n7104));
  jand g07038(.dina(n7104), .dinb(n1036), .dout(n7105));
  jand g07039(.dina(n7105), .dinb(n3242), .dout(n7106));
  jand g07040(.dina(n7106), .dinb(n1476), .dout(n7107));
  jand g07041(.dina(n7107), .dinb(n7103), .dout(n7108));
  jand g07042(.dina(n7108), .dinb(n7101), .dout(n7109));
  jand g07043(.dina(n2373), .dinb(n1578), .dout(n7110));
  jand g07044(.dina(n1327), .dinb(n1270), .dout(n7111));
  jand g07045(.dina(n7111), .dinb(n454), .dout(n7112));
  jand g07046(.dina(n7112), .dinb(n7110), .dout(n7113));
  jand g07047(.dina(n1375), .dinb(n481), .dout(n7114));
  jand g07048(.dina(n7114), .dinb(n1698), .dout(n7115));
  jand g07049(.dina(n7115), .dinb(n1366), .dout(n7116));
  jand g07050(.dina(n7116), .dinb(n7113), .dout(n7117));
  jand g07051(.dina(n7117), .dinb(n480), .dout(n7118));
  jand g07052(.dina(n7118), .dinb(n2114), .dout(n7119));
  jand g07053(.dina(n7119), .dinb(n7109), .dout(n7120));
  jand g07054(.dina(n7120), .dinb(n7100), .dout(n7121));
  jxor g07055(.dina(n7121), .dinb(n7073), .dout(n7122));
  jxor g07056(.dina(n7122), .dinb(n7071), .dout(n7123));
  jor  g07057(.dina(n4343), .dinb(n2208), .dout(n7124));
  jor  g07058(.dina(n4346), .dinb(n1790), .dout(n7125));
  jor  g07059(.dina(n3683), .dinb(n1606), .dout(n7126));
  jor  g07060(.dina(n4348), .dinb(n2057), .dout(n7127));
  jand g07061(.dina(n7127), .dinb(n7126), .dout(n7128));
  jand g07062(.dina(n7128), .dinb(n7125), .dout(n7129));
  jand g07063(.dina(n7129), .dinb(n7124), .dout(n7130));
  jxor g07064(.dina(n7130), .dinb(n93), .dout(n7131));
  jxor g07065(.dina(n7131), .dinb(n7123), .dout(n7132));
  jxor g07066(.dina(n7132), .dinb(n7060), .dout(n7133));
  jor  g07067(.dina(n2430), .dinb(n2303), .dout(n7134));
  jor  g07068(.dina(n2174), .dinb(n2306), .dout(n7135));
  jor  g07069(.dina(n2428), .dinb(n2309), .dout(n7136));
  jor  g07070(.dina(n1954), .dinb(n1805), .dout(n7137));
  jand g07071(.dina(n7137), .dinb(n7136), .dout(n7138));
  jand g07072(.dina(n7138), .dinb(n7135), .dout(n7139));
  jand g07073(.dina(n7139), .dinb(n7134), .dout(n7140));
  jxor g07074(.dina(n7140), .dinb(n77), .dout(n7141));
  jxor g07075(.dina(n7141), .dinb(n7133), .dout(n7142));
  jxor g07076(.dina(n7142), .dinb(n7057), .dout(n7143));
  jnot g07077(.din(n7143), .dout(n7144));
  jor  g07078(.dina(n2740), .dinb(n807), .dout(n7145));
  jor  g07079(.dina(n2553), .dinb(n1613), .dout(n7146));
  jor  g07080(.dina(n2629), .dinb(n1617), .dout(n7147));
  jand g07081(.dina(n7147), .dinb(n7146), .dout(n7148));
  jor  g07082(.dina(n2738), .dinb(n1621), .dout(n7149));
  jand g07083(.dina(n7149), .dinb(n7148), .dout(n7150));
  jand g07084(.dina(n7150), .dinb(n7145), .dout(n7151));
  jxor g07085(.dina(n7151), .dinb(\a[23] ), .dout(n7152));
  jxor g07086(.dina(n7152), .dinb(n7144), .dout(n7153));
  jxor g07087(.dina(n7153), .dinb(n7054), .dout(n7154));
  jnot g07088(.din(n7154), .dout(n7155));
  jor  g07089(.dina(n3440), .dinb(n1820), .dout(n7156));
  jor  g07090(.dina(n3203), .dinb(n2181), .dout(n7157));
  jor  g07091(.dina(n3286), .dinb(n2189), .dout(n7158));
  jand g07092(.dina(n7158), .dinb(n7157), .dout(n7159));
  jor  g07093(.dina(n3072), .dinb(n2186), .dout(n7160));
  jand g07094(.dina(n7160), .dinb(n7159), .dout(n7161));
  jand g07095(.dina(n7161), .dinb(n7156), .dout(n7162));
  jxor g07096(.dina(n7162), .dinb(\a[20] ), .dout(n7163));
  jxor g07097(.dina(n7163), .dinb(n7155), .dout(n7164));
  jxor g07098(.dina(n7164), .dinb(n7051), .dout(n7165));
  jor  g07099(.dina(n4051), .dinb(n2744), .dout(n7166));
  jor  g07100(.dina(n3787), .dinb(n2749), .dout(n7167));
  jor  g07101(.dina(n3863), .dinb(n2753), .dout(n7168));
  jor  g07102(.dina(n3420), .dinb(n2758), .dout(n7169));
  jand g07103(.dina(n7169), .dinb(n7168), .dout(n7170));
  jand g07104(.dina(n7170), .dinb(n7167), .dout(n7171));
  jand g07105(.dina(n7171), .dinb(n7166), .dout(n7172));
  jxor g07106(.dina(n7172), .dinb(n2441), .dout(n7173));
  jxor g07107(.dina(n7173), .dinb(n7165), .dout(n7174));
  jxor g07108(.dina(n7174), .dinb(n7046), .dout(n7175));
  jor  g07109(.dina(n4473), .dinb(n3424), .dout(n7176));
  jor  g07110(.dina(n4019), .dinb(n3429), .dout(n7177));
  jor  g07111(.dina(n3929), .dinb(n3211), .dout(n7178));
  jand g07112(.dina(n7178), .dinb(n7177), .dout(n7179));
  jor  g07113(.dina(n4471), .dinb(n3426), .dout(n7180));
  jand g07114(.dina(n7180), .dinb(n7179), .dout(n7181));
  jand g07115(.dina(n7181), .dinb(n7176), .dout(n7182));
  jxor g07116(.dina(n7182), .dinb(\a[14] ), .dout(n7183));
  jxor g07117(.dina(n7183), .dinb(n7175), .dout(n7184));
  jnot g07118(.din(n7184), .dout(n7185));
  jxor g07119(.dina(n7185), .dinb(n7042), .dout(n7186));
  jor  g07120(.dina(n4688), .dinb(n4023), .dout(n7187));
  jor  g07121(.dina(n4526), .dinb(n4028), .dout(n7188));
  jor  g07122(.dina(n4596), .dinb(n3871), .dout(n7189));
  jor  g07123(.dina(n4686), .dinb(n4025), .dout(n7190));
  jand g07124(.dina(n7190), .dinb(n7189), .dout(n7191));
  jand g07125(.dina(n7191), .dinb(n7188), .dout(n7192));
  jand g07126(.dina(n7192), .dinb(n7187), .dout(n7193));
  jxor g07127(.dina(n7193), .dinb(n4050), .dout(n7194));
  jxor g07128(.dina(n7194), .dinb(n7186), .dout(n7195));
  jxor g07129(.dina(n7195), .dinb(n7039), .dout(n7196));
  jnot g07130(.din(n7196), .dout(n7197));
  jor  g07131(.dina(n5549), .dinb(n4692), .dout(n7198));
  jor  g07132(.dina(n5422), .dinb(n4697), .dout(n7199));
  jor  g07133(.dina(n5264), .dinb(n4702), .dout(n7200));
  jand g07134(.dina(n7200), .dinb(n7199), .dout(n7201));
  jor  g07135(.dina(n5364), .dinb(n4705), .dout(n7202));
  jand g07136(.dina(n7202), .dinb(n7201), .dout(n7203));
  jand g07137(.dina(n7203), .dinb(n7198), .dout(n7204));
  jxor g07138(.dina(n7204), .dinb(\a[8] ), .dout(n7205));
  jxor g07139(.dina(n7205), .dinb(n7197), .dout(n7206));
  jxor g07140(.dina(n7206), .dinb(n7036), .dout(n7207));
  jor  g07141(.dina(n6516), .dinb(n5281), .dout(n7208));
  jor  g07142(.dina(n6205), .dinb(n5532), .dout(n7209));
  jor  g07143(.dina(n5537), .dinb(n5525), .dout(n7210));
  jor  g07144(.dina(n6390), .dinb(n5539), .dout(n7211));
  jand g07145(.dina(n7211), .dinb(n7210), .dout(n7212));
  jand g07146(.dina(n7212), .dinb(n7209), .dout(n7213));
  jand g07147(.dina(n7213), .dinb(n7208), .dout(n7214));
  jxor g07148(.dina(n7214), .dinb(n5277), .dout(n7215));
  jxor g07149(.dina(n7215), .dinb(n7207), .dout(n7216));
  jxor g07150(.dina(n7216), .dinb(n7033), .dout(n7217));
  jnot g07151(.din(n6489), .dout(n7218));
  jand g07152(.dina(n7218), .dinb(n6298), .dout(n7219));
  jnot g07153(.din(n7219), .dout(n7220));
  jnot g07154(.din(n6490), .dout(n7221));
  jor  g07155(.dina(n7221), .dinb(n6409), .dout(n7222));
  jand g07156(.dina(n7222), .dinb(n7220), .dout(n7223));
  jand g07157(.dina(n6462), .dinb(n6428), .dout(n7224));
  jand g07158(.dina(n2462), .dinb(n543), .dout(n7225));
  jand g07159(.dina(n1738), .dinb(n132), .dout(n7226));
  jand g07160(.dina(n1451), .dinb(n1583), .dout(n7227));
  jand g07161(.dina(n7227), .dinb(n7226), .dout(n7228));
  jand g07162(.dina(n7228), .dinb(n7225), .dout(n7229));
  jand g07163(.dina(n1834), .dinb(n1713), .dout(n7230));
  jand g07164(.dina(n695), .dinb(n1317), .dout(n7231));
  jand g07165(.dina(n7231), .dinb(n6464), .dout(n7232));
  jand g07166(.dina(n7232), .dinb(n7230), .dout(n7233));
  jand g07167(.dina(n7233), .dinb(n7229), .dout(n7234));
  jand g07168(.dina(n7234), .dinb(n7224), .dout(n7235));
  jand g07169(.dina(n7235), .dinb(n1316), .dout(n7236));
  jand g07170(.dina(n2529), .dinb(n1429), .dout(n7237));
  jand g07171(.dina(n7237), .dinb(n6339), .dout(n7238));
  jand g07172(.dina(n3760), .dinb(n1292), .dout(n7239));
  jand g07173(.dina(n7239), .dinb(n1977), .dout(n7240));
  jand g07174(.dina(n7240), .dinb(n7238), .dout(n7241));
  jand g07175(.dina(n2124), .dinb(n848), .dout(n7242));
  jand g07176(.dina(n1867), .dinb(n1349), .dout(n7243));
  jand g07177(.dina(n7243), .dinb(n7242), .dout(n7244));
  jand g07178(.dina(n1437), .dinb(n676), .dout(n7245));
  jand g07179(.dina(n7245), .dinb(n3814), .dout(n7246));
  jand g07180(.dina(n7246), .dinb(n7244), .dout(n7247));
  jand g07181(.dina(n5285), .dinb(n2500), .dout(n7248));
  jand g07182(.dina(n7248), .dinb(n1593), .dout(n7249));
  jand g07183(.dina(n7249), .dinb(n7247), .dout(n7250));
  jand g07184(.dina(n7250), .dinb(n7241), .dout(n7251));
  jand g07185(.dina(n7251), .dinb(n1365), .dout(n7252));
  jand g07186(.dina(n5351), .dinb(n929), .dout(n7253));
  jand g07187(.dina(n7253), .dinb(n647), .dout(n7254));
  jand g07188(.dina(n2526), .dinb(n982), .dout(n7255));
  jand g07189(.dina(n461), .dinb(n168), .dout(n7256));
  jand g07190(.dina(n7256), .dinb(n681), .dout(n7257));
  jand g07191(.dina(n7257), .dinb(n7255), .dout(n7258));
  jnot g07192(.din(n615), .dout(n7259));
  jand g07193(.dina(n7259), .dinb(n1289), .dout(n7260));
  jand g07194(.dina(n7260), .dinb(n7258), .dout(n7261));
  jand g07195(.dina(n2331), .dinb(n1903), .dout(n7262));
  jand g07196(.dina(n7262), .dinb(n6325), .dout(n7263));
  jand g07197(.dina(n7263), .dinb(n7261), .dout(n7264));
  jand g07198(.dina(n7264), .dinb(n7254), .dout(n7265));
  jand g07199(.dina(n7265), .dinb(n7252), .dout(n7266));
  jand g07200(.dina(n3392), .dinb(n3176), .dout(n7267));
  jand g07201(.dina(n266), .dinb(n1701), .dout(n7268));
  jand g07202(.dina(n1522), .dinb(n463), .dout(n7269));
  jand g07203(.dina(n7269), .dinb(n7268), .dout(n7270));
  jand g07204(.dina(n7270), .dinb(n672), .dout(n7271));
  jand g07205(.dina(n7271), .dinb(n7267), .dout(n7272));
  jand g07206(.dina(n7272), .dinb(n456), .dout(n7273));
  jand g07207(.dina(n7273), .dinb(n7266), .dout(n7274));
  jand g07208(.dina(n7274), .dinb(n7236), .dout(n7275));
  jand g07209(.dina(n715), .dinb(n1203), .dout(n7276));
  jand g07210(.dina(n7276), .dinb(n1169), .dout(n7277));
  jand g07211(.dina(n7277), .dinb(n562), .dout(n7278));
  jand g07212(.dina(n7278), .dinb(n1858), .dout(n7279));
  jand g07213(.dina(n1582), .dinb(n893), .dout(n7280));
  jand g07214(.dina(n4448), .dinb(n1168), .dout(n7281));
  jand g07215(.dina(n7281), .dinb(n7280), .dout(n7282));
  jand g07216(.dina(n7282), .dinb(n1768), .dout(n7283));
  jand g07217(.dina(n7283), .dinb(n6276), .dout(n7284));
  jand g07218(.dina(n7284), .dinb(n7279), .dout(n7285));
  jand g07219(.dina(n1467), .dinb(n1233), .dout(n7286));
  jand g07220(.dina(n1577), .dinb(n445), .dout(n7287));
  jand g07221(.dina(n1476), .dinb(n619), .dout(n7288));
  jand g07222(.dina(n630), .dinb(n499), .dout(n7289));
  jand g07223(.dina(n7289), .dinb(n7288), .dout(n7290));
  jand g07224(.dina(n7290), .dinb(n7287), .dout(n7291));
  jand g07225(.dina(n7291), .dinb(n7286), .dout(n7292));
  jand g07226(.dina(n7292), .dinb(n1016), .dout(n7293));
  jand g07227(.dina(n1310), .dinb(n1432), .dout(n7294));
  jand g07228(.dina(n503), .dinb(n1682), .dout(n7295));
  jand g07229(.dina(n7295), .dinb(n811), .dout(n7296));
  jand g07230(.dina(n7296), .dinb(n7294), .dout(n7297));
  jand g07231(.dina(n7297), .dinb(n6335), .dout(n7298));
  jand g07232(.dina(n7298), .dinb(n7293), .dout(n7299));
  jand g07233(.dina(n7299), .dinb(n7285), .dout(n7300));
  jand g07234(.dina(n7300), .dinb(n7275), .dout(n7301));
  jxor g07235(.dina(n7301), .dinb(n6489), .dout(n7302));
  jxor g07236(.dina(n7302), .dinb(n7223), .dout(n7303));
  jor  g07237(.dina(n7303), .dinb(n6496), .dout(n7304));
  jor  g07238(.dina(n7301), .dinb(n6504), .dout(n7305));
  jor  g07239(.dina(n6501), .dinb(n6297), .dout(n7306));
  jand g07240(.dina(n7306), .dinb(n7305), .dout(n7307));
  jor  g07241(.dina(n6507), .dinb(n6489), .dout(n7308));
  jand g07242(.dina(n7308), .dinb(n7307), .dout(n7309));
  jand g07243(.dina(n7309), .dinb(n7304), .dout(n7310));
  jxor g07244(.dina(n7310), .dinb(\a[2] ), .dout(n7311));
  jxor g07245(.dina(n7311), .dinb(n7217), .dout(n7312));
  jxor g07246(.dina(n7312), .dinb(n7028), .dout(n7313));
  jxor g07247(.dina(n7313), .dinb(n7021), .dout(n7314));
  jnot g07248(.din(n7314), .dout(n7315));
  jand g07249(.dina(n7315), .dinb(n806), .dout(n7316));
  jand g07250(.dina(n7019), .dinb(n1612), .dout(n7317));
  jand g07251(.dina(n7313), .dinb(n1620), .dout(n7318));
  jor  g07252(.dina(n7318), .dinb(n7317), .dout(n7319));
  jor  g07253(.dina(n7319), .dinb(n7316), .dout(n7320));
  jnot g07254(.din(n7320), .dout(n7321));
  jand g07255(.dina(n7019), .dinb(n804), .dout(n7322));
  jnot g07256(.din(n7322), .dout(n7323));
  jand g07257(.dina(n7323), .dinb(\a[23] ), .dout(n7324));
  jand g07258(.dina(n7324), .dinb(n7321), .dout(n7325));
  jand g07259(.dina(n7313), .dinb(n7021), .dout(n7326));
  jor  g07260(.dina(n6216), .dinb(n5936), .dout(n7327));
  jand g07261(.dina(n7327), .dinb(n7030), .dout(n7328));
  jxor g07262(.dina(n7216), .dinb(n7328), .dout(n7329));
  jor  g07263(.dina(n7311), .dinb(n7329), .dout(n7330));
  jnot g07264(.din(n7330), .dout(n7331));
  jxor g07265(.dina(n6512), .dinb(n7024), .dout(n7332));
  jor  g07266(.dina(n6524), .dinb(n6515), .dout(n7333));
  jor  g07267(.dina(n6537), .dinb(n6529), .dout(n7334));
  jor  g07268(.dina(n6551), .dinb(n6543), .dout(n7335));
  jor  g07269(.dina(n6565), .dinb(n6557), .dout(n7336));
  jor  g07270(.dina(n6579), .dinb(n6571), .dout(n7337));
  jor  g07271(.dina(n6593), .dinb(n6585), .dout(n7338));
  jor  g07272(.dina(n6607), .dinb(n6599), .dout(n7339));
  jnot g07273(.din(n6623), .dout(n7340));
  jor  g07274(.dina(n6634), .dinb(n6626), .dout(n7341));
  jor  g07275(.dina(n6648), .dinb(n6640), .dout(n7342));
  jor  g07276(.dina(n6662), .dinb(n6654), .dout(n7343));
  jand g07277(.dina(n6706), .dinb(n6219), .dout(n7344));
  jnot g07278(.din(n6708), .dout(n7345));
  jand g07279(.dina(n7345), .dinb(n6675), .dout(n7346));
  jor  g07280(.dina(n7346), .dinb(n7344), .dout(n7347));
  jand g07281(.dina(n7347), .dinb(n6668), .dout(n7348));
  jor  g07282(.dina(n7347), .dinb(n6668), .dout(n7349));
  jxor g07283(.dina(n6721), .dinb(n6219), .dout(n7350));
  jand g07284(.dina(n7350), .dinb(n6713), .dout(n7351));
  jor  g07285(.dina(n7350), .dinb(n6713), .dout(n7352));
  jnot g07286(.din(n6735), .dout(n7353));
  jxor g07287(.dina(n6733), .dinb(n6219), .dout(n7354));
  jand g07288(.dina(n7354), .dinb(n6725), .dout(n7355));
  jor  g07289(.dina(n6745), .dinb(n6737), .dout(n7356));
  jor  g07290(.dina(n6759), .dinb(n6751), .dout(n7357));
  jor  g07291(.dina(n6773), .dinb(n6765), .dout(n7358));
  jor  g07292(.dina(n6787), .dinb(n6779), .dout(n7359));
  jor  g07293(.dina(n6801), .dinb(n6800), .dout(n7360));
  jor  g07294(.dina(n6815), .dinb(n6814), .dout(n7361));
  jor  g07295(.dina(n6829), .dinb(n6821), .dout(n7362));
  jxor g07296(.dina(n6843), .dinb(n6219), .dout(n7363));
  jand g07297(.dina(n7363), .dinb(n6835), .dout(n7364));
  jor  g07298(.dina(n6868), .dinb(n5819), .dout(n7365));
  jxor g07299(.dina(n6884), .dinb(n6219), .dout(n7366));
  jand g07300(.dina(n7366), .dinb(n7365), .dout(n7367));
  jnot g07301(.din(n6889), .dout(n7369));
  jand g07302(.dina(n7369), .dinb(n7367), .dout(n7370));
  jor  g07303(.dina(n7369), .dinb(n7367), .dout(n7371));
  jxor g07304(.dina(n6898), .dinb(n6219), .dout(n7372));
  jand g07305(.dina(n7372), .dinb(n7371), .dout(n7373));
  jor  g07306(.dina(n7373), .dinb(n7370), .dout(n7374));
  jand g07307(.dina(n6904), .dinb(n7374), .dout(n7375));
  jor  g07308(.dina(n7375), .dinb(n6853), .dout(n7376));
  jor  g07309(.dina(n6904), .dinb(n7374), .dout(n7377));
  jand g07310(.dina(n7377), .dinb(n7376), .dout(n7378));
  jor  g07311(.dina(n7363), .dinb(n6835), .dout(n7379));
  jand g07312(.dina(n7379), .dinb(n7378), .dout(n7380));
  jor  g07313(.dina(n7380), .dinb(n7364), .dout(n7381));
  jand g07314(.dina(n7381), .dinb(n7362), .dout(n7382));
  jor  g07315(.dina(n7382), .dinb(n6830), .dout(n7383));
  jand g07316(.dina(n7383), .dinb(n7361), .dout(n7384));
  jor  g07317(.dina(n7384), .dinb(n6816), .dout(n7385));
  jand g07318(.dina(n7385), .dinb(n7360), .dout(n7386));
  jor  g07319(.dina(n7386), .dinb(n6802), .dout(n7387));
  jand g07320(.dina(n7387), .dinb(n7359), .dout(n7388));
  jor  g07321(.dina(n7388), .dinb(n6788), .dout(n7389));
  jand g07322(.dina(n7389), .dinb(n7358), .dout(n7390));
  jor  g07323(.dina(n7390), .dinb(n6774), .dout(n7391));
  jand g07324(.dina(n7391), .dinb(n7357), .dout(n7392));
  jor  g07325(.dina(n7392), .dinb(n6760), .dout(n7393));
  jand g07326(.dina(n7393), .dinb(n7356), .dout(n7394));
  jor  g07327(.dina(n7394), .dinb(n6746), .dout(n7395));
  jor  g07328(.dina(n7395), .dinb(n7355), .dout(n7396));
  jand g07329(.dina(n7396), .dinb(n7353), .dout(n7397));
  jand g07330(.dina(n7397), .dinb(n7352), .dout(n7398));
  jor  g07331(.dina(n7398), .dinb(n7351), .dout(n7399));
  jand g07332(.dina(n7399), .dinb(n7349), .dout(n7400));
  jor  g07333(.dina(n7400), .dinb(n7348), .dout(n7401));
  jand g07334(.dina(n7401), .dinb(n7343), .dout(n7402));
  jor  g07335(.dina(n7402), .dinb(n6663), .dout(n7403));
  jand g07336(.dina(n7403), .dinb(n7342), .dout(n7404));
  jor  g07337(.dina(n7404), .dinb(n6649), .dout(n7405));
  jand g07338(.dina(n7405), .dinb(n7341), .dout(n7406));
  jor  g07339(.dina(n7406), .dinb(n6635), .dout(n7407));
  jor  g07340(.dina(n7407), .dinb(n6624), .dout(n7408));
  jand g07341(.dina(n7407), .dinb(n6624), .dout(n7409));
  jnot g07342(.din(n6948), .dout(n7410));
  jor  g07343(.dina(n7410), .dinb(n7409), .dout(n7411));
  jand g07344(.dina(n7411), .dinb(n7408), .dout(n7412));
  jor  g07345(.dina(n6960), .dinb(n7412), .dout(n7413));
  jand g07346(.dina(n6963), .dinb(n7413), .dout(n7414));
  jand g07347(.dina(n6975), .dinb(n7414), .dout(n7415));
  jxor g07348(.dina(n5907), .dinb(n5906), .dout(n7416));
  jxor g07349(.dina(n6621), .dinb(n6219), .dout(n7417));
  jand g07350(.dina(n7417), .dinb(n7416), .dout(n7418));
  jor  g07351(.dina(n6979), .dinb(n7418), .dout(n7419));
  jor  g07352(.dina(n7419), .dinb(n7415), .dout(n7420));
  jand g07353(.dina(n7420), .dinb(n7340), .dout(n7421));
  jand g07354(.dina(n7421), .dinb(n7339), .dout(n7422));
  jor  g07355(.dina(n7422), .dinb(n6608), .dout(n7423));
  jand g07356(.dina(n7423), .dinb(n7338), .dout(n7424));
  jor  g07357(.dina(n7424), .dinb(n6594), .dout(n7425));
  jand g07358(.dina(n7425), .dinb(n7337), .dout(n7426));
  jor  g07359(.dina(n7426), .dinb(n6580), .dout(n7427));
  jand g07360(.dina(n7427), .dinb(n7336), .dout(n7428));
  jor  g07361(.dina(n7428), .dinb(n6566), .dout(n7429));
  jand g07362(.dina(n7429), .dinb(n7335), .dout(n7430));
  jor  g07363(.dina(n7430), .dinb(n6552), .dout(n7431));
  jand g07364(.dina(n7431), .dinb(n7334), .dout(n7432));
  jor  g07365(.dina(n7432), .dinb(n6538), .dout(n7433));
  jand g07366(.dina(n7433), .dinb(n7333), .dout(n7434));
  jor  g07367(.dina(n7434), .dinb(n6525), .dout(n7435));
  jor  g07368(.dina(n7015), .dinb(n7014), .dout(n7436));
  jand g07369(.dina(n7436), .dinb(n7435), .dout(n7437));
  jor  g07370(.dina(n7016), .dinb(n7437), .dout(n7438));
  jand g07371(.dina(n7438), .dinb(n7332), .dout(n7439));
  jor  g07372(.dina(n7439), .dinb(n7025), .dout(n7440));
  jxor g07373(.dina(n7311), .dinb(n7329), .dout(n7441));
  jand g07374(.dina(n7441), .dinb(n7440), .dout(n7442));
  jor  g07375(.dina(n7442), .dinb(n7331), .dout(n7443));
  jand g07376(.dina(n7215), .dinb(n7207), .dout(n7444));
  jnot g07377(.din(n7444), .dout(n7445));
  jnot g07378(.din(n7216), .dout(n7446));
  jor  g07379(.dina(n7446), .dinb(n7328), .dout(n7447));
  jand g07380(.dina(n7447), .dinb(n7445), .dout(n7448));
  jor  g07381(.dina(n7205), .dinb(n7197), .dout(n7449));
  jnot g07382(.din(n7449), .dout(n7450));
  jand g07383(.dina(n7206), .dinb(n7036), .dout(n7451));
  jor  g07384(.dina(n7451), .dinb(n7450), .dout(n7452));
  jand g07385(.dina(n7194), .dinb(n7186), .dout(n7453));
  jand g07386(.dina(n7195), .dinb(n7039), .dout(n7454));
  jor  g07387(.dina(n7454), .dinb(n7453), .dout(n7455));
  jnot g07388(.din(n7175), .dout(n7456));
  jor  g07389(.dina(n7183), .dinb(n7456), .dout(n7457));
  jnot g07390(.din(n7457), .dout(n7458));
  jand g07391(.dina(n7185), .dinb(n7042), .dout(n7459));
  jor  g07392(.dina(n7459), .dinb(n7458), .dout(n7460));
  jand g07393(.dina(n7173), .dinb(n7165), .dout(n7461));
  jand g07394(.dina(n7174), .dinb(n7046), .dout(n7462));
  jor  g07395(.dina(n7462), .dinb(n7461), .dout(n7463));
  jor  g07396(.dina(n7163), .dinb(n7155), .dout(n7464));
  jand g07397(.dina(n7164), .dinb(n7051), .dout(n7465));
  jnot g07398(.din(n7465), .dout(n7466));
  jand g07399(.dina(n7466), .dinb(n7464), .dout(n7467));
  jnot g07400(.din(n7467), .dout(n7468));
  jor  g07401(.dina(n7152), .dinb(n7144), .dout(n7469));
  jand g07402(.dina(n7153), .dinb(n7054), .dout(n7470));
  jnot g07403(.din(n7470), .dout(n7471));
  jand g07404(.dina(n7471), .dinb(n7469), .dout(n7472));
  jnot g07405(.din(n7472), .dout(n7473));
  jand g07406(.dina(n7141), .dinb(n7133), .dout(n7474));
  jand g07407(.dina(n7142), .dinb(n7057), .dout(n7475));
  jor  g07408(.dina(n7475), .dinb(n7474), .dout(n7476));
  jand g07409(.dina(n7131), .dinb(n7123), .dout(n7477));
  jand g07410(.dina(n7132), .dinb(n7060), .dout(n7478));
  jor  g07411(.dina(n7478), .dinb(n7477), .dout(n7479));
  jor  g07412(.dina(n7121), .dinb(n7073), .dout(n7480));
  jand g07413(.dina(n7122), .dinb(n7071), .dout(n7481));
  jnot g07414(.din(n7481), .dout(n7482));
  jand g07415(.dina(n7482), .dinb(n7480), .dout(n7483));
  jnot g07416(.din(n7483), .dout(n7484));
  jand g07417(.dina(n3323), .dinb(n503), .dout(n7485));
  jand g07418(.dina(n6343), .dinb(n6158), .dout(n7486));
  jand g07419(.dina(n7486), .dinb(n121), .dout(n7487));
  jand g07420(.dina(n7487), .dinb(n7485), .dout(n7488));
  jand g07421(.dina(n492), .dinb(n560), .dout(n7489));
  jand g07422(.dina(n7489), .dinb(n553), .dout(n7490));
  jand g07423(.dina(n1738), .dinb(n838), .dout(n7491));
  jand g07424(.dina(n7491), .dinb(n3841), .dout(n7492));
  jand g07425(.dina(n7492), .dinb(n843), .dout(n7493));
  jand g07426(.dina(n7493), .dinb(n7490), .dout(n7494));
  jand g07427(.dina(n7494), .dinb(n7488), .dout(n7495));
  jand g07428(.dina(n693), .dinb(n696), .dout(n7496));
  jand g07429(.dina(n7496), .dinb(n7495), .dout(n7497));
  jand g07430(.dina(n1167), .dinb(n991), .dout(n7498));
  jand g07431(.dina(n514), .dinb(n132), .dout(n7499));
  jand g07432(.dina(n7499), .dinb(n1772), .dout(n7500));
  jand g07433(.dina(n7500), .dinb(n1976), .dout(n7501));
  jand g07434(.dina(n7501), .dinb(n7498), .dout(n7502));
  jnot g07435(.din(n961), .dout(n7503));
  jand g07436(.dina(n1169), .dinb(n7503), .dout(n7504));
  jand g07437(.dina(n7504), .dinb(n7502), .dout(n7505));
  jand g07438(.dina(n7505), .dinb(n1852), .dout(n7506));
  jand g07439(.dina(n7506), .dinb(n7497), .dout(n7507));
  jnot g07440(.din(n218), .dout(n7508));
  jand g07441(.dina(n447), .dinb(n108), .dout(n7509));
  jand g07442(.dina(n7509), .dinb(n7508), .dout(n7510));
  jand g07443(.dina(n4422), .dinb(n2149), .dout(n7511));
  jand g07444(.dina(n1437), .dinb(n1708), .dout(n7512));
  jand g07445(.dina(n7512), .dinb(n3136), .dout(n7513));
  jand g07446(.dina(n7513), .dinb(n7511), .dout(n7514));
  jand g07447(.dina(n7514), .dinb(n7510), .dout(n7515));
  jand g07448(.dina(n718), .dinb(n532), .dout(n7516));
  jand g07449(.dina(n641), .dinb(n1213), .dout(n7517));
  jand g07450(.dina(n7517), .dinb(n7516), .dout(n7518));
  jand g07451(.dina(n7518), .dinb(n490), .dout(n7519));
  jand g07452(.dina(n7519), .dinb(n6021), .dout(n7520));
  jand g07453(.dina(n7520), .dinb(n7515), .dout(n7521));
  jand g07454(.dina(n7521), .dinb(n1952), .dout(n7522));
  jand g07455(.dina(n7522), .dinb(n7507), .dout(n7523));
  jor  g07456(.dina(n7061), .dinb(n1608), .dout(n7524));
  jand g07457(.dina(n6050), .dinb(n1175), .dout(n7525));
  jand g07458(.dina(n5082), .dinb(n1024), .dout(n7526));
  jand g07459(.dina(n5084), .dinb(n1673), .dout(n7527));
  jor  g07460(.dina(n7527), .dinb(n7526), .dout(n7528));
  jor  g07461(.dina(n7528), .dinb(n7525), .dout(n7529));
  jnot g07462(.din(n7529), .dout(n7530));
  jand g07463(.dina(n7530), .dinb(n7524), .dout(n7531));
  jxor g07464(.dina(n7531), .dinb(n7523), .dout(n7532));
  jxor g07465(.dina(n7532), .dinb(n7484), .dout(n7533));
  jor  g07466(.dina(n4343), .dinb(n2197), .dout(n7534));
  jor  g07467(.dina(n3683), .dinb(n1790), .dout(n7535));
  jor  g07468(.dina(n4348), .dinb(n1954), .dout(n7536));
  jor  g07469(.dina(n4346), .dinb(n2057), .dout(n7537));
  jand g07470(.dina(n7537), .dinb(n7536), .dout(n7538));
  jand g07471(.dina(n7538), .dinb(n7535), .dout(n7539));
  jand g07472(.dina(n7539), .dinb(n7534), .dout(n7540));
  jxor g07473(.dina(n7540), .dinb(n93), .dout(n7541));
  jxor g07474(.dina(n7541), .dinb(n7533), .dout(n7542));
  jxor g07475(.dina(n7542), .dinb(n7479), .dout(n7543));
  jnot g07476(.din(n7543), .dout(n7544));
  jor  g07477(.dina(n2174), .dinb(n1805), .dout(n7545));
  jor  g07478(.dina(n2779), .dinb(n2303), .dout(n7546));
  jor  g07479(.dina(n2629), .dinb(n2309), .dout(n7547));
  jor  g07480(.dina(n2428), .dinb(n2306), .dout(n7548));
  jand g07481(.dina(n7548), .dinb(n7547), .dout(n7549));
  jand g07482(.dina(n7549), .dinb(n7546), .dout(n7550));
  jand g07483(.dina(n7550), .dinb(n7545), .dout(n7551));
  jxor g07484(.dina(n7551), .dinb(\a[26] ), .dout(n7552));
  jxor g07485(.dina(n7552), .dinb(n7544), .dout(n7553));
  jxor g07486(.dina(n7553), .dinb(n7476), .dout(n7554));
  jnot g07487(.din(n7554), .dout(n7555));
  jor  g07488(.dina(n3081), .dinb(n807), .dout(n7556));
  jor  g07489(.dina(n2553), .dinb(n1617), .dout(n7557));
  jor  g07490(.dina(n2738), .dinb(n1613), .dout(n7558));
  jand g07491(.dina(n7558), .dinb(n7557), .dout(n7559));
  jor  g07492(.dina(n3072), .dinb(n1621), .dout(n7560));
  jand g07493(.dina(n7560), .dinb(n7559), .dout(n7561));
  jand g07494(.dina(n7561), .dinb(n7556), .dout(n7562));
  jxor g07495(.dina(n7562), .dinb(\a[23] ), .dout(n7563));
  jxor g07496(.dina(n7563), .dinb(n7555), .dout(n7564));
  jxor g07497(.dina(n7564), .dinb(n7473), .dout(n7565));
  jnot g07498(.din(n7565), .dout(n7566));
  jor  g07499(.dina(n3203), .dinb(n2186), .dout(n7567));
  jor  g07500(.dina(n3422), .dinb(n1820), .dout(n7568));
  jor  g07501(.dina(n3420), .dinb(n2189), .dout(n7569));
  jor  g07502(.dina(n3286), .dinb(n2181), .dout(n7570));
  jand g07503(.dina(n7570), .dinb(n7569), .dout(n7571));
  jand g07504(.dina(n7571), .dinb(n7568), .dout(n7572));
  jand g07505(.dina(n7572), .dinb(n7567), .dout(n7573));
  jxor g07506(.dina(n7573), .dinb(\a[20] ), .dout(n7574));
  jxor g07507(.dina(n7574), .dinb(n7566), .dout(n7575));
  jxor g07508(.dina(n7575), .dinb(n7468), .dout(n7576));
  jnot g07509(.din(n7576), .dout(n7577));
  jor  g07510(.dina(n4038), .dinb(n2744), .dout(n7578));
  jor  g07511(.dina(n3863), .dinb(n2749), .dout(n7579));
  jor  g07512(.dina(n3929), .dinb(n2753), .dout(n7580));
  jand g07513(.dina(n7580), .dinb(n7579), .dout(n7581));
  jor  g07514(.dina(n3787), .dinb(n2758), .dout(n7582));
  jand g07515(.dina(n7582), .dinb(n7581), .dout(n7583));
  jand g07516(.dina(n7583), .dinb(n7578), .dout(n7584));
  jxor g07517(.dina(n7584), .dinb(\a[17] ), .dout(n7585));
  jxor g07518(.dina(n7585), .dinb(n7577), .dout(n7586));
  jxor g07519(.dina(n7586), .dinb(n7463), .dout(n7587));
  jor  g07520(.dina(n4726), .dinb(n3424), .dout(n7588));
  jor  g07521(.dina(n4471), .dinb(n3429), .dout(n7589));
  jor  g07522(.dina(n4019), .dinb(n3211), .dout(n7590));
  jor  g07523(.dina(n4596), .dinb(n3426), .dout(n7591));
  jand g07524(.dina(n7591), .dinb(n7590), .dout(n7592));
  jand g07525(.dina(n7592), .dinb(n7589), .dout(n7593));
  jand g07526(.dina(n7593), .dinb(n7588), .dout(n7594));
  jxor g07527(.dina(n7594), .dinb(n3473), .dout(n7595));
  jxor g07528(.dina(n7595), .dinb(n7587), .dout(n7596));
  jxor g07529(.dina(n7596), .dinb(n7460), .dout(n7597));
  jor  g07530(.dina(n5266), .dinb(n4023), .dout(n7598));
  jor  g07531(.dina(n4686), .dinb(n4028), .dout(n7599));
  jor  g07532(.dina(n4526), .dinb(n3871), .dout(n7600));
  jor  g07533(.dina(n5264), .dinb(n4025), .dout(n7601));
  jand g07534(.dina(n7601), .dinb(n7600), .dout(n7602));
  jand g07535(.dina(n7602), .dinb(n7599), .dout(n7603));
  jand g07536(.dina(n7603), .dinb(n7598), .dout(n7604));
  jxor g07537(.dina(n7604), .dinb(n4050), .dout(n7605));
  jxor g07538(.dina(n7605), .dinb(n7597), .dout(n7606));
  jxor g07539(.dina(n7606), .dinb(n7455), .dout(n7607));
  jor  g07540(.dina(n5527), .dinb(n4692), .dout(n7608));
  jor  g07541(.dina(n5364), .dinb(n4697), .dout(n7609));
  jor  g07542(.dina(n5525), .dinb(n4705), .dout(n7610));
  jand g07543(.dina(n7610), .dinb(n7609), .dout(n7611));
  jor  g07544(.dina(n5422), .dinb(n4702), .dout(n7612));
  jand g07545(.dina(n7612), .dinb(n7611), .dout(n7613));
  jand g07546(.dina(n7613), .dinb(n7608), .dout(n7614));
  jxor g07547(.dina(n7614), .dinb(\a[8] ), .dout(n7615));
  jnot g07548(.din(n7615), .dout(n7616));
  jxor g07549(.dina(n7616), .dinb(n7607), .dout(n7617));
  jxor g07550(.dina(n7617), .dinb(n7452), .dout(n7618));
  jor  g07551(.dina(n6999), .dinb(n5281), .dout(n7619));
  jor  g07552(.dina(n6390), .dinb(n5532), .dout(n7620));
  jor  g07553(.dina(n6205), .dinb(n5537), .dout(n7621));
  jor  g07554(.dina(n6297), .dinb(n5539), .dout(n7622));
  jand g07555(.dina(n7622), .dinb(n7621), .dout(n7623));
  jand g07556(.dina(n7623), .dinb(n7620), .dout(n7624));
  jand g07557(.dina(n7624), .dinb(n7619), .dout(n7625));
  jxor g07558(.dina(n7625), .dinb(n5277), .dout(n7626));
  jxor g07559(.dina(n7626), .dinb(n7618), .dout(n7627));
  jxor g07560(.dina(n7627), .dinb(n7448), .dout(n7628));
  jnot g07561(.din(n7301), .dout(n7629));
  jand g07562(.dina(n7629), .dinb(n7218), .dout(n7630));
  jnot g07563(.din(n7630), .dout(n7631));
  jnot g07564(.din(n7302), .dout(n7632));
  jor  g07565(.dina(n7632), .dinb(n7223), .dout(n7633));
  jand g07566(.dina(n7633), .dinb(n7631), .dout(n7634));
  jand g07567(.dina(n1273), .dinb(n175), .dout(n7635));
  jand g07568(.dina(n7635), .dinb(n517), .dout(n7636));
  jand g07569(.dina(n7288), .dinb(n2597), .dout(n7637));
  jand g07570(.dina(n7637), .dinb(n7636), .dout(n7638));
  jand g07571(.dina(n6335), .dinb(n1976), .dout(n7639));
  jand g07572(.dina(n532), .dinb(n1188), .dout(n7640));
  jand g07573(.dina(n7640), .dinb(n82), .dout(n7641));
  jand g07574(.dina(n7641), .dinb(n7639), .dout(n7642));
  jand g07575(.dina(n7642), .dinb(n7638), .dout(n7643));
  jand g07576(.dina(n7643), .dinb(n983), .dout(n7644));
  jand g07577(.dina(n7644), .dinb(n7279), .dout(n7645));
  jand g07578(.dina(n7645), .dinb(n1559), .dout(n7646));
  jand g07579(.dina(n7646), .dinb(n1897), .dout(n7647));
  jand g07580(.dina(n2100), .dinb(n537), .dout(n7648));
  jand g07581(.dina(n703), .dinb(n1325), .dout(n7649));
  jand g07582(.dina(n7649), .dinb(n7648), .dout(n7650));
  jand g07583(.dina(n7650), .dinb(n5340), .dout(n7651));
  jand g07584(.dina(n7651), .dinb(n1367), .dout(n7652));
  jand g07585(.dina(n3264), .dinb(n1753), .dout(n7653));
  jand g07586(.dina(n7653), .dinb(n694), .dout(n7654));
  jand g07587(.dina(n7654), .dinb(n902), .dout(n7655));
  jand g07588(.dina(n7655), .dinb(n7652), .dout(n7656));
  jand g07589(.dina(n1042), .dinb(n1218), .dout(n7657));
  jand g07590(.dina(n7657), .dinb(n3150), .dout(n7658));
  jand g07591(.dina(n7658), .dinb(n2148), .dout(n7659));
  jand g07592(.dina(n7659), .dinb(n465), .dout(n7660));
  jand g07593(.dina(n7660), .dinb(n7656), .dout(n7661));
  jand g07594(.dina(n6169), .dinb(n4417), .dout(n7662));
  jand g07595(.dina(n7662), .dinb(n6472), .dout(n7663));
  jand g07596(.dina(n7663), .dinb(n7661), .dout(n7664));
  jand g07597(.dina(n7664), .dinb(n7647), .dout(n7665));
  jand g07598(.dina(n1731), .dinb(n1309), .dout(n7666));
  jand g07599(.dina(n7666), .dinb(n6360), .dout(n7667));
  jand g07600(.dina(n1553), .dinb(n650), .dout(n7668));
  jand g07601(.dina(n7668), .dinb(n2693), .dout(n7669));
  jand g07602(.dina(n7669), .dinb(n7667), .dout(n7670));
  jand g07603(.dina(n7287), .dinb(n653), .dout(n7671));
  jand g07604(.dina(n5285), .dinb(n456), .dout(n7672));
  jand g07605(.dina(n7672), .dinb(n7671), .dout(n7673));
  jand g07606(.dina(n4528), .dinb(n2077), .dout(n7674));
  jand g07607(.dina(n7674), .dinb(n1207), .dout(n7675));
  jand g07608(.dina(n7675), .dinb(n7673), .dout(n7676));
  jand g07609(.dina(n7676), .dinb(n7670), .dout(n7677));
  jand g07610(.dina(n7677), .dinb(n843), .dout(n7678));
  jand g07611(.dina(n7678), .dinb(n1560), .dout(n7679));
  jand g07612(.dina(n7679), .dinb(n7665), .dout(n7680));
  jxor g07613(.dina(n7680), .dinb(n7301), .dout(n7681));
  jxor g07614(.dina(n7681), .dinb(n7634), .dout(n7682));
  jor  g07615(.dina(n7682), .dinb(n6496), .dout(n7683));
  jor  g07616(.dina(n7301), .dinb(n6507), .dout(n7684));
  jor  g07617(.dina(n7680), .dinb(n6504), .dout(n7685));
  jand g07618(.dina(n7685), .dinb(n7684), .dout(n7686));
  jor  g07619(.dina(n6501), .dinb(n6489), .dout(n7687));
  jand g07620(.dina(n7687), .dinb(n7686), .dout(n7688));
  jand g07621(.dina(n7688), .dinb(n7683), .dout(n7689));
  jxor g07622(.dina(n7689), .dinb(\a[2] ), .dout(n7690));
  jxor g07623(.dina(n7690), .dinb(n7628), .dout(n7691));
  jxor g07624(.dina(n7691), .dinb(n7443), .dout(n7692));
  jxor g07625(.dina(n7692), .dinb(n7326), .dout(n7693));
  jand g07626(.dina(n7693), .dinb(n806), .dout(n7694));
  jand g07627(.dina(n7019), .dinb(n1644), .dout(n7695));
  jor  g07628(.dina(n7695), .dinb(n7694), .dout(n7696));
  jand g07629(.dina(n7692), .dinb(n1620), .dout(n7697));
  jand g07630(.dina(n7313), .dinb(n1612), .dout(n7698));
  jor  g07631(.dina(n7698), .dinb(n7697), .dout(n7699));
  jor  g07632(.dina(n7699), .dinb(n7696), .dout(n7700));
  jnot g07633(.din(n7700), .dout(n7701));
  jand g07634(.dina(n7701), .dinb(n7325), .dout(n7702));
  jand g07635(.dina(n7702), .dinb(n7020), .dout(n7703));
  jnot g07636(.din(n7703), .dout(n7704));
  jxor g07637(.dina(n7702), .dinb(n7020), .dout(n7705));
  jnot g07638(.din(n7705), .dout(n7706));
  jor  g07639(.dina(n7690), .dinb(n7628), .dout(n7707));
  jnot g07640(.din(n7707), .dout(n7708));
  jand g07641(.dina(n7691), .dinb(n7443), .dout(n7709));
  jor  g07642(.dina(n7709), .dinb(n7708), .dout(n7710));
  jand g07643(.dina(n7626), .dinb(n7618), .dout(n7711));
  jand g07644(.dina(n7216), .dinb(n7033), .dout(n7712));
  jor  g07645(.dina(n7712), .dinb(n7444), .dout(n7713));
  jand g07646(.dina(n7627), .dinb(n7713), .dout(n7714));
  jor  g07647(.dina(n7714), .dinb(n7711), .dout(n7715));
  jand g07648(.dina(n7616), .dinb(n7607), .dout(n7716));
  jand g07649(.dina(n7617), .dinb(n7452), .dout(n7717));
  jor  g07650(.dina(n7717), .dinb(n7716), .dout(n7718));
  jand g07651(.dina(n7605), .dinb(n7597), .dout(n7719));
  jand g07652(.dina(n7606), .dinb(n7455), .dout(n7720));
  jor  g07653(.dina(n7720), .dinb(n7719), .dout(n7721));
  jand g07654(.dina(n7595), .dinb(n7587), .dout(n7722));
  jnot g07655(.din(n7722), .dout(n7723));
  jnot g07656(.din(n7460), .dout(n7724));
  jnot g07657(.din(n7596), .dout(n7725));
  jor  g07658(.dina(n7725), .dinb(n7724), .dout(n7726));
  jand g07659(.dina(n7726), .dinb(n7723), .dout(n7727));
  jor  g07660(.dina(n7585), .dinb(n7577), .dout(n7728));
  jnot g07661(.din(n7728), .dout(n7729));
  jand g07662(.dina(n7586), .dinb(n7463), .dout(n7730));
  jor  g07663(.dina(n7730), .dinb(n7729), .dout(n7731));
  jor  g07664(.dina(n7574), .dinb(n7566), .dout(n7732));
  jand g07665(.dina(n7575), .dinb(n7468), .dout(n7733));
  jnot g07666(.din(n7733), .dout(n7734));
  jand g07667(.dina(n7734), .dinb(n7732), .dout(n7735));
  jnot g07668(.din(n7735), .dout(n7736));
  jor  g07669(.dina(n7563), .dinb(n7555), .dout(n7737));
  jand g07670(.dina(n7564), .dinb(n7473), .dout(n7738));
  jnot g07671(.din(n7738), .dout(n7739));
  jand g07672(.dina(n7739), .dinb(n7737), .dout(n7740));
  jnot g07673(.din(n7740), .dout(n7741));
  jor  g07674(.dina(n7552), .dinb(n7544), .dout(n7742));
  jand g07675(.dina(n7553), .dinb(n7476), .dout(n7743));
  jnot g07676(.din(n7743), .dout(n7744));
  jand g07677(.dina(n7744), .dinb(n7742), .dout(n7745));
  jnot g07678(.din(n7745), .dout(n7746));
  jand g07679(.dina(n7541), .dinb(n7533), .dout(n7747));
  jand g07680(.dina(n7542), .dinb(n7479), .dout(n7748));
  jor  g07681(.dina(n7748), .dinb(n7747), .dout(n7749));
  jor  g07682(.dina(n4343), .dinb(n2176), .dout(n7750));
  jor  g07683(.dina(n4348), .dinb(n2174), .dout(n7751));
  jor  g07684(.dina(n3683), .dinb(n2057), .dout(n7752));
  jor  g07685(.dina(n4346), .dinb(n1954), .dout(n7753));
  jand g07686(.dina(n7753), .dinb(n7752), .dout(n7754));
  jand g07687(.dina(n7754), .dinb(n7751), .dout(n7755));
  jand g07688(.dina(n7755), .dinb(n7750), .dout(n7756));
  jxor g07689(.dina(n7756), .dinb(n93), .dout(n7757));
  jor  g07690(.dina(n7531), .dinb(n7523), .dout(n7758));
  jand g07691(.dina(n7532), .dinb(n7484), .dout(n7759));
  jnot g07692(.din(n7759), .dout(n7760));
  jand g07693(.dina(n7760), .dinb(n7758), .dout(n7761));
  jnot g07694(.din(n7761), .dout(n7762));
  jand g07695(.dina(n445), .dinb(n454), .dout(n7763));
  jand g07696(.dina(n7763), .dinb(n921), .dout(n7764));
  jand g07697(.dina(n718), .dinb(n1378), .dout(n7765));
  jand g07698(.dina(n7765), .dinb(n2023), .dout(n7766));
  jand g07699(.dina(n7766), .dinb(n1945), .dout(n7767));
  jand g07700(.dina(n7767), .dinb(n7764), .dout(n7768));
  jand g07701(.dina(n6474), .dinb(n901), .dout(n7769));
  jand g07702(.dina(n7769), .dinb(n1498), .dout(n7770));
  jand g07703(.dina(n1743), .dinb(n929), .dout(n7771));
  jand g07704(.dina(n7771), .dinb(n685), .dout(n7772));
  jand g07705(.dina(n4669), .dinb(n3385), .dout(n7773));
  jand g07706(.dina(n7773), .dinb(n7772), .dout(n7774));
  jand g07707(.dina(n7774), .dinb(n7770), .dout(n7775));
  jand g07708(.dina(n691), .dinb(n696), .dout(n7776));
  jand g07709(.dina(n7776), .dinb(n1583), .dout(n7777));
  jand g07710(.dina(n7777), .dinb(n501), .dout(n7778));
  jand g07711(.dina(n7778), .dinb(n2690), .dout(n7779));
  jand g07712(.dina(n7779), .dinb(n7775), .dout(n7780));
  jand g07713(.dina(n481), .dinb(n542), .dout(n7781));
  jand g07714(.dina(n1903), .dinb(n411), .dout(n7782));
  jand g07715(.dina(n7782), .dinb(n7781), .dout(n7783));
  jand g07716(.dina(n547), .dinb(n560), .dout(n7784));
  jand g07717(.dina(n7784), .dinb(n920), .dout(n7785));
  jand g07718(.dina(n7785), .dinb(n7783), .dout(n7786));
  jand g07719(.dina(n1708), .dinb(n1226), .dout(n7787));
  jand g07720(.dina(n7787), .dinb(n6010), .dout(n7788));
  jand g07721(.dina(n7788), .dinb(n7786), .dout(n7789));
  jand g07722(.dina(n7789), .dinb(n1977), .dout(n7790));
  jand g07723(.dina(n7790), .dinb(n7780), .dout(n7791));
  jand g07724(.dina(n7791), .dinb(n7768), .dout(n7792));
  jand g07725(.dina(n1522), .dinb(n1534), .dout(n7793));
  jand g07726(.dina(n7793), .dinb(n1237), .dout(n7794));
  jand g07727(.dina(n7794), .dinb(n1965), .dout(n7795));
  jand g07728(.dina(n7795), .dinb(n3363), .dout(n7796));
  jand g07729(.dina(n895), .dinb(n693), .dout(n7797));
  jand g07730(.dina(n7797), .dinb(n493), .dout(n7798));
  jand g07731(.dina(n7798), .dinb(n7796), .dout(n7799));
  jand g07732(.dina(n7799), .dinb(n6258), .dout(n7800));
  jand g07733(.dina(n7800), .dinb(n7792), .dout(n7801));
  jand g07734(.dina(n2708), .dinb(n1375), .dout(n7802));
  jand g07735(.dina(n7802), .dinb(n178), .dout(n7803));
  jand g07736(.dina(n461), .dinb(n699), .dout(n7804));
  jand g07737(.dina(n1506), .dinb(n668), .dout(n7805));
  jand g07738(.dina(n7805), .dinb(n7804), .dout(n7806));
  jand g07739(.dina(n7806), .dinb(n554), .dout(n7807));
  jand g07740(.dina(n7807), .dinb(n7803), .dout(n7808));
  jand g07741(.dina(n7808), .dinb(n2578), .dout(n7809));
  jand g07742(.dina(n1460), .dinb(n843), .dout(n7810));
  jand g07743(.dina(n7810), .dinb(n2350), .dout(n7811));
  jand g07744(.dina(n3007), .dinb(n1203), .dout(n7812));
  jand g07745(.dina(n7812), .dinb(n979), .dout(n7813));
  jand g07746(.dina(n7813), .dinb(n7811), .dout(n7814));
  jand g07747(.dina(n1756), .dinb(n900), .dout(n7815));
  jand g07748(.dina(n495), .dinb(n349), .dout(n7816));
  jand g07749(.dina(n7816), .dinb(n639), .dout(n7817));
  jand g07750(.dina(n7817), .dinb(n7815), .dout(n7818));
  jand g07751(.dina(n2086), .dinb(n1247), .dout(n7819));
  jand g07752(.dina(n7819), .dinb(n7818), .dout(n7820));
  jand g07753(.dina(n7820), .dinb(n1306), .dout(n7821));
  jand g07754(.dina(n7821), .dinb(n7814), .dout(n7822));
  jand g07755(.dina(n7822), .dinb(n7809), .dout(n7823));
  jand g07756(.dina(n5395), .dinb(n948), .dout(n7824));
  jand g07757(.dina(n7824), .dinb(n2345), .dout(n7825));
  jand g07758(.dina(n1865), .dinb(n470), .dout(n7826));
  jand g07759(.dina(n2100), .dinb(n965), .dout(n7827));
  jand g07760(.dina(n7827), .dinb(n660), .dout(n7828));
  jand g07761(.dina(n7828), .dinb(n7826), .dout(n7829));
  jand g07762(.dina(n7829), .dinb(n5415), .dout(n7830));
  jand g07763(.dina(n7830), .dinb(n7825), .dout(n7831));
  jand g07764(.dina(n2444), .dinb(n1449), .dout(n7832));
  jand g07765(.dina(n7832), .dinb(n1207), .dout(n7833));
  jand g07766(.dina(n7833), .dinb(n1316), .dout(n7834));
  jand g07767(.dina(n7834), .dinb(n2046), .dout(n7835));
  jand g07768(.dina(n7835), .dinb(n7831), .dout(n7836));
  jand g07769(.dina(n7836), .dinb(n7823), .dout(n7837));
  jand g07770(.dina(n7837), .dinb(n7801), .dout(n7838));
  jor  g07771(.dina(n7061), .dinb(n1792), .dout(n7839));
  jand g07772(.dina(n5084), .dinb(n2061), .dout(n7840));
  jand g07773(.dina(n5082), .dinb(n1673), .dout(n7841));
  jor  g07774(.dina(n7841), .dinb(n7840), .dout(n7842));
  jand g07775(.dina(n6050), .dinb(n1024), .dout(n7843));
  jor  g07776(.dina(n7843), .dinb(n7842), .dout(n7844));
  jnot g07777(.din(n7844), .dout(n7845));
  jand g07778(.dina(n7845), .dinb(n7839), .dout(n7846));
  jxor g07779(.dina(n7846), .dinb(n7838), .dout(n7847));
  jxor g07780(.dina(n7847), .dinb(n7762), .dout(n7848));
  jxor g07781(.dina(n7848), .dinb(n7757), .dout(n7849));
  jxor g07782(.dina(n7849), .dinb(n7749), .dout(n7850));
  jor  g07783(.dina(n2768), .dinb(n2303), .dout(n7851));
  jor  g07784(.dina(n2553), .dinb(n2309), .dout(n7852));
  jor  g07785(.dina(n2428), .dinb(n1805), .dout(n7853));
  jor  g07786(.dina(n2629), .dinb(n2306), .dout(n7854));
  jand g07787(.dina(n7854), .dinb(n7853), .dout(n7855));
  jand g07788(.dina(n7855), .dinb(n7852), .dout(n7856));
  jand g07789(.dina(n7856), .dinb(n7851), .dout(n7857));
  jxor g07790(.dina(n7857), .dinb(n77), .dout(n7858));
  jxor g07791(.dina(n7858), .dinb(n7850), .dout(n7859));
  jxor g07792(.dina(n7859), .dinb(n7746), .dout(n7860));
  jnot g07793(.din(n7860), .dout(n7861));
  jor  g07794(.dina(n3451), .dinb(n807), .dout(n7862));
  jor  g07795(.dina(n3072), .dinb(n1613), .dout(n7863));
  jor  g07796(.dina(n2738), .dinb(n1617), .dout(n7864));
  jand g07797(.dina(n7864), .dinb(n7863), .dout(n7865));
  jor  g07798(.dina(n3203), .dinb(n1621), .dout(n7866));
  jand g07799(.dina(n7866), .dinb(n7865), .dout(n7867));
  jand g07800(.dina(n7867), .dinb(n7862), .dout(n7868));
  jxor g07801(.dina(n7868), .dinb(\a[23] ), .dout(n7869));
  jxor g07802(.dina(n7869), .dinb(n7861), .dout(n7870));
  jxor g07803(.dina(n7870), .dinb(n7741), .dout(n7871));
  jnot g07804(.din(n7871), .dout(n7872));
  jor  g07805(.dina(n3789), .dinb(n1820), .dout(n7873));
  jor  g07806(.dina(n3420), .dinb(n2181), .dout(n7874));
  jor  g07807(.dina(n3286), .dinb(n2186), .dout(n7875));
  jand g07808(.dina(n7875), .dinb(n7874), .dout(n7876));
  jor  g07809(.dina(n3787), .dinb(n2189), .dout(n7877));
  jand g07810(.dina(n7877), .dinb(n7876), .dout(n7878));
  jand g07811(.dina(n7878), .dinb(n7873), .dout(n7879));
  jxor g07812(.dina(n7879), .dinb(\a[20] ), .dout(n7880));
  jxor g07813(.dina(n7880), .dinb(n7872), .dout(n7881));
  jxor g07814(.dina(n7881), .dinb(n7736), .dout(n7882));
  jnot g07815(.din(n7882), .dout(n7883));
  jor  g07816(.dina(n3863), .dinb(n2758), .dout(n7884));
  jor  g07817(.dina(n4021), .dinb(n2744), .dout(n7885));
  jor  g07818(.dina(n4019), .dinb(n2753), .dout(n7886));
  jor  g07819(.dina(n3929), .dinb(n2749), .dout(n7887));
  jand g07820(.dina(n7887), .dinb(n7886), .dout(n7888));
  jand g07821(.dina(n7888), .dinb(n7885), .dout(n7889));
  jand g07822(.dina(n7889), .dinb(n7884), .dout(n7890));
  jxor g07823(.dina(n7890), .dinb(\a[17] ), .dout(n7891));
  jxor g07824(.dina(n7891), .dinb(n7883), .dout(n7892));
  jxor g07825(.dina(n7892), .dinb(n7731), .dout(n7893));
  jor  g07826(.dina(n4714), .dinb(n3424), .dout(n7894));
  jor  g07827(.dina(n4596), .dinb(n3429), .dout(n7895));
  jor  g07828(.dina(n4471), .dinb(n3211), .dout(n7896));
  jor  g07829(.dina(n4526), .dinb(n3426), .dout(n7897));
  jand g07830(.dina(n7897), .dinb(n7896), .dout(n7898));
  jand g07831(.dina(n7898), .dinb(n7895), .dout(n7899));
  jand g07832(.dina(n7899), .dinb(n7894), .dout(n7900));
  jxor g07833(.dina(n7900), .dinb(n3473), .dout(n7901));
  jxor g07834(.dina(n7901), .dinb(n7893), .dout(n7902));
  jnot g07835(.din(n7902), .dout(n7903));
  jxor g07836(.dina(n7903), .dinb(n7727), .dout(n7904));
  jor  g07837(.dina(n5560), .dinb(n4023), .dout(n7905));
  jor  g07838(.dina(n5264), .dinb(n4028), .dout(n7906));
  jor  g07839(.dina(n4686), .dinb(n3871), .dout(n7907));
  jor  g07840(.dina(n5422), .dinb(n4025), .dout(n7908));
  jand g07841(.dina(n7908), .dinb(n7907), .dout(n7909));
  jand g07842(.dina(n7909), .dinb(n7906), .dout(n7910));
  jand g07843(.dina(n7910), .dinb(n7905), .dout(n7911));
  jxor g07844(.dina(n7911), .dinb(n4050), .dout(n7912));
  jxor g07845(.dina(n7912), .dinb(n7904), .dout(n7913));
  jxor g07846(.dina(n7913), .dinb(n7721), .dout(n7914));
  jor  g07847(.dina(n6207), .dinb(n4692), .dout(n7915));
  jor  g07848(.dina(n5525), .dinb(n4697), .dout(n7916));
  jor  g07849(.dina(n6205), .dinb(n4705), .dout(n7917));
  jor  g07850(.dina(n5364), .dinb(n4702), .dout(n7918));
  jand g07851(.dina(n7918), .dinb(n7917), .dout(n7919));
  jand g07852(.dina(n7919), .dinb(n7916), .dout(n7920));
  jand g07853(.dina(n7920), .dinb(n7915), .dout(n7921));
  jxor g07854(.dina(n7921), .dinb(n4713), .dout(n7922));
  jxor g07855(.dina(n7922), .dinb(n7914), .dout(n7923));
  jxor g07856(.dina(n7923), .dinb(n7718), .dout(n7924));
  jor  g07857(.dina(n6491), .dinb(n5281), .dout(n7925));
  jor  g07858(.dina(n6297), .dinb(n5532), .dout(n7926));
  jor  g07859(.dina(n6390), .dinb(n5537), .dout(n7927));
  jand g07860(.dina(n7927), .dinb(n7926), .dout(n7928));
  jor  g07861(.dina(n6489), .dinb(n5539), .dout(n7929));
  jand g07862(.dina(n7929), .dinb(n7928), .dout(n7930));
  jand g07863(.dina(n7930), .dinb(n7925), .dout(n7931));
  jxor g07864(.dina(n7931), .dinb(\a[5] ), .dout(n7932));
  jxor g07865(.dina(n7932), .dinb(n7924), .dout(n7933));
  jxor g07866(.dina(n7933), .dinb(n7715), .dout(n7934));
  jnot g07867(.din(n7680), .dout(n7935));
  jand g07868(.dina(n7935), .dinb(n7629), .dout(n7936));
  jand g07869(.dina(n3421), .dinb(n6703), .dout(n7937));
  jor  g07870(.dina(n7937), .dinb(n3730), .dout(n7938));
  jand g07871(.dina(n3788), .dinb(n7938), .dout(n7939));
  jor  g07872(.dina(n7939), .dinb(n3936), .dout(n7940));
  jand g07873(.dina(n3941), .dinb(n7940), .dout(n7941));
  jor  g07874(.dina(n7941), .dinb(n3934), .dout(n7942));
  jand g07875(.dina(n3945), .dinb(n7942), .dout(n7943));
  jor  g07876(.dina(n7943), .dinb(n3931), .dout(n7944));
  jand g07877(.dina(n4020), .dinb(n7944), .dout(n7945));
  jor  g07878(.dina(n7945), .dinb(n4407), .dout(n7946));
  jand g07879(.dina(n4472), .dinb(n7946), .dout(n7947));
  jor  g07880(.dina(n7947), .dinb(n4603), .dout(n7948));
  jand g07881(.dina(n4608), .dinb(n7948), .dout(n7949));
  jor  g07882(.dina(n7949), .dinb(n4601), .dout(n7950));
  jand g07883(.dina(n4612), .dinb(n7950), .dout(n7951));
  jor  g07884(.dina(n7951), .dinb(n4598), .dout(n7952));
  jand g07885(.dina(n4687), .dinb(n7952), .dout(n7953));
  jor  g07886(.dina(n7953), .dinb(n5164), .dout(n7954));
  jand g07887(.dina(n5265), .dinb(n7954), .dout(n7955));
  jor  g07888(.dina(n7955), .dinb(n5429), .dout(n7956));
  jand g07889(.dina(n5434), .dinb(n7956), .dout(n7957));
  jor  g07890(.dina(n7957), .dinb(n5427), .dout(n7958));
  jand g07891(.dina(n5438), .dinb(n7958), .dout(n7959));
  jor  g07892(.dina(n7959), .dinb(n5424), .dout(n7960));
  jand g07893(.dina(n5526), .dinb(n7960), .dout(n7961));
  jor  g07894(.dina(n7961), .dinb(n6141), .dout(n7962));
  jand g07895(.dina(n6206), .dinb(n7962), .dout(n7963));
  jor  g07896(.dina(n7963), .dinb(n6397), .dout(n7964));
  jand g07897(.dina(n6402), .dinb(n7964), .dout(n7965));
  jor  g07898(.dina(n7965), .dinb(n6395), .dout(n7966));
  jand g07899(.dina(n6406), .dinb(n7966), .dout(n7967));
  jor  g07900(.dina(n7967), .dinb(n6392), .dout(n7968));
  jand g07901(.dina(n6490), .dinb(n7968), .dout(n7969));
  jor  g07902(.dina(n7969), .dinb(n7219), .dout(n7970));
  jand g07903(.dina(n7302), .dinb(n7970), .dout(n7971));
  jor  g07904(.dina(n7971), .dinb(n7630), .dout(n7972));
  jand g07905(.dina(n7681), .dinb(n7972), .dout(n7973));
  jor  g07906(.dina(n7973), .dinb(n7936), .dout(n7974));
  jand g07907(.dina(n7297), .dinb(n1560), .dout(n7975));
  jand g07908(.dina(n3014), .dinb(n1427), .dout(n7976));
  jand g07909(.dina(n1227), .dinb(n1040), .dout(n7977));
  jand g07910(.dina(n7977), .dinb(n994), .dout(n7978));
  jand g07911(.dina(n7978), .dinb(n7976), .dout(n7979));
  jand g07912(.dina(n3752), .dinb(n1768), .dout(n7980));
  jand g07913(.dina(n7980), .dinb(n1863), .dout(n7981));
  jand g07914(.dina(n7981), .dinb(n7979), .dout(n7982));
  jand g07915(.dina(n1238), .dinb(n920), .dout(n7983));
  jand g07916(.dina(n7983), .dinb(n948), .dout(n7984));
  jand g07917(.dina(n1506), .dinb(n469), .dout(n7985));
  jand g07918(.dina(n7985), .dinb(n2595), .dout(n7986));
  jand g07919(.dina(n7986), .dinb(n7984), .dout(n7987));
  jand g07920(.dina(n4448), .dinb(n3782), .dout(n7988));
  jand g07921(.dina(n7988), .dinb(n7987), .dout(n7989));
  jand g07922(.dina(n7989), .dinb(n7982), .dout(n7990));
  jand g07923(.dina(n1460), .dinb(n1016), .dout(n7991));
  jand g07924(.dina(n7991), .dinb(n1361), .dout(n7992));
  jand g07925(.dina(n2024), .dinb(n1735), .dout(n7993));
  jand g07926(.dina(n7993), .dinb(n7992), .dout(n7994));
  jand g07927(.dina(n7994), .dinb(n1900), .dout(n7995));
  jand g07928(.dina(n7995), .dinb(n7990), .dout(n7996));
  jand g07929(.dina(n7996), .dinb(n583), .dout(n7997));
  jand g07930(.dina(n7997), .dinb(n7975), .dout(n7998));
  jand g07931(.dina(n7998), .dinb(n7677), .dout(n7999));
  jnot g07932(.din(n7999), .dout(n8000));
  jxor g07933(.dina(n8000), .dinb(n7680), .dout(n8001));
  jxor g07934(.dina(n8001), .dinb(n7974), .dout(n8002));
  jor  g07935(.dina(n8002), .dinb(n6496), .dout(n8003));
  jand g07936(.dina(n8000), .dinb(n6503), .dout(n8004));
  jand g07937(.dina(n7935), .dinb(n6506), .dout(n8005));
  jor  g07938(.dina(n8005), .dinb(n8004), .dout(n8006));
  jnot g07939(.din(n8006), .dout(n8007));
  jand g07940(.dina(n8007), .dinb(n8003), .dout(n8008));
  jor  g07941(.dina(n8008), .dinb(\a[2] ), .dout(n8009));
  jnot g07942(.din(n7936), .dout(n8010));
  jnot g07943(.din(n7681), .dout(n8011));
  jor  g07944(.dina(n8011), .dinb(n7634), .dout(n8012));
  jand g07945(.dina(n8012), .dinb(n8010), .dout(n8013));
  jxor g07946(.dina(n8001), .dinb(n8013), .dout(n8014));
  jand g07947(.dina(n8014), .dinb(n6495), .dout(n8015));
  jor  g07948(.dina(n8006), .dinb(n8015), .dout(n8016));
  jand g07949(.dina(n7629), .dinb(n6500), .dout(n8017));
  jor  g07950(.dina(n8017), .dinb(n6219), .dout(n8018));
  jor  g07951(.dina(n8018), .dinb(n8016), .dout(n8019));
  jand g07952(.dina(n8019), .dinb(n8009), .dout(n8020));
  jxor g07953(.dina(n8020), .dinb(n7934), .dout(n8021));
  jxor g07954(.dina(n8021), .dinb(n7710), .dout(n8022));
  jxor g07955(.dina(n8022), .dinb(n7692), .dout(n8023));
  jnot g07956(.din(n7313), .dout(n8024));
  jnot g07957(.din(n7692), .dout(n8025));
  jand g07958(.dina(n8025), .dinb(n7021), .dout(n8026));
  jor  g07959(.dina(n8026), .dinb(n8024), .dout(n8027));
  jnot g07960(.din(n8027), .dout(n8028));
  jxor g07961(.dina(n8028), .dinb(n8023), .dout(n8029));
  jand g07962(.dina(n8029), .dinb(n806), .dout(n8030));
  jand g07963(.dina(n7692), .dinb(n1612), .dout(n8031));
  jand g07964(.dina(n8022), .dinb(n1620), .dout(n8032));
  jor  g07965(.dina(n8032), .dinb(n8031), .dout(n8033));
  jand g07966(.dina(n7313), .dinb(n1644), .dout(n8034));
  jor  g07967(.dina(n8034), .dinb(n8033), .dout(n8035));
  jor  g07968(.dina(n8035), .dinb(n8030), .dout(n8036));
  jxor g07969(.dina(n8036), .dinb(n65), .dout(n8037));
  jor  g07970(.dina(n8037), .dinb(n7706), .dout(n8038));
  jand g07971(.dina(n8038), .dinb(n7704), .dout(n8039));
  jnot g07972(.din(n8039), .dout(n8040));
  jand g07973(.dina(n7315), .dinb(n71), .dout(n8041));
  jand g07974(.dina(n7313), .dinb(n796), .dout(n8042));
  jand g07975(.dina(n7019), .dinb(n731), .dout(n8043));
  jor  g07976(.dina(n8043), .dinb(n8042), .dout(n8044));
  jor  g07977(.dina(n8044), .dinb(n8041), .dout(n8045));
  jnot g07978(.din(n7020), .dout(n8046));
  jor  g07979(.dina(n8046), .dinb(n77), .dout(n8047));
  jxor g07980(.dina(n8047), .dinb(n8045), .dout(n8048));
  jand g07981(.dina(n8022), .dinb(n7692), .dout(n8049));
  jand g07982(.dina(n8028), .dinb(n8023), .dout(n8050));
  jor  g07983(.dina(n8050), .dinb(n8049), .dout(n8051));
  jnot g07984(.din(n7932), .dout(n8052));
  jxor g07985(.dina(n8052), .dinb(n7924), .dout(n8053));
  jxor g07986(.dina(n8053), .dinb(n7715), .dout(n8054));
  jand g07987(.dina(n8016), .dinb(n6219), .dout(n8055));
  jnot g07988(.din(n8018), .dout(n8056));
  jand g07989(.dina(n8056), .dinb(n8008), .dout(n8057));
  jor  g07990(.dina(n8057), .dinb(n8055), .dout(n8058));
  jand g07991(.dina(n8058), .dinb(n8054), .dout(n8059));
  jand g07992(.dina(n8021), .dinb(n7710), .dout(n8060));
  jor  g07993(.dina(n8060), .dinb(n8059), .dout(n8061));
  jand g07994(.dina(n8052), .dinb(n7924), .dout(n8062));
  jand g07995(.dina(n8053), .dinb(n7715), .dout(n8063));
  jor  g07996(.dina(n8063), .dinb(n8062), .dout(n8064));
  jand g07997(.dina(n7922), .dinb(n7914), .dout(n8065));
  jand g07998(.dina(n7923), .dinb(n7718), .dout(n8066));
  jor  g07999(.dina(n8066), .dinb(n8065), .dout(n8067));
  jand g08000(.dina(n7912), .dinb(n7904), .dout(n8068));
  jand g08001(.dina(n7913), .dinb(n7721), .dout(n8069));
  jor  g08002(.dina(n8069), .dinb(n8068), .dout(n8070));
  jand g08003(.dina(n7901), .dinb(n7893), .dout(n8071));
  jnot g08004(.din(n8071), .dout(n8072));
  jor  g08005(.dina(n7903), .dinb(n7727), .dout(n8073));
  jand g08006(.dina(n8073), .dinb(n8072), .dout(n8074));
  jor  g08007(.dina(n7891), .dinb(n7883), .dout(n8075));
  jand g08008(.dina(n7892), .dinb(n7731), .dout(n8076));
  jnot g08009(.din(n8076), .dout(n8077));
  jand g08010(.dina(n8077), .dinb(n8075), .dout(n8078));
  jor  g08011(.dina(n7880), .dinb(n7872), .dout(n8079));
  jand g08012(.dina(n7881), .dinb(n7736), .dout(n8080));
  jnot g08013(.din(n8080), .dout(n8081));
  jand g08014(.dina(n8081), .dinb(n8079), .dout(n8082));
  jnot g08015(.din(n8082), .dout(n8083));
  jor  g08016(.dina(n7869), .dinb(n7861), .dout(n8084));
  jand g08017(.dina(n7870), .dinb(n7741), .dout(n8085));
  jnot g08018(.din(n8085), .dout(n8086));
  jand g08019(.dina(n8086), .dinb(n8084), .dout(n8087));
  jnot g08020(.din(n8087), .dout(n8088));
  jand g08021(.dina(n7858), .dinb(n7850), .dout(n8089));
  jand g08022(.dina(n7859), .dinb(n7746), .dout(n8090));
  jor  g08023(.dina(n8090), .dinb(n8089), .dout(n8091));
  jand g08024(.dina(n7848), .dinb(n7757), .dout(n8092));
  jand g08025(.dina(n7849), .dinb(n7749), .dout(n8093));
  jor  g08026(.dina(n8093), .dinb(n8092), .dout(n8094));
  jor  g08027(.dina(n7846), .dinb(n7838), .dout(n8095));
  jand g08028(.dina(n7847), .dinb(n7762), .dout(n8096));
  jnot g08029(.din(n8096), .dout(n8097));
  jand g08030(.dina(n8097), .dinb(n8095), .dout(n8098));
  jnot g08031(.din(n8098), .dout(n8099));
  jand g08032(.dina(n4639), .dinb(n3179), .dout(n8100));
  jand g08033(.dina(n8100), .dinb(n1358), .dout(n8101));
  jand g08034(.dina(n3985), .dinb(n2400), .dout(n8102));
  jand g08035(.dina(n8102), .dinb(n2152), .dout(n8103));
  jand g08036(.dina(n8103), .dinb(n1936), .dout(n8104));
  jand g08037(.dina(n548), .dinb(n2117), .dout(n8105));
  jand g08038(.dina(n8105), .dinb(n1367), .dout(n8106));
  jand g08039(.dina(n3217), .dinb(n1735), .dout(n8107));
  jand g08040(.dina(n8107), .dinb(n3116), .dout(n8108));
  jand g08041(.dina(n8108), .dinb(n8106), .dout(n8109));
  jand g08042(.dina(n8109), .dinb(n8104), .dout(n8110));
  jand g08043(.dina(n8110), .dinb(n5382), .dout(n8111));
  jand g08044(.dina(n8111), .dinb(n8101), .dout(n8112));
  jand g08045(.dina(n1107), .dinb(n542), .dout(n8113));
  jand g08046(.dina(n480), .dinb(n1225), .dout(n8114));
  jand g08047(.dina(n8114), .dinb(n8113), .dout(n8115));
  jnot g08048(.din(n1086), .dout(n8116));
  jand g08049(.dina(n1867), .dinb(n639), .dout(n8117));
  jand g08050(.dina(n8117), .dinb(n873), .dout(n8118));
  jand g08051(.dina(n8118), .dinb(n8116), .dout(n8119));
  jand g08052(.dina(n1159), .dinb(n826), .dout(n8120));
  jand g08053(.dina(n8120), .dinb(n1562), .dout(n8121));
  jand g08054(.dina(n8121), .dinb(n1580), .dout(n8122));
  jand g08055(.dina(n8122), .dinb(n8119), .dout(n8123));
  jand g08056(.dina(n8123), .dinb(n8115), .dout(n8124));
  jand g08057(.dina(n472), .dinb(n676), .dout(n8125));
  jand g08058(.dina(n8125), .dinb(n114), .dout(n8126));
  jand g08059(.dina(n1316), .dinb(n135), .dout(n8127));
  jand g08060(.dina(n8127), .dinb(n1846), .dout(n8128));
  jand g08061(.dina(n8128), .dinb(n8126), .dout(n8129));
  jand g08062(.dina(n5415), .dinb(n2588), .dout(n8130));
  jand g08063(.dina(n3014), .dinb(n697), .dout(n8131));
  jand g08064(.dina(n8131), .dinb(n8130), .dout(n8132));
  jand g08065(.dina(n8132), .dinb(n8129), .dout(n8133));
  jand g08066(.dina(n1756), .dinb(n171), .dout(n8134));
  jand g08067(.dina(n452), .dinb(n699), .dout(n8135));
  jand g08068(.dina(n8135), .dinb(n8134), .dout(n8136));
  jand g08069(.dina(n621), .dinb(n461), .dout(n8137));
  jand g08070(.dina(n8137), .dinb(n917), .dout(n8138));
  jand g08071(.dina(n8138), .dinb(n8136), .dout(n8139));
  jand g08072(.dina(n8139), .dinb(n5994), .dout(n8140));
  jand g08073(.dina(n8140), .dinb(n8133), .dout(n8141));
  jand g08074(.dina(n2521), .dinb(n320), .dout(n8142));
  jand g08075(.dina(n647), .dinb(n541), .dout(n8143));
  jand g08076(.dina(n8143), .dinb(n8142), .dout(n8144));
  jand g08077(.dina(n8144), .dinb(n6334), .dout(n8145));
  jand g08078(.dina(n1214), .dinb(n818), .dout(n8146));
  jand g08079(.dina(n8146), .dinb(n8145), .dout(n8147));
  jand g08080(.dina(n8147), .dinb(n8141), .dout(n8148));
  jand g08081(.dina(n8148), .dinb(n8124), .dout(n8149));
  jand g08082(.dina(n8149), .dinb(n8112), .dout(n8150));
  jor  g08083(.dina(n7061), .dinb(n2208), .dout(n8151));
  jand g08084(.dina(n5082), .dinb(n2061), .dout(n8152));
  jand g08085(.dina(n5084), .dinb(n2058), .dout(n8153));
  jor  g08086(.dina(n8153), .dinb(n8152), .dout(n8154));
  jand g08087(.dina(n6050), .dinb(n1673), .dout(n8155));
  jor  g08088(.dina(n8155), .dinb(n8154), .dout(n8156));
  jnot g08089(.din(n8156), .dout(n8157));
  jand g08090(.dina(n8157), .dinb(n8151), .dout(n8158));
  jxor g08091(.dina(n8158), .dinb(n8150), .dout(n8159));
  jxor g08092(.dina(n8159), .dinb(n8099), .dout(n8160));
  jor  g08093(.dina(n4343), .dinb(n2430), .dout(n8161));
  jor  g08094(.dina(n4346), .dinb(n2174), .dout(n8162));
  jor  g08095(.dina(n4348), .dinb(n2428), .dout(n8163));
  jor  g08096(.dina(n3683), .dinb(n1954), .dout(n8164));
  jand g08097(.dina(n8164), .dinb(n8163), .dout(n8165));
  jand g08098(.dina(n8165), .dinb(n8162), .dout(n8166));
  jand g08099(.dina(n8166), .dinb(n8161), .dout(n8167));
  jxor g08100(.dina(n8167), .dinb(n93), .dout(n8168));
  jxor g08101(.dina(n8168), .dinb(n8160), .dout(n8169));
  jxor g08102(.dina(n8169), .dinb(n8094), .dout(n8170));
  jnot g08103(.din(n8170), .dout(n8171));
  jor  g08104(.dina(n2740), .dinb(n2303), .dout(n8172));
  jor  g08105(.dina(n2553), .dinb(n2306), .dout(n8173));
  jor  g08106(.dina(n2629), .dinb(n1805), .dout(n8174));
  jand g08107(.dina(n8174), .dinb(n8173), .dout(n8175));
  jor  g08108(.dina(n2738), .dinb(n2309), .dout(n8176));
  jand g08109(.dina(n8176), .dinb(n8175), .dout(n8177));
  jand g08110(.dina(n8177), .dinb(n8172), .dout(n8178));
  jxor g08111(.dina(n8178), .dinb(\a[26] ), .dout(n8179));
  jxor g08112(.dina(n8179), .dinb(n8171), .dout(n8180));
  jxor g08113(.dina(n8180), .dinb(n8091), .dout(n8181));
  jnot g08114(.din(n8181), .dout(n8182));
  jor  g08115(.dina(n3440), .dinb(n807), .dout(n8183));
  jor  g08116(.dina(n3203), .dinb(n1613), .dout(n8184));
  jor  g08117(.dina(n3286), .dinb(n1621), .dout(n8185));
  jand g08118(.dina(n8185), .dinb(n8184), .dout(n8186));
  jor  g08119(.dina(n3072), .dinb(n1617), .dout(n8187));
  jand g08120(.dina(n8187), .dinb(n8186), .dout(n8188));
  jand g08121(.dina(n8188), .dinb(n8183), .dout(n8189));
  jxor g08122(.dina(n8189), .dinb(\a[23] ), .dout(n8190));
  jxor g08123(.dina(n8190), .dinb(n8182), .dout(n8191));
  jxor g08124(.dina(n8191), .dinb(n8088), .dout(n8192));
  jor  g08125(.dina(n4051), .dinb(n1820), .dout(n8193));
  jor  g08126(.dina(n3787), .dinb(n2181), .dout(n8194));
  jor  g08127(.dina(n3863), .dinb(n2189), .dout(n8195));
  jor  g08128(.dina(n3420), .dinb(n2186), .dout(n8196));
  jand g08129(.dina(n8196), .dinb(n8195), .dout(n8197));
  jand g08130(.dina(n8197), .dinb(n8194), .dout(n8198));
  jand g08131(.dina(n8198), .dinb(n8193), .dout(n8199));
  jxor g08132(.dina(n8199), .dinb(n2196), .dout(n8200));
  jxor g08133(.dina(n8200), .dinb(n8192), .dout(n8201));
  jxor g08134(.dina(n8201), .dinb(n8083), .dout(n8202));
  jor  g08135(.dina(n4473), .dinb(n2744), .dout(n8203));
  jor  g08136(.dina(n4019), .dinb(n2749), .dout(n8204));
  jor  g08137(.dina(n3929), .dinb(n2758), .dout(n8205));
  jor  g08138(.dina(n4471), .dinb(n2753), .dout(n8206));
  jand g08139(.dina(n8206), .dinb(n8205), .dout(n8207));
  jand g08140(.dina(n8207), .dinb(n8204), .dout(n8208));
  jand g08141(.dina(n8208), .dinb(n8203), .dout(n8209));
  jxor g08142(.dina(n8209), .dinb(n2441), .dout(n8210));
  jxor g08143(.dina(n8210), .dinb(n8202), .dout(n8211));
  jxor g08144(.dina(n8211), .dinb(n8078), .dout(n8212));
  jor  g08145(.dina(n4688), .dinb(n3424), .dout(n8213));
  jor  g08146(.dina(n4526), .dinb(n3429), .dout(n8214));
  jor  g08147(.dina(n4596), .dinb(n3211), .dout(n8215));
  jand g08148(.dina(n8215), .dinb(n8214), .dout(n8216));
  jor  g08149(.dina(n4686), .dinb(n3426), .dout(n8217));
  jand g08150(.dina(n8217), .dinb(n8216), .dout(n8218));
  jand g08151(.dina(n8218), .dinb(n8213), .dout(n8219));
  jxor g08152(.dina(n8219), .dinb(\a[14] ), .dout(n8220));
  jxor g08153(.dina(n8220), .dinb(n8212), .dout(n8221));
  jxor g08154(.dina(n8221), .dinb(n8074), .dout(n8222));
  jor  g08155(.dina(n5549), .dinb(n4023), .dout(n8223));
  jor  g08156(.dina(n5422), .dinb(n4028), .dout(n8224));
  jor  g08157(.dina(n5264), .dinb(n3871), .dout(n8225));
  jand g08158(.dina(n8225), .dinb(n8224), .dout(n8226));
  jor  g08159(.dina(n5364), .dinb(n4025), .dout(n8227));
  jand g08160(.dina(n8227), .dinb(n8226), .dout(n8228));
  jand g08161(.dina(n8228), .dinb(n8223), .dout(n8229));
  jxor g08162(.dina(n8229), .dinb(\a[11] ), .dout(n8230));
  jxor g08163(.dina(n8230), .dinb(n8222), .dout(n8231));
  jxor g08164(.dina(n8231), .dinb(n8070), .dout(n8232));
  jor  g08165(.dina(n6516), .dinb(n4692), .dout(n8233));
  jor  g08166(.dina(n6205), .dinb(n4697), .dout(n8234));
  jor  g08167(.dina(n5525), .dinb(n4702), .dout(n8235));
  jor  g08168(.dina(n6390), .dinb(n4705), .dout(n8236));
  jand g08169(.dina(n8236), .dinb(n8235), .dout(n8237));
  jand g08170(.dina(n8237), .dinb(n8234), .dout(n8238));
  jand g08171(.dina(n8238), .dinb(n8233), .dout(n8239));
  jxor g08172(.dina(n8239), .dinb(n4713), .dout(n8240));
  jxor g08173(.dina(n8240), .dinb(n8232), .dout(n8241));
  jxor g08174(.dina(n8241), .dinb(n8067), .dout(n8242));
  jor  g08175(.dina(n7303), .dinb(n5281), .dout(n8243));
  jor  g08176(.dina(n7301), .dinb(n5539), .dout(n8244));
  jor  g08177(.dina(n6297), .dinb(n5537), .dout(n8245));
  jor  g08178(.dina(n6489), .dinb(n5532), .dout(n8246));
  jand g08179(.dina(n8246), .dinb(n8245), .dout(n8247));
  jand g08180(.dina(n8247), .dinb(n8244), .dout(n8248));
  jand g08181(.dina(n8248), .dinb(n8243), .dout(n8249));
  jxor g08182(.dina(n8249), .dinb(n5277), .dout(n8250));
  jxor g08183(.dina(n8250), .dinb(n8242), .dout(n8251));
  jnot g08184(.din(n8251), .dout(n8252));
  jxor g08185(.dina(n8252), .dinb(n8064), .dout(n8253));
  jnot g08186(.din(n8001), .dout(n8254));
  jand g08187(.dina(n8254), .dinb(n7974), .dout(n8255));
  jor  g08188(.dina(n8255), .dinb(n7935), .dout(n8256));
  jand g08189(.dina(n8256), .dinb(n8000), .dout(n8257));
  jor  g08190(.dina(n8001), .dinb(n8013), .dout(n8258));
  jand g08191(.dina(n8258), .dinb(n7999), .dout(n8259));
  jor  g08192(.dina(n8259), .dinb(n8257), .dout(n8260));
  jor  g08193(.dina(n8260), .dinb(n6496), .dout(n8261));
  jor  g08194(.dina(n7680), .dinb(n6501), .dout(n8262));
  jor  g08195(.dina(n7999), .dinb(n6507), .dout(n8263));
  jand g08196(.dina(n8263), .dinb(n8262), .dout(n8264));
  jand g08197(.dina(n8264), .dinb(n8261), .dout(n8265));
  jxor g08198(.dina(n8265), .dinb(\a[2] ), .dout(n8266));
  jxor g08199(.dina(n8266), .dinb(n8253), .dout(n8267));
  jxor g08200(.dina(n8267), .dinb(n8061), .dout(n8268));
  jxor g08201(.dina(n8268), .dinb(n8022), .dout(n8269));
  jxor g08202(.dina(n8269), .dinb(n8051), .dout(n8270));
  jand g08203(.dina(n8270), .dinb(n806), .dout(n8271));
  jand g08204(.dina(n8022), .dinb(n1612), .dout(n8272));
  jand g08205(.dina(n8268), .dinb(n1620), .dout(n8273));
  jor  g08206(.dina(n8273), .dinb(n8272), .dout(n8274));
  jand g08207(.dina(n7692), .dinb(n1644), .dout(n8275));
  jor  g08208(.dina(n8275), .dinb(n8274), .dout(n8276));
  jor  g08209(.dina(n8276), .dinb(n8271), .dout(n8277));
  jxor g08210(.dina(n8277), .dinb(n65), .dout(n8278));
  jxor g08211(.dina(n8278), .dinb(n8048), .dout(n8279));
  jxor g08212(.dina(n8279), .dinb(n8040), .dout(n8280));
  jnot g08213(.din(n8280), .dout(n8281));
  jand g08214(.dina(n8250), .dinb(n8242), .dout(n8282));
  jand g08215(.dina(n8251), .dinb(n8064), .dout(n8283));
  jor  g08216(.dina(n8283), .dinb(n8282), .dout(n8284));
  jor  g08217(.dina(n7682), .dinb(n5281), .dout(n8285));
  jor  g08218(.dina(n7301), .dinb(n5532), .dout(n8286));
  jor  g08219(.dina(n6489), .dinb(n5537), .dout(n8287));
  jor  g08220(.dina(n7680), .dinb(n5539), .dout(n8288));
  jand g08221(.dina(n8288), .dinb(n8287), .dout(n8289));
  jand g08222(.dina(n8289), .dinb(n8286), .dout(n8290));
  jand g08223(.dina(n8290), .dinb(n8285), .dout(n8291));
  jxor g08224(.dina(n8291), .dinb(n5277), .dout(n8292));
  jnot g08225(.din(n8292), .dout(n8293));
  jand g08226(.dina(n8258), .dinb(n7680), .dout(n8294));
  jor  g08227(.dina(n8294), .dinb(n7999), .dout(n8295));
  jor  g08228(.dina(n8295), .dinb(n6496), .dout(n8296));
  jor  g08229(.dina(n8296), .dinb(\a[2] ), .dout(n8297));
  jand g08230(.dina(n8257), .dinb(n6495), .dout(n8298));
  jand g08231(.dina(n8000), .dinb(n6499), .dout(n8299));
  jor  g08232(.dina(n8299), .dinb(n6219), .dout(n8300));
  jor  g08233(.dina(n8300), .dinb(n8298), .dout(n8301));
  jand g08234(.dina(n8301), .dinb(n8297), .dout(n8302));
  jxor g08235(.dina(n8302), .dinb(n8293), .dout(n8303));
  jand g08236(.dina(n8240), .dinb(n8232), .dout(n8304));
  jand g08237(.dina(n8241), .dinb(n8067), .dout(n8305));
  jor  g08238(.dina(n8305), .dinb(n8304), .dout(n8306));
  jor  g08239(.dina(n8230), .dinb(n8222), .dout(n8307));
  jnot g08240(.din(n8307), .dout(n8308));
  jand g08241(.dina(n8231), .dinb(n8070), .dout(n8309));
  jor  g08242(.dina(n8309), .dinb(n8308), .dout(n8310));
  jor  g08243(.dina(n8220), .dinb(n8212), .dout(n8311));
  jnot g08244(.din(n8311), .dout(n8312));
  jnot g08245(.din(n8074), .dout(n8313));
  jand g08246(.dina(n8221), .dinb(n8313), .dout(n8314));
  jor  g08247(.dina(n8314), .dinb(n8312), .dout(n8315));
  jand g08248(.dina(n8210), .dinb(n8202), .dout(n8316));
  jnot g08249(.din(n8316), .dout(n8317));
  jnot g08250(.din(n8211), .dout(n8318));
  jor  g08251(.dina(n8318), .dinb(n8078), .dout(n8319));
  jand g08252(.dina(n8319), .dinb(n8317), .dout(n8320));
  jand g08253(.dina(n8200), .dinb(n8192), .dout(n8321));
  jand g08254(.dina(n8201), .dinb(n8083), .dout(n8322));
  jor  g08255(.dina(n8322), .dinb(n8321), .dout(n8323));
  jor  g08256(.dina(n8190), .dinb(n8182), .dout(n8324));
  jand g08257(.dina(n8191), .dinb(n8088), .dout(n8325));
  jnot g08258(.din(n8325), .dout(n8326));
  jand g08259(.dina(n8326), .dinb(n8324), .dout(n8327));
  jnot g08260(.din(n8327), .dout(n8328));
  jor  g08261(.dina(n8179), .dinb(n8171), .dout(n8329));
  jand g08262(.dina(n8180), .dinb(n8091), .dout(n8330));
  jnot g08263(.din(n8330), .dout(n8331));
  jand g08264(.dina(n8331), .dinb(n8329), .dout(n8332));
  jnot g08265(.din(n8332), .dout(n8333));
  jand g08266(.dina(n8168), .dinb(n8160), .dout(n8334));
  jand g08267(.dina(n8169), .dinb(n8094), .dout(n8335));
  jor  g08268(.dina(n8335), .dinb(n8334), .dout(n8336));
  jor  g08269(.dina(n8158), .dinb(n8150), .dout(n8337));
  jand g08270(.dina(n8159), .dinb(n8099), .dout(n8338));
  jnot g08271(.din(n8338), .dout(n8339));
  jand g08272(.dina(n8339), .dinb(n8337), .dout(n8340));
  jnot g08273(.din(n8340), .dout(n8341));
  jand g08274(.dina(n5395), .dinb(n1040), .dout(n8342));
  jand g08275(.dina(n8342), .dinb(n1016), .dout(n8343));
  jand g08276(.dina(n826), .dinb(n100), .dout(n8344));
  jand g08277(.dina(n8344), .dinb(n553), .dout(n8345));
  jand g08278(.dina(n8345), .dinb(n8343), .dout(n8346));
  jand g08279(.dina(n1827), .dinb(n431), .dout(n8347));
  jand g08280(.dina(n4585), .dinb(n2390), .dout(n8348));
  jand g08281(.dina(n8348), .dinb(n8347), .dout(n8349));
  jand g08282(.dina(n8349), .dinb(n3217), .dout(n8350));
  jand g08283(.dina(n8350), .dinb(n8346), .dout(n8351));
  jand g08284(.dina(n4678), .dinb(n1358), .dout(n8352));
  jand g08285(.dina(n8352), .dinb(n2077), .dout(n8353));
  jand g08286(.dina(n993), .dinb(n2148), .dout(n8354));
  jand g08287(.dina(n8354), .dinb(n7226), .dout(n8355));
  jand g08288(.dina(n8355), .dinb(n3392), .dout(n8356));
  jand g08289(.dina(n8356), .dinb(n8353), .dout(n8357));
  jand g08290(.dina(n8357), .dinb(n8351), .dout(n8358));
  jand g08291(.dina(n1867), .dinb(n1305), .dout(n8359));
  jand g08292(.dina(n8359), .dinb(n4644), .dout(n8360));
  jand g08293(.dina(n8360), .dinb(n4418), .dout(n8361));
  jand g08294(.dina(n2124), .dinb(n1682), .dout(n8362));
  jand g08295(.dina(n8362), .dinb(n2106), .dout(n8363));
  jand g08296(.dina(n8363), .dinb(n8361), .dout(n8364));
  jand g08297(.dina(n8364), .dinb(n8116), .dout(n8365));
  jand g08298(.dina(n2483), .dinb(n954), .dout(n8366));
  jand g08299(.dina(n933), .dinb(n178), .dout(n8367));
  jand g08300(.dina(n8367), .dinb(n1915), .dout(n8368));
  jand g08301(.dina(n8368), .dinb(n8366), .dout(n8369));
  jand g08302(.dina(n2023), .dinb(n881), .dout(n8370));
  jand g08303(.dina(n8370), .dinb(n662), .dout(n8371));
  jand g08304(.dina(n3819), .dinb(n1205), .dout(n8372));
  jand g08305(.dina(n8372), .dinb(n8371), .dout(n8373));
  jand g08306(.dina(n8373), .dinb(n8369), .dout(n8374));
  jand g08307(.dina(n8374), .dinb(n5351), .dout(n8375));
  jand g08308(.dina(n8375), .dinb(n3024), .dout(n8376));
  jand g08309(.dina(n8376), .dinb(n8365), .dout(n8377));
  jand g08310(.dina(n1189), .dinb(n495), .dout(n8378));
  jand g08311(.dina(n445), .dinb(n463), .dout(n8379));
  jand g08312(.dina(n8379), .dinb(n8378), .dout(n8380));
  jand g08313(.dina(n641), .dinb(n880), .dout(n8381));
  jand g08314(.dina(n8381), .dinb(n1247), .dout(n8382));
  jand g08315(.dina(n8382), .dinb(n8380), .dout(n8383));
  jand g08316(.dina(n452), .dinb(n1283), .dout(n8384));
  jand g08317(.dina(n4422), .dinb(n1536), .dout(n8385));
  jand g08318(.dina(n8385), .dinb(n8384), .dout(n8386));
  jand g08319(.dina(n8386), .dinb(n3150), .dout(n8387));
  jand g08320(.dina(n8387), .dinb(n8383), .dout(n8388));
  jand g08321(.dina(n1714), .dinb(n1976), .dout(n8389));
  jand g08322(.dina(n8389), .dinb(n4668), .dout(n8390));
  jand g08323(.dina(n8390), .dinb(n1959), .dout(n8391));
  jand g08324(.dina(n1225), .dinb(n1429), .dout(n8392));
  jand g08325(.dina(n718), .dinb(n92), .dout(n8393));
  jand g08326(.dina(n8393), .dinb(n8392), .dout(n8394));
  jand g08327(.dina(n5180), .dinb(n583), .dout(n8395));
  jand g08328(.dina(n8395), .dinb(n8394), .dout(n8396));
  jand g08329(.dina(n8396), .dinb(n3765), .dout(n8397));
  jand g08330(.dina(n8397), .dinb(n8391), .dout(n8398));
  jand g08331(.dina(n8398), .dinb(n8388), .dout(n8399));
  jand g08332(.dina(n1541), .dinb(n510), .dout(n8400));
  jand g08333(.dina(n8400), .dinb(n588), .dout(n8401));
  jand g08334(.dina(n8401), .dinb(n5304), .dout(n8402));
  jand g08335(.dina(n503), .dinb(n831), .dout(n8403));
  jand g08336(.dina(n8403), .dinb(n714), .dout(n8404));
  jand g08337(.dina(n1345), .dinb(n493), .dout(n8405));
  jand g08338(.dina(n8405), .dinb(n2165), .dout(n8406));
  jand g08339(.dina(n8406), .dinb(n8404), .dout(n8407));
  jand g08340(.dina(n5515), .dinb(n1495), .dout(n8408));
  jand g08341(.dina(n8408), .dinb(n2587), .dout(n8409));
  jand g08342(.dina(n8409), .dinb(n8407), .dout(n8410));
  jand g08343(.dina(n8410), .dinb(n8402), .dout(n8411));
  jand g08344(.dina(n8411), .dinb(n8399), .dout(n8412));
  jand g08345(.dina(n8412), .dinb(n8377), .dout(n8413));
  jand g08346(.dina(n8413), .dinb(n8358), .dout(n8414));
  jor  g08347(.dina(n7061), .dinb(n2197), .dout(n8415));
  jand g08348(.dina(n6050), .dinb(n2061), .dout(n8416));
  jand g08349(.dina(n5084), .dinb(n1955), .dout(n8417));
  jor  g08350(.dina(n8417), .dinb(n8416), .dout(n8418));
  jand g08351(.dina(n5082), .dinb(n2058), .dout(n8419));
  jor  g08352(.dina(n8419), .dinb(n8418), .dout(n8420));
  jnot g08353(.din(n8420), .dout(n8421));
  jand g08354(.dina(n8421), .dinb(n8415), .dout(n8422));
  jxor g08355(.dina(n8422), .dinb(n8414), .dout(n8423));
  jxor g08356(.dina(n8423), .dinb(n8341), .dout(n8424));
  jnot g08357(.din(n8424), .dout(n8425));
  jor  g08358(.dina(n4343), .dinb(n2779), .dout(n8426));
  jor  g08359(.dina(n4346), .dinb(n2428), .dout(n8427));
  jor  g08360(.dina(n4348), .dinb(n2629), .dout(n8428));
  jand g08361(.dina(n8428), .dinb(n8427), .dout(n8429));
  jor  g08362(.dina(n3683), .dinb(n2174), .dout(n8430));
  jand g08363(.dina(n8430), .dinb(n8429), .dout(n8431));
  jand g08364(.dina(n8431), .dinb(n8426), .dout(n8432));
  jxor g08365(.dina(n8432), .dinb(\a[29] ), .dout(n8433));
  jxor g08366(.dina(n8433), .dinb(n8425), .dout(n8434));
  jxor g08367(.dina(n8434), .dinb(n8336), .dout(n8435));
  jnot g08368(.din(n8435), .dout(n8436));
  jor  g08369(.dina(n3081), .dinb(n2303), .dout(n8437));
  jor  g08370(.dina(n2553), .dinb(n1805), .dout(n8438));
  jor  g08371(.dina(n2738), .dinb(n2306), .dout(n8439));
  jand g08372(.dina(n8439), .dinb(n8438), .dout(n8440));
  jor  g08373(.dina(n3072), .dinb(n2309), .dout(n8441));
  jand g08374(.dina(n8441), .dinb(n8440), .dout(n8442));
  jand g08375(.dina(n8442), .dinb(n8437), .dout(n8443));
  jxor g08376(.dina(n8443), .dinb(\a[26] ), .dout(n8444));
  jxor g08377(.dina(n8444), .dinb(n8436), .dout(n8445));
  jxor g08378(.dina(n8445), .dinb(n8333), .dout(n8446));
  jnot g08379(.din(n8446), .dout(n8447));
  jor  g08380(.dina(n3203), .dinb(n1617), .dout(n8448));
  jor  g08381(.dina(n3422), .dinb(n807), .dout(n8449));
  jor  g08382(.dina(n3420), .dinb(n1621), .dout(n8450));
  jor  g08383(.dina(n3286), .dinb(n1613), .dout(n8451));
  jand g08384(.dina(n8451), .dinb(n8450), .dout(n8452));
  jand g08385(.dina(n8452), .dinb(n8449), .dout(n8453));
  jand g08386(.dina(n8453), .dinb(n8448), .dout(n8454));
  jxor g08387(.dina(n8454), .dinb(\a[23] ), .dout(n8455));
  jxor g08388(.dina(n8455), .dinb(n8447), .dout(n8456));
  jxor g08389(.dina(n8456), .dinb(n8328), .dout(n8457));
  jnot g08390(.din(n8457), .dout(n8458));
  jor  g08391(.dina(n4038), .dinb(n1820), .dout(n8459));
  jor  g08392(.dina(n3863), .dinb(n2181), .dout(n8460));
  jor  g08393(.dina(n3929), .dinb(n2189), .dout(n8461));
  jand g08394(.dina(n8461), .dinb(n8460), .dout(n8462));
  jor  g08395(.dina(n3787), .dinb(n2186), .dout(n8463));
  jand g08396(.dina(n8463), .dinb(n8462), .dout(n8464));
  jand g08397(.dina(n8464), .dinb(n8459), .dout(n8465));
  jxor g08398(.dina(n8465), .dinb(\a[20] ), .dout(n8466));
  jxor g08399(.dina(n8466), .dinb(n8458), .dout(n8467));
  jxor g08400(.dina(n8467), .dinb(n8323), .dout(n8468));
  jor  g08401(.dina(n4726), .dinb(n2744), .dout(n8469));
  jor  g08402(.dina(n4471), .dinb(n2749), .dout(n8470));
  jor  g08403(.dina(n4596), .dinb(n2753), .dout(n8471));
  jor  g08404(.dina(n4019), .dinb(n2758), .dout(n8472));
  jand g08405(.dina(n8472), .dinb(n8471), .dout(n8473));
  jand g08406(.dina(n8473), .dinb(n8470), .dout(n8474));
  jand g08407(.dina(n8474), .dinb(n8469), .dout(n8475));
  jxor g08408(.dina(n8475), .dinb(n2441), .dout(n8476));
  jxor g08409(.dina(n8476), .dinb(n8468), .dout(n8477));
  jxor g08410(.dina(n8477), .dinb(n8320), .dout(n8478));
  jor  g08411(.dina(n5266), .dinb(n3424), .dout(n8479));
  jor  g08412(.dina(n4686), .dinb(n3429), .dout(n8480));
  jor  g08413(.dina(n5264), .dinb(n3426), .dout(n8481));
  jand g08414(.dina(n8481), .dinb(n8480), .dout(n8482));
  jor  g08415(.dina(n4526), .dinb(n3211), .dout(n8483));
  jand g08416(.dina(n8483), .dinb(n8482), .dout(n8484));
  jand g08417(.dina(n8484), .dinb(n8479), .dout(n8485));
  jxor g08418(.dina(n8485), .dinb(\a[14] ), .dout(n8486));
  jxor g08419(.dina(n8486), .dinb(n8478), .dout(n8487));
  jxor g08420(.dina(n8487), .dinb(n8315), .dout(n8488));
  jor  g08421(.dina(n5527), .dinb(n4023), .dout(n8489));
  jor  g08422(.dina(n5364), .dinb(n4028), .dout(n8490));
  jor  g08423(.dina(n5422), .dinb(n3871), .dout(n8491));
  jor  g08424(.dina(n5525), .dinb(n4025), .dout(n8492));
  jand g08425(.dina(n8492), .dinb(n8491), .dout(n8493));
  jand g08426(.dina(n8493), .dinb(n8490), .dout(n8494));
  jand g08427(.dina(n8494), .dinb(n8489), .dout(n8495));
  jxor g08428(.dina(n8495), .dinb(n4050), .dout(n8496));
  jxor g08429(.dina(n8496), .dinb(n8488), .dout(n8497));
  jxor g08430(.dina(n8497), .dinb(n8310), .dout(n8498));
  jor  g08431(.dina(n6999), .dinb(n4692), .dout(n8499));
  jor  g08432(.dina(n6390), .dinb(n4697), .dout(n8500));
  jor  g08433(.dina(n6205), .dinb(n4702), .dout(n8501));
  jor  g08434(.dina(n6297), .dinb(n4705), .dout(n8502));
  jand g08435(.dina(n8502), .dinb(n8501), .dout(n8503));
  jand g08436(.dina(n8503), .dinb(n8500), .dout(n8504));
  jand g08437(.dina(n8504), .dinb(n8499), .dout(n8505));
  jxor g08438(.dina(n8505), .dinb(n4713), .dout(n8506));
  jxor g08439(.dina(n8506), .dinb(n8498), .dout(n8507));
  jxor g08440(.dina(n8507), .dinb(n8306), .dout(n8508));
  jxor g08441(.dina(n8508), .dinb(n8303), .dout(n8509));
  jand g08442(.dina(n8509), .dinb(n8284), .dout(n8510));
  jxor g08443(.dina(n8509), .dinb(n8284), .dout(n8511));
  jxor g08444(.dina(n8251), .dinb(n8064), .dout(n8512));
  jxor g08445(.dina(n8265), .dinb(n6219), .dout(n8513));
  jand g08446(.dina(n8513), .dinb(n8512), .dout(n8514));
  jand g08447(.dina(n8267), .dinb(n8061), .dout(n8515));
  jor  g08448(.dina(n8515), .dinb(n8514), .dout(n8516));
  jand g08449(.dina(n8516), .dinb(n8511), .dout(n8517));
  jor  g08450(.dina(n8517), .dinb(n8510), .dout(n8518));
  jor  g08451(.dina(n8302), .dinb(n8293), .dout(n8519));
  jnot g08452(.din(n8519), .dout(n8520));
  jand g08453(.dina(n8508), .dinb(n8303), .dout(n8521));
  jor  g08454(.dina(n8521), .dinb(n8520), .dout(n8522));
  jand g08455(.dina(n8506), .dinb(n8498), .dout(n8523));
  jnot g08456(.din(n8523), .dout(n8524));
  jnot g08457(.din(n8306), .dout(n8525));
  jnot g08458(.din(n8507), .dout(n8526));
  jor  g08459(.dina(n8526), .dinb(n8525), .dout(n8527));
  jand g08460(.dina(n8527), .dinb(n8524), .dout(n8528));
  jand g08461(.dina(n8496), .dinb(n8488), .dout(n8529));
  jnot g08462(.din(n8529), .dout(n8530));
  jnot g08463(.din(n8310), .dout(n8531));
  jnot g08464(.din(n8497), .dout(n8532));
  jor  g08465(.dina(n8532), .dinb(n8531), .dout(n8533));
  jand g08466(.dina(n8533), .dinb(n8530), .dout(n8534));
  jor  g08467(.dina(n8486), .dinb(n8478), .dout(n8535));
  jnot g08468(.din(n8535), .dout(n8536));
  jand g08469(.dina(n8487), .dinb(n8315), .dout(n8537));
  jor  g08470(.dina(n8537), .dinb(n8536), .dout(n8538));
  jand g08471(.dina(n8476), .dinb(n8468), .dout(n8539));
  jnot g08472(.din(n8320), .dout(n8540));
  jand g08473(.dina(n8477), .dinb(n8540), .dout(n8541));
  jor  g08474(.dina(n8541), .dinb(n8539), .dout(n8542));
  jor  g08475(.dina(n8466), .dinb(n8458), .dout(n8543));
  jand g08476(.dina(n8467), .dinb(n8323), .dout(n8544));
  jnot g08477(.din(n8544), .dout(n8545));
  jand g08478(.dina(n8545), .dinb(n8543), .dout(n8546));
  jnot g08479(.din(n8546), .dout(n8547));
  jor  g08480(.dina(n8455), .dinb(n8447), .dout(n8548));
  jand g08481(.dina(n8456), .dinb(n8328), .dout(n8549));
  jnot g08482(.din(n8549), .dout(n8550));
  jand g08483(.dina(n8550), .dinb(n8548), .dout(n8551));
  jnot g08484(.din(n8551), .dout(n8552));
  jor  g08485(.dina(n8444), .dinb(n8436), .dout(n8553));
  jand g08486(.dina(n8445), .dinb(n8333), .dout(n8554));
  jnot g08487(.din(n8554), .dout(n8555));
  jand g08488(.dina(n8555), .dinb(n8553), .dout(n8556));
  jnot g08489(.din(n8556), .dout(n8557));
  jor  g08490(.dina(n8433), .dinb(n8425), .dout(n8558));
  jand g08491(.dina(n8434), .dinb(n8336), .dout(n8559));
  jnot g08492(.din(n8559), .dout(n8560));
  jand g08493(.dina(n8560), .dinb(n8558), .dout(n8561));
  jnot g08494(.din(n8561), .dout(n8562));
  jor  g08495(.dina(n8422), .dinb(n8414), .dout(n8563));
  jand g08496(.dina(n8423), .dinb(n8341), .dout(n8564));
  jnot g08497(.din(n8564), .dout(n8565));
  jand g08498(.dina(n8565), .dinb(n8563), .dout(n8566));
  jnot g08499(.din(n8566), .dout(n8567));
  jor  g08500(.dina(n7061), .dinb(n2176), .dout(n8568));
  jand g08501(.dina(n5082), .dinb(n1955), .dout(n8569));
  jand g08502(.dina(n6050), .dinb(n2058), .dout(n8570));
  jor  g08503(.dina(n8570), .dinb(n8569), .dout(n8571));
  jand g08504(.dina(n5084), .dinb(n2325), .dout(n8572));
  jor  g08505(.dina(n8572), .dinb(n8571), .dout(n8573));
  jnot g08506(.din(n8573), .dout(n8574));
  jand g08507(.dina(n8574), .dinb(n8568), .dout(n8575));
  jnot g08508(.din(n8575), .dout(n8576));
  jnot g08509(.din(n855), .dout(n8577));
  jand g08510(.dina(n3217), .dinb(n8577), .dout(n8578));
  jand g08511(.dina(n7512), .dinb(n1527), .dout(n8579));
  jand g08512(.dina(n1524), .dinb(n1449), .dout(n8580));
  jand g08513(.dina(n8580), .dinb(n8579), .dout(n8581));
  jand g08514(.dina(n8581), .dinb(n8578), .dout(n8582));
  jand g08515(.dina(n1378), .dinb(n699), .dout(n8583));
  jand g08516(.dina(n325), .dinb(n1203), .dout(n8584));
  jand g08517(.dina(n8584), .dinb(n8583), .dout(n8585));
  jand g08518(.dina(n8585), .dinb(n8582), .dout(n8586));
  jand g08519(.dina(n8586), .dinb(n3861), .dout(n8587));
  jand g08520(.dina(n694), .dinb(n1325), .dout(n8588));
  jand g08521(.dina(n1721), .dinb(n586), .dout(n8589));
  jand g08522(.dina(n8589), .dinb(n2077), .dout(n8590));
  jand g08523(.dina(n8590), .dinb(n2716), .dout(n8591));
  jand g08524(.dina(n8591), .dinb(n8588), .dout(n8592));
  jand g08525(.dina(n680), .dinb(n1476), .dout(n8593));
  jand g08526(.dina(n647), .dinb(n440), .dout(n8594));
  jand g08527(.dina(n8594), .dinb(n8593), .dout(n8595));
  jand g08528(.dina(n8595), .dinb(n511), .dout(n8596));
  jand g08529(.dina(n8596), .dinb(n2100), .dout(n8597));
  jand g08530(.dina(n8597), .dinb(n8592), .dout(n8598));
  jand g08531(.dina(n3322), .dinb(n2148), .dout(n8599));
  jand g08532(.dina(n8599), .dinb(n1772), .dout(n8600));
  jand g08533(.dina(n1731), .dinb(n100), .dout(n8601));
  jand g08534(.dina(n8601), .dinb(n1451), .dout(n8602));
  jand g08535(.dina(n1522), .dinb(n1317), .dout(n8603));
  jand g08536(.dina(n8603), .dinb(n1512), .dout(n8604));
  jand g08537(.dina(n8604), .dinb(n8602), .dout(n8605));
  jnot g08538(.din(n1032), .dout(n8606));
  jand g08539(.dina(n2701), .dinb(n8606), .dout(n8607));
  jand g08540(.dina(n8607), .dinb(n8605), .dout(n8608));
  jand g08541(.dina(n8608), .dinb(n8600), .dout(n8609));
  jand g08542(.dina(n8609), .dinb(n8598), .dout(n8610));
  jand g08543(.dina(n1352), .dinb(n92), .dout(n8611));
  jand g08544(.dina(n8611), .dinb(n2680), .dout(n8612));
  jand g08545(.dina(n826), .dinb(n908), .dout(n8613));
  jand g08546(.dina(n8613), .dinb(n1315), .dout(n8614));
  jand g08547(.dina(n8614), .dinb(n3261), .dout(n8615));
  jand g08548(.dina(n8615), .dinb(n8612), .dout(n8616));
  jand g08549(.dina(n1912), .dinb(n431), .dout(n8617));
  jand g08550(.dina(n670), .dinb(n1344), .dout(n8618));
  jand g08551(.dina(n8618), .dinb(n521), .dout(n8619));
  jand g08552(.dina(n1470), .dinb(n1238), .dout(n8620));
  jand g08553(.dina(n8620), .dinb(n2406), .dout(n8621));
  jand g08554(.dina(n8621), .dinb(n8619), .dout(n8622));
  jand g08555(.dina(n8622), .dinb(n8617), .dout(n8623));
  jand g08556(.dina(n8623), .dinb(n8616), .dout(n8624));
  jand g08557(.dina(n8624), .dinb(n8610), .dout(n8625));
  jand g08558(.dina(n8625), .dinb(n1298), .dout(n8626));
  jand g08559(.dina(n8626), .dinb(n8587), .dout(n8627));
  jxor g08560(.dina(n8627), .dinb(n6219), .dout(n8628));
  jxor g08561(.dina(n8628), .dinb(n8576), .dout(n8629));
  jxor g08562(.dina(n8629), .dinb(n8567), .dout(n8630));
  jor  g08563(.dina(n4343), .dinb(n2768), .dout(n8631));
  jor  g08564(.dina(n4348), .dinb(n2553), .dout(n8632));
  jor  g08565(.dina(n3683), .dinb(n2428), .dout(n8633));
  jor  g08566(.dina(n4346), .dinb(n2629), .dout(n8634));
  jand g08567(.dina(n8634), .dinb(n8633), .dout(n8635));
  jand g08568(.dina(n8635), .dinb(n8632), .dout(n8636));
  jand g08569(.dina(n8636), .dinb(n8631), .dout(n8637));
  jxor g08570(.dina(n8637), .dinb(n93), .dout(n8638));
  jxor g08571(.dina(n8638), .dinb(n8630), .dout(n8639));
  jxor g08572(.dina(n8639), .dinb(n8562), .dout(n8640));
  jor  g08573(.dina(n3451), .dinb(n2303), .dout(n8641));
  jor  g08574(.dina(n3072), .dinb(n2306), .dout(n8642));
  jor  g08575(.dina(n3203), .dinb(n2309), .dout(n8643));
  jor  g08576(.dina(n2738), .dinb(n1805), .dout(n8644));
  jand g08577(.dina(n8644), .dinb(n8643), .dout(n8645));
  jand g08578(.dina(n8645), .dinb(n8642), .dout(n8646));
  jand g08579(.dina(n8646), .dinb(n8641), .dout(n8647));
  jxor g08580(.dina(n8647), .dinb(n77), .dout(n8648));
  jxor g08581(.dina(n8648), .dinb(n8640), .dout(n8649));
  jxor g08582(.dina(n8649), .dinb(n8557), .dout(n8650));
  jnot g08583(.din(n8650), .dout(n8651));
  jor  g08584(.dina(n3789), .dinb(n807), .dout(n8652));
  jor  g08585(.dina(n3420), .dinb(n1613), .dout(n8653));
  jor  g08586(.dina(n3286), .dinb(n1617), .dout(n8654));
  jand g08587(.dina(n8654), .dinb(n8653), .dout(n8655));
  jor  g08588(.dina(n3787), .dinb(n1621), .dout(n8656));
  jand g08589(.dina(n8656), .dinb(n8655), .dout(n8657));
  jand g08590(.dina(n8657), .dinb(n8652), .dout(n8658));
  jxor g08591(.dina(n8658), .dinb(\a[23] ), .dout(n8659));
  jxor g08592(.dina(n8659), .dinb(n8651), .dout(n8660));
  jxor g08593(.dina(n8660), .dinb(n8552), .dout(n8661));
  jnot g08594(.din(n8661), .dout(n8662));
  jor  g08595(.dina(n3863), .dinb(n2186), .dout(n8663));
  jor  g08596(.dina(n4021), .dinb(n1820), .dout(n8664));
  jor  g08597(.dina(n4019), .dinb(n2189), .dout(n8665));
  jor  g08598(.dina(n3929), .dinb(n2181), .dout(n8666));
  jand g08599(.dina(n8666), .dinb(n8665), .dout(n8667));
  jand g08600(.dina(n8667), .dinb(n8664), .dout(n8668));
  jand g08601(.dina(n8668), .dinb(n8663), .dout(n8669));
  jxor g08602(.dina(n8669), .dinb(\a[20] ), .dout(n8670));
  jxor g08603(.dina(n8670), .dinb(n8662), .dout(n8671));
  jxor g08604(.dina(n8671), .dinb(n8547), .dout(n8672));
  jor  g08605(.dina(n4714), .dinb(n2744), .dout(n8673));
  jor  g08606(.dina(n4596), .dinb(n2749), .dout(n8674));
  jor  g08607(.dina(n4471), .dinb(n2758), .dout(n8675));
  jor  g08608(.dina(n4526), .dinb(n2753), .dout(n8676));
  jand g08609(.dina(n8676), .dinb(n8675), .dout(n8677));
  jand g08610(.dina(n8677), .dinb(n8674), .dout(n8678));
  jand g08611(.dina(n8678), .dinb(n8673), .dout(n8679));
  jxor g08612(.dina(n8679), .dinb(n2441), .dout(n8680));
  jxor g08613(.dina(n8680), .dinb(n8672), .dout(n8681));
  jxor g08614(.dina(n8681), .dinb(n8542), .dout(n8682));
  jor  g08615(.dina(n5560), .dinb(n3424), .dout(n8683));
  jor  g08616(.dina(n5264), .dinb(n3429), .dout(n8684));
  jor  g08617(.dina(n4686), .dinb(n3211), .dout(n8685));
  jor  g08618(.dina(n5422), .dinb(n3426), .dout(n8686));
  jand g08619(.dina(n8686), .dinb(n8685), .dout(n8687));
  jand g08620(.dina(n8687), .dinb(n8684), .dout(n8688));
  jand g08621(.dina(n8688), .dinb(n8683), .dout(n8689));
  jxor g08622(.dina(n8689), .dinb(n3473), .dout(n8690));
  jxor g08623(.dina(n8690), .dinb(n8682), .dout(n8691));
  jxor g08624(.dina(n8691), .dinb(n8538), .dout(n8692));
  jor  g08625(.dina(n6207), .dinb(n4023), .dout(n8693));
  jor  g08626(.dina(n5525), .dinb(n4028), .dout(n8694));
  jor  g08627(.dina(n5364), .dinb(n3871), .dout(n8695));
  jor  g08628(.dina(n6205), .dinb(n4025), .dout(n8696));
  jand g08629(.dina(n8696), .dinb(n8695), .dout(n8697));
  jand g08630(.dina(n8697), .dinb(n8694), .dout(n8698));
  jand g08631(.dina(n8698), .dinb(n8693), .dout(n8699));
  jxor g08632(.dina(n8699), .dinb(n4050), .dout(n8700));
  jxor g08633(.dina(n8700), .dinb(n8692), .dout(n8701));
  jxor g08634(.dina(n8701), .dinb(n8534), .dout(n8702));
  jor  g08635(.dina(n6491), .dinb(n4692), .dout(n8703));
  jor  g08636(.dina(n6297), .dinb(n4697), .dout(n8704));
  jor  g08637(.dina(n6489), .dinb(n4705), .dout(n8705));
  jand g08638(.dina(n8705), .dinb(n8704), .dout(n8706));
  jor  g08639(.dina(n6390), .dinb(n4702), .dout(n8707));
  jand g08640(.dina(n8707), .dinb(n8706), .dout(n8708));
  jand g08641(.dina(n8708), .dinb(n8703), .dout(n8709));
  jxor g08642(.dina(n8709), .dinb(\a[8] ), .dout(n8710));
  jxor g08643(.dina(n8710), .dinb(n8702), .dout(n8711));
  jxor g08644(.dina(n8711), .dinb(n8528), .dout(n8712));
  jor  g08645(.dina(n7301), .dinb(n5537), .dout(n8713));
  jor  g08646(.dina(n8002), .dinb(n5281), .dout(n8714));
  jor  g08647(.dina(n7999), .dinb(n5539), .dout(n8715));
  jor  g08648(.dina(n7680), .dinb(n5532), .dout(n8716));
  jand g08649(.dina(n8716), .dinb(n8715), .dout(n8717));
  jand g08650(.dina(n8717), .dinb(n8714), .dout(n8718));
  jand g08651(.dina(n8718), .dinb(n8713), .dout(n8719));
  jxor g08652(.dina(n8719), .dinb(\a[5] ), .dout(n8720));
  jxor g08653(.dina(n8720), .dinb(n8712), .dout(n8721));
  jxor g08654(.dina(n8721), .dinb(n8522), .dout(n8722));
  jxor g08655(.dina(n8722), .dinb(n8518), .dout(n8723));
  jnot g08656(.din(n8284), .dout(n8724));
  jxor g08657(.dina(n8509), .dinb(n8724), .dout(n8725));
  jor  g08658(.dina(n8266), .dinb(n8253), .dout(n8726));
  jor  g08659(.dina(n8020), .dinb(n7934), .dout(n8727));
  jor  g08660(.dina(n7312), .dinb(n7028), .dout(n8728));
  jand g08661(.dina(n8728), .dinb(n7330), .dout(n8729));
  jxor g08662(.dina(n7627), .dinb(n7713), .dout(n8730));
  jxor g08663(.dina(n7690), .dinb(n8730), .dout(n8731));
  jor  g08664(.dina(n8731), .dinb(n8729), .dout(n8732));
  jand g08665(.dina(n8732), .dinb(n7707), .dout(n8733));
  jxor g08666(.dina(n8020), .dinb(n8054), .dout(n8734));
  jor  g08667(.dina(n8734), .dinb(n8733), .dout(n8735));
  jand g08668(.dina(n8735), .dinb(n8727), .dout(n8736));
  jxor g08669(.dina(n8266), .dinb(n8512), .dout(n8737));
  jor  g08670(.dina(n8737), .dinb(n8736), .dout(n8738));
  jand g08671(.dina(n8738), .dinb(n8726), .dout(n8739));
  jxor g08672(.dina(n8739), .dinb(n8725), .dout(n8740));
  jand g08673(.dina(n8740), .dinb(n8723), .dout(n8741));
  jand g08674(.dina(n8740), .dinb(n8268), .dout(n8742));
  jand g08675(.dina(n8268), .dinb(n8022), .dout(n8743));
  jand g08676(.dina(n8269), .dinb(n8051), .dout(n8744));
  jor  g08677(.dina(n8744), .dinb(n8743), .dout(n8745));
  jxor g08678(.dina(n8740), .dinb(n8268), .dout(n8746));
  jand g08679(.dina(n8746), .dinb(n8745), .dout(n8747));
  jor  g08680(.dina(n8747), .dinb(n8742), .dout(n8748));
  jxor g08681(.dina(n8740), .dinb(n8723), .dout(n8749));
  jand g08682(.dina(n8749), .dinb(n8748), .dout(n8750));
  jor  g08683(.dina(n8750), .dinb(n8741), .dout(n8751));
  jand g08684(.dina(n8721), .dinb(n8522), .dout(n8752));
  jand g08685(.dina(n8722), .dinb(n8518), .dout(n8753));
  jor  g08686(.dina(n8753), .dinb(n8752), .dout(n8754));
  jnot g08687(.din(n8528), .dout(n8755));
  jand g08688(.dina(n8711), .dinb(n8755), .dout(n8756));
  jor  g08689(.dina(n8720), .dinb(n8712), .dout(n8757));
  jnot g08690(.din(n8757), .dout(n8758));
  jor  g08691(.dina(n8758), .dinb(n8756), .dout(n8759));
  jnot g08692(.din(n8534), .dout(n8760));
  jand g08693(.dina(n8701), .dinb(n8760), .dout(n8761));
  jnot g08694(.din(n8761), .dout(n8762));
  jor  g08695(.dina(n8710), .dinb(n8702), .dout(n8763));
  jand g08696(.dina(n8763), .dinb(n8762), .dout(n8764));
  jor  g08697(.dina(n7999), .dinb(n5532), .dout(n8765));
  jor  g08698(.dina(n8260), .dinb(n5281), .dout(n8766));
  jor  g08699(.dina(n7680), .dinb(n5537), .dout(n8767));
  jand g08700(.dina(n8767), .dinb(n8766), .dout(n8768));
  jand g08701(.dina(n8768), .dinb(n8765), .dout(n8769));
  jxor g08702(.dina(n8769), .dinb(\a[5] ), .dout(n8770));
  jxor g08703(.dina(n8770), .dinb(n8764), .dout(n8771));
  jand g08704(.dina(n8691), .dinb(n8538), .dout(n8772));
  jand g08705(.dina(n8700), .dinb(n8692), .dout(n8773));
  jor  g08706(.dina(n8773), .dinb(n8772), .dout(n8774));
  jand g08707(.dina(n8681), .dinb(n8542), .dout(n8775));
  jand g08708(.dina(n8690), .dinb(n8682), .dout(n8776));
  jor  g08709(.dina(n8776), .dinb(n8775), .dout(n8777));
  jand g08710(.dina(n8671), .dinb(n8547), .dout(n8778));
  jand g08711(.dina(n8680), .dinb(n8672), .dout(n8779));
  jor  g08712(.dina(n8779), .dinb(n8778), .dout(n8780));
  jand g08713(.dina(n8660), .dinb(n8552), .dout(n8781));
  jnot g08714(.din(n8781), .dout(n8782));
  jor  g08715(.dina(n8670), .dinb(n8662), .dout(n8783));
  jand g08716(.dina(n8783), .dinb(n8782), .dout(n8784));
  jnot g08717(.din(n8784), .dout(n8785));
  jand g08718(.dina(n8649), .dinb(n8557), .dout(n8786));
  jnot g08719(.din(n8786), .dout(n8787));
  jor  g08720(.dina(n8659), .dinb(n8651), .dout(n8788));
  jand g08721(.dina(n8788), .dinb(n8787), .dout(n8789));
  jnot g08722(.din(n8789), .dout(n8790));
  jand g08723(.dina(n8639), .dinb(n8562), .dout(n8791));
  jand g08724(.dina(n8648), .dinb(n8640), .dout(n8792));
  jor  g08725(.dina(n8792), .dinb(n8791), .dout(n8793));
  jand g08726(.dina(n8629), .dinb(n8567), .dout(n8794));
  jand g08727(.dina(n8638), .dinb(n8630), .dout(n8795));
  jor  g08728(.dina(n8795), .dinb(n8794), .dout(n8796));
  jor  g08729(.dina(n7061), .dinb(n2430), .dout(n8797));
  jand g08730(.dina(n6050), .dinb(n1955), .dout(n8798));
  jand g08731(.dina(n5084), .dinb(n2633), .dout(n8799));
  jor  g08732(.dina(n8799), .dinb(n8798), .dout(n8800));
  jand g08733(.dina(n5082), .dinb(n2325), .dout(n8801));
  jor  g08734(.dina(n8801), .dinb(n8800), .dout(n8802));
  jnot g08735(.din(n8802), .dout(n8803));
  jand g08736(.dina(n8803), .dinb(n8797), .dout(n8804));
  jnot g08737(.din(n8804), .dout(n8805));
  jor  g08738(.dina(n8627), .dinb(n6219), .dout(n8806));
  jand g08739(.dina(n8628), .dinb(n8576), .dout(n8807));
  jnot g08740(.din(n8807), .dout(n8808));
  jand g08741(.dina(n8808), .dinb(n8806), .dout(n8809));
  jnot g08742(.din(n8809), .dout(n8810));
  jand g08743(.dina(n5375), .dinb(n503), .dout(n8811));
  jand g08744(.dina(n8811), .dinb(n838), .dout(n8812));
  jand g08745(.dina(n1772), .dinb(n440), .dout(n8813));
  jand g08746(.dina(n8813), .dinb(n7512), .dout(n8814));
  jand g08747(.dina(n8814), .dinb(n8812), .dout(n8815));
  jand g08748(.dina(n2587), .dinb(n882), .dout(n8816));
  jand g08749(.dina(n8816), .dinb(n931), .dout(n8817));
  jand g08750(.dina(n8817), .dinb(n2152), .dout(n8818));
  jand g08751(.dina(n8818), .dinb(n8815), .dout(n8819));
  jand g08752(.dina(n700), .dinb(n511), .dout(n8820));
  jand g08753(.dina(n4675), .dinb(n1834), .dout(n8821));
  jand g08754(.dina(n8821), .dinb(n8820), .dout(n8822));
  jand g08755(.dina(n8822), .dinb(n2077), .dout(n8823));
  jand g08756(.dina(n8823), .dinb(n8819), .dout(n8824));
  jand g08757(.dina(n650), .dinb(n929), .dout(n8825));
  jand g08758(.dina(n8825), .dinb(n7983), .dout(n8826));
  jand g08759(.dina(n951), .dinb(n639), .dout(n8827));
  jand g08760(.dina(n811), .dinb(n130), .dout(n8828));
  jand g08761(.dina(n8828), .dinb(n3238), .dout(n8829));
  jand g08762(.dina(n8829), .dinb(n8827), .dout(n8830));
  jand g08763(.dina(n680), .dinb(n1334), .dout(n8831));
  jand g08764(.dina(n8831), .dinb(n964), .dout(n8832));
  jand g08765(.dina(n8832), .dinb(n8830), .dout(n8833));
  jand g08766(.dina(n8833), .dinb(n8826), .dout(n8834));
  jand g08767(.dina(n8362), .dinb(n965), .dout(n8835));
  jand g08768(.dina(n1511), .dinb(n619), .dout(n8836));
  jand g08769(.dina(n8836), .dinb(n1768), .dout(n8837));
  jand g08770(.dina(n8837), .dinb(n329), .dout(n8838));
  jand g08771(.dina(n8838), .dinb(n8835), .dout(n8839));
  jand g08772(.dina(n8839), .dinb(n5329), .dout(n8840));
  jand g08773(.dina(n8840), .dinb(n8834), .dout(n8841));
  jand g08774(.dina(n8841), .dinb(n8824), .dout(n8842));
  jand g08775(.dina(n1378), .dinb(n662), .dout(n8843));
  jand g08776(.dina(n8843), .dinb(n5401), .dout(n8844));
  jand g08777(.dina(n8844), .dinb(n8842), .dout(n8845));
  jand g08778(.dina(n8845), .dinb(n1202), .dout(n8846));
  jxor g08779(.dina(n8846), .dinb(n6219), .dout(n8847));
  jxor g08780(.dina(n8847), .dinb(n8810), .dout(n8848));
  jxor g08781(.dina(n8848), .dinb(n8805), .dout(n8849));
  jxor g08782(.dina(n8849), .dinb(n8796), .dout(n8850));
  jnot g08783(.din(n8850), .dout(n8851));
  jor  g08784(.dina(n4343), .dinb(n2740), .dout(n8852));
  jor  g08785(.dina(n4346), .dinb(n2553), .dout(n8853));
  jor  g08786(.dina(n4348), .dinb(n2738), .dout(n8854));
  jand g08787(.dina(n8854), .dinb(n8853), .dout(n8855));
  jor  g08788(.dina(n3683), .dinb(n2629), .dout(n8856));
  jand g08789(.dina(n8856), .dinb(n8855), .dout(n8857));
  jand g08790(.dina(n8857), .dinb(n8852), .dout(n8858));
  jxor g08791(.dina(n8858), .dinb(\a[29] ), .dout(n8859));
  jxor g08792(.dina(n8859), .dinb(n8851), .dout(n8860));
  jnot g08793(.din(n8860), .dout(n8861));
  jor  g08794(.dina(n3440), .dinb(n2303), .dout(n8862));
  jor  g08795(.dina(n3203), .dinb(n2306), .dout(n8863));
  jor  g08796(.dina(n3286), .dinb(n2309), .dout(n8864));
  jand g08797(.dina(n8864), .dinb(n8863), .dout(n8865));
  jor  g08798(.dina(n3072), .dinb(n1805), .dout(n8866));
  jand g08799(.dina(n8866), .dinb(n8865), .dout(n8867));
  jand g08800(.dina(n8867), .dinb(n8862), .dout(n8868));
  jxor g08801(.dina(n8868), .dinb(\a[26] ), .dout(n8869));
  jxor g08802(.dina(n8869), .dinb(n8861), .dout(n8870));
  jxor g08803(.dina(n8870), .dinb(n8793), .dout(n8871));
  jor  g08804(.dina(n4051), .dinb(n807), .dout(n8872));
  jor  g08805(.dina(n3787), .dinb(n1613), .dout(n8873));
  jor  g08806(.dina(n3863), .dinb(n1621), .dout(n8874));
  jor  g08807(.dina(n3420), .dinb(n1617), .dout(n8875));
  jand g08808(.dina(n8875), .dinb(n8874), .dout(n8876));
  jand g08809(.dina(n8876), .dinb(n8873), .dout(n8877));
  jand g08810(.dina(n8877), .dinb(n8872), .dout(n8878));
  jxor g08811(.dina(n8878), .dinb(n65), .dout(n8879));
  jxor g08812(.dina(n8879), .dinb(n8871), .dout(n8880));
  jxor g08813(.dina(n8880), .dinb(n8790), .dout(n8881));
  jor  g08814(.dina(n4473), .dinb(n1820), .dout(n8882));
  jor  g08815(.dina(n4019), .dinb(n2181), .dout(n8883));
  jor  g08816(.dina(n3929), .dinb(n2186), .dout(n8884));
  jor  g08817(.dina(n4471), .dinb(n2189), .dout(n8885));
  jand g08818(.dina(n8885), .dinb(n8884), .dout(n8886));
  jand g08819(.dina(n8886), .dinb(n8883), .dout(n8887));
  jand g08820(.dina(n8887), .dinb(n8882), .dout(n8888));
  jxor g08821(.dina(n8888), .dinb(n2196), .dout(n8889));
  jxor g08822(.dina(n8889), .dinb(n8881), .dout(n8890));
  jxor g08823(.dina(n8890), .dinb(n8785), .dout(n8891));
  jor  g08824(.dina(n4688), .dinb(n2744), .dout(n8892));
  jor  g08825(.dina(n4526), .dinb(n2749), .dout(n8893));
  jor  g08826(.dina(n4596), .dinb(n2758), .dout(n8894));
  jor  g08827(.dina(n4686), .dinb(n2753), .dout(n8895));
  jand g08828(.dina(n8895), .dinb(n8894), .dout(n8896));
  jand g08829(.dina(n8896), .dinb(n8893), .dout(n8897));
  jand g08830(.dina(n8897), .dinb(n8892), .dout(n8898));
  jxor g08831(.dina(n8898), .dinb(n2441), .dout(n8899));
  jxor g08832(.dina(n8899), .dinb(n8891), .dout(n8900));
  jxor g08833(.dina(n8900), .dinb(n8780), .dout(n8901));
  jnot g08834(.din(n8901), .dout(n8902));
  jor  g08835(.dina(n5549), .dinb(n3424), .dout(n8903));
  jor  g08836(.dina(n5422), .dinb(n3429), .dout(n8904));
  jor  g08837(.dina(n5364), .dinb(n3426), .dout(n8905));
  jand g08838(.dina(n8905), .dinb(n8904), .dout(n8906));
  jor  g08839(.dina(n5264), .dinb(n3211), .dout(n8907));
  jand g08840(.dina(n8907), .dinb(n8906), .dout(n8908));
  jand g08841(.dina(n8908), .dinb(n8903), .dout(n8909));
  jxor g08842(.dina(n8909), .dinb(\a[14] ), .dout(n8910));
  jxor g08843(.dina(n8910), .dinb(n8902), .dout(n8911));
  jxor g08844(.dina(n8911), .dinb(n8777), .dout(n8912));
  jnot g08845(.din(n8912), .dout(n8913));
  jor  g08846(.dina(n6516), .dinb(n4023), .dout(n8914));
  jor  g08847(.dina(n6205), .dinb(n4028), .dout(n8915));
  jor  g08848(.dina(n6390), .dinb(n4025), .dout(n8916));
  jand g08849(.dina(n8916), .dinb(n8915), .dout(n8917));
  jor  g08850(.dina(n5525), .dinb(n3871), .dout(n8918));
  jand g08851(.dina(n8918), .dinb(n8917), .dout(n8919));
  jand g08852(.dina(n8919), .dinb(n8914), .dout(n8920));
  jxor g08853(.dina(n8920), .dinb(\a[11] ), .dout(n8921));
  jxor g08854(.dina(n8921), .dinb(n8913), .dout(n8922));
  jxor g08855(.dina(n8922), .dinb(n8774), .dout(n8923));
  jnot g08856(.din(n8923), .dout(n8924));
  jor  g08857(.dina(n7301), .dinb(n4705), .dout(n8925));
  jor  g08858(.dina(n7303), .dinb(n4692), .dout(n8926));
  jor  g08859(.dina(n6297), .dinb(n4702), .dout(n8927));
  jor  g08860(.dina(n6489), .dinb(n4697), .dout(n8928));
  jand g08861(.dina(n8928), .dinb(n8927), .dout(n8929));
  jand g08862(.dina(n8929), .dinb(n8926), .dout(n8930));
  jand g08863(.dina(n8930), .dinb(n8925), .dout(n8931));
  jxor g08864(.dina(n8931), .dinb(\a[8] ), .dout(n8932));
  jxor g08865(.dina(n8932), .dinb(n8924), .dout(n8933));
  jxor g08866(.dina(n8933), .dinb(n8771), .dout(n8934));
  jxor g08867(.dina(n8934), .dinb(n8759), .dout(n8935));
  jxor g08868(.dina(n8935), .dinb(n8754), .dout(n8936));
  jxor g08869(.dina(n8936), .dinb(n8723), .dout(n8937));
  jxor g08870(.dina(n8937), .dinb(n8751), .dout(n8938));
  jand g08871(.dina(n8938), .dinb(n1819), .dout(n8939));
  jand g08872(.dina(n8723), .dinb(n2180), .dout(n8940));
  jand g08873(.dina(n8936), .dinb(n2243), .dout(n8941));
  jor  g08874(.dina(n8941), .dinb(n8940), .dout(n8942));
  jand g08875(.dina(n8740), .dinb(n2185), .dout(n8943));
  jor  g08876(.dina(n8943), .dinb(n8942), .dout(n8944));
  jor  g08877(.dina(n8944), .dinb(n8939), .dout(n8945));
  jxor g08878(.dina(n8945), .dinb(n2196), .dout(n8946));
  jor  g08879(.dina(n8946), .dinb(n8281), .dout(n8947));
  jxor g08880(.dina(n8037), .dinb(n7706), .dout(n8948));
  jnot g08881(.din(n8948), .dout(n8949));
  jxor g08882(.dina(n8749), .dinb(n8748), .dout(n8950));
  jand g08883(.dina(n8950), .dinb(n1819), .dout(n8951));
  jand g08884(.dina(n8740), .dinb(n2180), .dout(n8952));
  jand g08885(.dina(n8723), .dinb(n2243), .dout(n8953));
  jor  g08886(.dina(n8953), .dinb(n8952), .dout(n8954));
  jand g08887(.dina(n8268), .dinb(n2185), .dout(n8955));
  jor  g08888(.dina(n8955), .dinb(n8954), .dout(n8956));
  jor  g08889(.dina(n8956), .dinb(n8951), .dout(n8957));
  jxor g08890(.dina(n8957), .dinb(n2196), .dout(n8958));
  jor  g08891(.dina(n8958), .dinb(n8949), .dout(n8959));
  jor  g08892(.dina(n7325), .dinb(n65), .dout(n8960));
  jxor g08893(.dina(n8960), .dinb(n7701), .dout(n8961));
  jxor g08894(.dina(n8746), .dinb(n8745), .dout(n8962));
  jand g08895(.dina(n8962), .dinb(n1819), .dout(n8963));
  jand g08896(.dina(n8740), .dinb(n2243), .dout(n8964));
  jand g08897(.dina(n8268), .dinb(n2180), .dout(n8965));
  jand g08898(.dina(n8022), .dinb(n2185), .dout(n8966));
  jor  g08899(.dina(n8966), .dinb(n8965), .dout(n8967));
  jor  g08900(.dina(n8967), .dinb(n8964), .dout(n8968));
  jor  g08901(.dina(n8968), .dinb(n8963), .dout(n8969));
  jxor g08902(.dina(n8969), .dinb(\a[20] ), .dout(n8970));
  jand g08903(.dina(n8970), .dinb(n8961), .dout(n8971));
  jand g08904(.dina(n7322), .dinb(\a[23] ), .dout(n8972));
  jxor g08905(.dina(n8972), .dinb(n7320), .dout(n8973));
  jnot g08906(.din(n8973), .dout(n8974));
  jand g08907(.dina(n8270), .dinb(n1819), .dout(n8975));
  jand g08908(.dina(n8022), .dinb(n2180), .dout(n8976));
  jand g08909(.dina(n8268), .dinb(n2243), .dout(n8977));
  jor  g08910(.dina(n8977), .dinb(n8976), .dout(n8978));
  jand g08911(.dina(n7692), .dinb(n2185), .dout(n8979));
  jor  g08912(.dina(n8979), .dinb(n8978), .dout(n8980));
  jor  g08913(.dina(n8980), .dinb(n8975), .dout(n8981));
  jxor g08914(.dina(n8981), .dinb(n2196), .dout(n8982));
  jor  g08915(.dina(n8982), .dinb(n8974), .dout(n8983));
  jand g08916(.dina(n7315), .dinb(n1819), .dout(n8984));
  jand g08917(.dina(n7019), .dinb(n2180), .dout(n8985));
  jand g08918(.dina(n7313), .dinb(n2243), .dout(n8986));
  jor  g08919(.dina(n8986), .dinb(n8985), .dout(n8987));
  jor  g08920(.dina(n8987), .dinb(n8984), .dout(n8988));
  jnot g08921(.din(n8988), .dout(n8989));
  jand g08922(.dina(n7019), .dinb(n1817), .dout(n8990));
  jnot g08923(.din(n8990), .dout(n8991));
  jand g08924(.dina(n8991), .dinb(\a[20] ), .dout(n8992));
  jand g08925(.dina(n8992), .dinb(n8989), .dout(n8993));
  jand g08926(.dina(n7693), .dinb(n1819), .dout(n8994));
  jand g08927(.dina(n7313), .dinb(n2180), .dout(n8995));
  jor  g08928(.dina(n8995), .dinb(n8994), .dout(n8996));
  jand g08929(.dina(n7692), .dinb(n2243), .dout(n8997));
  jand g08930(.dina(n7019), .dinb(n2185), .dout(n8998));
  jor  g08931(.dina(n8998), .dinb(n8997), .dout(n8999));
  jor  g08932(.dina(n8999), .dinb(n8996), .dout(n9000));
  jnot g08933(.din(n9000), .dout(n9001));
  jand g08934(.dina(n9001), .dinb(n8993), .dout(n9002));
  jand g08935(.dina(n9002), .dinb(n7322), .dout(n9003));
  jnot g08936(.din(n9003), .dout(n9004));
  jxor g08937(.dina(n9002), .dinb(n7322), .dout(n9005));
  jnot g08938(.din(n9005), .dout(n9006));
  jand g08939(.dina(n8029), .dinb(n1819), .dout(n9007));
  jand g08940(.dina(n7692), .dinb(n2180), .dout(n9008));
  jand g08941(.dina(n8022), .dinb(n2243), .dout(n9009));
  jor  g08942(.dina(n9009), .dinb(n9008), .dout(n9010));
  jand g08943(.dina(n7313), .dinb(n2185), .dout(n9011));
  jor  g08944(.dina(n9011), .dinb(n9010), .dout(n9012));
  jor  g08945(.dina(n9012), .dinb(n9007), .dout(n9013));
  jxor g08946(.dina(n9013), .dinb(n2196), .dout(n9014));
  jor  g08947(.dina(n9014), .dinb(n9006), .dout(n9015));
  jand g08948(.dina(n9015), .dinb(n9004), .dout(n9016));
  jnot g08949(.din(n9016), .dout(n9017));
  jxor g08950(.dina(n8982), .dinb(n8974), .dout(n9018));
  jand g08951(.dina(n9018), .dinb(n9017), .dout(n9019));
  jnot g08952(.din(n9019), .dout(n9020));
  jand g08953(.dina(n9020), .dinb(n8983), .dout(n9021));
  jnot g08954(.din(n9021), .dout(n9022));
  jxor g08955(.dina(n8970), .dinb(n8961), .dout(n9023));
  jand g08956(.dina(n9023), .dinb(n9022), .dout(n9024));
  jor  g08957(.dina(n9024), .dinb(n8971), .dout(n9025));
  jxor g08958(.dina(n8958), .dinb(n8949), .dout(n9026));
  jand g08959(.dina(n9026), .dinb(n9025), .dout(n9027));
  jnot g08960(.din(n9027), .dout(n9028));
  jand g08961(.dina(n9028), .dinb(n8959), .dout(n9029));
  jnot g08962(.din(n9029), .dout(n9030));
  jxor g08963(.dina(n8946), .dinb(n8281), .dout(n9031));
  jand g08964(.dina(n9031), .dinb(n9030), .dout(n9032));
  jnot g08965(.din(n9032), .dout(n9033));
  jand g08966(.dina(n9033), .dinb(n8947), .dout(n9034));
  jnot g08967(.din(n9034), .dout(n9035));
  jor  g08968(.dina(n8278), .dinb(n8048), .dout(n9036));
  jand g08969(.dina(n8279), .dinb(n8040), .dout(n9037));
  jnot g08970(.din(n9037), .dout(n9038));
  jand g08971(.dina(n9038), .dinb(n9036), .dout(n9039));
  jnot g08972(.din(n9039), .dout(n9040));
  jand g08973(.dina(n8962), .dinb(n806), .dout(n9041));
  jand g08974(.dina(n8268), .dinb(n1612), .dout(n9042));
  jand g08975(.dina(n8740), .dinb(n1620), .dout(n9043));
  jor  g08976(.dina(n9043), .dinb(n9042), .dout(n9044));
  jand g08977(.dina(n8022), .dinb(n1644), .dout(n9045));
  jor  g08978(.dina(n9045), .dinb(n9044), .dout(n9046));
  jor  g08979(.dina(n9046), .dinb(n9041), .dout(n9047));
  jxor g08980(.dina(n9047), .dinb(n65), .dout(n9048));
  jnot g08981(.din(n9048), .dout(n9049));
  jand g08982(.dina(n7693), .dinb(n71), .dout(n9050));
  jand g08983(.dina(n7313), .dinb(n731), .dout(n9051));
  jor  g08984(.dina(n9051), .dinb(n9050), .dout(n9052));
  jand g08985(.dina(n7692), .dinb(n796), .dout(n9053));
  jand g08986(.dina(n7019), .dinb(n1806), .dout(n9054));
  jor  g08987(.dina(n9054), .dinb(n9053), .dout(n9055));
  jor  g08988(.dina(n9055), .dinb(n9052), .dout(n9056));
  jor  g08989(.dina(n7020), .dinb(n77), .dout(n9057));
  jor  g08990(.dina(n9057), .dinb(n8045), .dout(n9058));
  jand g08991(.dina(n9058), .dinb(\a[26] ), .dout(n9059));
  jxor g08992(.dina(n9059), .dinb(n9056), .dout(n9060));
  jxor g08993(.dina(n9060), .dinb(n9049), .dout(n9061));
  jxor g08994(.dina(n9061), .dinb(n9040), .dout(n9062));
  jnot g08995(.din(n9062), .dout(n9063));
  jand g08996(.dina(n8936), .dinb(n8723), .dout(n9064));
  jand g08997(.dina(n8937), .dinb(n8751), .dout(n9065));
  jor  g08998(.dina(n9065), .dinb(n9064), .dout(n9066));
  jor  g08999(.dina(n8770), .dinb(n8764), .dout(n9067));
  jnot g09000(.din(n9067), .dout(n9068));
  jand g09001(.dina(n8933), .dinb(n8771), .dout(n9069));
  jor  g09002(.dina(n9069), .dinb(n9068), .dout(n9070));
  jand g09003(.dina(n8922), .dinb(n8774), .dout(n9071));
  jnot g09004(.din(n9071), .dout(n9072));
  jor  g09005(.dina(n8932), .dinb(n8924), .dout(n9073));
  jand g09006(.dina(n9073), .dinb(n9072), .dout(n9074));
  jand g09007(.dina(n8256), .dinb(n5280), .dout(n9075));
  jor  g09008(.dina(n9075), .dinb(n5536), .dout(n9076));
  jand g09009(.dina(n9076), .dinb(n8000), .dout(n9077));
  jxor g09010(.dina(n9077), .dinb(n5277), .dout(n9078));
  jxor g09011(.dina(n9078), .dinb(n9074), .dout(n9079));
  jand g09012(.dina(n8911), .dinb(n8777), .dout(n9080));
  jnot g09013(.din(n9080), .dout(n9081));
  jor  g09014(.dina(n8921), .dinb(n8913), .dout(n9082));
  jand g09015(.dina(n9082), .dinb(n9081), .dout(n9083));
  jnot g09016(.din(n9083), .dout(n9084));
  jand g09017(.dina(n8900), .dinb(n8780), .dout(n9085));
  jnot g09018(.din(n9085), .dout(n9086));
  jor  g09019(.dina(n8910), .dinb(n8902), .dout(n9087));
  jand g09020(.dina(n9087), .dinb(n9086), .dout(n9088));
  jnot g09021(.din(n9088), .dout(n9089));
  jand g09022(.dina(n8890), .dinb(n8785), .dout(n9090));
  jand g09023(.dina(n8899), .dinb(n8891), .dout(n9091));
  jor  g09024(.dina(n9091), .dinb(n9090), .dout(n9092));
  jand g09025(.dina(n8880), .dinb(n8790), .dout(n9093));
  jand g09026(.dina(n8889), .dinb(n8881), .dout(n9094));
  jor  g09027(.dina(n9094), .dinb(n9093), .dout(n9095));
  jand g09028(.dina(n8870), .dinb(n8793), .dout(n9096));
  jand g09029(.dina(n8879), .dinb(n8871), .dout(n9097));
  jor  g09030(.dina(n9097), .dinb(n9096), .dout(n9098));
  jor  g09031(.dina(n8859), .dinb(n8851), .dout(n9099));
  jor  g09032(.dina(n8869), .dinb(n8861), .dout(n9100));
  jand g09033(.dina(n9100), .dinb(n9099), .dout(n9101));
  jnot g09034(.din(n9101), .dout(n9102));
  jand g09035(.dina(n8848), .dinb(n8805), .dout(n9103));
  jand g09036(.dina(n8849), .dinb(n8796), .dout(n9104));
  jor  g09037(.dina(n9104), .dinb(n9103), .dout(n9105));
  jor  g09038(.dina(n7061), .dinb(n2779), .dout(n9106));
  jand g09039(.dina(n6050), .dinb(n2325), .dout(n9107));
  jand g09040(.dina(n5084), .dinb(n2630), .dout(n9108));
  jor  g09041(.dina(n9108), .dinb(n9107), .dout(n9109));
  jand g09042(.dina(n5082), .dinb(n2633), .dout(n9110));
  jor  g09043(.dina(n9110), .dinb(n9109), .dout(n9111));
  jnot g09044(.din(n9111), .dout(n9112));
  jand g09045(.dina(n9112), .dinb(n9106), .dout(n9113));
  jnot g09046(.din(n9113), .dout(n9114));
  jor  g09047(.dina(n8846), .dinb(n6219), .dout(n9115));
  jand g09048(.dina(n8847), .dinb(n8810), .dout(n9116));
  jnot g09049(.din(n9116), .dout(n9117));
  jand g09050(.dina(n9117), .dinb(n9115), .dout(n9118));
  jnot g09051(.din(n9118), .dout(n9119));
  jand g09052(.dina(n6183), .dinb(n920), .dout(n9120));
  jand g09053(.dina(n714), .dinb(n135), .dout(n9121));
  jand g09054(.dina(n9121), .dinb(n171), .dout(n9122));
  jand g09055(.dina(n9122), .dinb(n2384), .dout(n9123));
  jand g09056(.dina(n9123), .dinb(n9120), .dout(n9124));
  jand g09057(.dina(n1090), .dinb(n691), .dout(n9125));
  jand g09058(.dina(n9125), .dinb(n1040), .dout(n9126));
  jand g09059(.dina(n2100), .dinb(n718), .dout(n9127));
  jand g09060(.dina(n9127), .dinb(n1687), .dout(n9128));
  jand g09061(.dina(n9128), .dinb(n9126), .dout(n9129));
  jand g09062(.dina(n8580), .dinb(n1834), .dout(n9130));
  jand g09063(.dina(n9130), .dinb(n9129), .dout(n9131));
  jand g09064(.dina(n950), .dinb(n463), .dout(n9132));
  jand g09065(.dina(n9132), .dinb(n3977), .dout(n9133));
  jand g09066(.dina(n9133), .dinb(n9131), .dout(n9134));
  jand g09067(.dina(n909), .dinb(n1333), .dout(n9135));
  jand g09068(.dina(n2148), .dinb(n948), .dout(n9136));
  jand g09069(.dina(n9136), .dinb(n664), .dout(n9137));
  jand g09070(.dina(n9137), .dinb(n9135), .dout(n9138));
  jand g09071(.dina(n3117), .dinb(n589), .dout(n9139));
  jand g09072(.dina(n9139), .dinb(n9138), .dout(n9140));
  jand g09073(.dina(n1714), .dinb(n517), .dout(n9141));
  jand g09074(.dina(n9141), .dinb(n1096), .dout(n9142));
  jand g09075(.dina(n9142), .dinb(n8115), .dout(n9143));
  jand g09076(.dina(n9143), .dinb(n9140), .dout(n9144));
  jand g09077(.dina(n9144), .dinb(n2701), .dout(n9145));
  jand g09078(.dina(n9145), .dinb(n1521), .dout(n9146));
  jand g09079(.dina(n9146), .dinb(n9134), .dout(n9147));
  jand g09080(.dina(n9147), .dinb(n9124), .dout(n9148));
  jxor g09081(.dina(n9148), .dinb(n6219), .dout(n9149));
  jxor g09082(.dina(n9149), .dinb(n9119), .dout(n9150));
  jxor g09083(.dina(n9150), .dinb(n9114), .dout(n9151));
  jxor g09084(.dina(n9151), .dinb(n9105), .dout(n9152));
  jnot g09085(.din(n9152), .dout(n9153));
  jor  g09086(.dina(n3081), .dinb(n4343), .dout(n9154));
  jor  g09087(.dina(n3683), .dinb(n2553), .dout(n9155));
  jor  g09088(.dina(n4346), .dinb(n2738), .dout(n9156));
  jand g09089(.dina(n9156), .dinb(n9155), .dout(n9157));
  jor  g09090(.dina(n3072), .dinb(n4348), .dout(n9158));
  jand g09091(.dina(n9158), .dinb(n9157), .dout(n9159));
  jand g09092(.dina(n9159), .dinb(n9154), .dout(n9160));
  jxor g09093(.dina(n9160), .dinb(\a[29] ), .dout(n9161));
  jxor g09094(.dina(n9161), .dinb(n9153), .dout(n9162));
  jor  g09095(.dina(n3422), .dinb(n2303), .dout(n9163));
  jor  g09096(.dina(n3203), .dinb(n1805), .dout(n9164));
  jor  g09097(.dina(n3420), .dinb(n2309), .dout(n9165));
  jor  g09098(.dina(n3286), .dinb(n2306), .dout(n9166));
  jand g09099(.dina(n9166), .dinb(n9165), .dout(n9167));
  jand g09100(.dina(n9167), .dinb(n9164), .dout(n9168));
  jand g09101(.dina(n9168), .dinb(n9163), .dout(n9169));
  jxor g09102(.dina(n9169), .dinb(n77), .dout(n9170));
  jxor g09103(.dina(n9170), .dinb(n9162), .dout(n9171));
  jxor g09104(.dina(n9171), .dinb(n9102), .dout(n9172));
  jnot g09105(.din(n9172), .dout(n9173));
  jor  g09106(.dina(n4038), .dinb(n807), .dout(n9174));
  jor  g09107(.dina(n3863), .dinb(n1613), .dout(n9175));
  jor  g09108(.dina(n3929), .dinb(n1621), .dout(n9176));
  jand g09109(.dina(n9176), .dinb(n9175), .dout(n9177));
  jor  g09110(.dina(n3787), .dinb(n1617), .dout(n9178));
  jand g09111(.dina(n9178), .dinb(n9177), .dout(n9179));
  jand g09112(.dina(n9179), .dinb(n9174), .dout(n9180));
  jxor g09113(.dina(n9180), .dinb(\a[23] ), .dout(n9181));
  jxor g09114(.dina(n9181), .dinb(n9173), .dout(n9182));
  jxor g09115(.dina(n9182), .dinb(n9098), .dout(n9183));
  jor  g09116(.dina(n4726), .dinb(n1820), .dout(n9184));
  jor  g09117(.dina(n4471), .dinb(n2181), .dout(n9185));
  jor  g09118(.dina(n4019), .dinb(n2186), .dout(n9186));
  jor  g09119(.dina(n4596), .dinb(n2189), .dout(n9187));
  jand g09120(.dina(n9187), .dinb(n9186), .dout(n9188));
  jand g09121(.dina(n9188), .dinb(n9185), .dout(n9189));
  jand g09122(.dina(n9189), .dinb(n9184), .dout(n9190));
  jxor g09123(.dina(n9190), .dinb(n2196), .dout(n9191));
  jxor g09124(.dina(n9191), .dinb(n9183), .dout(n9192));
  jxor g09125(.dina(n9192), .dinb(n9095), .dout(n9193));
  jor  g09126(.dina(n5266), .dinb(n2744), .dout(n9194));
  jor  g09127(.dina(n4686), .dinb(n2749), .dout(n9195));
  jor  g09128(.dina(n5264), .dinb(n2753), .dout(n9196));
  jor  g09129(.dina(n4526), .dinb(n2758), .dout(n9197));
  jand g09130(.dina(n9197), .dinb(n9196), .dout(n9198));
  jand g09131(.dina(n9198), .dinb(n9195), .dout(n9199));
  jand g09132(.dina(n9199), .dinb(n9194), .dout(n9200));
  jxor g09133(.dina(n9200), .dinb(n2441), .dout(n9201));
  jxor g09134(.dina(n9201), .dinb(n9193), .dout(n9202));
  jxor g09135(.dina(n9202), .dinb(n9092), .dout(n9203));
  jor  g09136(.dina(n5527), .dinb(n3424), .dout(n9204));
  jor  g09137(.dina(n5364), .dinb(n3429), .dout(n9205));
  jor  g09138(.dina(n5422), .dinb(n3211), .dout(n9206));
  jor  g09139(.dina(n5525), .dinb(n3426), .dout(n9207));
  jand g09140(.dina(n9207), .dinb(n9206), .dout(n9208));
  jand g09141(.dina(n9208), .dinb(n9205), .dout(n9209));
  jand g09142(.dina(n9209), .dinb(n9204), .dout(n9210));
  jxor g09143(.dina(n9210), .dinb(n3473), .dout(n9211));
  jxor g09144(.dina(n9211), .dinb(n9203), .dout(n9212));
  jxor g09145(.dina(n9212), .dinb(n9089), .dout(n9213));
  jor  g09146(.dina(n6999), .dinb(n4023), .dout(n9214));
  jor  g09147(.dina(n6390), .dinb(n4028), .dout(n9215));
  jor  g09148(.dina(n6205), .dinb(n3871), .dout(n9216));
  jor  g09149(.dina(n6297), .dinb(n4025), .dout(n9217));
  jand g09150(.dina(n9217), .dinb(n9216), .dout(n9218));
  jand g09151(.dina(n9218), .dinb(n9215), .dout(n9219));
  jand g09152(.dina(n9219), .dinb(n9214), .dout(n9220));
  jxor g09153(.dina(n9220), .dinb(n4050), .dout(n9221));
  jxor g09154(.dina(n9221), .dinb(n9213), .dout(n9222));
  jxor g09155(.dina(n9222), .dinb(n9084), .dout(n9223));
  jor  g09156(.dina(n7682), .dinb(n4692), .dout(n9224));
  jor  g09157(.dina(n7301), .dinb(n4697), .dout(n9225));
  jor  g09158(.dina(n6489), .dinb(n4702), .dout(n9226));
  jor  g09159(.dina(n7680), .dinb(n4705), .dout(n9227));
  jand g09160(.dina(n9227), .dinb(n9226), .dout(n9228));
  jand g09161(.dina(n9228), .dinb(n9225), .dout(n9229));
  jand g09162(.dina(n9229), .dinb(n9224), .dout(n9230));
  jxor g09163(.dina(n9230), .dinb(n4713), .dout(n9231));
  jxor g09164(.dina(n9231), .dinb(n9223), .dout(n9232));
  jxor g09165(.dina(n9232), .dinb(n9079), .dout(n9233));
  jxor g09166(.dina(n9233), .dinb(n9070), .dout(n9234));
  jnot g09167(.din(n9234), .dout(n9235));
  jand g09168(.dina(n8934), .dinb(n8759), .dout(n9236));
  jnot g09169(.din(n9236), .dout(n9237));
  jnot g09170(.din(n8752), .dout(n9238));
  jnot g09171(.din(n8510), .dout(n9239));
  jor  g09172(.dina(n8739), .dinb(n8725), .dout(n9240));
  jand g09173(.dina(n9240), .dinb(n9239), .dout(n9241));
  jnot g09174(.din(n8522), .dout(n9242));
  jxor g09175(.dina(n8721), .dinb(n9242), .dout(n9243));
  jor  g09176(.dina(n9243), .dinb(n9241), .dout(n9244));
  jand g09177(.dina(n9244), .dinb(n9238), .dout(n9245));
  jnot g09178(.din(n8934), .dout(n9246));
  jxor g09179(.dina(n9246), .dinb(n8759), .dout(n9247));
  jor  g09180(.dina(n9247), .dinb(n9245), .dout(n9248));
  jand g09181(.dina(n9248), .dinb(n9237), .dout(n9249));
  jxor g09182(.dina(n9249), .dinb(n9235), .dout(n9250));
  jxor g09183(.dina(n9250), .dinb(n8936), .dout(n9251));
  jxor g09184(.dina(n9251), .dinb(n9066), .dout(n9252));
  jand g09185(.dina(n9252), .dinb(n1819), .dout(n9253));
  jand g09186(.dina(n8936), .dinb(n2180), .dout(n9254));
  jand g09187(.dina(n9250), .dinb(n2243), .dout(n9255));
  jor  g09188(.dina(n9255), .dinb(n9254), .dout(n9256));
  jand g09189(.dina(n8723), .dinb(n2185), .dout(n9257));
  jor  g09190(.dina(n9257), .dinb(n9256), .dout(n9258));
  jor  g09191(.dina(n9258), .dinb(n9253), .dout(n9259));
  jxor g09192(.dina(n9259), .dinb(n2196), .dout(n9260));
  jxor g09193(.dina(n9260), .dinb(n9063), .dout(n9261));
  jxor g09194(.dina(n9261), .dinb(n9035), .dout(n9262));
  jnot g09195(.din(n9262), .dout(n9263));
  jor  g09196(.dina(n9078), .dinb(n9074), .dout(n9264));
  jnot g09197(.din(n9264), .dout(n9265));
  jand g09198(.dina(n9232), .dinb(n9079), .dout(n9266));
  jor  g09199(.dina(n9266), .dinb(n9265), .dout(n9267));
  jand g09200(.dina(n9212), .dinb(n9089), .dout(n9268));
  jand g09201(.dina(n9221), .dinb(n9213), .dout(n9269));
  jor  g09202(.dina(n9269), .dinb(n9268), .dout(n9270));
  jnot g09203(.din(n9270), .dout(n9271));
  jor  g09204(.dina(n6491), .dinb(n4023), .dout(n9272));
  jor  g09205(.dina(n6297), .dinb(n4028), .dout(n9273));
  jor  g09206(.dina(n6390), .dinb(n3871), .dout(n9274));
  jand g09207(.dina(n9274), .dinb(n9273), .dout(n9275));
  jor  g09208(.dina(n6489), .dinb(n4025), .dout(n9276));
  jand g09209(.dina(n9276), .dinb(n9275), .dout(n9277));
  jand g09210(.dina(n9277), .dinb(n9272), .dout(n9278));
  jxor g09211(.dina(n9278), .dinb(\a[11] ), .dout(n9279));
  jxor g09212(.dina(n9279), .dinb(n9271), .dout(n9280));
  jand g09213(.dina(n9202), .dinb(n9092), .dout(n9281));
  jand g09214(.dina(n9211), .dinb(n9203), .dout(n9282));
  jor  g09215(.dina(n9282), .dinb(n9281), .dout(n9283));
  jand g09216(.dina(n9192), .dinb(n9095), .dout(n9284));
  jand g09217(.dina(n9201), .dinb(n9193), .dout(n9285));
  jor  g09218(.dina(n9285), .dinb(n9284), .dout(n9286));
  jand g09219(.dina(n9182), .dinb(n9098), .dout(n9287));
  jand g09220(.dina(n9191), .dinb(n9183), .dout(n9288));
  jor  g09221(.dina(n9288), .dinb(n9287), .dout(n9289));
  jand g09222(.dina(n9171), .dinb(n9102), .dout(n9290));
  jnot g09223(.din(n9290), .dout(n9291));
  jor  g09224(.dina(n9181), .dinb(n9173), .dout(n9292));
  jand g09225(.dina(n9292), .dinb(n9291), .dout(n9293));
  jnot g09226(.din(n9293), .dout(n9294));
  jor  g09227(.dina(n9161), .dinb(n9153), .dout(n9295));
  jand g09228(.dina(n9170), .dinb(n9162), .dout(n9296));
  jnot g09229(.din(n9296), .dout(n9297));
  jand g09230(.dina(n9297), .dinb(n9295), .dout(n9298));
  jnot g09231(.din(n9298), .dout(n9299));
  jand g09232(.dina(n9150), .dinb(n9114), .dout(n9300));
  jand g09233(.dina(n9151), .dinb(n9105), .dout(n9301));
  jor  g09234(.dina(n9301), .dinb(n9300), .dout(n9302));
  jor  g09235(.dina(n7061), .dinb(n2768), .dout(n9303));
  jand g09236(.dina(n5084), .dinb(n2554), .dout(n9304));
  jand g09237(.dina(n6050), .dinb(n2633), .dout(n9305));
  jor  g09238(.dina(n9305), .dinb(n9304), .dout(n9306));
  jand g09239(.dina(n5082), .dinb(n2630), .dout(n9307));
  jor  g09240(.dina(n9307), .dinb(n9306), .dout(n9308));
  jnot g09241(.din(n9308), .dout(n9309));
  jand g09242(.dina(n9309), .dinb(n9303), .dout(n9310));
  jnot g09243(.din(n9310), .dout(n9311));
  jor  g09244(.dina(n9148), .dinb(n6219), .dout(n9312));
  jand g09245(.dina(n9149), .dinb(n9119), .dout(n9313));
  jnot g09246(.din(n9313), .dout(n9314));
  jand g09247(.dina(n9314), .dinb(n9312), .dout(n9315));
  jnot g09248(.din(n9315), .dout(n9316));
  jand g09249(.dina(n6381), .dinb(n1872), .dout(n9317));
  jand g09250(.dina(n3829), .dinb(n3328), .dout(n9318));
  jand g09251(.dina(n9318), .dinb(n9317), .dout(n9319));
  jand g09252(.dina(n442), .dinb(n964), .dout(n9320));
  jand g09253(.dina(n9320), .dinb(n1360), .dout(n9321));
  jand g09254(.dina(n9321), .dinb(n1778), .dout(n9322));
  jand g09255(.dina(n833), .dinb(n325), .dout(n9323));
  jand g09256(.dina(n9323), .dinb(n5473), .dout(n9324));
  jand g09257(.dina(n9324), .dinb(n9322), .dout(n9325));
  jand g09258(.dina(n1471), .dinb(n683), .dout(n9326));
  jand g09259(.dina(n9326), .dinb(n1682), .dout(n9327));
  jand g09260(.dina(n9327), .dinb(n9325), .dout(n9328));
  jand g09261(.dina(n9328), .dinb(n8351), .dout(n9329));
  jand g09262(.dina(n9329), .dinb(n9319), .dout(n9330));
  jand g09263(.dina(n3363), .dinb(n1591), .dout(n9331));
  jand g09264(.dina(n547), .dinb(n916), .dout(n9332));
  jand g09265(.dina(n9332), .dinb(n3357), .dout(n9333));
  jand g09266(.dina(n9333), .dinb(n5515), .dout(n9334));
  jand g09267(.dina(n9334), .dinb(n9331), .dout(n9335));
  jand g09268(.dina(n965), .dinb(n171), .dout(n9336));
  jand g09269(.dina(n9336), .dinb(n1230), .dout(n9337));
  jand g09270(.dina(n1713), .dinb(n696), .dout(n9338));
  jand g09271(.dina(n548), .dinb(n654), .dout(n9339));
  jand g09272(.dina(n9339), .dinb(n9338), .dout(n9340));
  jand g09273(.dina(n9340), .dinb(n1542), .dout(n9341));
  jand g09274(.dina(n9341), .dinb(n9337), .dout(n9342));
  jand g09275(.dina(n1511), .dinb(n664), .dout(n9343));
  jand g09276(.dina(n9343), .dinb(n670), .dout(n9344));
  jand g09277(.dina(n1160), .dinb(n136), .dout(n9345));
  jand g09278(.dina(n9345), .dinb(n9344), .dout(n9346));
  jand g09279(.dina(n9346), .dinb(n5294), .dout(n9347));
  jand g09280(.dina(n9347), .dinb(n9342), .dout(n9348));
  jand g09281(.dina(n9348), .dinb(n1366), .dout(n9349));
  jand g09282(.dina(n9349), .dinb(n9335), .dout(n9350));
  jand g09283(.dina(n9350), .dinb(n9330), .dout(n9351));
  jand g09284(.dina(n1167), .dinb(n270), .dout(n9352));
  jand g09285(.dina(n9352), .dinb(n2124), .dout(n9353));
  jand g09286(.dina(n1559), .dinb(n445), .dout(n9354));
  jand g09287(.dina(n1096), .dinb(n672), .dout(n9355));
  jand g09288(.dina(n9355), .dinb(n9354), .dout(n9356));
  jand g09289(.dina(n9356), .dinb(n9353), .dout(n9357));
  jand g09290(.dina(n328), .dinb(n843), .dout(n9358));
  jand g09291(.dina(n9358), .dinb(n1162), .dout(n9359));
  jand g09292(.dina(n9359), .dinb(n8404), .dout(n9360));
  jand g09293(.dina(n9360), .dinb(n9357), .dout(n9361));
  jand g09294(.dina(n9361), .dinb(n3178), .dout(n9362));
  jand g09295(.dina(n3015), .dinb(n1188), .dout(n9363));
  jand g09296(.dina(n873), .dinb(n691), .dout(n9364));
  jand g09297(.dina(n9364), .dinb(n9363), .dout(n9365));
  jand g09298(.dina(n6012), .dinb(n2472), .dout(n9366));
  jand g09299(.dina(n9366), .dinb(n9365), .dout(n9367));
  jand g09300(.dina(n1098), .dinb(n495), .dout(n9368));
  jand g09301(.dina(n9368), .dinb(n1476), .dout(n9369));
  jand g09302(.dina(n1453), .dinb(n1225), .dout(n9370));
  jand g09303(.dina(n925), .dinb(n647), .dout(n9371));
  jand g09304(.dina(n9371), .dinb(n9370), .dout(n9372));
  jand g09305(.dina(n9372), .dinb(n9369), .dout(n9373));
  jand g09306(.dina(n1326), .dinb(n1277), .dout(n9374));
  jand g09307(.dina(n9374), .dinb(n9373), .dout(n9375));
  jand g09308(.dina(n9375), .dinb(n5415), .dout(n9376));
  jand g09309(.dina(n9376), .dinb(n9367), .dout(n9377));
  jand g09310(.dina(n9377), .dinb(n9362), .dout(n9378));
  jand g09311(.dina(n9378), .dinb(n5314), .dout(n9379));
  jand g09312(.dina(n9379), .dinb(n9351), .dout(n9380));
  jxor g09313(.dina(n9380), .dinb(\a[2] ), .dout(n9381));
  jxor g09314(.dina(n9381), .dinb(n5277), .dout(n9382));
  jxor g09315(.dina(n9382), .dinb(n9316), .dout(n9383));
  jxor g09316(.dina(n9383), .dinb(n9311), .dout(n9384));
  jxor g09317(.dina(n9384), .dinb(n9302), .dout(n9385));
  jnot g09318(.din(n9385), .dout(n9386));
  jor  g09319(.dina(n3451), .dinb(n4343), .dout(n9387));
  jor  g09320(.dina(n3072), .dinb(n4346), .dout(n9388));
  jor  g09321(.dina(n3683), .dinb(n2738), .dout(n9389));
  jand g09322(.dina(n9389), .dinb(n9388), .dout(n9390));
  jor  g09323(.dina(n3203), .dinb(n4348), .dout(n9391));
  jand g09324(.dina(n9391), .dinb(n9390), .dout(n9392));
  jand g09325(.dina(n9392), .dinb(n9387), .dout(n9393));
  jxor g09326(.dina(n9393), .dinb(\a[29] ), .dout(n9394));
  jxor g09327(.dina(n9394), .dinb(n9386), .dout(n9395));
  jnot g09328(.din(n9395), .dout(n9396));
  jor  g09329(.dina(n3789), .dinb(n2303), .dout(n9397));
  jor  g09330(.dina(n3420), .dinb(n2306), .dout(n9398));
  jor  g09331(.dina(n3286), .dinb(n1805), .dout(n9399));
  jand g09332(.dina(n9399), .dinb(n9398), .dout(n9400));
  jor  g09333(.dina(n3787), .dinb(n2309), .dout(n9401));
  jand g09334(.dina(n9401), .dinb(n9400), .dout(n9402));
  jand g09335(.dina(n9402), .dinb(n9397), .dout(n9403));
  jxor g09336(.dina(n9403), .dinb(\a[26] ), .dout(n9404));
  jxor g09337(.dina(n9404), .dinb(n9396), .dout(n9405));
  jxor g09338(.dina(n9405), .dinb(n9299), .dout(n9406));
  jor  g09339(.dina(n4021), .dinb(n807), .dout(n9407));
  jor  g09340(.dina(n3863), .dinb(n1617), .dout(n9408));
  jor  g09341(.dina(n4019), .dinb(n1621), .dout(n9409));
  jor  g09342(.dina(n3929), .dinb(n1613), .dout(n9410));
  jand g09343(.dina(n9410), .dinb(n9409), .dout(n9411));
  jand g09344(.dina(n9411), .dinb(n9408), .dout(n9412));
  jand g09345(.dina(n9412), .dinb(n9407), .dout(n9413));
  jxor g09346(.dina(n9413), .dinb(n65), .dout(n9414));
  jxor g09347(.dina(n9414), .dinb(n9406), .dout(n9415));
  jxor g09348(.dina(n9415), .dinb(n9294), .dout(n9416));
  jor  g09349(.dina(n4714), .dinb(n1820), .dout(n9417));
  jor  g09350(.dina(n4596), .dinb(n2181), .dout(n9418));
  jor  g09351(.dina(n4471), .dinb(n2186), .dout(n9419));
  jor  g09352(.dina(n4526), .dinb(n2189), .dout(n9420));
  jand g09353(.dina(n9420), .dinb(n9419), .dout(n9421));
  jand g09354(.dina(n9421), .dinb(n9418), .dout(n9422));
  jand g09355(.dina(n9422), .dinb(n9417), .dout(n9423));
  jxor g09356(.dina(n9423), .dinb(n2196), .dout(n9424));
  jxor g09357(.dina(n9424), .dinb(n9416), .dout(n9425));
  jxor g09358(.dina(n9425), .dinb(n9289), .dout(n9426));
  jor  g09359(.dina(n5560), .dinb(n2744), .dout(n9427));
  jor  g09360(.dina(n5264), .dinb(n2749), .dout(n9428));
  jor  g09361(.dina(n4686), .dinb(n2758), .dout(n9429));
  jor  g09362(.dina(n5422), .dinb(n2753), .dout(n9430));
  jand g09363(.dina(n9430), .dinb(n9429), .dout(n9431));
  jand g09364(.dina(n9431), .dinb(n9428), .dout(n9432));
  jand g09365(.dina(n9432), .dinb(n9427), .dout(n9433));
  jxor g09366(.dina(n9433), .dinb(n2441), .dout(n9434));
  jxor g09367(.dina(n9434), .dinb(n9426), .dout(n9435));
  jxor g09368(.dina(n9435), .dinb(n9286), .dout(n9436));
  jor  g09369(.dina(n6207), .dinb(n3424), .dout(n9437));
  jor  g09370(.dina(n5525), .dinb(n3429), .dout(n9438));
  jor  g09371(.dina(n5364), .dinb(n3211), .dout(n9439));
  jor  g09372(.dina(n6205), .dinb(n3426), .dout(n9440));
  jand g09373(.dina(n9440), .dinb(n9439), .dout(n9441));
  jand g09374(.dina(n9441), .dinb(n9438), .dout(n9442));
  jand g09375(.dina(n9442), .dinb(n9437), .dout(n9443));
  jxor g09376(.dina(n9443), .dinb(n3473), .dout(n9444));
  jxor g09377(.dina(n9444), .dinb(n9436), .dout(n9445));
  jxor g09378(.dina(n9445), .dinb(n9283), .dout(n9446));
  jxor g09379(.dina(n9446), .dinb(n9280), .dout(n9447));
  jand g09380(.dina(n9222), .dinb(n9084), .dout(n9448));
  jand g09381(.dina(n9231), .dinb(n9223), .dout(n9449));
  jor  g09382(.dina(n9449), .dinb(n9448), .dout(n9450));
  jnot g09383(.din(n9450), .dout(n9451));
  jor  g09384(.dina(n7301), .dinb(n4702), .dout(n9452));
  jor  g09385(.dina(n8002), .dinb(n4692), .dout(n9453));
  jor  g09386(.dina(n7999), .dinb(n4705), .dout(n9454));
  jor  g09387(.dina(n7680), .dinb(n4697), .dout(n9455));
  jand g09388(.dina(n9455), .dinb(n9454), .dout(n9456));
  jand g09389(.dina(n9456), .dinb(n9453), .dout(n9457));
  jand g09390(.dina(n9457), .dinb(n9452), .dout(n9458));
  jxor g09391(.dina(n9458), .dinb(\a[8] ), .dout(n9459));
  jxor g09392(.dina(n9459), .dinb(n9451), .dout(n9460));
  jxor g09393(.dina(n9460), .dinb(n9447), .dout(n9461));
  jand g09394(.dina(n9461), .dinb(n9267), .dout(n9462));
  jand g09395(.dina(n9233), .dinb(n9070), .dout(n9463));
  jand g09396(.dina(n8935), .dinb(n8754), .dout(n9464));
  jor  g09397(.dina(n9464), .dinb(n9236), .dout(n9465));
  jand g09398(.dina(n9465), .dinb(n9234), .dout(n9466));
  jor  g09399(.dina(n9466), .dinb(n9463), .dout(n9467));
  jxor g09400(.dina(n9461), .dinb(n9267), .dout(n9468));
  jand g09401(.dina(n9468), .dinb(n9467), .dout(n9469));
  jor  g09402(.dina(n9469), .dinb(n9462), .dout(n9470));
  jor  g09403(.dina(n9459), .dinb(n9451), .dout(n9471));
  jnot g09404(.din(n9471), .dout(n9472));
  jand g09405(.dina(n9460), .dinb(n9447), .dout(n9473));
  jor  g09406(.dina(n9473), .dinb(n9472), .dout(n9474));
  jor  g09407(.dina(n9279), .dinb(n9271), .dout(n9475));
  jand g09408(.dina(n9446), .dinb(n9280), .dout(n9476));
  jnot g09409(.din(n9476), .dout(n9477));
  jand g09410(.dina(n9477), .dinb(n9475), .dout(n9478));
  jor  g09411(.dina(n7999), .dinb(n4697), .dout(n9479));
  jor  g09412(.dina(n8260), .dinb(n4692), .dout(n9480));
  jor  g09413(.dina(n7680), .dinb(n4702), .dout(n9481));
  jand g09414(.dina(n9481), .dinb(n9480), .dout(n9482));
  jand g09415(.dina(n9482), .dinb(n9479), .dout(n9483));
  jxor g09416(.dina(n9483), .dinb(\a[8] ), .dout(n9484));
  jxor g09417(.dina(n9484), .dinb(n9478), .dout(n9485));
  jand g09418(.dina(n9444), .dinb(n9436), .dout(n9486));
  jand g09419(.dina(n9445), .dinb(n9283), .dout(n9487));
  jor  g09420(.dina(n9487), .dinb(n9486), .dout(n9488));
  jand g09421(.dina(n9434), .dinb(n9426), .dout(n9489));
  jand g09422(.dina(n9435), .dinb(n9286), .dout(n9490));
  jor  g09423(.dina(n9490), .dinb(n9489), .dout(n9491));
  jand g09424(.dina(n9424), .dinb(n9416), .dout(n9492));
  jand g09425(.dina(n9425), .dinb(n9289), .dout(n9493));
  jor  g09426(.dina(n9493), .dinb(n9492), .dout(n9494));
  jand g09427(.dina(n9414), .dinb(n9406), .dout(n9495));
  jand g09428(.dina(n9415), .dinb(n9294), .dout(n9496));
  jor  g09429(.dina(n9496), .dinb(n9495), .dout(n9497));
  jor  g09430(.dina(n9404), .dinb(n9396), .dout(n9498));
  jand g09431(.dina(n9405), .dinb(n9299), .dout(n9499));
  jnot g09432(.din(n9499), .dout(n9500));
  jand g09433(.dina(n9500), .dinb(n9498), .dout(n9501));
  jnot g09434(.din(n9501), .dout(n9502));
  jand g09435(.dina(n9384), .dinb(n9302), .dout(n9503));
  jnot g09436(.din(n9503), .dout(n9504));
  jor  g09437(.dina(n9394), .dinb(n9386), .dout(n9505));
  jand g09438(.dina(n9505), .dinb(n9504), .dout(n9506));
  jnot g09439(.din(n9506), .dout(n9507));
  jand g09440(.dina(n9382), .dinb(n9316), .dout(n9508));
  jand g09441(.dina(n9383), .dinb(n9311), .dout(n9509));
  jor  g09442(.dina(n9509), .dinb(n9508), .dout(n9510));
  jor  g09443(.dina(n7061), .dinb(n2740), .dout(n9511));
  jand g09444(.dina(n5082), .dinb(n2554), .dout(n9512));
  jand g09445(.dina(n5084), .dinb(n3074), .dout(n9513));
  jor  g09446(.dina(n9513), .dinb(n9512), .dout(n9514));
  jand g09447(.dina(n6050), .dinb(n2630), .dout(n9515));
  jor  g09448(.dina(n9515), .dinb(n9514), .dout(n9516));
  jnot g09449(.din(n9516), .dout(n9517));
  jand g09450(.dina(n9517), .dinb(n9511), .dout(n9518));
  jnot g09451(.din(n9518), .dout(n9519));
  jand g09452(.dina(n1167), .dinb(n1005), .dout(n9520));
  jand g09453(.dina(n9520), .dinb(n1159), .dout(n9521));
  jand g09454(.dina(n534), .dinb(n1575), .dout(n9522));
  jand g09455(.dina(n9522), .dinb(n9521), .dout(n9523));
  jand g09456(.dina(n3161), .dinb(n681), .dout(n9524));
  jand g09457(.dina(n9524), .dinb(n9523), .dout(n9525));
  jand g09458(.dina(n1713), .dinb(n838), .dout(n9526));
  jand g09459(.dina(n9526), .dinb(n641), .dout(n9527));
  jand g09460(.dina(n9527), .dinb(n325), .dout(n9528));
  jand g09461(.dina(n9528), .dinb(n9525), .dout(n9529));
  jand g09462(.dina(n9529), .dinb(n8605), .dout(n9530));
  jand g09463(.dina(n9530), .dinb(n7792), .dout(n9531));
  jand g09464(.dina(n1839), .dinb(n600), .dout(n9532));
  jand g09465(.dina(n9532), .dinb(n511), .dout(n9533));
  jand g09466(.dina(n672), .dinb(n2117), .dout(n9534));
  jand g09467(.dina(n9534), .dinb(n843), .dout(n9535));
  jand g09468(.dina(n1426), .dinb(n676), .dout(n9536));
  jand g09469(.dina(n9536), .dinb(n9535), .dout(n9537));
  jand g09470(.dina(n9537), .dinb(n9533), .dout(n9538));
  jand g09471(.dina(n3094), .dinb(n1098), .dout(n9539));
  jand g09472(.dina(n2100), .dinb(n1260), .dout(n9540));
  jand g09473(.dina(n9540), .dinb(n480), .dout(n9541));
  jand g09474(.dina(n9541), .dinb(n981), .dout(n9542));
  jand g09475(.dina(n9542), .dinb(n9539), .dout(n9543));
  jand g09476(.dina(n1739), .dinb(n586), .dout(n9544));
  jand g09477(.dina(n1096), .dinb(n811), .dout(n9545));
  jand g09478(.dina(n9545), .dinb(n9544), .dout(n9546));
  jand g09479(.dina(n2508), .dinb(n1753), .dout(n9547));
  jand g09480(.dina(n9547), .dinb(n9546), .dout(n9548));
  jand g09481(.dina(n4541), .dinb(n988), .dout(n9549));
  jand g09482(.dina(n9549), .dinb(n3747), .dout(n9550));
  jand g09483(.dina(n9550), .dinb(n9548), .dout(n9551));
  jand g09484(.dina(n9551), .dinb(n9543), .dout(n9552));
  jand g09485(.dina(n9552), .dinb(n9538), .dout(n9553));
  jand g09486(.dina(n664), .dinb(n114), .dout(n9554));
  jand g09487(.dina(n9554), .dinb(n1577), .dout(n9555));
  jand g09488(.dina(n893), .dinb(n171), .dout(n9556));
  jand g09489(.dina(n9556), .dinb(n2352), .dout(n9557));
  jand g09490(.dina(n9557), .dinb(n9555), .dout(n9558));
  jand g09491(.dina(n2379), .dinb(n1846), .dout(n9559));
  jand g09492(.dina(n870), .dinb(n1259), .dout(n9560));
  jand g09493(.dina(n9560), .dinb(n9559), .dout(n9561));
  jand g09494(.dina(n9561), .dinb(n9558), .dout(n9562));
  jand g09495(.dina(n6374), .dinb(n1532), .dout(n9563));
  jand g09496(.dina(n9563), .dinb(n4618), .dout(n9564));
  jand g09497(.dina(n9564), .dinb(n9562), .dout(n9565));
  jand g09498(.dina(n1212), .dinb(n1042), .dout(n9566));
  jand g09499(.dina(n9566), .dinb(n8400), .dout(n9567));
  jand g09500(.dina(n9567), .dinb(n3060), .dout(n9568));
  jand g09501(.dina(n9568), .dinb(n916), .dout(n9569));
  jand g09502(.dina(n9569), .dinb(n9565), .dout(n9570));
  jand g09503(.dina(n9570), .dinb(n9553), .dout(n9571));
  jand g09504(.dina(n9571), .dinb(n9531), .dout(n9572));
  jnot g09505(.din(n9572), .dout(n9573));
  jor  g09506(.dina(n9380), .dinb(\a[2] ), .dout(n9574));
  jand g09507(.dina(n9381), .dinb(n5277), .dout(n9575));
  jnot g09508(.din(n9575), .dout(n9576));
  jand g09509(.dina(n9576), .dinb(n9574), .dout(n9577));
  jxor g09510(.dina(n9577), .dinb(n9573), .dout(n9578));
  jxor g09511(.dina(n9578), .dinb(n9519), .dout(n9579));
  jxor g09512(.dina(n9579), .dinb(n9510), .dout(n9580));
  jnot g09513(.din(n9580), .dout(n9581));
  jor  g09514(.dina(n3440), .dinb(n4343), .dout(n9582));
  jor  g09515(.dina(n3203), .dinb(n4346), .dout(n9583));
  jor  g09516(.dina(n3286), .dinb(n4348), .dout(n9584));
  jand g09517(.dina(n9584), .dinb(n9583), .dout(n9585));
  jor  g09518(.dina(n3683), .dinb(n3072), .dout(n9586));
  jand g09519(.dina(n9586), .dinb(n9585), .dout(n9587));
  jand g09520(.dina(n9587), .dinb(n9582), .dout(n9588));
  jxor g09521(.dina(n9588), .dinb(\a[29] ), .dout(n9589));
  jxor g09522(.dina(n9589), .dinb(n9581), .dout(n9590));
  jxor g09523(.dina(n9590), .dinb(n9507), .dout(n9591));
  jor  g09524(.dina(n4051), .dinb(n2303), .dout(n9592));
  jor  g09525(.dina(n3787), .dinb(n2306), .dout(n9593));
  jor  g09526(.dina(n3863), .dinb(n2309), .dout(n9594));
  jor  g09527(.dina(n3420), .dinb(n1805), .dout(n9595));
  jand g09528(.dina(n9595), .dinb(n9594), .dout(n9596));
  jand g09529(.dina(n9596), .dinb(n9593), .dout(n9597));
  jand g09530(.dina(n9597), .dinb(n9592), .dout(n9598));
  jxor g09531(.dina(n9598), .dinb(n77), .dout(n9599));
  jxor g09532(.dina(n9599), .dinb(n9591), .dout(n9600));
  jxor g09533(.dina(n9600), .dinb(n9502), .dout(n9601));
  jor  g09534(.dina(n4473), .dinb(n807), .dout(n9602));
  jor  g09535(.dina(n4019), .dinb(n1613), .dout(n9603));
  jor  g09536(.dina(n3929), .dinb(n1617), .dout(n9604));
  jor  g09537(.dina(n4471), .dinb(n1621), .dout(n9605));
  jand g09538(.dina(n9605), .dinb(n9604), .dout(n9606));
  jand g09539(.dina(n9606), .dinb(n9603), .dout(n9607));
  jand g09540(.dina(n9607), .dinb(n9602), .dout(n9608));
  jxor g09541(.dina(n9608), .dinb(n65), .dout(n9609));
  jxor g09542(.dina(n9609), .dinb(n9601), .dout(n9610));
  jxor g09543(.dina(n9610), .dinb(n9497), .dout(n9611));
  jor  g09544(.dina(n4688), .dinb(n1820), .dout(n9612));
  jor  g09545(.dina(n4526), .dinb(n2181), .dout(n9613));
  jor  g09546(.dina(n4596), .dinb(n2186), .dout(n9614));
  jor  g09547(.dina(n4686), .dinb(n2189), .dout(n9615));
  jand g09548(.dina(n9615), .dinb(n9614), .dout(n9616));
  jand g09549(.dina(n9616), .dinb(n9613), .dout(n9617));
  jand g09550(.dina(n9617), .dinb(n9612), .dout(n9618));
  jxor g09551(.dina(n9618), .dinb(n2196), .dout(n9619));
  jxor g09552(.dina(n9619), .dinb(n9611), .dout(n9620));
  jxor g09553(.dina(n9620), .dinb(n9494), .dout(n9621));
  jnot g09554(.din(n9621), .dout(n9622));
  jor  g09555(.dina(n5549), .dinb(n2744), .dout(n9623));
  jor  g09556(.dina(n5422), .dinb(n2749), .dout(n9624));
  jor  g09557(.dina(n5364), .dinb(n2753), .dout(n9625));
  jand g09558(.dina(n9625), .dinb(n9624), .dout(n9626));
  jor  g09559(.dina(n5264), .dinb(n2758), .dout(n9627));
  jand g09560(.dina(n9627), .dinb(n9626), .dout(n9628));
  jand g09561(.dina(n9628), .dinb(n9623), .dout(n9629));
  jxor g09562(.dina(n9629), .dinb(\a[17] ), .dout(n9630));
  jxor g09563(.dina(n9630), .dinb(n9622), .dout(n9631));
  jxor g09564(.dina(n9631), .dinb(n9491), .dout(n9632));
  jnot g09565(.din(n9632), .dout(n9633));
  jor  g09566(.dina(n6516), .dinb(n3424), .dout(n9634));
  jor  g09567(.dina(n6205), .dinb(n3429), .dout(n9635));
  jor  g09568(.dina(n6390), .dinb(n3426), .dout(n9636));
  jand g09569(.dina(n9636), .dinb(n9635), .dout(n9637));
  jor  g09570(.dina(n5525), .dinb(n3211), .dout(n9638));
  jand g09571(.dina(n9638), .dinb(n9637), .dout(n9639));
  jand g09572(.dina(n9639), .dinb(n9634), .dout(n9640));
  jxor g09573(.dina(n9640), .dinb(\a[14] ), .dout(n9641));
  jxor g09574(.dina(n9641), .dinb(n9633), .dout(n9642));
  jxor g09575(.dina(n9642), .dinb(n9488), .dout(n9643));
  jor  g09576(.dina(n7303), .dinb(n4023), .dout(n9644));
  jor  g09577(.dina(n7301), .dinb(n4025), .dout(n9645));
  jor  g09578(.dina(n6297), .dinb(n3871), .dout(n9646));
  jor  g09579(.dina(n6489), .dinb(n4028), .dout(n9647));
  jand g09580(.dina(n9647), .dinb(n9646), .dout(n9648));
  jand g09581(.dina(n9648), .dinb(n9645), .dout(n9649));
  jand g09582(.dina(n9649), .dinb(n9644), .dout(n9650));
  jxor g09583(.dina(n9650), .dinb(n4050), .dout(n9651));
  jxor g09584(.dina(n9651), .dinb(n9643), .dout(n9652));
  jxor g09585(.dina(n9652), .dinb(n9485), .dout(n9653));
  jxor g09586(.dina(n9653), .dinb(n9474), .dout(n9654));
  jxor g09587(.dina(n9654), .dinb(n9470), .dout(n9655));
  jxor g09588(.dina(n9468), .dinb(n9467), .dout(n9656));
  jand g09589(.dina(n9656), .dinb(n9655), .dout(n9657));
  jand g09590(.dina(n9656), .dinb(n9250), .dout(n9658));
  jand g09591(.dina(n9250), .dinb(n8936), .dout(n9659));
  jand g09592(.dina(n9251), .dinb(n9066), .dout(n9660));
  jor  g09593(.dina(n9660), .dinb(n9659), .dout(n9661));
  jxor g09594(.dina(n9656), .dinb(n9250), .dout(n9662));
  jand g09595(.dina(n9662), .dinb(n9661), .dout(n9663));
  jor  g09596(.dina(n9663), .dinb(n9658), .dout(n9664));
  jxor g09597(.dina(n9656), .dinb(n9655), .dout(n9665));
  jand g09598(.dina(n9665), .dinb(n9664), .dout(n9666));
  jor  g09599(.dina(n9666), .dinb(n9657), .dout(n9667));
  jor  g09600(.dina(n9484), .dinb(n9478), .dout(n9668));
  jand g09601(.dina(n9652), .dinb(n9485), .dout(n9669));
  jnot g09602(.din(n9669), .dout(n9670));
  jand g09603(.dina(n9670), .dinb(n9668), .dout(n9671));
  jnot g09604(.din(n9671), .dout(n9672));
  jand g09605(.dina(n9642), .dinb(n9488), .dout(n9673));
  jand g09606(.dina(n9651), .dinb(n9643), .dout(n9674));
  jor  g09607(.dina(n9674), .dinb(n9673), .dout(n9675));
  jnot g09608(.din(n9675), .dout(n9676));
  jand g09609(.dina(n8256), .dinb(n4691), .dout(n9677));
  jor  g09610(.dina(n9677), .dinb(n4701), .dout(n9678));
  jand g09611(.dina(n9678), .dinb(n8000), .dout(n9679));
  jxor g09612(.dina(n9679), .dinb(n4713), .dout(n9680));
  jxor g09613(.dina(n9680), .dinb(n9676), .dout(n9681));
  jand g09614(.dina(n9631), .dinb(n9491), .dout(n9682));
  jnot g09615(.din(n9682), .dout(n9683));
  jor  g09616(.dina(n9641), .dinb(n9633), .dout(n9684));
  jand g09617(.dina(n9684), .dinb(n9683), .dout(n9685));
  jnot g09618(.din(n9685), .dout(n9686));
  jand g09619(.dina(n9620), .dinb(n9494), .dout(n9687));
  jnot g09620(.din(n9687), .dout(n9688));
  jor  g09621(.dina(n9630), .dinb(n9622), .dout(n9689));
  jand g09622(.dina(n9689), .dinb(n9688), .dout(n9690));
  jnot g09623(.din(n9690), .dout(n9691));
  jand g09624(.dina(n9610), .dinb(n9497), .dout(n9692));
  jand g09625(.dina(n9619), .dinb(n9611), .dout(n9693));
  jor  g09626(.dina(n9693), .dinb(n9692), .dout(n9694));
  jand g09627(.dina(n9600), .dinb(n9502), .dout(n9695));
  jand g09628(.dina(n9609), .dinb(n9601), .dout(n9696));
  jor  g09629(.dina(n9696), .dinb(n9695), .dout(n9697));
  jand g09630(.dina(n9590), .dinb(n9507), .dout(n9698));
  jand g09631(.dina(n9599), .dinb(n9591), .dout(n9699));
  jor  g09632(.dina(n9699), .dinb(n9698), .dout(n9700));
  jand g09633(.dina(n9579), .dinb(n9510), .dout(n9701));
  jnot g09634(.din(n9701), .dout(n9702));
  jor  g09635(.dina(n9589), .dinb(n9581), .dout(n9703));
  jand g09636(.dina(n9703), .dinb(n9702), .dout(n9704));
  jnot g09637(.din(n9704), .dout(n9705));
  jor  g09638(.dina(n7061), .dinb(n3081), .dout(n9706));
  jand g09639(.dina(n6050), .dinb(n2554), .dout(n9707));
  jand g09640(.dina(n5082), .dinb(n3074), .dout(n9708));
  jor  g09641(.dina(n9708), .dinb(n9707), .dout(n9709));
  jand g09642(.dina(n5084), .dinb(n3290), .dout(n9710));
  jor  g09643(.dina(n9710), .dinb(n9709), .dout(n9711));
  jnot g09644(.din(n9711), .dout(n9712));
  jand g09645(.dina(n9712), .dinb(n9706), .dout(n9713));
  jnot g09646(.din(n9713), .dout(n9714));
  jor  g09647(.dina(n9577), .dinb(n9573), .dout(n9715));
  jand g09648(.dina(n9578), .dinb(n9519), .dout(n9716));
  jnot g09649(.din(n9716), .dout(n9717));
  jand g09650(.dina(n9717), .dinb(n9715), .dout(n9718));
  jnot g09651(.din(n9718), .dout(n9719));
  jand g09652(.dina(n895), .dinb(n1345), .dout(n9720));
  jand g09653(.dina(n9720), .dinb(n1697), .dout(n9721));
  jand g09654(.dina(n1851), .dinb(n1583), .dout(n9722));
  jand g09655(.dina(n9722), .dinb(n5231), .dout(n9723));
  jand g09656(.dina(n9723), .dinb(n9721), .dout(n9724));
  jand g09657(.dina(n586), .dinb(n178), .dout(n9725));
  jand g09658(.dina(n2148), .dinb(n328), .dout(n9726));
  jand g09659(.dina(n9726), .dinb(n2142), .dout(n9727));
  jand g09660(.dina(n9727), .dinb(n9725), .dout(n9728));
  jand g09661(.dina(n9728), .dinb(n9724), .dout(n9729));
  jand g09662(.dina(n9729), .dinb(n2587), .dout(n9730));
  jand g09663(.dina(n2052), .dinb(n1868), .dout(n9731));
  jand g09664(.dina(n9731), .dinb(n3417), .dout(n9732));
  jand g09665(.dina(n1351), .dinb(n900), .dout(n9733));
  jand g09666(.dina(n9733), .dinb(n664), .dout(n9734));
  jand g09667(.dina(n9734), .dinb(n1189), .dout(n9735));
  jand g09668(.dina(n3771), .dinb(n456), .dout(n9736));
  jand g09669(.dina(n8603), .dinb(n172), .dout(n9737));
  jand g09670(.dina(n9737), .dinb(n9736), .dout(n9738));
  jand g09671(.dina(n9738), .dinb(n9735), .dout(n9739));
  jand g09672(.dina(n9739), .dinb(n1569), .dout(n9740));
  jand g09673(.dina(n9740), .dinb(n9732), .dout(n9741));
  jand g09674(.dina(n9741), .dinb(n9730), .dout(n9742));
  jand g09675(.dina(n9525), .dinb(n6441), .dout(n9743));
  jand g09676(.dina(n9743), .dinb(n938), .dout(n9744));
  jand g09677(.dina(n9744), .dinb(n9742), .dout(n9745));
  jand g09678(.dina(n1560), .dinb(n122), .dout(n9746));
  jand g09679(.dina(n9746), .dinb(n1686), .dout(n9747));
  jand g09680(.dina(n9747), .dinb(n716), .dout(n9748));
  jand g09681(.dina(n1744), .dinb(n1213), .dout(n9749));
  jand g09682(.dina(n9749), .dinb(n632), .dout(n9750));
  jand g09683(.dina(n1515), .dinb(n481), .dout(n9751));
  jand g09684(.dina(n9751), .dinb(n3276), .dout(n9752));
  jand g09685(.dina(n2086), .dinb(n1043), .dout(n9753));
  jand g09686(.dina(n9753), .dinb(n9752), .dout(n9754));
  jand g09687(.dina(n9754), .dinb(n9750), .dout(n9755));
  jand g09688(.dina(n660), .dinb(n430), .dout(n9756));
  jand g09689(.dina(n3840), .dinb(n1053), .dout(n9757));
  jand g09690(.dina(n9757), .dinb(n9756), .dout(n9758));
  jand g09691(.dina(n9758), .dinb(n6186), .dout(n9759));
  jand g09692(.dina(n9759), .dinb(n9755), .dout(n9760));
  jand g09693(.dina(n9760), .dinb(n9748), .dout(n9761));
  jand g09694(.dina(n2100), .dinb(n831), .dout(n9762));
  jand g09695(.dina(n9762), .dinb(n672), .dout(n9763));
  jand g09696(.dina(n516), .dinb(n349), .dout(n9764));
  jand g09697(.dina(n9764), .dinb(n9763), .dout(n9765));
  jand g09698(.dina(n668), .dinb(n829), .dout(n9766));
  jand g09699(.dina(n9766), .dinb(n1334), .dout(n9767));
  jand g09700(.dina(n700), .dinb(n583), .dout(n9768));
  jand g09701(.dina(n9768), .dinb(n1107), .dout(n9769));
  jand g09702(.dina(n9769), .dinb(n9767), .dout(n9770));
  jand g09703(.dina(n9770), .dinb(n9765), .dout(n9771));
  jand g09704(.dina(n3978), .dinb(n2357), .dout(n9772));
  jand g09705(.dina(n9772), .dinb(n2538), .dout(n9773));
  jand g09706(.dina(n647), .dinb(n1778), .dout(n9774));
  jand g09707(.dina(n9774), .dinb(n824), .dout(n9775));
  jand g09708(.dina(n9775), .dinb(n1219), .dout(n9776));
  jand g09709(.dina(n563), .dinb(n1306), .dout(n9777));
  jand g09710(.dina(n9777), .dinb(n9776), .dout(n9778));
  jand g09711(.dina(n9778), .dinb(n9773), .dout(n9779));
  jand g09712(.dina(n9779), .dinb(n9771), .dout(n9780));
  jand g09713(.dina(n9780), .dinb(n9761), .dout(n9781));
  jand g09714(.dina(n9781), .dinb(n9745), .dout(n9782));
  jxor g09715(.dina(n9782), .dinb(n9573), .dout(n9783));
  jxor g09716(.dina(n9783), .dinb(n9719), .dout(n9784));
  jxor g09717(.dina(n9784), .dinb(n9714), .dout(n9785));
  jxor g09718(.dina(n9785), .dinb(n9705), .dout(n9786));
  jor  g09719(.dina(n3422), .dinb(n4343), .dout(n9787));
  jor  g09720(.dina(n3683), .dinb(n3203), .dout(n9788));
  jor  g09721(.dina(n3420), .dinb(n4348), .dout(n9789));
  jor  g09722(.dina(n3286), .dinb(n4346), .dout(n9790));
  jand g09723(.dina(n9790), .dinb(n9789), .dout(n9791));
  jand g09724(.dina(n9791), .dinb(n9788), .dout(n9792));
  jand g09725(.dina(n9792), .dinb(n9787), .dout(n9793));
  jxor g09726(.dina(n9793), .dinb(n93), .dout(n9794));
  jxor g09727(.dina(n9794), .dinb(n9786), .dout(n9795));
  jnot g09728(.din(n9795), .dout(n9796));
  jor  g09729(.dina(n4038), .dinb(n2303), .dout(n9797));
  jor  g09730(.dina(n3863), .dinb(n2306), .dout(n9798));
  jor  g09731(.dina(n3929), .dinb(n2309), .dout(n9799));
  jand g09732(.dina(n9799), .dinb(n9798), .dout(n9800));
  jor  g09733(.dina(n3787), .dinb(n1805), .dout(n9801));
  jand g09734(.dina(n9801), .dinb(n9800), .dout(n9802));
  jand g09735(.dina(n9802), .dinb(n9797), .dout(n9803));
  jxor g09736(.dina(n9803), .dinb(\a[26] ), .dout(n9804));
  jxor g09737(.dina(n9804), .dinb(n9796), .dout(n9805));
  jxor g09738(.dina(n9805), .dinb(n9700), .dout(n9806));
  jor  g09739(.dina(n4726), .dinb(n807), .dout(n9807));
  jor  g09740(.dina(n4471), .dinb(n1613), .dout(n9808));
  jor  g09741(.dina(n4596), .dinb(n1621), .dout(n9809));
  jor  g09742(.dina(n4019), .dinb(n1617), .dout(n9810));
  jand g09743(.dina(n9810), .dinb(n9809), .dout(n9811));
  jand g09744(.dina(n9811), .dinb(n9808), .dout(n9812));
  jand g09745(.dina(n9812), .dinb(n9807), .dout(n9813));
  jxor g09746(.dina(n9813), .dinb(n65), .dout(n9814));
  jxor g09747(.dina(n9814), .dinb(n9806), .dout(n9815));
  jxor g09748(.dina(n9815), .dinb(n9697), .dout(n9816));
  jor  g09749(.dina(n5266), .dinb(n1820), .dout(n9817));
  jor  g09750(.dina(n4686), .dinb(n2181), .dout(n9818));
  jor  g09751(.dina(n5264), .dinb(n2189), .dout(n9819));
  jor  g09752(.dina(n4526), .dinb(n2186), .dout(n9820));
  jand g09753(.dina(n9820), .dinb(n9819), .dout(n9821));
  jand g09754(.dina(n9821), .dinb(n9818), .dout(n9822));
  jand g09755(.dina(n9822), .dinb(n9817), .dout(n9823));
  jxor g09756(.dina(n9823), .dinb(n2196), .dout(n9824));
  jxor g09757(.dina(n9824), .dinb(n9816), .dout(n9825));
  jxor g09758(.dina(n9825), .dinb(n9694), .dout(n9826));
  jor  g09759(.dina(n5527), .dinb(n2744), .dout(n9827));
  jor  g09760(.dina(n5364), .dinb(n2749), .dout(n9828));
  jor  g09761(.dina(n5422), .dinb(n2758), .dout(n9829));
  jor  g09762(.dina(n5525), .dinb(n2753), .dout(n9830));
  jand g09763(.dina(n9830), .dinb(n9829), .dout(n9831));
  jand g09764(.dina(n9831), .dinb(n9828), .dout(n9832));
  jand g09765(.dina(n9832), .dinb(n9827), .dout(n9833));
  jxor g09766(.dina(n9833), .dinb(n2441), .dout(n9834));
  jxor g09767(.dina(n9834), .dinb(n9826), .dout(n9835));
  jxor g09768(.dina(n9835), .dinb(n9691), .dout(n9836));
  jnot g09769(.din(n9836), .dout(n9837));
  jor  g09770(.dina(n6999), .dinb(n3424), .dout(n9838));
  jor  g09771(.dina(n6390), .dinb(n3429), .dout(n9839));
  jor  g09772(.dina(n6297), .dinb(n3426), .dout(n9840));
  jand g09773(.dina(n9840), .dinb(n9839), .dout(n9841));
  jor  g09774(.dina(n6205), .dinb(n3211), .dout(n9842));
  jand g09775(.dina(n9842), .dinb(n9841), .dout(n9843));
  jand g09776(.dina(n9843), .dinb(n9838), .dout(n9844));
  jxor g09777(.dina(n9844), .dinb(\a[14] ), .dout(n9845));
  jxor g09778(.dina(n9845), .dinb(n9837), .dout(n9846));
  jxor g09779(.dina(n9846), .dinb(n9686), .dout(n9847));
  jor  g09780(.dina(n7682), .dinb(n4023), .dout(n9848));
  jor  g09781(.dina(n7301), .dinb(n4028), .dout(n9849));
  jor  g09782(.dina(n7680), .dinb(n4025), .dout(n9850));
  jor  g09783(.dina(n6489), .dinb(n3871), .dout(n9851));
  jand g09784(.dina(n9851), .dinb(n9850), .dout(n9852));
  jand g09785(.dina(n9852), .dinb(n9849), .dout(n9853));
  jand g09786(.dina(n9853), .dinb(n9848), .dout(n9854));
  jxor g09787(.dina(n9854), .dinb(n4050), .dout(n9855));
  jxor g09788(.dina(n9855), .dinb(n9847), .dout(n9856));
  jxor g09789(.dina(n9856), .dinb(n9681), .dout(n9857));
  jxor g09790(.dina(n9857), .dinb(n9672), .dout(n9858));
  jnot g09791(.din(n9858), .dout(n9859));
  jand g09792(.dina(n9653), .dinb(n9474), .dout(n9860));
  jnot g09793(.din(n9860), .dout(n9861));
  jnot g09794(.din(n9462), .dout(n9862));
  jnot g09795(.din(n9463), .dout(n9863));
  jor  g09796(.dina(n9249), .dinb(n9235), .dout(n9864));
  jand g09797(.dina(n9864), .dinb(n9863), .dout(n9865));
  jnot g09798(.din(n9468), .dout(n9866));
  jor  g09799(.dina(n9866), .dinb(n9865), .dout(n9867));
  jand g09800(.dina(n9867), .dinb(n9862), .dout(n9868));
  jnot g09801(.din(n9654), .dout(n9869));
  jor  g09802(.dina(n9869), .dinb(n9868), .dout(n9870));
  jand g09803(.dina(n9870), .dinb(n9861), .dout(n9871));
  jxor g09804(.dina(n9871), .dinb(n9859), .dout(n9872));
  jxor g09805(.dina(n9872), .dinb(n9655), .dout(n9873));
  jxor g09806(.dina(n9873), .dinb(n9667), .dout(n9874));
  jand g09807(.dina(n9874), .dinb(n2743), .dout(n9875));
  jand g09808(.dina(n9872), .dinb(n2752), .dout(n9876));
  jand g09809(.dina(n9655), .dinb(n2748), .dout(n9877));
  jand g09810(.dina(n9656), .dinb(n2757), .dout(n9878));
  jor  g09811(.dina(n9878), .dinb(n9877), .dout(n9879));
  jor  g09812(.dina(n9879), .dinb(n9876), .dout(n9880));
  jor  g09813(.dina(n9880), .dinb(n9875), .dout(n9881));
  jxor g09814(.dina(n9881), .dinb(n2441), .dout(n9882));
  jor  g09815(.dina(n9882), .dinb(n9263), .dout(n9883));
  jxor g09816(.dina(n9031), .dinb(n9030), .dout(n9884));
  jnot g09817(.din(n9884), .dout(n9885));
  jxor g09818(.dina(n9665), .dinb(n9664), .dout(n9886));
  jand g09819(.dina(n9886), .dinb(n2743), .dout(n9887));
  jand g09820(.dina(n9655), .dinb(n2752), .dout(n9888));
  jand g09821(.dina(n9656), .dinb(n2748), .dout(n9889));
  jand g09822(.dina(n9250), .dinb(n2757), .dout(n9890));
  jor  g09823(.dina(n9890), .dinb(n9889), .dout(n9891));
  jor  g09824(.dina(n9891), .dinb(n9888), .dout(n9892));
  jor  g09825(.dina(n9892), .dinb(n9887), .dout(n9893));
  jxor g09826(.dina(n9893), .dinb(n2441), .dout(n9894));
  jor  g09827(.dina(n9894), .dinb(n9885), .dout(n9895));
  jxor g09828(.dina(n9026), .dinb(n9025), .dout(n9896));
  jnot g09829(.din(n9896), .dout(n9897));
  jxor g09830(.dina(n9662), .dinb(n9661), .dout(n9898));
  jand g09831(.dina(n9898), .dinb(n2743), .dout(n9899));
  jand g09832(.dina(n9656), .dinb(n2752), .dout(n9900));
  jand g09833(.dina(n9250), .dinb(n2748), .dout(n9901));
  jand g09834(.dina(n8936), .dinb(n2757), .dout(n9902));
  jor  g09835(.dina(n9902), .dinb(n9901), .dout(n9903));
  jor  g09836(.dina(n9903), .dinb(n9900), .dout(n9904));
  jor  g09837(.dina(n9904), .dinb(n9899), .dout(n9905));
  jxor g09838(.dina(n9905), .dinb(n2441), .dout(n9906));
  jor  g09839(.dina(n9906), .dinb(n9897), .dout(n9907));
  jxor g09840(.dina(n9023), .dinb(n9022), .dout(n9908));
  jnot g09841(.din(n9908), .dout(n9909));
  jand g09842(.dina(n9252), .dinb(n2743), .dout(n9910));
  jand g09843(.dina(n9250), .dinb(n2752), .dout(n9911));
  jand g09844(.dina(n8936), .dinb(n2748), .dout(n9912));
  jand g09845(.dina(n8723), .dinb(n2757), .dout(n9913));
  jor  g09846(.dina(n9913), .dinb(n9912), .dout(n9914));
  jor  g09847(.dina(n9914), .dinb(n9911), .dout(n9915));
  jor  g09848(.dina(n9915), .dinb(n9910), .dout(n9916));
  jxor g09849(.dina(n9916), .dinb(n2441), .dout(n9917));
  jor  g09850(.dina(n9917), .dinb(n9909), .dout(n9918));
  jxor g09851(.dina(n9018), .dinb(n9017), .dout(n9919));
  jnot g09852(.din(n9919), .dout(n9920));
  jand g09853(.dina(n8938), .dinb(n2743), .dout(n9921));
  jand g09854(.dina(n8936), .dinb(n2752), .dout(n9922));
  jand g09855(.dina(n8723), .dinb(n2748), .dout(n9923));
  jand g09856(.dina(n8740), .dinb(n2757), .dout(n9924));
  jor  g09857(.dina(n9924), .dinb(n9923), .dout(n9925));
  jor  g09858(.dina(n9925), .dinb(n9922), .dout(n9926));
  jor  g09859(.dina(n9926), .dinb(n9921), .dout(n9927));
  jxor g09860(.dina(n9927), .dinb(n2441), .dout(n9928));
  jor  g09861(.dina(n9928), .dinb(n9920), .dout(n9929));
  jxor g09862(.dina(n9014), .dinb(n9006), .dout(n9930));
  jnot g09863(.din(n9930), .dout(n9931));
  jand g09864(.dina(n8950), .dinb(n2743), .dout(n9932));
  jand g09865(.dina(n8723), .dinb(n2752), .dout(n9933));
  jand g09866(.dina(n8740), .dinb(n2748), .dout(n9934));
  jand g09867(.dina(n8268), .dinb(n2757), .dout(n9935));
  jor  g09868(.dina(n9935), .dinb(n9934), .dout(n9936));
  jor  g09869(.dina(n9936), .dinb(n9933), .dout(n9937));
  jor  g09870(.dina(n9937), .dinb(n9932), .dout(n9938));
  jxor g09871(.dina(n9938), .dinb(n2441), .dout(n9939));
  jor  g09872(.dina(n9939), .dinb(n9931), .dout(n9940));
  jand g09873(.dina(n8962), .dinb(n2743), .dout(n9941));
  jand g09874(.dina(n8740), .dinb(n2752), .dout(n9942));
  jand g09875(.dina(n8268), .dinb(n2748), .dout(n9943));
  jand g09876(.dina(n8022), .dinb(n2757), .dout(n9944));
  jor  g09877(.dina(n9944), .dinb(n9943), .dout(n9945));
  jor  g09878(.dina(n9945), .dinb(n9942), .dout(n9946));
  jor  g09879(.dina(n9946), .dinb(n9941), .dout(n9947));
  jxor g09880(.dina(n9947), .dinb(n2441), .dout(n9948));
  jnot g09881(.din(n9948), .dout(n9949));
  jor  g09882(.dina(n8993), .dinb(n2196), .dout(n9950));
  jxor g09883(.dina(n9950), .dinb(n9001), .dout(n9951));
  jand g09884(.dina(n9951), .dinb(n9949), .dout(n9952));
  jand g09885(.dina(n8990), .dinb(\a[20] ), .dout(n9953));
  jxor g09886(.dina(n9953), .dinb(n8988), .dout(n9954));
  jnot g09887(.din(n9954), .dout(n9955));
  jand g09888(.dina(n8270), .dinb(n2743), .dout(n9956));
  jand g09889(.dina(n8022), .dinb(n2748), .dout(n9957));
  jand g09890(.dina(n8268), .dinb(n2752), .dout(n9958));
  jor  g09891(.dina(n9958), .dinb(n9957), .dout(n9959));
  jand g09892(.dina(n7692), .dinb(n2757), .dout(n9960));
  jor  g09893(.dina(n9960), .dinb(n9959), .dout(n9961));
  jor  g09894(.dina(n9961), .dinb(n9956), .dout(n9962));
  jxor g09895(.dina(n9962), .dinb(n2441), .dout(n9963));
  jor  g09896(.dina(n9963), .dinb(n9955), .dout(n9964));
  jand g09897(.dina(n7315), .dinb(n2743), .dout(n9965));
  jand g09898(.dina(n7019), .dinb(n2748), .dout(n9966));
  jand g09899(.dina(n7313), .dinb(n2752), .dout(n9967));
  jor  g09900(.dina(n9967), .dinb(n9966), .dout(n9968));
  jor  g09901(.dina(n9968), .dinb(n9965), .dout(n9969));
  jnot g09902(.din(n9969), .dout(n9970));
  jand g09903(.dina(n7019), .dinb(n2741), .dout(n9971));
  jnot g09904(.din(n9971), .dout(n9972));
  jand g09905(.dina(n9972), .dinb(\a[17] ), .dout(n9973));
  jand g09906(.dina(n9973), .dinb(n9970), .dout(n9974));
  jand g09907(.dina(n7693), .dinb(n2743), .dout(n9975));
  jand g09908(.dina(n7313), .dinb(n2748), .dout(n9976));
  jor  g09909(.dina(n9976), .dinb(n9975), .dout(n9977));
  jand g09910(.dina(n7692), .dinb(n2752), .dout(n9978));
  jand g09911(.dina(n7019), .dinb(n2757), .dout(n9979));
  jor  g09912(.dina(n9979), .dinb(n9978), .dout(n9980));
  jor  g09913(.dina(n9980), .dinb(n9977), .dout(n9981));
  jnot g09914(.din(n9981), .dout(n9982));
  jand g09915(.dina(n9982), .dinb(n9974), .dout(n9983));
  jand g09916(.dina(n9983), .dinb(n8990), .dout(n9984));
  jnot g09917(.din(n9984), .dout(n9985));
  jxor g09918(.dina(n9983), .dinb(n8990), .dout(n9986));
  jnot g09919(.din(n9986), .dout(n9987));
  jand g09920(.dina(n8029), .dinb(n2743), .dout(n9988));
  jand g09921(.dina(n8022), .dinb(n2752), .dout(n9989));
  jand g09922(.dina(n7692), .dinb(n2748), .dout(n9990));
  jand g09923(.dina(n7313), .dinb(n2757), .dout(n9991));
  jor  g09924(.dina(n9991), .dinb(n9990), .dout(n9992));
  jor  g09925(.dina(n9992), .dinb(n9989), .dout(n9993));
  jor  g09926(.dina(n9993), .dinb(n9988), .dout(n9994));
  jxor g09927(.dina(n9994), .dinb(n2441), .dout(n9995));
  jor  g09928(.dina(n9995), .dinb(n9987), .dout(n9996));
  jand g09929(.dina(n9996), .dinb(n9985), .dout(n9997));
  jnot g09930(.din(n9997), .dout(n9998));
  jxor g09931(.dina(n9963), .dinb(n9955), .dout(n9999));
  jand g09932(.dina(n9999), .dinb(n9998), .dout(n10000));
  jnot g09933(.din(n10000), .dout(n10001));
  jand g09934(.dina(n10001), .dinb(n9964), .dout(n10002));
  jnot g09935(.din(n10002), .dout(n10003));
  jxor g09936(.dina(n9951), .dinb(n9949), .dout(n10004));
  jand g09937(.dina(n10004), .dinb(n10003), .dout(n10005));
  jor  g09938(.dina(n10005), .dinb(n9952), .dout(n10006));
  jxor g09939(.dina(n9939), .dinb(n9931), .dout(n10007));
  jand g09940(.dina(n10007), .dinb(n10006), .dout(n10008));
  jnot g09941(.din(n10008), .dout(n10009));
  jand g09942(.dina(n10009), .dinb(n9940), .dout(n10010));
  jnot g09943(.din(n10010), .dout(n10011));
  jxor g09944(.dina(n9928), .dinb(n9920), .dout(n10012));
  jand g09945(.dina(n10012), .dinb(n10011), .dout(n10013));
  jnot g09946(.din(n10013), .dout(n10014));
  jand g09947(.dina(n10014), .dinb(n9929), .dout(n10015));
  jnot g09948(.din(n10015), .dout(n10016));
  jxor g09949(.dina(n9917), .dinb(n9909), .dout(n10017));
  jand g09950(.dina(n10017), .dinb(n10016), .dout(n10018));
  jnot g09951(.din(n10018), .dout(n10019));
  jand g09952(.dina(n10019), .dinb(n9918), .dout(n10020));
  jnot g09953(.din(n10020), .dout(n10021));
  jxor g09954(.dina(n9906), .dinb(n9897), .dout(n10022));
  jand g09955(.dina(n10022), .dinb(n10021), .dout(n10023));
  jnot g09956(.din(n10023), .dout(n10024));
  jand g09957(.dina(n10024), .dinb(n9907), .dout(n10025));
  jnot g09958(.din(n10025), .dout(n10026));
  jxor g09959(.dina(n9894), .dinb(n9885), .dout(n10027));
  jand g09960(.dina(n10027), .dinb(n10026), .dout(n10028));
  jnot g09961(.din(n10028), .dout(n10029));
  jand g09962(.dina(n10029), .dinb(n9895), .dout(n10030));
  jnot g09963(.din(n10030), .dout(n10031));
  jxor g09964(.dina(n9882), .dinb(n9263), .dout(n10032));
  jand g09965(.dina(n10032), .dinb(n10031), .dout(n10033));
  jnot g09966(.din(n10033), .dout(n10034));
  jand g09967(.dina(n10034), .dinb(n9883), .dout(n10035));
  jnot g09968(.din(n10035), .dout(n10036));
  jor  g09969(.dina(n9260), .dinb(n9063), .dout(n10037));
  jand g09970(.dina(n9261), .dinb(n9035), .dout(n10038));
  jnot g09971(.din(n10038), .dout(n10039));
  jand g09972(.dina(n10039), .dinb(n10037), .dout(n10040));
  jnot g09973(.din(n10040), .dout(n10041));
  jand g09974(.dina(n9060), .dinb(n9049), .dout(n10042));
  jand g09975(.dina(n9061), .dinb(n9040), .dout(n10043));
  jor  g09976(.dina(n10043), .dinb(n10042), .dout(n10044));
  jand g09977(.dina(n7019), .dinb(n64), .dout(n10045));
  jnot g09978(.din(n10045), .dout(n10046));
  jor  g09979(.dina(n9058), .dinb(n9056), .dout(n10047));
  jxor g09980(.dina(n10047), .dinb(n10046), .dout(n10048));
  jnot g09981(.din(n10048), .dout(n10049));
  jand g09982(.dina(n8029), .dinb(n71), .dout(n10050));
  jand g09983(.dina(n7692), .dinb(n731), .dout(n10051));
  jand g09984(.dina(n8022), .dinb(n796), .dout(n10052));
  jor  g09985(.dina(n10052), .dinb(n10051), .dout(n10053));
  jand g09986(.dina(n7313), .dinb(n1806), .dout(n10054));
  jor  g09987(.dina(n10054), .dinb(n10053), .dout(n10055));
  jor  g09988(.dina(n10055), .dinb(n10050), .dout(n10056));
  jxor g09989(.dina(n10056), .dinb(n77), .dout(n10057));
  jxor g09990(.dina(n10057), .dinb(n10049), .dout(n10058));
  jnot g09991(.din(n10058), .dout(n10059));
  jand g09992(.dina(n8950), .dinb(n806), .dout(n10060));
  jand g09993(.dina(n8740), .dinb(n1612), .dout(n10061));
  jand g09994(.dina(n8723), .dinb(n1620), .dout(n10062));
  jor  g09995(.dina(n10062), .dinb(n10061), .dout(n10063));
  jand g09996(.dina(n8268), .dinb(n1644), .dout(n10064));
  jor  g09997(.dina(n10064), .dinb(n10063), .dout(n10065));
  jor  g09998(.dina(n10065), .dinb(n10060), .dout(n10066));
  jxor g09999(.dina(n10066), .dinb(n65), .dout(n10067));
  jxor g10000(.dina(n10067), .dinb(n10059), .dout(n10068));
  jxor g10001(.dina(n10068), .dinb(n10044), .dout(n10069));
  jnot g10002(.din(n10069), .dout(n10070));
  jand g10003(.dina(n9898), .dinb(n1819), .dout(n10071));
  jand g10004(.dina(n9250), .dinb(n2180), .dout(n10072));
  jand g10005(.dina(n9656), .dinb(n2243), .dout(n10073));
  jor  g10006(.dina(n10073), .dinb(n10072), .dout(n10074));
  jand g10007(.dina(n8936), .dinb(n2185), .dout(n10075));
  jor  g10008(.dina(n10075), .dinb(n10074), .dout(n10076));
  jor  g10009(.dina(n10076), .dinb(n10071), .dout(n10077));
  jxor g10010(.dina(n10077), .dinb(n2196), .dout(n10078));
  jxor g10011(.dina(n10078), .dinb(n10070), .dout(n10079));
  jxor g10012(.dina(n10079), .dinb(n10041), .dout(n10080));
  jnot g10013(.din(n10080), .dout(n10081));
  jand g10014(.dina(n9872), .dinb(n9655), .dout(n10082));
  jand g10015(.dina(n9873), .dinb(n9667), .dout(n10083));
  jor  g10016(.dina(n10083), .dinb(n10082), .dout(n10084));
  jor  g10017(.dina(n9680), .dinb(n9676), .dout(n10085));
  jand g10018(.dina(n9856), .dinb(n9681), .dout(n10086));
  jnot g10019(.din(n10086), .dout(n10087));
  jand g10020(.dina(n10087), .dinb(n10085), .dout(n10088));
  jnot g10021(.din(n10088), .dout(n10089));
  jand g10022(.dina(n9846), .dinb(n9686), .dout(n10090));
  jand g10023(.dina(n9855), .dinb(n9847), .dout(n10091));
  jor  g10024(.dina(n10091), .dinb(n10090), .dout(n10092));
  jor  g10025(.dina(n8002), .dinb(n4023), .dout(n10093));
  jor  g10026(.dina(n7301), .dinb(n3871), .dout(n10094));
  jor  g10027(.dina(n7999), .dinb(n4025), .dout(n10095));
  jor  g10028(.dina(n7680), .dinb(n4028), .dout(n10096));
  jand g10029(.dina(n10096), .dinb(n10095), .dout(n10097));
  jand g10030(.dina(n10097), .dinb(n10094), .dout(n10098));
  jand g10031(.dina(n10098), .dinb(n10093), .dout(n10099));
  jxor g10032(.dina(n10099), .dinb(n4050), .dout(n10100));
  jxor g10033(.dina(n10100), .dinb(n10092), .dout(n10101));
  jand g10034(.dina(n9835), .dinb(n9691), .dout(n10102));
  jnot g10035(.din(n10102), .dout(n10103));
  jor  g10036(.dina(n9845), .dinb(n9837), .dout(n10104));
  jand g10037(.dina(n10104), .dinb(n10103), .dout(n10105));
  jnot g10038(.din(n10105), .dout(n10106));
  jand g10039(.dina(n9825), .dinb(n9694), .dout(n10107));
  jand g10040(.dina(n9834), .dinb(n9826), .dout(n10108));
  jor  g10041(.dina(n10108), .dinb(n10107), .dout(n10109));
  jand g10042(.dina(n9815), .dinb(n9697), .dout(n10110));
  jand g10043(.dina(n9824), .dinb(n9816), .dout(n10111));
  jor  g10044(.dina(n10111), .dinb(n10110), .dout(n10112));
  jand g10045(.dina(n9805), .dinb(n9700), .dout(n10113));
  jand g10046(.dina(n9814), .dinb(n9806), .dout(n10114));
  jor  g10047(.dina(n10114), .dinb(n10113), .dout(n10115));
  jand g10048(.dina(n9794), .dinb(n9786), .dout(n10116));
  jnot g10049(.din(n10116), .dout(n10117));
  jor  g10050(.dina(n9804), .dinb(n9796), .dout(n10118));
  jand g10051(.dina(n10118), .dinb(n10117), .dout(n10119));
  jnot g10052(.din(n10119), .dout(n10120));
  jand g10053(.dina(n9784), .dinb(n9714), .dout(n10121));
  jand g10054(.dina(n9785), .dinb(n9705), .dout(n10122));
  jor  g10055(.dina(n10122), .dinb(n10121), .dout(n10123));
  jor  g10056(.dina(n7061), .dinb(n3451), .dout(n10124));
  jand g10057(.dina(n5082), .dinb(n3290), .dout(n10125));
  jand g10058(.dina(n5084), .dinb(n3213), .dout(n10126));
  jor  g10059(.dina(n10126), .dinb(n10125), .dout(n10127));
  jand g10060(.dina(n6050), .dinb(n3074), .dout(n10128));
  jor  g10061(.dina(n10128), .dinb(n10127), .dout(n10129));
  jnot g10062(.din(n10129), .dout(n10130));
  jand g10063(.dina(n10130), .dinb(n10124), .dout(n10131));
  jnot g10064(.din(n10131), .dout(n10132));
  jand g10065(.dina(n9778), .dinb(n1562), .dout(n10133));
  jand g10066(.dina(n3276), .dinb(n2570), .dout(n10134));
  jand g10067(.dina(n2087), .dinb(n2117), .dout(n10135));
  jand g10068(.dina(n10135), .dinb(n895), .dout(n10136));
  jand g10069(.dina(n10136), .dinb(n2024), .dout(n10137));
  jand g10070(.dina(n10137), .dinb(n10134), .dout(n10138));
  jand g10071(.dina(n10138), .dinb(n10133), .dout(n10139));
  jand g10072(.dina(n1772), .dinb(n678), .dout(n10140));
  jand g10073(.dina(n10140), .dinb(n326), .dout(n10141));
  jand g10074(.dina(n10141), .dinb(n4576), .dout(n10142));
  jand g10075(.dina(n881), .dinb(n811), .dout(n10143));
  jand g10076(.dina(n1207), .dinb(n1283), .dout(n10144));
  jand g10077(.dina(n668), .dinb(n831), .dout(n10145));
  jand g10078(.dina(n10145), .dinb(n10144), .dout(n10146));
  jand g10079(.dina(n3840), .dinb(n1698), .dout(n10147));
  jand g10080(.dina(n10147), .dinb(n10146), .dout(n10148));
  jand g10081(.dina(n685), .dinb(n900), .dout(n10149));
  jand g10082(.dina(n10149), .dinb(n1514), .dout(n10150));
  jand g10083(.dina(n10150), .dinb(n6269), .dout(n10151));
  jand g10084(.dina(n10151), .dinb(n10148), .dout(n10152));
  jand g10085(.dina(n1367), .dinb(n135), .dout(n10153));
  jand g10086(.dina(n10153), .dinb(n4669), .dout(n10154));
  jand g10087(.dina(n10154), .dinb(n994), .dout(n10155));
  jand g10088(.dina(n10155), .dinb(n10152), .dout(n10156));
  jand g10089(.dina(n10156), .dinb(n10143), .dout(n10157));
  jand g10090(.dina(n10157), .dinb(n10142), .dout(n10158));
  jand g10091(.dina(n10158), .dinb(n10139), .dout(n10159));
  jand g10092(.dina(n699), .dinb(n1233), .dout(n10160));
  jand g10093(.dina(n452), .dinb(n1346), .dout(n10161));
  jand g10094(.dina(n10161), .dinb(n10160), .dout(n10162));
  jand g10095(.dina(n1016), .dinb(n472), .dout(n10163));
  jand g10096(.dina(n1536), .dinb(n514), .dout(n10164));
  jand g10097(.dina(n10164), .dinb(n10163), .dout(n10165));
  jand g10098(.dina(n10165), .dinb(n2526), .dout(n10166));
  jand g10099(.dina(n10166), .dinb(n10162), .dout(n10167));
  jand g10100(.dina(n1240), .dinb(n1376), .dout(n10168));
  jand g10101(.dina(n349), .dinb(n916), .dout(n10169));
  jand g10102(.dina(n10169), .dinb(n1325), .dout(n10170));
  jand g10103(.dina(n10170), .dinb(n4528), .dout(n10171));
  jand g10104(.dina(n5415), .dinb(n3264), .dout(n10172));
  jand g10105(.dina(n10172), .dinb(n5378), .dout(n10173));
  jand g10106(.dina(n10173), .dinb(n10171), .dout(n10174));
  jand g10107(.dina(n650), .dinb(n838), .dout(n10175));
  jand g10108(.dina(n10175), .dinb(n1560), .dout(n10176));
  jand g10109(.dina(n10176), .dinb(n4668), .dout(n10177));
  jand g10110(.dina(n1042), .dinb(n1316), .dout(n10178));
  jand g10111(.dina(n10178), .dinb(n1524), .dout(n10179));
  jand g10112(.dina(n10179), .dinb(n10177), .dout(n10180));
  jand g10113(.dina(n10180), .dinb(n10174), .dout(n10181));
  jand g10114(.dina(n10181), .dinb(n10168), .dout(n10182));
  jand g10115(.dina(n10182), .dinb(n10167), .dout(n10183));
  jand g10116(.dina(n10183), .dinb(n10159), .dout(n10184));
  jand g10117(.dina(n1765), .dinb(n1315), .dout(n10185));
  jand g10118(.dina(n3857), .dinb(n1592), .dout(n10186));
  jand g10119(.dina(n10186), .dinb(n3214), .dout(n10187));
  jand g10120(.dina(n10187), .dinb(n10185), .dout(n10188));
  jand g10121(.dina(n461), .dinb(n1738), .dout(n10189));
  jand g10122(.dina(n1227), .dinb(n82), .dout(n10190));
  jand g10123(.dina(n672), .dinb(n447), .dout(n10191));
  jand g10124(.dina(n10191), .dinb(n10190), .dout(n10192));
  jand g10125(.dina(n10192), .dinb(n10189), .dout(n10193));
  jand g10126(.dina(n10193), .dinb(n10188), .dout(n10194));
  jand g10127(.dina(n660), .dinb(n1260), .dout(n10195));
  jand g10128(.dina(n537), .dinb(n907), .dout(n10196));
  jand g10129(.dina(n1159), .dinb(n1575), .dout(n10197));
  jand g10130(.dina(n10197), .dinb(n10196), .dout(n10198));
  jand g10131(.dina(n600), .dinb(n2148), .dout(n10199));
  jand g10132(.dina(n10199), .dinb(n555), .dout(n10200));
  jand g10133(.dina(n10200), .dinb(n10198), .dout(n10201));
  jand g10134(.dina(n10201), .dinb(n10195), .dout(n10202));
  jand g10135(.dina(n10202), .dinb(n715), .dout(n10203));
  jand g10136(.dina(n5506), .dinb(n3322), .dout(n10204));
  jand g10137(.dina(n10204), .dinb(n1218), .dout(n10205));
  jand g10138(.dina(n1721), .dinb(n1203), .dout(n10206));
  jand g10139(.dina(n10206), .dinb(n884), .dout(n10207));
  jand g10140(.dina(n1476), .dinb(n1304), .dout(n10208));
  jand g10141(.dina(n10208), .dinb(n10207), .dout(n10209));
  jand g10142(.dina(n10209), .dinb(n172), .dout(n10210));
  jand g10143(.dina(n10210), .dinb(n10205), .dout(n10211));
  jand g10144(.dina(n2587), .dinb(n2152), .dout(n10212));
  jand g10145(.dina(n10212), .dinb(n3397), .dout(n10213));
  jand g10146(.dina(n10213), .dinb(n8383), .dout(n10214));
  jand g10147(.dina(n10214), .dinb(n10211), .dout(n10215));
  jand g10148(.dina(n10215), .dinb(n10203), .dout(n10216));
  jand g10149(.dina(n10216), .dinb(n10194), .dout(n10217));
  jand g10150(.dina(n10217), .dinb(n10184), .dout(n10218));
  jand g10151(.dina(n10218), .dinb(n9572), .dout(n10219));
  jnot g10152(.din(n10219), .dout(n10220));
  jor  g10153(.dina(n10218), .dinb(n9572), .dout(n10221));
  jand g10154(.dina(n10221), .dinb(n4713), .dout(n10222));
  jand g10155(.dina(n10222), .dinb(n10220), .dout(n10223));
  jnot g10156(.din(n10223), .dout(n10224));
  jand g10157(.dina(n10224), .dinb(n4713), .dout(n10225));
  jand g10158(.dina(n10224), .dinb(n10221), .dout(n10226));
  jand g10159(.dina(n10226), .dinb(n10220), .dout(n10227));
  jor  g10160(.dina(n10227), .dinb(n10225), .dout(n10228));
  jnot g10161(.din(n10228), .dout(n10229));
  jor  g10162(.dina(n9782), .dinb(n9573), .dout(n10230));
  jand g10163(.dina(n9783), .dinb(n9719), .dout(n10231));
  jnot g10164(.din(n10231), .dout(n10232));
  jand g10165(.dina(n10232), .dinb(n10230), .dout(n10233));
  jxor g10166(.dina(n10233), .dinb(n10229), .dout(n10234));
  jxor g10167(.dina(n10234), .dinb(n10132), .dout(n10235));
  jnot g10168(.din(n10235), .dout(n10236));
  jor  g10169(.dina(n3789), .dinb(n4343), .dout(n10237));
  jor  g10170(.dina(n3420), .dinb(n4346), .dout(n10238));
  jor  g10171(.dina(n3683), .dinb(n3286), .dout(n10239));
  jand g10172(.dina(n10239), .dinb(n10238), .dout(n10240));
  jor  g10173(.dina(n3787), .dinb(n4348), .dout(n10241));
  jand g10174(.dina(n10241), .dinb(n10240), .dout(n10242));
  jand g10175(.dina(n10242), .dinb(n10237), .dout(n10243));
  jxor g10176(.dina(n10243), .dinb(\a[29] ), .dout(n10244));
  jxor g10177(.dina(n10244), .dinb(n10236), .dout(n10245));
  jxor g10178(.dina(n10245), .dinb(n10123), .dout(n10246));
  jor  g10179(.dina(n4021), .dinb(n2303), .dout(n10247));
  jor  g10180(.dina(n3863), .dinb(n1805), .dout(n10248));
  jor  g10181(.dina(n4019), .dinb(n2309), .dout(n10249));
  jor  g10182(.dina(n3929), .dinb(n2306), .dout(n10250));
  jand g10183(.dina(n10250), .dinb(n10249), .dout(n10251));
  jand g10184(.dina(n10251), .dinb(n10248), .dout(n10252));
  jand g10185(.dina(n10252), .dinb(n10247), .dout(n10253));
  jxor g10186(.dina(n10253), .dinb(n77), .dout(n10254));
  jxor g10187(.dina(n10254), .dinb(n10246), .dout(n10255));
  jxor g10188(.dina(n10255), .dinb(n10120), .dout(n10256));
  jnot g10189(.din(n10256), .dout(n10257));
  jor  g10190(.dina(n4714), .dinb(n807), .dout(n10258));
  jor  g10191(.dina(n4596), .dinb(n1613), .dout(n10259));
  jor  g10192(.dina(n4526), .dinb(n1621), .dout(n10260));
  jand g10193(.dina(n10260), .dinb(n10259), .dout(n10261));
  jor  g10194(.dina(n4471), .dinb(n1617), .dout(n10262));
  jand g10195(.dina(n10262), .dinb(n10261), .dout(n10263));
  jand g10196(.dina(n10263), .dinb(n10258), .dout(n10264));
  jxor g10197(.dina(n10264), .dinb(\a[23] ), .dout(n10265));
  jxor g10198(.dina(n10265), .dinb(n10257), .dout(n10266));
  jxor g10199(.dina(n10266), .dinb(n10115), .dout(n10267));
  jor  g10200(.dina(n5560), .dinb(n1820), .dout(n10268));
  jor  g10201(.dina(n5264), .dinb(n2181), .dout(n10269));
  jor  g10202(.dina(n4686), .dinb(n2186), .dout(n10270));
  jor  g10203(.dina(n5422), .dinb(n2189), .dout(n10271));
  jand g10204(.dina(n10271), .dinb(n10270), .dout(n10272));
  jand g10205(.dina(n10272), .dinb(n10269), .dout(n10273));
  jand g10206(.dina(n10273), .dinb(n10268), .dout(n10274));
  jxor g10207(.dina(n10274), .dinb(n2196), .dout(n10275));
  jxor g10208(.dina(n10275), .dinb(n10267), .dout(n10276));
  jxor g10209(.dina(n10276), .dinb(n10112), .dout(n10277));
  jor  g10210(.dina(n6207), .dinb(n2744), .dout(n10278));
  jor  g10211(.dina(n5525), .dinb(n2749), .dout(n10279));
  jor  g10212(.dina(n5364), .dinb(n2758), .dout(n10280));
  jor  g10213(.dina(n6205), .dinb(n2753), .dout(n10281));
  jand g10214(.dina(n10281), .dinb(n10280), .dout(n10282));
  jand g10215(.dina(n10282), .dinb(n10279), .dout(n10283));
  jand g10216(.dina(n10283), .dinb(n10278), .dout(n10284));
  jxor g10217(.dina(n10284), .dinb(n2441), .dout(n10285));
  jxor g10218(.dina(n10285), .dinb(n10277), .dout(n10286));
  jxor g10219(.dina(n10286), .dinb(n10109), .dout(n10287));
  jor  g10220(.dina(n6491), .dinb(n3424), .dout(n10288));
  jor  g10221(.dina(n6297), .dinb(n3429), .dout(n10289));
  jor  g10222(.dina(n6390), .dinb(n3211), .dout(n10290));
  jor  g10223(.dina(n6489), .dinb(n3426), .dout(n10291));
  jand g10224(.dina(n10291), .dinb(n10290), .dout(n10292));
  jand g10225(.dina(n10292), .dinb(n10289), .dout(n10293));
  jand g10226(.dina(n10293), .dinb(n10288), .dout(n10294));
  jxor g10227(.dina(n10294), .dinb(n3473), .dout(n10295));
  jxor g10228(.dina(n10295), .dinb(n10287), .dout(n10296));
  jxor g10229(.dina(n10296), .dinb(n10106), .dout(n10297));
  jxor g10230(.dina(n10297), .dinb(n10101), .dout(n10298));
  jxor g10231(.dina(n10298), .dinb(n10089), .dout(n10299));
  jnot g10232(.din(n10299), .dout(n10300));
  jand g10233(.dina(n9857), .dinb(n9672), .dout(n10301));
  jnot g10234(.din(n10301), .dout(n10302));
  jor  g10235(.dina(n9871), .dinb(n9859), .dout(n10303));
  jand g10236(.dina(n10303), .dinb(n10302), .dout(n10304));
  jxor g10237(.dina(n10304), .dinb(n10300), .dout(n10305));
  jxor g10238(.dina(n10305), .dinb(n9872), .dout(n10306));
  jxor g10239(.dina(n10306), .dinb(n10084), .dout(n10307));
  jand g10240(.dina(n10307), .dinb(n2743), .dout(n10308));
  jand g10241(.dina(n10305), .dinb(n2752), .dout(n10309));
  jand g10242(.dina(n9872), .dinb(n2748), .dout(n10310));
  jand g10243(.dina(n9655), .dinb(n2757), .dout(n10311));
  jor  g10244(.dina(n10311), .dinb(n10310), .dout(n10312));
  jor  g10245(.dina(n10312), .dinb(n10309), .dout(n10313));
  jor  g10246(.dina(n10313), .dinb(n10308), .dout(n10314));
  jxor g10247(.dina(n10314), .dinb(n2441), .dout(n10315));
  jxor g10248(.dina(n10315), .dinb(n10081), .dout(n10316));
  jxor g10249(.dina(n10316), .dinb(n10036), .dout(n10317));
  jnot g10250(.din(n10317), .dout(n10318));
  jand g10251(.dina(n10295), .dinb(n10287), .dout(n10319));
  jand g10252(.dina(n10296), .dinb(n10106), .dout(n10320));
  jor  g10253(.dina(n10320), .dinb(n10319), .dout(n10321));
  jnot g10254(.din(n10321), .dout(n10322));
  jor  g10255(.dina(n8260), .dinb(n4023), .dout(n10323));
  jor  g10256(.dina(n7680), .dinb(n3871), .dout(n10324));
  jor  g10257(.dina(n7999), .dinb(n4028), .dout(n10325));
  jand g10258(.dina(n10325), .dinb(n10324), .dout(n10326));
  jand g10259(.dina(n10326), .dinb(n10323), .dout(n10327));
  jxor g10260(.dina(n10327), .dinb(\a[11] ), .dout(n10328));
  jor  g10261(.dina(n10328), .dinb(n10322), .dout(n10329));
  jxor g10262(.dina(n10328), .dinb(n10322), .dout(n10330));
  jand g10263(.dina(n10285), .dinb(n10277), .dout(n10331));
  jand g10264(.dina(n10286), .dinb(n10109), .dout(n10332));
  jor  g10265(.dina(n10332), .dinb(n10331), .dout(n10333));
  jand g10266(.dina(n10275), .dinb(n10267), .dout(n10334));
  jand g10267(.dina(n10276), .dinb(n10112), .dout(n10335));
  jor  g10268(.dina(n10335), .dinb(n10334), .dout(n10336));
  jor  g10269(.dina(n10265), .dinb(n10257), .dout(n10337));
  jand g10270(.dina(n10266), .dinb(n10115), .dout(n10338));
  jnot g10271(.din(n10338), .dout(n10339));
  jand g10272(.dina(n10339), .dinb(n10337), .dout(n10340));
  jnot g10273(.din(n10340), .dout(n10341));
  jand g10274(.dina(n10254), .dinb(n10246), .dout(n10342));
  jand g10275(.dina(n10255), .dinb(n10120), .dout(n10343));
  jor  g10276(.dina(n10343), .dinb(n10342), .dout(n10344));
  jor  g10277(.dina(n10244), .dinb(n10236), .dout(n10345));
  jand g10278(.dina(n10245), .dinb(n10123), .dout(n10346));
  jnot g10279(.din(n10346), .dout(n10347));
  jand g10280(.dina(n10347), .dinb(n10345), .dout(n10348));
  jnot g10281(.din(n10348), .dout(n10349));
  jor  g10282(.dina(n10233), .dinb(n10229), .dout(n10350));
  jand g10283(.dina(n10234), .dinb(n10132), .dout(n10351));
  jnot g10284(.din(n10351), .dout(n10352));
  jand g10285(.dina(n10352), .dinb(n10350), .dout(n10353));
  jnot g10286(.din(n10353), .dout(n10354));
  jor  g10287(.dina(n7061), .dinb(n3440), .dout(n10355));
  jand g10288(.dina(n6050), .dinb(n3290), .dout(n10356));
  jand g10289(.dina(n5084), .dinb(n3287), .dout(n10357));
  jor  g10290(.dina(n10357), .dinb(n10356), .dout(n10358));
  jand g10291(.dina(n5082), .dinb(n3213), .dout(n10359));
  jor  g10292(.dina(n10359), .dinb(n10358), .dout(n10360));
  jnot g10293(.din(n10360), .dout(n10361));
  jand g10294(.dina(n10361), .dinb(n10355), .dout(n10362));
  jnot g10295(.din(n10362), .dout(n10363));
  jand g10296(.dina(n848), .dinb(n838), .dout(n10364));
  jand g10297(.dina(n10364), .dinb(n2666), .dout(n10365));
  jand g10298(.dina(n10365), .dinb(n1228), .dout(n10366));
  jand g10299(.dina(n1218), .dinb(n901), .dout(n10367));
  jand g10300(.dina(n10367), .dinb(n479), .dout(n10368));
  jand g10301(.dina(n10368), .dinb(n1470), .dout(n10369));
  jand g10302(.dina(n9545), .dinb(n1327), .dout(n10370));
  jand g10303(.dina(n10370), .dinb(n10369), .dout(n10371));
  jand g10304(.dina(n10371), .dinb(n10366), .dout(n10372));
  jand g10305(.dina(n3031), .dinb(n1346), .dout(n10373));
  jand g10306(.dina(n10373), .dinb(n8128), .dout(n10374));
  jand g10307(.dina(n1167), .dinb(n430), .dout(n10375));
  jand g10308(.dina(n1693), .dinb(n893), .dout(n10376));
  jand g10309(.dina(n1037), .dinb(n1358), .dout(n10377));
  jand g10310(.dina(n10377), .dinb(n10376), .dout(n10378));
  jand g10311(.dina(n10378), .dinb(n10375), .dout(n10379));
  jand g10312(.dina(n10379), .dinb(n10374), .dout(n10380));
  jand g10313(.dina(n10380), .dinb(n10372), .dout(n10381));
  jand g10314(.dina(n1107), .dinb(n1430), .dout(n10382));
  jand g10315(.dina(n10382), .dinb(n1534), .dout(n10383));
  jand g10316(.dina(n503), .dinb(n676), .dout(n10384));
  jand g10317(.dina(n10384), .dinb(n440), .dout(n10385));
  jand g10318(.dina(n10385), .dinb(n10383), .dout(n10386));
  jand g10319(.dina(n1361), .dinb(n465), .dout(n10387));
  jand g10320(.dina(n10387), .dinb(n1822), .dout(n10388));
  jand g10321(.dina(n10388), .dinb(n1225), .dout(n10389));
  jand g10322(.dina(n1288), .dinb(n1273), .dout(n10390));
  jand g10323(.dina(n10390), .dinb(n101), .dout(n10391));
  jand g10324(.dina(n10391), .dinb(n1236), .dout(n10392));
  jand g10325(.dina(n10392), .dinb(n10389), .dout(n10393));
  jand g10326(.dina(n10393), .dinb(n10386), .dout(n10394));
  jand g10327(.dina(n10394), .dinb(n325), .dout(n10395));
  jand g10328(.dina(n10395), .dinb(n10381), .dout(n10396));
  jand g10329(.dina(n694), .dinb(n1344), .dout(n10397));
  jand g10330(.dina(n10397), .dinb(n1763), .dout(n10398));
  jand g10331(.dina(n678), .dinb(n869), .dout(n10399));
  jand g10332(.dina(n10399), .dinb(n1246), .dout(n10400));
  jand g10333(.dina(n10400), .dinb(n480), .dout(n10401));
  jand g10334(.dina(n10401), .dinb(n10398), .dout(n10402));
  jand g10335(.dina(n10402), .dinb(n3221), .dout(n10403));
  jand g10336(.dina(n932), .dinb(n510), .dout(n10404));
  jand g10337(.dina(n993), .dinb(n808), .dout(n10405));
  jand g10338(.dina(n10405), .dinb(n1433), .dout(n10406));
  jand g10339(.dina(n6439), .dinb(n683), .dout(n10407));
  jand g10340(.dina(n10407), .dinb(n10406), .dout(n10408));
  jand g10341(.dina(n1326), .dinb(n1315), .dout(n10409));
  jand g10342(.dina(n8370), .dinb(n6368), .dout(n10410));
  jand g10343(.dina(n10410), .dinb(n10409), .dout(n10411));
  jand g10344(.dina(n10411), .dinb(n10408), .dout(n10412));
  jand g10345(.dina(n680), .dinb(n1040), .dout(n10413));
  jand g10346(.dina(n7991), .dinb(n1365), .dout(n10414));
  jand g10347(.dina(n10414), .dinb(n10413), .dout(n10415));
  jand g10348(.dina(n10415), .dinb(n10412), .dout(n10416));
  jand g10349(.dina(n10416), .dinb(n10404), .dout(n10417));
  jand g10350(.dina(n10417), .dinb(n10403), .dout(n10418));
  jand g10351(.dina(n10418), .dinb(n10396), .dout(n10419));
  jand g10352(.dina(n10419), .dinb(n5347), .dout(n10420));
  jnot g10353(.din(n10420), .dout(n10421));
  jxor g10354(.dina(n10421), .dinb(n10226), .dout(n10422));
  jxor g10355(.dina(n10422), .dinb(n10363), .dout(n10423));
  jxor g10356(.dina(n10423), .dinb(n10354), .dout(n10424));
  jor  g10357(.dina(n4051), .dinb(n4343), .dout(n10425));
  jor  g10358(.dina(n3787), .dinb(n4346), .dout(n10426));
  jor  g10359(.dina(n3863), .dinb(n4348), .dout(n10427));
  jor  g10360(.dina(n3683), .dinb(n3420), .dout(n10428));
  jand g10361(.dina(n10428), .dinb(n10427), .dout(n10429));
  jand g10362(.dina(n10429), .dinb(n10426), .dout(n10430));
  jand g10363(.dina(n10430), .dinb(n10425), .dout(n10431));
  jxor g10364(.dina(n10431), .dinb(n93), .dout(n10432));
  jxor g10365(.dina(n10432), .dinb(n10424), .dout(n10433));
  jxor g10366(.dina(n10433), .dinb(n10349), .dout(n10434));
  jnot g10367(.din(n10434), .dout(n10435));
  jor  g10368(.dina(n4473), .dinb(n2303), .dout(n10436));
  jor  g10369(.dina(n4019), .dinb(n2306), .dout(n10437));
  jor  g10370(.dina(n4471), .dinb(n2309), .dout(n10438));
  jand g10371(.dina(n10438), .dinb(n10437), .dout(n10439));
  jor  g10372(.dina(n3929), .dinb(n1805), .dout(n10440));
  jand g10373(.dina(n10440), .dinb(n10439), .dout(n10441));
  jand g10374(.dina(n10441), .dinb(n10436), .dout(n10442));
  jxor g10375(.dina(n10442), .dinb(\a[26] ), .dout(n10443));
  jxor g10376(.dina(n10443), .dinb(n10435), .dout(n10444));
  jxor g10377(.dina(n10444), .dinb(n10344), .dout(n10445));
  jor  g10378(.dina(n4688), .dinb(n807), .dout(n10446));
  jor  g10379(.dina(n4526), .dinb(n1613), .dout(n10447));
  jor  g10380(.dina(n4596), .dinb(n1617), .dout(n10448));
  jor  g10381(.dina(n4686), .dinb(n1621), .dout(n10449));
  jand g10382(.dina(n10449), .dinb(n10448), .dout(n10450));
  jand g10383(.dina(n10450), .dinb(n10447), .dout(n10451));
  jand g10384(.dina(n10451), .dinb(n10446), .dout(n10452));
  jxor g10385(.dina(n10452), .dinb(n65), .dout(n10453));
  jxor g10386(.dina(n10453), .dinb(n10445), .dout(n10454));
  jxor g10387(.dina(n10454), .dinb(n10341), .dout(n10455));
  jor  g10388(.dina(n5549), .dinb(n1820), .dout(n10456));
  jor  g10389(.dina(n5422), .dinb(n2181), .dout(n10457));
  jor  g10390(.dina(n5364), .dinb(n2189), .dout(n10458));
  jor  g10391(.dina(n5264), .dinb(n2186), .dout(n10459));
  jand g10392(.dina(n10459), .dinb(n10458), .dout(n10460));
  jand g10393(.dina(n10460), .dinb(n10457), .dout(n10461));
  jand g10394(.dina(n10461), .dinb(n10456), .dout(n10462));
  jxor g10395(.dina(n10462), .dinb(n2196), .dout(n10463));
  jxor g10396(.dina(n10463), .dinb(n10455), .dout(n10464));
  jxor g10397(.dina(n10464), .dinb(n10336), .dout(n10465));
  jor  g10398(.dina(n6516), .dinb(n2744), .dout(n10466));
  jor  g10399(.dina(n6205), .dinb(n2749), .dout(n10467));
  jor  g10400(.dina(n5525), .dinb(n2758), .dout(n10468));
  jor  g10401(.dina(n6390), .dinb(n2753), .dout(n10469));
  jand g10402(.dina(n10469), .dinb(n10468), .dout(n10470));
  jand g10403(.dina(n10470), .dinb(n10467), .dout(n10471));
  jand g10404(.dina(n10471), .dinb(n10466), .dout(n10472));
  jxor g10405(.dina(n10472), .dinb(n2441), .dout(n10473));
  jxor g10406(.dina(n10473), .dinb(n10465), .dout(n10474));
  jxor g10407(.dina(n10474), .dinb(n10333), .dout(n10475));
  jnot g10408(.din(n10475), .dout(n10476));
  jor  g10409(.dina(n7301), .dinb(n3426), .dout(n10477));
  jor  g10410(.dina(n7303), .dinb(n3424), .dout(n10478));
  jor  g10411(.dina(n6297), .dinb(n3211), .dout(n10479));
  jor  g10412(.dina(n6489), .dinb(n3429), .dout(n10480));
  jand g10413(.dina(n10480), .dinb(n10479), .dout(n10481));
  jand g10414(.dina(n10481), .dinb(n10478), .dout(n10482));
  jand g10415(.dina(n10482), .dinb(n10477), .dout(n10483));
  jxor g10416(.dina(n10483), .dinb(\a[14] ), .dout(n10484));
  jxor g10417(.dina(n10484), .dinb(n10476), .dout(n10485));
  jand g10418(.dina(n10485), .dinb(n10330), .dout(n10486));
  jnot g10419(.din(n10486), .dout(n10487));
  jand g10420(.dina(n10487), .dinb(n10329), .dout(n10488));
  jnot g10421(.din(n10488), .dout(n10489));
  jand g10422(.dina(n10474), .dinb(n10333), .dout(n10490));
  jnot g10423(.din(n10490), .dout(n10491));
  jor  g10424(.dina(n10484), .dinb(n10476), .dout(n10492));
  jand g10425(.dina(n10492), .dinb(n10491), .dout(n10493));
  jand g10426(.dina(n8256), .dinb(n4022), .dout(n10494));
  jor  g10427(.dina(n10494), .dinb(n3870), .dout(n10495));
  jand g10428(.dina(n10495), .dinb(n8000), .dout(n10496));
  jxor g10429(.dina(n10496), .dinb(n4050), .dout(n10497));
  jxor g10430(.dina(n10497), .dinb(n10493), .dout(n10498));
  jand g10431(.dina(n10464), .dinb(n10336), .dout(n10499));
  jand g10432(.dina(n10473), .dinb(n10465), .dout(n10500));
  jor  g10433(.dina(n10500), .dinb(n10499), .dout(n10501));
  jand g10434(.dina(n10454), .dinb(n10341), .dout(n10502));
  jand g10435(.dina(n10463), .dinb(n10455), .dout(n10503));
  jor  g10436(.dina(n10503), .dinb(n10502), .dout(n10504));
  jand g10437(.dina(n10444), .dinb(n10344), .dout(n10505));
  jand g10438(.dina(n10453), .dinb(n10445), .dout(n10506));
  jor  g10439(.dina(n10506), .dinb(n10505), .dout(n10507));
  jand g10440(.dina(n10433), .dinb(n10349), .dout(n10508));
  jnot g10441(.din(n10508), .dout(n10509));
  jor  g10442(.dina(n10443), .dinb(n10435), .dout(n10510));
  jand g10443(.dina(n10510), .dinb(n10509), .dout(n10511));
  jnot g10444(.din(n10511), .dout(n10512));
  jand g10445(.dina(n10423), .dinb(n10354), .dout(n10513));
  jand g10446(.dina(n10432), .dinb(n10424), .dout(n10514));
  jor  g10447(.dina(n10514), .dinb(n10513), .dout(n10515));
  jand g10448(.dina(n5076), .dinb(n6704), .dout(n10516));
  jand g10449(.dina(n6050), .dinb(n3213), .dout(n10517));
  jand g10450(.dina(n5084), .dinb(n3729), .dout(n10518));
  jor  g10451(.dina(n10518), .dinb(n10517), .dout(n10519));
  jand g10452(.dina(n5082), .dinb(n3287), .dout(n10520));
  jor  g10453(.dina(n10520), .dinb(n10519), .dout(n10521));
  jor  g10454(.dina(n10521), .dinb(n10516), .dout(n10522));
  jnot g10455(.din(n10226), .dout(n10523));
  jand g10456(.dina(n10420), .dinb(n10523), .dout(n10524));
  jand g10457(.dina(n10422), .dinb(n10363), .dout(n10525));
  jor  g10458(.dina(n10525), .dinb(n10524), .dout(n10526));
  jand g10459(.dina(n1697), .dinb(n428), .dout(n10527));
  jand g10460(.dina(n10527), .dinb(n326), .dout(n10528));
  jand g10461(.dina(n10528), .dinb(n920), .dout(n10529));
  jand g10462(.dina(n983), .dinb(n537), .dout(n10530));
  jand g10463(.dina(n693), .dinb(n588), .dout(n10531));
  jand g10464(.dina(n10531), .dinb(n10530), .dout(n10532));
  jand g10465(.dina(n10532), .dinb(n10529), .dout(n10533));
  jand g10466(.dina(n848), .dinb(n1316), .dout(n10534));
  jand g10467(.dina(n10534), .dinb(n8600), .dout(n10535));
  jand g10468(.dina(n10535), .dinb(n10533), .dout(n10536));
  jand g10469(.dina(n1579), .dinb(n1569), .dout(n10537));
  jand g10470(.dina(n10537), .dinb(n504), .dout(n10538));
  jand g10471(.dina(n10538), .dinb(n10536), .dout(n10539));
  jand g10472(.dina(n4556), .dinb(n1344), .dout(n10540));
  jand g10473(.dina(n10540), .dinb(n9142), .dout(n10541));
  jand g10474(.dina(n2023), .dinb(n1053), .dout(n10542));
  jand g10475(.dina(n10542), .dinb(n430), .dout(n10543));
  jand g10476(.dina(n10543), .dinb(n10541), .dout(n10544));
  jand g10477(.dina(n10544), .dinb(n7807), .dout(n10545));
  jand g10478(.dina(n10545), .dinb(n10539), .dout(n10546));
  jand g10479(.dina(n10546), .dinb(n3246), .dout(n10547));
  jand g10480(.dina(n10547), .dinb(n4507), .dout(n10548));
  jxor g10481(.dina(n10548), .dinb(n10421), .dout(n10549));
  jor  g10482(.dina(n10549), .dinb(n10526), .dout(n10550));
  jnot g10483(.din(n10548), .dout(n10551));
  jand g10484(.dina(n10551), .dinb(n10420), .dout(n10552));
  jnot g10485(.din(n10552), .dout(n10553));
  jand g10486(.dina(n10548), .dinb(n10421), .dout(n10554));
  jnot g10487(.din(n10554), .dout(n10555));
  jand g10488(.dina(n10555), .dinb(n10526), .dout(n10556));
  jand g10489(.dina(n10556), .dinb(n10553), .dout(n10557));
  jnot g10490(.din(n10557), .dout(n10558));
  jand g10491(.dina(n10558), .dinb(n10550), .dout(n10559));
  jxor g10492(.dina(n10559), .dinb(n10522), .dout(n10560));
  jnot g10493(.din(n10560), .dout(n10561));
  jor  g10494(.dina(n4038), .dinb(n4343), .dout(n10562));
  jor  g10495(.dina(n3863), .dinb(n4346), .dout(n10563));
  jor  g10496(.dina(n3929), .dinb(n4348), .dout(n10564));
  jand g10497(.dina(n10564), .dinb(n10563), .dout(n10565));
  jor  g10498(.dina(n3787), .dinb(n3683), .dout(n10566));
  jand g10499(.dina(n10566), .dinb(n10565), .dout(n10567));
  jand g10500(.dina(n10567), .dinb(n10562), .dout(n10568));
  jxor g10501(.dina(n10568), .dinb(\a[29] ), .dout(n10569));
  jxor g10502(.dina(n10569), .dinb(n10561), .dout(n10570));
  jxor g10503(.dina(n10570), .dinb(n10515), .dout(n10571));
  jnot g10504(.din(n10571), .dout(n10572));
  jor  g10505(.dina(n4726), .dinb(n2303), .dout(n10573));
  jor  g10506(.dina(n4471), .dinb(n2306), .dout(n10574));
  jor  g10507(.dina(n4596), .dinb(n2309), .dout(n10575));
  jand g10508(.dina(n10575), .dinb(n10574), .dout(n10576));
  jor  g10509(.dina(n4019), .dinb(n1805), .dout(n10577));
  jand g10510(.dina(n10577), .dinb(n10576), .dout(n10578));
  jand g10511(.dina(n10578), .dinb(n10573), .dout(n10579));
  jxor g10512(.dina(n10579), .dinb(\a[26] ), .dout(n10580));
  jxor g10513(.dina(n10580), .dinb(n10572), .dout(n10581));
  jxor g10514(.dina(n10581), .dinb(n10512), .dout(n10582));
  jor  g10515(.dina(n5266), .dinb(n807), .dout(n10583));
  jor  g10516(.dina(n4686), .dinb(n1613), .dout(n10584));
  jor  g10517(.dina(n4526), .dinb(n1617), .dout(n10585));
  jor  g10518(.dina(n5264), .dinb(n1621), .dout(n10586));
  jand g10519(.dina(n10586), .dinb(n10585), .dout(n10587));
  jand g10520(.dina(n10587), .dinb(n10584), .dout(n10588));
  jand g10521(.dina(n10588), .dinb(n10583), .dout(n10589));
  jxor g10522(.dina(n10589), .dinb(n65), .dout(n10590));
  jxor g10523(.dina(n10590), .dinb(n10582), .dout(n10591));
  jxor g10524(.dina(n10591), .dinb(n10507), .dout(n10592));
  jor  g10525(.dina(n5527), .dinb(n1820), .dout(n10593));
  jor  g10526(.dina(n5364), .dinb(n2181), .dout(n10594));
  jor  g10527(.dina(n5422), .dinb(n2186), .dout(n10595));
  jor  g10528(.dina(n5525), .dinb(n2189), .dout(n10596));
  jand g10529(.dina(n10596), .dinb(n10595), .dout(n10597));
  jand g10530(.dina(n10597), .dinb(n10594), .dout(n10598));
  jand g10531(.dina(n10598), .dinb(n10593), .dout(n10599));
  jxor g10532(.dina(n10599), .dinb(n2196), .dout(n10600));
  jxor g10533(.dina(n10600), .dinb(n10592), .dout(n10601));
  jxor g10534(.dina(n10601), .dinb(n10504), .dout(n10602));
  jor  g10535(.dina(n6999), .dinb(n2744), .dout(n10603));
  jor  g10536(.dina(n6390), .dinb(n2749), .dout(n10604));
  jor  g10537(.dina(n6297), .dinb(n2753), .dout(n10605));
  jor  g10538(.dina(n6205), .dinb(n2758), .dout(n10606));
  jand g10539(.dina(n10606), .dinb(n10605), .dout(n10607));
  jand g10540(.dina(n10607), .dinb(n10604), .dout(n10608));
  jand g10541(.dina(n10608), .dinb(n10603), .dout(n10609));
  jxor g10542(.dina(n10609), .dinb(n2441), .dout(n10610));
  jxor g10543(.dina(n10610), .dinb(n10602), .dout(n10611));
  jxor g10544(.dina(n10611), .dinb(n10501), .dout(n10612));
  jnot g10545(.din(n10612), .dout(n10613));
  jor  g10546(.dina(n7682), .dinb(n3424), .dout(n10614));
  jor  g10547(.dina(n7301), .dinb(n3429), .dout(n10615));
  jor  g10548(.dina(n6489), .dinb(n3211), .dout(n10616));
  jand g10549(.dina(n10616), .dinb(n10615), .dout(n10617));
  jor  g10550(.dina(n7680), .dinb(n3426), .dout(n10618));
  jand g10551(.dina(n10618), .dinb(n10617), .dout(n10619));
  jand g10552(.dina(n10619), .dinb(n10614), .dout(n10620));
  jxor g10553(.dina(n10620), .dinb(\a[14] ), .dout(n10621));
  jxor g10554(.dina(n10621), .dinb(n10613), .dout(n10622));
  jxor g10555(.dina(n10622), .dinb(n10498), .dout(n10623));
  jxor g10556(.dina(n10623), .dinb(n10489), .dout(n10624));
  jnot g10557(.din(n10624), .dout(n10625));
  jand g10558(.dina(n10100), .dinb(n10092), .dout(n10626));
  jand g10559(.dina(n10297), .dinb(n10101), .dout(n10627));
  jor  g10560(.dina(n10627), .dinb(n10626), .dout(n10628));
  jxor g10561(.dina(n10485), .dinb(n10330), .dout(n10629));
  jand g10562(.dina(n10629), .dinb(n10628), .dout(n10630));
  jnot g10563(.din(n10630), .dout(n10631));
  jand g10564(.dina(n10298), .dinb(n10089), .dout(n10632));
  jnot g10565(.din(n10632), .dout(n10633));
  jor  g10566(.dina(n10304), .dinb(n10300), .dout(n10634));
  jand g10567(.dina(n10634), .dinb(n10633), .dout(n10635));
  jxor g10568(.dina(n10629), .dinb(n10628), .dout(n10636));
  jnot g10569(.din(n10636), .dout(n10637));
  jor  g10570(.dina(n10637), .dinb(n10635), .dout(n10638));
  jand g10571(.dina(n10638), .dinb(n10631), .dout(n10639));
  jxor g10572(.dina(n10639), .dinb(n10625), .dout(n10640));
  jand g10573(.dina(n9654), .dinb(n9470), .dout(n10641));
  jor  g10574(.dina(n10641), .dinb(n9860), .dout(n10642));
  jand g10575(.dina(n10642), .dinb(n9858), .dout(n10643));
  jor  g10576(.dina(n10643), .dinb(n10301), .dout(n10644));
  jand g10577(.dina(n10644), .dinb(n10299), .dout(n10645));
  jor  g10578(.dina(n10645), .dinb(n10632), .dout(n10646));
  jxor g10579(.dina(n10636), .dinb(n10646), .dout(n10647));
  jand g10580(.dina(n10647), .dinb(n10640), .dout(n10648));
  jand g10581(.dina(n10647), .dinb(n10305), .dout(n10649));
  jand g10582(.dina(n10305), .dinb(n9872), .dout(n10650));
  jand g10583(.dina(n10306), .dinb(n10084), .dout(n10651));
  jor  g10584(.dina(n10651), .dinb(n10650), .dout(n10652));
  jxor g10585(.dina(n10647), .dinb(n10305), .dout(n10653));
  jand g10586(.dina(n10653), .dinb(n10652), .dout(n10654));
  jor  g10587(.dina(n10654), .dinb(n10649), .dout(n10655));
  jxor g10588(.dina(n10647), .dinb(n10640), .dout(n10656));
  jand g10589(.dina(n10656), .dinb(n10655), .dout(n10657));
  jor  g10590(.dina(n10657), .dinb(n10648), .dout(n10658));
  jand g10591(.dina(n10623), .dinb(n10489), .dout(n10659));
  jand g10592(.dina(n10636), .dinb(n10646), .dout(n10660));
  jor  g10593(.dina(n10660), .dinb(n10630), .dout(n10661));
  jand g10594(.dina(n10661), .dinb(n10624), .dout(n10662));
  jor  g10595(.dina(n10662), .dinb(n10659), .dout(n10663));
  jor  g10596(.dina(n10497), .dinb(n10493), .dout(n10664));
  jand g10597(.dina(n10622), .dinb(n10498), .dout(n10665));
  jnot g10598(.din(n10665), .dout(n10666));
  jand g10599(.dina(n10666), .dinb(n10664), .dout(n10667));
  jnot g10600(.din(n10667), .dout(n10668));
  jand g10601(.dina(n10601), .dinb(n10504), .dout(n10669));
  jand g10602(.dina(n10610), .dinb(n10602), .dout(n10670));
  jor  g10603(.dina(n10670), .dinb(n10669), .dout(n10671));
  jand g10604(.dina(n10591), .dinb(n10507), .dout(n10672));
  jand g10605(.dina(n10600), .dinb(n10592), .dout(n10673));
  jor  g10606(.dina(n10673), .dinb(n10672), .dout(n10674));
  jand g10607(.dina(n10581), .dinb(n10512), .dout(n10675));
  jand g10608(.dina(n10590), .dinb(n10582), .dout(n10676));
  jor  g10609(.dina(n10676), .dinb(n10675), .dout(n10677));
  jand g10610(.dina(n10570), .dinb(n10515), .dout(n10678));
  jnot g10611(.din(n10678), .dout(n10679));
  jor  g10612(.dina(n10580), .dinb(n10572), .dout(n10680));
  jand g10613(.dina(n10680), .dinb(n10679), .dout(n10681));
  jnot g10614(.din(n10681), .dout(n10682));
  jand g10615(.dina(n10559), .dinb(n10522), .dout(n10683));
  jnot g10616(.din(n10683), .dout(n10684));
  jor  g10617(.dina(n10569), .dinb(n10561), .dout(n10685));
  jand g10618(.dina(n10685), .dinb(n10684), .dout(n10686));
  jnot g10619(.din(n10686), .dout(n10687));
  jor  g10620(.dina(n10556), .dinb(n10552), .dout(n10688));
  jand g10621(.dina(n1167), .dinb(n1227), .dout(n10689));
  jand g10622(.dina(n10689), .dinb(n2386), .dout(n10690));
  jand g10623(.dina(n1205), .dinb(n100), .dout(n10691));
  jand g10624(.dina(n10691), .dinb(n3026), .dout(n10692));
  jand g10625(.dina(n10692), .dinb(n10690), .dout(n10693));
  jand g10626(.dina(n9527), .dinb(n1779), .dout(n10694));
  jand g10627(.dina(n10694), .dinb(n10693), .dout(n10695));
  jand g10628(.dina(n1524), .dinb(n703), .dout(n10696));
  jand g10629(.dina(n660), .dinb(n716), .dout(n10697));
  jand g10630(.dina(n10697), .dinb(n10696), .dout(n10698));
  jand g10631(.dina(n978), .dinb(n895), .dout(n10699));
  jand g10632(.dina(n10699), .dinb(n1753), .dout(n10700));
  jand g10633(.dina(n10700), .dinb(n10698), .dout(n10701));
  jand g10634(.dina(n10701), .dinb(n1702), .dout(n10702));
  jand g10635(.dina(n10702), .dinb(n10695), .dout(n10703));
  jand g10636(.dina(n10703), .dinb(n4634), .dout(n10704));
  jand g10637(.dina(n10704), .dinb(n8124), .dout(n10705));
  jand g10638(.dina(n8820), .dinb(n467), .dout(n10706));
  jand g10639(.dina(n10706), .dinb(n3766), .dout(n10707));
  jand g10640(.dina(n829), .dinb(n654), .dout(n10708));
  jand g10641(.dina(n1228), .dinb(n178), .dout(n10709));
  jand g10642(.dina(n10709), .dinb(n10708), .dout(n10710));
  jand g10643(.dina(n9522), .dinb(n6196), .dout(n10711));
  jand g10644(.dina(n10711), .dinb(n10710), .dout(n10712));
  jand g10645(.dina(n10712), .dinb(n5492), .dout(n10713));
  jand g10646(.dina(n10713), .dinb(n10707), .dout(n10714));
  jand g10647(.dina(n901), .dinb(n1260), .dout(n10715));
  jand g10648(.dina(n1189), .dinb(n848), .dout(n10716));
  jand g10649(.dina(n10716), .dinb(n10715), .dout(n10717));
  jand g10650(.dina(n662), .dinb(n114), .dout(n10718));
  jand g10651(.dina(n10718), .dinb(n9358), .dout(n10719));
  jand g10652(.dina(n10719), .dinb(n10717), .dout(n10720));
  jand g10653(.dina(n514), .dinb(n445), .dout(n10721));
  jand g10654(.dina(n10721), .dinb(n3324), .dout(n10722));
  jand g10655(.dina(n10722), .dinb(n4668), .dout(n10723));
  jand g10656(.dina(n10723), .dinb(n10720), .dout(n10724));
  jand g10657(.dina(n10724), .dinb(n3954), .dout(n10725));
  jand g10658(.dina(n10725), .dinb(n10714), .dout(n10726));
  jand g10659(.dina(n10726), .dinb(n10416), .dout(n10727));
  jand g10660(.dina(n10727), .dinb(n10705), .dout(n10728));
  jand g10661(.dina(n1429), .dinb(n168), .dout(n10729));
  jand g10662(.dina(n10729), .dinb(n1533), .dout(n10730));
  jand g10663(.dina(n3356), .dinb(n453), .dout(n10731));
  jand g10664(.dina(n2154), .dinb(n479), .dout(n10732));
  jand g10665(.dina(n1915), .dinb(n495), .dout(n10733));
  jand g10666(.dina(n10733), .dinb(n1427), .dout(n10734));
  jand g10667(.dina(n10734), .dinb(n10732), .dout(n10735));
  jand g10668(.dina(n2367), .dinb(n1308), .dout(n10736));
  jand g10669(.dina(n1577), .dinb(n893), .dout(n10737));
  jand g10670(.dina(n1316), .dinb(n1213), .dout(n10738));
  jand g10671(.dina(n10738), .dinb(n10737), .dout(n10739));
  jand g10672(.dina(n1731), .dinb(n472), .dout(n10740));
  jand g10673(.dina(n10740), .dinb(n10739), .dout(n10741));
  jand g10674(.dina(n10741), .dinb(n10736), .dout(n10742));
  jand g10675(.dina(n10742), .dinb(n10735), .dout(n10743));
  jand g10676(.dina(n10743), .dinb(n10731), .dout(n10744));
  jand g10677(.dina(n10744), .dinb(n10730), .dout(n10745));
  jand g10678(.dina(n10745), .dinb(n10728), .dout(n10746));
  jand g10679(.dina(n10746), .dinb(n10420), .dout(n10747));
  jnot g10680(.din(n10747), .dout(n10748));
  jor  g10681(.dina(n10746), .dinb(n10420), .dout(n10749));
  jand g10682(.dina(n10749), .dinb(n4050), .dout(n10750));
  jand g10683(.dina(n10750), .dinb(n10748), .dout(n10751));
  jnot g10684(.din(n10751), .dout(n10752));
  jand g10685(.dina(n10752), .dinb(n4050), .dout(n10753));
  jand g10686(.dina(n10752), .dinb(n10749), .dout(n10754));
  jand g10687(.dina(n10754), .dinb(n10748), .dout(n10755));
  jor  g10688(.dina(n10755), .dinb(n10753), .dout(n10756));
  jnot g10689(.din(n10756), .dout(n10757));
  jor  g10690(.dina(n7061), .dinb(n3789), .dout(n10758));
  jand g10691(.dina(n5082), .dinb(n3729), .dout(n10759));
  jand g10692(.dina(n6050), .dinb(n3287), .dout(n10760));
  jor  g10693(.dina(n10760), .dinb(n10759), .dout(n10761));
  jand g10694(.dina(n5084), .dinb(n3933), .dout(n10762));
  jor  g10695(.dina(n10762), .dinb(n10761), .dout(n10763));
  jnot g10696(.din(n10763), .dout(n10764));
  jand g10697(.dina(n10764), .dinb(n10758), .dout(n10765));
  jxor g10698(.dina(n10765), .dinb(n10757), .dout(n10766));
  jxor g10699(.dina(n10766), .dinb(n10688), .dout(n10767));
  jxor g10700(.dina(n10767), .dinb(n10687), .dout(n10768));
  jor  g10701(.dina(n4021), .dinb(n4343), .dout(n10769));
  jor  g10702(.dina(n3863), .dinb(n3683), .dout(n10770));
  jor  g10703(.dina(n4019), .dinb(n4348), .dout(n10771));
  jor  g10704(.dina(n3929), .dinb(n4346), .dout(n10772));
  jand g10705(.dina(n10772), .dinb(n10771), .dout(n10773));
  jand g10706(.dina(n10773), .dinb(n10770), .dout(n10774));
  jand g10707(.dina(n10774), .dinb(n10769), .dout(n10775));
  jxor g10708(.dina(n10775), .dinb(n93), .dout(n10776));
  jxor g10709(.dina(n10776), .dinb(n10768), .dout(n10777));
  jnot g10710(.din(n10777), .dout(n10778));
  jor  g10711(.dina(n4714), .dinb(n2303), .dout(n10779));
  jor  g10712(.dina(n4596), .dinb(n2306), .dout(n10780));
  jor  g10713(.dina(n4471), .dinb(n1805), .dout(n10781));
  jand g10714(.dina(n10781), .dinb(n10780), .dout(n10782));
  jor  g10715(.dina(n4526), .dinb(n2309), .dout(n10783));
  jand g10716(.dina(n10783), .dinb(n10782), .dout(n10784));
  jand g10717(.dina(n10784), .dinb(n10779), .dout(n10785));
  jxor g10718(.dina(n10785), .dinb(\a[26] ), .dout(n10786));
  jxor g10719(.dina(n10786), .dinb(n10778), .dout(n10787));
  jxor g10720(.dina(n10787), .dinb(n10682), .dout(n10788));
  jnot g10721(.din(n10788), .dout(n10789));
  jor  g10722(.dina(n5560), .dinb(n807), .dout(n10790));
  jor  g10723(.dina(n5264), .dinb(n1613), .dout(n10791));
  jor  g10724(.dina(n5422), .dinb(n1621), .dout(n10792));
  jand g10725(.dina(n10792), .dinb(n10791), .dout(n10793));
  jor  g10726(.dina(n4686), .dinb(n1617), .dout(n10794));
  jand g10727(.dina(n10794), .dinb(n10793), .dout(n10795));
  jand g10728(.dina(n10795), .dinb(n10790), .dout(n10796));
  jxor g10729(.dina(n10796), .dinb(\a[23] ), .dout(n10797));
  jxor g10730(.dina(n10797), .dinb(n10789), .dout(n10798));
  jxor g10731(.dina(n10798), .dinb(n10677), .dout(n10799));
  jor  g10732(.dina(n6207), .dinb(n1820), .dout(n10800));
  jor  g10733(.dina(n5525), .dinb(n2181), .dout(n10801));
  jor  g10734(.dina(n5364), .dinb(n2186), .dout(n10802));
  jor  g10735(.dina(n6205), .dinb(n2189), .dout(n10803));
  jand g10736(.dina(n10803), .dinb(n10802), .dout(n10804));
  jand g10737(.dina(n10804), .dinb(n10801), .dout(n10805));
  jand g10738(.dina(n10805), .dinb(n10800), .dout(n10806));
  jxor g10739(.dina(n10806), .dinb(n2196), .dout(n10807));
  jxor g10740(.dina(n10807), .dinb(n10799), .dout(n10808));
  jxor g10741(.dina(n10808), .dinb(n10674), .dout(n10809));
  jor  g10742(.dina(n6491), .dinb(n2744), .dout(n10810));
  jor  g10743(.dina(n6297), .dinb(n2749), .dout(n10811));
  jor  g10744(.dina(n6390), .dinb(n2758), .dout(n10812));
  jor  g10745(.dina(n6489), .dinb(n2753), .dout(n10813));
  jand g10746(.dina(n10813), .dinb(n10812), .dout(n10814));
  jand g10747(.dina(n10814), .dinb(n10811), .dout(n10815));
  jand g10748(.dina(n10815), .dinb(n10810), .dout(n10816));
  jxor g10749(.dina(n10816), .dinb(n2441), .dout(n10817));
  jxor g10750(.dina(n10817), .dinb(n10809), .dout(n10818));
  jxor g10751(.dina(n10818), .dinb(n10671), .dout(n10819));
  jand g10752(.dina(n10611), .dinb(n10501), .dout(n10820));
  jnot g10753(.din(n10820), .dout(n10821));
  jor  g10754(.dina(n10621), .dinb(n10613), .dout(n10822));
  jand g10755(.dina(n10822), .dinb(n10821), .dout(n10823));
  jnot g10756(.din(n10823), .dout(n10824));
  jor  g10757(.dina(n8002), .dinb(n3424), .dout(n10825));
  jor  g10758(.dina(n7301), .dinb(n3211), .dout(n10826));
  jor  g10759(.dina(n7999), .dinb(n3426), .dout(n10827));
  jor  g10760(.dina(n7680), .dinb(n3429), .dout(n10828));
  jand g10761(.dina(n10828), .dinb(n10827), .dout(n10829));
  jand g10762(.dina(n10829), .dinb(n10826), .dout(n10830));
  jand g10763(.dina(n10830), .dinb(n10825), .dout(n10831));
  jxor g10764(.dina(n10831), .dinb(n3473), .dout(n10832));
  jxor g10765(.dina(n10832), .dinb(n10824), .dout(n10833));
  jxor g10766(.dina(n10833), .dinb(n10819), .dout(n10834));
  jxor g10767(.dina(n10834), .dinb(n10668), .dout(n10835));
  jxor g10768(.dina(n10835), .dinb(n10663), .dout(n10836));
  jxor g10769(.dina(n10836), .dinb(n10640), .dout(n10837));
  jxor g10770(.dina(n10837), .dinb(n10658), .dout(n10838));
  jand g10771(.dina(n10838), .dinb(n3423), .dout(n10839));
  jand g10772(.dina(n10836), .dinb(n3569), .dout(n10840));
  jand g10773(.dina(n10640), .dinb(n3428), .dout(n10841));
  jand g10774(.dina(n10647), .dinb(n3210), .dout(n10842));
  jor  g10775(.dina(n10842), .dinb(n10841), .dout(n10843));
  jor  g10776(.dina(n10843), .dinb(n10840), .dout(n10844));
  jor  g10777(.dina(n10844), .dinb(n10839), .dout(n10845));
  jxor g10778(.dina(n10845), .dinb(n3473), .dout(n10846));
  jor  g10779(.dina(n10846), .dinb(n10318), .dout(n10847));
  jxor g10780(.dina(n10032), .dinb(n10031), .dout(n10848));
  jnot g10781(.din(n10848), .dout(n10849));
  jxor g10782(.dina(n10656), .dinb(n10655), .dout(n10850));
  jand g10783(.dina(n10850), .dinb(n3423), .dout(n10851));
  jand g10784(.dina(n10640), .dinb(n3569), .dout(n10852));
  jand g10785(.dina(n10647), .dinb(n3428), .dout(n10853));
  jand g10786(.dina(n10305), .dinb(n3210), .dout(n10854));
  jor  g10787(.dina(n10854), .dinb(n10853), .dout(n10855));
  jor  g10788(.dina(n10855), .dinb(n10852), .dout(n10856));
  jor  g10789(.dina(n10856), .dinb(n10851), .dout(n10857));
  jxor g10790(.dina(n10857), .dinb(n3473), .dout(n10858));
  jor  g10791(.dina(n10858), .dinb(n10849), .dout(n10859));
  jxor g10792(.dina(n10027), .dinb(n10026), .dout(n10860));
  jnot g10793(.din(n10860), .dout(n10861));
  jxor g10794(.dina(n10653), .dinb(n10652), .dout(n10862));
  jand g10795(.dina(n10862), .dinb(n3423), .dout(n10863));
  jand g10796(.dina(n10647), .dinb(n3569), .dout(n10864));
  jand g10797(.dina(n10305), .dinb(n3428), .dout(n10865));
  jand g10798(.dina(n9872), .dinb(n3210), .dout(n10866));
  jor  g10799(.dina(n10866), .dinb(n10865), .dout(n10867));
  jor  g10800(.dina(n10867), .dinb(n10864), .dout(n10868));
  jor  g10801(.dina(n10868), .dinb(n10863), .dout(n10869));
  jxor g10802(.dina(n10869), .dinb(n3473), .dout(n10870));
  jor  g10803(.dina(n10870), .dinb(n10861), .dout(n10871));
  jxor g10804(.dina(n10022), .dinb(n10021), .dout(n10872));
  jand g10805(.dina(n10307), .dinb(n3423), .dout(n10873));
  jand g10806(.dina(n10305), .dinb(n3569), .dout(n10874));
  jand g10807(.dina(n9872), .dinb(n3428), .dout(n10875));
  jand g10808(.dina(n9655), .dinb(n3210), .dout(n10876));
  jor  g10809(.dina(n10876), .dinb(n10875), .dout(n10877));
  jor  g10810(.dina(n10877), .dinb(n10874), .dout(n10878));
  jor  g10811(.dina(n10878), .dinb(n10873), .dout(n10879));
  jxor g10812(.dina(n10879), .dinb(\a[14] ), .dout(n10880));
  jand g10813(.dina(n10880), .dinb(n10872), .dout(n10881));
  jxor g10814(.dina(n10017), .dinb(n10016), .dout(n10882));
  jnot g10815(.din(n10882), .dout(n10883));
  jand g10816(.dina(n9874), .dinb(n3423), .dout(n10884));
  jand g10817(.dina(n9655), .dinb(n3428), .dout(n10885));
  jand g10818(.dina(n9872), .dinb(n3569), .dout(n10886));
  jor  g10819(.dina(n10886), .dinb(n10885), .dout(n10887));
  jand g10820(.dina(n9656), .dinb(n3210), .dout(n10888));
  jor  g10821(.dina(n10888), .dinb(n10887), .dout(n10889));
  jor  g10822(.dina(n10889), .dinb(n10884), .dout(n10890));
  jxor g10823(.dina(n10890), .dinb(n3473), .dout(n10891));
  jor  g10824(.dina(n10891), .dinb(n10883), .dout(n10892));
  jxor g10825(.dina(n10012), .dinb(n10011), .dout(n10893));
  jnot g10826(.din(n10893), .dout(n10894));
  jand g10827(.dina(n9886), .dinb(n3423), .dout(n10895));
  jand g10828(.dina(n9656), .dinb(n3428), .dout(n10896));
  jand g10829(.dina(n9655), .dinb(n3569), .dout(n10897));
  jor  g10830(.dina(n10897), .dinb(n10896), .dout(n10898));
  jand g10831(.dina(n9250), .dinb(n3210), .dout(n10899));
  jor  g10832(.dina(n10899), .dinb(n10898), .dout(n10900));
  jor  g10833(.dina(n10900), .dinb(n10895), .dout(n10901));
  jxor g10834(.dina(n10901), .dinb(n3473), .dout(n10902));
  jor  g10835(.dina(n10902), .dinb(n10894), .dout(n10903));
  jxor g10836(.dina(n10007), .dinb(n10006), .dout(n10904));
  jnot g10837(.din(n10904), .dout(n10905));
  jand g10838(.dina(n9898), .dinb(n3423), .dout(n10906));
  jand g10839(.dina(n9656), .dinb(n3569), .dout(n10907));
  jand g10840(.dina(n9250), .dinb(n3428), .dout(n10908));
  jand g10841(.dina(n8936), .dinb(n3210), .dout(n10909));
  jor  g10842(.dina(n10909), .dinb(n10908), .dout(n10910));
  jor  g10843(.dina(n10910), .dinb(n10907), .dout(n10911));
  jor  g10844(.dina(n10911), .dinb(n10906), .dout(n10912));
  jxor g10845(.dina(n10912), .dinb(n3473), .dout(n10913));
  jor  g10846(.dina(n10913), .dinb(n10905), .dout(n10914));
  jxor g10847(.dina(n10004), .dinb(n10003), .dout(n10915));
  jnot g10848(.din(n10915), .dout(n10916));
  jand g10849(.dina(n9252), .dinb(n3423), .dout(n10917));
  jand g10850(.dina(n9250), .dinb(n3569), .dout(n10918));
  jand g10851(.dina(n8936), .dinb(n3428), .dout(n10919));
  jand g10852(.dina(n8723), .dinb(n3210), .dout(n10920));
  jor  g10853(.dina(n10920), .dinb(n10919), .dout(n10921));
  jor  g10854(.dina(n10921), .dinb(n10918), .dout(n10922));
  jor  g10855(.dina(n10922), .dinb(n10917), .dout(n10923));
  jxor g10856(.dina(n10923), .dinb(n3473), .dout(n10924));
  jor  g10857(.dina(n10924), .dinb(n10916), .dout(n10925));
  jxor g10858(.dina(n9999), .dinb(n9998), .dout(n10926));
  jnot g10859(.din(n10926), .dout(n10927));
  jand g10860(.dina(n8938), .dinb(n3423), .dout(n10928));
  jand g10861(.dina(n8723), .dinb(n3428), .dout(n10929));
  jand g10862(.dina(n8936), .dinb(n3569), .dout(n10930));
  jor  g10863(.dina(n10930), .dinb(n10929), .dout(n10931));
  jand g10864(.dina(n8740), .dinb(n3210), .dout(n10932));
  jor  g10865(.dina(n10932), .dinb(n10931), .dout(n10933));
  jor  g10866(.dina(n10933), .dinb(n10928), .dout(n10934));
  jxor g10867(.dina(n10934), .dinb(n3473), .dout(n10935));
  jor  g10868(.dina(n10935), .dinb(n10927), .dout(n10936));
  jxor g10869(.dina(n9995), .dinb(n9987), .dout(n10937));
  jnot g10870(.din(n10937), .dout(n10938));
  jand g10871(.dina(n8950), .dinb(n3423), .dout(n10939));
  jand g10872(.dina(n8723), .dinb(n3569), .dout(n10940));
  jand g10873(.dina(n8740), .dinb(n3428), .dout(n10941));
  jand g10874(.dina(n8268), .dinb(n3210), .dout(n10942));
  jor  g10875(.dina(n10942), .dinb(n10941), .dout(n10943));
  jor  g10876(.dina(n10943), .dinb(n10940), .dout(n10944));
  jor  g10877(.dina(n10944), .dinb(n10939), .dout(n10945));
  jxor g10878(.dina(n10945), .dinb(n3473), .dout(n10946));
  jor  g10879(.dina(n10946), .dinb(n10938), .dout(n10947));
  jor  g10880(.dina(n9974), .dinb(n2441), .dout(n10948));
  jxor g10881(.dina(n10948), .dinb(n9982), .dout(n10949));
  jand g10882(.dina(n8962), .dinb(n3423), .dout(n10950));
  jand g10883(.dina(n8740), .dinb(n3569), .dout(n10951));
  jand g10884(.dina(n8268), .dinb(n3428), .dout(n10952));
  jand g10885(.dina(n8022), .dinb(n3210), .dout(n10953));
  jor  g10886(.dina(n10953), .dinb(n10952), .dout(n10954));
  jor  g10887(.dina(n10954), .dinb(n10951), .dout(n10955));
  jor  g10888(.dina(n10955), .dinb(n10950), .dout(n10956));
  jxor g10889(.dina(n10956), .dinb(\a[14] ), .dout(n10957));
  jand g10890(.dina(n10957), .dinb(n10949), .dout(n10958));
  jand g10891(.dina(n9971), .dinb(\a[17] ), .dout(n10959));
  jxor g10892(.dina(n10959), .dinb(n9969), .dout(n10960));
  jnot g10893(.din(n10960), .dout(n10961));
  jand g10894(.dina(n8270), .dinb(n3423), .dout(n10962));
  jand g10895(.dina(n8022), .dinb(n3428), .dout(n10963));
  jand g10896(.dina(n8268), .dinb(n3569), .dout(n10964));
  jor  g10897(.dina(n10964), .dinb(n10963), .dout(n10965));
  jand g10898(.dina(n7692), .dinb(n3210), .dout(n10966));
  jor  g10899(.dina(n10966), .dinb(n10965), .dout(n10967));
  jor  g10900(.dina(n10967), .dinb(n10962), .dout(n10968));
  jxor g10901(.dina(n10968), .dinb(n3473), .dout(n10969));
  jor  g10902(.dina(n10969), .dinb(n10961), .dout(n10970));
  jand g10903(.dina(n7315), .dinb(n3423), .dout(n10971));
  jand g10904(.dina(n7019), .dinb(n3428), .dout(n10972));
  jand g10905(.dina(n7313), .dinb(n3569), .dout(n10973));
  jor  g10906(.dina(n10973), .dinb(n10972), .dout(n10974));
  jor  g10907(.dina(n10974), .dinb(n10971), .dout(n10975));
  jnot g10908(.din(n10975), .dout(n10976));
  jand g10909(.dina(n7019), .dinb(n3205), .dout(n10977));
  jnot g10910(.din(n10977), .dout(n10978));
  jand g10911(.dina(n10978), .dinb(\a[14] ), .dout(n10979));
  jand g10912(.dina(n10979), .dinb(n10976), .dout(n10980));
  jand g10913(.dina(n7693), .dinb(n3423), .dout(n10981));
  jand g10914(.dina(n7313), .dinb(n3428), .dout(n10982));
  jand g10915(.dina(n7692), .dinb(n3569), .dout(n10983));
  jor  g10916(.dina(n10983), .dinb(n10982), .dout(n10984));
  jand g10917(.dina(n7019), .dinb(n3210), .dout(n10985));
  jor  g10918(.dina(n10985), .dinb(n10984), .dout(n10986));
  jor  g10919(.dina(n10986), .dinb(n10981), .dout(n10987));
  jnot g10920(.din(n10987), .dout(n10988));
  jand g10921(.dina(n10988), .dinb(n10980), .dout(n10989));
  jand g10922(.dina(n10989), .dinb(n9971), .dout(n10990));
  jnot g10923(.din(n10990), .dout(n10991));
  jxor g10924(.dina(n10989), .dinb(n9971), .dout(n10992));
  jnot g10925(.din(n10992), .dout(n10993));
  jand g10926(.dina(n8029), .dinb(n3423), .dout(n10994));
  jand g10927(.dina(n8022), .dinb(n3569), .dout(n10995));
  jand g10928(.dina(n7313), .dinb(n3210), .dout(n10996));
  jand g10929(.dina(n7692), .dinb(n3428), .dout(n10997));
  jor  g10930(.dina(n10997), .dinb(n10996), .dout(n10998));
  jor  g10931(.dina(n10998), .dinb(n10995), .dout(n10999));
  jor  g10932(.dina(n10999), .dinb(n10994), .dout(n11000));
  jxor g10933(.dina(n11000), .dinb(n3473), .dout(n11001));
  jor  g10934(.dina(n11001), .dinb(n10993), .dout(n11002));
  jand g10935(.dina(n11002), .dinb(n10991), .dout(n11003));
  jnot g10936(.din(n11003), .dout(n11004));
  jxor g10937(.dina(n10969), .dinb(n10961), .dout(n11005));
  jand g10938(.dina(n11005), .dinb(n11004), .dout(n11006));
  jnot g10939(.din(n11006), .dout(n11007));
  jand g10940(.dina(n11007), .dinb(n10970), .dout(n11008));
  jnot g10941(.din(n11008), .dout(n11009));
  jxor g10942(.dina(n10957), .dinb(n10949), .dout(n11010));
  jand g10943(.dina(n11010), .dinb(n11009), .dout(n11011));
  jor  g10944(.dina(n11011), .dinb(n10958), .dout(n11012));
  jxor g10945(.dina(n10946), .dinb(n10938), .dout(n11013));
  jand g10946(.dina(n11013), .dinb(n11012), .dout(n11014));
  jnot g10947(.din(n11014), .dout(n11015));
  jand g10948(.dina(n11015), .dinb(n10947), .dout(n11016));
  jnot g10949(.din(n11016), .dout(n11017));
  jxor g10950(.dina(n10935), .dinb(n10927), .dout(n11018));
  jand g10951(.dina(n11018), .dinb(n11017), .dout(n11019));
  jnot g10952(.din(n11019), .dout(n11020));
  jand g10953(.dina(n11020), .dinb(n10936), .dout(n11021));
  jnot g10954(.din(n11021), .dout(n11022));
  jxor g10955(.dina(n10924), .dinb(n10916), .dout(n11023));
  jand g10956(.dina(n11023), .dinb(n11022), .dout(n11024));
  jnot g10957(.din(n11024), .dout(n11025));
  jand g10958(.dina(n11025), .dinb(n10925), .dout(n11026));
  jnot g10959(.din(n11026), .dout(n11027));
  jxor g10960(.dina(n10913), .dinb(n10905), .dout(n11028));
  jand g10961(.dina(n11028), .dinb(n11027), .dout(n11029));
  jnot g10962(.din(n11029), .dout(n11030));
  jand g10963(.dina(n11030), .dinb(n10914), .dout(n11031));
  jnot g10964(.din(n11031), .dout(n11032));
  jxor g10965(.dina(n10902), .dinb(n10894), .dout(n11033));
  jand g10966(.dina(n11033), .dinb(n11032), .dout(n11034));
  jnot g10967(.din(n11034), .dout(n11035));
  jand g10968(.dina(n11035), .dinb(n10903), .dout(n11036));
  jnot g10969(.din(n11036), .dout(n11037));
  jxor g10970(.dina(n10891), .dinb(n10883), .dout(n11038));
  jand g10971(.dina(n11038), .dinb(n11037), .dout(n11039));
  jnot g10972(.din(n11039), .dout(n11040));
  jand g10973(.dina(n11040), .dinb(n10892), .dout(n11041));
  jnot g10974(.din(n11041), .dout(n11042));
  jxor g10975(.dina(n10880), .dinb(n10872), .dout(n11043));
  jand g10976(.dina(n11043), .dinb(n11042), .dout(n11044));
  jor  g10977(.dina(n11044), .dinb(n10881), .dout(n11045));
  jxor g10978(.dina(n10870), .dinb(n10861), .dout(n11046));
  jand g10979(.dina(n11046), .dinb(n11045), .dout(n11047));
  jnot g10980(.din(n11047), .dout(n11048));
  jand g10981(.dina(n11048), .dinb(n10871), .dout(n11049));
  jnot g10982(.din(n11049), .dout(n11050));
  jxor g10983(.dina(n10858), .dinb(n10849), .dout(n11051));
  jand g10984(.dina(n11051), .dinb(n11050), .dout(n11052));
  jnot g10985(.din(n11052), .dout(n11053));
  jand g10986(.dina(n11053), .dinb(n10859), .dout(n11054));
  jxor g10987(.dina(n10846), .dinb(n10318), .dout(n11055));
  jnot g10988(.din(n11055), .dout(n11056));
  jor  g10989(.dina(n11056), .dinb(n11054), .dout(n11057));
  jand g10990(.dina(n11057), .dinb(n10847), .dout(n11058));
  jor  g10991(.dina(n10315), .dinb(n10081), .dout(n11059));
  jand g10992(.dina(n10316), .dinb(n10036), .dout(n11060));
  jnot g10993(.din(n11060), .dout(n11061));
  jand g10994(.dina(n11061), .dinb(n11059), .dout(n11062));
  jnot g10995(.din(n11062), .dout(n11063));
  jor  g10996(.dina(n10078), .dinb(n10070), .dout(n11064));
  jand g10997(.dina(n10079), .dinb(n10041), .dout(n11065));
  jnot g10998(.din(n11065), .dout(n11066));
  jand g10999(.dina(n11066), .dinb(n11064), .dout(n11067));
  jnot g11000(.din(n11067), .dout(n11068));
  jor  g11001(.dina(n10067), .dinb(n10059), .dout(n11069));
  jand g11002(.dina(n10068), .dinb(n10044), .dout(n11070));
  jnot g11003(.din(n11070), .dout(n11071));
  jand g11004(.dina(n11071), .dinb(n11069), .dout(n11072));
  jnot g11005(.din(n11072), .dout(n11073));
  jnot g11006(.din(n10047), .dout(n11074));
  jand g11007(.dina(n11074), .dinb(n10045), .dout(n11075));
  jnot g11008(.din(n11075), .dout(n11076));
  jor  g11009(.dina(n10057), .dinb(n10049), .dout(n11077));
  jand g11010(.dina(n11077), .dinb(n11076), .dout(n11078));
  jnot g11011(.din(n11078), .dout(n11079));
  jand g11012(.dina(n7315), .dinb(n2936), .dout(n11080));
  jand g11013(.dina(n7019), .dinb(n2940), .dout(n11081));
  jand g11014(.dina(n7313), .dinb(n2943), .dout(n11082));
  jor  g11015(.dina(n11082), .dinb(n11081), .dout(n11083));
  jor  g11016(.dina(n11083), .dinb(n11080), .dout(n11084));
  jor  g11017(.dina(n10046), .dinb(n93), .dout(n11085));
  jxor g11018(.dina(n11085), .dinb(n11084), .dout(n11086));
  jand g11019(.dina(n8270), .dinb(n71), .dout(n11087));
  jand g11020(.dina(n8022), .dinb(n731), .dout(n11088));
  jand g11021(.dina(n8268), .dinb(n796), .dout(n11089));
  jor  g11022(.dina(n11089), .dinb(n11088), .dout(n11090));
  jand g11023(.dina(n7692), .dinb(n1806), .dout(n11091));
  jor  g11024(.dina(n11091), .dinb(n11090), .dout(n11092));
  jor  g11025(.dina(n11092), .dinb(n11087), .dout(n11093));
  jxor g11026(.dina(n11093), .dinb(n77), .dout(n11094));
  jxor g11027(.dina(n11094), .dinb(n11086), .dout(n11095));
  jxor g11028(.dina(n11095), .dinb(n11079), .dout(n11096));
  jnot g11029(.din(n11096), .dout(n11097));
  jand g11030(.dina(n8938), .dinb(n806), .dout(n11098));
  jand g11031(.dina(n8723), .dinb(n1612), .dout(n11099));
  jand g11032(.dina(n8936), .dinb(n1620), .dout(n11100));
  jor  g11033(.dina(n11100), .dinb(n11099), .dout(n11101));
  jand g11034(.dina(n8740), .dinb(n1644), .dout(n11102));
  jor  g11035(.dina(n11102), .dinb(n11101), .dout(n11103));
  jor  g11036(.dina(n11103), .dinb(n11098), .dout(n11104));
  jxor g11037(.dina(n11104), .dinb(n65), .dout(n11105));
  jxor g11038(.dina(n11105), .dinb(n11097), .dout(n11106));
  jxor g11039(.dina(n11106), .dinb(n11073), .dout(n11107));
  jnot g11040(.din(n11107), .dout(n11108));
  jand g11041(.dina(n9886), .dinb(n1819), .dout(n11109));
  jand g11042(.dina(n9655), .dinb(n2243), .dout(n11110));
  jand g11043(.dina(n9656), .dinb(n2180), .dout(n11111));
  jand g11044(.dina(n9250), .dinb(n2185), .dout(n11112));
  jor  g11045(.dina(n11112), .dinb(n11111), .dout(n11113));
  jor  g11046(.dina(n11113), .dinb(n11110), .dout(n11114));
  jor  g11047(.dina(n11114), .dinb(n11109), .dout(n11115));
  jxor g11048(.dina(n11115), .dinb(n2196), .dout(n11116));
  jxor g11049(.dina(n11116), .dinb(n11108), .dout(n11117));
  jxor g11050(.dina(n11117), .dinb(n11068), .dout(n11118));
  jnot g11051(.din(n11118), .dout(n11119));
  jand g11052(.dina(n10862), .dinb(n2743), .dout(n11120));
  jand g11053(.dina(n10647), .dinb(n2752), .dout(n11121));
  jand g11054(.dina(n10305), .dinb(n2748), .dout(n11122));
  jand g11055(.dina(n9872), .dinb(n2757), .dout(n11123));
  jor  g11056(.dina(n11123), .dinb(n11122), .dout(n11124));
  jor  g11057(.dina(n11124), .dinb(n11121), .dout(n11125));
  jor  g11058(.dina(n11125), .dinb(n11120), .dout(n11126));
  jxor g11059(.dina(n11126), .dinb(n2441), .dout(n11127));
  jxor g11060(.dina(n11127), .dinb(n11119), .dout(n11128));
  jxor g11061(.dina(n11128), .dinb(n11063), .dout(n11129));
  jnot g11062(.din(n11129), .dout(n11130));
  jand g11063(.dina(n10836), .dinb(n10640), .dout(n11131));
  jand g11064(.dina(n10837), .dinb(n10658), .dout(n11132));
  jor  g11065(.dina(n11132), .dinb(n11131), .dout(n11133));
  jand g11066(.dina(n10834), .dinb(n10668), .dout(n11134));
  jand g11067(.dina(n10835), .dinb(n10663), .dout(n11135));
  jor  g11068(.dina(n11135), .dinb(n11134), .dout(n11136));
  jand g11069(.dina(n10832), .dinb(n10824), .dout(n11137));
  jand g11070(.dina(n10833), .dinb(n10819), .dout(n11138));
  jor  g11071(.dina(n11138), .dinb(n11137), .dout(n11139));
  jand g11072(.dina(n10817), .dinb(n10809), .dout(n11140));
  jand g11073(.dina(n10818), .dinb(n10671), .dout(n11141));
  jor  g11074(.dina(n11141), .dinb(n11140), .dout(n11142));
  jnot g11075(.din(n11142), .dout(n11143));
  jor  g11076(.dina(n8260), .dinb(n3424), .dout(n11144));
  jor  g11077(.dina(n7680), .dinb(n3211), .dout(n11145));
  jor  g11078(.dina(n7999), .dinb(n3429), .dout(n11146));
  jand g11079(.dina(n11146), .dinb(n11145), .dout(n11147));
  jand g11080(.dina(n11147), .dinb(n11144), .dout(n11148));
  jxor g11081(.dina(n11148), .dinb(\a[14] ), .dout(n11149));
  jxor g11082(.dina(n11149), .dinb(n11143), .dout(n11150));
  jand g11083(.dina(n10807), .dinb(n10799), .dout(n11151));
  jand g11084(.dina(n10808), .dinb(n10674), .dout(n11152));
  jor  g11085(.dina(n11152), .dinb(n11151), .dout(n11153));
  jor  g11086(.dina(n10797), .dinb(n10789), .dout(n11154));
  jand g11087(.dina(n10798), .dinb(n10677), .dout(n11155));
  jnot g11088(.din(n11155), .dout(n11156));
  jand g11089(.dina(n11156), .dinb(n11154), .dout(n11157));
  jnot g11090(.din(n11157), .dout(n11158));
  jor  g11091(.dina(n10786), .dinb(n10778), .dout(n11159));
  jand g11092(.dina(n10787), .dinb(n10682), .dout(n11160));
  jnot g11093(.din(n11160), .dout(n11161));
  jand g11094(.dina(n11161), .dinb(n11159), .dout(n11162));
  jnot g11095(.din(n11162), .dout(n11163));
  jand g11096(.dina(n10767), .dinb(n10687), .dout(n11164));
  jand g11097(.dina(n10776), .dinb(n10768), .dout(n11165));
  jor  g11098(.dina(n11165), .dinb(n11164), .dout(n11166));
  jor  g11099(.dina(n10765), .dinb(n10757), .dout(n11167));
  jand g11100(.dina(n10766), .dinb(n10688), .dout(n11168));
  jnot g11101(.din(n11168), .dout(n11169));
  jand g11102(.dina(n11169), .dinb(n11167), .dout(n11170));
  jnot g11103(.din(n11170), .dout(n11171));
  jor  g11104(.dina(n7061), .dinb(n4051), .dout(n11172));
  jand g11105(.dina(n6050), .dinb(n3729), .dout(n11173));
  jand g11106(.dina(n5084), .dinb(n3873), .dout(n11174));
  jor  g11107(.dina(n11174), .dinb(n11173), .dout(n11175));
  jand g11108(.dina(n5082), .dinb(n3933), .dout(n11176));
  jor  g11109(.dina(n11176), .dinb(n11175), .dout(n11177));
  jnot g11110(.din(n11177), .dout(n11178));
  jand g11111(.dina(n11178), .dinb(n11172), .dout(n11179));
  jnot g11112(.din(n11179), .dout(n11180));
  jand g11113(.dina(n1577), .dinb(n1037), .dout(n11181));
  jand g11114(.dina(n11181), .dinb(n454), .dout(n11182));
  jand g11115(.dina(n11182), .dinb(n352), .dout(n11183));
  jand g11116(.dina(n630), .dinb(n1346), .dout(n11184));
  jand g11117(.dina(n11184), .dinb(n4590), .dout(n11185));
  jand g11118(.dina(n11185), .dinb(n7769), .dout(n11186));
  jand g11119(.dina(n11186), .dinb(n11183), .dout(n11187));
  jand g11120(.dina(n1756), .dinb(n1429), .dout(n11188));
  jand g11121(.dina(n11188), .dinb(n811), .dout(n11189));
  jand g11122(.dina(n11189), .dinb(n676), .dout(n11190));
  jand g11123(.dina(n11190), .dinb(n662), .dout(n11191));
  jand g11124(.dina(n11191), .dinb(n11187), .dout(n11192));
  jand g11125(.dina(n2025), .dinb(n647), .dout(n11193));
  jand g11126(.dina(n11193), .dinb(n1088), .dout(n11194));
  jand g11127(.dina(n10393), .dinb(n82), .dout(n11195));
  jand g11128(.dina(n11195), .dinb(n11194), .dout(n11196));
  jand g11129(.dina(n11196), .dinb(n11192), .dout(n11197));
  jand g11130(.dina(n8361), .dinb(n1380), .dout(n11198));
  jand g11131(.dina(n5282), .dinb(n1326), .dout(n11199));
  jand g11132(.dina(n11199), .dinb(n11198), .dout(n11200));
  jand g11133(.dina(n8815), .dinb(n827), .dout(n11201));
  jand g11134(.dina(n11201), .dinb(n11200), .dout(n11202));
  jand g11135(.dina(n1190), .dinb(n638), .dout(n11203));
  jand g11136(.dina(n11203), .dinb(n1511), .dout(n11204));
  jand g11137(.dina(n11204), .dinb(n1098), .dout(n11205));
  jand g11138(.dina(n1461), .dinb(n1043), .dout(n11206));
  jand g11139(.dina(n11206), .dinb(n1544), .dout(n11207));
  jand g11140(.dina(n11207), .dinb(n11205), .dout(n11208));
  jand g11141(.dina(n495), .dinb(n1360), .dout(n11209));
  jand g11142(.dina(n11209), .dinb(n472), .dout(n11210));
  jand g11143(.dina(n2491), .dinb(n674), .dout(n11211));
  jand g11144(.dina(n11211), .dinb(n11210), .dout(n11212));
  jand g11145(.dina(n11212), .dinb(n5355), .dout(n11213));
  jand g11146(.dina(n11213), .dinb(n11208), .dout(n11214));
  jand g11147(.dina(n11214), .dinb(n11202), .dout(n11215));
  jand g11148(.dina(n11215), .dinb(n1559), .dout(n11216));
  jand g11149(.dina(n11216), .dinb(n11197), .dout(n11217));
  jand g11150(.dina(n5248), .dinb(n704), .dout(n11218));
  jand g11151(.dina(n11218), .dinb(n1965), .dout(n11219));
  jand g11152(.dina(n1470), .dinb(n470), .dout(n11220));
  jand g11153(.dina(n11220), .dinb(n4511), .dout(n11221));
  jand g11154(.dina(n11221), .dinb(n9132), .dout(n11222));
  jand g11155(.dina(n11222), .dinb(n11219), .dout(n11223));
  jand g11156(.dina(n1537), .dinb(n1228), .dout(n11224));
  jand g11157(.dina(n11224), .dinb(n699), .dout(n11225));
  jand g11158(.dina(n1345), .dinb(n1738), .dout(n11226));
  jand g11159(.dina(n11226), .dinb(n11225), .dout(n11227));
  jand g11160(.dina(n1591), .dinb(n1261), .dout(n11228));
  jand g11161(.dina(n1159), .dinb(n1237), .dout(n11229));
  jand g11162(.dina(n11229), .dinb(n931), .dout(n11230));
  jand g11163(.dina(n11230), .dinb(n11228), .dout(n11231));
  jand g11164(.dina(n11231), .dinb(n523), .dout(n11232));
  jand g11165(.dina(n11232), .dinb(n11227), .dout(n11233));
  jand g11166(.dina(n2612), .dinb(n547), .dout(n11234));
  jand g11167(.dina(n2119), .dinb(n456), .dout(n11235));
  jand g11168(.dina(n11235), .dinb(n664), .dout(n11236));
  jand g11169(.dina(n11236), .dinb(n5504), .dout(n11237));
  jand g11170(.dina(n11237), .dinb(n11234), .dout(n11238));
  jand g11171(.dina(n11238), .dinb(n4449), .dout(n11239));
  jand g11172(.dina(n11239), .dinb(n11233), .dout(n11240));
  jand g11173(.dina(n695), .dinb(n121), .dout(n11241));
  jand g11174(.dina(n11241), .dinb(n650), .dout(n11242));
  jand g11175(.dina(n11242), .dinb(n654), .dout(n11243));
  jand g11176(.dina(n11243), .dinb(n11240), .dout(n11244));
  jand g11177(.dina(n11244), .dinb(n11223), .dout(n11245));
  jand g11178(.dina(n11245), .dinb(n11217), .dout(n11246));
  jnot g11179(.din(n11246), .dout(n11247));
  jxor g11180(.dina(n11247), .dinb(n10754), .dout(n11248));
  jxor g11181(.dina(n11248), .dinb(n11180), .dout(n11249));
  jxor g11182(.dina(n11249), .dinb(n11171), .dout(n11250));
  jnot g11183(.din(n11250), .dout(n11251));
  jor  g11184(.dina(n4473), .dinb(n4343), .dout(n11252));
  jor  g11185(.dina(n4019), .dinb(n4346), .dout(n11253));
  jor  g11186(.dina(n3929), .dinb(n3683), .dout(n11254));
  jand g11187(.dina(n11254), .dinb(n11253), .dout(n11255));
  jor  g11188(.dina(n4471), .dinb(n4348), .dout(n11256));
  jand g11189(.dina(n11256), .dinb(n11255), .dout(n11257));
  jand g11190(.dina(n11257), .dinb(n11252), .dout(n11258));
  jxor g11191(.dina(n11258), .dinb(\a[29] ), .dout(n11259));
  jxor g11192(.dina(n11259), .dinb(n11251), .dout(n11260));
  jxor g11193(.dina(n11260), .dinb(n11166), .dout(n11261));
  jnot g11194(.din(n11261), .dout(n11262));
  jor  g11195(.dina(n4688), .dinb(n2303), .dout(n11263));
  jor  g11196(.dina(n4526), .dinb(n2306), .dout(n11264));
  jor  g11197(.dina(n4686), .dinb(n2309), .dout(n11265));
  jand g11198(.dina(n11265), .dinb(n11264), .dout(n11266));
  jor  g11199(.dina(n4596), .dinb(n1805), .dout(n11267));
  jand g11200(.dina(n11267), .dinb(n11266), .dout(n11268));
  jand g11201(.dina(n11268), .dinb(n11263), .dout(n11269));
  jxor g11202(.dina(n11269), .dinb(\a[26] ), .dout(n11270));
  jxor g11203(.dina(n11270), .dinb(n11262), .dout(n11271));
  jxor g11204(.dina(n11271), .dinb(n11163), .dout(n11272));
  jnot g11205(.din(n11272), .dout(n11273));
  jor  g11206(.dina(n5549), .dinb(n807), .dout(n11274));
  jor  g11207(.dina(n5422), .dinb(n1613), .dout(n11275));
  jor  g11208(.dina(n5264), .dinb(n1617), .dout(n11276));
  jand g11209(.dina(n11276), .dinb(n11275), .dout(n11277));
  jor  g11210(.dina(n5364), .dinb(n1621), .dout(n11278));
  jand g11211(.dina(n11278), .dinb(n11277), .dout(n11279));
  jand g11212(.dina(n11279), .dinb(n11274), .dout(n11280));
  jxor g11213(.dina(n11280), .dinb(\a[23] ), .dout(n11281));
  jxor g11214(.dina(n11281), .dinb(n11273), .dout(n11282));
  jxor g11215(.dina(n11282), .dinb(n11158), .dout(n11283));
  jor  g11216(.dina(n6516), .dinb(n1820), .dout(n11284));
  jor  g11217(.dina(n6205), .dinb(n2181), .dout(n11285));
  jor  g11218(.dina(n5525), .dinb(n2186), .dout(n11286));
  jor  g11219(.dina(n6390), .dinb(n2189), .dout(n11287));
  jand g11220(.dina(n11287), .dinb(n11286), .dout(n11288));
  jand g11221(.dina(n11288), .dinb(n11285), .dout(n11289));
  jand g11222(.dina(n11289), .dinb(n11284), .dout(n11290));
  jxor g11223(.dina(n11290), .dinb(n2196), .dout(n11291));
  jxor g11224(.dina(n11291), .dinb(n11283), .dout(n11292));
  jxor g11225(.dina(n11292), .dinb(n11153), .dout(n11293));
  jnot g11226(.din(n11293), .dout(n11294));
  jor  g11227(.dina(n7301), .dinb(n2753), .dout(n11295));
  jor  g11228(.dina(n7303), .dinb(n2744), .dout(n11296));
  jor  g11229(.dina(n6297), .dinb(n2758), .dout(n11297));
  jor  g11230(.dina(n6489), .dinb(n2749), .dout(n11298));
  jand g11231(.dina(n11298), .dinb(n11297), .dout(n11299));
  jand g11232(.dina(n11299), .dinb(n11296), .dout(n11300));
  jand g11233(.dina(n11300), .dinb(n11295), .dout(n11301));
  jxor g11234(.dina(n11301), .dinb(\a[17] ), .dout(n11302));
  jxor g11235(.dina(n11302), .dinb(n11294), .dout(n11303));
  jxor g11236(.dina(n11303), .dinb(n11150), .dout(n11304));
  jxor g11237(.dina(n11304), .dinb(n11139), .dout(n11305));
  jxor g11238(.dina(n11305), .dinb(n11136), .dout(n11306));
  jxor g11239(.dina(n11306), .dinb(n10836), .dout(n11307));
  jxor g11240(.dina(n11307), .dinb(n11133), .dout(n11308));
  jand g11241(.dina(n11308), .dinb(n3423), .dout(n11309));
  jand g11242(.dina(n11306), .dinb(n3569), .dout(n11310));
  jand g11243(.dina(n10836), .dinb(n3428), .dout(n11311));
  jand g11244(.dina(n10640), .dinb(n3210), .dout(n11312));
  jor  g11245(.dina(n11312), .dinb(n11311), .dout(n11313));
  jor  g11246(.dina(n11313), .dinb(n11310), .dout(n11314));
  jor  g11247(.dina(n11314), .dinb(n11309), .dout(n11315));
  jxor g11248(.dina(n11315), .dinb(n3473), .dout(n11316));
  jxor g11249(.dina(n11316), .dinb(n11130), .dout(n11317));
  jnot g11250(.din(n11317), .dout(n11318));
  jxor g11251(.dina(n11318), .dinb(n11058), .dout(n11319));
  jnot g11252(.din(n11319), .dout(n11320));
  jand g11253(.dina(n11292), .dinb(n11153), .dout(n11321));
  jnot g11254(.din(n11321), .dout(n11322));
  jor  g11255(.dina(n11302), .dinb(n11294), .dout(n11323));
  jand g11256(.dina(n11323), .dinb(n11322), .dout(n11324));
  jor  g11257(.dina(n7999), .dinb(n3211), .dout(n11325));
  jor  g11258(.dina(n8295), .dinb(n3424), .dout(n11326));
  jand g11259(.dina(n11326), .dinb(n11325), .dout(n11327));
  jxor g11260(.dina(n11327), .dinb(\a[14] ), .dout(n11328));
  jor  g11261(.dina(n11328), .dinb(n11324), .dout(n11329));
  jxor g11262(.dina(n11328), .dinb(n11324), .dout(n11330));
  jand g11263(.dina(n11282), .dinb(n11158), .dout(n11331));
  jand g11264(.dina(n11291), .dinb(n11283), .dout(n11332));
  jor  g11265(.dina(n11332), .dinb(n11331), .dout(n11333));
  jand g11266(.dina(n11271), .dinb(n11163), .dout(n11334));
  jnot g11267(.din(n11334), .dout(n11335));
  jor  g11268(.dina(n11281), .dinb(n11273), .dout(n11336));
  jand g11269(.dina(n11336), .dinb(n11335), .dout(n11337));
  jnot g11270(.din(n11337), .dout(n11338));
  jand g11271(.dina(n11260), .dinb(n11166), .dout(n11339));
  jnot g11272(.din(n11339), .dout(n11340));
  jor  g11273(.dina(n11270), .dinb(n11262), .dout(n11341));
  jand g11274(.dina(n11341), .dinb(n11340), .dout(n11342));
  jnot g11275(.din(n11342), .dout(n11343));
  jnot g11276(.din(n10754), .dout(n11344));
  jand g11277(.dina(n11246), .dinb(n11344), .dout(n11345));
  jand g11278(.dina(n11248), .dinb(n11180), .dout(n11346));
  jor  g11279(.dina(n11346), .dinb(n11345), .dout(n11347));
  jor  g11280(.dina(n7061), .dinb(n4038), .dout(n11348));
  jand g11281(.dina(n5082), .dinb(n3873), .dout(n11349));
  jand g11282(.dina(n5084), .dinb(n3930), .dout(n11350));
  jor  g11283(.dina(n11350), .dinb(n11349), .dout(n11351));
  jand g11284(.dina(n6050), .dinb(n3933), .dout(n11352));
  jor  g11285(.dina(n11352), .dinb(n11351), .dout(n11353));
  jnot g11286(.din(n11353), .dout(n11354));
  jand g11287(.dina(n11354), .dinb(n11348), .dout(n11355));
  jnot g11288(.din(n11355), .dout(n11356));
  jand g11289(.dina(n1227), .dinb(n1225), .dout(n11357));
  jand g11290(.dina(n11357), .dinb(n869), .dout(n11358));
  jand g11291(.dina(n11358), .dinb(n6421), .dout(n11359));
  jand g11292(.dina(n1861), .dinb(n351), .dout(n11360));
  jand g11293(.dina(n950), .dinb(n621), .dout(n11361));
  jand g11294(.dina(n11361), .dinb(n11360), .dout(n11362));
  jand g11295(.dina(n11362), .dinb(n11359), .dout(n11363));
  jand g11296(.dina(n3328), .dinb(n1351), .dout(n11364));
  jand g11297(.dina(n11364), .dinb(n2096), .dout(n11365));
  jand g11298(.dina(n11365), .dinb(n1917), .dout(n11366));
  jand g11299(.dina(n8107), .dinb(n463), .dout(n11367));
  jand g11300(.dina(n11367), .dinb(n11366), .dout(n11368));
  jand g11301(.dina(n11368), .dinb(n11363), .dout(n11369));
  jand g11302(.dina(n9774), .dinb(n445), .dout(n11370));
  jand g11303(.dina(n11370), .dinb(n1506), .dout(n11371));
  jand g11304(.dina(n1207), .dinb(n662), .dout(n11372));
  jand g11305(.dina(n2620), .dinb(n496), .dout(n11373));
  jand g11306(.dina(n2131), .dinb(n639), .dout(n11374));
  jand g11307(.dina(n11374), .dinb(n11373), .dout(n11375));
  jand g11308(.dina(n8580), .dinb(n1515), .dout(n11376));
  jand g11309(.dina(n11376), .dinb(n537), .dout(n11377));
  jand g11310(.dina(n11377), .dinb(n11375), .dout(n11378));
  jand g11311(.dina(n11378), .dinb(n11372), .dout(n11379));
  jand g11312(.dina(n11379), .dinb(n11371), .dout(n11380));
  jand g11313(.dina(n11380), .dinb(n11369), .dout(n11381));
  jand g11314(.dina(n8120), .dinb(n1205), .dout(n11382));
  jand g11315(.dina(n11382), .dinb(n843), .dout(n11383));
  jand g11316(.dina(n1346), .dinb(n1040), .dout(n11384));
  jand g11317(.dina(n11384), .dinb(n918), .dout(n11385));
  jand g11318(.dina(n11385), .dinb(n11383), .dout(n11386));
  jand g11319(.dina(n11386), .dinb(n2152), .dout(n11387));
  jand g11320(.dina(n11387), .dinb(n2586), .dout(n11388));
  jand g11321(.dina(n11388), .dinb(n11381), .dout(n11389));
  jand g11322(.dina(n8601), .dinb(n2042), .dout(n11390));
  jand g11323(.dina(n1016), .dinb(n517), .dout(n11391));
  jand g11324(.dina(n11391), .dinb(n697), .dout(n11392));
  jand g11325(.dina(n11392), .dinb(n11390), .dout(n11393));
  jand g11326(.dina(n1721), .dinb(n1429), .dout(n11394));
  jand g11327(.dina(n11394), .dinb(n1832), .dout(n11395));
  jand g11328(.dina(n11395), .dinb(n11393), .dout(n11396));
  jand g11329(.dina(n1527), .dinb(n982), .dout(n11397));
  jand g11330(.dina(n11397), .dinb(n1511), .dout(n11398));
  jand g11331(.dina(n11398), .dinb(n2571), .dout(n11399));
  jand g11332(.dina(n11399), .dinb(n11396), .dout(n11400));
  jand g11333(.dina(n8583), .dinb(n5456), .dout(n11401));
  jand g11334(.dina(n4417), .dinb(n2483), .dout(n11402));
  jand g11335(.dina(n11402), .dinb(n11401), .dout(n11403));
  jand g11336(.dina(n11403), .dinb(n8820), .dout(n11404));
  jand g11337(.dina(n11404), .dinb(n5406), .dout(n11405));
  jand g11338(.dina(n11405), .dinb(n11400), .dout(n11406));
  jnot g11339(.din(n1083), .dout(n11407));
  jand g11340(.dina(n11407), .dinb(n848), .dout(n11408));
  jand g11341(.dina(n11408), .dinb(n6478), .dout(n11409));
  jand g11342(.dina(n3176), .dinb(n1304), .dout(n11410));
  jand g11343(.dina(n11410), .dinb(n3978), .dout(n11411));
  jand g11344(.dina(n11411), .dinb(n11409), .dout(n11412));
  jand g11345(.dina(n320), .dinb(n108), .dout(n11413));
  jand g11346(.dina(n1237), .dinb(n1053), .dout(n11414));
  jand g11347(.dina(n11414), .dinb(n470), .dout(n11415));
  jand g11348(.dina(n11415), .dinb(n11413), .dout(n11416));
  jand g11349(.dina(n11416), .dinb(n598), .dout(n11417));
  jand g11350(.dina(n11417), .dinb(n11412), .dout(n11418));
  jand g11351(.dina(n8362), .dinb(n1701), .dout(n11419));
  jand g11352(.dina(n11419), .dinb(n2499), .dout(n11420));
  jand g11353(.dina(n11420), .dinb(n2528), .dout(n11421));
  jand g11354(.dina(n1107), .dinb(n1036), .dout(n11422));
  jand g11355(.dina(n11422), .dinb(n452), .dout(n11423));
  jand g11356(.dina(n499), .dinb(n442), .dout(n11424));
  jand g11357(.dina(n11424), .dinb(n920), .dout(n11425));
  jand g11358(.dina(n11425), .dinb(n11423), .dout(n11426));
  jand g11359(.dina(n11426), .dinb(n1477), .dout(n11427));
  jand g11360(.dina(n11427), .dinb(n11421), .dout(n11428));
  jand g11361(.dina(n11428), .dinb(n11418), .dout(n11429));
  jand g11362(.dina(n11429), .dinb(n11406), .dout(n11430));
  jand g11363(.dina(n11430), .dinb(n11389), .dout(n11431));
  jxor g11364(.dina(n11431), .dinb(n11247), .dout(n11432));
  jxor g11365(.dina(n11432), .dinb(n11356), .dout(n11433));
  jxor g11366(.dina(n11433), .dinb(n11347), .dout(n11434));
  jnot g11367(.din(n11434), .dout(n11435));
  jand g11368(.dina(n11249), .dinb(n11171), .dout(n11436));
  jnot g11369(.din(n11436), .dout(n11437));
  jor  g11370(.dina(n11259), .dinb(n11251), .dout(n11438));
  jand g11371(.dina(n11438), .dinb(n11437), .dout(n11439));
  jxor g11372(.dina(n11439), .dinb(n11435), .dout(n11440));
  jor  g11373(.dina(n4726), .dinb(n4343), .dout(n11441));
  jor  g11374(.dina(n4471), .dinb(n4346), .dout(n11442));
  jor  g11375(.dina(n4019), .dinb(n3683), .dout(n11443));
  jor  g11376(.dina(n4596), .dinb(n4348), .dout(n11444));
  jand g11377(.dina(n11444), .dinb(n11443), .dout(n11445));
  jand g11378(.dina(n11445), .dinb(n11442), .dout(n11446));
  jand g11379(.dina(n11446), .dinb(n11441), .dout(n11447));
  jxor g11380(.dina(n11447), .dinb(n93), .dout(n11448));
  jxor g11381(.dina(n11448), .dinb(n11440), .dout(n11449));
  jnot g11382(.din(n11449), .dout(n11450));
  jor  g11383(.dina(n5266), .dinb(n2303), .dout(n11451));
  jor  g11384(.dina(n4686), .dinb(n2306), .dout(n11452));
  jor  g11385(.dina(n4526), .dinb(n1805), .dout(n11453));
  jand g11386(.dina(n11453), .dinb(n11452), .dout(n11454));
  jor  g11387(.dina(n5264), .dinb(n2309), .dout(n11455));
  jand g11388(.dina(n11455), .dinb(n11454), .dout(n11456));
  jand g11389(.dina(n11456), .dinb(n11451), .dout(n11457));
  jxor g11390(.dina(n11457), .dinb(\a[26] ), .dout(n11458));
  jxor g11391(.dina(n11458), .dinb(n11450), .dout(n11459));
  jxor g11392(.dina(n11459), .dinb(n11343), .dout(n11460));
  jor  g11393(.dina(n5527), .dinb(n807), .dout(n11461));
  jor  g11394(.dina(n5364), .dinb(n1613), .dout(n11462));
  jor  g11395(.dina(n5525), .dinb(n1621), .dout(n11463));
  jor  g11396(.dina(n5422), .dinb(n1617), .dout(n11464));
  jand g11397(.dina(n11464), .dinb(n11463), .dout(n11465));
  jand g11398(.dina(n11465), .dinb(n11462), .dout(n11466));
  jand g11399(.dina(n11466), .dinb(n11461), .dout(n11467));
  jxor g11400(.dina(n11467), .dinb(n65), .dout(n11468));
  jxor g11401(.dina(n11468), .dinb(n11460), .dout(n11469));
  jxor g11402(.dina(n11469), .dinb(n11338), .dout(n11470));
  jnot g11403(.din(n11470), .dout(n11471));
  jor  g11404(.dina(n6999), .dinb(n1820), .dout(n11472));
  jor  g11405(.dina(n6390), .dinb(n2181), .dout(n11473));
  jor  g11406(.dina(n6297), .dinb(n2189), .dout(n11474));
  jand g11407(.dina(n11474), .dinb(n11473), .dout(n11475));
  jor  g11408(.dina(n6205), .dinb(n2186), .dout(n11476));
  jand g11409(.dina(n11476), .dinb(n11475), .dout(n11477));
  jand g11410(.dina(n11477), .dinb(n11472), .dout(n11478));
  jxor g11411(.dina(n11478), .dinb(\a[20] ), .dout(n11479));
  jxor g11412(.dina(n11479), .dinb(n11471), .dout(n11480));
  jxor g11413(.dina(n11480), .dinb(n11333), .dout(n11481));
  jor  g11414(.dina(n7682), .dinb(n2744), .dout(n11482));
  jor  g11415(.dina(n7301), .dinb(n2749), .dout(n11483));
  jor  g11416(.dina(n6489), .dinb(n2758), .dout(n11484));
  jor  g11417(.dina(n7680), .dinb(n2753), .dout(n11485));
  jand g11418(.dina(n11485), .dinb(n11484), .dout(n11486));
  jand g11419(.dina(n11486), .dinb(n11483), .dout(n11487));
  jand g11420(.dina(n11487), .dinb(n11482), .dout(n11488));
  jxor g11421(.dina(n11488), .dinb(n2441), .dout(n11489));
  jxor g11422(.dina(n11489), .dinb(n11481), .dout(n11490));
  jand g11423(.dina(n11490), .dinb(n11330), .dout(n11491));
  jnot g11424(.din(n11491), .dout(n11492));
  jand g11425(.dina(n11492), .dinb(n11329), .dout(n11493));
  jnot g11426(.din(n11493), .dout(n11494));
  jand g11427(.dina(n11480), .dinb(n11333), .dout(n11495));
  jand g11428(.dina(n11489), .dinb(n11481), .dout(n11496));
  jor  g11429(.dina(n11496), .dinb(n11495), .dout(n11497));
  jor  g11430(.dina(n8002), .dinb(n2744), .dout(n11498));
  jor  g11431(.dina(n7301), .dinb(n2758), .dout(n11499));
  jor  g11432(.dina(n7999), .dinb(n2753), .dout(n11500));
  jor  g11433(.dina(n7680), .dinb(n2749), .dout(n11501));
  jand g11434(.dina(n11501), .dinb(n11500), .dout(n11502));
  jand g11435(.dina(n11502), .dinb(n11499), .dout(n11503));
  jand g11436(.dina(n11503), .dinb(n11498), .dout(n11504));
  jxor g11437(.dina(n11504), .dinb(n2441), .dout(n11505));
  jxor g11438(.dina(n11505), .dinb(n11497), .dout(n11506));
  jand g11439(.dina(n11469), .dinb(n11338), .dout(n11507));
  jnot g11440(.din(n11507), .dout(n11508));
  jor  g11441(.dina(n11479), .dinb(n11471), .dout(n11509));
  jand g11442(.dina(n11509), .dinb(n11508), .dout(n11510));
  jnot g11443(.din(n11510), .dout(n11511));
  jand g11444(.dina(n11459), .dinb(n11343), .dout(n11512));
  jand g11445(.dina(n11468), .dinb(n11460), .dout(n11513));
  jor  g11446(.dina(n11513), .dinb(n11512), .dout(n11514));
  jand g11447(.dina(n11448), .dinb(n11440), .dout(n11515));
  jnot g11448(.din(n11515), .dout(n11516));
  jor  g11449(.dina(n11458), .dinb(n11450), .dout(n11517));
  jand g11450(.dina(n11517), .dinb(n11516), .dout(n11518));
  jnot g11451(.din(n11518), .dout(n11519));
  jand g11452(.dina(n11433), .dinb(n11347), .dout(n11520));
  jnot g11453(.din(n11520), .dout(n11521));
  jor  g11454(.dina(n11439), .dinb(n11435), .dout(n11522));
  jand g11455(.dina(n11522), .dinb(n11521), .dout(n11523));
  jnot g11456(.din(n11523), .dout(n11524));
  jor  g11457(.dina(n7061), .dinb(n4021), .dout(n11525));
  jand g11458(.dina(n6050), .dinb(n3873), .dout(n11526));
  jand g11459(.dina(n5084), .dinb(n4406), .dout(n11527));
  jor  g11460(.dina(n11527), .dinb(n11526), .dout(n11528));
  jand g11461(.dina(n5082), .dinb(n3930), .dout(n11529));
  jor  g11462(.dina(n11529), .dinb(n11528), .dout(n11530));
  jnot g11463(.din(n11530), .dout(n11531));
  jand g11464(.dina(n11531), .dinb(n11525), .dout(n11532));
  jnot g11465(.din(n11532), .dout(n11533));
  jand g11466(.dina(n3885), .dinb(n933), .dout(n11534));
  jand g11467(.dina(n908), .dinb(n328), .dout(n11535));
  jand g11468(.dina(n11535), .dinb(n8370), .dout(n11536));
  jand g11469(.dina(n11536), .dinb(n11534), .dout(n11537));
  jand g11470(.dina(n1005), .dinb(n517), .dout(n11538));
  jand g11471(.dina(n11538), .dinb(n1995), .dout(n11539));
  jand g11472(.dina(n534), .dinb(n411), .dout(n11540));
  jand g11473(.dina(n11540), .dinb(n11539), .dout(n11541));
  jand g11474(.dina(n11541), .dinb(n3026), .dout(n11542));
  jand g11475(.dina(n11542), .dinb(n11537), .dout(n11543));
  jand g11476(.dina(n11543), .dinb(n3812), .dout(n11544));
  jand g11477(.dina(n11544), .dinb(n8399), .dout(n11545));
  jand g11478(.dina(n547), .dinb(n1334), .dout(n11546));
  jand g11479(.dina(n11546), .dinb(n492), .dout(n11547));
  jand g11480(.dina(n11547), .dinb(n4429), .dout(n11548));
  jand g11481(.dina(n839), .dinb(n1203), .dout(n11549));
  jand g11482(.dina(n2595), .dinb(n558), .dout(n11550));
  jand g11483(.dina(n11550), .dinb(n11549), .dout(n11551));
  jand g11484(.dina(n11551), .dinb(n3014), .dout(n11552));
  jand g11485(.dina(n11552), .dinb(n11548), .dout(n11553));
  jand g11486(.dina(n6334), .dinb(n3827), .dout(n11554));
  jand g11487(.dina(n11554), .dinb(n9543), .dout(n11555));
  jand g11488(.dina(n11555), .dinb(n1524), .dout(n11556));
  jand g11489(.dina(n11556), .dinb(n11553), .dout(n11557));
  jand g11490(.dina(n11557), .dinb(n11545), .dout(n11558));
  jand g11491(.dina(n11558), .dinb(n9330), .dout(n11559));
  jand g11492(.dina(n11559), .dinb(n11246), .dout(n11560));
  jnot g11493(.din(n11560), .dout(n11561));
  jor  g11494(.dina(n11559), .dinb(n11246), .dout(n11562));
  jand g11495(.dina(n11562), .dinb(n3473), .dout(n11563));
  jand g11496(.dina(n11563), .dinb(n11561), .dout(n11564));
  jnot g11497(.din(n11564), .dout(n11565));
  jand g11498(.dina(n11565), .dinb(n3473), .dout(n11566));
  jand g11499(.dina(n11565), .dinb(n11562), .dout(n11567));
  jand g11500(.dina(n11567), .dinb(n11561), .dout(n11568));
  jor  g11501(.dina(n11568), .dinb(n11566), .dout(n11569));
  jnot g11502(.din(n11569), .dout(n11570));
  jor  g11503(.dina(n11431), .dinb(n11247), .dout(n11571));
  jand g11504(.dina(n11432), .dinb(n11356), .dout(n11572));
  jnot g11505(.din(n11572), .dout(n11573));
  jand g11506(.dina(n11573), .dinb(n11571), .dout(n11574));
  jxor g11507(.dina(n11574), .dinb(n11570), .dout(n11575));
  jxor g11508(.dina(n11575), .dinb(n11533), .dout(n11576));
  jnot g11509(.din(n11576), .dout(n11577));
  jor  g11510(.dina(n4714), .dinb(n4343), .dout(n11578));
  jor  g11511(.dina(n4596), .dinb(n4346), .dout(n11579));
  jor  g11512(.dina(n4526), .dinb(n4348), .dout(n11580));
  jand g11513(.dina(n11580), .dinb(n11579), .dout(n11581));
  jor  g11514(.dina(n4471), .dinb(n3683), .dout(n11582));
  jand g11515(.dina(n11582), .dinb(n11581), .dout(n11583));
  jand g11516(.dina(n11583), .dinb(n11578), .dout(n11584));
  jxor g11517(.dina(n11584), .dinb(\a[29] ), .dout(n11585));
  jxor g11518(.dina(n11585), .dinb(n11577), .dout(n11586));
  jxor g11519(.dina(n11586), .dinb(n11524), .dout(n11587));
  jnot g11520(.din(n11587), .dout(n11588));
  jor  g11521(.dina(n5560), .dinb(n2303), .dout(n11589));
  jor  g11522(.dina(n5264), .dinb(n2306), .dout(n11590));
  jor  g11523(.dina(n5422), .dinb(n2309), .dout(n11591));
  jand g11524(.dina(n11591), .dinb(n11590), .dout(n11592));
  jor  g11525(.dina(n4686), .dinb(n1805), .dout(n11593));
  jand g11526(.dina(n11593), .dinb(n11592), .dout(n11594));
  jand g11527(.dina(n11594), .dinb(n11589), .dout(n11595));
  jxor g11528(.dina(n11595), .dinb(\a[26] ), .dout(n11596));
  jxor g11529(.dina(n11596), .dinb(n11588), .dout(n11597));
  jxor g11530(.dina(n11597), .dinb(n11519), .dout(n11598));
  jor  g11531(.dina(n6207), .dinb(n807), .dout(n11599));
  jor  g11532(.dina(n5525), .dinb(n1613), .dout(n11600));
  jor  g11533(.dina(n5364), .dinb(n1617), .dout(n11601));
  jor  g11534(.dina(n6205), .dinb(n1621), .dout(n11602));
  jand g11535(.dina(n11602), .dinb(n11601), .dout(n11603));
  jand g11536(.dina(n11603), .dinb(n11600), .dout(n11604));
  jand g11537(.dina(n11604), .dinb(n11599), .dout(n11605));
  jxor g11538(.dina(n11605), .dinb(n65), .dout(n11606));
  jxor g11539(.dina(n11606), .dinb(n11598), .dout(n11607));
  jxor g11540(.dina(n11607), .dinb(n11514), .dout(n11608));
  jor  g11541(.dina(n6491), .dinb(n1820), .dout(n11609));
  jor  g11542(.dina(n6297), .dinb(n2181), .dout(n11610));
  jor  g11543(.dina(n6390), .dinb(n2186), .dout(n11611));
  jor  g11544(.dina(n6489), .dinb(n2189), .dout(n11612));
  jand g11545(.dina(n11612), .dinb(n11611), .dout(n11613));
  jand g11546(.dina(n11613), .dinb(n11610), .dout(n11614));
  jand g11547(.dina(n11614), .dinb(n11609), .dout(n11615));
  jxor g11548(.dina(n11615), .dinb(n2196), .dout(n11616));
  jxor g11549(.dina(n11616), .dinb(n11608), .dout(n11617));
  jxor g11550(.dina(n11617), .dinb(n11511), .dout(n11618));
  jxor g11551(.dina(n11618), .dinb(n11506), .dout(n11619));
  jxor g11552(.dina(n11619), .dinb(n11494), .dout(n11620));
  jnot g11553(.din(n11620), .dout(n11621));
  jor  g11554(.dina(n11149), .dinb(n11143), .dout(n11622));
  jand g11555(.dina(n11303), .dinb(n11150), .dout(n11623));
  jnot g11556(.din(n11623), .dout(n11624));
  jand g11557(.dina(n11624), .dinb(n11622), .dout(n11625));
  jnot g11558(.din(n11625), .dout(n11626));
  jxor g11559(.dina(n11490), .dinb(n11330), .dout(n11627));
  jand g11560(.dina(n11627), .dinb(n11626), .dout(n11628));
  jnot g11561(.din(n11628), .dout(n11629));
  jxor g11562(.dina(n11627), .dinb(n11626), .dout(n11630));
  jnot g11563(.din(n11630), .dout(n11631));
  jand g11564(.dina(n11304), .dinb(n11139), .dout(n11632));
  jnot g11565(.din(n11632), .dout(n11633));
  jnot g11566(.din(n11134), .dout(n11634));
  jnot g11567(.din(n10659), .dout(n11635));
  jor  g11568(.dina(n10639), .dinb(n10625), .dout(n11636));
  jand g11569(.dina(n11636), .dinb(n11635), .dout(n11637));
  jnot g11570(.din(n10835), .dout(n11638));
  jor  g11571(.dina(n11638), .dinb(n11637), .dout(n11639));
  jand g11572(.dina(n11639), .dinb(n11634), .dout(n11640));
  jnot g11573(.din(n11305), .dout(n11641));
  jor  g11574(.dina(n11641), .dinb(n11640), .dout(n11642));
  jand g11575(.dina(n11642), .dinb(n11633), .dout(n11643));
  jor  g11576(.dina(n11643), .dinb(n11631), .dout(n11644));
  jand g11577(.dina(n11644), .dinb(n11629), .dout(n11645));
  jxor g11578(.dina(n11645), .dinb(n11621), .dout(n11646));
  jxor g11579(.dina(n11643), .dinb(n11631), .dout(n11647));
  jand g11580(.dina(n11647), .dinb(n11646), .dout(n11648));
  jand g11581(.dina(n11647), .dinb(n11306), .dout(n11649));
  jand g11582(.dina(n11306), .dinb(n10836), .dout(n11650));
  jand g11583(.dina(n11307), .dinb(n11133), .dout(n11651));
  jor  g11584(.dina(n11651), .dinb(n11650), .dout(n11652));
  jxor g11585(.dina(n11647), .dinb(n11306), .dout(n11653));
  jand g11586(.dina(n11653), .dinb(n11652), .dout(n11654));
  jor  g11587(.dina(n11654), .dinb(n11649), .dout(n11655));
  jxor g11588(.dina(n11647), .dinb(n11646), .dout(n11656));
  jand g11589(.dina(n11656), .dinb(n11655), .dout(n11657));
  jor  g11590(.dina(n11657), .dinb(n11648), .dout(n11658));
  jand g11591(.dina(n11505), .dinb(n11497), .dout(n11659));
  jand g11592(.dina(n11618), .dinb(n11506), .dout(n11660));
  jor  g11593(.dina(n11660), .dinb(n11659), .dout(n11661));
  jand g11594(.dina(n11616), .dinb(n11608), .dout(n11662));
  jand g11595(.dina(n11617), .dinb(n11511), .dout(n11663));
  jor  g11596(.dina(n11663), .dinb(n11662), .dout(n11664));
  jand g11597(.dina(n11606), .dinb(n11598), .dout(n11665));
  jand g11598(.dina(n11607), .dinb(n11514), .dout(n11666));
  jor  g11599(.dina(n11666), .dinb(n11665), .dout(n11667));
  jor  g11600(.dina(n11596), .dinb(n11588), .dout(n11668));
  jand g11601(.dina(n11597), .dinb(n11519), .dout(n11669));
  jnot g11602(.din(n11669), .dout(n11670));
  jand g11603(.dina(n11670), .dinb(n11668), .dout(n11671));
  jnot g11604(.din(n11671), .dout(n11672));
  jor  g11605(.dina(n11585), .dinb(n11577), .dout(n11673));
  jand g11606(.dina(n11586), .dinb(n11524), .dout(n11674));
  jnot g11607(.din(n11674), .dout(n11675));
  jand g11608(.dina(n11675), .dinb(n11673), .dout(n11676));
  jnot g11609(.din(n11676), .dout(n11677));
  jor  g11610(.dina(n11574), .dinb(n11570), .dout(n11678));
  jand g11611(.dina(n11575), .dinb(n11533), .dout(n11679));
  jnot g11612(.din(n11679), .dout(n11680));
  jand g11613(.dina(n11680), .dinb(n11678), .dout(n11681));
  jnot g11614(.din(n11681), .dout(n11682));
  jor  g11615(.dina(n7061), .dinb(n4473), .dout(n11683));
  jand g11616(.dina(n6050), .dinb(n3930), .dout(n11684));
  jand g11617(.dina(n5084), .dinb(n4600), .dout(n11685));
  jor  g11618(.dina(n11685), .dinb(n11684), .dout(n11686));
  jand g11619(.dina(n5082), .dinb(n4406), .dout(n11687));
  jor  g11620(.dina(n11687), .dinb(n11686), .dout(n11688));
  jnot g11621(.din(n11688), .dout(n11689));
  jand g11622(.dina(n11689), .dinb(n11683), .dout(n11690));
  jnot g11623(.din(n11690), .dout(n11691));
  jand g11624(.dina(n621), .dinb(n452), .dout(n11692));
  jand g11625(.dina(n11692), .dinb(n1327), .dout(n11693));
  jand g11626(.dina(n11693), .dinb(n4544), .dout(n11694));
  jand g11627(.dina(n11694), .dinb(n2423), .dout(n11695));
  jand g11628(.dina(n11695), .dinb(n7503), .dout(n11696));
  jand g11629(.dina(n11696), .dinb(n1876), .dout(n11697));
  jand g11630(.dina(n1453), .dinb(n328), .dout(n11698));
  jand g11631(.dina(n11698), .dinb(n10384), .dout(n11699));
  jand g11632(.dina(n10718), .dinb(n3178), .dout(n11700));
  jand g11633(.dina(n11700), .dinb(n11699), .dout(n11701));
  jand g11634(.dina(n1981), .dinb(n1233), .dout(n11702));
  jand g11635(.dina(n11702), .dinb(n11701), .dout(n11703));
  jand g11636(.dina(n11703), .dinb(n11234), .dout(n11704));
  jand g11637(.dina(n11704), .dinb(n11697), .dout(n11705));
  jand g11638(.dina(n11705), .dinb(n2413), .dout(n11706));
  jand g11639(.dina(n1731), .dinb(n560), .dout(n11707));
  jand g11640(.dina(n11707), .dinb(n9327), .dout(n11708));
  jand g11641(.dina(n950), .dinb(n811), .dout(n11709));
  jand g11642(.dina(n11709), .dinb(n1438), .dout(n11710));
  jand g11643(.dina(n1393), .dinb(n456), .dout(n11711));
  jand g11644(.dina(n11711), .dinb(n11710), .dout(n11712));
  jand g11645(.dina(n11712), .dinb(n2599), .dout(n11713));
  jand g11646(.dina(n991), .dinb(n1291), .dout(n11714));
  jand g11647(.dina(n668), .dinb(n600), .dout(n11715));
  jand g11648(.dina(n11715), .dinb(n693), .dout(n11716));
  jand g11649(.dina(n11716), .dinb(n11714), .dout(n11717));
  jand g11650(.dina(n11717), .dinb(n1738), .dout(n11718));
  jand g11651(.dina(n11718), .dinb(n11713), .dout(n11719));
  jand g11652(.dina(n11719), .dinb(n11708), .dout(n11720));
  jand g11653(.dina(n925), .dinb(n916), .dout(n11721));
  jand g11654(.dina(n2659), .dinb(n721), .dout(n11722));
  jand g11655(.dina(n11722), .dinb(n11721), .dout(n11723));
  jand g11656(.dina(n11723), .dinb(n11720), .dout(n11724));
  jand g11657(.dina(n11724), .dinb(n1721), .dout(n11725));
  jand g11658(.dina(n11725), .dinb(n11706), .dout(n11726));
  jand g11659(.dina(n5170), .dinb(n833), .dout(n11727));
  jand g11660(.dina(n11727), .dinb(n519), .dout(n11728));
  jand g11661(.dina(n1912), .dinb(n175), .dout(n11729));
  jand g11662(.dina(n3066), .dinb(n1378), .dout(n11730));
  jand g11663(.dina(n11730), .dinb(n11729), .dout(n11731));
  jand g11664(.dina(n11731), .dinb(n1992), .dout(n11732));
  jand g11665(.dina(n11732), .dinb(n1596), .dout(n11733));
  jand g11666(.dina(n11733), .dinb(n11728), .dout(n11734));
  jand g11667(.dina(n11734), .dinb(n11208), .dout(n11735));
  jand g11668(.dina(n11735), .dinb(n11726), .dout(n11736));
  jnot g11669(.din(n11736), .dout(n11737));
  jxor g11670(.dina(n11737), .dinb(n11567), .dout(n11738));
  jxor g11671(.dina(n11738), .dinb(n11691), .dout(n11739));
  jxor g11672(.dina(n11739), .dinb(n11682), .dout(n11740));
  jnot g11673(.din(n11740), .dout(n11741));
  jor  g11674(.dina(n4688), .dinb(n4343), .dout(n11742));
  jor  g11675(.dina(n4526), .dinb(n4346), .dout(n11743));
  jor  g11676(.dina(n4686), .dinb(n4348), .dout(n11744));
  jand g11677(.dina(n11744), .dinb(n11743), .dout(n11745));
  jor  g11678(.dina(n4596), .dinb(n3683), .dout(n11746));
  jand g11679(.dina(n11746), .dinb(n11745), .dout(n11747));
  jand g11680(.dina(n11747), .dinb(n11742), .dout(n11748));
  jxor g11681(.dina(n11748), .dinb(\a[29] ), .dout(n11749));
  jxor g11682(.dina(n11749), .dinb(n11741), .dout(n11750));
  jxor g11683(.dina(n11750), .dinb(n11677), .dout(n11751));
  jnot g11684(.din(n11751), .dout(n11752));
  jor  g11685(.dina(n5264), .dinb(n1805), .dout(n11753));
  jor  g11686(.dina(n5549), .dinb(n2303), .dout(n11754));
  jor  g11687(.dina(n5364), .dinb(n2309), .dout(n11755));
  jor  g11688(.dina(n5422), .dinb(n2306), .dout(n11756));
  jand g11689(.dina(n11756), .dinb(n11755), .dout(n11757));
  jand g11690(.dina(n11757), .dinb(n11754), .dout(n11758));
  jand g11691(.dina(n11758), .dinb(n11753), .dout(n11759));
  jxor g11692(.dina(n11759), .dinb(\a[26] ), .dout(n11760));
  jxor g11693(.dina(n11760), .dinb(n11752), .dout(n11761));
  jxor g11694(.dina(n11761), .dinb(n11672), .dout(n11762));
  jor  g11695(.dina(n6516), .dinb(n807), .dout(n11763));
  jor  g11696(.dina(n6205), .dinb(n1613), .dout(n11764));
  jor  g11697(.dina(n6390), .dinb(n1621), .dout(n11765));
  jor  g11698(.dina(n5525), .dinb(n1617), .dout(n11766));
  jand g11699(.dina(n11766), .dinb(n11765), .dout(n11767));
  jand g11700(.dina(n11767), .dinb(n11764), .dout(n11768));
  jand g11701(.dina(n11768), .dinb(n11763), .dout(n11769));
  jxor g11702(.dina(n11769), .dinb(n65), .dout(n11770));
  jxor g11703(.dina(n11770), .dinb(n11762), .dout(n11771));
  jxor g11704(.dina(n11771), .dinb(n11667), .dout(n11772));
  jnot g11705(.din(n11772), .dout(n11773));
  jor  g11706(.dina(n7301), .dinb(n2189), .dout(n11774));
  jor  g11707(.dina(n7303), .dinb(n1820), .dout(n11775));
  jor  g11708(.dina(n6297), .dinb(n2186), .dout(n11776));
  jor  g11709(.dina(n6489), .dinb(n2181), .dout(n11777));
  jand g11710(.dina(n11777), .dinb(n11776), .dout(n11778));
  jand g11711(.dina(n11778), .dinb(n11775), .dout(n11779));
  jand g11712(.dina(n11779), .dinb(n11774), .dout(n11780));
  jxor g11713(.dina(n11780), .dinb(\a[20] ), .dout(n11781));
  jxor g11714(.dina(n11781), .dinb(n11773), .dout(n11782));
  jxor g11715(.dina(n11782), .dinb(n11664), .dout(n11783));
  jnot g11716(.din(n11783), .dout(n11784));
  jor  g11717(.dina(n8260), .dinb(n2744), .dout(n11785));
  jor  g11718(.dina(n7680), .dinb(n2758), .dout(n11786));
  jor  g11719(.dina(n7999), .dinb(n2749), .dout(n11787));
  jand g11720(.dina(n11787), .dinb(n11786), .dout(n11788));
  jand g11721(.dina(n11788), .dinb(n11785), .dout(n11789));
  jxor g11722(.dina(n11789), .dinb(\a[17] ), .dout(n11790));
  jxor g11723(.dina(n11790), .dinb(n11784), .dout(n11791));
  jxor g11724(.dina(n11791), .dinb(n11661), .dout(n11792));
  jnot g11725(.din(n11792), .dout(n11793));
  jand g11726(.dina(n11619), .dinb(n11494), .dout(n11794));
  jnot g11727(.din(n11794), .dout(n11795));
  jor  g11728(.dina(n11645), .dinb(n11621), .dout(n11796));
  jand g11729(.dina(n11796), .dinb(n11795), .dout(n11797));
  jxor g11730(.dina(n11797), .dinb(n11793), .dout(n11798));
  jxor g11731(.dina(n11798), .dinb(n11646), .dout(n11799));
  jxor g11732(.dina(n11799), .dinb(n11658), .dout(n11800));
  jand g11733(.dina(n11800), .dinb(n4022), .dout(n11801));
  jand g11734(.dina(n11798), .dinb(n4220), .dout(n11802));
  jand g11735(.dina(n11646), .dinb(n4027), .dout(n11803));
  jand g11736(.dina(n11647), .dinb(n3870), .dout(n11804));
  jor  g11737(.dina(n11804), .dinb(n11803), .dout(n11805));
  jor  g11738(.dina(n11805), .dinb(n11802), .dout(n11806));
  jor  g11739(.dina(n11806), .dinb(n11801), .dout(n11807));
  jxor g11740(.dina(n11807), .dinb(n4050), .dout(n11808));
  jor  g11741(.dina(n11808), .dinb(n11320), .dout(n11809));
  jxor g11742(.dina(n11056), .dinb(n11054), .dout(n11810));
  jnot g11743(.din(n11810), .dout(n11811));
  jxor g11744(.dina(n11656), .dinb(n11655), .dout(n11812));
  jand g11745(.dina(n11812), .dinb(n4022), .dout(n11813));
  jand g11746(.dina(n11646), .dinb(n4220), .dout(n11814));
  jand g11747(.dina(n11647), .dinb(n4027), .dout(n11815));
  jand g11748(.dina(n11306), .dinb(n3870), .dout(n11816));
  jor  g11749(.dina(n11816), .dinb(n11815), .dout(n11817));
  jor  g11750(.dina(n11817), .dinb(n11814), .dout(n11818));
  jor  g11751(.dina(n11818), .dinb(n11813), .dout(n11819));
  jxor g11752(.dina(n11819), .dinb(n4050), .dout(n11820));
  jor  g11753(.dina(n11820), .dinb(n11811), .dout(n11821));
  jxor g11754(.dina(n11051), .dinb(n11050), .dout(n11822));
  jnot g11755(.din(n11822), .dout(n11823));
  jxor g11756(.dina(n11653), .dinb(n11652), .dout(n11824));
  jand g11757(.dina(n11824), .dinb(n4022), .dout(n11825));
  jand g11758(.dina(n11647), .dinb(n4220), .dout(n11826));
  jand g11759(.dina(n11306), .dinb(n4027), .dout(n11827));
  jand g11760(.dina(n10836), .dinb(n3870), .dout(n11828));
  jor  g11761(.dina(n11828), .dinb(n11827), .dout(n11829));
  jor  g11762(.dina(n11829), .dinb(n11826), .dout(n11830));
  jor  g11763(.dina(n11830), .dinb(n11825), .dout(n11831));
  jxor g11764(.dina(n11831), .dinb(n4050), .dout(n11832));
  jor  g11765(.dina(n11832), .dinb(n11823), .dout(n11833));
  jxor g11766(.dina(n11046), .dinb(n11045), .dout(n11834));
  jnot g11767(.din(n11834), .dout(n11835));
  jand g11768(.dina(n11308), .dinb(n4022), .dout(n11836));
  jand g11769(.dina(n10836), .dinb(n4027), .dout(n11837));
  jand g11770(.dina(n11306), .dinb(n4220), .dout(n11838));
  jor  g11771(.dina(n11838), .dinb(n11837), .dout(n11839));
  jand g11772(.dina(n10640), .dinb(n3870), .dout(n11840));
  jor  g11773(.dina(n11840), .dinb(n11839), .dout(n11841));
  jor  g11774(.dina(n11841), .dinb(n11836), .dout(n11842));
  jxor g11775(.dina(n11842), .dinb(n4050), .dout(n11843));
  jor  g11776(.dina(n11843), .dinb(n11835), .dout(n11844));
  jxor g11777(.dina(n11043), .dinb(n11042), .dout(n11845));
  jnot g11778(.din(n11845), .dout(n11846));
  jand g11779(.dina(n10838), .dinb(n4022), .dout(n11847));
  jand g11780(.dina(n10640), .dinb(n4027), .dout(n11848));
  jand g11781(.dina(n10836), .dinb(n4220), .dout(n11849));
  jor  g11782(.dina(n11849), .dinb(n11848), .dout(n11850));
  jand g11783(.dina(n10647), .dinb(n3870), .dout(n11851));
  jor  g11784(.dina(n11851), .dinb(n11850), .dout(n11852));
  jor  g11785(.dina(n11852), .dinb(n11847), .dout(n11853));
  jxor g11786(.dina(n11853), .dinb(n4050), .dout(n11854));
  jor  g11787(.dina(n11854), .dinb(n11846), .dout(n11855));
  jxor g11788(.dina(n11038), .dinb(n11037), .dout(n11856));
  jnot g11789(.din(n11856), .dout(n11857));
  jand g11790(.dina(n10850), .dinb(n4022), .dout(n11858));
  jand g11791(.dina(n10647), .dinb(n4027), .dout(n11859));
  jand g11792(.dina(n10640), .dinb(n4220), .dout(n11860));
  jor  g11793(.dina(n11860), .dinb(n11859), .dout(n11861));
  jand g11794(.dina(n10305), .dinb(n3870), .dout(n11862));
  jor  g11795(.dina(n11862), .dinb(n11861), .dout(n11863));
  jor  g11796(.dina(n11863), .dinb(n11858), .dout(n11864));
  jxor g11797(.dina(n11864), .dinb(n4050), .dout(n11865));
  jor  g11798(.dina(n11865), .dinb(n11857), .dout(n11866));
  jxor g11799(.dina(n11033), .dinb(n11032), .dout(n11867));
  jnot g11800(.din(n11867), .dout(n11868));
  jand g11801(.dina(n10862), .dinb(n4022), .dout(n11869));
  jand g11802(.dina(n10305), .dinb(n4027), .dout(n11870));
  jand g11803(.dina(n10647), .dinb(n4220), .dout(n11871));
  jor  g11804(.dina(n11871), .dinb(n11870), .dout(n11872));
  jand g11805(.dina(n9872), .dinb(n3870), .dout(n11873));
  jor  g11806(.dina(n11873), .dinb(n11872), .dout(n11874));
  jor  g11807(.dina(n11874), .dinb(n11869), .dout(n11875));
  jxor g11808(.dina(n11875), .dinb(n4050), .dout(n11876));
  jor  g11809(.dina(n11876), .dinb(n11868), .dout(n11877));
  jxor g11810(.dina(n11028), .dinb(n11027), .dout(n11878));
  jnot g11811(.din(n11878), .dout(n11879));
  jand g11812(.dina(n10307), .dinb(n4022), .dout(n11880));
  jand g11813(.dina(n10305), .dinb(n4220), .dout(n11881));
  jand g11814(.dina(n9872), .dinb(n4027), .dout(n11882));
  jand g11815(.dina(n9655), .dinb(n3870), .dout(n11883));
  jor  g11816(.dina(n11883), .dinb(n11882), .dout(n11884));
  jor  g11817(.dina(n11884), .dinb(n11881), .dout(n11885));
  jor  g11818(.dina(n11885), .dinb(n11880), .dout(n11886));
  jxor g11819(.dina(n11886), .dinb(n4050), .dout(n11887));
  jor  g11820(.dina(n11887), .dinb(n11879), .dout(n11888));
  jxor g11821(.dina(n11023), .dinb(n11022), .dout(n11889));
  jnot g11822(.din(n11889), .dout(n11890));
  jand g11823(.dina(n9874), .dinb(n4022), .dout(n11891));
  jand g11824(.dina(n9655), .dinb(n4027), .dout(n11892));
  jand g11825(.dina(n9872), .dinb(n4220), .dout(n11893));
  jor  g11826(.dina(n11893), .dinb(n11892), .dout(n11894));
  jand g11827(.dina(n9656), .dinb(n3870), .dout(n11895));
  jor  g11828(.dina(n11895), .dinb(n11894), .dout(n11896));
  jor  g11829(.dina(n11896), .dinb(n11891), .dout(n11897));
  jxor g11830(.dina(n11897), .dinb(n4050), .dout(n11898));
  jor  g11831(.dina(n11898), .dinb(n11890), .dout(n11899));
  jxor g11832(.dina(n11018), .dinb(n11017), .dout(n11900));
  jnot g11833(.din(n11900), .dout(n11901));
  jand g11834(.dina(n9886), .dinb(n4022), .dout(n11902));
  jand g11835(.dina(n9655), .dinb(n4220), .dout(n11903));
  jand g11836(.dina(n9656), .dinb(n4027), .dout(n11904));
  jand g11837(.dina(n9250), .dinb(n3870), .dout(n11905));
  jor  g11838(.dina(n11905), .dinb(n11904), .dout(n11906));
  jor  g11839(.dina(n11906), .dinb(n11903), .dout(n11907));
  jor  g11840(.dina(n11907), .dinb(n11902), .dout(n11908));
  jxor g11841(.dina(n11908), .dinb(n4050), .dout(n11909));
  jor  g11842(.dina(n11909), .dinb(n11901), .dout(n11910));
  jxor g11843(.dina(n11013), .dinb(n11012), .dout(n11911));
  jnot g11844(.din(n11911), .dout(n11912));
  jand g11845(.dina(n9898), .dinb(n4022), .dout(n11913));
  jand g11846(.dina(n9250), .dinb(n4027), .dout(n11914));
  jand g11847(.dina(n9656), .dinb(n4220), .dout(n11915));
  jor  g11848(.dina(n11915), .dinb(n11914), .dout(n11916));
  jand g11849(.dina(n8936), .dinb(n3870), .dout(n11917));
  jor  g11850(.dina(n11917), .dinb(n11916), .dout(n11918));
  jor  g11851(.dina(n11918), .dinb(n11913), .dout(n11919));
  jxor g11852(.dina(n11919), .dinb(n4050), .dout(n11920));
  jor  g11853(.dina(n11920), .dinb(n11912), .dout(n11921));
  jxor g11854(.dina(n11010), .dinb(n11009), .dout(n11922));
  jnot g11855(.din(n11922), .dout(n11923));
  jand g11856(.dina(n9252), .dinb(n4022), .dout(n11924));
  jand g11857(.dina(n9250), .dinb(n4220), .dout(n11925));
  jand g11858(.dina(n8936), .dinb(n4027), .dout(n11926));
  jand g11859(.dina(n8723), .dinb(n3870), .dout(n11927));
  jor  g11860(.dina(n11927), .dinb(n11926), .dout(n11928));
  jor  g11861(.dina(n11928), .dinb(n11925), .dout(n11929));
  jor  g11862(.dina(n11929), .dinb(n11924), .dout(n11930));
  jxor g11863(.dina(n11930), .dinb(n4050), .dout(n11931));
  jor  g11864(.dina(n11931), .dinb(n11923), .dout(n11932));
  jxor g11865(.dina(n11005), .dinb(n11004), .dout(n11933));
  jnot g11866(.din(n11933), .dout(n11934));
  jand g11867(.dina(n8938), .dinb(n4022), .dout(n11935));
  jand g11868(.dina(n8723), .dinb(n4027), .dout(n11936));
  jand g11869(.dina(n8936), .dinb(n4220), .dout(n11937));
  jor  g11870(.dina(n11937), .dinb(n11936), .dout(n11938));
  jand g11871(.dina(n8740), .dinb(n3870), .dout(n11939));
  jor  g11872(.dina(n11939), .dinb(n11938), .dout(n11940));
  jor  g11873(.dina(n11940), .dinb(n11935), .dout(n11941));
  jxor g11874(.dina(n11941), .dinb(n4050), .dout(n11942));
  jor  g11875(.dina(n11942), .dinb(n11934), .dout(n11943));
  jxor g11876(.dina(n11001), .dinb(n10993), .dout(n11944));
  jnot g11877(.din(n11944), .dout(n11945));
  jand g11878(.dina(n8950), .dinb(n4022), .dout(n11946));
  jand g11879(.dina(n8740), .dinb(n4027), .dout(n11947));
  jand g11880(.dina(n8723), .dinb(n4220), .dout(n11948));
  jor  g11881(.dina(n11948), .dinb(n11947), .dout(n11949));
  jand g11882(.dina(n8268), .dinb(n3870), .dout(n11950));
  jor  g11883(.dina(n11950), .dinb(n11949), .dout(n11951));
  jor  g11884(.dina(n11951), .dinb(n11946), .dout(n11952));
  jxor g11885(.dina(n11952), .dinb(n4050), .dout(n11953));
  jor  g11886(.dina(n11953), .dinb(n11945), .dout(n11954));
  jor  g11887(.dina(n10980), .dinb(n3473), .dout(n11955));
  jxor g11888(.dina(n11955), .dinb(n10988), .dout(n11956));
  jand g11889(.dina(n8962), .dinb(n4022), .dout(n11957));
  jand g11890(.dina(n8740), .dinb(n4220), .dout(n11958));
  jand g11891(.dina(n8268), .dinb(n4027), .dout(n11959));
  jand g11892(.dina(n8022), .dinb(n3870), .dout(n11960));
  jor  g11893(.dina(n11960), .dinb(n11959), .dout(n11961));
  jor  g11894(.dina(n11961), .dinb(n11958), .dout(n11962));
  jor  g11895(.dina(n11962), .dinb(n11957), .dout(n11963));
  jxor g11896(.dina(n11963), .dinb(\a[11] ), .dout(n11964));
  jand g11897(.dina(n11964), .dinb(n11956), .dout(n11965));
  jand g11898(.dina(n10977), .dinb(\a[14] ), .dout(n11966));
  jxor g11899(.dina(n11966), .dinb(n10975), .dout(n11967));
  jnot g11900(.din(n11967), .dout(n11968));
  jand g11901(.dina(n8270), .dinb(n4022), .dout(n11969));
  jand g11902(.dina(n8022), .dinb(n4027), .dout(n11970));
  jand g11903(.dina(n8268), .dinb(n4220), .dout(n11971));
  jor  g11904(.dina(n11971), .dinb(n11970), .dout(n11972));
  jand g11905(.dina(n7692), .dinb(n3870), .dout(n11973));
  jor  g11906(.dina(n11973), .dinb(n11972), .dout(n11974));
  jor  g11907(.dina(n11974), .dinb(n11969), .dout(n11975));
  jxor g11908(.dina(n11975), .dinb(n4050), .dout(n11976));
  jor  g11909(.dina(n11976), .dinb(n11968), .dout(n11977));
  jand g11910(.dina(n7315), .dinb(n4022), .dout(n11978));
  jand g11911(.dina(n7019), .dinb(n4027), .dout(n11979));
  jand g11912(.dina(n7313), .dinb(n4220), .dout(n11980));
  jor  g11913(.dina(n11980), .dinb(n11979), .dout(n11981));
  jor  g11914(.dina(n11981), .dinb(n11978), .dout(n11982));
  jnot g11915(.din(n11982), .dout(n11983));
  jand g11916(.dina(n7019), .dinb(n3865), .dout(n11984));
  jnot g11917(.din(n11984), .dout(n11985));
  jand g11918(.dina(n11985), .dinb(\a[11] ), .dout(n11986));
  jand g11919(.dina(n11986), .dinb(n11983), .dout(n11987));
  jand g11920(.dina(n7693), .dinb(n4022), .dout(n11988));
  jand g11921(.dina(n7313), .dinb(n4027), .dout(n11989));
  jor  g11922(.dina(n11989), .dinb(n11988), .dout(n11990));
  jand g11923(.dina(n7692), .dinb(n4220), .dout(n11991));
  jand g11924(.dina(n7019), .dinb(n3870), .dout(n11992));
  jor  g11925(.dina(n11992), .dinb(n11991), .dout(n11993));
  jor  g11926(.dina(n11993), .dinb(n11990), .dout(n11994));
  jnot g11927(.din(n11994), .dout(n11995));
  jand g11928(.dina(n11995), .dinb(n11987), .dout(n11996));
  jand g11929(.dina(n11996), .dinb(n10977), .dout(n11997));
  jnot g11930(.din(n11997), .dout(n11998));
  jxor g11931(.dina(n11996), .dinb(n10977), .dout(n11999));
  jnot g11932(.din(n11999), .dout(n12000));
  jand g11933(.dina(n8029), .dinb(n4022), .dout(n12001));
  jand g11934(.dina(n7692), .dinb(n4027), .dout(n12002));
  jand g11935(.dina(n8022), .dinb(n4220), .dout(n12003));
  jor  g11936(.dina(n12003), .dinb(n12002), .dout(n12004));
  jand g11937(.dina(n7313), .dinb(n3870), .dout(n12005));
  jor  g11938(.dina(n12005), .dinb(n12004), .dout(n12006));
  jor  g11939(.dina(n12006), .dinb(n12001), .dout(n12007));
  jxor g11940(.dina(n12007), .dinb(n4050), .dout(n12008));
  jor  g11941(.dina(n12008), .dinb(n12000), .dout(n12009));
  jand g11942(.dina(n12009), .dinb(n11998), .dout(n12010));
  jnot g11943(.din(n12010), .dout(n12011));
  jxor g11944(.dina(n11976), .dinb(n11968), .dout(n12012));
  jand g11945(.dina(n12012), .dinb(n12011), .dout(n12013));
  jnot g11946(.din(n12013), .dout(n12014));
  jand g11947(.dina(n12014), .dinb(n11977), .dout(n12015));
  jnot g11948(.din(n12015), .dout(n12016));
  jxor g11949(.dina(n11964), .dinb(n11956), .dout(n12017));
  jand g11950(.dina(n12017), .dinb(n12016), .dout(n12018));
  jor  g11951(.dina(n12018), .dinb(n11965), .dout(n12019));
  jxor g11952(.dina(n11953), .dinb(n11945), .dout(n12020));
  jand g11953(.dina(n12020), .dinb(n12019), .dout(n12021));
  jnot g11954(.din(n12021), .dout(n12022));
  jand g11955(.dina(n12022), .dinb(n11954), .dout(n12023));
  jnot g11956(.din(n12023), .dout(n12024));
  jxor g11957(.dina(n11942), .dinb(n11934), .dout(n12025));
  jand g11958(.dina(n12025), .dinb(n12024), .dout(n12026));
  jnot g11959(.din(n12026), .dout(n12027));
  jand g11960(.dina(n12027), .dinb(n11943), .dout(n12028));
  jnot g11961(.din(n12028), .dout(n12029));
  jxor g11962(.dina(n11931), .dinb(n11923), .dout(n12030));
  jand g11963(.dina(n12030), .dinb(n12029), .dout(n12031));
  jnot g11964(.din(n12031), .dout(n12032));
  jand g11965(.dina(n12032), .dinb(n11932), .dout(n12033));
  jnot g11966(.din(n12033), .dout(n12034));
  jxor g11967(.dina(n11920), .dinb(n11912), .dout(n12035));
  jand g11968(.dina(n12035), .dinb(n12034), .dout(n12036));
  jnot g11969(.din(n12036), .dout(n12037));
  jand g11970(.dina(n12037), .dinb(n11921), .dout(n12038));
  jnot g11971(.din(n12038), .dout(n12039));
  jxor g11972(.dina(n11909), .dinb(n11901), .dout(n12040));
  jand g11973(.dina(n12040), .dinb(n12039), .dout(n12041));
  jnot g11974(.din(n12041), .dout(n12042));
  jand g11975(.dina(n12042), .dinb(n11910), .dout(n12043));
  jnot g11976(.din(n12043), .dout(n12044));
  jxor g11977(.dina(n11898), .dinb(n11890), .dout(n12045));
  jand g11978(.dina(n12045), .dinb(n12044), .dout(n12046));
  jnot g11979(.din(n12046), .dout(n12047));
  jand g11980(.dina(n12047), .dinb(n11899), .dout(n12048));
  jxor g11981(.dina(n11887), .dinb(n11879), .dout(n12049));
  jnot g11982(.din(n12049), .dout(n12050));
  jor  g11983(.dina(n12050), .dinb(n12048), .dout(n12051));
  jand g11984(.dina(n12051), .dinb(n11888), .dout(n12052));
  jxor g11985(.dina(n11876), .dinb(n11868), .dout(n12053));
  jnot g11986(.din(n12053), .dout(n12054));
  jor  g11987(.dina(n12054), .dinb(n12052), .dout(n12055));
  jand g11988(.dina(n12055), .dinb(n11877), .dout(n12056));
  jxor g11989(.dina(n11865), .dinb(n11857), .dout(n12057));
  jnot g11990(.din(n12057), .dout(n12058));
  jor  g11991(.dina(n12058), .dinb(n12056), .dout(n12059));
  jand g11992(.dina(n12059), .dinb(n11866), .dout(n12060));
  jxor g11993(.dina(n11854), .dinb(n11846), .dout(n12061));
  jnot g11994(.din(n12061), .dout(n12062));
  jor  g11995(.dina(n12062), .dinb(n12060), .dout(n12063));
  jand g11996(.dina(n12063), .dinb(n11855), .dout(n12064));
  jxor g11997(.dina(n11843), .dinb(n11835), .dout(n12065));
  jnot g11998(.din(n12065), .dout(n12066));
  jor  g11999(.dina(n12066), .dinb(n12064), .dout(n12067));
  jand g12000(.dina(n12067), .dinb(n11844), .dout(n12068));
  jxor g12001(.dina(n11832), .dinb(n11823), .dout(n12069));
  jnot g12002(.din(n12069), .dout(n12070));
  jor  g12003(.dina(n12070), .dinb(n12068), .dout(n12071));
  jand g12004(.dina(n12071), .dinb(n11833), .dout(n12072));
  jxor g12005(.dina(n11820), .dinb(n11810), .dout(n12073));
  jor  g12006(.dina(n12073), .dinb(n12072), .dout(n12074));
  jand g12007(.dina(n12074), .dinb(n11821), .dout(n12075));
  jxor g12008(.dina(n11808), .dinb(n11319), .dout(n12076));
  jor  g12009(.dina(n12076), .dinb(n12075), .dout(n12077));
  jand g12010(.dina(n12077), .dinb(n11809), .dout(n12078));
  jor  g12011(.dina(n11316), .dinb(n11130), .dout(n12079));
  jor  g12012(.dina(n11318), .dinb(n11058), .dout(n12080));
  jand g12013(.dina(n12080), .dinb(n12079), .dout(n12081));
  jor  g12014(.dina(n11127), .dinb(n11119), .dout(n12082));
  jand g12015(.dina(n11128), .dinb(n11063), .dout(n12083));
  jnot g12016(.din(n12083), .dout(n12084));
  jand g12017(.dina(n12084), .dinb(n12082), .dout(n12085));
  jnot g12018(.din(n12085), .dout(n12086));
  jor  g12019(.dina(n11116), .dinb(n11108), .dout(n12087));
  jand g12020(.dina(n11117), .dinb(n11068), .dout(n12088));
  jnot g12021(.din(n12088), .dout(n12089));
  jand g12022(.dina(n12089), .dinb(n12087), .dout(n12090));
  jnot g12023(.din(n12090), .dout(n12091));
  jor  g12024(.dina(n11105), .dinb(n11097), .dout(n12092));
  jand g12025(.dina(n11106), .dinb(n11073), .dout(n12093));
  jnot g12026(.din(n12093), .dout(n12094));
  jand g12027(.dina(n12094), .dinb(n12092), .dout(n12095));
  jnot g12028(.din(n12095), .dout(n12096));
  jor  g12029(.dina(n11094), .dinb(n11086), .dout(n12097));
  jand g12030(.dina(n11095), .dinb(n11079), .dout(n12098));
  jnot g12031(.din(n12098), .dout(n12099));
  jand g12032(.dina(n12099), .dinb(n12097), .dout(n12100));
  jnot g12033(.din(n12100), .dout(n12101));
  jand g12034(.dina(n7693), .dinb(n2936), .dout(n12102));
  jand g12035(.dina(n7313), .dinb(n2940), .dout(n12103));
  jand g12036(.dina(n7692), .dinb(n2943), .dout(n12104));
  jor  g12037(.dina(n12104), .dinb(n12103), .dout(n12105));
  jand g12038(.dina(n7019), .dinb(n3684), .dout(n12106));
  jor  g12039(.dina(n12106), .dinb(n12105), .dout(n12107));
  jor  g12040(.dina(n12107), .dinb(n12102), .dout(n12108));
  jnot g12041(.din(n11084), .dout(n12109));
  jand g12042(.dina(n10046), .dinb(\a[29] ), .dout(n12110));
  jand g12043(.dina(n12110), .dinb(n12109), .dout(n12111));
  jnot g12044(.din(n12111), .dout(n12112));
  jand g12045(.dina(n12112), .dinb(\a[29] ), .dout(n12113));
  jxor g12046(.dina(n12113), .dinb(n12108), .dout(n12114));
  jand g12047(.dina(n8962), .dinb(n71), .dout(n12115));
  jand g12048(.dina(n8740), .dinb(n796), .dout(n12116));
  jand g12049(.dina(n8268), .dinb(n731), .dout(n12117));
  jand g12050(.dina(n8022), .dinb(n1806), .dout(n12118));
  jor  g12051(.dina(n12118), .dinb(n12117), .dout(n12119));
  jor  g12052(.dina(n12119), .dinb(n12116), .dout(n12120));
  jor  g12053(.dina(n12120), .dinb(n12115), .dout(n12121));
  jxor g12054(.dina(n12121), .dinb(\a[26] ), .dout(n12122));
  jxor g12055(.dina(n12122), .dinb(n12114), .dout(n12123));
  jxor g12056(.dina(n12123), .dinb(n12101), .dout(n12124));
  jnot g12057(.din(n12124), .dout(n12125));
  jand g12058(.dina(n9252), .dinb(n806), .dout(n12126));
  jand g12059(.dina(n9250), .dinb(n1620), .dout(n12127));
  jand g12060(.dina(n8936), .dinb(n1612), .dout(n12128));
  jand g12061(.dina(n8723), .dinb(n1644), .dout(n12129));
  jor  g12062(.dina(n12129), .dinb(n12128), .dout(n12130));
  jor  g12063(.dina(n12130), .dinb(n12127), .dout(n12131));
  jor  g12064(.dina(n12131), .dinb(n12126), .dout(n12132));
  jxor g12065(.dina(n12132), .dinb(n65), .dout(n12133));
  jxor g12066(.dina(n12133), .dinb(n12125), .dout(n12134));
  jxor g12067(.dina(n12134), .dinb(n12096), .dout(n12135));
  jand g12068(.dina(n9874), .dinb(n1819), .dout(n12136));
  jand g12069(.dina(n9872), .dinb(n2243), .dout(n12137));
  jand g12070(.dina(n9655), .dinb(n2180), .dout(n12138));
  jand g12071(.dina(n9656), .dinb(n2185), .dout(n12139));
  jor  g12072(.dina(n12139), .dinb(n12138), .dout(n12140));
  jor  g12073(.dina(n12140), .dinb(n12137), .dout(n12141));
  jor  g12074(.dina(n12141), .dinb(n12136), .dout(n12142));
  jxor g12075(.dina(n12142), .dinb(\a[20] ), .dout(n12143));
  jxor g12076(.dina(n12143), .dinb(n12135), .dout(n12144));
  jxor g12077(.dina(n12144), .dinb(n12091), .dout(n12145));
  jnot g12078(.din(n12145), .dout(n12146));
  jand g12079(.dina(n10850), .dinb(n2743), .dout(n12147));
  jand g12080(.dina(n10640), .dinb(n2752), .dout(n12148));
  jand g12081(.dina(n10647), .dinb(n2748), .dout(n12149));
  jand g12082(.dina(n10305), .dinb(n2757), .dout(n12150));
  jor  g12083(.dina(n12150), .dinb(n12149), .dout(n12151));
  jor  g12084(.dina(n12151), .dinb(n12148), .dout(n12152));
  jor  g12085(.dina(n12152), .dinb(n12147), .dout(n12153));
  jxor g12086(.dina(n12153), .dinb(n2441), .dout(n12154));
  jxor g12087(.dina(n12154), .dinb(n12146), .dout(n12155));
  jxor g12088(.dina(n12155), .dinb(n12086), .dout(n12156));
  jnot g12089(.din(n12156), .dout(n12157));
  jand g12090(.dina(n11824), .dinb(n3423), .dout(n12158));
  jand g12091(.dina(n11306), .dinb(n3428), .dout(n12159));
  jand g12092(.dina(n11647), .dinb(n3569), .dout(n12160));
  jor  g12093(.dina(n12160), .dinb(n12159), .dout(n12161));
  jand g12094(.dina(n10836), .dinb(n3210), .dout(n12162));
  jor  g12095(.dina(n12162), .dinb(n12161), .dout(n12163));
  jor  g12096(.dina(n12163), .dinb(n12158), .dout(n12164));
  jxor g12097(.dina(n12164), .dinb(n3473), .dout(n12165));
  jxor g12098(.dina(n12165), .dinb(n12157), .dout(n12166));
  jxor g12099(.dina(n12166), .dinb(n12081), .dout(n12167));
  jand g12100(.dina(n11798), .dinb(n11646), .dout(n12168));
  jand g12101(.dina(n11799), .dinb(n11658), .dout(n12169));
  jor  g12102(.dina(n12169), .dinb(n12168), .dout(n12170));
  jand g12103(.dina(n11782), .dinb(n11664), .dout(n12171));
  jnot g12104(.din(n12171), .dout(n12172));
  jor  g12105(.dina(n11790), .dinb(n11784), .dout(n12173));
  jand g12106(.dina(n12173), .dinb(n12172), .dout(n12174));
  jnot g12107(.din(n12174), .dout(n12175));
  jand g12108(.dina(n11771), .dinb(n11667), .dout(n12176));
  jnot g12109(.din(n12176), .dout(n12177));
  jor  g12110(.dina(n11781), .dinb(n11773), .dout(n12178));
  jand g12111(.dina(n12178), .dinb(n12177), .dout(n12179));
  jand g12112(.dina(n8256), .dinb(n2743), .dout(n12180));
  jor  g12113(.dina(n12180), .dinb(n2757), .dout(n12181));
  jand g12114(.dina(n12181), .dinb(n8000), .dout(n12182));
  jxor g12115(.dina(n12182), .dinb(n2441), .dout(n12183));
  jxor g12116(.dina(n12183), .dinb(n12179), .dout(n12184));
  jand g12117(.dina(n11761), .dinb(n11672), .dout(n12185));
  jand g12118(.dina(n11770), .dinb(n11762), .dout(n12186));
  jor  g12119(.dina(n12186), .dinb(n12185), .dout(n12187));
  jand g12120(.dina(n11750), .dinb(n11677), .dout(n12188));
  jnot g12121(.din(n12188), .dout(n12189));
  jor  g12122(.dina(n11760), .dinb(n11752), .dout(n12190));
  jand g12123(.dina(n12190), .dinb(n12189), .dout(n12191));
  jnot g12124(.din(n12191), .dout(n12192));
  jand g12125(.dina(n11739), .dinb(n11682), .dout(n12193));
  jnot g12126(.din(n12193), .dout(n12194));
  jor  g12127(.dina(n11749), .dinb(n11741), .dout(n12195));
  jand g12128(.dina(n12195), .dinb(n12194), .dout(n12196));
  jnot g12129(.din(n12196), .dout(n12197));
  jor  g12130(.dina(n7061), .dinb(n4726), .dout(n12198));
  jand g12131(.dina(n6050), .dinb(n4406), .dout(n12199));
  jand g12132(.dina(n5084), .dinb(n4597), .dout(n12200));
  jor  g12133(.dina(n12200), .dinb(n12199), .dout(n12201));
  jand g12134(.dina(n5082), .dinb(n4600), .dout(n12202));
  jor  g12135(.dina(n12202), .dinb(n12201), .dout(n12203));
  jnot g12136(.din(n12203), .dout(n12204));
  jand g12137(.dina(n12204), .dinb(n12198), .dout(n12205));
  jnot g12138(.din(n12205), .dout(n12206));
  jnot g12139(.din(n11567), .dout(n12207));
  jand g12140(.dina(n11736), .dinb(n12207), .dout(n12208));
  jand g12141(.dina(n11738), .dinb(n11691), .dout(n12209));
  jor  g12142(.dina(n12209), .dinb(n12208), .dout(n12210));
  jand g12143(.dina(n11394), .dinb(n172), .dout(n12211));
  jand g12144(.dina(n12211), .dinb(n5300), .dout(n12212));
  jand g12145(.dina(n12212), .dinb(n1831), .dout(n12213));
  jand g12146(.dina(n5375), .dinb(n3900), .dout(n12214));
  jand g12147(.dina(n12214), .dinb(n1588), .dout(n12215));
  jand g12148(.dina(n12215), .dinb(n12213), .dout(n12216));
  jand g12149(.dina(n9764), .dinb(n1449), .dout(n12217));
  jand g12150(.dina(n12217), .dinb(n1317), .dout(n12218));
  jand g12151(.dina(n873), .dinb(n510), .dout(n12219));
  jand g12152(.dina(n12219), .dinb(n3195), .dout(n12220));
  jand g12153(.dina(n5206), .dinb(n554), .dout(n12221));
  jand g12154(.dina(n12221), .dinb(n12220), .dout(n12222));
  jand g12155(.dina(n12222), .dinb(n12218), .dout(n12223));
  jand g12156(.dina(n685), .dinb(n664), .dout(n12224));
  jand g12157(.dina(n12224), .dinb(n7269), .dout(n12225));
  jand g12158(.dina(n12225), .dinb(n12223), .dout(n12226));
  jand g12159(.dina(n12226), .dinb(n6447), .dout(n12227));
  jand g12160(.dina(n12227), .dinb(n6323), .dout(n12228));
  jand g12161(.dina(n12228), .dinb(n12216), .dout(n12229));
  jxor g12162(.dina(n12229), .dinb(n11737), .dout(n12230));
  jxor g12163(.dina(n12230), .dinb(n12210), .dout(n12231));
  jxor g12164(.dina(n12231), .dinb(n12206), .dout(n12232));
  jnot g12165(.din(n12232), .dout(n12233));
  jor  g12166(.dina(n5266), .dinb(n4343), .dout(n12234));
  jor  g12167(.dina(n4686), .dinb(n4346), .dout(n12235));
  jor  g12168(.dina(n5264), .dinb(n4348), .dout(n12236));
  jand g12169(.dina(n12236), .dinb(n12235), .dout(n12237));
  jor  g12170(.dina(n4526), .dinb(n3683), .dout(n12238));
  jand g12171(.dina(n12238), .dinb(n12237), .dout(n12239));
  jand g12172(.dina(n12239), .dinb(n12234), .dout(n12240));
  jxor g12173(.dina(n12240), .dinb(\a[29] ), .dout(n12241));
  jxor g12174(.dina(n12241), .dinb(n12233), .dout(n12242));
  jxor g12175(.dina(n12242), .dinb(n12197), .dout(n12243));
  jor  g12176(.dina(n5527), .dinb(n2303), .dout(n12244));
  jor  g12177(.dina(n5364), .dinb(n2306), .dout(n12245));
  jor  g12178(.dina(n5525), .dinb(n2309), .dout(n12246));
  jor  g12179(.dina(n5422), .dinb(n1805), .dout(n12247));
  jand g12180(.dina(n12247), .dinb(n12246), .dout(n12248));
  jand g12181(.dina(n12248), .dinb(n12245), .dout(n12249));
  jand g12182(.dina(n12249), .dinb(n12244), .dout(n12250));
  jxor g12183(.dina(n12250), .dinb(n77), .dout(n12251));
  jxor g12184(.dina(n12251), .dinb(n12243), .dout(n12252));
  jxor g12185(.dina(n12252), .dinb(n12192), .dout(n12253));
  jnot g12186(.din(n12253), .dout(n12254));
  jor  g12187(.dina(n6999), .dinb(n807), .dout(n12255));
  jor  g12188(.dina(n6390), .dinb(n1613), .dout(n12256));
  jor  g12189(.dina(n6297), .dinb(n1621), .dout(n12257));
  jand g12190(.dina(n12257), .dinb(n12256), .dout(n12258));
  jor  g12191(.dina(n6205), .dinb(n1617), .dout(n12259));
  jand g12192(.dina(n12259), .dinb(n12258), .dout(n12260));
  jand g12193(.dina(n12260), .dinb(n12255), .dout(n12261));
  jxor g12194(.dina(n12261), .dinb(\a[23] ), .dout(n12262));
  jxor g12195(.dina(n12262), .dinb(n12254), .dout(n12263));
  jxor g12196(.dina(n12263), .dinb(n12187), .dout(n12264));
  jnot g12197(.din(n12264), .dout(n12265));
  jor  g12198(.dina(n7682), .dinb(n1820), .dout(n12266));
  jor  g12199(.dina(n7301), .dinb(n2181), .dout(n12267));
  jor  g12200(.dina(n7680), .dinb(n2189), .dout(n12268));
  jand g12201(.dina(n12268), .dinb(n12267), .dout(n12269));
  jor  g12202(.dina(n6489), .dinb(n2186), .dout(n12270));
  jand g12203(.dina(n12270), .dinb(n12269), .dout(n12271));
  jand g12204(.dina(n12271), .dinb(n12266), .dout(n12272));
  jxor g12205(.dina(n12272), .dinb(\a[20] ), .dout(n12273));
  jxor g12206(.dina(n12273), .dinb(n12265), .dout(n12274));
  jxor g12207(.dina(n12274), .dinb(n12184), .dout(n12275));
  jxor g12208(.dina(n12275), .dinb(n12175), .dout(n12276));
  jnot g12209(.din(n12276), .dout(n12277));
  jand g12210(.dina(n11791), .dinb(n11661), .dout(n12278));
  jnot g12211(.din(n12278), .dout(n12279));
  jor  g12212(.dina(n11797), .dinb(n11793), .dout(n12280));
  jand g12213(.dina(n12280), .dinb(n12279), .dout(n12281));
  jxor g12214(.dina(n12281), .dinb(n12277), .dout(n12282));
  jxor g12215(.dina(n12282), .dinb(n11798), .dout(n12283));
  jxor g12216(.dina(n12283), .dinb(n12170), .dout(n12284));
  jand g12217(.dina(n12284), .dinb(n4022), .dout(n12285));
  jand g12218(.dina(n12282), .dinb(n4220), .dout(n12286));
  jand g12219(.dina(n11798), .dinb(n4027), .dout(n12287));
  jand g12220(.dina(n11646), .dinb(n3870), .dout(n12288));
  jor  g12221(.dina(n12288), .dinb(n12287), .dout(n12289));
  jor  g12222(.dina(n12289), .dinb(n12286), .dout(n12290));
  jor  g12223(.dina(n12290), .dinb(n12285), .dout(n12291));
  jxor g12224(.dina(n12291), .dinb(n4050), .dout(n12292));
  jxor g12225(.dina(n12292), .dinb(n12167), .dout(n12293));
  jxor g12226(.dina(n12293), .dinb(n12078), .dout(n12294));
  jand g12227(.dina(n12263), .dinb(n12187), .dout(n12295));
  jnot g12228(.din(n12295), .dout(n12296));
  jor  g12229(.dina(n12273), .dinb(n12265), .dout(n12297));
  jand g12230(.dina(n12297), .dinb(n12296), .dout(n12298));
  jnot g12231(.din(n12298), .dout(n12299));
  jor  g12232(.dina(n8002), .dinb(n1820), .dout(n12300));
  jor  g12233(.dina(n7301), .dinb(n2186), .dout(n12301));
  jor  g12234(.dina(n7999), .dinb(n2189), .dout(n12302));
  jor  g12235(.dina(n7680), .dinb(n2181), .dout(n12303));
  jand g12236(.dina(n12303), .dinb(n12302), .dout(n12304));
  jand g12237(.dina(n12304), .dinb(n12301), .dout(n12305));
  jand g12238(.dina(n12305), .dinb(n12300), .dout(n12306));
  jxor g12239(.dina(n12306), .dinb(n2196), .dout(n12307));
  jand g12240(.dina(n12307), .dinb(n12299), .dout(n12308));
  jand g12241(.dina(n12252), .dinb(n12192), .dout(n12309));
  jnot g12242(.din(n12309), .dout(n12310));
  jor  g12243(.dina(n12262), .dinb(n12254), .dout(n12311));
  jand g12244(.dina(n12311), .dinb(n12310), .dout(n12312));
  jnot g12245(.din(n12312), .dout(n12313));
  jand g12246(.dina(n12242), .dinb(n12197), .dout(n12314));
  jand g12247(.dina(n12251), .dinb(n12243), .dout(n12315));
  jor  g12248(.dina(n12315), .dinb(n12314), .dout(n12316));
  jand g12249(.dina(n12231), .dinb(n12206), .dout(n12317));
  jnot g12250(.din(n12317), .dout(n12318));
  jor  g12251(.dina(n12241), .dinb(n12233), .dout(n12319));
  jand g12252(.dina(n12319), .dinb(n12318), .dout(n12320));
  jnot g12253(.din(n12320), .dout(n12321));
  jand g12254(.dina(n12229), .dinb(n11737), .dout(n12322));
  jand g12255(.dina(n12230), .dinb(n12210), .dout(n12323));
  jor  g12256(.dina(n12323), .dinb(n12322), .dout(n12324));
  jand g12257(.dina(n7489), .dinb(n3318), .dout(n12325));
  jand g12258(.dina(n1236), .dinb(n827), .dout(n12326));
  jand g12259(.dina(n12326), .dinb(n12325), .dout(n12327));
  jand g12260(.dina(n12327), .dinb(n3026), .dout(n12328));
  jand g12261(.dina(n3739), .dinb(n454), .dout(n12329));
  jand g12262(.dina(n12329), .dinb(n2077), .dout(n12330));
  jand g12263(.dina(n12330), .dinb(n6325), .dout(n12331));
  jand g12264(.dina(n1219), .dinb(n1096), .dout(n12332));
  jand g12265(.dina(n1378), .dinb(n716), .dout(n12333));
  jand g12266(.dina(n12333), .dinb(n12332), .dout(n12334));
  jand g12267(.dina(n12334), .dinb(n349), .dout(n12335));
  jand g12268(.dina(n1522), .dinb(n325), .dout(n12336));
  jand g12269(.dina(n12336), .dinb(n12335), .dout(n12337));
  jand g12270(.dina(n12337), .dinb(n8343), .dout(n12338));
  jand g12271(.dina(n12338), .dinb(n12331), .dout(n12339));
  jand g12272(.dina(n12339), .dinb(n2567), .dout(n12340));
  jand g12273(.dina(n12340), .dinb(n12328), .dout(n12341));
  jand g12274(.dina(n5998), .dinb(n5472), .dout(n12342));
  jand g12275(.dina(n12342), .dinb(n12341), .dout(n12343));
  jand g12276(.dina(n12343), .dinb(n12229), .dout(n12344));
  jnot g12277(.din(n12344), .dout(n12345));
  jor  g12278(.dina(n12343), .dinb(n12229), .dout(n12346));
  jand g12279(.dina(n12346), .dinb(n2441), .dout(n12347));
  jand g12280(.dina(n12347), .dinb(n12345), .dout(n12348));
  jnot g12281(.din(n12348), .dout(n12349));
  jand g12282(.dina(n12349), .dinb(n2441), .dout(n12350));
  jand g12283(.dina(n12349), .dinb(n12346), .dout(n12351));
  jand g12284(.dina(n12351), .dinb(n12345), .dout(n12352));
  jor  g12285(.dina(n12352), .dinb(n12350), .dout(n12353));
  jnot g12286(.din(n12353), .dout(n12354));
  jor  g12287(.dina(n7061), .dinb(n4714), .dout(n12355));
  jand g12288(.dina(n6050), .dinb(n4600), .dout(n12356));
  jand g12289(.dina(n5084), .dinb(n4527), .dout(n12357));
  jor  g12290(.dina(n12357), .dinb(n12356), .dout(n12358));
  jand g12291(.dina(n5082), .dinb(n4597), .dout(n12359));
  jor  g12292(.dina(n12359), .dinb(n12358), .dout(n12360));
  jnot g12293(.din(n12360), .dout(n12361));
  jand g12294(.dina(n12361), .dinb(n12355), .dout(n12362));
  jxor g12295(.dina(n12362), .dinb(n12354), .dout(n12363));
  jxor g12296(.dina(n12363), .dinb(n12324), .dout(n12364));
  jxor g12297(.dina(n12364), .dinb(n12321), .dout(n12365));
  jnot g12298(.din(n12365), .dout(n12366));
  jor  g12299(.dina(n5560), .dinb(n4343), .dout(n12367));
  jor  g12300(.dina(n5264), .dinb(n4346), .dout(n12368));
  jor  g12301(.dina(n5422), .dinb(n4348), .dout(n12369));
  jand g12302(.dina(n12369), .dinb(n12368), .dout(n12370));
  jor  g12303(.dina(n4686), .dinb(n3683), .dout(n12371));
  jand g12304(.dina(n12371), .dinb(n12370), .dout(n12372));
  jand g12305(.dina(n12372), .dinb(n12367), .dout(n12373));
  jxor g12306(.dina(n12373), .dinb(\a[29] ), .dout(n12374));
  jxor g12307(.dina(n12374), .dinb(n12366), .dout(n12375));
  jor  g12308(.dina(n6207), .dinb(n2303), .dout(n12376));
  jor  g12309(.dina(n5364), .dinb(n1805), .dout(n12377));
  jor  g12310(.dina(n6205), .dinb(n2309), .dout(n12378));
  jor  g12311(.dina(n5525), .dinb(n2306), .dout(n12379));
  jand g12312(.dina(n12379), .dinb(n12378), .dout(n12380));
  jand g12313(.dina(n12380), .dinb(n12377), .dout(n12381));
  jand g12314(.dina(n12381), .dinb(n12376), .dout(n12382));
  jxor g12315(.dina(n12382), .dinb(n77), .dout(n12383));
  jxor g12316(.dina(n12383), .dinb(n12375), .dout(n12384));
  jxor g12317(.dina(n12384), .dinb(n12316), .dout(n12385));
  jnot g12318(.din(n12385), .dout(n12386));
  jor  g12319(.dina(n6491), .dinb(n807), .dout(n12387));
  jor  g12320(.dina(n6297), .dinb(n1613), .dout(n12388));
  jor  g12321(.dina(n6489), .dinb(n1621), .dout(n12389));
  jand g12322(.dina(n12389), .dinb(n12388), .dout(n12390));
  jor  g12323(.dina(n6390), .dinb(n1617), .dout(n12391));
  jand g12324(.dina(n12391), .dinb(n12390), .dout(n12392));
  jand g12325(.dina(n12392), .dinb(n12387), .dout(n12393));
  jxor g12326(.dina(n12393), .dinb(\a[23] ), .dout(n12394));
  jxor g12327(.dina(n12394), .dinb(n12386), .dout(n12395));
  jxor g12328(.dina(n12395), .dinb(n12313), .dout(n12396));
  jxor g12329(.dina(n12307), .dinb(n12299), .dout(n12397));
  jand g12330(.dina(n12397), .dinb(n12396), .dout(n12398));
  jor  g12331(.dina(n12398), .dinb(n12308), .dout(n12399));
  jor  g12332(.dina(n12394), .dinb(n12386), .dout(n12400));
  jand g12333(.dina(n12395), .dinb(n12313), .dout(n12401));
  jnot g12334(.din(n12401), .dout(n12402));
  jand g12335(.dina(n12402), .dinb(n12400), .dout(n12403));
  jnot g12336(.din(n12403), .dout(n12404));
  jand g12337(.dina(n12383), .dinb(n12375), .dout(n12405));
  jand g12338(.dina(n12384), .dinb(n12316), .dout(n12406));
  jor  g12339(.dina(n12406), .dinb(n12405), .dout(n12407));
  jand g12340(.dina(n12364), .dinb(n12321), .dout(n12408));
  jnot g12341(.din(n12408), .dout(n12409));
  jor  g12342(.dina(n12374), .dinb(n12366), .dout(n12410));
  jand g12343(.dina(n12410), .dinb(n12409), .dout(n12411));
  jnot g12344(.din(n12411), .dout(n12412));
  jor  g12345(.dina(n12362), .dinb(n12354), .dout(n12413));
  jand g12346(.dina(n12363), .dinb(n12324), .dout(n12414));
  jnot g12347(.din(n12414), .dout(n12415));
  jand g12348(.dina(n12415), .dinb(n12413), .dout(n12416));
  jnot g12349(.din(n12416), .dout(n12417));
  jor  g12350(.dina(n7061), .dinb(n4688), .dout(n12418));
  jand g12351(.dina(n6050), .dinb(n4597), .dout(n12419));
  jand g12352(.dina(n5084), .dinb(n5163), .dout(n12420));
  jor  g12353(.dina(n12420), .dinb(n12419), .dout(n12421));
  jand g12354(.dina(n5082), .dinb(n4527), .dout(n12422));
  jor  g12355(.dina(n12422), .dinb(n12421), .dout(n12423));
  jnot g12356(.din(n12423), .dout(n12424));
  jand g12357(.dina(n12424), .dinb(n12418), .dout(n12425));
  jnot g12358(.din(n12425), .dout(n12426));
  jand g12359(.dina(n6254), .dinb(n270), .dout(n12427));
  jand g12360(.dina(n1207), .dinb(n1380), .dout(n12428));
  jand g12361(.dina(n12428), .dinb(n2343), .dout(n12429));
  jand g12362(.dina(n12429), .dinb(n12427), .dout(n12430));
  jand g12363(.dina(n5339), .dinb(n700), .dout(n12431));
  jand g12364(.dina(n1451), .dinb(n716), .dout(n12432));
  jand g12365(.dina(n12432), .dinb(n1865), .dout(n12433));
  jand g12366(.dina(n12433), .dinb(n12431), .dout(n12434));
  jand g12367(.dina(n3758), .dinb(n714), .dout(n12435));
  jand g12368(.dina(n3066), .dinb(n2526), .dout(n12436));
  jand g12369(.dina(n12436), .dinb(n12435), .dout(n12437));
  jand g12370(.dina(n12437), .dinb(n12434), .dout(n12438));
  jnot g12371(.din(n608), .dout(n12439));
  jand g12372(.dina(n2675), .dinb(n12439), .dout(n12440));
  jand g12373(.dina(n12440), .dinb(n11193), .dout(n12441));
  jand g12374(.dina(n12441), .dinb(n12438), .dout(n12442));
  jand g12375(.dina(n12442), .dinb(n12430), .dout(n12443));
  jand g12376(.dina(n4541), .dinb(n1326), .dout(n12444));
  jand g12377(.dina(n6433), .dinb(n981), .dout(n12445));
  jand g12378(.dina(n2508), .dinb(n1867), .dout(n12446));
  jand g12379(.dina(n12446), .dinb(n12445), .dout(n12447));
  jand g12380(.dina(n12447), .dinb(n12444), .dout(n12448));
  jand g12381(.dina(n12448), .dinb(n3966), .dout(n12449));
  jand g12382(.dina(n12449), .dinb(n3375), .dout(n12450));
  jand g12383(.dina(n12450), .dinb(n12443), .dout(n12451));
  jand g12384(.dina(n1832), .dinb(n1169), .dout(n12452));
  jand g12385(.dina(n5253), .dinb(n4670), .dout(n12453));
  jand g12386(.dina(n12453), .dinb(n12452), .dout(n12454));
  jand g12387(.dina(n440), .dinb(n92), .dout(n12455));
  jand g12388(.dina(n12455), .dinb(n917), .dout(n12456));
  jand g12389(.dina(n12456), .dinb(n558), .dout(n12457));
  jand g12390(.dina(n12457), .dinb(n12454), .dout(n12458));
  jand g12391(.dina(n12458), .dinb(n2712), .dout(n12459));
  jand g12392(.dina(n672), .dinb(n1432), .dout(n12460));
  jand g12393(.dina(n11721), .dinb(n1846), .dout(n12461));
  jand g12394(.dina(n12461), .dinb(n1088), .dout(n12462));
  jand g12395(.dina(n12462), .dinb(n12460), .dout(n12463));
  jand g12396(.dina(n12463), .dinb(n10724), .dout(n12464));
  jand g12397(.dina(n12464), .dinb(n12459), .dout(n12465));
  jand g12398(.dina(n1968), .dinb(n1328), .dout(n12466));
  jand g12399(.dina(n4675), .dinb(n3328), .dout(n12467));
  jand g12400(.dina(n12467), .dinb(n7230), .dout(n12468));
  jand g12401(.dina(n12468), .dinb(n12466), .dout(n12469));
  jand g12402(.dina(n12469), .dinb(n2132), .dout(n12470));
  jand g12403(.dina(n12470), .dinb(n881), .dout(n12471));
  jand g12404(.dina(n12471), .dinb(n12465), .dout(n12472));
  jand g12405(.dina(n12472), .dinb(n12451), .dout(n12473));
  jnot g12406(.din(n12473), .dout(n12474));
  jxor g12407(.dina(n12474), .dinb(n12351), .dout(n12475));
  jxor g12408(.dina(n12475), .dinb(n12426), .dout(n12476));
  jxor g12409(.dina(n12476), .dinb(n12417), .dout(n12477));
  jnot g12410(.din(n12477), .dout(n12478));
  jor  g12411(.dina(n5549), .dinb(n4343), .dout(n12479));
  jor  g12412(.dina(n5422), .dinb(n4346), .dout(n12480));
  jor  g12413(.dina(n5364), .dinb(n4348), .dout(n12481));
  jand g12414(.dina(n12481), .dinb(n12480), .dout(n12482));
  jor  g12415(.dina(n5264), .dinb(n3683), .dout(n12483));
  jand g12416(.dina(n12483), .dinb(n12482), .dout(n12484));
  jand g12417(.dina(n12484), .dinb(n12479), .dout(n12485));
  jxor g12418(.dina(n12485), .dinb(\a[29] ), .dout(n12486));
  jxor g12419(.dina(n12486), .dinb(n12478), .dout(n12487));
  jxor g12420(.dina(n12487), .dinb(n12412), .dout(n12488));
  jor  g12421(.dina(n6516), .dinb(n2303), .dout(n12489));
  jor  g12422(.dina(n6205), .dinb(n2306), .dout(n12490));
  jor  g12423(.dina(n5525), .dinb(n1805), .dout(n12491));
  jor  g12424(.dina(n6390), .dinb(n2309), .dout(n12492));
  jand g12425(.dina(n12492), .dinb(n12491), .dout(n12493));
  jand g12426(.dina(n12493), .dinb(n12490), .dout(n12494));
  jand g12427(.dina(n12494), .dinb(n12489), .dout(n12495));
  jxor g12428(.dina(n12495), .dinb(n77), .dout(n12496));
  jxor g12429(.dina(n12496), .dinb(n12488), .dout(n12497));
  jxor g12430(.dina(n12497), .dinb(n12407), .dout(n12498));
  jnot g12431(.din(n12498), .dout(n12499));
  jor  g12432(.dina(n7301), .dinb(n1621), .dout(n12500));
  jor  g12433(.dina(n7303), .dinb(n807), .dout(n12501));
  jor  g12434(.dina(n6297), .dinb(n1617), .dout(n12502));
  jor  g12435(.dina(n6489), .dinb(n1613), .dout(n12503));
  jand g12436(.dina(n12503), .dinb(n12502), .dout(n12504));
  jand g12437(.dina(n12504), .dinb(n12501), .dout(n12505));
  jand g12438(.dina(n12505), .dinb(n12500), .dout(n12506));
  jxor g12439(.dina(n12506), .dinb(\a[23] ), .dout(n12507));
  jxor g12440(.dina(n12507), .dinb(n12499), .dout(n12508));
  jxor g12441(.dina(n12508), .dinb(n12404), .dout(n12509));
  jnot g12442(.din(n12509), .dout(n12510));
  jor  g12443(.dina(n7999), .dinb(n2181), .dout(n12511));
  jor  g12444(.dina(n8260), .dinb(n1820), .dout(n12512));
  jor  g12445(.dina(n7680), .dinb(n2186), .dout(n12513));
  jand g12446(.dina(n12513), .dinb(n12512), .dout(n12514));
  jand g12447(.dina(n12514), .dinb(n12511), .dout(n12515));
  jxor g12448(.dina(n12515), .dinb(\a[20] ), .dout(n12516));
  jxor g12449(.dina(n12516), .dinb(n12510), .dout(n12517));
  jxor g12450(.dina(n12517), .dinb(n12399), .dout(n12518));
  jnot g12451(.din(n12518), .dout(n12519));
  jor  g12452(.dina(n12183), .dinb(n12179), .dout(n12520));
  jand g12453(.dina(n12274), .dinb(n12184), .dout(n12521));
  jnot g12454(.din(n12521), .dout(n12522));
  jand g12455(.dina(n12522), .dinb(n12520), .dout(n12523));
  jnot g12456(.din(n12523), .dout(n12524));
  jxor g12457(.dina(n12397), .dinb(n12396), .dout(n12525));
  jand g12458(.dina(n12525), .dinb(n12524), .dout(n12526));
  jnot g12459(.din(n12526), .dout(n12527));
  jand g12460(.dina(n12275), .dinb(n12175), .dout(n12528));
  jnot g12461(.din(n12528), .dout(n12529));
  jor  g12462(.dina(n12281), .dinb(n12277), .dout(n12530));
  jand g12463(.dina(n12530), .dinb(n12529), .dout(n12531));
  jxor g12464(.dina(n12525), .dinb(n12524), .dout(n12532));
  jnot g12465(.din(n12532), .dout(n12533));
  jor  g12466(.dina(n12533), .dinb(n12531), .dout(n12534));
  jand g12467(.dina(n12534), .dinb(n12527), .dout(n12535));
  jxor g12468(.dina(n12535), .dinb(n12519), .dout(n12536));
  jand g12469(.dina(n11305), .dinb(n11136), .dout(n12537));
  jor  g12470(.dina(n12537), .dinb(n11632), .dout(n12538));
  jand g12471(.dina(n12538), .dinb(n11630), .dout(n12539));
  jor  g12472(.dina(n12539), .dinb(n11628), .dout(n12540));
  jand g12473(.dina(n12540), .dinb(n11620), .dout(n12541));
  jor  g12474(.dina(n12541), .dinb(n11794), .dout(n12542));
  jand g12475(.dina(n12542), .dinb(n11792), .dout(n12543));
  jor  g12476(.dina(n12543), .dinb(n12278), .dout(n12544));
  jand g12477(.dina(n12544), .dinb(n12276), .dout(n12545));
  jor  g12478(.dina(n12545), .dinb(n12528), .dout(n12546));
  jxor g12479(.dina(n12532), .dinb(n12546), .dout(n12547));
  jand g12480(.dina(n12547), .dinb(n12536), .dout(n12548));
  jand g12481(.dina(n12547), .dinb(n12282), .dout(n12549));
  jand g12482(.dina(n12282), .dinb(n11798), .dout(n12550));
  jand g12483(.dina(n12283), .dinb(n12170), .dout(n12551));
  jor  g12484(.dina(n12551), .dinb(n12550), .dout(n12552));
  jxor g12485(.dina(n12547), .dinb(n12282), .dout(n12553));
  jand g12486(.dina(n12553), .dinb(n12552), .dout(n12554));
  jor  g12487(.dina(n12554), .dinb(n12549), .dout(n12555));
  jxor g12488(.dina(n12547), .dinb(n12536), .dout(n12556));
  jand g12489(.dina(n12556), .dinb(n12555), .dout(n12557));
  jor  g12490(.dina(n12557), .dinb(n12548), .dout(n12558));
  jand g12491(.dina(n12508), .dinb(n12404), .dout(n12559));
  jnot g12492(.din(n12559), .dout(n12560));
  jor  g12493(.dina(n12516), .dinb(n12510), .dout(n12561));
  jand g12494(.dina(n12561), .dinb(n12560), .dout(n12562));
  jnot g12495(.din(n12562), .dout(n12563));
  jand g12496(.dina(n12497), .dinb(n12407), .dout(n12564));
  jnot g12497(.din(n12564), .dout(n12565));
  jor  g12498(.dina(n12507), .dinb(n12499), .dout(n12566));
  jand g12499(.dina(n12566), .dinb(n12565), .dout(n12567));
  jor  g12500(.dina(n7999), .dinb(n2186), .dout(n12568));
  jor  g12501(.dina(n8295), .dinb(n1820), .dout(n12569));
  jand g12502(.dina(n12569), .dinb(n12568), .dout(n12570));
  jxor g12503(.dina(n12570), .dinb(\a[20] ), .dout(n12571));
  jxor g12504(.dina(n12571), .dinb(n12567), .dout(n12572));
  jand g12505(.dina(n12487), .dinb(n12412), .dout(n12573));
  jand g12506(.dina(n12496), .dinb(n12488), .dout(n12574));
  jor  g12507(.dina(n12574), .dinb(n12573), .dout(n12575));
  jnot g12508(.din(n12351), .dout(n12576));
  jand g12509(.dina(n12473), .dinb(n12576), .dout(n12577));
  jand g12510(.dina(n12475), .dinb(n12426), .dout(n12578));
  jor  g12511(.dina(n12578), .dinb(n12577), .dout(n12579));
  jor  g12512(.dina(n5266), .dinb(n7061), .dout(n12580));
  jand g12513(.dina(n6050), .dinb(n4527), .dout(n12581));
  jand g12514(.dina(n5426), .dinb(n5084), .dout(n12582));
  jor  g12515(.dina(n12582), .dinb(n12581), .dout(n12583));
  jand g12516(.dina(n5082), .dinb(n5163), .dout(n12584));
  jor  g12517(.dina(n12584), .dinb(n12583), .dout(n12585));
  jnot g12518(.din(n12585), .dout(n12586));
  jand g12519(.dina(n12586), .dinb(n12580), .dout(n12587));
  jnot g12520(.din(n12587), .dout(n12588));
  jand g12521(.dina(n950), .dinb(n1284), .dout(n12589));
  jand g12522(.dina(n8820), .dinb(n3978), .dout(n12590));
  jand g12523(.dina(n12590), .dinb(n3995), .dout(n12591));
  jand g12524(.dina(n12591), .dinb(n2476), .dout(n12592));
  jand g12525(.dina(n12592), .dinb(n12589), .dout(n12593));
  jand g12526(.dina(n12593), .dinb(n1907), .dout(n12594));
  jand g12527(.dina(n12594), .dinb(n10216), .dout(n12595));
  jand g12528(.dina(n3740), .dinb(n1345), .dout(n12596));
  jand g12529(.dina(n12596), .dinb(n1005), .dout(n12597));
  jand g12530(.dina(n1219), .dinb(n1334), .dout(n12598));
  jand g12531(.dina(n12598), .dinb(n5306), .dout(n12599));
  jand g12532(.dina(n6337), .dinb(n917), .dout(n12600));
  jand g12533(.dina(n5396), .dinb(n827), .dout(n12601));
  jand g12534(.dina(n12601), .dinb(n12600), .dout(n12602));
  jand g12535(.dina(n12602), .dinb(n12599), .dout(n12603));
  jand g12536(.dina(n12603), .dinb(n12597), .dout(n12604));
  jand g12537(.dina(n2367), .dinb(n465), .dout(n12605));
  jand g12538(.dina(n12605), .dinb(n1752), .dout(n12606));
  jand g12539(.dina(n12606), .dinb(n10136), .dout(n12607));
  jand g12540(.dina(n589), .dinb(n1430), .dout(n12608));
  jand g12541(.dina(n12608), .dinb(n2039), .dout(n12609));
  jand g12542(.dina(n1288), .dinb(n92), .dout(n12610));
  jand g12543(.dina(n12610), .dinb(n1346), .dout(n12611));
  jand g12544(.dina(n12611), .dinb(n650), .dout(n12612));
  jand g12545(.dina(n12612), .dinb(n12609), .dout(n12613));
  jand g12546(.dina(n12613), .dinb(n12607), .dout(n12614));
  jand g12547(.dina(n12614), .dinb(n10171), .dout(n12615));
  jand g12548(.dina(n12615), .dinb(n12604), .dout(n12616));
  jand g12549(.dina(n1167), .dinb(n1429), .dout(n12617));
  jand g12550(.dina(n12617), .dinb(n4576), .dout(n12618));
  jand g12551(.dina(n7490), .dinb(n5191), .dout(n12619));
  jand g12552(.dina(n12619), .dinb(n12618), .dout(n12620));
  jand g12553(.dina(n12620), .dinb(n12616), .dout(n12621));
  jand g12554(.dina(n12621), .dinb(n12595), .dout(n12622));
  jxor g12555(.dina(n12622), .dinb(n12474), .dout(n12623));
  jxor g12556(.dina(n12623), .dinb(n12588), .dout(n12624));
  jxor g12557(.dina(n12624), .dinb(n12579), .dout(n12625));
  jnot g12558(.din(n12625), .dout(n12626));
  jand g12559(.dina(n12476), .dinb(n12417), .dout(n12627));
  jnot g12560(.din(n12627), .dout(n12628));
  jor  g12561(.dina(n12486), .dinb(n12478), .dout(n12629));
  jand g12562(.dina(n12629), .dinb(n12628), .dout(n12630));
  jxor g12563(.dina(n12630), .dinb(n12626), .dout(n12631));
  jnot g12564(.din(n12631), .dout(n12632));
  jor  g12565(.dina(n5527), .dinb(n4343), .dout(n12633));
  jor  g12566(.dina(n5364), .dinb(n4346), .dout(n12634));
  jor  g12567(.dina(n5525), .dinb(n4348), .dout(n12635));
  jand g12568(.dina(n12635), .dinb(n12634), .dout(n12636));
  jor  g12569(.dina(n5422), .dinb(n3683), .dout(n12637));
  jand g12570(.dina(n12637), .dinb(n12636), .dout(n12638));
  jand g12571(.dina(n12638), .dinb(n12633), .dout(n12639));
  jxor g12572(.dina(n12639), .dinb(\a[29] ), .dout(n12640));
  jxor g12573(.dina(n12640), .dinb(n12632), .dout(n12641));
  jor  g12574(.dina(n6999), .dinb(n2303), .dout(n12642));
  jor  g12575(.dina(n6390), .dinb(n2306), .dout(n12643));
  jor  g12576(.dina(n6205), .dinb(n1805), .dout(n12644));
  jor  g12577(.dina(n6297), .dinb(n2309), .dout(n12645));
  jand g12578(.dina(n12645), .dinb(n12644), .dout(n12646));
  jand g12579(.dina(n12646), .dinb(n12643), .dout(n12647));
  jand g12580(.dina(n12647), .dinb(n12642), .dout(n12648));
  jxor g12581(.dina(n12648), .dinb(n77), .dout(n12649));
  jxor g12582(.dina(n12649), .dinb(n12641), .dout(n12650));
  jxor g12583(.dina(n12650), .dinb(n12575), .dout(n12651));
  jnot g12584(.din(n12651), .dout(n12652));
  jor  g12585(.dina(n7682), .dinb(n807), .dout(n12653));
  jor  g12586(.dina(n7301), .dinb(n1613), .dout(n12654));
  jor  g12587(.dina(n6489), .dinb(n1617), .dout(n12655));
  jand g12588(.dina(n12655), .dinb(n12654), .dout(n12656));
  jor  g12589(.dina(n7680), .dinb(n1621), .dout(n12657));
  jand g12590(.dina(n12657), .dinb(n12656), .dout(n12658));
  jand g12591(.dina(n12658), .dinb(n12653), .dout(n12659));
  jxor g12592(.dina(n12659), .dinb(\a[23] ), .dout(n12660));
  jxor g12593(.dina(n12660), .dinb(n12652), .dout(n12661));
  jxor g12594(.dina(n12661), .dinb(n12572), .dout(n12662));
  jxor g12595(.dina(n12662), .dinb(n12563), .dout(n12663));
  jnot g12596(.din(n12663), .dout(n12664));
  jand g12597(.dina(n12517), .dinb(n12399), .dout(n12665));
  jnot g12598(.din(n12665), .dout(n12666));
  jor  g12599(.dina(n12535), .dinb(n12519), .dout(n12667));
  jand g12600(.dina(n12667), .dinb(n12666), .dout(n12668));
  jxor g12601(.dina(n12668), .dinb(n12664), .dout(n12669));
  jxor g12602(.dina(n12669), .dinb(n12536), .dout(n12670));
  jxor g12603(.dina(n12670), .dinb(n12558), .dout(n12671));
  jand g12604(.dina(n12671), .dinb(n4691), .dout(n12672));
  jand g12605(.dina(n12669), .dinb(n4941), .dout(n12673));
  jand g12606(.dina(n12536), .dinb(n4696), .dout(n12674));
  jand g12607(.dina(n12547), .dinb(n4701), .dout(n12675));
  jor  g12608(.dina(n12675), .dinb(n12674), .dout(n12676));
  jor  g12609(.dina(n12676), .dinb(n12673), .dout(n12677));
  jor  g12610(.dina(n12677), .dinb(n12672), .dout(n12678));
  jxor g12611(.dina(n12678), .dinb(n4713), .dout(n12679));
  jor  g12612(.dina(n12679), .dinb(n12294), .dout(n12680));
  jnot g12613(.din(n12680), .dout(n12681));
  jxor g12614(.dina(n12076), .dinb(n12075), .dout(n12682));
  jnot g12615(.din(n12682), .dout(n12683));
  jxor g12616(.dina(n12556), .dinb(n12555), .dout(n12684));
  jand g12617(.dina(n12684), .dinb(n4691), .dout(n12685));
  jand g12618(.dina(n12536), .dinb(n4941), .dout(n12686));
  jand g12619(.dina(n12547), .dinb(n4696), .dout(n12687));
  jand g12620(.dina(n12282), .dinb(n4701), .dout(n12688));
  jor  g12621(.dina(n12688), .dinb(n12687), .dout(n12689));
  jor  g12622(.dina(n12689), .dinb(n12686), .dout(n12690));
  jor  g12623(.dina(n12690), .dinb(n12685), .dout(n12691));
  jxor g12624(.dina(n12691), .dinb(n4713), .dout(n12692));
  jor  g12625(.dina(n12692), .dinb(n12683), .dout(n12693));
  jxor g12626(.dina(n12073), .dinb(n12072), .dout(n12694));
  jnot g12627(.din(n12694), .dout(n12695));
  jxor g12628(.dina(n12553), .dinb(n12552), .dout(n12696));
  jand g12629(.dina(n12696), .dinb(n4691), .dout(n12697));
  jand g12630(.dina(n12547), .dinb(n4941), .dout(n12698));
  jand g12631(.dina(n12282), .dinb(n4696), .dout(n12699));
  jand g12632(.dina(n11798), .dinb(n4701), .dout(n12700));
  jor  g12633(.dina(n12700), .dinb(n12699), .dout(n12701));
  jor  g12634(.dina(n12701), .dinb(n12698), .dout(n12702));
  jor  g12635(.dina(n12702), .dinb(n12697), .dout(n12703));
  jxor g12636(.dina(n12703), .dinb(n4713), .dout(n12704));
  jor  g12637(.dina(n12704), .dinb(n12695), .dout(n12705));
  jxor g12638(.dina(n12069), .dinb(n12068), .dout(n12706));
  jand g12639(.dina(n12284), .dinb(n4691), .dout(n12707));
  jand g12640(.dina(n12282), .dinb(n4941), .dout(n12708));
  jand g12641(.dina(n11798), .dinb(n4696), .dout(n12709));
  jand g12642(.dina(n11646), .dinb(n4701), .dout(n12710));
  jor  g12643(.dina(n12710), .dinb(n12709), .dout(n12711));
  jor  g12644(.dina(n12711), .dinb(n12708), .dout(n12712));
  jor  g12645(.dina(n12712), .dinb(n12707), .dout(n12713));
  jxor g12646(.dina(n12713), .dinb(n4713), .dout(n12714));
  jor  g12647(.dina(n12714), .dinb(n12706), .dout(n12715));
  jxor g12648(.dina(n12066), .dinb(n12064), .dout(n12716));
  jnot g12649(.din(n12716), .dout(n12717));
  jand g12650(.dina(n11800), .dinb(n4691), .dout(n12718));
  jand g12651(.dina(n11646), .dinb(n4696), .dout(n12719));
  jand g12652(.dina(n11798), .dinb(n4941), .dout(n12720));
  jor  g12653(.dina(n12720), .dinb(n12719), .dout(n12721));
  jand g12654(.dina(n11647), .dinb(n4701), .dout(n12722));
  jor  g12655(.dina(n12722), .dinb(n12721), .dout(n12723));
  jor  g12656(.dina(n12723), .dinb(n12718), .dout(n12724));
  jxor g12657(.dina(n12724), .dinb(n4713), .dout(n12725));
  jor  g12658(.dina(n12725), .dinb(n12717), .dout(n12726));
  jxor g12659(.dina(n12062), .dinb(n12060), .dout(n12727));
  jnot g12660(.din(n12727), .dout(n12728));
  jand g12661(.dina(n11812), .dinb(n4691), .dout(n12729));
  jand g12662(.dina(n11646), .dinb(n4941), .dout(n12730));
  jand g12663(.dina(n11647), .dinb(n4696), .dout(n12731));
  jand g12664(.dina(n11306), .dinb(n4701), .dout(n12732));
  jor  g12665(.dina(n12732), .dinb(n12731), .dout(n12733));
  jor  g12666(.dina(n12733), .dinb(n12730), .dout(n12734));
  jor  g12667(.dina(n12734), .dinb(n12729), .dout(n12735));
  jxor g12668(.dina(n12735), .dinb(n4713), .dout(n12736));
  jor  g12669(.dina(n12736), .dinb(n12728), .dout(n12737));
  jxor g12670(.dina(n12058), .dinb(n12056), .dout(n12738));
  jnot g12671(.din(n12738), .dout(n12739));
  jand g12672(.dina(n11824), .dinb(n4691), .dout(n12740));
  jand g12673(.dina(n11306), .dinb(n4696), .dout(n12741));
  jand g12674(.dina(n11647), .dinb(n4941), .dout(n12742));
  jor  g12675(.dina(n12742), .dinb(n12741), .dout(n12743));
  jand g12676(.dina(n10836), .dinb(n4701), .dout(n12744));
  jor  g12677(.dina(n12744), .dinb(n12743), .dout(n12745));
  jor  g12678(.dina(n12745), .dinb(n12740), .dout(n12746));
  jxor g12679(.dina(n12746), .dinb(n4713), .dout(n12747));
  jor  g12680(.dina(n12747), .dinb(n12739), .dout(n12748));
  jxor g12681(.dina(n12054), .dinb(n12052), .dout(n12749));
  jnot g12682(.din(n12749), .dout(n12750));
  jand g12683(.dina(n11308), .dinb(n4691), .dout(n12751));
  jand g12684(.dina(n11306), .dinb(n4941), .dout(n12752));
  jand g12685(.dina(n10836), .dinb(n4696), .dout(n12753));
  jand g12686(.dina(n10640), .dinb(n4701), .dout(n12754));
  jor  g12687(.dina(n12754), .dinb(n12753), .dout(n12755));
  jor  g12688(.dina(n12755), .dinb(n12752), .dout(n12756));
  jor  g12689(.dina(n12756), .dinb(n12751), .dout(n12757));
  jxor g12690(.dina(n12757), .dinb(n4713), .dout(n12758));
  jor  g12691(.dina(n12758), .dinb(n12750), .dout(n12759));
  jxor g12692(.dina(n12050), .dinb(n12048), .dout(n12760));
  jnot g12693(.din(n12760), .dout(n12761));
  jand g12694(.dina(n10838), .dinb(n4691), .dout(n12762));
  jand g12695(.dina(n10836), .dinb(n4941), .dout(n12763));
  jand g12696(.dina(n10640), .dinb(n4696), .dout(n12764));
  jand g12697(.dina(n10647), .dinb(n4701), .dout(n12765));
  jor  g12698(.dina(n12765), .dinb(n12764), .dout(n12766));
  jor  g12699(.dina(n12766), .dinb(n12763), .dout(n12767));
  jor  g12700(.dina(n12767), .dinb(n12762), .dout(n12768));
  jxor g12701(.dina(n12768), .dinb(n4713), .dout(n12769));
  jor  g12702(.dina(n12769), .dinb(n12761), .dout(n12770));
  jxor g12703(.dina(n12045), .dinb(n12044), .dout(n12771));
  jnot g12704(.din(n12771), .dout(n12772));
  jand g12705(.dina(n10850), .dinb(n4691), .dout(n12773));
  jand g12706(.dina(n10640), .dinb(n4941), .dout(n12774));
  jand g12707(.dina(n10647), .dinb(n4696), .dout(n12775));
  jand g12708(.dina(n10305), .dinb(n4701), .dout(n12776));
  jor  g12709(.dina(n12776), .dinb(n12775), .dout(n12777));
  jor  g12710(.dina(n12777), .dinb(n12774), .dout(n12778));
  jor  g12711(.dina(n12778), .dinb(n12773), .dout(n12779));
  jxor g12712(.dina(n12779), .dinb(n4713), .dout(n12780));
  jor  g12713(.dina(n12780), .dinb(n12772), .dout(n12781));
  jxor g12714(.dina(n12040), .dinb(n12039), .dout(n12782));
  jnot g12715(.din(n12782), .dout(n12783));
  jand g12716(.dina(n10862), .dinb(n4691), .dout(n12784));
  jand g12717(.dina(n10647), .dinb(n4941), .dout(n12785));
  jand g12718(.dina(n10305), .dinb(n4696), .dout(n12786));
  jand g12719(.dina(n9872), .dinb(n4701), .dout(n12787));
  jor  g12720(.dina(n12787), .dinb(n12786), .dout(n12788));
  jor  g12721(.dina(n12788), .dinb(n12785), .dout(n12789));
  jor  g12722(.dina(n12789), .dinb(n12784), .dout(n12790));
  jxor g12723(.dina(n12790), .dinb(n4713), .dout(n12791));
  jor  g12724(.dina(n12791), .dinb(n12783), .dout(n12792));
  jxor g12725(.dina(n12035), .dinb(n12034), .dout(n12793));
  jnot g12726(.din(n12793), .dout(n12794));
  jand g12727(.dina(n10307), .dinb(n4691), .dout(n12795));
  jand g12728(.dina(n9872), .dinb(n4696), .dout(n12796));
  jand g12729(.dina(n10305), .dinb(n4941), .dout(n12797));
  jor  g12730(.dina(n12797), .dinb(n12796), .dout(n12798));
  jand g12731(.dina(n9655), .dinb(n4701), .dout(n12799));
  jor  g12732(.dina(n12799), .dinb(n12798), .dout(n12800));
  jor  g12733(.dina(n12800), .dinb(n12795), .dout(n12801));
  jxor g12734(.dina(n12801), .dinb(n4713), .dout(n12802));
  jor  g12735(.dina(n12802), .dinb(n12794), .dout(n12803));
  jxor g12736(.dina(n12030), .dinb(n12029), .dout(n12804));
  jnot g12737(.din(n12804), .dout(n12805));
  jand g12738(.dina(n9874), .dinb(n4691), .dout(n12806));
  jand g12739(.dina(n9872), .dinb(n4941), .dout(n12807));
  jand g12740(.dina(n9655), .dinb(n4696), .dout(n12808));
  jand g12741(.dina(n9656), .dinb(n4701), .dout(n12809));
  jor  g12742(.dina(n12809), .dinb(n12808), .dout(n12810));
  jor  g12743(.dina(n12810), .dinb(n12807), .dout(n12811));
  jor  g12744(.dina(n12811), .dinb(n12806), .dout(n12812));
  jxor g12745(.dina(n12812), .dinb(n4713), .dout(n12813));
  jor  g12746(.dina(n12813), .dinb(n12805), .dout(n12814));
  jxor g12747(.dina(n12025), .dinb(n12024), .dout(n12815));
  jnot g12748(.din(n12815), .dout(n12816));
  jand g12749(.dina(n9886), .dinb(n4691), .dout(n12817));
  jand g12750(.dina(n9655), .dinb(n4941), .dout(n12818));
  jand g12751(.dina(n9656), .dinb(n4696), .dout(n12819));
  jand g12752(.dina(n9250), .dinb(n4701), .dout(n12820));
  jor  g12753(.dina(n12820), .dinb(n12819), .dout(n12821));
  jor  g12754(.dina(n12821), .dinb(n12818), .dout(n12822));
  jor  g12755(.dina(n12822), .dinb(n12817), .dout(n12823));
  jxor g12756(.dina(n12823), .dinb(n4713), .dout(n12824));
  jor  g12757(.dina(n12824), .dinb(n12816), .dout(n12825));
  jxor g12758(.dina(n12020), .dinb(n12019), .dout(n12826));
  jnot g12759(.din(n12826), .dout(n12827));
  jand g12760(.dina(n9898), .dinb(n4691), .dout(n12828));
  jand g12761(.dina(n9656), .dinb(n4941), .dout(n12829));
  jand g12762(.dina(n9250), .dinb(n4696), .dout(n12830));
  jand g12763(.dina(n8936), .dinb(n4701), .dout(n12831));
  jor  g12764(.dina(n12831), .dinb(n12830), .dout(n12832));
  jor  g12765(.dina(n12832), .dinb(n12829), .dout(n12833));
  jor  g12766(.dina(n12833), .dinb(n12828), .dout(n12834));
  jxor g12767(.dina(n12834), .dinb(n4713), .dout(n12835));
  jor  g12768(.dina(n12835), .dinb(n12827), .dout(n12836));
  jxor g12769(.dina(n12017), .dinb(n12016), .dout(n12837));
  jnot g12770(.din(n12837), .dout(n12838));
  jand g12771(.dina(n9252), .dinb(n4691), .dout(n12839));
  jand g12772(.dina(n8936), .dinb(n4696), .dout(n12840));
  jand g12773(.dina(n9250), .dinb(n4941), .dout(n12841));
  jor  g12774(.dina(n12841), .dinb(n12840), .dout(n12842));
  jand g12775(.dina(n8723), .dinb(n4701), .dout(n12843));
  jor  g12776(.dina(n12843), .dinb(n12842), .dout(n12844));
  jor  g12777(.dina(n12844), .dinb(n12839), .dout(n12845));
  jxor g12778(.dina(n12845), .dinb(n4713), .dout(n12846));
  jor  g12779(.dina(n12846), .dinb(n12838), .dout(n12847));
  jxor g12780(.dina(n12012), .dinb(n12011), .dout(n12848));
  jnot g12781(.din(n12848), .dout(n12849));
  jand g12782(.dina(n8938), .dinb(n4691), .dout(n12850));
  jand g12783(.dina(n8723), .dinb(n4696), .dout(n12851));
  jand g12784(.dina(n8936), .dinb(n4941), .dout(n12852));
  jor  g12785(.dina(n12852), .dinb(n12851), .dout(n12853));
  jand g12786(.dina(n8740), .dinb(n4701), .dout(n12854));
  jor  g12787(.dina(n12854), .dinb(n12853), .dout(n12855));
  jor  g12788(.dina(n12855), .dinb(n12850), .dout(n12856));
  jxor g12789(.dina(n12856), .dinb(n4713), .dout(n12857));
  jor  g12790(.dina(n12857), .dinb(n12849), .dout(n12858));
  jxor g12791(.dina(n12008), .dinb(n12000), .dout(n12859));
  jnot g12792(.din(n12859), .dout(n12860));
  jand g12793(.dina(n8950), .dinb(n4691), .dout(n12861));
  jand g12794(.dina(n8723), .dinb(n4941), .dout(n12862));
  jand g12795(.dina(n8740), .dinb(n4696), .dout(n12863));
  jand g12796(.dina(n8268), .dinb(n4701), .dout(n12864));
  jor  g12797(.dina(n12864), .dinb(n12863), .dout(n12865));
  jor  g12798(.dina(n12865), .dinb(n12862), .dout(n12866));
  jor  g12799(.dina(n12866), .dinb(n12861), .dout(n12867));
  jxor g12800(.dina(n12867), .dinb(n4713), .dout(n12868));
  jor  g12801(.dina(n12868), .dinb(n12860), .dout(n12869));
  jand g12802(.dina(n8962), .dinb(n4691), .dout(n12870));
  jand g12803(.dina(n8740), .dinb(n4941), .dout(n12871));
  jand g12804(.dina(n8268), .dinb(n4696), .dout(n12872));
  jand g12805(.dina(n8022), .dinb(n4701), .dout(n12873));
  jor  g12806(.dina(n12873), .dinb(n12872), .dout(n12874));
  jor  g12807(.dina(n12874), .dinb(n12871), .dout(n12875));
  jor  g12808(.dina(n12875), .dinb(n12870), .dout(n12876));
  jxor g12809(.dina(n12876), .dinb(n4713), .dout(n12877));
  jnot g12810(.din(n12877), .dout(n12878));
  jor  g12811(.dina(n11987), .dinb(n4050), .dout(n12879));
  jxor g12812(.dina(n12879), .dinb(n11995), .dout(n12880));
  jand g12813(.dina(n12880), .dinb(n12878), .dout(n12881));
  jand g12814(.dina(n11984), .dinb(\a[11] ), .dout(n12882));
  jxor g12815(.dina(n12882), .dinb(n11982), .dout(n12883));
  jnot g12816(.din(n12883), .dout(n12884));
  jand g12817(.dina(n8270), .dinb(n4691), .dout(n12885));
  jand g12818(.dina(n8022), .dinb(n4696), .dout(n12886));
  jand g12819(.dina(n8268), .dinb(n4941), .dout(n12887));
  jor  g12820(.dina(n12887), .dinb(n12886), .dout(n12888));
  jand g12821(.dina(n7692), .dinb(n4701), .dout(n12889));
  jor  g12822(.dina(n12889), .dinb(n12888), .dout(n12890));
  jor  g12823(.dina(n12890), .dinb(n12885), .dout(n12891));
  jxor g12824(.dina(n12891), .dinb(n4713), .dout(n12892));
  jor  g12825(.dina(n12892), .dinb(n12884), .dout(n12893));
  jand g12826(.dina(n7315), .dinb(n4691), .dout(n12894));
  jand g12827(.dina(n7019), .dinb(n4696), .dout(n12895));
  jand g12828(.dina(n7313), .dinb(n4941), .dout(n12896));
  jor  g12829(.dina(n12896), .dinb(n12895), .dout(n12897));
  jor  g12830(.dina(n12897), .dinb(n12894), .dout(n12898));
  jnot g12831(.din(n12898), .dout(n12899));
  jand g12832(.dina(n7019), .dinb(n4689), .dout(n12900));
  jnot g12833(.din(n12900), .dout(n12901));
  jand g12834(.dina(n12901), .dinb(\a[8] ), .dout(n12902));
  jand g12835(.dina(n12902), .dinb(n12899), .dout(n12903));
  jand g12836(.dina(n7693), .dinb(n4691), .dout(n12904));
  jand g12837(.dina(n7313), .dinb(n4696), .dout(n12905));
  jor  g12838(.dina(n12905), .dinb(n12904), .dout(n12906));
  jand g12839(.dina(n7692), .dinb(n4941), .dout(n12907));
  jand g12840(.dina(n7019), .dinb(n4701), .dout(n12908));
  jor  g12841(.dina(n12908), .dinb(n12907), .dout(n12909));
  jor  g12842(.dina(n12909), .dinb(n12906), .dout(n12910));
  jnot g12843(.din(n12910), .dout(n12911));
  jand g12844(.dina(n12911), .dinb(n12903), .dout(n12912));
  jand g12845(.dina(n12912), .dinb(n11984), .dout(n12913));
  jnot g12846(.din(n12913), .dout(n12914));
  jxor g12847(.dina(n12912), .dinb(n11984), .dout(n12915));
  jnot g12848(.din(n12915), .dout(n12916));
  jand g12849(.dina(n8029), .dinb(n4691), .dout(n12917));
  jand g12850(.dina(n8022), .dinb(n4941), .dout(n12918));
  jand g12851(.dina(n7313), .dinb(n4701), .dout(n12919));
  jand g12852(.dina(n7692), .dinb(n4696), .dout(n12920));
  jor  g12853(.dina(n12920), .dinb(n12919), .dout(n12921));
  jor  g12854(.dina(n12921), .dinb(n12918), .dout(n12922));
  jor  g12855(.dina(n12922), .dinb(n12917), .dout(n12923));
  jxor g12856(.dina(n12923), .dinb(n4713), .dout(n12924));
  jor  g12857(.dina(n12924), .dinb(n12916), .dout(n12925));
  jand g12858(.dina(n12925), .dinb(n12914), .dout(n12926));
  jnot g12859(.din(n12926), .dout(n12927));
  jxor g12860(.dina(n12892), .dinb(n12884), .dout(n12928));
  jand g12861(.dina(n12928), .dinb(n12927), .dout(n12929));
  jnot g12862(.din(n12929), .dout(n12930));
  jand g12863(.dina(n12930), .dinb(n12893), .dout(n12931));
  jnot g12864(.din(n12931), .dout(n12932));
  jxor g12865(.dina(n12880), .dinb(n12878), .dout(n12933));
  jand g12866(.dina(n12933), .dinb(n12932), .dout(n12934));
  jor  g12867(.dina(n12934), .dinb(n12881), .dout(n12935));
  jxor g12868(.dina(n12868), .dinb(n12860), .dout(n12936));
  jand g12869(.dina(n12936), .dinb(n12935), .dout(n12937));
  jnot g12870(.din(n12937), .dout(n12938));
  jand g12871(.dina(n12938), .dinb(n12869), .dout(n12939));
  jnot g12872(.din(n12939), .dout(n12940));
  jxor g12873(.dina(n12857), .dinb(n12849), .dout(n12941));
  jand g12874(.dina(n12941), .dinb(n12940), .dout(n12942));
  jnot g12875(.din(n12942), .dout(n12943));
  jand g12876(.dina(n12943), .dinb(n12858), .dout(n12944));
  jnot g12877(.din(n12944), .dout(n12945));
  jxor g12878(.dina(n12846), .dinb(n12838), .dout(n12946));
  jand g12879(.dina(n12946), .dinb(n12945), .dout(n12947));
  jnot g12880(.din(n12947), .dout(n12948));
  jand g12881(.dina(n12948), .dinb(n12847), .dout(n12949));
  jnot g12882(.din(n12949), .dout(n12950));
  jxor g12883(.dina(n12835), .dinb(n12827), .dout(n12951));
  jand g12884(.dina(n12951), .dinb(n12950), .dout(n12952));
  jnot g12885(.din(n12952), .dout(n12953));
  jand g12886(.dina(n12953), .dinb(n12836), .dout(n12954));
  jxor g12887(.dina(n12824), .dinb(n12816), .dout(n12955));
  jnot g12888(.din(n12955), .dout(n12956));
  jor  g12889(.dina(n12956), .dinb(n12954), .dout(n12957));
  jand g12890(.dina(n12957), .dinb(n12825), .dout(n12958));
  jxor g12891(.dina(n12813), .dinb(n12805), .dout(n12959));
  jnot g12892(.din(n12959), .dout(n12960));
  jor  g12893(.dina(n12960), .dinb(n12958), .dout(n12961));
  jand g12894(.dina(n12961), .dinb(n12814), .dout(n12962));
  jxor g12895(.dina(n12802), .dinb(n12794), .dout(n12963));
  jnot g12896(.din(n12963), .dout(n12964));
  jor  g12897(.dina(n12964), .dinb(n12962), .dout(n12965));
  jand g12898(.dina(n12965), .dinb(n12803), .dout(n12966));
  jxor g12899(.dina(n12791), .dinb(n12783), .dout(n12967));
  jnot g12900(.din(n12967), .dout(n12968));
  jor  g12901(.dina(n12968), .dinb(n12966), .dout(n12969));
  jand g12902(.dina(n12969), .dinb(n12792), .dout(n12970));
  jxor g12903(.dina(n12780), .dinb(n12772), .dout(n12971));
  jnot g12904(.din(n12971), .dout(n12972));
  jor  g12905(.dina(n12972), .dinb(n12970), .dout(n12973));
  jand g12906(.dina(n12973), .dinb(n12781), .dout(n12974));
  jxor g12907(.dina(n12769), .dinb(n12760), .dout(n12975));
  jor  g12908(.dina(n12975), .dinb(n12974), .dout(n12976));
  jand g12909(.dina(n12976), .dinb(n12770), .dout(n12977));
  jxor g12910(.dina(n12758), .dinb(n12749), .dout(n12978));
  jor  g12911(.dina(n12978), .dinb(n12977), .dout(n12979));
  jand g12912(.dina(n12979), .dinb(n12759), .dout(n12980));
  jxor g12913(.dina(n12747), .dinb(n12738), .dout(n12981));
  jor  g12914(.dina(n12981), .dinb(n12980), .dout(n12982));
  jand g12915(.dina(n12982), .dinb(n12748), .dout(n12983));
  jxor g12916(.dina(n12736), .dinb(n12727), .dout(n12984));
  jor  g12917(.dina(n12984), .dinb(n12983), .dout(n12985));
  jand g12918(.dina(n12985), .dinb(n12737), .dout(n12986));
  jxor g12919(.dina(n12725), .dinb(n12716), .dout(n12987));
  jor  g12920(.dina(n12987), .dinb(n12986), .dout(n12988));
  jand g12921(.dina(n12988), .dinb(n12726), .dout(n12989));
  jxor g12922(.dina(n12714), .dinb(n12706), .dout(n12990));
  jnot g12923(.din(n12990), .dout(n12991));
  jor  g12924(.dina(n12991), .dinb(n12989), .dout(n12992));
  jand g12925(.dina(n12992), .dinb(n12715), .dout(n12993));
  jxor g12926(.dina(n12704), .dinb(n12695), .dout(n12994));
  jnot g12927(.din(n12994), .dout(n12995));
  jor  g12928(.dina(n12995), .dinb(n12993), .dout(n12996));
  jand g12929(.dina(n12996), .dinb(n12705), .dout(n12997));
  jxor g12930(.dina(n12692), .dinb(n12683), .dout(n12998));
  jnot g12931(.din(n12998), .dout(n12999));
  jor  g12932(.dina(n12999), .dinb(n12997), .dout(n13000));
  jand g12933(.dina(n13000), .dinb(n12693), .dout(n13001));
  jnot g12934(.din(n13001), .dout(n13002));
  jxor g12935(.dina(n12679), .dinb(n12294), .dout(n13003));
  jand g12936(.dina(n13003), .dinb(n13002), .dout(n13004));
  jor  g12937(.dina(n13004), .dinb(n12681), .dout(n13005));
  jor  g12938(.dina(n12292), .dinb(n12167), .dout(n13006));
  jnot g12939(.din(n12293), .dout(n13007));
  jor  g12940(.dina(n13007), .dinb(n12078), .dout(n13008));
  jand g12941(.dina(n13008), .dinb(n13006), .dout(n13009));
  jor  g12942(.dina(n12165), .dinb(n12157), .dout(n13010));
  jnot g12943(.din(n13010), .dout(n13011));
  jnot g12944(.din(n12081), .dout(n13012));
  jand g12945(.dina(n12166), .dinb(n13012), .dout(n13013));
  jor  g12946(.dina(n13013), .dinb(n13011), .dout(n13014));
  jor  g12947(.dina(n12154), .dinb(n12146), .dout(n13015));
  jand g12948(.dina(n12155), .dinb(n12086), .dout(n13016));
  jnot g12949(.din(n13016), .dout(n13017));
  jand g12950(.dina(n13017), .dinb(n13015), .dout(n13018));
  jnot g12951(.din(n13018), .dout(n13019));
  jand g12952(.dina(n12143), .dinb(n12135), .dout(n13020));
  jand g12953(.dina(n12144), .dinb(n12091), .dout(n13021));
  jor  g12954(.dina(n13021), .dinb(n13020), .dout(n13022));
  jor  g12955(.dina(n12133), .dinb(n12125), .dout(n13023));
  jand g12956(.dina(n12134), .dinb(n12096), .dout(n13024));
  jnot g12957(.din(n13024), .dout(n13025));
  jand g12958(.dina(n13025), .dinb(n13023), .dout(n13026));
  jnot g12959(.din(n13026), .dout(n13027));
  jand g12960(.dina(n12122), .dinb(n12114), .dout(n13028));
  jand g12961(.dina(n12123), .dinb(n12101), .dout(n13029));
  jor  g12962(.dina(n13029), .dinb(n13028), .dout(n13030));
  jand g12963(.dina(n7019), .dinb(n4338), .dout(n13031));
  jor  g12964(.dina(n12112), .dinb(n12108), .dout(n13032));
  jnot g12965(.din(n13032), .dout(n13033));
  jxor g12966(.dina(n13033), .dinb(n13031), .dout(n13034));
  jnot g12967(.din(n13034), .dout(n13035));
  jand g12968(.dina(n8029), .dinb(n2936), .dout(n13036));
  jand g12969(.dina(n7692), .dinb(n2940), .dout(n13037));
  jand g12970(.dina(n8022), .dinb(n2943), .dout(n13038));
  jor  g12971(.dina(n13038), .dinb(n13037), .dout(n13039));
  jand g12972(.dina(n7313), .dinb(n3684), .dout(n13040));
  jor  g12973(.dina(n13040), .dinb(n13039), .dout(n13041));
  jor  g12974(.dina(n13041), .dinb(n13036), .dout(n13042));
  jxor g12975(.dina(n13042), .dinb(n93), .dout(n13043));
  jxor g12976(.dina(n13043), .dinb(n13035), .dout(n13044));
  jand g12977(.dina(n8950), .dinb(n71), .dout(n13045));
  jand g12978(.dina(n8723), .dinb(n796), .dout(n13046));
  jand g12979(.dina(n8268), .dinb(n1806), .dout(n13047));
  jand g12980(.dina(n8740), .dinb(n731), .dout(n13048));
  jor  g12981(.dina(n13048), .dinb(n13047), .dout(n13049));
  jor  g12982(.dina(n13049), .dinb(n13046), .dout(n13050));
  jor  g12983(.dina(n13050), .dinb(n13045), .dout(n13051));
  jxor g12984(.dina(n13051), .dinb(\a[26] ), .dout(n13052));
  jxor g12985(.dina(n13052), .dinb(n13044), .dout(n13053));
  jxor g12986(.dina(n13053), .dinb(n13030), .dout(n13054));
  jnot g12987(.din(n13054), .dout(n13055));
  jand g12988(.dina(n9898), .dinb(n806), .dout(n13056));
  jand g12989(.dina(n9656), .dinb(n1620), .dout(n13057));
  jand g12990(.dina(n9250), .dinb(n1612), .dout(n13058));
  jand g12991(.dina(n8936), .dinb(n1644), .dout(n13059));
  jor  g12992(.dina(n13059), .dinb(n13058), .dout(n13060));
  jor  g12993(.dina(n13060), .dinb(n13057), .dout(n13061));
  jor  g12994(.dina(n13061), .dinb(n13056), .dout(n13062));
  jxor g12995(.dina(n13062), .dinb(n65), .dout(n13063));
  jxor g12996(.dina(n13063), .dinb(n13055), .dout(n13064));
  jxor g12997(.dina(n13064), .dinb(n13027), .dout(n13065));
  jnot g12998(.din(n13065), .dout(n13066));
  jand g12999(.dina(n10307), .dinb(n1819), .dout(n13067));
  jand g13000(.dina(n10305), .dinb(n2243), .dout(n13068));
  jand g13001(.dina(n9872), .dinb(n2180), .dout(n13069));
  jand g13002(.dina(n9655), .dinb(n2185), .dout(n13070));
  jor  g13003(.dina(n13070), .dinb(n13069), .dout(n13071));
  jor  g13004(.dina(n13071), .dinb(n13068), .dout(n13072));
  jor  g13005(.dina(n13072), .dinb(n13067), .dout(n13073));
  jxor g13006(.dina(n13073), .dinb(n2196), .dout(n13074));
  jxor g13007(.dina(n13074), .dinb(n13066), .dout(n13075));
  jxor g13008(.dina(n13075), .dinb(n13022), .dout(n13076));
  jnot g13009(.din(n13076), .dout(n13077));
  jand g13010(.dina(n10838), .dinb(n2743), .dout(n13078));
  jand g13011(.dina(n10836), .dinb(n2752), .dout(n13079));
  jand g13012(.dina(n10640), .dinb(n2748), .dout(n13080));
  jand g13013(.dina(n10647), .dinb(n2757), .dout(n13081));
  jor  g13014(.dina(n13081), .dinb(n13080), .dout(n13082));
  jor  g13015(.dina(n13082), .dinb(n13079), .dout(n13083));
  jor  g13016(.dina(n13083), .dinb(n13078), .dout(n13084));
  jxor g13017(.dina(n13084), .dinb(n2441), .dout(n13085));
  jxor g13018(.dina(n13085), .dinb(n13077), .dout(n13086));
  jxor g13019(.dina(n13086), .dinb(n13019), .dout(n13087));
  jnot g13020(.din(n13087), .dout(n13088));
  jand g13021(.dina(n11812), .dinb(n3423), .dout(n13089));
  jand g13022(.dina(n11646), .dinb(n3569), .dout(n13090));
  jand g13023(.dina(n11647), .dinb(n3428), .dout(n13091));
  jand g13024(.dina(n11306), .dinb(n3210), .dout(n13092));
  jor  g13025(.dina(n13092), .dinb(n13091), .dout(n13093));
  jor  g13026(.dina(n13093), .dinb(n13090), .dout(n13094));
  jor  g13027(.dina(n13094), .dinb(n13089), .dout(n13095));
  jxor g13028(.dina(n13095), .dinb(n3473), .dout(n13096));
  jxor g13029(.dina(n13096), .dinb(n13088), .dout(n13097));
  jxor g13030(.dina(n13097), .dinb(n13014), .dout(n13098));
  jand g13031(.dina(n12696), .dinb(n4022), .dout(n13099));
  jand g13032(.dina(n12547), .dinb(n4220), .dout(n13100));
  jand g13033(.dina(n12282), .dinb(n4027), .dout(n13101));
  jand g13034(.dina(n11798), .dinb(n3870), .dout(n13102));
  jor  g13035(.dina(n13102), .dinb(n13101), .dout(n13103));
  jor  g13036(.dina(n13103), .dinb(n13100), .dout(n13104));
  jor  g13037(.dina(n13104), .dinb(n13099), .dout(n13105));
  jxor g13038(.dina(n13105), .dinb(n4050), .dout(n13106));
  jxor g13039(.dina(n13106), .dinb(n13098), .dout(n13107));
  jxor g13040(.dina(n13107), .dinb(n13009), .dout(n13108));
  jand g13041(.dina(n12669), .dinb(n12536), .dout(n13109));
  jand g13042(.dina(n12670), .dinb(n12558), .dout(n13110));
  jor  g13043(.dina(n13110), .dinb(n13109), .dout(n13111));
  jor  g13044(.dina(n12571), .dinb(n12567), .dout(n13112));
  jand g13045(.dina(n12661), .dinb(n12572), .dout(n13113));
  jnot g13046(.din(n13113), .dout(n13114));
  jand g13047(.dina(n13114), .dinb(n13112), .dout(n13115));
  jnot g13048(.din(n13115), .dout(n13116));
  jand g13049(.dina(n12650), .dinb(n12575), .dout(n13117));
  jnot g13050(.din(n13117), .dout(n13118));
  jor  g13051(.dina(n12660), .dinb(n12652), .dout(n13119));
  jand g13052(.dina(n13119), .dinb(n13118), .dout(n13120));
  jor  g13053(.dina(n7301), .dinb(n1617), .dout(n13121));
  jor  g13054(.dina(n8002), .dinb(n807), .dout(n13122));
  jor  g13055(.dina(n7999), .dinb(n1621), .dout(n13123));
  jor  g13056(.dina(n7680), .dinb(n1613), .dout(n13124));
  jand g13057(.dina(n13124), .dinb(n13123), .dout(n13125));
  jand g13058(.dina(n13125), .dinb(n13122), .dout(n13126));
  jand g13059(.dina(n13126), .dinb(n13121), .dout(n13127));
  jxor g13060(.dina(n13127), .dinb(\a[23] ), .dout(n13128));
  jxor g13061(.dina(n13128), .dinb(n13120), .dout(n13129));
  jor  g13062(.dina(n12640), .dinb(n12632), .dout(n13130));
  jand g13063(.dina(n12649), .dinb(n12641), .dout(n13131));
  jnot g13064(.din(n13131), .dout(n13132));
  jand g13065(.dina(n13132), .dinb(n13130), .dout(n13133));
  jnot g13066(.din(n13133), .dout(n13134));
  jand g13067(.dina(n12624), .dinb(n12579), .dout(n13135));
  jnot g13068(.din(n13135), .dout(n13136));
  jor  g13069(.dina(n12630), .dinb(n12626), .dout(n13137));
  jand g13070(.dina(n13137), .dinb(n13136), .dout(n13138));
  jnot g13071(.din(n13138), .dout(n13139));
  jor  g13072(.dina(n5560), .dinb(n7061), .dout(n13140));
  jand g13073(.dina(n6050), .dinb(n5163), .dout(n13141));
  jand g13074(.dina(n5423), .dinb(n5084), .dout(n13142));
  jor  g13075(.dina(n13142), .dinb(n13141), .dout(n13143));
  jand g13076(.dina(n5426), .dinb(n5082), .dout(n13144));
  jor  g13077(.dina(n13144), .dinb(n13143), .dout(n13145));
  jnot g13078(.din(n13145), .dout(n13146));
  jand g13079(.dina(n13146), .dinb(n13140), .dout(n13147));
  jnot g13080(.din(n13147), .dout(n13148));
  jor  g13081(.dina(n12622), .dinb(n12474), .dout(n13149));
  jand g13082(.dina(n12623), .dinb(n12588), .dout(n13150));
  jnot g13083(.din(n13150), .dout(n13151));
  jand g13084(.dina(n13151), .dinb(n13149), .dout(n13152));
  jnot g13085(.din(n13152), .dout(n13153));
  jand g13086(.dina(n440), .dinb(n964), .dout(n13154));
  jand g13087(.dina(n13154), .dinb(n6192), .dout(n13155));
  jand g13088(.dina(n7649), .dinb(n4428), .dout(n13156));
  jand g13089(.dina(n1536), .dinb(n501), .dout(n13157));
  jand g13090(.dina(n619), .dinb(n266), .dout(n13158));
  jand g13091(.dina(n13158), .dinb(n13157), .dout(n13159));
  jand g13092(.dina(n13159), .dinb(n13156), .dout(n13160));
  jand g13093(.dina(n1219), .dinb(n1495), .dout(n13161));
  jand g13094(.dina(n13161), .dinb(n662), .dout(n13162));
  jand g13095(.dina(n13162), .dinb(n13160), .dout(n13163));
  jand g13096(.dina(n13163), .dinb(n13155), .dout(n13164));
  jand g13097(.dina(n5487), .dinb(n2409), .dout(n13165));
  jand g13098(.dina(n13165), .dinb(n1562), .dout(n13166));
  jand g13099(.dina(n13166), .dinb(n514), .dout(n13167));
  jand g13100(.dina(n13167), .dinb(n6359), .dout(n13168));
  jand g13101(.dina(n13168), .dinb(n13164), .dout(n13169));
  jand g13102(.dina(n1765), .dinb(n1288), .dout(n13170));
  jand g13103(.dina(n5499), .dinb(n809), .dout(n13171));
  jand g13104(.dina(n13171), .dinb(n13170), .dout(n13172));
  jand g13105(.dina(n1005), .dinb(n929), .dout(n13173));
  jand g13106(.dina(n13173), .dinb(n6441), .dout(n13174));
  jand g13107(.dina(n13174), .dinb(n1453), .dout(n13175));
  jand g13108(.dina(n9545), .dinb(n670), .dout(n13176));
  jand g13109(.dina(n13176), .dinb(n1743), .dout(n13177));
  jand g13110(.dina(n13177), .dinb(n13175), .dout(n13178));
  jand g13111(.dina(n13178), .dinb(n13172), .dout(n13179));
  jand g13112(.dina(n2106), .dinb(n934), .dout(n13180));
  jand g13113(.dina(n2087), .dinb(n1284), .dout(n13181));
  jand g13114(.dina(n13181), .dinb(n13180), .dout(n13182));
  jand g13115(.dina(n4585), .dinb(n838), .dout(n13183));
  jand g13116(.dina(n1577), .dinb(n548), .dout(n13184));
  jand g13117(.dina(n13184), .dinb(n1379), .dout(n13185));
  jand g13118(.dina(n13185), .dinb(n13183), .dout(n13186));
  jand g13119(.dina(n9756), .dinb(n2019), .dout(n13187));
  jand g13120(.dina(n13187), .dinb(n2131), .dout(n13188));
  jand g13121(.dina(n13188), .dinb(n13186), .dout(n13189));
  jand g13122(.dina(n13189), .dinb(n13182), .dout(n13190));
  jand g13123(.dina(n13190), .dinb(n13179), .dout(n13191));
  jand g13124(.dina(n1167), .dinb(n1541), .dout(n13192));
  jand g13125(.dina(n13192), .dinb(n1998), .dout(n13193));
  jand g13126(.dina(n1451), .dinb(n880), .dout(n13194));
  jand g13127(.dina(n13194), .dinb(n907), .dout(n13195));
  jand g13128(.dina(n13195), .dinb(n135), .dout(n13196));
  jand g13129(.dina(n1246), .dinb(n1098), .dout(n13197));
  jand g13130(.dina(n13197), .dinb(n1477), .dout(n13198));
  jand g13131(.dina(n948), .dinb(n1432), .dout(n13199));
  jand g13132(.dina(n13199), .dinb(n715), .dout(n13200));
  jand g13133(.dina(n13200), .dinb(n13198), .dout(n13201));
  jand g13134(.dina(n13201), .dinb(n13196), .dout(n13202));
  jand g13135(.dina(n2522), .dinb(n1778), .dout(n13203));
  jand g13136(.dina(n13203), .dinb(n13202), .dout(n13204));
  jand g13137(.dina(n13204), .dinb(n13193), .dout(n13205));
  jand g13138(.dina(n13205), .dinb(n13191), .dout(n13206));
  jand g13139(.dina(n13206), .dinb(n9742), .dout(n13207));
  jand g13140(.dina(n13207), .dinb(n13169), .dout(n13208));
  jand g13141(.dina(n13208), .dinb(n12473), .dout(n13209));
  jnot g13142(.din(n13209), .dout(n13210));
  jor  g13143(.dina(n13208), .dinb(n12473), .dout(n13211));
  jand g13144(.dina(n13211), .dinb(n2196), .dout(n13212));
  jand g13145(.dina(n13212), .dinb(n13210), .dout(n13213));
  jnot g13146(.din(n13213), .dout(n13214));
  jand g13147(.dina(n13214), .dinb(n2196), .dout(n13215));
  jand g13148(.dina(n13214), .dinb(n13211), .dout(n13216));
  jand g13149(.dina(n13216), .dinb(n13210), .dout(n13217));
  jor  g13150(.dina(n13217), .dinb(n13215), .dout(n13218));
  jxor g13151(.dina(n13218), .dinb(n13153), .dout(n13219));
  jxor g13152(.dina(n13219), .dinb(n13148), .dout(n13220));
  jor  g13153(.dina(n6207), .dinb(n4343), .dout(n13221));
  jor  g13154(.dina(n5525), .dinb(n4346), .dout(n13222));
  jor  g13155(.dina(n5364), .dinb(n3683), .dout(n13223));
  jor  g13156(.dina(n6205), .dinb(n4348), .dout(n13224));
  jand g13157(.dina(n13224), .dinb(n13223), .dout(n13225));
  jand g13158(.dina(n13225), .dinb(n13222), .dout(n13226));
  jand g13159(.dina(n13226), .dinb(n13221), .dout(n13227));
  jxor g13160(.dina(n13227), .dinb(n93), .dout(n13228));
  jxor g13161(.dina(n13228), .dinb(n13220), .dout(n13229));
  jxor g13162(.dina(n13229), .dinb(n13139), .dout(n13230));
  jor  g13163(.dina(n6491), .dinb(n2303), .dout(n13231));
  jor  g13164(.dina(n6297), .dinb(n2306), .dout(n13232));
  jor  g13165(.dina(n6390), .dinb(n1805), .dout(n13233));
  jor  g13166(.dina(n6489), .dinb(n2309), .dout(n13234));
  jand g13167(.dina(n13234), .dinb(n13233), .dout(n13235));
  jand g13168(.dina(n13235), .dinb(n13232), .dout(n13236));
  jand g13169(.dina(n13236), .dinb(n13231), .dout(n13237));
  jxor g13170(.dina(n13237), .dinb(n77), .dout(n13238));
  jxor g13171(.dina(n13238), .dinb(n13230), .dout(n13239));
  jxor g13172(.dina(n13239), .dinb(n13134), .dout(n13240));
  jxor g13173(.dina(n13240), .dinb(n13129), .dout(n13241));
  jxor g13174(.dina(n13241), .dinb(n13116), .dout(n13242));
  jnot g13175(.din(n13242), .dout(n13243));
  jand g13176(.dina(n12662), .dinb(n12563), .dout(n13244));
  jnot g13177(.din(n13244), .dout(n13245));
  jor  g13178(.dina(n12668), .dinb(n12664), .dout(n13246));
  jand g13179(.dina(n13246), .dinb(n13245), .dout(n13247));
  jxor g13180(.dina(n13247), .dinb(n13243), .dout(n13248));
  jxor g13181(.dina(n13248), .dinb(n12669), .dout(n13249));
  jxor g13182(.dina(n13249), .dinb(n13111), .dout(n13250));
  jand g13183(.dina(n13250), .dinb(n4691), .dout(n13251));
  jand g13184(.dina(n13248), .dinb(n4941), .dout(n13252));
  jand g13185(.dina(n12669), .dinb(n4696), .dout(n13253));
  jand g13186(.dina(n12536), .dinb(n4701), .dout(n13254));
  jor  g13187(.dina(n13254), .dinb(n13253), .dout(n13255));
  jor  g13188(.dina(n13255), .dinb(n13252), .dout(n13256));
  jor  g13189(.dina(n13256), .dinb(n13251), .dout(n13257));
  jxor g13190(.dina(n13257), .dinb(n4713), .dout(n13258));
  jxor g13191(.dina(n13258), .dinb(n13108), .dout(n13259));
  jnot g13192(.din(n13259), .dout(n13260));
  jxor g13193(.dina(n13260), .dinb(n13005), .dout(n13261));
  jnot g13194(.din(n13261), .dout(n13262));
  jand g13195(.dina(n13238), .dinb(n13230), .dout(n13263));
  jand g13196(.dina(n13239), .dinb(n13134), .dout(n13264));
  jor  g13197(.dina(n13264), .dinb(n13263), .dout(n13265));
  jand g13198(.dina(n13228), .dinb(n13220), .dout(n13266));
  jand g13199(.dina(n13229), .dinb(n13139), .dout(n13267));
  jor  g13200(.dina(n13267), .dinb(n13266), .dout(n13268));
  jand g13201(.dina(n13218), .dinb(n13153), .dout(n13269));
  jand g13202(.dina(n13219), .dinb(n13148), .dout(n13270));
  jor  g13203(.dina(n13270), .dinb(n13269), .dout(n13271));
  jor  g13204(.dina(n5549), .dinb(n7061), .dout(n13272));
  jand g13205(.dina(n6050), .dinb(n5426), .dout(n13273));
  jand g13206(.dina(n5365), .dinb(n5084), .dout(n13274));
  jor  g13207(.dina(n13274), .dinb(n13273), .dout(n13275));
  jand g13208(.dina(n5423), .dinb(n5082), .dout(n13276));
  jor  g13209(.dina(n13276), .dinb(n13275), .dout(n13277));
  jnot g13210(.din(n13277), .dout(n13278));
  jand g13211(.dina(n13278), .dinb(n13272), .dout(n13279));
  jnot g13212(.din(n13279), .dout(n13280));
  jand g13213(.dina(n4629), .dinb(n328), .dout(n13281));
  jand g13214(.dina(n2101), .dinb(n824), .dout(n13282));
  jand g13215(.dina(n13282), .dinb(n5408), .dout(n13283));
  jand g13216(.dina(n13283), .dinb(n13281), .dout(n13284));
  jand g13217(.dina(n1327), .dinb(n1284), .dout(n13285));
  jand g13218(.dina(n13285), .dinb(n1160), .dout(n13286));
  jand g13219(.dina(n13286), .dinb(n1257), .dout(n13287));
  jand g13220(.dina(n13287), .dinb(n13284), .dout(n13288));
  jand g13221(.dina(n12456), .dinb(n447), .dout(n13289));
  jand g13222(.dina(n1351), .dinb(n351), .dout(n13290));
  jand g13223(.dina(n320), .dinb(n492), .dout(n13291));
  jand g13224(.dina(n13291), .dinb(n13290), .dout(n13292));
  jand g13225(.dina(n13292), .dinb(n632), .dout(n13293));
  jand g13226(.dina(n13293), .dinb(n13289), .dout(n13294));
  jand g13227(.dina(n6441), .dinb(n480), .dout(n13295));
  jand g13228(.dina(n13295), .dinb(n10715), .dout(n13296));
  jand g13229(.dina(n13296), .dinb(n13294), .dout(n13297));
  jand g13230(.dina(n13297), .dinb(n4566), .dout(n13298));
  jand g13231(.dina(n13298), .dinb(n5247), .dout(n13299));
  jand g13232(.dina(n13299), .dinb(n13288), .dout(n13300));
  jand g13233(.dina(n1541), .dinb(n130), .dout(n13301));
  jand g13234(.dina(n13301), .dinb(n1207), .dout(n13302));
  jand g13235(.dina(n13302), .dinb(n6269), .dout(n13303));
  jand g13236(.dina(n3066), .dinb(n695), .dout(n13304));
  jand g13237(.dina(n6443), .dinb(n3827), .dout(n13305));
  jand g13238(.dina(n13305), .dinb(n13304), .dout(n13306));
  jand g13239(.dina(n13306), .dinb(n13303), .dout(n13307));
  jand g13240(.dina(n696), .dinb(n1279), .dout(n13308));
  jand g13241(.dina(n829), .dinb(n1309), .dout(n13309));
  jand g13242(.dina(n13309), .dinb(n648), .dout(n13310));
  jand g13243(.dina(n13310), .dinb(n3167), .dout(n13311));
  jand g13244(.dina(n13311), .dinb(n13308), .dout(n13312));
  jand g13245(.dina(n1219), .dinb(n1288), .dout(n13313));
  jand g13246(.dina(n2149), .dinb(n122), .dout(n13314));
  jand g13247(.dina(n452), .dinb(n1334), .dout(n13315));
  jand g13248(.dina(n13315), .dinb(n8120), .dout(n13316));
  jand g13249(.dina(n13316), .dinb(n13314), .dout(n13317));
  jand g13250(.dina(n13317), .dinb(n13313), .dout(n13318));
  jand g13251(.dina(n13318), .dinb(n13312), .dout(n13319));
  jand g13252(.dina(n13319), .dinb(n13307), .dout(n13320));
  jand g13253(.dina(n13320), .dinb(n1986), .dout(n13321));
  jand g13254(.dina(n13321), .dinb(n13300), .dout(n13322));
  jnot g13255(.din(n13322), .dout(n13323));
  jxor g13256(.dina(n13323), .dinb(n13216), .dout(n13324));
  jxor g13257(.dina(n13324), .dinb(n13280), .dout(n13325));
  jxor g13258(.dina(n13325), .dinb(n13271), .dout(n13326));
  jor  g13259(.dina(n6516), .dinb(n4343), .dout(n13327));
  jor  g13260(.dina(n6205), .dinb(n4346), .dout(n13328));
  jor  g13261(.dina(n5525), .dinb(n3683), .dout(n13329));
  jor  g13262(.dina(n6390), .dinb(n4348), .dout(n13330));
  jand g13263(.dina(n13330), .dinb(n13329), .dout(n13331));
  jand g13264(.dina(n13331), .dinb(n13328), .dout(n13332));
  jand g13265(.dina(n13332), .dinb(n13327), .dout(n13333));
  jxor g13266(.dina(n13333), .dinb(n93), .dout(n13334));
  jxor g13267(.dina(n13334), .dinb(n13326), .dout(n13335));
  jxor g13268(.dina(n13335), .dinb(n13268), .dout(n13336));
  jor  g13269(.dina(n7303), .dinb(n2303), .dout(n13337));
  jor  g13270(.dina(n7301), .dinb(n2309), .dout(n13338));
  jor  g13271(.dina(n6297), .dinb(n1805), .dout(n13339));
  jor  g13272(.dina(n6489), .dinb(n2306), .dout(n13340));
  jand g13273(.dina(n13340), .dinb(n13339), .dout(n13341));
  jand g13274(.dina(n13341), .dinb(n13338), .dout(n13342));
  jand g13275(.dina(n13342), .dinb(n13337), .dout(n13343));
  jxor g13276(.dina(n13343), .dinb(n77), .dout(n13344));
  jxor g13277(.dina(n13344), .dinb(n13336), .dout(n13345));
  jand g13278(.dina(n13345), .dinb(n13265), .dout(n13346));
  jnot g13279(.din(n13346), .dout(n13347));
  jxor g13280(.dina(n13345), .dinb(n13265), .dout(n13348));
  jnot g13281(.din(n13348), .dout(n13349));
  jor  g13282(.dina(n7999), .dinb(n1613), .dout(n13350));
  jor  g13283(.dina(n8260), .dinb(n807), .dout(n13351));
  jor  g13284(.dina(n7680), .dinb(n1617), .dout(n13352));
  jand g13285(.dina(n13352), .dinb(n13351), .dout(n13353));
  jand g13286(.dina(n13353), .dinb(n13350), .dout(n13354));
  jxor g13287(.dina(n13354), .dinb(\a[23] ), .dout(n13355));
  jor  g13288(.dina(n13355), .dinb(n13349), .dout(n13356));
  jand g13289(.dina(n13356), .dinb(n13347), .dout(n13357));
  jnot g13290(.din(n13357), .dout(n13358));
  jand g13291(.dina(n13335), .dinb(n13268), .dout(n13359));
  jand g13292(.dina(n13344), .dinb(n13336), .dout(n13360));
  jor  g13293(.dina(n13360), .dinb(n13359), .dout(n13361));
  jnot g13294(.din(n13361), .dout(n13362));
  jand g13295(.dina(n8256), .dinb(n806), .dout(n13363));
  jor  g13296(.dina(n13363), .dinb(n1644), .dout(n13364));
  jand g13297(.dina(n13364), .dinb(n8000), .dout(n13365));
  jxor g13298(.dina(n13365), .dinb(n65), .dout(n13366));
  jxor g13299(.dina(n13366), .dinb(n13362), .dout(n13367));
  jand g13300(.dina(n13325), .dinb(n13271), .dout(n13368));
  jand g13301(.dina(n13334), .dinb(n13326), .dout(n13369));
  jor  g13302(.dina(n13369), .dinb(n13368), .dout(n13370));
  jor  g13303(.dina(n5527), .dinb(n7061), .dout(n13371));
  jand g13304(.dina(n6050), .dinb(n5423), .dout(n13372));
  jand g13305(.dina(n6140), .dinb(n5084), .dout(n13373));
  jor  g13306(.dina(n13373), .dinb(n13372), .dout(n13374));
  jand g13307(.dina(n5365), .dinb(n5082), .dout(n13375));
  jor  g13308(.dina(n13375), .dinb(n13374), .dout(n13376));
  jnot g13309(.din(n13376), .dout(n13377));
  jand g13310(.dina(n13377), .dinb(n13371), .dout(n13378));
  jnot g13311(.din(n13378), .dout(n13379));
  jnot g13312(.din(n13216), .dout(n13380));
  jand g13313(.dina(n13322), .dinb(n13380), .dout(n13381));
  jand g13314(.dina(n13324), .dinb(n13280), .dout(n13382));
  jor  g13315(.dina(n13382), .dinb(n13381), .dout(n13383));
  jand g13316(.dina(n10714), .dinb(n10533), .dout(n13384));
  jand g13317(.dina(n557), .dinb(n811), .dout(n13385));
  jand g13318(.dina(n13385), .dinb(n6031), .dout(n13386));
  jand g13319(.dina(n13386), .dinb(n1453), .dout(n13387));
  jand g13320(.dina(n13387), .dinb(n1211), .dout(n13388));
  jand g13321(.dina(n5487), .dinb(n1225), .dout(n13389));
  jand g13322(.dina(n931), .dinb(n680), .dout(n13390));
  jand g13323(.dina(n13390), .dinb(n1288), .dout(n13391));
  jand g13324(.dina(n13391), .dinb(n13389), .dout(n13392));
  jand g13325(.dina(n3306), .dinb(n1933), .dout(n13393));
  jand g13326(.dina(n13393), .dinb(n13392), .dout(n13394));
  jand g13327(.dina(n1361), .dinb(n948), .dout(n13395));
  jand g13328(.dina(n1536), .dinb(n481), .dout(n13396));
  jand g13329(.dina(n13396), .dinb(n2020), .dout(n13397));
  jand g13330(.dina(n13397), .dinb(n13395), .dout(n13398));
  jand g13331(.dina(n13398), .dinb(n13394), .dout(n13399));
  jand g13332(.dina(n13399), .dinb(n13388), .dout(n13400));
  jand g13333(.dina(n13400), .dinb(n13384), .dout(n13401));
  jand g13334(.dina(n670), .dinb(n1591), .dout(n13402));
  jand g13335(.dina(n1375), .dinb(n991), .dout(n13403));
  jand g13336(.dina(n13403), .dinb(n13402), .dout(n13404));
  jand g13337(.dina(n13404), .dinb(n917), .dout(n13405));
  jand g13338(.dina(n716), .dinb(n639), .dout(n13406));
  jand g13339(.dina(n13406), .dinb(n981), .dout(n13407));
  jand g13340(.dina(n1344), .dinb(n517), .dout(n13408));
  jand g13341(.dina(n647), .dinb(n1226), .dout(n13409));
  jand g13342(.dina(n13409), .dinb(n13408), .dout(n13410));
  jand g13343(.dina(n13410), .dinb(n13407), .dout(n13411));
  jand g13344(.dina(n13411), .dinb(n13405), .dout(n13412));
  jand g13345(.dina(n4448), .dinb(n3758), .dout(n13413));
  jand g13346(.dina(n13413), .dinb(n1579), .dout(n13414));
  jand g13347(.dina(n13414), .dinb(n13412), .dout(n13415));
  jand g13348(.dina(n3324), .dinb(n541), .dout(n13416));
  jand g13349(.dina(n13416), .dinb(n100), .dout(n13417));
  jand g13350(.dina(n13417), .dinb(n9750), .dout(n13418));
  jand g13351(.dina(n1713), .dinb(n521), .dout(n13419));
  jand g13352(.dina(n884), .dinb(n1088), .dout(n13420));
  jand g13353(.dina(n13420), .dinb(n13419), .dout(n13421));
  jand g13354(.dina(n13421), .dinb(n1439), .dout(n13422));
  jand g13355(.dina(n13422), .dinb(n2665), .dout(n13423));
  jand g13356(.dina(n13423), .dinb(n13418), .dout(n13424));
  jand g13357(.dina(n13424), .dinb(n13415), .dout(n13425));
  jand g13358(.dina(n13425), .dinb(n13401), .dout(n13426));
  jxor g13359(.dina(n13426), .dinb(n13323), .dout(n13427));
  jxor g13360(.dina(n13427), .dinb(n13383), .dout(n13428));
  jxor g13361(.dina(n13428), .dinb(n13379), .dout(n13429));
  jxor g13362(.dina(n13429), .dinb(n13370), .dout(n13430));
  jnot g13363(.din(n13430), .dout(n13431));
  jor  g13364(.dina(n6999), .dinb(n4343), .dout(n13432));
  jor  g13365(.dina(n6390), .dinb(n4346), .dout(n13433));
  jor  g13366(.dina(n6297), .dinb(n4348), .dout(n13434));
  jand g13367(.dina(n13434), .dinb(n13433), .dout(n13435));
  jor  g13368(.dina(n6205), .dinb(n3683), .dout(n13436));
  jand g13369(.dina(n13436), .dinb(n13435), .dout(n13437));
  jand g13370(.dina(n13437), .dinb(n13432), .dout(n13438));
  jxor g13371(.dina(n13438), .dinb(\a[29] ), .dout(n13439));
  jxor g13372(.dina(n13439), .dinb(n13431), .dout(n13440));
  jor  g13373(.dina(n7682), .dinb(n2303), .dout(n13441));
  jor  g13374(.dina(n7301), .dinb(n2306), .dout(n13442));
  jor  g13375(.dina(n7680), .dinb(n2309), .dout(n13443));
  jor  g13376(.dina(n6489), .dinb(n1805), .dout(n13444));
  jand g13377(.dina(n13444), .dinb(n13443), .dout(n13445));
  jand g13378(.dina(n13445), .dinb(n13442), .dout(n13446));
  jand g13379(.dina(n13446), .dinb(n13441), .dout(n13447));
  jxor g13380(.dina(n13447), .dinb(n77), .dout(n13448));
  jxor g13381(.dina(n13448), .dinb(n13440), .dout(n13449));
  jxor g13382(.dina(n13449), .dinb(n13367), .dout(n13450));
  jxor g13383(.dina(n13450), .dinb(n13358), .dout(n13451));
  jnot g13384(.din(n13451), .dout(n13452));
  jor  g13385(.dina(n13128), .dinb(n13120), .dout(n13453));
  jand g13386(.dina(n13240), .dinb(n13129), .dout(n13454));
  jnot g13387(.din(n13454), .dout(n13455));
  jand g13388(.dina(n13455), .dinb(n13453), .dout(n13456));
  jnot g13389(.din(n13456), .dout(n13457));
  jxor g13390(.dina(n13355), .dinb(n13349), .dout(n13458));
  jand g13391(.dina(n13458), .dinb(n13457), .dout(n13459));
  jnot g13392(.din(n13459), .dout(n13460));
  jand g13393(.dina(n13241), .dinb(n13116), .dout(n13461));
  jnot g13394(.din(n13461), .dout(n13462));
  jor  g13395(.dina(n13247), .dinb(n13243), .dout(n13463));
  jand g13396(.dina(n13463), .dinb(n13462), .dout(n13464));
  jxor g13397(.dina(n13458), .dinb(n13457), .dout(n13465));
  jnot g13398(.din(n13465), .dout(n13466));
  jor  g13399(.dina(n13466), .dinb(n13464), .dout(n13467));
  jand g13400(.dina(n13467), .dinb(n13460), .dout(n13468));
  jxor g13401(.dina(n13468), .dinb(n13452), .dout(n13469));
  jand g13402(.dina(n12532), .dinb(n12546), .dout(n13470));
  jor  g13403(.dina(n13470), .dinb(n12526), .dout(n13471));
  jand g13404(.dina(n13471), .dinb(n12518), .dout(n13472));
  jor  g13405(.dina(n13472), .dinb(n12665), .dout(n13473));
  jand g13406(.dina(n13473), .dinb(n12663), .dout(n13474));
  jor  g13407(.dina(n13474), .dinb(n13244), .dout(n13475));
  jand g13408(.dina(n13475), .dinb(n13242), .dout(n13476));
  jor  g13409(.dina(n13476), .dinb(n13461), .dout(n13477));
  jxor g13410(.dina(n13465), .dinb(n13477), .dout(n13478));
  jand g13411(.dina(n13478), .dinb(n13469), .dout(n13479));
  jand g13412(.dina(n13478), .dinb(n13248), .dout(n13480));
  jand g13413(.dina(n13248), .dinb(n12669), .dout(n13481));
  jand g13414(.dina(n13249), .dinb(n13111), .dout(n13482));
  jor  g13415(.dina(n13482), .dinb(n13481), .dout(n13483));
  jxor g13416(.dina(n13478), .dinb(n13248), .dout(n13484));
  jand g13417(.dina(n13484), .dinb(n13483), .dout(n13485));
  jor  g13418(.dina(n13485), .dinb(n13480), .dout(n13486));
  jxor g13419(.dina(n13478), .dinb(n13469), .dout(n13487));
  jand g13420(.dina(n13487), .dinb(n13486), .dout(n13488));
  jor  g13421(.dina(n13488), .dinb(n13479), .dout(n13489));
  jand g13422(.dina(n13450), .dinb(n13358), .dout(n13490));
  jand g13423(.dina(n13465), .dinb(n13477), .dout(n13491));
  jor  g13424(.dina(n13491), .dinb(n13459), .dout(n13492));
  jand g13425(.dina(n13492), .dinb(n13451), .dout(n13493));
  jor  g13426(.dina(n13493), .dinb(n13490), .dout(n13494));
  jor  g13427(.dina(n13366), .dinb(n13362), .dout(n13495));
  jand g13428(.dina(n13449), .dinb(n13367), .dout(n13496));
  jnot g13429(.din(n13496), .dout(n13497));
  jand g13430(.dina(n13497), .dinb(n13495), .dout(n13498));
  jnot g13431(.din(n13498), .dout(n13499));
  jand g13432(.dina(n13428), .dinb(n13379), .dout(n13500));
  jand g13433(.dina(n13429), .dinb(n13370), .dout(n13501));
  jor  g13434(.dina(n13501), .dinb(n13500), .dout(n13502));
  jand g13435(.dina(n13426), .dinb(n13323), .dout(n13503));
  jand g13436(.dina(n13427), .dinb(n13383), .dout(n13504));
  jor  g13437(.dina(n13504), .dinb(n13503), .dout(n13505));
  jand g13438(.dina(n6028), .dinb(n479), .dout(n13506));
  jand g13439(.dina(n1713), .dinb(n1476), .dout(n13507));
  jand g13440(.dina(n13507), .dinb(n5329), .dout(n13508));
  jand g13441(.dina(n13508), .dinb(n3384), .dout(n13509));
  jand g13442(.dina(n1351), .dinb(n1701), .dout(n13510));
  jand g13443(.dina(n13510), .dinb(n1328), .dout(n13511));
  jand g13444(.dina(n1305), .dinb(n171), .dout(n13512));
  jand g13445(.dina(n13512), .dinb(n179), .dout(n13513));
  jand g13446(.dina(n13513), .dinb(n1283), .dout(n13514));
  jand g13447(.dina(n13514), .dinb(n13511), .dout(n13515));
  jand g13448(.dina(n13515), .dinb(n13509), .dout(n13516));
  jand g13449(.dina(n3261), .dinb(n1561), .dout(n13517));
  jand g13450(.dina(n7243), .dinb(n328), .dout(n13518));
  jand g13451(.dina(n3995), .dinb(n818), .dout(n13519));
  jand g13452(.dina(n13519), .dinb(n122), .dout(n13520));
  jand g13453(.dina(n13520), .dinb(n13518), .dout(n13521));
  jand g13454(.dina(n884), .dinb(n991), .dout(n13522));
  jand g13455(.dina(n13522), .dinb(n848), .dout(n13523));
  jand g13456(.dina(n13523), .dinb(n2024), .dout(n13524));
  jand g13457(.dina(n13524), .dinb(n13521), .dout(n13525));
  jand g13458(.dina(n13525), .dinb(n13517), .dout(n13526));
  jand g13459(.dina(n13526), .dinb(n839), .dout(n13527));
  jand g13460(.dina(n13527), .dinb(n13516), .dout(n13528));
  jand g13461(.dina(n13528), .dinb(n13506), .dout(n13529));
  jand g13462(.dina(n1697), .dinb(n654), .dout(n13530));
  jand g13463(.dina(n1099), .dinb(n1037), .dout(n13531));
  jand g13464(.dina(n13531), .dinb(n11407), .dout(n13532));
  jand g13465(.dina(n13532), .dinb(n13530), .dout(n13533));
  jand g13466(.dina(n1465), .dinb(n1449), .dout(n13534));
  jand g13467(.dina(n13534), .dinb(n2154), .dout(n13535));
  jand g13468(.dina(n13535), .dinb(n1506), .dout(n13536));
  jand g13469(.dina(n6236), .dinb(n1370), .dout(n13537));
  jand g13470(.dina(n13537), .dinb(n1732), .dout(n13538));
  jand g13471(.dina(n13538), .dinb(n13536), .dout(n13539));
  jand g13472(.dina(n13539), .dinb(n13533), .dout(n13540));
  jand g13473(.dina(n442), .dinb(n450), .dout(n13541));
  jand g13474(.dina(n13541), .dinb(n1872), .dout(n13542));
  jand g13475(.dina(n13542), .dinb(n1583), .dout(n13543));
  jand g13476(.dina(n716), .dinb(n130), .dout(n13544));
  jand g13477(.dina(n495), .dinb(n1822), .dout(n13545));
  jand g13478(.dina(n13545), .dinb(n2100), .dout(n13546));
  jand g13479(.dina(n13546), .dinb(n13544), .dout(n13547));
  jand g13480(.dina(n13547), .dinb(n13543), .dout(n13548));
  jand g13481(.dina(n1189), .dinb(n699), .dout(n13549));
  jand g13482(.dina(n465), .dinb(n1270), .dout(n13550));
  jand g13483(.dina(n13550), .dinb(n13549), .dout(n13551));
  jand g13484(.dina(n13551), .dinb(n3969), .dout(n13552));
  jand g13485(.dina(n13552), .dinb(n13548), .dout(n13553));
  jand g13486(.dina(n562), .dinb(n534), .dout(n13554));
  jand g13487(.dina(n13554), .dinb(n9545), .dout(n13555));
  jand g13488(.dina(n13555), .dinb(n829), .dout(n13556));
  jand g13489(.dina(n13556), .dinb(n13553), .dout(n13557));
  jand g13490(.dina(n13557), .dinb(n13540), .dout(n13558));
  jand g13491(.dina(n988), .dinb(n1288), .dout(n13559));
  jand g13492(.dina(n13559), .dinb(n1245), .dout(n13560));
  jand g13493(.dina(n1042), .dinb(n983), .dout(n13561));
  jand g13494(.dina(n13561), .dinb(n3371), .dout(n13562));
  jand g13495(.dina(n13562), .dinb(n13560), .dout(n13563));
  jand g13496(.dina(n13563), .dinb(n881), .dout(n13564));
  jand g13497(.dina(n13564), .dinb(n13558), .dout(n13565));
  jand g13498(.dina(n13565), .dinb(n4488), .dout(n13566));
  jand g13499(.dina(n13566), .dinb(n13529), .dout(n13567));
  jand g13500(.dina(n13567), .dinb(n13426), .dout(n13568));
  jnot g13501(.din(n13568), .dout(n13569));
  jor  g13502(.dina(n13567), .dinb(n13426), .dout(n13570));
  jand g13503(.dina(n13570), .dinb(n65), .dout(n13571));
  jand g13504(.dina(n13571), .dinb(n13569), .dout(n13572));
  jnot g13505(.din(n13572), .dout(n13573));
  jand g13506(.dina(n13573), .dinb(n65), .dout(n13574));
  jand g13507(.dina(n13573), .dinb(n13570), .dout(n13575));
  jand g13508(.dina(n13575), .dinb(n13569), .dout(n13576));
  jor  g13509(.dina(n13576), .dinb(n13574), .dout(n13577));
  jnot g13510(.din(n13577), .dout(n13578));
  jor  g13511(.dina(n6207), .dinb(n7061), .dout(n13579));
  jand g13512(.dina(n6050), .dinb(n5365), .dout(n13580));
  jand g13513(.dina(n6394), .dinb(n5084), .dout(n13581));
  jor  g13514(.dina(n13581), .dinb(n13580), .dout(n13582));
  jand g13515(.dina(n6140), .dinb(n5082), .dout(n13583));
  jor  g13516(.dina(n13583), .dinb(n13582), .dout(n13584));
  jnot g13517(.din(n13584), .dout(n13585));
  jand g13518(.dina(n13585), .dinb(n13579), .dout(n13586));
  jxor g13519(.dina(n13586), .dinb(n13578), .dout(n13587));
  jxor g13520(.dina(n13587), .dinb(n13505), .dout(n13588));
  jxor g13521(.dina(n13588), .dinb(n13502), .dout(n13589));
  jor  g13522(.dina(n6491), .dinb(n4343), .dout(n13590));
  jor  g13523(.dina(n6297), .dinb(n4346), .dout(n13591));
  jor  g13524(.dina(n6390), .dinb(n3683), .dout(n13592));
  jor  g13525(.dina(n6489), .dinb(n4348), .dout(n13593));
  jand g13526(.dina(n13593), .dinb(n13592), .dout(n13594));
  jand g13527(.dina(n13594), .dinb(n13591), .dout(n13595));
  jand g13528(.dina(n13595), .dinb(n13590), .dout(n13596));
  jxor g13529(.dina(n13596), .dinb(n93), .dout(n13597));
  jxor g13530(.dina(n13597), .dinb(n13589), .dout(n13598));
  jor  g13531(.dina(n13439), .dinb(n13431), .dout(n13599));
  jand g13532(.dina(n13448), .dinb(n13440), .dout(n13600));
  jnot g13533(.din(n13600), .dout(n13601));
  jand g13534(.dina(n13601), .dinb(n13599), .dout(n13602));
  jor  g13535(.dina(n7301), .dinb(n1805), .dout(n13603));
  jor  g13536(.dina(n8002), .dinb(n2303), .dout(n13604));
  jor  g13537(.dina(n7999), .dinb(n2309), .dout(n13605));
  jor  g13538(.dina(n7680), .dinb(n2306), .dout(n13606));
  jand g13539(.dina(n13606), .dinb(n13605), .dout(n13607));
  jand g13540(.dina(n13607), .dinb(n13604), .dout(n13608));
  jand g13541(.dina(n13608), .dinb(n13603), .dout(n13609));
  jxor g13542(.dina(n13609), .dinb(\a[26] ), .dout(n13610));
  jxor g13543(.dina(n13610), .dinb(n13602), .dout(n13611));
  jxor g13544(.dina(n13611), .dinb(n13598), .dout(n13612));
  jxor g13545(.dina(n13612), .dinb(n13499), .dout(n13613));
  jxor g13546(.dina(n13613), .dinb(n13494), .dout(n13614));
  jxor g13547(.dina(n13614), .dinb(n13469), .dout(n13615));
  jxor g13548(.dina(n13615), .dinb(n13489), .dout(n13616));
  jand g13549(.dina(n13616), .dinb(n5280), .dout(n13617));
  jand g13550(.dina(n13614), .dinb(n5814), .dout(n13618));
  jand g13551(.dina(n13469), .dinb(n5531), .dout(n13619));
  jand g13552(.dina(n13478), .dinb(n5536), .dout(n13620));
  jor  g13553(.dina(n13620), .dinb(n13619), .dout(n13621));
  jor  g13554(.dina(n13621), .dinb(n13618), .dout(n13622));
  jor  g13555(.dina(n13622), .dinb(n13617), .dout(n13623));
  jxor g13556(.dina(n13623), .dinb(n5277), .dout(n13624));
  jor  g13557(.dina(n13624), .dinb(n13262), .dout(n13625));
  jxor g13558(.dina(n13003), .dinb(n13001), .dout(n13626));
  jxor g13559(.dina(n13487), .dinb(n13486), .dout(n13627));
  jand g13560(.dina(n13627), .dinb(n5280), .dout(n13628));
  jand g13561(.dina(n13469), .dinb(n5814), .dout(n13629));
  jand g13562(.dina(n13478), .dinb(n5531), .dout(n13630));
  jand g13563(.dina(n13248), .dinb(n5536), .dout(n13631));
  jor  g13564(.dina(n13631), .dinb(n13630), .dout(n13632));
  jor  g13565(.dina(n13632), .dinb(n13629), .dout(n13633));
  jor  g13566(.dina(n13633), .dinb(n13628), .dout(n13634));
  jxor g13567(.dina(n13634), .dinb(n5277), .dout(n13635));
  jor  g13568(.dina(n13635), .dinb(n13626), .dout(n13636));
  jnot g13569(.din(n13636), .dout(n13637));
  jxor g13570(.dina(n12998), .dinb(n12997), .dout(n13638));
  jxor g13571(.dina(n13484), .dinb(n13483), .dout(n13639));
  jand g13572(.dina(n13639), .dinb(n5280), .dout(n13640));
  jand g13573(.dina(n13248), .dinb(n5531), .dout(n13641));
  jand g13574(.dina(n13478), .dinb(n5814), .dout(n13642));
  jor  g13575(.dina(n13642), .dinb(n13641), .dout(n13643));
  jand g13576(.dina(n12669), .dinb(n5536), .dout(n13644));
  jor  g13577(.dina(n13644), .dinb(n13643), .dout(n13645));
  jor  g13578(.dina(n13645), .dinb(n13640), .dout(n13646));
  jxor g13579(.dina(n13646), .dinb(n5277), .dout(n13647));
  jor  g13580(.dina(n13647), .dinb(n13638), .dout(n13648));
  jnot g13581(.din(n13648), .dout(n13649));
  jxor g13582(.dina(n12994), .dinb(n12993), .dout(n13650));
  jand g13583(.dina(n13250), .dinb(n5280), .dout(n13651));
  jand g13584(.dina(n12669), .dinb(n5531), .dout(n13652));
  jand g13585(.dina(n13248), .dinb(n5814), .dout(n13653));
  jor  g13586(.dina(n13653), .dinb(n13652), .dout(n13654));
  jand g13587(.dina(n12536), .dinb(n5536), .dout(n13655));
  jor  g13588(.dina(n13655), .dinb(n13654), .dout(n13656));
  jor  g13589(.dina(n13656), .dinb(n13651), .dout(n13657));
  jxor g13590(.dina(n13657), .dinb(n5277), .dout(n13658));
  jor  g13591(.dina(n13658), .dinb(n13650), .dout(n13659));
  jnot g13592(.din(n13659), .dout(n13660));
  jxor g13593(.dina(n12991), .dinb(n12989), .dout(n13661));
  jand g13594(.dina(n12671), .dinb(n5280), .dout(n13662));
  jand g13595(.dina(n12669), .dinb(n5814), .dout(n13663));
  jand g13596(.dina(n12536), .dinb(n5531), .dout(n13664));
  jand g13597(.dina(n12547), .dinb(n5536), .dout(n13665));
  jor  g13598(.dina(n13665), .dinb(n13664), .dout(n13666));
  jor  g13599(.dina(n13666), .dinb(n13663), .dout(n13667));
  jor  g13600(.dina(n13667), .dinb(n13662), .dout(n13668));
  jxor g13601(.dina(n13668), .dinb(\a[5] ), .dout(n13669));
  jand g13602(.dina(n13669), .dinb(n13661), .dout(n13670));
  jnot g13603(.din(n12987), .dout(n13671));
  jxor g13604(.dina(n13671), .dinb(n12986), .dout(n13672));
  jand g13605(.dina(n12684), .dinb(n5280), .dout(n13673));
  jand g13606(.dina(n12547), .dinb(n5531), .dout(n13674));
  jand g13607(.dina(n12536), .dinb(n5814), .dout(n13675));
  jor  g13608(.dina(n13675), .dinb(n13674), .dout(n13676));
  jand g13609(.dina(n12282), .dinb(n5536), .dout(n13677));
  jor  g13610(.dina(n13677), .dinb(n13676), .dout(n13678));
  jor  g13611(.dina(n13678), .dinb(n13673), .dout(n13679));
  jxor g13612(.dina(n13679), .dinb(n5277), .dout(n13680));
  jor  g13613(.dina(n13680), .dinb(n13672), .dout(n13681));
  jnot g13614(.din(n13681), .dout(n13682));
  jnot g13615(.din(n12984), .dout(n13683));
  jxor g13616(.dina(n13683), .dinb(n12983), .dout(n13684));
  jand g13617(.dina(n12696), .dinb(n5280), .dout(n13685));
  jand g13618(.dina(n12547), .dinb(n5814), .dout(n13686));
  jand g13619(.dina(n12282), .dinb(n5531), .dout(n13687));
  jand g13620(.dina(n11798), .dinb(n5536), .dout(n13688));
  jor  g13621(.dina(n13688), .dinb(n13687), .dout(n13689));
  jor  g13622(.dina(n13689), .dinb(n13686), .dout(n13690));
  jor  g13623(.dina(n13690), .dinb(n13685), .dout(n13691));
  jxor g13624(.dina(n13691), .dinb(n5277), .dout(n13692));
  jor  g13625(.dina(n13692), .dinb(n13684), .dout(n13693));
  jnot g13626(.din(n13693), .dout(n13694));
  jnot g13627(.din(n12981), .dout(n13695));
  jxor g13628(.dina(n13695), .dinb(n12980), .dout(n13696));
  jand g13629(.dina(n12284), .dinb(n5280), .dout(n13697));
  jand g13630(.dina(n12282), .dinb(n5814), .dout(n13698));
  jand g13631(.dina(n11798), .dinb(n5531), .dout(n13699));
  jand g13632(.dina(n11646), .dinb(n5536), .dout(n13700));
  jor  g13633(.dina(n13700), .dinb(n13699), .dout(n13701));
  jor  g13634(.dina(n13701), .dinb(n13698), .dout(n13702));
  jor  g13635(.dina(n13702), .dinb(n13697), .dout(n13703));
  jxor g13636(.dina(n13703), .dinb(n5277), .dout(n13704));
  jor  g13637(.dina(n13704), .dinb(n13696), .dout(n13705));
  jnot g13638(.din(n13705), .dout(n13706));
  jnot g13639(.din(n12978), .dout(n13707));
  jxor g13640(.dina(n13707), .dinb(n12977), .dout(n13708));
  jand g13641(.dina(n11800), .dinb(n5280), .dout(n13709));
  jand g13642(.dina(n11646), .dinb(n5531), .dout(n13710));
  jand g13643(.dina(n11798), .dinb(n5814), .dout(n13711));
  jor  g13644(.dina(n13711), .dinb(n13710), .dout(n13712));
  jand g13645(.dina(n11647), .dinb(n5536), .dout(n13713));
  jor  g13646(.dina(n13713), .dinb(n13712), .dout(n13714));
  jor  g13647(.dina(n13714), .dinb(n13709), .dout(n13715));
  jxor g13648(.dina(n13715), .dinb(n5277), .dout(n13716));
  jor  g13649(.dina(n13716), .dinb(n13708), .dout(n13717));
  jnot g13650(.din(n13717), .dout(n13718));
  jnot g13651(.din(n12975), .dout(n13719));
  jxor g13652(.dina(n13719), .dinb(n12974), .dout(n13720));
  jand g13653(.dina(n11812), .dinb(n5280), .dout(n13721));
  jand g13654(.dina(n11646), .dinb(n5814), .dout(n13722));
  jand g13655(.dina(n11647), .dinb(n5531), .dout(n13723));
  jand g13656(.dina(n11306), .dinb(n5536), .dout(n13724));
  jor  g13657(.dina(n13724), .dinb(n13723), .dout(n13725));
  jor  g13658(.dina(n13725), .dinb(n13722), .dout(n13726));
  jor  g13659(.dina(n13726), .dinb(n13721), .dout(n13727));
  jxor g13660(.dina(n13727), .dinb(n5277), .dout(n13728));
  jor  g13661(.dina(n13728), .dinb(n13720), .dout(n13729));
  jnot g13662(.din(n13729), .dout(n13730));
  jxor g13663(.dina(n12971), .dinb(n12970), .dout(n13731));
  jnot g13664(.din(n13731), .dout(n13732));
  jand g13665(.dina(n11824), .dinb(n5280), .dout(n13733));
  jand g13666(.dina(n11647), .dinb(n5814), .dout(n13734));
  jand g13667(.dina(n11306), .dinb(n5531), .dout(n13735));
  jand g13668(.dina(n10836), .dinb(n5536), .dout(n13736));
  jor  g13669(.dina(n13736), .dinb(n13735), .dout(n13737));
  jor  g13670(.dina(n13737), .dinb(n13734), .dout(n13738));
  jor  g13671(.dina(n13738), .dinb(n13733), .dout(n13739));
  jxor g13672(.dina(n13739), .dinb(\a[5] ), .dout(n13740));
  jand g13673(.dina(n13740), .dinb(n13732), .dout(n13741));
  jxor g13674(.dina(n12968), .dinb(n12966), .dout(n13742));
  jnot g13675(.din(n13742), .dout(n13743));
  jand g13676(.dina(n11308), .dinb(n5280), .dout(n13744));
  jand g13677(.dina(n10836), .dinb(n5531), .dout(n13745));
  jand g13678(.dina(n11306), .dinb(n5814), .dout(n13746));
  jor  g13679(.dina(n13746), .dinb(n13745), .dout(n13747));
  jand g13680(.dina(n10640), .dinb(n5536), .dout(n13748));
  jor  g13681(.dina(n13748), .dinb(n13747), .dout(n13749));
  jor  g13682(.dina(n13749), .dinb(n13744), .dout(n13750));
  jxor g13683(.dina(n13750), .dinb(n5277), .dout(n13751));
  jor  g13684(.dina(n13751), .dinb(n13743), .dout(n13752));
  jxor g13685(.dina(n12964), .dinb(n12962), .dout(n13753));
  jnot g13686(.din(n13753), .dout(n13754));
  jand g13687(.dina(n10838), .dinb(n5280), .dout(n13755));
  jand g13688(.dina(n10640), .dinb(n5531), .dout(n13756));
  jand g13689(.dina(n10836), .dinb(n5814), .dout(n13757));
  jor  g13690(.dina(n13757), .dinb(n13756), .dout(n13758));
  jand g13691(.dina(n10647), .dinb(n5536), .dout(n13759));
  jor  g13692(.dina(n13759), .dinb(n13758), .dout(n13760));
  jor  g13693(.dina(n13760), .dinb(n13755), .dout(n13761));
  jxor g13694(.dina(n13761), .dinb(n5277), .dout(n13762));
  jor  g13695(.dina(n13762), .dinb(n13754), .dout(n13763));
  jxor g13696(.dina(n12960), .dinb(n12958), .dout(n13764));
  jnot g13697(.din(n13764), .dout(n13765));
  jand g13698(.dina(n10850), .dinb(n5280), .dout(n13766));
  jand g13699(.dina(n10640), .dinb(n5814), .dout(n13767));
  jand g13700(.dina(n10647), .dinb(n5531), .dout(n13768));
  jand g13701(.dina(n10305), .dinb(n5536), .dout(n13769));
  jor  g13702(.dina(n13769), .dinb(n13768), .dout(n13770));
  jor  g13703(.dina(n13770), .dinb(n13767), .dout(n13771));
  jor  g13704(.dina(n13771), .dinb(n13766), .dout(n13772));
  jxor g13705(.dina(n13772), .dinb(n5277), .dout(n13773));
  jor  g13706(.dina(n13773), .dinb(n13765), .dout(n13774));
  jxor g13707(.dina(n12956), .dinb(n12954), .dout(n13775));
  jnot g13708(.din(n13775), .dout(n13776));
  jand g13709(.dina(n10862), .dinb(n5280), .dout(n13777));
  jand g13710(.dina(n10305), .dinb(n5531), .dout(n13778));
  jand g13711(.dina(n10647), .dinb(n5814), .dout(n13779));
  jor  g13712(.dina(n13779), .dinb(n13778), .dout(n13780));
  jand g13713(.dina(n9872), .dinb(n5536), .dout(n13781));
  jor  g13714(.dina(n13781), .dinb(n13780), .dout(n13782));
  jor  g13715(.dina(n13782), .dinb(n13777), .dout(n13783));
  jxor g13716(.dina(n13783), .dinb(n5277), .dout(n13784));
  jor  g13717(.dina(n13784), .dinb(n13776), .dout(n13785));
  jxor g13718(.dina(n12951), .dinb(n12950), .dout(n13786));
  jand g13719(.dina(n10307), .dinb(n5280), .dout(n13787));
  jand g13720(.dina(n10305), .dinb(n5814), .dout(n13788));
  jand g13721(.dina(n9872), .dinb(n5531), .dout(n13789));
  jand g13722(.dina(n9655), .dinb(n5536), .dout(n13790));
  jor  g13723(.dina(n13790), .dinb(n13789), .dout(n13791));
  jor  g13724(.dina(n13791), .dinb(n13788), .dout(n13792));
  jor  g13725(.dina(n13792), .dinb(n13787), .dout(n13793));
  jxor g13726(.dina(n13793), .dinb(\a[5] ), .dout(n13794));
  jand g13727(.dina(n13794), .dinb(n13786), .dout(n13795));
  jnot g13728(.din(n13795), .dout(n13796));
  jxor g13729(.dina(n12946), .dinb(n12945), .dout(n13797));
  jnot g13730(.din(n13797), .dout(n13798));
  jand g13731(.dina(n9874), .dinb(n5280), .dout(n13799));
  jand g13732(.dina(n9655), .dinb(n5531), .dout(n13800));
  jand g13733(.dina(n9872), .dinb(n5814), .dout(n13801));
  jor  g13734(.dina(n13801), .dinb(n13800), .dout(n13802));
  jand g13735(.dina(n9656), .dinb(n5536), .dout(n13803));
  jor  g13736(.dina(n13803), .dinb(n13802), .dout(n13804));
  jor  g13737(.dina(n13804), .dinb(n13799), .dout(n13805));
  jxor g13738(.dina(n13805), .dinb(n5277), .dout(n13806));
  jor  g13739(.dina(n13806), .dinb(n13798), .dout(n13807));
  jxor g13740(.dina(n12941), .dinb(n12940), .dout(n13808));
  jnot g13741(.din(n13808), .dout(n13809));
  jand g13742(.dina(n9886), .dinb(n5280), .dout(n13810));
  jand g13743(.dina(n9655), .dinb(n5814), .dout(n13811));
  jand g13744(.dina(n9656), .dinb(n5531), .dout(n13812));
  jand g13745(.dina(n9250), .dinb(n5536), .dout(n13813));
  jor  g13746(.dina(n13813), .dinb(n13812), .dout(n13814));
  jor  g13747(.dina(n13814), .dinb(n13811), .dout(n13815));
  jor  g13748(.dina(n13815), .dinb(n13810), .dout(n13816));
  jxor g13749(.dina(n13816), .dinb(n5277), .dout(n13817));
  jor  g13750(.dina(n13817), .dinb(n13809), .dout(n13818));
  jxor g13751(.dina(n12936), .dinb(n12935), .dout(n13819));
  jnot g13752(.din(n13819), .dout(n13820));
  jand g13753(.dina(n9898), .dinb(n5280), .dout(n13821));
  jand g13754(.dina(n9250), .dinb(n5531), .dout(n13822));
  jand g13755(.dina(n9656), .dinb(n5814), .dout(n13823));
  jor  g13756(.dina(n13823), .dinb(n13822), .dout(n13824));
  jand g13757(.dina(n8936), .dinb(n5536), .dout(n13825));
  jor  g13758(.dina(n13825), .dinb(n13824), .dout(n13826));
  jor  g13759(.dina(n13826), .dinb(n13821), .dout(n13827));
  jxor g13760(.dina(n13827), .dinb(n5277), .dout(n13828));
  jor  g13761(.dina(n13828), .dinb(n13820), .dout(n13829));
  jxor g13762(.dina(n12933), .dinb(n12932), .dout(n13830));
  jnot g13763(.din(n13830), .dout(n13831));
  jand g13764(.dina(n9252), .dinb(n5280), .dout(n13832));
  jand g13765(.dina(n9250), .dinb(n5814), .dout(n13833));
  jand g13766(.dina(n8936), .dinb(n5531), .dout(n13834));
  jand g13767(.dina(n8723), .dinb(n5536), .dout(n13835));
  jor  g13768(.dina(n13835), .dinb(n13834), .dout(n13836));
  jor  g13769(.dina(n13836), .dinb(n13833), .dout(n13837));
  jor  g13770(.dina(n13837), .dinb(n13832), .dout(n13838));
  jxor g13771(.dina(n13838), .dinb(n5277), .dout(n13839));
  jor  g13772(.dina(n13839), .dinb(n13831), .dout(n13840));
  jxor g13773(.dina(n12928), .dinb(n12927), .dout(n13841));
  jnot g13774(.din(n13841), .dout(n13842));
  jand g13775(.dina(n8938), .dinb(n5280), .dout(n13843));
  jand g13776(.dina(n8723), .dinb(n5531), .dout(n13844));
  jand g13777(.dina(n8936), .dinb(n5814), .dout(n13845));
  jor  g13778(.dina(n13845), .dinb(n13844), .dout(n13846));
  jand g13779(.dina(n8740), .dinb(n5536), .dout(n13847));
  jor  g13780(.dina(n13847), .dinb(n13846), .dout(n13848));
  jor  g13781(.dina(n13848), .dinb(n13843), .dout(n13849));
  jxor g13782(.dina(n13849), .dinb(n5277), .dout(n13850));
  jor  g13783(.dina(n13850), .dinb(n13842), .dout(n13851));
  jxor g13784(.dina(n12924), .dinb(n12916), .dout(n13852));
  jnot g13785(.din(n13852), .dout(n13853));
  jand g13786(.dina(n8950), .dinb(n5280), .dout(n13854));
  jand g13787(.dina(n8740), .dinb(n5531), .dout(n13855));
  jand g13788(.dina(n8723), .dinb(n5814), .dout(n13856));
  jor  g13789(.dina(n13856), .dinb(n13855), .dout(n13857));
  jand g13790(.dina(n8268), .dinb(n5536), .dout(n13858));
  jor  g13791(.dina(n13858), .dinb(n13857), .dout(n13859));
  jor  g13792(.dina(n13859), .dinb(n13854), .dout(n13860));
  jxor g13793(.dina(n13860), .dinb(n5277), .dout(n13861));
  jor  g13794(.dina(n13861), .dinb(n13853), .dout(n13862));
  jand g13795(.dina(n8962), .dinb(n5280), .dout(n13863));
  jand g13796(.dina(n8740), .dinb(n5814), .dout(n13864));
  jand g13797(.dina(n8268), .dinb(n5531), .dout(n13865));
  jand g13798(.dina(n8022), .dinb(n5536), .dout(n13866));
  jor  g13799(.dina(n13866), .dinb(n13865), .dout(n13867));
  jor  g13800(.dina(n13867), .dinb(n13864), .dout(n13868));
  jor  g13801(.dina(n13868), .dinb(n13863), .dout(n13869));
  jxor g13802(.dina(n13869), .dinb(n5277), .dout(n13870));
  jnot g13803(.din(n13870), .dout(n13871));
  jor  g13804(.dina(n12903), .dinb(n4713), .dout(n13872));
  jxor g13805(.dina(n13872), .dinb(n12911), .dout(n13873));
  jand g13806(.dina(n13873), .dinb(n13871), .dout(n13874));
  jand g13807(.dina(n12900), .dinb(\a[8] ), .dout(n13875));
  jxor g13808(.dina(n13875), .dinb(n12898), .dout(n13876));
  jnot g13809(.din(n13876), .dout(n13877));
  jand g13810(.dina(n8270), .dinb(n5280), .dout(n13878));
  jand g13811(.dina(n8022), .dinb(n5531), .dout(n13879));
  jand g13812(.dina(n8268), .dinb(n5814), .dout(n13880));
  jor  g13813(.dina(n13880), .dinb(n13879), .dout(n13881));
  jand g13814(.dina(n7692), .dinb(n5536), .dout(n13882));
  jor  g13815(.dina(n13882), .dinb(n13881), .dout(n13883));
  jor  g13816(.dina(n13883), .dinb(n13878), .dout(n13884));
  jxor g13817(.dina(n13884), .dinb(n5277), .dout(n13885));
  jor  g13818(.dina(n13885), .dinb(n13877), .dout(n13886));
  jand g13819(.dina(n7315), .dinb(n5280), .dout(n13887));
  jand g13820(.dina(n7019), .dinb(n5531), .dout(n13888));
  jand g13821(.dina(n7313), .dinb(n5814), .dout(n13889));
  jor  g13822(.dina(n13889), .dinb(n13888), .dout(n13890));
  jor  g13823(.dina(n13890), .dinb(n13887), .dout(n13891));
  jnot g13824(.din(n13891), .dout(n13892));
  jand g13825(.dina(n7019), .dinb(n5279), .dout(n13893));
  jnot g13826(.din(n13893), .dout(n13894));
  jand g13827(.dina(n13894), .dinb(\a[5] ), .dout(n13895));
  jand g13828(.dina(n13895), .dinb(n13892), .dout(n13896));
  jand g13829(.dina(n7693), .dinb(n5280), .dout(n13897));
  jand g13830(.dina(n7313), .dinb(n5531), .dout(n13898));
  jand g13831(.dina(n7692), .dinb(n5814), .dout(n13899));
  jor  g13832(.dina(n13899), .dinb(n13898), .dout(n13900));
  jand g13833(.dina(n7019), .dinb(n5536), .dout(n13901));
  jor  g13834(.dina(n13901), .dinb(n13900), .dout(n13902));
  jor  g13835(.dina(n13902), .dinb(n13897), .dout(n13903));
  jnot g13836(.din(n13903), .dout(n13904));
  jand g13837(.dina(n13904), .dinb(n13896), .dout(n13905));
  jand g13838(.dina(n13905), .dinb(n12900), .dout(n13906));
  jnot g13839(.din(n13906), .dout(n13907));
  jxor g13840(.dina(n13905), .dinb(n12900), .dout(n13908));
  jnot g13841(.din(n13908), .dout(n13909));
  jand g13842(.dina(n8029), .dinb(n5280), .dout(n13910));
  jand g13843(.dina(n7692), .dinb(n5531), .dout(n13911));
  jand g13844(.dina(n8022), .dinb(n5814), .dout(n13912));
  jor  g13845(.dina(n13912), .dinb(n13911), .dout(n13913));
  jand g13846(.dina(n7313), .dinb(n5536), .dout(n13914));
  jor  g13847(.dina(n13914), .dinb(n13913), .dout(n13915));
  jor  g13848(.dina(n13915), .dinb(n13910), .dout(n13916));
  jxor g13849(.dina(n13916), .dinb(n5277), .dout(n13917));
  jor  g13850(.dina(n13917), .dinb(n13909), .dout(n13918));
  jand g13851(.dina(n13918), .dinb(n13907), .dout(n13919));
  jnot g13852(.din(n13919), .dout(n13920));
  jxor g13853(.dina(n13885), .dinb(n13877), .dout(n13921));
  jand g13854(.dina(n13921), .dinb(n13920), .dout(n13922));
  jnot g13855(.din(n13922), .dout(n13923));
  jand g13856(.dina(n13923), .dinb(n13886), .dout(n13924));
  jnot g13857(.din(n13924), .dout(n13925));
  jxor g13858(.dina(n13873), .dinb(n13871), .dout(n13926));
  jand g13859(.dina(n13926), .dinb(n13925), .dout(n13927));
  jor  g13860(.dina(n13927), .dinb(n13874), .dout(n13928));
  jxor g13861(.dina(n13861), .dinb(n13853), .dout(n13929));
  jand g13862(.dina(n13929), .dinb(n13928), .dout(n13930));
  jnot g13863(.din(n13930), .dout(n13931));
  jand g13864(.dina(n13931), .dinb(n13862), .dout(n13932));
  jnot g13865(.din(n13932), .dout(n13933));
  jxor g13866(.dina(n13850), .dinb(n13842), .dout(n13934));
  jand g13867(.dina(n13934), .dinb(n13933), .dout(n13935));
  jnot g13868(.din(n13935), .dout(n13936));
  jand g13869(.dina(n13936), .dinb(n13851), .dout(n13937));
  jxor g13870(.dina(n13839), .dinb(n13831), .dout(n13938));
  jnot g13871(.din(n13938), .dout(n13939));
  jor  g13872(.dina(n13939), .dinb(n13937), .dout(n13940));
  jand g13873(.dina(n13940), .dinb(n13840), .dout(n13941));
  jxor g13874(.dina(n13828), .dinb(n13820), .dout(n13942));
  jnot g13875(.din(n13942), .dout(n13943));
  jor  g13876(.dina(n13943), .dinb(n13941), .dout(n13944));
  jand g13877(.dina(n13944), .dinb(n13829), .dout(n13945));
  jxor g13878(.dina(n13817), .dinb(n13809), .dout(n13946));
  jnot g13879(.din(n13946), .dout(n13947));
  jor  g13880(.dina(n13947), .dinb(n13945), .dout(n13948));
  jand g13881(.dina(n13948), .dinb(n13818), .dout(n13949));
  jxor g13882(.dina(n13806), .dinb(n13798), .dout(n13950));
  jnot g13883(.din(n13950), .dout(n13951));
  jor  g13884(.dina(n13951), .dinb(n13949), .dout(n13952));
  jand g13885(.dina(n13952), .dinb(n13807), .dout(n13953));
  jxor g13886(.dina(n13794), .dinb(n13786), .dout(n13954));
  jnot g13887(.din(n13954), .dout(n13955));
  jor  g13888(.dina(n13955), .dinb(n13953), .dout(n13956));
  jand g13889(.dina(n13956), .dinb(n13796), .dout(n13957));
  jxor g13890(.dina(n13784), .dinb(n13775), .dout(n13958));
  jor  g13891(.dina(n13958), .dinb(n13957), .dout(n13959));
  jand g13892(.dina(n13959), .dinb(n13785), .dout(n13960));
  jxor g13893(.dina(n13773), .dinb(n13764), .dout(n13961));
  jor  g13894(.dina(n13961), .dinb(n13960), .dout(n13962));
  jand g13895(.dina(n13962), .dinb(n13774), .dout(n13963));
  jxor g13896(.dina(n13762), .dinb(n13753), .dout(n13964));
  jor  g13897(.dina(n13964), .dinb(n13963), .dout(n13965));
  jand g13898(.dina(n13965), .dinb(n13763), .dout(n13966));
  jxor g13899(.dina(n13751), .dinb(n13742), .dout(n13967));
  jor  g13900(.dina(n13967), .dinb(n13966), .dout(n13968));
  jand g13901(.dina(n13968), .dinb(n13752), .dout(n13969));
  jxor g13902(.dina(n13740), .dinb(n13731), .dout(n13970));
  jor  g13903(.dina(n13970), .dinb(n13969), .dout(n13971));
  jnot g13904(.din(n13971), .dout(n13972));
  jor  g13905(.dina(n13972), .dinb(n13741), .dout(n13973));
  jxor g13906(.dina(n13728), .dinb(n13720), .dout(n13974));
  jand g13907(.dina(n13974), .dinb(n13973), .dout(n13975));
  jor  g13908(.dina(n13975), .dinb(n13730), .dout(n13976));
  jxor g13909(.dina(n13716), .dinb(n13708), .dout(n13977));
  jand g13910(.dina(n13977), .dinb(n13976), .dout(n13978));
  jor  g13911(.dina(n13978), .dinb(n13718), .dout(n13979));
  jxor g13912(.dina(n13704), .dinb(n13696), .dout(n13980));
  jand g13913(.dina(n13980), .dinb(n13979), .dout(n13981));
  jor  g13914(.dina(n13981), .dinb(n13706), .dout(n13982));
  jxor g13915(.dina(n13692), .dinb(n13684), .dout(n13983));
  jand g13916(.dina(n13983), .dinb(n13982), .dout(n13984));
  jor  g13917(.dina(n13984), .dinb(n13694), .dout(n13985));
  jxor g13918(.dina(n13680), .dinb(n13672), .dout(n13986));
  jand g13919(.dina(n13986), .dinb(n13985), .dout(n13987));
  jor  g13920(.dina(n13987), .dinb(n13682), .dout(n13988));
  jxor g13921(.dina(n13669), .dinb(n13661), .dout(n13989));
  jand g13922(.dina(n13989), .dinb(n13988), .dout(n13990));
  jor  g13923(.dina(n13990), .dinb(n13670), .dout(n13991));
  jxor g13924(.dina(n13658), .dinb(n13650), .dout(n13992));
  jand g13925(.dina(n13992), .dinb(n13991), .dout(n13993));
  jor  g13926(.dina(n13993), .dinb(n13660), .dout(n13994));
  jxor g13927(.dina(n13647), .dinb(n13638), .dout(n13995));
  jand g13928(.dina(n13995), .dinb(n13994), .dout(n13996));
  jor  g13929(.dina(n13996), .dinb(n13649), .dout(n13997));
  jxor g13930(.dina(n13635), .dinb(n13626), .dout(n13998));
  jand g13931(.dina(n13998), .dinb(n13997), .dout(n13999));
  jor  g13932(.dina(n13999), .dinb(n13637), .dout(n14000));
  jnot g13933(.din(n14000), .dout(n14001));
  jxor g13934(.dina(n13624), .dinb(n13261), .dout(n14002));
  jor  g13935(.dina(n14002), .dinb(n14001), .dout(n14003));
  jand g13936(.dina(n14003), .dinb(n13625), .dout(n14004));
  jnot g13937(.din(n13108), .dout(n14005));
  jor  g13938(.dina(n13258), .dinb(n14005), .dout(n14006));
  jnot g13939(.din(n14006), .dout(n14007));
  jand g13940(.dina(n13260), .dinb(n13005), .dout(n14008));
  jor  g13941(.dina(n14008), .dinb(n14007), .dout(n14009));
  jnot g13942(.din(n13098), .dout(n14010));
  jor  g13943(.dina(n13106), .dinb(n14010), .dout(n14011));
  jor  g13944(.dina(n13107), .dinb(n13009), .dout(n14012));
  jand g13945(.dina(n14012), .dinb(n14011), .dout(n14013));
  jor  g13946(.dina(n13096), .dinb(n13088), .dout(n14014));
  jnot g13947(.din(n14014), .dout(n14015));
  jand g13948(.dina(n13097), .dinb(n13014), .dout(n14016));
  jor  g13949(.dina(n14016), .dinb(n14015), .dout(n14017));
  jor  g13950(.dina(n13085), .dinb(n13077), .dout(n14018));
  jand g13951(.dina(n13086), .dinb(n13019), .dout(n14019));
  jnot g13952(.din(n14019), .dout(n14020));
  jand g13953(.dina(n14020), .dinb(n14018), .dout(n14021));
  jnot g13954(.din(n14021), .dout(n14022));
  jor  g13955(.dina(n13074), .dinb(n13066), .dout(n14023));
  jand g13956(.dina(n13075), .dinb(n13022), .dout(n14024));
  jnot g13957(.din(n14024), .dout(n14025));
  jand g13958(.dina(n14025), .dinb(n14023), .dout(n14026));
  jnot g13959(.din(n14026), .dout(n14027));
  jor  g13960(.dina(n13063), .dinb(n13055), .dout(n14028));
  jand g13961(.dina(n13064), .dinb(n13027), .dout(n14029));
  jnot g13962(.din(n14029), .dout(n14030));
  jand g13963(.dina(n14030), .dinb(n14028), .dout(n14031));
  jnot g13964(.din(n14031), .dout(n14032));
  jand g13965(.dina(n13052), .dinb(n13044), .dout(n14033));
  jand g13966(.dina(n13053), .dinb(n13030), .dout(n14034));
  jor  g13967(.dina(n14034), .dinb(n14033), .dout(n14035));
  jand g13968(.dina(n13033), .dinb(n13031), .dout(n14036));
  jnot g13969(.din(n14036), .dout(n14037));
  jor  g13970(.dina(n13043), .dinb(n13035), .dout(n14038));
  jand g13971(.dina(n14038), .dinb(n14037), .dout(n14039));
  jnot g13972(.din(n14039), .dout(n14040));
  jand g13973(.dina(n2337), .dinb(n645), .dout(n14041));
  jand g13974(.dina(n14041), .dinb(n7495), .dout(n14042));
  jand g13975(.dina(n14042), .dinb(n3261), .dout(n14043));
  jand g13976(.dina(n14043), .dinb(n1734), .dout(n14044));
  jand g13977(.dina(n326), .dinb(n831), .dout(n14045));
  jand g13978(.dina(n14045), .dinb(n895), .dout(n14046));
  jand g13979(.dina(n1534), .dinb(n1213), .dout(n14047));
  jand g13980(.dina(n14047), .dinb(n2521), .dout(n14048));
  jand g13981(.dina(n14048), .dinb(n14046), .dout(n14049));
  jand g13982(.dina(n14049), .dinb(n171), .dout(n14050));
  jand g13983(.dina(n1865), .dinb(n351), .dout(n14051));
  jand g13984(.dina(n14051), .dinb(n4008), .dout(n14052));
  jand g13985(.dina(n908), .dinb(n1360), .dout(n14053));
  jand g13986(.dina(n14053), .dinb(n440), .dout(n14054));
  jand g13987(.dina(n14054), .dinb(n884), .dout(n14055));
  jand g13988(.dina(n14055), .dinb(n14052), .dout(n14056));
  jand g13989(.dina(n461), .dinb(n454), .dout(n14057));
  jand g13990(.dina(n14057), .dinb(n1163), .dout(n14058));
  jand g13991(.dina(n14058), .dinb(n7230), .dout(n14059));
  jand g13992(.dina(n2600), .dinb(n1782), .dout(n14060));
  jand g13993(.dina(n14060), .dinb(n1976), .dout(n14061));
  jand g13994(.dina(n14061), .dinb(n14059), .dout(n14062));
  jand g13995(.dina(n14062), .dinb(n14056), .dout(n14063));
  jand g13996(.dina(n921), .dinb(n713), .dout(n14064));
  jand g13997(.dina(n14064), .dinb(n3150), .dout(n14065));
  jand g13998(.dina(n14065), .dinb(n1772), .dout(n14066));
  jand g13999(.dina(n14066), .dinb(n6418), .dout(n14067));
  jand g14000(.dina(n14067), .dinb(n1218), .dout(n14068));
  jand g14001(.dina(n14068), .dinb(n14063), .dout(n14069));
  jand g14002(.dina(n14069), .dinb(n14050), .dout(n14070));
  jand g14003(.dina(n445), .dinb(n465), .dout(n14071));
  jand g14004(.dina(n14071), .dinb(n493), .dout(n14072));
  jand g14005(.dina(n2364), .dinb(n2159), .dout(n14073));
  jand g14006(.dina(n6262), .dinb(n4435), .dout(n14074));
  jand g14007(.dina(n14074), .dinb(n14073), .dout(n14075));
  jand g14008(.dina(n14075), .dinb(n14072), .dout(n14076));
  jand g14009(.dina(n2024), .dinb(n542), .dout(n14077));
  jand g14010(.dina(n14077), .dinb(n14076), .dout(n14078));
  jand g14011(.dina(n14078), .dinb(n14070), .dout(n14079));
  jand g14012(.dina(n14079), .dinb(n14044), .dout(n14080));
  jnot g14013(.din(n14080), .dout(n14081));
  jand g14014(.dina(n7315), .dinb(n5076), .dout(n14082));
  jand g14015(.dina(n7313), .dinb(n5084), .dout(n14083));
  jand g14016(.dina(n7019), .dinb(n5082), .dout(n14084));
  jor  g14017(.dina(n14084), .dinb(n14083), .dout(n14085));
  jor  g14018(.dina(n14085), .dinb(n14082), .dout(n14086));
  jxor g14019(.dina(n14086), .dinb(n14081), .dout(n14087));
  jnot g14020(.din(n14087), .dout(n14088));
  jand g14021(.dina(n8270), .dinb(n2936), .dout(n14089));
  jand g14022(.dina(n8022), .dinb(n2940), .dout(n14090));
  jand g14023(.dina(n8268), .dinb(n2943), .dout(n14091));
  jor  g14024(.dina(n14091), .dinb(n14090), .dout(n14092));
  jand g14025(.dina(n7692), .dinb(n3684), .dout(n14093));
  jor  g14026(.dina(n14093), .dinb(n14092), .dout(n14094));
  jor  g14027(.dina(n14094), .dinb(n14089), .dout(n14095));
  jxor g14028(.dina(n14095), .dinb(n93), .dout(n14096));
  jxor g14029(.dina(n14096), .dinb(n14088), .dout(n14097));
  jxor g14030(.dina(n14097), .dinb(n14040), .dout(n14098));
  jnot g14031(.din(n14098), .dout(n14099));
  jand g14032(.dina(n8938), .dinb(n71), .dout(n14100));
  jand g14033(.dina(n8723), .dinb(n731), .dout(n14101));
  jand g14034(.dina(n8936), .dinb(n796), .dout(n14102));
  jor  g14035(.dina(n14102), .dinb(n14101), .dout(n14103));
  jand g14036(.dina(n8740), .dinb(n1806), .dout(n14104));
  jor  g14037(.dina(n14104), .dinb(n14103), .dout(n14105));
  jor  g14038(.dina(n14105), .dinb(n14100), .dout(n14106));
  jxor g14039(.dina(n14106), .dinb(n77), .dout(n14107));
  jxor g14040(.dina(n14107), .dinb(n14099), .dout(n14108));
  jxor g14041(.dina(n14108), .dinb(n14035), .dout(n14109));
  jnot g14042(.din(n14109), .dout(n14110));
  jand g14043(.dina(n9886), .dinb(n806), .dout(n14111));
  jand g14044(.dina(n9656), .dinb(n1612), .dout(n14112));
  jand g14045(.dina(n9655), .dinb(n1620), .dout(n14113));
  jor  g14046(.dina(n14113), .dinb(n14112), .dout(n14114));
  jand g14047(.dina(n9250), .dinb(n1644), .dout(n14115));
  jor  g14048(.dina(n14115), .dinb(n14114), .dout(n14116));
  jor  g14049(.dina(n14116), .dinb(n14111), .dout(n14117));
  jxor g14050(.dina(n14117), .dinb(n65), .dout(n14118));
  jxor g14051(.dina(n14118), .dinb(n14110), .dout(n14119));
  jxor g14052(.dina(n14119), .dinb(n14032), .dout(n14120));
  jnot g14053(.din(n14120), .dout(n14121));
  jand g14054(.dina(n10862), .dinb(n1819), .dout(n14122));
  jand g14055(.dina(n10647), .dinb(n2243), .dout(n14123));
  jand g14056(.dina(n10305), .dinb(n2180), .dout(n14124));
  jand g14057(.dina(n9872), .dinb(n2185), .dout(n14125));
  jor  g14058(.dina(n14125), .dinb(n14124), .dout(n14126));
  jor  g14059(.dina(n14126), .dinb(n14123), .dout(n14127));
  jor  g14060(.dina(n14127), .dinb(n14122), .dout(n14128));
  jxor g14061(.dina(n14128), .dinb(n2196), .dout(n14129));
  jxor g14062(.dina(n14129), .dinb(n14121), .dout(n14130));
  jxor g14063(.dina(n14130), .dinb(n14027), .dout(n14131));
  jnot g14064(.din(n14131), .dout(n14132));
  jand g14065(.dina(n11308), .dinb(n2743), .dout(n14133));
  jand g14066(.dina(n11306), .dinb(n2752), .dout(n14134));
  jand g14067(.dina(n10836), .dinb(n2748), .dout(n14135));
  jand g14068(.dina(n10640), .dinb(n2757), .dout(n14136));
  jor  g14069(.dina(n14136), .dinb(n14135), .dout(n14137));
  jor  g14070(.dina(n14137), .dinb(n14134), .dout(n14138));
  jor  g14071(.dina(n14138), .dinb(n14133), .dout(n14139));
  jxor g14072(.dina(n14139), .dinb(n2441), .dout(n14140));
  jxor g14073(.dina(n14140), .dinb(n14132), .dout(n14141));
  jxor g14074(.dina(n14141), .dinb(n14022), .dout(n14142));
  jand g14075(.dina(n11800), .dinb(n3423), .dout(n14143));
  jand g14076(.dina(n11646), .dinb(n3428), .dout(n14144));
  jand g14077(.dina(n11798), .dinb(n3569), .dout(n14145));
  jor  g14078(.dina(n14145), .dinb(n14144), .dout(n14146));
  jand g14079(.dina(n11647), .dinb(n3210), .dout(n14147));
  jor  g14080(.dina(n14147), .dinb(n14146), .dout(n14148));
  jor  g14081(.dina(n14148), .dinb(n14143), .dout(n14149));
  jxor g14082(.dina(n14149), .dinb(n3473), .dout(n14150));
  jxor g14083(.dina(n14150), .dinb(n14142), .dout(n14151));
  jxor g14084(.dina(n14151), .dinb(n14017), .dout(n14152));
  jand g14085(.dina(n12684), .dinb(n4022), .dout(n14153));
  jand g14086(.dina(n12536), .dinb(n4220), .dout(n14154));
  jand g14087(.dina(n12547), .dinb(n4027), .dout(n14155));
  jand g14088(.dina(n12282), .dinb(n3870), .dout(n14156));
  jor  g14089(.dina(n14156), .dinb(n14155), .dout(n14157));
  jor  g14090(.dina(n14157), .dinb(n14154), .dout(n14158));
  jor  g14091(.dina(n14158), .dinb(n14153), .dout(n14159));
  jxor g14092(.dina(n14159), .dinb(\a[11] ), .dout(n14160));
  jxor g14093(.dina(n14160), .dinb(n14152), .dout(n14161));
  jxor g14094(.dina(n14161), .dinb(n14013), .dout(n14162));
  jand g14095(.dina(n13639), .dinb(n4691), .dout(n14163));
  jand g14096(.dina(n13478), .dinb(n4941), .dout(n14164));
  jand g14097(.dina(n13248), .dinb(n4696), .dout(n14165));
  jand g14098(.dina(n12669), .dinb(n4701), .dout(n14166));
  jor  g14099(.dina(n14166), .dinb(n14165), .dout(n14167));
  jor  g14100(.dina(n14167), .dinb(n14164), .dout(n14168));
  jor  g14101(.dina(n14168), .dinb(n14163), .dout(n14169));
  jxor g14102(.dina(n14169), .dinb(n4713), .dout(n14170));
  jxor g14103(.dina(n14170), .dinb(n14162), .dout(n14171));
  jnot g14104(.din(n14171), .dout(n14172));
  jxor g14105(.dina(n14172), .dinb(n14009), .dout(n14173));
  jand g14106(.dina(n13614), .dinb(n13469), .dout(n14174));
  jand g14107(.dina(n13615), .dinb(n13489), .dout(n14175));
  jor  g14108(.dina(n14175), .dinb(n14174), .dout(n14176));
  jand g14109(.dina(n13612), .dinb(n13499), .dout(n14177));
  jand g14110(.dina(n13613), .dinb(n13494), .dout(n14178));
  jor  g14111(.dina(n14178), .dinb(n14177), .dout(n14179));
  jor  g14112(.dina(n13610), .dinb(n13602), .dout(n14180));
  jand g14113(.dina(n13611), .dinb(n13598), .dout(n14181));
  jnot g14114(.din(n14181), .dout(n14182));
  jand g14115(.dina(n14182), .dinb(n14180), .dout(n14183));
  jnot g14116(.din(n14183), .dout(n14184));
  jand g14117(.dina(n13588), .dinb(n13502), .dout(n14185));
  jand g14118(.dina(n13597), .dinb(n13589), .dout(n14186));
  jor  g14119(.dina(n14186), .dinb(n14185), .dout(n14187));
  jor  g14120(.dina(n13586), .dinb(n13578), .dout(n14188));
  jand g14121(.dina(n13587), .dinb(n13505), .dout(n14189));
  jnot g14122(.din(n14189), .dout(n14190));
  jand g14123(.dina(n14190), .dinb(n14188), .dout(n14191));
  jnot g14124(.din(n14191), .dout(n14192));
  jor  g14125(.dina(n6516), .dinb(n7061), .dout(n14193));
  jand g14126(.dina(n6050), .dinb(n6140), .dout(n14194));
  jand g14127(.dina(n6391), .dinb(n5084), .dout(n14195));
  jor  g14128(.dina(n14195), .dinb(n14194), .dout(n14196));
  jand g14129(.dina(n6394), .dinb(n5082), .dout(n14197));
  jor  g14130(.dina(n14197), .dinb(n14196), .dout(n14198));
  jnot g14131(.din(n14198), .dout(n14199));
  jand g14132(.dina(n14199), .dinb(n14193), .dout(n14200));
  jnot g14133(.din(n14200), .dout(n14201));
  jand g14134(.dina(n2135), .dinb(n510), .dout(n14202));
  jand g14135(.dina(n14202), .dinb(n1273), .dout(n14203));
  jand g14136(.dina(n551), .dinb(n1040), .dout(n14204));
  jand g14137(.dina(n14204), .dinb(n2442), .dout(n14205));
  jand g14138(.dina(n14205), .dinb(n14203), .dout(n14206));
  jand g14139(.dina(n14206), .dinb(n8834), .dout(n14207));
  jand g14140(.dina(n14207), .dinb(n9378), .dout(n14208));
  jand g14141(.dina(n8580), .dinb(n2042), .dout(n14209));
  jand g14142(.dina(n1915), .dinb(n1376), .dout(n14210));
  jand g14143(.dina(n14210), .dinb(n14209), .dout(n14211));
  jand g14144(.dina(n2410), .dinb(n1596), .dout(n14212));
  jand g14145(.dina(n14212), .dinb(n1169), .dout(n14213));
  jand g14146(.dina(n14213), .dinb(n14211), .dout(n14214));
  jand g14147(.dina(n2148), .dinb(n82), .dout(n14215));
  jand g14148(.dina(n1346), .dinb(n463), .dout(n14216));
  jand g14149(.dina(n14216), .dinb(n14215), .dout(n14217));
  jand g14150(.dina(n887), .dinb(n266), .dout(n14218));
  jand g14151(.dina(n534), .dinb(n1304), .dout(n14219));
  jand g14152(.dina(n14219), .dinb(n325), .dout(n14220));
  jand g14153(.dina(n14220), .dinb(n14218), .dout(n14221));
  jand g14154(.dina(n14221), .dinb(n14217), .dout(n14222));
  jand g14155(.dina(n14222), .dinb(n14214), .dout(n14223));
  jand g14156(.dina(n14223), .dinb(n3342), .dout(n14224));
  jand g14157(.dina(n14224), .dinb(n14208), .dout(n14225));
  jnot g14158(.din(n14225), .dout(n14226));
  jxor g14159(.dina(n14226), .dinb(n13575), .dout(n14227));
  jxor g14160(.dina(n14227), .dinb(n14201), .dout(n14228));
  jxor g14161(.dina(n14228), .dinb(n14192), .dout(n14229));
  jor  g14162(.dina(n7303), .dinb(n4343), .dout(n14230));
  jor  g14163(.dina(n7301), .dinb(n4348), .dout(n14231));
  jor  g14164(.dina(n6297), .dinb(n3683), .dout(n14232));
  jor  g14165(.dina(n6489), .dinb(n4346), .dout(n14233));
  jand g14166(.dina(n14233), .dinb(n14232), .dout(n14234));
  jand g14167(.dina(n14234), .dinb(n14231), .dout(n14235));
  jand g14168(.dina(n14235), .dinb(n14230), .dout(n14236));
  jxor g14169(.dina(n14236), .dinb(n93), .dout(n14237));
  jxor g14170(.dina(n14237), .dinb(n14229), .dout(n14238));
  jxor g14171(.dina(n14238), .dinb(n14187), .dout(n14239));
  jnot g14172(.din(n14239), .dout(n14240));
  jor  g14173(.dina(n8260), .dinb(n2303), .dout(n14241));
  jor  g14174(.dina(n7680), .dinb(n1805), .dout(n14242));
  jor  g14175(.dina(n7999), .dinb(n2306), .dout(n14243));
  jand g14176(.dina(n14243), .dinb(n14242), .dout(n14244));
  jand g14177(.dina(n14244), .dinb(n14241), .dout(n14245));
  jxor g14178(.dina(n14245), .dinb(\a[26] ), .dout(n14246));
  jxor g14179(.dina(n14246), .dinb(n14240), .dout(n14247));
  jxor g14180(.dina(n14247), .dinb(n14184), .dout(n14248));
  jxor g14181(.dina(n14248), .dinb(n14179), .dout(n14249));
  jxor g14182(.dina(n14249), .dinb(n13614), .dout(n14250));
  jxor g14183(.dina(n14250), .dinb(n14176), .dout(n14251));
  jand g14184(.dina(n14251), .dinb(n5280), .dout(n14252));
  jand g14185(.dina(n13614), .dinb(n5531), .dout(n14253));
  jand g14186(.dina(n14249), .dinb(n5814), .dout(n14254));
  jor  g14187(.dina(n14254), .dinb(n14253), .dout(n14255));
  jand g14188(.dina(n13469), .dinb(n5536), .dout(n14256));
  jor  g14189(.dina(n14256), .dinb(n14255), .dout(n14257));
  jor  g14190(.dina(n14257), .dinb(n14252), .dout(n14258));
  jxor g14191(.dina(n14258), .dinb(n5277), .dout(n14259));
  jxor g14192(.dina(n14259), .dinb(n14173), .dout(n14260));
  jxor g14193(.dina(n14260), .dinb(n14004), .dout(n14261));
  jnot g14194(.din(n14261), .dout(n14262));
  jand g14195(.dina(n14238), .dinb(n14187), .dout(n14263));
  jnot g14196(.din(n14263), .dout(n14264));
  jor  g14197(.dina(n14246), .dinb(n14240), .dout(n14265));
  jand g14198(.dina(n14265), .dinb(n14264), .dout(n14266));
  jnot g14199(.din(n14266), .dout(n14267));
  jnot g14200(.din(n13575), .dout(n14268));
  jand g14201(.dina(n14225), .dinb(n14268), .dout(n14269));
  jand g14202(.dina(n14227), .dinb(n14201), .dout(n14270));
  jor  g14203(.dina(n14270), .dinb(n14269), .dout(n14271));
  jor  g14204(.dina(n6999), .dinb(n7061), .dout(n14272));
  jand g14205(.dina(n6394), .dinb(n6050), .dout(n14273));
  jand g14206(.dina(n6298), .dinb(n5084), .dout(n14274));
  jor  g14207(.dina(n14274), .dinb(n14273), .dout(n14275));
  jand g14208(.dina(n6391), .dinb(n5082), .dout(n14276));
  jor  g14209(.dina(n14276), .dinb(n14275), .dout(n14277));
  jnot g14210(.din(n14277), .dout(n14278));
  jand g14211(.dina(n14278), .dinb(n14272), .dout(n14279));
  jnot g14212(.din(n14279), .dout(n14280));
  jand g14213(.dina(n1099), .dinb(n548), .dout(n14281));
  jand g14214(.dina(n495), .dinb(n1351), .dout(n14282));
  jand g14215(.dina(n14282), .dinb(n1233), .dout(n14283));
  jand g14216(.dina(n14283), .dinb(n14281), .dout(n14284));
  jand g14217(.dina(n1325), .dinb(n1238), .dout(n14285));
  jand g14218(.dina(n14285), .dinb(n1315), .dout(n14286));
  jand g14219(.dina(n14286), .dinb(n1169), .dout(n14287));
  jand g14220(.dina(n9720), .dinb(n1218), .dout(n14288));
  jand g14221(.dina(n14288), .dinb(n14287), .dout(n14289));
  jand g14222(.dina(n14289), .dinb(n14284), .dout(n14290));
  jand g14223(.dina(n14290), .dinb(n4628), .dout(n14291));
  jand g14224(.dina(n685), .dinb(n880), .dout(n14292));
  jand g14225(.dina(n14292), .dinb(n1427), .dout(n14293));
  jand g14226(.dina(n14293), .dinb(n9344), .dout(n14294));
  jand g14227(.dina(n14294), .dinb(n5241), .dout(n14295));
  jand g14228(.dina(n2023), .dinb(n521), .dout(n14296));
  jand g14229(.dina(n14296), .dinb(n1516), .dout(n14297));
  jand g14230(.dina(n1163), .dinb(n535), .dout(n14298));
  jand g14231(.dina(n14298), .dinb(n14297), .dout(n14299));
  jand g14232(.dina(n14299), .dinb(n4417), .dout(n14300));
  jand g14233(.dina(n14300), .dinb(n14295), .dout(n14301));
  jand g14234(.dina(n442), .dinb(n135), .dout(n14302));
  jand g14235(.dina(n14302), .dinb(n1835), .dout(n14303));
  jand g14236(.dina(n808), .dinb(n920), .dout(n14304));
  jand g14237(.dina(n14304), .dinb(n14303), .dout(n14305));
  jand g14238(.dina(n1037), .dinb(n826), .dout(n14306));
  jand g14239(.dina(n14306), .dinb(n14305), .dout(n14307));
  jand g14240(.dina(n452), .dinb(n713), .dout(n14308));
  jand g14241(.dina(n14308), .dinb(n8593), .dout(n14309));
  jand g14242(.dina(n14309), .dinb(n6292), .dout(n14310));
  jand g14243(.dina(n1005), .dinb(n838), .dout(n14311));
  jand g14244(.dina(n14311), .dinb(n672), .dout(n14312));
  jand g14245(.dina(n1867), .dinb(n168), .dout(n14313));
  jand g14246(.dina(n14313), .dinb(n583), .dout(n14314));
  jand g14247(.dina(n14314), .dinb(n14312), .dout(n14315));
  jand g14248(.dina(n14315), .dinb(n14310), .dout(n14316));
  jand g14249(.dina(n14316), .dinb(n14307), .dout(n14317));
  jand g14250(.dina(n3320), .dinb(n326), .dout(n14318));
  jand g14251(.dina(n14318), .dinb(n11363), .dout(n14319));
  jand g14252(.dina(n14319), .dinb(n14317), .dout(n14320));
  jand g14253(.dina(n14320), .dinb(n14301), .dout(n14321));
  jand g14254(.dina(n1779), .dinb(n1168), .dout(n14322));
  jand g14255(.dina(n1207), .dinb(n884), .dout(n14323));
  jand g14256(.dina(n14323), .dinb(n3397), .dout(n14324));
  jand g14257(.dina(n14324), .dinb(n14322), .dout(n14325));
  jand g14258(.dina(n907), .dinb(n517), .dout(n14326));
  jand g14259(.dina(n14326), .dinb(n553), .dout(n14327));
  jand g14260(.dina(n14327), .dinb(n11707), .dout(n14328));
  jand g14261(.dina(n14328), .dinb(n14325), .dout(n14329));
  jand g14262(.dina(n1743), .dinb(n1367), .dout(n14330));
  jand g14263(.dina(n14330), .dinb(n8589), .dout(n14331));
  jand g14264(.dina(n14331), .dinb(n3978), .dout(n14332));
  jand g14265(.dina(n14332), .dinb(n14329), .dout(n14333));
  jand g14266(.dina(n14333), .dinb(n14321), .dout(n14334));
  jand g14267(.dina(n14334), .dinb(n14291), .dout(n14335));
  jxor g14268(.dina(n14335), .dinb(n14226), .dout(n14336));
  jxor g14269(.dina(n14336), .dinb(n14280), .dout(n14337));
  jxor g14270(.dina(n14337), .dinb(n14271), .dout(n14338));
  jand g14271(.dina(n14228), .dinb(n14192), .dout(n14339));
  jand g14272(.dina(n14237), .dinb(n14229), .dout(n14340));
  jor  g14273(.dina(n14340), .dinb(n14339), .dout(n14341));
  jxor g14274(.dina(n14341), .dinb(n14338), .dout(n14342));
  jor  g14275(.dina(n7999), .dinb(n1805), .dout(n14343));
  jor  g14276(.dina(n8295), .dinb(n2303), .dout(n14344));
  jand g14277(.dina(n14344), .dinb(n14343), .dout(n14345));
  jxor g14278(.dina(n14345), .dinb(\a[26] ), .dout(n14346));
  jor  g14279(.dina(n7682), .dinb(n4343), .dout(n14347));
  jor  g14280(.dina(n7301), .dinb(n4346), .dout(n14348));
  jor  g14281(.dina(n7680), .dinb(n4348), .dout(n14349));
  jand g14282(.dina(n14349), .dinb(n14348), .dout(n14350));
  jor  g14283(.dina(n6489), .dinb(n3683), .dout(n14351));
  jand g14284(.dina(n14351), .dinb(n14350), .dout(n14352));
  jand g14285(.dina(n14352), .dinb(n14347), .dout(n14353));
  jxor g14286(.dina(n14353), .dinb(\a[29] ), .dout(n14354));
  jxor g14287(.dina(n14354), .dinb(n14346), .dout(n14355));
  jxor g14288(.dina(n14355), .dinb(n14342), .dout(n14356));
  jand g14289(.dina(n14356), .dinb(n14267), .dout(n14357));
  jand g14290(.dina(n14247), .dinb(n14184), .dout(n14358));
  jand g14291(.dina(n14248), .dinb(n14179), .dout(n14359));
  jor  g14292(.dina(n14359), .dinb(n14358), .dout(n14360));
  jxor g14293(.dina(n14356), .dinb(n14267), .dout(n14361));
  jand g14294(.dina(n14361), .dinb(n14360), .dout(n14362));
  jor  g14295(.dina(n14362), .dinb(n14357), .dout(n14363));
  jor  g14296(.dina(n14354), .dinb(n14346), .dout(n14364));
  jand g14297(.dina(n14355), .dinb(n14342), .dout(n14365));
  jnot g14298(.din(n14365), .dout(n14366));
  jand g14299(.dina(n14366), .dinb(n14364), .dout(n14367));
  jnot g14300(.din(n14367), .dout(n14368));
  jand g14301(.dina(n14337), .dinb(n14271), .dout(n14369));
  jand g14302(.dina(n14341), .dinb(n14338), .dout(n14370));
  jor  g14303(.dina(n14370), .dinb(n14369), .dout(n14371));
  jor  g14304(.dina(n6491), .dinb(n7061), .dout(n14372));
  jand g14305(.dina(n6391), .dinb(n6050), .dout(n14373));
  jand g14306(.dina(n7218), .dinb(n5084), .dout(n14374));
  jor  g14307(.dina(n14374), .dinb(n14373), .dout(n14375));
  jand g14308(.dina(n6298), .dinb(n5082), .dout(n14376));
  jor  g14309(.dina(n14376), .dinb(n14375), .dout(n14377));
  jnot g14310(.din(n14377), .dout(n14378));
  jand g14311(.dina(n14378), .dinb(n14372), .dout(n14379));
  jnot g14312(.din(n14379), .dout(n14380));
  jor  g14313(.dina(n14335), .dinb(n14226), .dout(n14381));
  jand g14314(.dina(n14336), .dinb(n14280), .dout(n14382));
  jnot g14315(.din(n14382), .dout(n14383));
  jand g14316(.dina(n14383), .dinb(n14381), .dout(n14384));
  jnot g14317(.din(n14384), .dout(n14385));
  jand g14318(.dina(n965), .dinb(n650), .dout(n14386));
  jand g14319(.dina(n14386), .dinb(n3827), .dout(n14387));
  jand g14320(.dina(n14387), .dinb(n9332), .dout(n14388));
  jand g14321(.dina(n4678), .dinb(n1868), .dout(n14389));
  jand g14322(.dina(n14389), .dinb(n14388), .dout(n14390));
  jand g14323(.dina(n881), .dinb(n1327), .dout(n14391));
  jand g14324(.dina(n14391), .dinb(n10191), .dout(n14392));
  jand g14325(.dina(n8589), .dinb(n6151), .dout(n14393));
  jand g14326(.dina(n14393), .dinb(n14392), .dout(n14394));
  jand g14327(.dina(n1541), .dinb(n714), .dout(n14395));
  jand g14328(.dina(n14395), .dinb(n1360), .dout(n14396));
  jand g14329(.dina(n3819), .dinb(n3758), .dout(n14397));
  jand g14330(.dina(n14397), .dinb(n14396), .dout(n14398));
  jand g14331(.dina(n14398), .dinb(n14394), .dout(n14399));
  jand g14332(.dina(n14399), .dinb(n8616), .dout(n14400));
  jand g14333(.dina(n14400), .dinb(n14390), .dout(n14401));
  jand g14334(.dina(n14066), .dinb(n886), .dout(n14402));
  jand g14335(.dina(n1511), .dinb(n430), .dout(n14403));
  jand g14336(.dina(n14403), .dinb(n873), .dout(n14404));
  jand g14337(.dina(n2993), .dinb(n1090), .dout(n14405));
  jand g14338(.dina(n14405), .dinb(n1308), .dout(n14406));
  jand g14339(.dina(n14406), .dinb(n14404), .dout(n14407));
  jand g14340(.dina(n13524), .dinb(n11371), .dout(n14408));
  jand g14341(.dina(n14408), .dinb(n14407), .dout(n14409));
  jand g14342(.dina(n5395), .dinb(n1714), .dout(n14410));
  jand g14343(.dina(n14410), .dinb(n1763), .dout(n14411));
  jand g14344(.dina(n10527), .dinb(n2477), .dout(n14412));
  jand g14345(.dina(n14412), .dinb(n1438), .dout(n14413));
  jand g14346(.dina(n14413), .dinb(n14411), .dout(n14414));
  jand g14347(.dina(n534), .dinb(n469), .dout(n14415));
  jand g14348(.dina(n14415), .dinb(n1190), .dout(n14416));
  jand g14349(.dina(n14416), .dinb(n8578), .dout(n14417));
  jand g14350(.dina(n14417), .dinb(n1522), .dout(n14418));
  jand g14351(.dina(n14418), .dinb(n14414), .dout(n14419));
  jand g14352(.dina(n14419), .dinb(n14409), .dout(n14420));
  jand g14353(.dina(n14420), .dinb(n14402), .dout(n14421));
  jand g14354(.dina(n14421), .dinb(n1300), .dout(n14422));
  jand g14355(.dina(n14422), .dinb(n14401), .dout(n14423));
  jand g14356(.dina(n14423), .dinb(n14225), .dout(n14424));
  jnot g14357(.din(n14424), .dout(n14425));
  jor  g14358(.dina(n14423), .dinb(n14225), .dout(n14426));
  jand g14359(.dina(n14426), .dinb(n77), .dout(n14427));
  jand g14360(.dina(n14427), .dinb(n14425), .dout(n14428));
  jnot g14361(.din(n14428), .dout(n14429));
  jand g14362(.dina(n14429), .dinb(n77), .dout(n14430));
  jand g14363(.dina(n14429), .dinb(n14426), .dout(n14431));
  jand g14364(.dina(n14431), .dinb(n14425), .dout(n14432));
  jor  g14365(.dina(n14432), .dinb(n14430), .dout(n14433));
  jxor g14366(.dina(n14433), .dinb(n14385), .dout(n14434));
  jxor g14367(.dina(n14434), .dinb(n14380), .dout(n14435));
  jxor g14368(.dina(n14435), .dinb(n14371), .dout(n14436));
  jor  g14369(.dina(n8002), .dinb(n4343), .dout(n14437));
  jor  g14370(.dina(n7301), .dinb(n3683), .dout(n14438));
  jor  g14371(.dina(n7999), .dinb(n4348), .dout(n14439));
  jor  g14372(.dina(n7680), .dinb(n4346), .dout(n14440));
  jand g14373(.dina(n14440), .dinb(n14439), .dout(n14441));
  jand g14374(.dina(n14441), .dinb(n14438), .dout(n14442));
  jand g14375(.dina(n14442), .dinb(n14437), .dout(n14443));
  jxor g14376(.dina(n14443), .dinb(n93), .dout(n14444));
  jxor g14377(.dina(n14444), .dinb(n14436), .dout(n14445));
  jxor g14378(.dina(n14445), .dinb(n14368), .dout(n14446));
  jxor g14379(.dina(n14446), .dinb(n14363), .dout(n14447));
  jxor g14380(.dina(n14361), .dinb(n14360), .dout(n14448));
  jand g14381(.dina(n14448), .dinb(n14447), .dout(n14449));
  jand g14382(.dina(n14448), .dinb(n14249), .dout(n14450));
  jand g14383(.dina(n14249), .dinb(n13614), .dout(n14451));
  jand g14384(.dina(n14250), .dinb(n14176), .dout(n14452));
  jor  g14385(.dina(n14452), .dinb(n14451), .dout(n14453));
  jxor g14386(.dina(n14448), .dinb(n14249), .dout(n14454));
  jand g14387(.dina(n14454), .dinb(n14453), .dout(n14455));
  jor  g14388(.dina(n14455), .dinb(n14450), .dout(n14456));
  jxor g14389(.dina(n14448), .dinb(n14447), .dout(n14457));
  jand g14390(.dina(n14457), .dinb(n14456), .dout(n14458));
  jor  g14391(.dina(n14458), .dinb(n14449), .dout(n14459));
  jand g14392(.dina(n14435), .dinb(n14371), .dout(n14460));
  jand g14393(.dina(n14444), .dinb(n14436), .dout(n14461));
  jor  g14394(.dina(n14461), .dinb(n14460), .dout(n14462));
  jand g14395(.dina(n14433), .dinb(n14385), .dout(n14463));
  jand g14396(.dina(n14434), .dinb(n14380), .dout(n14464));
  jor  g14397(.dina(n14464), .dinb(n14463), .dout(n14465));
  jor  g14398(.dina(n7303), .dinb(n7061), .dout(n14466));
  jand g14399(.dina(n7629), .dinb(n5084), .dout(n14467));
  jand g14400(.dina(n6298), .dinb(n6050), .dout(n14468));
  jor  g14401(.dina(n14468), .dinb(n14467), .dout(n14469));
  jand g14402(.dina(n7218), .dinb(n5082), .dout(n14470));
  jor  g14403(.dina(n14470), .dinb(n14469), .dout(n14471));
  jnot g14404(.din(n14471), .dout(n14472));
  jand g14405(.dina(n14472), .dinb(n14466), .dout(n14473));
  jnot g14406(.din(n14473), .dout(n14474));
  jand g14407(.dina(n5501), .dinb(n966), .dout(n14475));
  jand g14408(.dina(n14475), .dinb(n1562), .dout(n14476));
  jand g14409(.dina(n1449), .dinb(n1701), .dout(n14477));
  jand g14410(.dina(n929), .dinb(n541), .dout(n14478));
  jand g14411(.dina(n14478), .dinb(n3967), .dout(n14479));
  jand g14412(.dina(n14479), .dinb(n14477), .dout(n14480));
  jand g14413(.dina(n1541), .dinb(n320), .dout(n14481));
  jand g14414(.dina(n14481), .dinb(n843), .dout(n14482));
  jand g14415(.dina(n14482), .dinb(n14480), .dout(n14483));
  jand g14416(.dina(n14483), .dinb(n14476), .dout(n14484));
  jand g14417(.dina(n1846), .dinb(n1325), .dout(n14485));
  jand g14418(.dina(n14485), .dinb(n1257), .dout(n14486));
  jand g14419(.dina(n14486), .dinb(n3264), .dout(n14487));
  jand g14420(.dina(n7105), .dinb(n463), .dout(n14488));
  jand g14421(.dina(n14488), .dinb(n14487), .dout(n14489));
  jand g14422(.dina(n14489), .dinb(n6254), .dout(n14490));
  jand g14423(.dina(n14490), .dinb(n14484), .dout(n14491));
  jand g14424(.dina(n1732), .dinb(n349), .dout(n14492));
  jand g14425(.dina(n6335), .dinb(n3888), .dout(n14493));
  jand g14426(.dina(n834), .dinb(n638), .dout(n14494));
  jand g14427(.dina(n14494), .dinb(n3026), .dout(n14495));
  jand g14428(.dina(n14495), .dinb(n14493), .dout(n14496));
  jand g14429(.dina(n532), .dinb(n445), .dout(n14497));
  jand g14430(.dina(n14497), .dinb(n838), .dout(n14498));
  jand g14431(.dina(n14498), .dinb(n10207), .dout(n14499));
  jand g14432(.dina(n13199), .dinb(n440), .dout(n14500));
  jand g14433(.dina(n14500), .dinb(n3176), .dout(n14501));
  jand g14434(.dina(n14501), .dinb(n14499), .dout(n14502));
  jand g14435(.dina(n14502), .dinb(n14496), .dout(n14503));
  jand g14436(.dina(n14503), .dinb(n14492), .dout(n14504));
  jand g14437(.dina(n1903), .dinb(n871), .dout(n14505));
  jand g14438(.dina(n14505), .dinb(n1852), .dout(n14506));
  jand g14439(.dina(n14506), .dinb(n1310), .dout(n14507));
  jand g14440(.dina(n902), .dinb(n1591), .dout(n14508));
  jand g14441(.dina(n14508), .dinb(n9369), .dout(n14509));
  jand g14442(.dina(n14509), .dinb(n5289), .dout(n14510));
  jand g14443(.dina(n14510), .dinb(n14507), .dout(n14511));
  jand g14444(.dina(n14511), .dinb(n14504), .dout(n14512));
  jand g14445(.dina(n14512), .dinb(n11705), .dout(n14513));
  jand g14446(.dina(n14513), .dinb(n14491), .dout(n14514));
  jnot g14447(.din(n14514), .dout(n14515));
  jxor g14448(.dina(n14515), .dinb(n14431), .dout(n14516));
  jxor g14449(.dina(n14516), .dinb(n14474), .dout(n14517));
  jxor g14450(.dina(n14517), .dinb(n14465), .dout(n14518));
  jnot g14451(.din(n14518), .dout(n14519));
  jor  g14452(.dina(n8260), .dinb(n4343), .dout(n14520));
  jor  g14453(.dina(n7680), .dinb(n3683), .dout(n14521));
  jor  g14454(.dina(n7999), .dinb(n4346), .dout(n14522));
  jand g14455(.dina(n14522), .dinb(n14521), .dout(n14523));
  jand g14456(.dina(n14523), .dinb(n14520), .dout(n14524));
  jxor g14457(.dina(n14524), .dinb(\a[29] ), .dout(n14525));
  jxor g14458(.dina(n14525), .dinb(n14519), .dout(n14526));
  jxor g14459(.dina(n14526), .dinb(n14462), .dout(n14527));
  jnot g14460(.din(n14527), .dout(n14528));
  jand g14461(.dina(n14445), .dinb(n14368), .dout(n14529));
  jnot g14462(.din(n14529), .dout(n14530));
  jnot g14463(.din(n14357), .dout(n14531));
  jnot g14464(.din(n14358), .dout(n14532));
  jnot g14465(.din(n14177), .dout(n14533));
  jnot g14466(.din(n13490), .dout(n14534));
  jor  g14467(.dina(n13468), .dinb(n13452), .dout(n14535));
  jand g14468(.dina(n14535), .dinb(n14534), .dout(n14536));
  jnot g14469(.din(n13613), .dout(n14537));
  jor  g14470(.dina(n14537), .dinb(n14536), .dout(n14538));
  jand g14471(.dina(n14538), .dinb(n14533), .dout(n14539));
  jnot g14472(.din(n14248), .dout(n14540));
  jor  g14473(.dina(n14540), .dinb(n14539), .dout(n14541));
  jand g14474(.dina(n14541), .dinb(n14532), .dout(n14542));
  jnot g14475(.din(n14361), .dout(n14543));
  jor  g14476(.dina(n14543), .dinb(n14542), .dout(n14544));
  jand g14477(.dina(n14544), .dinb(n14531), .dout(n14545));
  jnot g14478(.din(n14446), .dout(n14546));
  jor  g14479(.dina(n14546), .dinb(n14545), .dout(n14547));
  jand g14480(.dina(n14547), .dinb(n14530), .dout(n14548));
  jxor g14481(.dina(n14548), .dinb(n14528), .dout(n14549));
  jxor g14482(.dina(n14549), .dinb(n14447), .dout(n14550));
  jxor g14483(.dina(n14550), .dinb(n14459), .dout(n14551));
  jand g14484(.dina(n14551), .dinb(n6495), .dout(n14552));
  jand g14485(.dina(n14549), .dinb(n6503), .dout(n14553));
  jand g14486(.dina(n14447), .dinb(n6506), .dout(n14554));
  jand g14487(.dina(n14448), .dinb(n6500), .dout(n14555));
  jor  g14488(.dina(n14555), .dinb(n14554), .dout(n14556));
  jor  g14489(.dina(n14556), .dinb(n14553), .dout(n14557));
  jor  g14490(.dina(n14557), .dinb(n14552), .dout(n14558));
  jxor g14491(.dina(n14558), .dinb(n6219), .dout(n14559));
  jxor g14492(.dina(n14559), .dinb(n14262), .dout(n14560));
  jxor g14493(.dina(n14002), .dinb(n14001), .dout(n14561));
  jxor g14494(.dina(n14457), .dinb(n14456), .dout(n14562));
  jnot g14495(.din(n14562), .dout(n14563));
  jor  g14496(.dina(n14563), .dinb(n6496), .dout(n14564));
  jnot g14497(.din(n14447), .dout(n14565));
  jor  g14498(.dina(n14565), .dinb(n6504), .dout(n14566));
  jnot g14499(.din(n14448), .dout(n14567));
  jor  g14500(.dina(n14567), .dinb(n6507), .dout(n14568));
  jnot g14501(.din(n14249), .dout(n14569));
  jor  g14502(.dina(n14569), .dinb(n6501), .dout(n14570));
  jand g14503(.dina(n14570), .dinb(n14568), .dout(n14571));
  jand g14504(.dina(n14571), .dinb(n14566), .dout(n14572));
  jand g14505(.dina(n14572), .dinb(n14564), .dout(n14573));
  jxor g14506(.dina(n14573), .dinb(n6219), .dout(n14574));
  jand g14507(.dina(n14574), .dinb(n14561), .dout(n14575));
  jor  g14508(.dina(n14574), .dinb(n14561), .dout(n14576));
  jxor g14509(.dina(n13998), .dinb(n13997), .dout(n14577));
  jnot g14510(.din(n14577), .dout(n14578));
  jxor g14511(.dina(n14454), .dinb(n14453), .dout(n14579));
  jnot g14512(.din(n14579), .dout(n14580));
  jor  g14513(.dina(n14580), .dinb(n6496), .dout(n14581));
  jor  g14514(.dina(n14567), .dinb(n6504), .dout(n14582));
  jor  g14515(.dina(n14569), .dinb(n6507), .dout(n14583));
  jnot g14516(.din(n13614), .dout(n14584));
  jor  g14517(.dina(n14584), .dinb(n6501), .dout(n14585));
  jand g14518(.dina(n14585), .dinb(n14583), .dout(n14586));
  jand g14519(.dina(n14586), .dinb(n14582), .dout(n14587));
  jand g14520(.dina(n14587), .dinb(n14581), .dout(n14588));
  jxor g14521(.dina(n14588), .dinb(n6219), .dout(n14589));
  jnot g14522(.din(n14589), .dout(n14590));
  jand g14523(.dina(n14590), .dinb(n14578), .dout(n14591));
  jnot g14524(.din(n14591), .dout(n14592));
  jxor g14525(.dina(n13992), .dinb(n13991), .dout(n14593));
  jnot g14526(.din(n14593), .dout(n14594));
  jxor g14527(.dina(n13989), .dinb(n13988), .dout(n14595));
  jand g14528(.dina(n13627), .dinb(n6495), .dout(n14596));
  jand g14529(.dina(n13469), .dinb(n6503), .dout(n14597));
  jand g14530(.dina(n13478), .dinb(n6506), .dout(n14598));
  jand g14531(.dina(n13248), .dinb(n6500), .dout(n14599));
  jor  g14532(.dina(n14599), .dinb(n14598), .dout(n14600));
  jor  g14533(.dina(n14600), .dinb(n14597), .dout(n14601));
  jor  g14534(.dina(n14601), .dinb(n14596), .dout(n14602));
  jxor g14535(.dina(n14602), .dinb(n6219), .dout(n14603));
  jnot g14536(.din(n14603), .dout(n14604));
  jand g14537(.dina(n14604), .dinb(n14595), .dout(n14605));
  jnot g14538(.din(n14605), .dout(n14606));
  jor  g14539(.dina(n14604), .dinb(n14595), .dout(n14607));
  jnot g14540(.din(n14607), .dout(n14608));
  jxor g14541(.dina(n13986), .dinb(n13985), .dout(n14609));
  jand g14542(.dina(n13639), .dinb(n6495), .dout(n14610));
  jand g14543(.dina(n13478), .dinb(n6503), .dout(n14611));
  jand g14544(.dina(n13248), .dinb(n6506), .dout(n14612));
  jand g14545(.dina(n12669), .dinb(n6500), .dout(n14613));
  jor  g14546(.dina(n14613), .dinb(n14612), .dout(n14614));
  jor  g14547(.dina(n14614), .dinb(n14611), .dout(n14615));
  jor  g14548(.dina(n14615), .dinb(n14610), .dout(n14616));
  jxor g14549(.dina(n14616), .dinb(\a[2] ), .dout(n14617));
  jand g14550(.dina(n14617), .dinb(n14609), .dout(n14618));
  jnot g14551(.din(n14618), .dout(n14619));
  jor  g14552(.dina(n14617), .dinb(n14609), .dout(n14620));
  jnot g14553(.din(n14620), .dout(n14621));
  jxor g14554(.dina(n13983), .dinb(n13982), .dout(n14622));
  jand g14555(.dina(n13250), .dinb(n6495), .dout(n14623));
  jand g14556(.dina(n13248), .dinb(n6503), .dout(n14624));
  jand g14557(.dina(n12669), .dinb(n6506), .dout(n14625));
  jand g14558(.dina(n12536), .dinb(n6500), .dout(n14626));
  jor  g14559(.dina(n14626), .dinb(n14625), .dout(n14627));
  jor  g14560(.dina(n14627), .dinb(n14624), .dout(n14628));
  jor  g14561(.dina(n14628), .dinb(n14623), .dout(n14629));
  jxor g14562(.dina(n14629), .dinb(\a[2] ), .dout(n14630));
  jand g14563(.dina(n14630), .dinb(n14622), .dout(n14631));
  jnot g14564(.din(n14631), .dout(n14632));
  jor  g14565(.dina(n14630), .dinb(n14622), .dout(n14633));
  jnot g14566(.din(n14633), .dout(n14634));
  jxor g14567(.dina(n13980), .dinb(n13979), .dout(n14635));
  jand g14568(.dina(n12671), .dinb(n6495), .dout(n14636));
  jand g14569(.dina(n12669), .dinb(n6503), .dout(n14637));
  jand g14570(.dina(n12536), .dinb(n6506), .dout(n14638));
  jand g14571(.dina(n12547), .dinb(n6500), .dout(n14639));
  jor  g14572(.dina(n14639), .dinb(n14638), .dout(n14640));
  jor  g14573(.dina(n14640), .dinb(n14637), .dout(n14641));
  jor  g14574(.dina(n14641), .dinb(n14636), .dout(n14642));
  jxor g14575(.dina(n14642), .dinb(n6219), .dout(n14643));
  jnot g14576(.din(n14643), .dout(n14644));
  jand g14577(.dina(n14644), .dinb(n14635), .dout(n14645));
  jnot g14578(.din(n14645), .dout(n14646));
  jor  g14579(.dina(n14644), .dinb(n14635), .dout(n14647));
  jnot g14580(.din(n14647), .dout(n14648));
  jxor g14581(.dina(n13977), .dinb(n13976), .dout(n14649));
  jand g14582(.dina(n12684), .dinb(n6495), .dout(n14650));
  jand g14583(.dina(n12536), .dinb(n6503), .dout(n14651));
  jand g14584(.dina(n12547), .dinb(n6506), .dout(n14652));
  jand g14585(.dina(n12282), .dinb(n6500), .dout(n14653));
  jor  g14586(.dina(n14653), .dinb(n14652), .dout(n14654));
  jor  g14587(.dina(n14654), .dinb(n14651), .dout(n14655));
  jor  g14588(.dina(n14655), .dinb(n14650), .dout(n14656));
  jxor g14589(.dina(n14656), .dinb(n6219), .dout(n14657));
  jnot g14590(.din(n14657), .dout(n14658));
  jand g14591(.dina(n14658), .dinb(n14649), .dout(n14659));
  jnot g14592(.din(n14659), .dout(n14660));
  jor  g14593(.dina(n14658), .dinb(n14649), .dout(n14661));
  jnot g14594(.din(n14661), .dout(n14662));
  jxor g14595(.dina(n13974), .dinb(n13973), .dout(n14663));
  jand g14596(.dina(n12696), .dinb(n6495), .dout(n14664));
  jand g14597(.dina(n12547), .dinb(n6503), .dout(n14665));
  jand g14598(.dina(n12282), .dinb(n6506), .dout(n14666));
  jand g14599(.dina(n11798), .dinb(n6500), .dout(n14667));
  jor  g14600(.dina(n14667), .dinb(n14666), .dout(n14668));
  jor  g14601(.dina(n14668), .dinb(n14665), .dout(n14669));
  jor  g14602(.dina(n14669), .dinb(n14664), .dout(n14670));
  jxor g14603(.dina(n14670), .dinb(n6219), .dout(n14671));
  jnot g14604(.din(n14671), .dout(n14672));
  jand g14605(.dina(n14672), .dinb(n14663), .dout(n14673));
  jnot g14606(.din(n14673), .dout(n14674));
  jor  g14607(.dina(n14672), .dinb(n14663), .dout(n14675));
  jnot g14608(.din(n14675), .dout(n14676));
  jxor g14609(.dina(n13970), .dinb(n13969), .dout(n14677));
  jand g14610(.dina(n12284), .dinb(n6495), .dout(n14678));
  jand g14611(.dina(n12282), .dinb(n6503), .dout(n14679));
  jand g14612(.dina(n11798), .dinb(n6506), .dout(n14680));
  jand g14613(.dina(n11646), .dinb(n6500), .dout(n14681));
  jor  g14614(.dina(n14681), .dinb(n14680), .dout(n14682));
  jor  g14615(.dina(n14682), .dinb(n14679), .dout(n14683));
  jor  g14616(.dina(n14683), .dinb(n14678), .dout(n14684));
  jxor g14617(.dina(n14684), .dinb(n6219), .dout(n14685));
  jnot g14618(.din(n14685), .dout(n14686));
  jand g14619(.dina(n14686), .dinb(n14677), .dout(n14687));
  jnot g14620(.din(n14687), .dout(n14688));
  jor  g14621(.dina(n14686), .dinb(n14677), .dout(n14689));
  jnot g14622(.din(n14689), .dout(n14690));
  jxor g14623(.dina(n13967), .dinb(n13966), .dout(n14691));
  jand g14624(.dina(n11800), .dinb(n6495), .dout(n14692));
  jand g14625(.dina(n11798), .dinb(n6503), .dout(n14693));
  jand g14626(.dina(n11646), .dinb(n6506), .dout(n14694));
  jand g14627(.dina(n11647), .dinb(n6500), .dout(n14695));
  jor  g14628(.dina(n14695), .dinb(n14694), .dout(n14696));
  jor  g14629(.dina(n14696), .dinb(n14693), .dout(n14697));
  jor  g14630(.dina(n14697), .dinb(n14692), .dout(n14698));
  jxor g14631(.dina(n14698), .dinb(n6219), .dout(n14699));
  jnot g14632(.din(n14699), .dout(n14700));
  jand g14633(.dina(n14700), .dinb(n14691), .dout(n14701));
  jnot g14634(.din(n14701), .dout(n14702));
  jor  g14635(.dina(n14700), .dinb(n14691), .dout(n14703));
  jnot g14636(.din(n14703), .dout(n14704));
  jxor g14637(.dina(n13964), .dinb(n13963), .dout(n14705));
  jand g14638(.dina(n11812), .dinb(n6495), .dout(n14706));
  jand g14639(.dina(n11646), .dinb(n6503), .dout(n14707));
  jand g14640(.dina(n11647), .dinb(n6506), .dout(n14708));
  jand g14641(.dina(n11306), .dinb(n6500), .dout(n14709));
  jor  g14642(.dina(n14709), .dinb(n14708), .dout(n14710));
  jor  g14643(.dina(n14710), .dinb(n14707), .dout(n14711));
  jor  g14644(.dina(n14711), .dinb(n14706), .dout(n14712));
  jxor g14645(.dina(n14712), .dinb(\a[2] ), .dout(n14713));
  jand g14646(.dina(n14713), .dinb(n14705), .dout(n14714));
  jnot g14647(.din(n14714), .dout(n14715));
  jor  g14648(.dina(n14713), .dinb(n14705), .dout(n14716));
  jnot g14649(.din(n14716), .dout(n14717));
  jxor g14650(.dina(n13961), .dinb(n13960), .dout(n14718));
  jand g14651(.dina(n11824), .dinb(n6495), .dout(n14719));
  jand g14652(.dina(n11647), .dinb(n6503), .dout(n14720));
  jand g14653(.dina(n11306), .dinb(n6506), .dout(n14721));
  jand g14654(.dina(n10836), .dinb(n6500), .dout(n14722));
  jor  g14655(.dina(n14722), .dinb(n14721), .dout(n14723));
  jor  g14656(.dina(n14723), .dinb(n14720), .dout(n14724));
  jor  g14657(.dina(n14724), .dinb(n14719), .dout(n14725));
  jxor g14658(.dina(n14725), .dinb(\a[2] ), .dout(n14726));
  jand g14659(.dina(n14726), .dinb(n14718), .dout(n14727));
  jnot g14660(.din(n14727), .dout(n14728));
  jor  g14661(.dina(n14726), .dinb(n14718), .dout(n14729));
  jnot g14662(.din(n14729), .dout(n14730));
  jxor g14663(.dina(n13958), .dinb(n13957), .dout(n14731));
  jnot g14664(.din(n14731), .dout(n14732));
  jxor g14665(.dina(n13955), .dinb(n13953), .dout(n14733));
  jand g14666(.dina(n10838), .dinb(n6495), .dout(n14734));
  jand g14667(.dina(n10836), .dinb(n6503), .dout(n14735));
  jand g14668(.dina(n10640), .dinb(n6506), .dout(n14736));
  jand g14669(.dina(n10647), .dinb(n6500), .dout(n14737));
  jor  g14670(.dina(n14737), .dinb(n14736), .dout(n14738));
  jor  g14671(.dina(n14738), .dinb(n14735), .dout(n14739));
  jor  g14672(.dina(n14739), .dinb(n14734), .dout(n14740));
  jxor g14673(.dina(n14740), .dinb(n6219), .dout(n14741));
  jnot g14674(.din(n14741), .dout(n14742));
  jand g14675(.dina(n14742), .dinb(n14733), .dout(n14743));
  jor  g14676(.dina(n14742), .dinb(n14733), .dout(n14744));
  jxor g14677(.dina(n13951), .dinb(n13949), .dout(n14745));
  jand g14678(.dina(n10850), .dinb(n6495), .dout(n14746));
  jand g14679(.dina(n10640), .dinb(n6503), .dout(n14747));
  jand g14680(.dina(n10647), .dinb(n6506), .dout(n14748));
  jand g14681(.dina(n10305), .dinb(n6500), .dout(n14749));
  jor  g14682(.dina(n14749), .dinb(n14748), .dout(n14750));
  jor  g14683(.dina(n14750), .dinb(n14747), .dout(n14751));
  jor  g14684(.dina(n14751), .dinb(n14746), .dout(n14752));
  jxor g14685(.dina(n14752), .dinb(\a[2] ), .dout(n14753));
  jand g14686(.dina(n14753), .dinb(n14745), .dout(n14754));
  jxor g14687(.dina(n13947), .dinb(n13945), .dout(n14755));
  jand g14688(.dina(n10862), .dinb(n6495), .dout(n14756));
  jand g14689(.dina(n10647), .dinb(n6503), .dout(n14757));
  jand g14690(.dina(n10305), .dinb(n6506), .dout(n14758));
  jand g14691(.dina(n9872), .dinb(n6500), .dout(n14759));
  jor  g14692(.dina(n14759), .dinb(n14758), .dout(n14760));
  jor  g14693(.dina(n14760), .dinb(n14757), .dout(n14761));
  jor  g14694(.dina(n14761), .dinb(n14756), .dout(n14762));
  jxor g14695(.dina(n14762), .dinb(n6219), .dout(n14763));
  jnot g14696(.din(n14763), .dout(n14764));
  jand g14697(.dina(n14764), .dinb(n14755), .dout(n14765));
  jor  g14698(.dina(n14764), .dinb(n14755), .dout(n14766));
  jxor g14699(.dina(n13943), .dinb(n13941), .dout(n14767));
  jnot g14700(.din(n14767), .dout(n14768));
  jnot g14701(.din(n10307), .dout(n14769));
  jor  g14702(.dina(n14769), .dinb(n6496), .dout(n14770));
  jnot g14703(.din(n10305), .dout(n14771));
  jor  g14704(.dina(n14771), .dinb(n6504), .dout(n14772));
  jnot g14705(.din(n9872), .dout(n14773));
  jor  g14706(.dina(n14773), .dinb(n6507), .dout(n14774));
  jnot g14707(.din(n9655), .dout(n14775));
  jor  g14708(.dina(n14775), .dinb(n6501), .dout(n14776));
  jand g14709(.dina(n14776), .dinb(n14774), .dout(n14777));
  jand g14710(.dina(n14777), .dinb(n14772), .dout(n14778));
  jand g14711(.dina(n14778), .dinb(n14770), .dout(n14779));
  jxor g14712(.dina(n14779), .dinb(n6219), .dout(n14780));
  jnot g14713(.din(n14780), .dout(n14781));
  jand g14714(.dina(n14781), .dinb(n14768), .dout(n14782));
  jand g14715(.dina(n14780), .dinb(n14767), .dout(n14783));
  jnot g14716(.din(n14783), .dout(n14784));
  jxor g14717(.dina(n13939), .dinb(n13937), .dout(n14785));
  jnot g14718(.din(n14785), .dout(n14786));
  jnot g14719(.din(n9874), .dout(n14787));
  jor  g14720(.dina(n14787), .dinb(n6496), .dout(n14788));
  jor  g14721(.dina(n14773), .dinb(n6504), .dout(n14789));
  jor  g14722(.dina(n14775), .dinb(n6507), .dout(n14790));
  jnot g14723(.din(n9656), .dout(n14791));
  jor  g14724(.dina(n14791), .dinb(n6501), .dout(n14792));
  jand g14725(.dina(n14792), .dinb(n14790), .dout(n14793));
  jand g14726(.dina(n14793), .dinb(n14789), .dout(n14794));
  jand g14727(.dina(n14794), .dinb(n14788), .dout(n14795));
  jxor g14728(.dina(n14795), .dinb(n6219), .dout(n14796));
  jnot g14729(.din(n14796), .dout(n14797));
  jand g14730(.dina(n14797), .dinb(n14786), .dout(n14798));
  jand g14731(.dina(n14796), .dinb(n14785), .dout(n14799));
  jnot g14732(.din(n14799), .dout(n14800));
  jxor g14733(.dina(n13934), .dinb(n13933), .dout(n14801));
  jnot g14734(.din(n14801), .dout(n14802));
  jand g14735(.dina(n9886), .dinb(n6495), .dout(n14803));
  jand g14736(.dina(n9655), .dinb(n6503), .dout(n14804));
  jand g14737(.dina(n9656), .dinb(n6506), .dout(n14805));
  jand g14738(.dina(n9250), .dinb(n6500), .dout(n14806));
  jor  g14739(.dina(n14806), .dinb(n14805), .dout(n14807));
  jor  g14740(.dina(n14807), .dinb(n14804), .dout(n14808));
  jor  g14741(.dina(n14808), .dinb(n14803), .dout(n14809));
  jxor g14742(.dina(n14809), .dinb(n6219), .dout(n14810));
  jand g14743(.dina(n14810), .dinb(n14802), .dout(n14811));
  jor  g14744(.dina(n14810), .dinb(n14802), .dout(n14812));
  jxor g14745(.dina(n13929), .dinb(n13928), .dout(n14813));
  jnot g14746(.din(n14813), .dout(n14814));
  jand g14747(.dina(n9898), .dinb(n6495), .dout(n14815));
  jand g14748(.dina(n9656), .dinb(n6503), .dout(n14816));
  jand g14749(.dina(n9250), .dinb(n6506), .dout(n14817));
  jand g14750(.dina(n8936), .dinb(n6500), .dout(n14818));
  jor  g14751(.dina(n14818), .dinb(n14817), .dout(n14819));
  jor  g14752(.dina(n14819), .dinb(n14816), .dout(n14820));
  jor  g14753(.dina(n14820), .dinb(n14815), .dout(n14821));
  jxor g14754(.dina(n14821), .dinb(n6219), .dout(n14822));
  jand g14755(.dina(n14822), .dinb(n14814), .dout(n14823));
  jnot g14756(.din(n14823), .dout(n14824));
  jor  g14757(.dina(n14822), .dinb(n14814), .dout(n14825));
  jnot g14758(.din(n14825), .dout(n14826));
  jxor g14759(.dina(n13926), .dinb(n13925), .dout(n14827));
  jnot g14760(.din(n14827), .dout(n14828));
  jand g14761(.dina(n9252), .dinb(n6495), .dout(n14829));
  jand g14762(.dina(n9250), .dinb(n6503), .dout(n14830));
  jand g14763(.dina(n8936), .dinb(n6506), .dout(n14831));
  jand g14764(.dina(n8723), .dinb(n6500), .dout(n14832));
  jor  g14765(.dina(n14832), .dinb(n14831), .dout(n14833));
  jor  g14766(.dina(n14833), .dinb(n14830), .dout(n14834));
  jor  g14767(.dina(n14834), .dinb(n14829), .dout(n14835));
  jxor g14768(.dina(n14835), .dinb(n6219), .dout(n14836));
  jand g14769(.dina(n14836), .dinb(n14828), .dout(n14837));
  jnot g14770(.din(n14837), .dout(n14838));
  jor  g14771(.dina(n14836), .dinb(n14828), .dout(n14839));
  jnot g14772(.din(n14839), .dout(n14840));
  jxor g14773(.dina(n13921), .dinb(n13920), .dout(n14841));
  jand g14774(.dina(n8938), .dinb(n6495), .dout(n14842));
  jand g14775(.dina(n8936), .dinb(n6503), .dout(n14843));
  jand g14776(.dina(n8723), .dinb(n6506), .dout(n14844));
  jand g14777(.dina(n8740), .dinb(n6500), .dout(n14845));
  jor  g14778(.dina(n14845), .dinb(n14844), .dout(n14846));
  jor  g14779(.dina(n14846), .dinb(n14843), .dout(n14847));
  jor  g14780(.dina(n14847), .dinb(n14842), .dout(n14848));
  jxor g14781(.dina(n14848), .dinb(\a[2] ), .dout(n14849));
  jand g14782(.dina(n14849), .dinb(n14841), .dout(n14850));
  jxor g14783(.dina(n13917), .dinb(n13909), .dout(n14851));
  jnot g14784(.din(n14851), .dout(n14852));
  jand g14785(.dina(n8950), .dinb(n6495), .dout(n14853));
  jand g14786(.dina(n8723), .dinb(n6503), .dout(n14854));
  jand g14787(.dina(n8740), .dinb(n6506), .dout(n14855));
  jand g14788(.dina(n8268), .dinb(n6500), .dout(n14856));
  jor  g14789(.dina(n14856), .dinb(n14855), .dout(n14857));
  jor  g14790(.dina(n14857), .dinb(n14854), .dout(n14858));
  jor  g14791(.dina(n14858), .dinb(n14853), .dout(n14859));
  jxor g14792(.dina(n14859), .dinb(n6219), .dout(n14860));
  jand g14793(.dina(n14860), .dinb(n14852), .dout(n14861));
  jnot g14794(.din(n14861), .dout(n14862));
  jor  g14795(.dina(n14860), .dinb(n14852), .dout(n14863));
  jnot g14796(.din(n14863), .dout(n14864));
  jor  g14797(.dina(n13896), .dinb(n5277), .dout(n14865));
  jxor g14798(.dina(n14865), .dinb(n13904), .dout(n14866));
  jand g14799(.dina(n8962), .dinb(n6495), .dout(n14867));
  jand g14800(.dina(n8740), .dinb(n6503), .dout(n14868));
  jand g14801(.dina(n8268), .dinb(n6506), .dout(n14869));
  jand g14802(.dina(n8022), .dinb(n6500), .dout(n14870));
  jor  g14803(.dina(n14870), .dinb(n14869), .dout(n14871));
  jor  g14804(.dina(n14871), .dinb(n14868), .dout(n14872));
  jor  g14805(.dina(n14872), .dinb(n14867), .dout(n14873));
  jxor g14806(.dina(n14873), .dinb(\a[2] ), .dout(n14874));
  jand g14807(.dina(n14874), .dinb(n14866), .dout(n14875));
  jand g14808(.dina(n7692), .dinb(n6503), .dout(n14876));
  jnot g14809(.din(n14876), .dout(n14877));
  jand g14810(.dina(n8024), .dinb(n7019), .dout(n14878));
  jnot g14811(.din(n14878), .dout(n14879));
  jnot g14812(.din(n7326), .dout(n14880));
  jand g14813(.dina(n8025), .dinb(n14880), .dout(n14881));
  jand g14814(.dina(n14881), .dinb(n14879), .dout(n14882));
  jor  g14815(.dina(n14882), .dinb(n6861), .dout(n14883));
  jand g14816(.dina(n7021), .dinb(\a[2] ), .dout(n14884));
  jand g14817(.dina(n7313), .dinb(n6856), .dout(n14885));
  jnot g14818(.din(n14885), .dout(n14886));
  jand g14819(.dina(n14886), .dinb(n14884), .dout(n14887));
  jand g14820(.dina(n14887), .dinb(n14883), .dout(n14888));
  jand g14821(.dina(n14888), .dinb(n14877), .dout(n14889));
  jor  g14822(.dina(n14889), .dinb(n13893), .dout(n14891));
  jand g14823(.dina(n8029), .dinb(n6495), .dout(n14892));
  jand g14824(.dina(n8022), .dinb(n6503), .dout(n14893));
  jand g14825(.dina(n7692), .dinb(n6506), .dout(n14894));
  jand g14826(.dina(n7313), .dinb(n6500), .dout(n14895));
  jor  g14827(.dina(n14895), .dinb(n14894), .dout(n14896));
  jor  g14828(.dina(n14896), .dinb(n14893), .dout(n14897));
  jor  g14829(.dina(n14897), .dinb(n14892), .dout(n14898));
  jxor g14830(.dina(n14898), .dinb(n6219), .dout(n14899));
  jnot g14831(.din(n14899), .dout(n14900));
  jand g14832(.dina(n14900), .dinb(n14891), .dout(n14901));
  jand g14833(.dina(n8270), .dinb(n6495), .dout(n14903));
  jand g14834(.dina(n8268), .dinb(n6503), .dout(n14904));
  jand g14835(.dina(n8022), .dinb(n6506), .dout(n14905));
  jand g14836(.dina(n7692), .dinb(n6500), .dout(n14906));
  jor  g14837(.dina(n14906), .dinb(n14905), .dout(n14907));
  jor  g14838(.dina(n14907), .dinb(n14904), .dout(n14908));
  jor  g14839(.dina(n14908), .dinb(n14903), .dout(n14909));
  jxor g14840(.dina(n14909), .dinb(n6219), .dout(n14910));
  jnot g14841(.din(n14910), .dout(n14911));
  jand g14842(.dina(n14911), .dinb(n14901), .dout(n14912));
  jor  g14843(.dina(n14911), .dinb(n14901), .dout(n14913));
  jand g14844(.dina(n13893), .dinb(\a[5] ), .dout(n14914));
  jxor g14845(.dina(n14914), .dinb(n13891), .dout(n14915));
  jand g14846(.dina(n14915), .dinb(n14913), .dout(n14916));
  jor  g14847(.dina(n14916), .dinb(n14912), .dout(n14917));
  jor  g14848(.dina(n14874), .dinb(n14866), .dout(n14918));
  jand g14849(.dina(n14918), .dinb(n14917), .dout(n14919));
  jor  g14850(.dina(n14919), .dinb(n14875), .dout(n14920));
  jor  g14851(.dina(n14920), .dinb(n14864), .dout(n14921));
  jand g14852(.dina(n14921), .dinb(n14862), .dout(n14922));
  jor  g14853(.dina(n14849), .dinb(n14841), .dout(n14923));
  jand g14854(.dina(n14923), .dinb(n14922), .dout(n14924));
  jor  g14855(.dina(n14924), .dinb(n14850), .dout(n14925));
  jor  g14856(.dina(n14925), .dinb(n14840), .dout(n14926));
  jand g14857(.dina(n14926), .dinb(n14838), .dout(n14927));
  jor  g14858(.dina(n14927), .dinb(n14826), .dout(n14928));
  jand g14859(.dina(n14928), .dinb(n14824), .dout(n14929));
  jnot g14860(.din(n14929), .dout(n14930));
  jand g14861(.dina(n14930), .dinb(n14812), .dout(n14931));
  jor  g14862(.dina(n14931), .dinb(n14811), .dout(n14932));
  jand g14863(.dina(n14932), .dinb(n14800), .dout(n14933));
  jor  g14864(.dina(n14933), .dinb(n14798), .dout(n14934));
  jand g14865(.dina(n14934), .dinb(n14784), .dout(n14935));
  jor  g14866(.dina(n14935), .dinb(n14782), .dout(n14936));
  jnot g14867(.din(n14936), .dout(n14937));
  jand g14868(.dina(n14937), .dinb(n14766), .dout(n14938));
  jor  g14869(.dina(n14938), .dinb(n14765), .dout(n14939));
  jor  g14870(.dina(n14753), .dinb(n14745), .dout(n14940));
  jand g14871(.dina(n14940), .dinb(n14939), .dout(n14941));
  jor  g14872(.dina(n14941), .dinb(n14754), .dout(n14942));
  jand g14873(.dina(n14942), .dinb(n14744), .dout(n14943));
  jor  g14874(.dina(n14943), .dinb(n14743), .dout(n14944));
  jnot g14875(.din(n14944), .dout(n14945));
  jand g14876(.dina(n14945), .dinb(n14732), .dout(n14946));
  jand g14877(.dina(n14944), .dinb(n14731), .dout(n14947));
  jnot g14878(.din(n14947), .dout(n14948));
  jnot g14879(.din(n11308), .dout(n14949));
  jor  g14880(.dina(n14949), .dinb(n6496), .dout(n14950));
  jnot g14881(.din(n11306), .dout(n14951));
  jor  g14882(.dina(n14951), .dinb(n6504), .dout(n14952));
  jnot g14883(.din(n10836), .dout(n14953));
  jor  g14884(.dina(n14953), .dinb(n6507), .dout(n14954));
  jnot g14885(.din(n10640), .dout(n14955));
  jor  g14886(.dina(n14955), .dinb(n6501), .dout(n14956));
  jand g14887(.dina(n14956), .dinb(n14954), .dout(n14957));
  jand g14888(.dina(n14957), .dinb(n14952), .dout(n14958));
  jand g14889(.dina(n14958), .dinb(n14950), .dout(n14959));
  jxor g14890(.dina(n14959), .dinb(\a[2] ), .dout(n14960));
  jand g14891(.dina(n14960), .dinb(n14948), .dout(n14961));
  jor  g14892(.dina(n14961), .dinb(n14946), .dout(n14962));
  jor  g14893(.dina(n14962), .dinb(n14730), .dout(n14963));
  jand g14894(.dina(n14963), .dinb(n14728), .dout(n14964));
  jor  g14895(.dina(n14964), .dinb(n14717), .dout(n14965));
  jand g14896(.dina(n14965), .dinb(n14715), .dout(n14966));
  jor  g14897(.dina(n14966), .dinb(n14704), .dout(n14967));
  jand g14898(.dina(n14967), .dinb(n14702), .dout(n14968));
  jor  g14899(.dina(n14968), .dinb(n14690), .dout(n14969));
  jand g14900(.dina(n14969), .dinb(n14688), .dout(n14970));
  jor  g14901(.dina(n14970), .dinb(n14676), .dout(n14971));
  jand g14902(.dina(n14971), .dinb(n14674), .dout(n14972));
  jor  g14903(.dina(n14972), .dinb(n14662), .dout(n14973));
  jand g14904(.dina(n14973), .dinb(n14660), .dout(n14974));
  jor  g14905(.dina(n14974), .dinb(n14648), .dout(n14975));
  jand g14906(.dina(n14975), .dinb(n14646), .dout(n14976));
  jor  g14907(.dina(n14976), .dinb(n14634), .dout(n14977));
  jand g14908(.dina(n14977), .dinb(n14632), .dout(n14978));
  jor  g14909(.dina(n14978), .dinb(n14621), .dout(n14979));
  jand g14910(.dina(n14979), .dinb(n14619), .dout(n14980));
  jor  g14911(.dina(n14980), .dinb(n14608), .dout(n14981));
  jand g14912(.dina(n14981), .dinb(n14606), .dout(n14982));
  jand g14913(.dina(n14982), .dinb(n14594), .dout(n14983));
  jor  g14914(.dina(n14982), .dinb(n14594), .dout(n14984));
  jnot g14915(.din(n13616), .dout(n14985));
  jor  g14916(.dina(n14985), .dinb(n6496), .dout(n14986));
  jor  g14917(.dina(n14584), .dinb(n6504), .dout(n14987));
  jnot g14918(.din(n13469), .dout(n14988));
  jor  g14919(.dina(n14988), .dinb(n6507), .dout(n14989));
  jnot g14920(.din(n13478), .dout(n14990));
  jor  g14921(.dina(n14990), .dinb(n6501), .dout(n14991));
  jand g14922(.dina(n14991), .dinb(n14989), .dout(n14992));
  jand g14923(.dina(n14992), .dinb(n14987), .dout(n14993));
  jand g14924(.dina(n14993), .dinb(n14986), .dout(n14994));
  jxor g14925(.dina(n14994), .dinb(\a[2] ), .dout(n14995));
  jand g14926(.dina(n14995), .dinb(n14984), .dout(n14996));
  jor  g14927(.dina(n14996), .dinb(n14983), .dout(n14997));
  jxor g14928(.dina(n13995), .dinb(n13994), .dout(n14998));
  jnot g14929(.din(n14998), .dout(n14999));
  jnot g14930(.din(n14251), .dout(n15000));
  jor  g14931(.dina(n15000), .dinb(n6496), .dout(n15001));
  jor  g14932(.dina(n14569), .dinb(n6504), .dout(n15002));
  jor  g14933(.dina(n14584), .dinb(n6507), .dout(n15003));
  jor  g14934(.dina(n14988), .dinb(n6501), .dout(n15004));
  jand g14935(.dina(n15004), .dinb(n15003), .dout(n15005));
  jand g14936(.dina(n15005), .dinb(n15002), .dout(n15006));
  jand g14937(.dina(n15006), .dinb(n15001), .dout(n15007));
  jxor g14938(.dina(n15007), .dinb(n6219), .dout(n15008));
  jnot g14939(.din(n15008), .dout(n15009));
  jand g14940(.dina(n15009), .dinb(n14999), .dout(n15010));
  jor  g14941(.dina(n15010), .dinb(n14997), .dout(n15011));
  jnot g14942(.din(n15011), .dout(n15012));
  jand g14943(.dina(n14589), .dinb(n14577), .dout(n15013));
  jand g14944(.dina(n15008), .dinb(n14998), .dout(n15014));
  jor  g14945(.dina(n15014), .dinb(n15013), .dout(n15015));
  jor  g14946(.dina(n15015), .dinb(n15012), .dout(n15016));
  jand g14947(.dina(n15016), .dinb(n14592), .dout(n15017));
  jand g14948(.dina(n15017), .dinb(n14576), .dout(n15018));
  jor  g14949(.dina(n15018), .dinb(n14575), .dout(n15019));
  jxor g14950(.dina(n15019), .dinb(n14560), .dout(n15020));
  jand g14951(.dina(n15020), .dinb(n64), .dout(n15021));
  jnot g14952(.din(n15020), .dout(n15022));
  jor  g14953(.dina(n14559), .dinb(n14262), .dout(n15023));
  jnot g14954(.din(n15023), .dout(n15024));
  jand g14955(.dina(n15019), .dinb(n14560), .dout(n15025));
  jor  g14956(.dina(n15025), .dinb(n15024), .dout(n15026));
  jnot g14957(.din(n14173), .dout(n15027));
  jor  g14958(.dina(n14259), .dinb(n15027), .dout(n15028));
  jor  g14959(.dina(n14260), .dinb(n14004), .dout(n15029));
  jand g14960(.dina(n15029), .dinb(n15028), .dout(n15030));
  jnot g14961(.din(n14162), .dout(n15031));
  jor  g14962(.dina(n14170), .dinb(n15031), .dout(n15032));
  jnot g14963(.din(n15032), .dout(n15033));
  jand g14964(.dina(n14172), .dinb(n14009), .dout(n15034));
  jor  g14965(.dina(n15034), .dinb(n15033), .dout(n15035));
  jnot g14966(.din(n14152), .dout(n15036));
  jand g14967(.dina(n14160), .dinb(n15036), .dout(n15037));
  jnot g14968(.din(n15037), .dout(n15038));
  jor  g14969(.dina(n14161), .dinb(n14013), .dout(n15039));
  jand g14970(.dina(n15039), .dinb(n15038), .dout(n15040));
  jnot g14971(.din(n15040), .dout(n15041));
  jnot g14972(.din(n14142), .dout(n15042));
  jor  g14973(.dina(n14150), .dinb(n15042), .dout(n15043));
  jnot g14974(.din(n14151), .dout(n15044));
  jand g14975(.dina(n15044), .dinb(n14017), .dout(n15045));
  jnot g14976(.din(n15045), .dout(n15046));
  jand g14977(.dina(n15046), .dinb(n15043), .dout(n15047));
  jor  g14978(.dina(n14140), .dinb(n14132), .dout(n15048));
  jnot g14979(.din(n15048), .dout(n15049));
  jand g14980(.dina(n14141), .dinb(n14022), .dout(n15050));
  jor  g14981(.dina(n15050), .dinb(n15049), .dout(n15051));
  jor  g14982(.dina(n14129), .dinb(n14121), .dout(n15052));
  jand g14983(.dina(n14130), .dinb(n14027), .dout(n15053));
  jnot g14984(.din(n15053), .dout(n15054));
  jand g14985(.dina(n15054), .dinb(n15052), .dout(n15055));
  jnot g14986(.din(n15055), .dout(n15056));
  jor  g14987(.dina(n14118), .dinb(n14110), .dout(n15057));
  jand g14988(.dina(n14119), .dinb(n14032), .dout(n15058));
  jnot g14989(.din(n15058), .dout(n15059));
  jand g14990(.dina(n15059), .dinb(n15057), .dout(n15060));
  jnot g14991(.din(n15060), .dout(n15061));
  jor  g14992(.dina(n14107), .dinb(n14099), .dout(n15062));
  jand g14993(.dina(n14108), .dinb(n14035), .dout(n15063));
  jnot g14994(.din(n15063), .dout(n15064));
  jand g14995(.dina(n15064), .dinb(n15062), .dout(n15065));
  jnot g14996(.din(n15065), .dout(n15066));
  jor  g14997(.dina(n14096), .dinb(n14088), .dout(n15067));
  jand g14998(.dina(n14097), .dinb(n14040), .dout(n15068));
  jnot g14999(.din(n15068), .dout(n15069));
  jand g15000(.dina(n15069), .dinb(n15067), .dout(n15070));
  jnot g15001(.din(n15070), .dout(n15071));
  jand g15002(.dina(n7693), .dinb(n5076), .dout(n15072));
  jand g15003(.dina(n7313), .dinb(n5082), .dout(n15073));
  jor  g15004(.dina(n15073), .dinb(n15072), .dout(n15074));
  jand g15005(.dina(n7692), .dinb(n5084), .dout(n15075));
  jand g15006(.dina(n7019), .dinb(n6050), .dout(n15076));
  jor  g15007(.dina(n15076), .dinb(n15075), .dout(n15077));
  jor  g15008(.dina(n15077), .dinb(n15074), .dout(n15078));
  jand g15009(.dina(n14086), .dinb(n14081), .dout(n15079));
  jnot g15010(.din(n15079), .dout(n15080));
  jand g15011(.dina(n978), .dinb(n645), .dout(n15081));
  jand g15012(.dina(n15081), .dinb(n1516), .dout(n15082));
  jand g15013(.dina(n15082), .dinb(n1721), .dout(n15083));
  jand g15014(.dina(n10739), .dinb(n678), .dout(n15084));
  jand g15015(.dina(n15084), .dinb(n15083), .dout(n15085));
  jand g15016(.dina(n15085), .dinb(n5349), .dout(n15086));
  jand g15017(.dina(n1714), .dinb(n492), .dout(n15087));
  jand g15018(.dina(n3762), .dinb(n713), .dout(n15088));
  jand g15019(.dina(n15088), .dinb(n15087), .dout(n15089));
  jand g15020(.dina(n15089), .dinb(n2465), .dout(n15090));
  jand g15021(.dina(n472), .dinb(n638), .dout(n15091));
  jand g15022(.dina(n15091), .dinb(n1260), .dout(n15092));
  jand g15023(.dina(n15092), .dinb(n1744), .dout(n15093));
  jand g15024(.dina(n15093), .dinb(n3819), .dout(n15094));
  jand g15025(.dina(n15094), .dinb(n15090), .dout(n15095));
  jand g15026(.dina(n15095), .dinb(n2487), .dout(n15096));
  jand g15027(.dina(n1305), .dinb(n871), .dout(n15097));
  jand g15028(.dina(n15097), .dinb(n933), .dout(n15098));
  jand g15029(.dina(n15098), .dinb(n1851), .dout(n15099));
  jand g15030(.dina(n15099), .dinb(n1165), .dout(n15100));
  jand g15031(.dina(n6158), .dinb(n1976), .dout(n15101));
  jand g15032(.dina(n1246), .dinb(n2148), .dout(n15102));
  jand g15033(.dina(n583), .dinb(n510), .dout(n15103));
  jand g15034(.dina(n15103), .dinb(n15102), .dout(n15104));
  jand g15035(.dina(n15104), .dinb(n2089), .dout(n15105));
  jand g15036(.dina(n15105), .dinb(n15101), .dout(n15106));
  jand g15037(.dina(n15106), .dinb(n15100), .dout(n15107));
  jand g15038(.dina(n15107), .dinb(n15096), .dout(n15108));
  jand g15039(.dina(n1522), .dinb(n503), .dout(n15109));
  jand g15040(.dina(n15109), .dinb(n1373), .dout(n15110));
  jand g15041(.dina(n14071), .dinb(n2587), .dout(n15111));
  jand g15042(.dina(n3857), .dinb(n1042), .dout(n15112));
  jand g15043(.dina(n15112), .dinb(n15111), .dout(n15113));
  jand g15044(.dina(n15113), .dinb(n15110), .dout(n15114));
  jnot g15045(.din(n943), .dout(n15115));
  jand g15046(.dina(n5232), .dinb(n2580), .dout(n15116));
  jand g15047(.dina(n15116), .dinb(n15115), .dout(n15117));
  jand g15048(.dina(n1541), .dinb(n1708), .dout(n15118));
  jand g15049(.dina(n15118), .dinb(n1016), .dout(n15119));
  jand g15050(.dina(n15119), .dinb(n2521), .dout(n15120));
  jand g15051(.dina(n15120), .dinb(n15117), .dout(n15121));
  jand g15052(.dina(n15121), .dinb(n15114), .dout(n15122));
  jand g15053(.dina(n843), .dinb(n493), .dout(n15123));
  jand g15054(.dina(n15123), .dinb(n6241), .dout(n15124));
  jand g15055(.dina(n2538), .dinb(n670), .dout(n15125));
  jand g15056(.dina(n15125), .dinb(n15124), .dout(n15126));
  jand g15057(.dina(n6343), .dinb(n1308), .dout(n15127));
  jand g15058(.dina(n15127), .dinb(n14286), .dout(n15128));
  jand g15059(.dina(n15128), .dinb(n15126), .dout(n15129));
  jand g15060(.dina(n534), .dinb(n495), .dout(n15130));
  jand g15061(.dina(n15130), .dinb(n1309), .dout(n15131));
  jand g15062(.dina(n881), .dinb(n542), .dout(n15132));
  jand g15063(.dina(n15132), .dinb(n2454), .dout(n15133));
  jand g15064(.dina(n15133), .dinb(n6299), .dout(n15134));
  jand g15065(.dina(n15134), .dinb(n15131), .dout(n15135));
  jand g15066(.dina(n15135), .dinb(n15129), .dout(n15136));
  jand g15067(.dina(n15136), .dinb(n15122), .dout(n15137));
  jand g15068(.dina(n15137), .dinb(n15108), .dout(n15138));
  jand g15069(.dina(n15138), .dinb(n15086), .dout(n15139));
  jxor g15070(.dina(n15139), .dinb(n15080), .dout(n15140));
  jxor g15071(.dina(n15140), .dinb(n15078), .dout(n15141));
  jnot g15072(.din(n15141), .dout(n15142));
  jand g15073(.dina(n8962), .dinb(n2936), .dout(n15143));
  jand g15074(.dina(n8268), .dinb(n2940), .dout(n15144));
  jand g15075(.dina(n8740), .dinb(n2943), .dout(n15145));
  jor  g15076(.dina(n15145), .dinb(n15144), .dout(n15146));
  jand g15077(.dina(n8022), .dinb(n3684), .dout(n15147));
  jor  g15078(.dina(n15147), .dinb(n15146), .dout(n15148));
  jor  g15079(.dina(n15148), .dinb(n15143), .dout(n15149));
  jxor g15080(.dina(n15149), .dinb(n93), .dout(n15150));
  jxor g15081(.dina(n15150), .dinb(n15142), .dout(n15151));
  jxor g15082(.dina(n15151), .dinb(n15071), .dout(n15152));
  jnot g15083(.din(n15152), .dout(n15153));
  jand g15084(.dina(n9252), .dinb(n71), .dout(n15154));
  jand g15085(.dina(n9250), .dinb(n796), .dout(n15155));
  jand g15086(.dina(n8723), .dinb(n1806), .dout(n15156));
  jand g15087(.dina(n8936), .dinb(n731), .dout(n15157));
  jor  g15088(.dina(n15157), .dinb(n15156), .dout(n15158));
  jor  g15089(.dina(n15158), .dinb(n15155), .dout(n15159));
  jor  g15090(.dina(n15159), .dinb(n15154), .dout(n15160));
  jxor g15091(.dina(n15160), .dinb(n77), .dout(n15161));
  jxor g15092(.dina(n15161), .dinb(n15153), .dout(n15162));
  jxor g15093(.dina(n15162), .dinb(n15066), .dout(n15163));
  jnot g15094(.din(n15163), .dout(n15164));
  jand g15095(.dina(n9874), .dinb(n806), .dout(n15165));
  jand g15096(.dina(n9655), .dinb(n1612), .dout(n15166));
  jand g15097(.dina(n9872), .dinb(n1620), .dout(n15167));
  jor  g15098(.dina(n15167), .dinb(n15166), .dout(n15168));
  jand g15099(.dina(n9656), .dinb(n1644), .dout(n15169));
  jor  g15100(.dina(n15169), .dinb(n15168), .dout(n15170));
  jor  g15101(.dina(n15170), .dinb(n15165), .dout(n15171));
  jxor g15102(.dina(n15171), .dinb(n65), .dout(n15172));
  jxor g15103(.dina(n15172), .dinb(n15164), .dout(n15173));
  jxor g15104(.dina(n15173), .dinb(n15061), .dout(n15174));
  jnot g15105(.din(n15174), .dout(n15175));
  jand g15106(.dina(n10850), .dinb(n1819), .dout(n15176));
  jand g15107(.dina(n10640), .dinb(n2243), .dout(n15177));
  jand g15108(.dina(n10647), .dinb(n2180), .dout(n15178));
  jand g15109(.dina(n10305), .dinb(n2185), .dout(n15179));
  jor  g15110(.dina(n15179), .dinb(n15178), .dout(n15180));
  jor  g15111(.dina(n15180), .dinb(n15177), .dout(n15181));
  jor  g15112(.dina(n15181), .dinb(n15176), .dout(n15182));
  jxor g15113(.dina(n15182), .dinb(n2196), .dout(n15183));
  jxor g15114(.dina(n15183), .dinb(n15175), .dout(n15184));
  jxor g15115(.dina(n15184), .dinb(n15056), .dout(n15185));
  jnot g15116(.din(n15185), .dout(n15186));
  jand g15117(.dina(n11824), .dinb(n2743), .dout(n15187));
  jand g15118(.dina(n11647), .dinb(n2752), .dout(n15188));
  jand g15119(.dina(n11306), .dinb(n2748), .dout(n15189));
  jand g15120(.dina(n10836), .dinb(n2757), .dout(n15190));
  jor  g15121(.dina(n15190), .dinb(n15189), .dout(n15191));
  jor  g15122(.dina(n15191), .dinb(n15188), .dout(n15192));
  jor  g15123(.dina(n15192), .dinb(n15187), .dout(n15193));
  jxor g15124(.dina(n15193), .dinb(n2441), .dout(n15194));
  jxor g15125(.dina(n15194), .dinb(n15186), .dout(n15195));
  jxor g15126(.dina(n15195), .dinb(n15051), .dout(n15196));
  jand g15127(.dina(n12284), .dinb(n3423), .dout(n15197));
  jand g15128(.dina(n12282), .dinb(n3569), .dout(n15198));
  jand g15129(.dina(n11798), .dinb(n3428), .dout(n15199));
  jand g15130(.dina(n11646), .dinb(n3210), .dout(n15200));
  jor  g15131(.dina(n15200), .dinb(n15199), .dout(n15201));
  jor  g15132(.dina(n15201), .dinb(n15198), .dout(n15202));
  jor  g15133(.dina(n15202), .dinb(n15197), .dout(n15203));
  jxor g15134(.dina(n15203), .dinb(n3473), .dout(n15204));
  jxor g15135(.dina(n15204), .dinb(n15196), .dout(n15205));
  jxor g15136(.dina(n15205), .dinb(n15047), .dout(n15206));
  jnot g15137(.din(n15206), .dout(n15207));
  jand g15138(.dina(n12671), .dinb(n4022), .dout(n15208));
  jand g15139(.dina(n12669), .dinb(n4220), .dout(n15209));
  jand g15140(.dina(n12536), .dinb(n4027), .dout(n15210));
  jand g15141(.dina(n12547), .dinb(n3870), .dout(n15211));
  jor  g15142(.dina(n15211), .dinb(n15210), .dout(n15212));
  jor  g15143(.dina(n15212), .dinb(n15209), .dout(n15213));
  jor  g15144(.dina(n15213), .dinb(n15208), .dout(n15214));
  jxor g15145(.dina(n15214), .dinb(n4050), .dout(n15215));
  jxor g15146(.dina(n15215), .dinb(n15207), .dout(n15216));
  jxor g15147(.dina(n15216), .dinb(n15041), .dout(n15217));
  jand g15148(.dina(n13627), .dinb(n4691), .dout(n15218));
  jand g15149(.dina(n13469), .dinb(n4941), .dout(n15219));
  jand g15150(.dina(n13478), .dinb(n4696), .dout(n15220));
  jand g15151(.dina(n13248), .dinb(n4701), .dout(n15221));
  jor  g15152(.dina(n15221), .dinb(n15220), .dout(n15222));
  jor  g15153(.dina(n15222), .dinb(n15219), .dout(n15223));
  jor  g15154(.dina(n15223), .dinb(n15218), .dout(n15224));
  jxor g15155(.dina(n15224), .dinb(n4713), .dout(n15225));
  jxor g15156(.dina(n15225), .dinb(n15217), .dout(n15226));
  jxor g15157(.dina(n15226), .dinb(n15035), .dout(n15227));
  jand g15158(.dina(n14579), .dinb(n5280), .dout(n15228));
  jand g15159(.dina(n14249), .dinb(n5531), .dout(n15229));
  jand g15160(.dina(n14448), .dinb(n5814), .dout(n15230));
  jor  g15161(.dina(n15230), .dinb(n15229), .dout(n15231));
  jand g15162(.dina(n13614), .dinb(n5536), .dout(n15232));
  jor  g15163(.dina(n15232), .dinb(n15231), .dout(n15233));
  jor  g15164(.dina(n15233), .dinb(n15228), .dout(n15234));
  jxor g15165(.dina(n15234), .dinb(n5277), .dout(n15235));
  jxor g15166(.dina(n15235), .dinb(n15227), .dout(n15236));
  jxor g15167(.dina(n15236), .dinb(n15030), .dout(n15237));
  jand g15168(.dina(n14549), .dinb(n14447), .dout(n15238));
  jand g15169(.dina(n14550), .dinb(n14459), .dout(n15239));
  jor  g15170(.dina(n15239), .dinb(n15238), .dout(n15240));
  jand g15171(.dina(n14526), .dinb(n14462), .dout(n15241));
  jand g15172(.dina(n14446), .dinb(n14363), .dout(n15242));
  jor  g15173(.dina(n15242), .dinb(n14529), .dout(n15243));
  jand g15174(.dina(n15243), .dinb(n14527), .dout(n15244));
  jor  g15175(.dina(n15244), .dinb(n15241), .dout(n15245));
  jand g15176(.dina(n14517), .dinb(n14465), .dout(n15246));
  jnot g15177(.din(n15246), .dout(n15247));
  jor  g15178(.dina(n14525), .dinb(n14519), .dout(n15248));
  jand g15179(.dina(n15248), .dinb(n15247), .dout(n15249));
  jnot g15180(.din(n15249), .dout(n15250));
  jor  g15181(.dina(n7682), .dinb(n7061), .dout(n15251));
  jand g15182(.dina(n7629), .dinb(n5082), .dout(n15252));
  jand g15183(.dina(n7935), .dinb(n5084), .dout(n15253));
  jor  g15184(.dina(n15253), .dinb(n15252), .dout(n15254));
  jand g15185(.dina(n7218), .dinb(n6050), .dout(n15255));
  jor  g15186(.dina(n15255), .dinb(n15254), .dout(n15256));
  jnot g15187(.din(n15256), .dout(n15257));
  jand g15188(.dina(n15257), .dinb(n15251), .dout(n15258));
  jand g15189(.dina(n8256), .dinb(n2936), .dout(n15259));
  jor  g15190(.dina(n15259), .dinb(n3684), .dout(n15260));
  jand g15191(.dina(n15260), .dinb(n8000), .dout(n15261));
  jxor g15192(.dina(n15261), .dinb(n93), .dout(n15262));
  jxor g15193(.dina(n15262), .dinb(n15258), .dout(n15263));
  jnot g15194(.din(n14431), .dout(n15264));
  jand g15195(.dina(n14514), .dinb(n15264), .dout(n15265));
  jand g15196(.dina(n14516), .dinb(n14474), .dout(n15266));
  jor  g15197(.dina(n15266), .dinb(n15265), .dout(n15267));
  jand g15198(.dina(n6169), .dinb(n1762), .dout(n15268));
  jand g15199(.dina(n447), .dinb(n511), .dout(n15269));
  jand g15200(.dina(n15269), .dinb(n1291), .dout(n15270));
  jand g15201(.dina(n15270), .dinb(n1682), .dout(n15271));
  jand g15202(.dina(n15271), .dinb(n15268), .dout(n15272));
  jand g15203(.dina(n2100), .dinb(n1559), .dout(n15273));
  jand g15204(.dina(n931), .dinb(n534), .dout(n15274));
  jand g15205(.dina(n15274), .dinb(n15273), .dout(n15275));
  jand g15206(.dina(n15275), .dinb(n5171), .dout(n15276));
  jand g15207(.dina(n15276), .dinb(n175), .dout(n15277));
  jand g15208(.dina(n15277), .dinb(n15272), .dout(n15278));
  jand g15209(.dina(n2445), .dinb(n1167), .dout(n15279));
  jand g15210(.dina(n15279), .dinb(n15278), .dout(n15280));
  jand g15211(.dina(n1107), .dinb(n881), .dout(n15281));
  jand g15212(.dina(n15281), .dinb(n1778), .dout(n15282));
  jand g15213(.dina(n1867), .dinb(n965), .dout(n15283));
  jand g15214(.dina(n15283), .dinb(n135), .dout(n15284));
  jand g15215(.dina(n15284), .dinb(n15282), .dout(n15285));
  jand g15216(.dina(n13544), .dinb(n713), .dout(n15286));
  jand g15217(.dina(n10384), .dinb(n2529), .dout(n15287));
  jand g15218(.dina(n15287), .dinb(n15286), .dout(n15288));
  jand g15219(.dina(n15288), .dinb(n15285), .dout(n15289));
  jand g15220(.dina(n15289), .dinb(n4007), .dout(n15290));
  jand g15221(.dina(n4012), .dinb(n1367), .dout(n15291));
  jand g15222(.dina(n15291), .dinb(n1449), .dout(n15292));
  jand g15223(.dina(n15292), .dinb(n15290), .dout(n15293));
  jand g15224(.dina(n1713), .dinb(n645), .dout(n15294));
  jand g15225(.dina(n15294), .dinb(n10739), .dout(n15295));
  jand g15226(.dina(n15295), .dinb(n519), .dout(n15296));
  jand g15227(.dina(n15296), .dinb(n4494), .dout(n15297));
  jand g15228(.dina(n470), .dinb(n1431), .dout(n15298));
  jand g15229(.dina(n3758), .dinb(n555), .dout(n15299));
  jand g15230(.dina(n15299), .dinb(n15298), .dout(n15300));
  jand g15231(.dina(n4422), .dinb(n2052), .dout(n15301));
  jand g15232(.dina(n1361), .dinb(n1738), .dout(n15302));
  jand g15233(.dina(n15302), .dinb(n1462), .dout(n15303));
  jand g15234(.dina(n15303), .dinb(n15301), .dout(n15304));
  jand g15235(.dina(n15304), .dinb(n3163), .dout(n15305));
  jand g15236(.dina(n15305), .dinb(n15300), .dout(n15306));
  jand g15237(.dina(n15306), .dinb(n15297), .dout(n15307));
  jand g15238(.dina(n15307), .dinb(n15293), .dout(n15308));
  jand g15239(.dina(n15308), .dinb(n15280), .dout(n15309));
  jand g15240(.dina(n15309), .dinb(n1406), .dout(n15310));
  jxor g15241(.dina(n15310), .dinb(n14515), .dout(n15311));
  jxor g15242(.dina(n15311), .dinb(n15267), .dout(n15312));
  jxor g15243(.dina(n15312), .dinb(n15263), .dout(n15313));
  jxor g15244(.dina(n15313), .dinb(n15250), .dout(n15314));
  jxor g15245(.dina(n15314), .dinb(n15245), .dout(n15315));
  jxor g15246(.dina(n15315), .dinb(n14549), .dout(n15316));
  jxor g15247(.dina(n15316), .dinb(n15240), .dout(n15317));
  jand g15248(.dina(n15317), .dinb(n6495), .dout(n15318));
  jand g15249(.dina(n15315), .dinb(n6503), .dout(n15319));
  jand g15250(.dina(n14549), .dinb(n6506), .dout(n15320));
  jand g15251(.dina(n14447), .dinb(n6500), .dout(n15321));
  jor  g15252(.dina(n15321), .dinb(n15320), .dout(n15322));
  jor  g15253(.dina(n15322), .dinb(n15319), .dout(n15323));
  jor  g15254(.dina(n15323), .dinb(n15318), .dout(n15324));
  jxor g15255(.dina(n15324), .dinb(n6219), .dout(n15325));
  jxor g15256(.dina(n15325), .dinb(n15237), .dout(n15326));
  jxor g15257(.dina(n15326), .dinb(n15026), .dout(n15327));
  jxor g15258(.dina(n15327), .dinb(n15022), .dout(n15328));
  jnot g15259(.din(n15328), .dout(n15329));
  jand g15260(.dina(n15329), .dinb(n71), .dout(n15330));
  jand g15261(.dina(n15020), .dinb(n731), .dout(n15331));
  jand g15262(.dina(n15327), .dinb(n796), .dout(n15332));
  jor  g15263(.dina(n15332), .dinb(n15331), .dout(n15333));
  jor  g15264(.dina(n15333), .dinb(n15330), .dout(n15334));
  jnot g15265(.din(n15334), .dout(n15335));
  jand g15266(.dina(n15020), .dinb(n67), .dout(n15336));
  jnot g15267(.din(n15336), .dout(n15337));
  jand g15268(.dina(n15337), .dinb(\a[26] ), .dout(n15338));
  jand g15269(.dina(n15338), .dinb(n15335), .dout(n15339));
  jand g15270(.dina(n15327), .dinb(n15022), .dout(n15340));
  jor  g15271(.dina(n15325), .dinb(n15237), .dout(n15341));
  jnot g15272(.din(n15341), .dout(n15342));
  jand g15273(.dina(n15326), .dinb(n15026), .dout(n15343));
  jor  g15274(.dina(n15343), .dinb(n15342), .dout(n15344));
  jor  g15275(.dina(n15235), .dinb(n15227), .dout(n15345));
  jnot g15276(.din(n15236), .dout(n15346));
  jor  g15277(.dina(n15346), .dinb(n15030), .dout(n15347));
  jand g15278(.dina(n15347), .dinb(n15345), .dout(n15348));
  jnot g15279(.din(n15217), .dout(n15349));
  jor  g15280(.dina(n15225), .dinb(n15349), .dout(n15350));
  jnot g15281(.din(n15035), .dout(n15351));
  jor  g15282(.dina(n15226), .dinb(n15351), .dout(n15352));
  jand g15283(.dina(n15352), .dinb(n15350), .dout(n15353));
  jor  g15284(.dina(n15215), .dinb(n15207), .dout(n15354));
  jand g15285(.dina(n15216), .dinb(n15041), .dout(n15355));
  jnot g15286(.din(n15355), .dout(n15356));
  jand g15287(.dina(n15356), .dinb(n15354), .dout(n15357));
  jnot g15288(.din(n15196), .dout(n15358));
  jor  g15289(.dina(n15204), .dinb(n15358), .dout(n15359));
  jnot g15290(.din(n15047), .dout(n15360));
  jnot g15291(.din(n15205), .dout(n15361));
  jand g15292(.dina(n15361), .dinb(n15360), .dout(n15362));
  jnot g15293(.din(n15362), .dout(n15363));
  jand g15294(.dina(n15363), .dinb(n15359), .dout(n15364));
  jor  g15295(.dina(n15194), .dinb(n15186), .dout(n15365));
  jnot g15296(.din(n15365), .dout(n15366));
  jand g15297(.dina(n15195), .dinb(n15051), .dout(n15367));
  jor  g15298(.dina(n15367), .dinb(n15366), .dout(n15368));
  jor  g15299(.dina(n15183), .dinb(n15175), .dout(n15369));
  jand g15300(.dina(n15184), .dinb(n15056), .dout(n15370));
  jnot g15301(.din(n15370), .dout(n15371));
  jand g15302(.dina(n15371), .dinb(n15369), .dout(n15372));
  jnot g15303(.din(n15372), .dout(n15373));
  jor  g15304(.dina(n15172), .dinb(n15164), .dout(n15374));
  jand g15305(.dina(n15173), .dinb(n15061), .dout(n15375));
  jnot g15306(.din(n15375), .dout(n15376));
  jand g15307(.dina(n15376), .dinb(n15374), .dout(n15377));
  jnot g15308(.din(n15377), .dout(n15378));
  jor  g15309(.dina(n15161), .dinb(n15153), .dout(n15379));
  jand g15310(.dina(n15162), .dinb(n15066), .dout(n15380));
  jnot g15311(.din(n15380), .dout(n15381));
  jand g15312(.dina(n15381), .dinb(n15379), .dout(n15382));
  jnot g15313(.din(n15382), .dout(n15383));
  jor  g15314(.dina(n15150), .dinb(n15142), .dout(n15384));
  jand g15315(.dina(n15151), .dinb(n15071), .dout(n15385));
  jnot g15316(.din(n15385), .dout(n15386));
  jand g15317(.dina(n15386), .dinb(n15384), .dout(n15387));
  jnot g15318(.din(n15387), .dout(n15388));
  jor  g15319(.dina(n15139), .dinb(n15080), .dout(n15389));
  jand g15320(.dina(n15140), .dinb(n15078), .dout(n15390));
  jnot g15321(.din(n15390), .dout(n15391));
  jand g15322(.dina(n15391), .dinb(n15389), .dout(n15392));
  jnot g15323(.din(n15392), .dout(n15393));
  jand g15324(.dina(n10167), .dinb(n978), .dout(n15394));
  jand g15325(.dina(n15394), .dinb(n15278), .dout(n15395));
  jand g15326(.dina(n13195), .dinb(n1929), .dout(n15396));
  jand g15327(.dina(n15396), .dinb(n101), .dout(n15397));
  jand g15328(.dina(n15397), .dinb(n1460), .dout(n15398));
  jand g15329(.dina(n2529), .dinb(n1708), .dout(n15399));
  jand g15330(.dina(n15399), .dinb(n1334), .dout(n15400));
  jand g15331(.dina(n15400), .dinb(n15398), .dout(n15401));
  jand g15332(.dina(n15401), .dinb(n15395), .dout(n15402));
  jand g15333(.dina(n6426), .dinb(n1232), .dout(n15403));
  jand g15334(.dina(n15403), .dinb(n8103), .dout(n15404));
  jand g15335(.dina(n15404), .dinb(n14504), .dout(n15405));
  jand g15336(.dina(n15405), .dinb(n9742), .dout(n15406));
  jand g15337(.dina(n15406), .dinb(n15402), .dout(n15407));
  jnot g15338(.din(n15407), .dout(n15408));
  jand g15339(.dina(n8029), .dinb(n5076), .dout(n15409));
  jand g15340(.dina(n8022), .dinb(n5084), .dout(n15410));
  jand g15341(.dina(n7313), .dinb(n6050), .dout(n15411));
  jand g15342(.dina(n7692), .dinb(n5082), .dout(n15412));
  jor  g15343(.dina(n15412), .dinb(n15411), .dout(n15413));
  jor  g15344(.dina(n15413), .dinb(n15410), .dout(n15414));
  jor  g15345(.dina(n15414), .dinb(n15409), .dout(n15415));
  jxor g15346(.dina(n15415), .dinb(n15408), .dout(n15416));
  jxor g15347(.dina(n15416), .dinb(n15393), .dout(n15417));
  jnot g15348(.din(n15417), .dout(n15418));
  jand g15349(.dina(n8950), .dinb(n2936), .dout(n15419));
  jand g15350(.dina(n8740), .dinb(n2940), .dout(n15420));
  jand g15351(.dina(n8723), .dinb(n2943), .dout(n15421));
  jor  g15352(.dina(n15421), .dinb(n15420), .dout(n15422));
  jand g15353(.dina(n8268), .dinb(n3684), .dout(n15423));
  jor  g15354(.dina(n15423), .dinb(n15422), .dout(n15424));
  jor  g15355(.dina(n15424), .dinb(n15419), .dout(n15425));
  jxor g15356(.dina(n15425), .dinb(n93), .dout(n15426));
  jxor g15357(.dina(n15426), .dinb(n15418), .dout(n15427));
  jxor g15358(.dina(n15427), .dinb(n15388), .dout(n15428));
  jnot g15359(.din(n15428), .dout(n15429));
  jand g15360(.dina(n9898), .dinb(n71), .dout(n15430));
  jand g15361(.dina(n9656), .dinb(n796), .dout(n15431));
  jand g15362(.dina(n9250), .dinb(n731), .dout(n15432));
  jand g15363(.dina(n8936), .dinb(n1806), .dout(n15433));
  jor  g15364(.dina(n15433), .dinb(n15432), .dout(n15434));
  jor  g15365(.dina(n15434), .dinb(n15431), .dout(n15435));
  jor  g15366(.dina(n15435), .dinb(n15430), .dout(n15436));
  jxor g15367(.dina(n15436), .dinb(n77), .dout(n15437));
  jxor g15368(.dina(n15437), .dinb(n15429), .dout(n15438));
  jxor g15369(.dina(n15438), .dinb(n15383), .dout(n15439));
  jnot g15370(.din(n15439), .dout(n15440));
  jand g15371(.dina(n10307), .dinb(n806), .dout(n15441));
  jand g15372(.dina(n10305), .dinb(n1620), .dout(n15442));
  jand g15373(.dina(n9872), .dinb(n1612), .dout(n15443));
  jand g15374(.dina(n9655), .dinb(n1644), .dout(n15444));
  jor  g15375(.dina(n15444), .dinb(n15443), .dout(n15445));
  jor  g15376(.dina(n15445), .dinb(n15442), .dout(n15446));
  jor  g15377(.dina(n15446), .dinb(n15441), .dout(n15447));
  jxor g15378(.dina(n15447), .dinb(n65), .dout(n15448));
  jxor g15379(.dina(n15448), .dinb(n15440), .dout(n15449));
  jxor g15380(.dina(n15449), .dinb(n15378), .dout(n15450));
  jnot g15381(.din(n15450), .dout(n15451));
  jand g15382(.dina(n10838), .dinb(n1819), .dout(n15452));
  jand g15383(.dina(n10640), .dinb(n2180), .dout(n15453));
  jand g15384(.dina(n10836), .dinb(n2243), .dout(n15454));
  jor  g15385(.dina(n15454), .dinb(n15453), .dout(n15455));
  jand g15386(.dina(n10647), .dinb(n2185), .dout(n15456));
  jor  g15387(.dina(n15456), .dinb(n15455), .dout(n15457));
  jor  g15388(.dina(n15457), .dinb(n15452), .dout(n15458));
  jxor g15389(.dina(n15458), .dinb(n2196), .dout(n15459));
  jxor g15390(.dina(n15459), .dinb(n15451), .dout(n15460));
  jxor g15391(.dina(n15460), .dinb(n15373), .dout(n15461));
  jand g15392(.dina(n11812), .dinb(n2743), .dout(n15462));
  jand g15393(.dina(n11646), .dinb(n2752), .dout(n15463));
  jand g15394(.dina(n11647), .dinb(n2748), .dout(n15464));
  jand g15395(.dina(n11306), .dinb(n2757), .dout(n15465));
  jor  g15396(.dina(n15465), .dinb(n15464), .dout(n15466));
  jor  g15397(.dina(n15466), .dinb(n15463), .dout(n15467));
  jor  g15398(.dina(n15467), .dinb(n15462), .dout(n15468));
  jxor g15399(.dina(n15468), .dinb(\a[17] ), .dout(n15469));
  jxor g15400(.dina(n15469), .dinb(n15461), .dout(n15470));
  jxor g15401(.dina(n15470), .dinb(n15368), .dout(n15471));
  jand g15402(.dina(n12696), .dinb(n3423), .dout(n15472));
  jand g15403(.dina(n12547), .dinb(n3569), .dout(n15473));
  jand g15404(.dina(n12282), .dinb(n3428), .dout(n15474));
  jand g15405(.dina(n11798), .dinb(n3210), .dout(n15475));
  jor  g15406(.dina(n15475), .dinb(n15474), .dout(n15476));
  jor  g15407(.dina(n15476), .dinb(n15473), .dout(n15477));
  jor  g15408(.dina(n15477), .dinb(n15472), .dout(n15478));
  jxor g15409(.dina(n15478), .dinb(n3473), .dout(n15479));
  jxor g15410(.dina(n15479), .dinb(n15471), .dout(n15480));
  jnot g15411(.din(n15480), .dout(n15481));
  jxor g15412(.dina(n15481), .dinb(n15364), .dout(n15482));
  jand g15413(.dina(n13250), .dinb(n4022), .dout(n15483));
  jand g15414(.dina(n12669), .dinb(n4027), .dout(n15484));
  jand g15415(.dina(n13248), .dinb(n4220), .dout(n15485));
  jor  g15416(.dina(n15485), .dinb(n15484), .dout(n15486));
  jand g15417(.dina(n12536), .dinb(n3870), .dout(n15487));
  jor  g15418(.dina(n15487), .dinb(n15486), .dout(n15488));
  jor  g15419(.dina(n15488), .dinb(n15483), .dout(n15489));
  jxor g15420(.dina(n15489), .dinb(n4050), .dout(n15490));
  jxor g15421(.dina(n15490), .dinb(n15482), .dout(n15491));
  jxor g15422(.dina(n15491), .dinb(n15357), .dout(n15492));
  jand g15423(.dina(n13616), .dinb(n4691), .dout(n15493));
  jand g15424(.dina(n13469), .dinb(n4696), .dout(n15494));
  jand g15425(.dina(n13614), .dinb(n4941), .dout(n15495));
  jor  g15426(.dina(n15495), .dinb(n15494), .dout(n15496));
  jand g15427(.dina(n13478), .dinb(n4701), .dout(n15497));
  jor  g15428(.dina(n15497), .dinb(n15496), .dout(n15498));
  jor  g15429(.dina(n15498), .dinb(n15493), .dout(n15499));
  jxor g15430(.dina(n15499), .dinb(n4713), .dout(n15500));
  jxor g15431(.dina(n15500), .dinb(n15492), .dout(n15501));
  jxor g15432(.dina(n15501), .dinb(n15353), .dout(n15502));
  jand g15433(.dina(n14562), .dinb(n5280), .dout(n15503));
  jand g15434(.dina(n14447), .dinb(n5814), .dout(n15504));
  jand g15435(.dina(n14448), .dinb(n5531), .dout(n15505));
  jand g15436(.dina(n14249), .dinb(n5536), .dout(n15506));
  jor  g15437(.dina(n15506), .dinb(n15505), .dout(n15507));
  jor  g15438(.dina(n15507), .dinb(n15504), .dout(n15508));
  jor  g15439(.dina(n15508), .dinb(n15503), .dout(n15509));
  jxor g15440(.dina(n15509), .dinb(n5277), .dout(n15510));
  jxor g15441(.dina(n15510), .dinb(n15502), .dout(n15511));
  jxor g15442(.dina(n15511), .dinb(n15348), .dout(n15512));
  jand g15443(.dina(n15315), .dinb(n14549), .dout(n15513));
  jand g15444(.dina(n15316), .dinb(n15240), .dout(n15514));
  jor  g15445(.dina(n15514), .dinb(n15513), .dout(n15515));
  jand g15446(.dina(n15313), .dinb(n15250), .dout(n15516));
  jand g15447(.dina(n15314), .dinb(n15245), .dout(n15517));
  jor  g15448(.dina(n15517), .dinb(n15516), .dout(n15518));
  jor  g15449(.dina(n15262), .dinb(n15258), .dout(n15519));
  jand g15450(.dina(n15312), .dinb(n15263), .dout(n15520));
  jnot g15451(.din(n15520), .dout(n15521));
  jand g15452(.dina(n15521), .dinb(n15519), .dout(n15522));
  jnot g15453(.din(n15522), .dout(n15523));
  jand g15454(.dina(n8014), .dinb(n5076), .dout(n15524));
  jand g15455(.dina(n7629), .dinb(n6050), .dout(n15525));
  jand g15456(.dina(n7935), .dinb(n5082), .dout(n15528));
  jor  g15457(.dina(n15528), .dinb(n15525), .dout(n15529));
  jor  g15458(.dina(n15529), .dinb(n15524), .dout(n15530));
  jand g15459(.dina(n10699), .dinb(n7102), .dout(n15531));
  jand g15460(.dina(n15531), .dinb(n6454), .dout(n15532));
  jand g15461(.dina(n3066), .dinb(n1511), .dout(n15533));
  jand g15462(.dina(n15533), .dinb(n3847), .dout(n15534));
  jand g15463(.dina(n15534), .dinb(n1016), .dout(n15535));
  jand g15464(.dina(n15535), .dinb(n7272), .dout(n15536));
  jand g15465(.dina(n3179), .dinb(n555), .dout(n15537));
  jand g15466(.dina(n15537), .dinb(n6462), .dout(n15538));
  jand g15467(.dina(n14386), .dinb(n2080), .dout(n15539));
  jand g15468(.dina(n15539), .dinb(n2089), .dout(n15540));
  jand g15469(.dina(n6169), .dinb(n1903), .dout(n15541));
  jand g15470(.dina(n7287), .dinb(n4417), .dout(n15542));
  jand g15471(.dina(n15542), .dinb(n4528), .dout(n15543));
  jand g15472(.dina(n15543), .dinb(n15541), .dout(n15544));
  jand g15473(.dina(n15544), .dinb(n15540), .dout(n15545));
  jand g15474(.dina(n15545), .dinb(n7088), .dout(n15546));
  jand g15475(.dina(n15546), .dinb(n15538), .dout(n15547));
  jand g15476(.dina(n15547), .dinb(n15536), .dout(n15548));
  jand g15477(.dina(n15548), .dinb(n7261), .dout(n15549));
  jand g15478(.dina(n15549), .dinb(n15532), .dout(n15550));
  jand g15479(.dina(n15550), .dinb(n15310), .dout(n15551));
  jnot g15480(.din(n15551), .dout(n15552));
  jor  g15481(.dina(n15550), .dinb(n15310), .dout(n15553));
  jand g15482(.dina(n15553), .dinb(n93), .dout(n15554));
  jand g15483(.dina(n15554), .dinb(n15552), .dout(n15555));
  jnot g15484(.din(n15555), .dout(n15556));
  jand g15485(.dina(n15556), .dinb(n93), .dout(n15557));
  jand g15486(.dina(n15556), .dinb(n15553), .dout(n15558));
  jand g15487(.dina(n15558), .dinb(n15552), .dout(n15559));
  jor  g15488(.dina(n15559), .dinb(n15557), .dout(n15560));
  jand g15489(.dina(n15310), .dinb(n14515), .dout(n15561));
  jand g15490(.dina(n15311), .dinb(n15267), .dout(n15562));
  jor  g15491(.dina(n15562), .dinb(n15561), .dout(n15563));
  jxor g15492(.dina(n15563), .dinb(n15560), .dout(n15564));
  jxor g15493(.dina(n15564), .dinb(n15530), .dout(n15565));
  jxor g15494(.dina(n15565), .dinb(n15523), .dout(n15566));
  jxor g15495(.dina(n15566), .dinb(n15518), .dout(n15567));
  jxor g15496(.dina(n15567), .dinb(n15315), .dout(n15568));
  jxor g15497(.dina(n15568), .dinb(n15515), .dout(n15569));
  jand g15498(.dina(n15569), .dinb(n6495), .dout(n15570));
  jand g15499(.dina(n15567), .dinb(n6503), .dout(n15571));
  jand g15500(.dina(n15315), .dinb(n6506), .dout(n15572));
  jand g15501(.dina(n14549), .dinb(n6500), .dout(n15573));
  jor  g15502(.dina(n15573), .dinb(n15572), .dout(n15574));
  jor  g15503(.dina(n15574), .dinb(n15571), .dout(n15575));
  jor  g15504(.dina(n15575), .dinb(n15570), .dout(n15576));
  jxor g15505(.dina(n15576), .dinb(n6219), .dout(n15577));
  jxor g15506(.dina(n15577), .dinb(n15512), .dout(n15578));
  jxor g15507(.dina(n15578), .dinb(n15344), .dout(n15579));
  jxor g15508(.dina(n15579), .dinb(n15340), .dout(n15580));
  jand g15509(.dina(n15580), .dinb(n71), .dout(n15581));
  jand g15510(.dina(n15327), .dinb(n731), .dout(n15582));
  jor  g15511(.dina(n15582), .dinb(n15581), .dout(n15583));
  jand g15512(.dina(n15579), .dinb(n796), .dout(n15584));
  jand g15513(.dina(n15020), .dinb(n1806), .dout(n15585));
  jor  g15514(.dina(n15585), .dinb(n15584), .dout(n15586));
  jor  g15515(.dina(n15586), .dinb(n15583), .dout(n15587));
  jnot g15516(.din(n15587), .dout(n15588));
  jand g15517(.dina(n15588), .dinb(n15339), .dout(n15589));
  jxor g15518(.dina(n15589), .dinb(n15021), .dout(n15590));
  jnot g15519(.din(n15590), .dout(n15591));
  jor  g15520(.dina(n15577), .dinb(n15512), .dout(n15592));
  jnot g15521(.din(n15592), .dout(n15593));
  jand g15522(.dina(n15578), .dinb(n15344), .dout(n15594));
  jor  g15523(.dina(n15594), .dinb(n15593), .dout(n15595));
  jor  g15524(.dina(n15510), .dinb(n15502), .dout(n15596));
  jnot g15525(.din(n15511), .dout(n15597));
  jor  g15526(.dina(n15597), .dinb(n15348), .dout(n15598));
  jand g15527(.dina(n15598), .dinb(n15596), .dout(n15599));
  jor  g15528(.dina(n15500), .dinb(n15492), .dout(n15600));
  jnot g15529(.din(n15600), .dout(n15601));
  jnot g15530(.din(n15353), .dout(n15602));
  jand g15531(.dina(n15501), .dinb(n15602), .dout(n15603));
  jor  g15532(.dina(n15603), .dinb(n15601), .dout(n15604));
  jor  g15533(.dina(n15490), .dinb(n15482), .dout(n15605));
  jnot g15534(.din(n15491), .dout(n15606));
  jor  g15535(.dina(n15606), .dinb(n15357), .dout(n15607));
  jand g15536(.dina(n15607), .dinb(n15605), .dout(n15608));
  jnot g15537(.din(n15471), .dout(n15609));
  jor  g15538(.dina(n15479), .dinb(n15609), .dout(n15610));
  jor  g15539(.dina(n15480), .dinb(n15364), .dout(n15611));
  jand g15540(.dina(n15611), .dinb(n15610), .dout(n15612));
  jand g15541(.dina(n15469), .dinb(n15461), .dout(n15613));
  jand g15542(.dina(n15470), .dinb(n15368), .dout(n15614));
  jor  g15543(.dina(n15614), .dinb(n15613), .dout(n15615));
  jor  g15544(.dina(n15459), .dinb(n15451), .dout(n15616));
  jand g15545(.dina(n15460), .dinb(n15373), .dout(n15617));
  jnot g15546(.din(n15617), .dout(n15618));
  jand g15547(.dina(n15618), .dinb(n15616), .dout(n15619));
  jnot g15548(.din(n15619), .dout(n15620));
  jor  g15549(.dina(n15448), .dinb(n15440), .dout(n15621));
  jand g15550(.dina(n15449), .dinb(n15378), .dout(n15622));
  jnot g15551(.din(n15622), .dout(n15623));
  jand g15552(.dina(n15623), .dinb(n15621), .dout(n15624));
  jnot g15553(.din(n15624), .dout(n15625));
  jor  g15554(.dina(n15437), .dinb(n15429), .dout(n15626));
  jand g15555(.dina(n15438), .dinb(n15383), .dout(n15627));
  jnot g15556(.din(n15627), .dout(n15628));
  jand g15557(.dina(n15628), .dinb(n15626), .dout(n15629));
  jnot g15558(.din(n15629), .dout(n15630));
  jor  g15559(.dina(n15426), .dinb(n15418), .dout(n15631));
  jand g15560(.dina(n15427), .dinb(n15388), .dout(n15632));
  jnot g15561(.din(n15632), .dout(n15633));
  jand g15562(.dina(n15633), .dinb(n15631), .dout(n15634));
  jnot g15563(.din(n15634), .dout(n15635));
  jand g15564(.dina(n15415), .dinb(n15408), .dout(n15636));
  jand g15565(.dina(n15416), .dinb(n15393), .dout(n15637));
  jor  g15566(.dina(n15637), .dinb(n15636), .dout(n15638));
  jand g15567(.dina(n12219), .dinb(n5210), .dout(n15639));
  jand g15568(.dina(n11416), .dinb(n929), .dout(n15640));
  jand g15569(.dina(n15640), .dinb(n3752), .dout(n15641));
  jand g15570(.dina(n15641), .dinb(n15639), .dout(n15642));
  jand g15571(.dina(n1682), .dinb(n179), .dout(n15643));
  jand g15572(.dina(n15643), .dinb(n2036), .dout(n15644));
  jand g15573(.dina(n917), .dinb(n901), .dout(n15645));
  jand g15574(.dina(n15645), .dinb(n3108), .dout(n15646));
  jand g15575(.dina(n15646), .dinb(n1498), .dout(n15647));
  jand g15576(.dina(n15647), .dinb(n1238), .dout(n15648));
  jand g15577(.dina(n15648), .dinb(n15644), .dout(n15649));
  jand g15578(.dina(n15649), .dinb(n15642), .dout(n15650));
  jand g15579(.dina(n9756), .dinb(n1317), .dout(n15651));
  jand g15580(.dina(n1096), .dinb(n1310), .dout(n15652));
  jand g15581(.dina(n15652), .dinb(n15651), .dout(n15653));
  jand g15582(.dina(n15653), .dinb(n6312), .dout(n15654));
  jnot g15583(.din(n969), .dout(n15655));
  jand g15584(.dina(n1090), .dinb(n664), .dout(n15656));
  jand g15585(.dina(n15656), .dinb(n15655), .dout(n15657));
  jand g15586(.dina(n15657), .dinb(n700), .dout(n15658));
  jand g15587(.dina(n15658), .dinb(n7639), .dout(n15659));
  jand g15588(.dina(n15659), .dinb(n15654), .dout(n15660));
  jand g15589(.dina(n542), .dinb(n1272), .dout(n15661));
  jand g15590(.dina(n15661), .dinb(n15660), .dout(n15662));
  jand g15591(.dina(n1861), .dinb(n1765), .dout(n15663));
  jand g15592(.dina(n447), .dinb(n1205), .dout(n15664));
  jand g15593(.dina(n452), .dinb(n838), .dout(n15665));
  jand g15594(.dina(n15665), .dinb(n1582), .dout(n15666));
  jand g15595(.dina(n15666), .dinb(n15664), .dout(n15667));
  jand g15596(.dina(n1228), .dinb(n428), .dout(n15668));
  jand g15597(.dina(n15668), .dinb(n100), .dout(n15669));
  jand g15598(.dina(n15669), .dinb(n15667), .dout(n15670));
  jand g15599(.dina(n15670), .dinb(n15663), .dout(n15671));
  jand g15600(.dina(n808), .dinb(n92), .dout(n15672));
  jand g15601(.dina(n15672), .dinb(n1709), .dout(n15673));
  jand g15602(.dina(n15673), .dinb(n1098), .dout(n15674));
  jand g15603(.dina(n696), .dinb(n1346), .dout(n15675));
  jand g15604(.dina(n15675), .dinb(n13395), .dout(n15676));
  jand g15605(.dina(n15676), .dinb(n15674), .dout(n15677));
  jand g15606(.dina(n15677), .dinb(n15671), .dout(n15678));
  jand g15607(.dina(n15678), .dinb(n15662), .dout(n15679));
  jand g15608(.dina(n15679), .dinb(n3342), .dout(n15680));
  jand g15609(.dina(n15680), .dinb(n15650), .dout(n15681));
  jnot g15610(.din(n15681), .dout(n15682));
  jand g15611(.dina(n8270), .dinb(n5076), .dout(n15683));
  jand g15612(.dina(n8268), .dinb(n5084), .dout(n15684));
  jand g15613(.dina(n7692), .dinb(n6050), .dout(n15685));
  jand g15614(.dina(n8022), .dinb(n5082), .dout(n15686));
  jor  g15615(.dina(n15686), .dinb(n15685), .dout(n15687));
  jor  g15616(.dina(n15687), .dinb(n15684), .dout(n15688));
  jor  g15617(.dina(n15688), .dinb(n15683), .dout(n15689));
  jxor g15618(.dina(n15689), .dinb(n15682), .dout(n15690));
  jxor g15619(.dina(n15690), .dinb(n15638), .dout(n15691));
  jnot g15620(.din(n15691), .dout(n15692));
  jand g15621(.dina(n8938), .dinb(n2936), .dout(n15693));
  jand g15622(.dina(n8723), .dinb(n2940), .dout(n15694));
  jand g15623(.dina(n8936), .dinb(n2943), .dout(n15695));
  jor  g15624(.dina(n15695), .dinb(n15694), .dout(n15696));
  jand g15625(.dina(n8740), .dinb(n3684), .dout(n15697));
  jor  g15626(.dina(n15697), .dinb(n15696), .dout(n15698));
  jor  g15627(.dina(n15698), .dinb(n15693), .dout(n15699));
  jxor g15628(.dina(n15699), .dinb(n93), .dout(n15700));
  jxor g15629(.dina(n15700), .dinb(n15692), .dout(n15701));
  jxor g15630(.dina(n15701), .dinb(n15635), .dout(n15702));
  jnot g15631(.din(n15702), .dout(n15703));
  jand g15632(.dina(n9886), .dinb(n71), .dout(n15704));
  jand g15633(.dina(n9655), .dinb(n796), .dout(n15705));
  jand g15634(.dina(n9656), .dinb(n731), .dout(n15706));
  jand g15635(.dina(n9250), .dinb(n1806), .dout(n15707));
  jor  g15636(.dina(n15707), .dinb(n15706), .dout(n15708));
  jor  g15637(.dina(n15708), .dinb(n15705), .dout(n15709));
  jor  g15638(.dina(n15709), .dinb(n15704), .dout(n15710));
  jxor g15639(.dina(n15710), .dinb(n77), .dout(n15711));
  jxor g15640(.dina(n15711), .dinb(n15703), .dout(n15712));
  jxor g15641(.dina(n15712), .dinb(n15630), .dout(n15713));
  jnot g15642(.din(n15713), .dout(n15714));
  jand g15643(.dina(n10862), .dinb(n806), .dout(n15715));
  jand g15644(.dina(n10305), .dinb(n1612), .dout(n15716));
  jand g15645(.dina(n10647), .dinb(n1620), .dout(n15717));
  jor  g15646(.dina(n15717), .dinb(n15716), .dout(n15718));
  jand g15647(.dina(n9872), .dinb(n1644), .dout(n15719));
  jor  g15648(.dina(n15719), .dinb(n15718), .dout(n15720));
  jor  g15649(.dina(n15720), .dinb(n15715), .dout(n15721));
  jxor g15650(.dina(n15721), .dinb(n65), .dout(n15722));
  jxor g15651(.dina(n15722), .dinb(n15714), .dout(n15723));
  jxor g15652(.dina(n15723), .dinb(n15625), .dout(n15724));
  jnot g15653(.din(n15724), .dout(n15725));
  jand g15654(.dina(n11308), .dinb(n1819), .dout(n15726));
  jand g15655(.dina(n11306), .dinb(n2243), .dout(n15727));
  jand g15656(.dina(n10836), .dinb(n2180), .dout(n15728));
  jand g15657(.dina(n10640), .dinb(n2185), .dout(n15729));
  jor  g15658(.dina(n15729), .dinb(n15728), .dout(n15730));
  jor  g15659(.dina(n15730), .dinb(n15727), .dout(n15731));
  jor  g15660(.dina(n15731), .dinb(n15726), .dout(n15732));
  jxor g15661(.dina(n15732), .dinb(n2196), .dout(n15733));
  jxor g15662(.dina(n15733), .dinb(n15725), .dout(n15734));
  jxor g15663(.dina(n15734), .dinb(n15620), .dout(n15735));
  jnot g15664(.din(n15735), .dout(n15736));
  jand g15665(.dina(n11800), .dinb(n2743), .dout(n15737));
  jand g15666(.dina(n11798), .dinb(n2752), .dout(n15738));
  jand g15667(.dina(n11646), .dinb(n2748), .dout(n15739));
  jand g15668(.dina(n11647), .dinb(n2757), .dout(n15740));
  jor  g15669(.dina(n15740), .dinb(n15739), .dout(n15741));
  jor  g15670(.dina(n15741), .dinb(n15738), .dout(n15742));
  jor  g15671(.dina(n15742), .dinb(n15737), .dout(n15743));
  jxor g15672(.dina(n15743), .dinb(n2441), .dout(n15744));
  jxor g15673(.dina(n15744), .dinb(n15736), .dout(n15745));
  jxor g15674(.dina(n15745), .dinb(n15615), .dout(n15746));
  jand g15675(.dina(n12684), .dinb(n3423), .dout(n15747));
  jand g15676(.dina(n12536), .dinb(n3569), .dout(n15748));
  jand g15677(.dina(n12547), .dinb(n3428), .dout(n15749));
  jand g15678(.dina(n12282), .dinb(n3210), .dout(n15750));
  jor  g15679(.dina(n15750), .dinb(n15749), .dout(n15751));
  jor  g15680(.dina(n15751), .dinb(n15748), .dout(n15752));
  jor  g15681(.dina(n15752), .dinb(n15747), .dout(n15753));
  jxor g15682(.dina(n15753), .dinb(n3473), .dout(n15754));
  jxor g15683(.dina(n15754), .dinb(n15746), .dout(n15755));
  jxor g15684(.dina(n15755), .dinb(n15612), .dout(n15756));
  jand g15685(.dina(n13639), .dinb(n4022), .dout(n15757));
  jand g15686(.dina(n13248), .dinb(n4027), .dout(n15758));
  jand g15687(.dina(n13478), .dinb(n4220), .dout(n15759));
  jor  g15688(.dina(n15759), .dinb(n15758), .dout(n15760));
  jand g15689(.dina(n12669), .dinb(n3870), .dout(n15761));
  jor  g15690(.dina(n15761), .dinb(n15760), .dout(n15762));
  jor  g15691(.dina(n15762), .dinb(n15757), .dout(n15763));
  jxor g15692(.dina(n15763), .dinb(n4050), .dout(n15764));
  jxor g15693(.dina(n15764), .dinb(n15756), .dout(n15765));
  jnot g15694(.din(n15765), .dout(n15766));
  jxor g15695(.dina(n15766), .dinb(n15608), .dout(n15767));
  jand g15696(.dina(n14251), .dinb(n4691), .dout(n15768));
  jand g15697(.dina(n14249), .dinb(n4941), .dout(n15769));
  jand g15698(.dina(n13614), .dinb(n4696), .dout(n15770));
  jand g15699(.dina(n13469), .dinb(n4701), .dout(n15771));
  jor  g15700(.dina(n15771), .dinb(n15770), .dout(n15772));
  jor  g15701(.dina(n15772), .dinb(n15769), .dout(n15773));
  jor  g15702(.dina(n15773), .dinb(n15768), .dout(n15774));
  jxor g15703(.dina(n15774), .dinb(n4713), .dout(n15775));
  jxor g15704(.dina(n15775), .dinb(n15767), .dout(n15776));
  jxor g15705(.dina(n15776), .dinb(n15604), .dout(n15777));
  jand g15706(.dina(n14551), .dinb(n5280), .dout(n15778));
  jand g15707(.dina(n14549), .dinb(n5814), .dout(n15779));
  jand g15708(.dina(n14447), .dinb(n5531), .dout(n15780));
  jand g15709(.dina(n14448), .dinb(n5536), .dout(n15781));
  jor  g15710(.dina(n15781), .dinb(n15780), .dout(n15782));
  jor  g15711(.dina(n15782), .dinb(n15779), .dout(n15783));
  jor  g15712(.dina(n15783), .dinb(n15778), .dout(n15784));
  jxor g15713(.dina(n15784), .dinb(\a[5] ), .dout(n15785));
  jxor g15714(.dina(n15785), .dinb(n15777), .dout(n15786));
  jxor g15715(.dina(n15786), .dinb(n15599), .dout(n15787));
  jand g15716(.dina(n15567), .dinb(n15315), .dout(n15788));
  jand g15717(.dina(n15568), .dinb(n15515), .dout(n15789));
  jor  g15718(.dina(n15789), .dinb(n15788), .dout(n15790));
  jand g15719(.dina(n15563), .dinb(n15560), .dout(n15791));
  jand g15720(.dina(n15564), .dinb(n15530), .dout(n15792));
  jor  g15721(.dina(n15792), .dinb(n15791), .dout(n15793));
  jor  g15722(.dina(n8260), .dinb(n7061), .dout(n15794));
  jand g15723(.dina(n8000), .dinb(n5082), .dout(n15796));
  jnot g15724(.din(n15796), .dout(n15798));
  jand g15725(.dina(n15798), .dinb(n15794), .dout(n15799));
  jnot g15726(.din(n15799), .dout(n15800));
  jand g15727(.dina(n7266), .dinb(n6183), .dout(n15801));
  jand g15728(.dina(n15536), .dinb(n1261), .dout(n15802));
  jand g15729(.dina(n15802), .dinb(n132), .dout(n15803));
  jand g15730(.dina(n7982), .dinb(n697), .dout(n15804));
  jand g15731(.dina(n6449), .dinb(n1883), .dout(n15805));
  jand g15732(.dina(n15805), .dinb(n270), .dout(n15806));
  jand g15733(.dina(n15806), .dinb(n7643), .dout(n15807));
  jand g15734(.dina(n15807), .dinb(n15804), .dout(n15808));
  jand g15735(.dina(n15808), .dinb(n9562), .dout(n15809));
  jand g15736(.dina(n15809), .dinb(n15803), .dout(n15810));
  jand g15737(.dina(n15810), .dinb(n15801), .dout(n15811));
  jnot g15738(.din(n15811), .dout(n15812));
  jxor g15739(.dina(n15812), .dinb(n15558), .dout(n15813));
  jxor g15740(.dina(n15813), .dinb(n15800), .dout(n15814));
  jxor g15741(.dina(n15814), .dinb(n15793), .dout(n15815));
  jnot g15742(.din(n15815), .dout(n15816));
  jand g15743(.dina(n15565), .dinb(n15523), .dout(n15817));
  jnot g15744(.din(n15817), .dout(n15818));
  jnot g15745(.din(n15516), .dout(n15819));
  jnot g15746(.din(n15241), .dout(n15820));
  jor  g15747(.dina(n14548), .dinb(n14528), .dout(n15821));
  jand g15748(.dina(n15821), .dinb(n15820), .dout(n15822));
  jnot g15749(.din(n15314), .dout(n15823));
  jor  g15750(.dina(n15823), .dinb(n15822), .dout(n15824));
  jand g15751(.dina(n15824), .dinb(n15819), .dout(n15825));
  jnot g15752(.din(n15566), .dout(n15826));
  jor  g15753(.dina(n15826), .dinb(n15825), .dout(n15827));
  jand g15754(.dina(n15827), .dinb(n15818), .dout(n15828));
  jxor g15755(.dina(n15828), .dinb(n15816), .dout(n15829));
  jxor g15756(.dina(n15829), .dinb(n15567), .dout(n15830));
  jxor g15757(.dina(n15830), .dinb(n15790), .dout(n15831));
  jand g15758(.dina(n15831), .dinb(n6495), .dout(n15832));
  jand g15759(.dina(n15829), .dinb(n6503), .dout(n15833));
  jand g15760(.dina(n15567), .dinb(n6506), .dout(n15834));
  jand g15761(.dina(n15315), .dinb(n6500), .dout(n15835));
  jor  g15762(.dina(n15835), .dinb(n15834), .dout(n15836));
  jor  g15763(.dina(n15836), .dinb(n15833), .dout(n15837));
  jor  g15764(.dina(n15837), .dinb(n15832), .dout(n15838));
  jxor g15765(.dina(n15838), .dinb(n6219), .dout(n15839));
  jxor g15766(.dina(n15839), .dinb(n15787), .dout(n15840));
  jxor g15767(.dina(n15840), .dinb(n15595), .dout(n15841));
  jxor g15768(.dina(n15841), .dinb(n15579), .dout(n15842));
  jnot g15769(.din(n15327), .dout(n15843));
  jnot g15770(.din(n15579), .dout(n15844));
  jand g15771(.dina(n15844), .dinb(n15022), .dout(n15845));
  jor  g15772(.dina(n15845), .dinb(n15843), .dout(n15846));
  jnot g15773(.din(n15846), .dout(n15847));
  jxor g15774(.dina(n15847), .dinb(n15842), .dout(n15848));
  jand g15775(.dina(n15848), .dinb(n71), .dout(n15849));
  jand g15776(.dina(n15841), .dinb(n796), .dout(n15850));
  jand g15777(.dina(n15327), .dinb(n1806), .dout(n15851));
  jand g15778(.dina(n15579), .dinb(n731), .dout(n15852));
  jor  g15779(.dina(n15852), .dinb(n15851), .dout(n15853));
  jor  g15780(.dina(n15853), .dinb(n15850), .dout(n15854));
  jor  g15781(.dina(n15854), .dinb(n15849), .dout(n15855));
  jxor g15782(.dina(n15855), .dinb(n77), .dout(n15856));
  jxor g15783(.dina(n15856), .dinb(n15591), .dout(n15857));
  jnot g15784(.din(n15857), .dout(n15858));
  jand g15785(.dina(n15785), .dinb(n15777), .dout(n15859));
  jnot g15786(.din(n15859), .dout(n15860));
  jnot g15787(.din(n15501), .dout(n15861));
  jor  g15788(.dina(n15861), .dinb(n15353), .dout(n15862));
  jand g15789(.dina(n15862), .dinb(n15600), .dout(n15863));
  jxor g15790(.dina(n15776), .dinb(n15863), .dout(n15864));
  jxor g15791(.dina(n15785), .dinb(n15864), .dout(n15865));
  jor  g15792(.dina(n15865), .dinb(n15599), .dout(n15866));
  jand g15793(.dina(n15866), .dinb(n15860), .dout(n15867));
  jor  g15794(.dina(n15775), .dinb(n15767), .dout(n15868));
  jnot g15795(.din(n15868), .dout(n15869));
  jand g15796(.dina(n15776), .dinb(n15604), .dout(n15870));
  jor  g15797(.dina(n15870), .dinb(n15869), .dout(n15871));
  jnot g15798(.din(n15756), .dout(n15872));
  jor  g15799(.dina(n15764), .dinb(n15872), .dout(n15873));
  jor  g15800(.dina(n15765), .dinb(n15608), .dout(n15874));
  jand g15801(.dina(n15874), .dinb(n15873), .dout(n15875));
  jnot g15802(.din(n15746), .dout(n15876));
  jor  g15803(.dina(n15754), .dinb(n15876), .dout(n15877));
  jor  g15804(.dina(n15755), .dinb(n15612), .dout(n15878));
  jand g15805(.dina(n15878), .dinb(n15877), .dout(n15879));
  jor  g15806(.dina(n15744), .dinb(n15736), .dout(n15880));
  jnot g15807(.din(n15880), .dout(n15881));
  jand g15808(.dina(n15745), .dinb(n15615), .dout(n15882));
  jor  g15809(.dina(n15882), .dinb(n15881), .dout(n15883));
  jor  g15810(.dina(n15733), .dinb(n15725), .dout(n15884));
  jand g15811(.dina(n15734), .dinb(n15620), .dout(n15885));
  jnot g15812(.din(n15885), .dout(n15886));
  jand g15813(.dina(n15886), .dinb(n15884), .dout(n15887));
  jnot g15814(.din(n15887), .dout(n15888));
  jor  g15815(.dina(n15722), .dinb(n15714), .dout(n15889));
  jand g15816(.dina(n15723), .dinb(n15625), .dout(n15890));
  jnot g15817(.din(n15890), .dout(n15891));
  jand g15818(.dina(n15891), .dinb(n15889), .dout(n15892));
  jnot g15819(.din(n15892), .dout(n15893));
  jor  g15820(.dina(n15711), .dinb(n15703), .dout(n15894));
  jand g15821(.dina(n15712), .dinb(n15630), .dout(n15895));
  jnot g15822(.din(n15895), .dout(n15896));
  jand g15823(.dina(n15896), .dinb(n15894), .dout(n15897));
  jnot g15824(.din(n15897), .dout(n15898));
  jor  g15825(.dina(n15700), .dinb(n15692), .dout(n15899));
  jand g15826(.dina(n15701), .dinb(n15635), .dout(n15900));
  jnot g15827(.din(n15900), .dout(n15901));
  jand g15828(.dina(n15901), .dinb(n15899), .dout(n15902));
  jnot g15829(.din(n15902), .dout(n15903));
  jand g15830(.dina(n15689), .dinb(n15682), .dout(n15904));
  jand g15831(.dina(n15690), .dinb(n15638), .dout(n15905));
  jor  g15832(.dina(n15905), .dinb(n15904), .dout(n15906));
  jand g15833(.dina(n2560), .dinb(n1682), .dout(n15907));
  jand g15834(.dina(n1731), .dinb(n541), .dout(n15908));
  jand g15835(.dina(n15908), .dinb(n1375), .dout(n15909));
  jand g15836(.dina(n15909), .dinb(n934), .dout(n15910));
  jand g15837(.dina(n15910), .dinb(n3110), .dout(n15911));
  jand g15838(.dina(n15911), .dinb(n352), .dout(n15912));
  jand g15839(.dina(n15912), .dinb(n15907), .dout(n15913));
  jand g15840(.dina(n3856), .dinb(n1477), .dout(n15914));
  jand g15841(.dina(n1283), .dinb(n662), .dout(n15915));
  jand g15842(.dina(n15915), .dinb(n3897), .dout(n15916));
  jand g15843(.dina(n15916), .dinb(n14314), .dout(n15917));
  jand g15844(.dina(n15917), .dinb(n2087), .dout(n15918));
  jand g15845(.dina(n1470), .dinb(n1040), .dout(n15919));
  jand g15846(.dina(n15919), .dinb(n3066), .dout(n15920));
  jand g15847(.dina(n15920), .dinb(n14396), .dout(n15921));
  jand g15848(.dina(n5378), .dinb(n554), .dout(n15922));
  jand g15849(.dina(n15922), .dinb(n15921), .dout(n15923));
  jand g15850(.dina(n15923), .dinb(n1306), .dout(n15924));
  jand g15851(.dina(n15924), .dinb(n15918), .dout(n15925));
  jand g15852(.dina(n15925), .dinb(n15914), .dout(n15926));
  jand g15853(.dina(n15926), .dinb(n15913), .dout(n15927));
  jand g15854(.dina(n12334), .dinb(n1686), .dout(n15928));
  jand g15855(.dina(n1373), .dinb(n929), .dout(n15929));
  jand g15856(.dina(n886), .dinb(n470), .dout(n15930));
  jand g15857(.dina(n15930), .dinb(n1288), .dout(n15931));
  jand g15858(.dina(n15931), .dinb(n15929), .dout(n15932));
  jand g15859(.dina(n4541), .dinb(n3345), .dout(n15933));
  jand g15860(.dina(n15933), .dinb(n5984), .dout(n15934));
  jand g15861(.dina(n15934), .dinb(n15932), .dout(n15935));
  jand g15862(.dina(n15935), .dinb(n15928), .dout(n15936));
  jand g15863(.dina(n1847), .dinb(n130), .dout(n15937));
  jand g15864(.dina(n2587), .dinb(n1271), .dout(n15938));
  jand g15865(.dina(n15938), .dinb(n15937), .dout(n15939));
  jand g15866(.dina(n1212), .dinb(n1260), .dout(n15940));
  jand g15867(.dina(n15940), .dinb(n4422), .dout(n15941));
  jand g15868(.dina(n650), .dinb(n547), .dout(n15942));
  jand g15869(.dina(n15942), .dinb(n15941), .dout(n15943));
  jand g15870(.dina(n15943), .dinb(n15939), .dout(n15944));
  jand g15871(.dina(n3041), .dinb(n1716), .dout(n15945));
  jand g15872(.dina(n15945), .dinb(n14301), .dout(n15946));
  jand g15873(.dina(n15946), .dinb(n15944), .dout(n15947));
  jand g15874(.dina(n15947), .dinb(n15936), .dout(n15948));
  jand g15875(.dina(n15948), .dinb(n15927), .dout(n15949));
  jnot g15876(.din(n15949), .dout(n15950));
  jand g15877(.dina(n8962), .dinb(n5076), .dout(n15951));
  jand g15878(.dina(n8740), .dinb(n5084), .dout(n15952));
  jand g15879(.dina(n8022), .dinb(n6050), .dout(n15953));
  jand g15880(.dina(n8268), .dinb(n5082), .dout(n15954));
  jor  g15881(.dina(n15954), .dinb(n15953), .dout(n15955));
  jor  g15882(.dina(n15955), .dinb(n15952), .dout(n15956));
  jor  g15883(.dina(n15956), .dinb(n15951), .dout(n15957));
  jxor g15884(.dina(n15957), .dinb(n15950), .dout(n15958));
  jxor g15885(.dina(n15958), .dinb(n15906), .dout(n15959));
  jand g15886(.dina(n9252), .dinb(n2936), .dout(n15960));
  jand g15887(.dina(n9250), .dinb(n2943), .dout(n15961));
  jand g15888(.dina(n8936), .dinb(n2940), .dout(n15962));
  jand g15889(.dina(n8723), .dinb(n3684), .dout(n15963));
  jor  g15890(.dina(n15963), .dinb(n15962), .dout(n15964));
  jor  g15891(.dina(n15964), .dinb(n15961), .dout(n15965));
  jor  g15892(.dina(n15965), .dinb(n15960), .dout(n15966));
  jxor g15893(.dina(n15966), .dinb(\a[29] ), .dout(n15967));
  jxor g15894(.dina(n15967), .dinb(n15959), .dout(n15968));
  jxor g15895(.dina(n15968), .dinb(n15903), .dout(n15969));
  jnot g15896(.din(n15969), .dout(n15970));
  jand g15897(.dina(n9874), .dinb(n71), .dout(n15971));
  jand g15898(.dina(n9872), .dinb(n796), .dout(n15972));
  jand g15899(.dina(n9655), .dinb(n731), .dout(n15973));
  jand g15900(.dina(n9656), .dinb(n1806), .dout(n15974));
  jor  g15901(.dina(n15974), .dinb(n15973), .dout(n15975));
  jor  g15902(.dina(n15975), .dinb(n15972), .dout(n15976));
  jor  g15903(.dina(n15976), .dinb(n15971), .dout(n15977));
  jxor g15904(.dina(n15977), .dinb(n77), .dout(n15978));
  jxor g15905(.dina(n15978), .dinb(n15970), .dout(n15979));
  jxor g15906(.dina(n15979), .dinb(n15898), .dout(n15980));
  jnot g15907(.din(n15980), .dout(n15981));
  jand g15908(.dina(n10850), .dinb(n806), .dout(n15982));
  jand g15909(.dina(n10647), .dinb(n1612), .dout(n15983));
  jand g15910(.dina(n10640), .dinb(n1620), .dout(n15984));
  jor  g15911(.dina(n15984), .dinb(n15983), .dout(n15985));
  jand g15912(.dina(n10305), .dinb(n1644), .dout(n15986));
  jor  g15913(.dina(n15986), .dinb(n15985), .dout(n15987));
  jor  g15914(.dina(n15987), .dinb(n15982), .dout(n15988));
  jxor g15915(.dina(n15988), .dinb(n65), .dout(n15989));
  jxor g15916(.dina(n15989), .dinb(n15981), .dout(n15990));
  jxor g15917(.dina(n15990), .dinb(n15893), .dout(n15991));
  jnot g15918(.din(n15991), .dout(n15992));
  jand g15919(.dina(n11824), .dinb(n1819), .dout(n15993));
  jand g15920(.dina(n11647), .dinb(n2243), .dout(n15994));
  jand g15921(.dina(n11306), .dinb(n2180), .dout(n15995));
  jand g15922(.dina(n10836), .dinb(n2185), .dout(n15996));
  jor  g15923(.dina(n15996), .dinb(n15995), .dout(n15997));
  jor  g15924(.dina(n15997), .dinb(n15994), .dout(n15998));
  jor  g15925(.dina(n15998), .dinb(n15993), .dout(n15999));
  jxor g15926(.dina(n15999), .dinb(n2196), .dout(n16000));
  jxor g15927(.dina(n16000), .dinb(n15992), .dout(n16001));
  jxor g15928(.dina(n16001), .dinb(n15888), .dout(n16002));
  jnot g15929(.din(n16002), .dout(n16003));
  jand g15930(.dina(n12284), .dinb(n2743), .dout(n16004));
  jand g15931(.dina(n12282), .dinb(n2752), .dout(n16005));
  jand g15932(.dina(n11798), .dinb(n2748), .dout(n16006));
  jand g15933(.dina(n11646), .dinb(n2757), .dout(n16007));
  jor  g15934(.dina(n16007), .dinb(n16006), .dout(n16008));
  jor  g15935(.dina(n16008), .dinb(n16005), .dout(n16009));
  jor  g15936(.dina(n16009), .dinb(n16004), .dout(n16010));
  jxor g15937(.dina(n16010), .dinb(n2441), .dout(n16011));
  jxor g15938(.dina(n16011), .dinb(n16003), .dout(n16012));
  jxor g15939(.dina(n16012), .dinb(n15883), .dout(n16013));
  jand g15940(.dina(n12671), .dinb(n3423), .dout(n16014));
  jand g15941(.dina(n12536), .dinb(n3428), .dout(n16015));
  jand g15942(.dina(n12669), .dinb(n3569), .dout(n16016));
  jor  g15943(.dina(n16016), .dinb(n16015), .dout(n16017));
  jand g15944(.dina(n12547), .dinb(n3210), .dout(n16018));
  jor  g15945(.dina(n16018), .dinb(n16017), .dout(n16019));
  jor  g15946(.dina(n16019), .dinb(n16014), .dout(n16020));
  jxor g15947(.dina(n16020), .dinb(n3473), .dout(n16021));
  jxor g15948(.dina(n16021), .dinb(n16013), .dout(n16022));
  jxor g15949(.dina(n16022), .dinb(n15879), .dout(n16023));
  jand g15950(.dina(n13627), .dinb(n4022), .dout(n16024));
  jand g15951(.dina(n13478), .dinb(n4027), .dout(n16025));
  jand g15952(.dina(n13469), .dinb(n4220), .dout(n16026));
  jor  g15953(.dina(n16026), .dinb(n16025), .dout(n16027));
  jand g15954(.dina(n13248), .dinb(n3870), .dout(n16028));
  jor  g15955(.dina(n16028), .dinb(n16027), .dout(n16029));
  jor  g15956(.dina(n16029), .dinb(n16024), .dout(n16030));
  jxor g15957(.dina(n16030), .dinb(n4050), .dout(n16031));
  jxor g15958(.dina(n16031), .dinb(n16023), .dout(n16032));
  jnot g15959(.din(n16032), .dout(n16033));
  jxor g15960(.dina(n16033), .dinb(n15875), .dout(n16034));
  jand g15961(.dina(n14579), .dinb(n4691), .dout(n16035));
  jand g15962(.dina(n14448), .dinb(n4941), .dout(n16036));
  jand g15963(.dina(n14249), .dinb(n4696), .dout(n16037));
  jand g15964(.dina(n13614), .dinb(n4701), .dout(n16038));
  jor  g15965(.dina(n16038), .dinb(n16037), .dout(n16039));
  jor  g15966(.dina(n16039), .dinb(n16036), .dout(n16040));
  jor  g15967(.dina(n16040), .dinb(n16035), .dout(n16041));
  jxor g15968(.dina(n16041), .dinb(n4713), .dout(n16042));
  jxor g15969(.dina(n16042), .dinb(n16034), .dout(n16043));
  jxor g15970(.dina(n16043), .dinb(n15871), .dout(n16044));
  jand g15971(.dina(n15317), .dinb(n5280), .dout(n16045));
  jand g15972(.dina(n15315), .dinb(n5814), .dout(n16046));
  jand g15973(.dina(n14549), .dinb(n5531), .dout(n16047));
  jand g15974(.dina(n14447), .dinb(n5536), .dout(n16048));
  jor  g15975(.dina(n16048), .dinb(n16047), .dout(n16049));
  jor  g15976(.dina(n16049), .dinb(n16046), .dout(n16050));
  jor  g15977(.dina(n16050), .dinb(n16045), .dout(n16051));
  jxor g15978(.dina(n16051), .dinb(\a[5] ), .dout(n16052));
  jxor g15979(.dina(n16052), .dinb(n16044), .dout(n16053));
  jxor g15980(.dina(n16053), .dinb(n15867), .dout(n16054));
  jand g15981(.dina(n15829), .dinb(n15567), .dout(n16055));
  jand g15982(.dina(n15830), .dinb(n15790), .dout(n16056));
  jor  g15983(.dina(n16056), .dinb(n16055), .dout(n16057));
  jnot g15984(.din(n15558), .dout(n16058));
  jand g15985(.dina(n15811), .dinb(n16058), .dout(n16059));
  jand g15986(.dina(n15813), .dinb(n15800), .dout(n16060));
  jor  g15987(.dina(n16060), .dinb(n16059), .dout(n16061));
  jand g15988(.dina(n6473), .dinb(n456), .dout(n16062));
  jand g15989(.dina(n7987), .dinb(n583), .dout(n16063));
  jand g15990(.dina(n16063), .dinb(n15544), .dout(n16064));
  jand g15991(.dina(n16064), .dinb(n16062), .dout(n16065));
  jand g15992(.dina(n1765), .dinb(n1735), .dout(n16066));
  jand g15993(.dina(n16066), .dinb(n2023), .dout(n16067));
  jand g15994(.dina(n16067), .dinb(n16065), .dout(n16068));
  jand g15995(.dina(n16068), .dinb(n7647), .dout(n16069));
  jnot g15996(.din(n16069), .dout(n16070));
  jxor g15997(.dina(n16070), .dinb(n15811), .dout(n16071));
  jxor g15998(.dina(n16071), .dinb(n16061), .dout(n16076));
  jnot g15999(.din(n16076), .dout(n16077));
  jand g16000(.dina(n15814), .dinb(n15793), .dout(n16078));
  jnot g16001(.din(n16078), .dout(n16079));
  jor  g16002(.dina(n15828), .dinb(n15816), .dout(n16080));
  jand g16003(.dina(n16080), .dinb(n16079), .dout(n16081));
  jxor g16004(.dina(n16081), .dinb(n16077), .dout(n16082));
  jxor g16005(.dina(n16082), .dinb(n15829), .dout(n16083));
  jxor g16006(.dina(n16083), .dinb(n16057), .dout(n16084));
  jand g16007(.dina(n16084), .dinb(n6495), .dout(n16085));
  jand g16008(.dina(n16082), .dinb(n6503), .dout(n16086));
  jand g16009(.dina(n15829), .dinb(n6506), .dout(n16087));
  jand g16010(.dina(n15567), .dinb(n6500), .dout(n16088));
  jor  g16011(.dina(n16088), .dinb(n16087), .dout(n16089));
  jor  g16012(.dina(n16089), .dinb(n16086), .dout(n16090));
  jor  g16013(.dina(n16090), .dinb(n16085), .dout(n16091));
  jxor g16014(.dina(n16091), .dinb(n6219), .dout(n16092));
  jor  g16015(.dina(n16092), .dinb(n16054), .dout(n16093));
  jor  g16016(.dina(n15839), .dinb(n15787), .dout(n16094));
  jnot g16017(.din(n15595), .dout(n16095));
  jnot g16018(.din(n15596), .dout(n16096));
  jnot g16019(.din(n15348), .dout(n16097));
  jand g16020(.dina(n15511), .dinb(n16097), .dout(n16098));
  jor  g16021(.dina(n16098), .dinb(n16096), .dout(n16099));
  jxor g16022(.dina(n15786), .dinb(n16099), .dout(n16100));
  jxor g16023(.dina(n15839), .dinb(n16100), .dout(n16101));
  jor  g16024(.dina(n16101), .dinb(n16095), .dout(n16102));
  jand g16025(.dina(n16102), .dinb(n16094), .dout(n16103));
  jand g16026(.dina(n15786), .dinb(n16099), .dout(n16104));
  jor  g16027(.dina(n16104), .dinb(n15859), .dout(n16105));
  jxor g16028(.dina(n16053), .dinb(n16105), .dout(n16106));
  jxor g16029(.dina(n16092), .dinb(n16106), .dout(n16107));
  jor  g16030(.dina(n16107), .dinb(n16103), .dout(n16108));
  jand g16031(.dina(n16108), .dinb(n16093), .dout(n16109));
  jand g16032(.dina(n16052), .dinb(n16044), .dout(n16110));
  jand g16033(.dina(n16053), .dinb(n16105), .dout(n16111));
  jor  g16034(.dina(n16111), .dinb(n16110), .dout(n16112));
  jor  g16035(.dina(n16042), .dinb(n16034), .dout(n16113));
  jnot g16036(.din(n15605), .dout(n16114));
  jnot g16037(.din(n15357), .dout(n16115));
  jand g16038(.dina(n15491), .dinb(n16115), .dout(n16116));
  jor  g16039(.dina(n16116), .dinb(n16114), .dout(n16117));
  jxor g16040(.dina(n15766), .dinb(n16117), .dout(n16118));
  jxor g16041(.dina(n15775), .dinb(n16118), .dout(n16119));
  jor  g16042(.dina(n16119), .dinb(n15863), .dout(n16120));
  jand g16043(.dina(n16120), .dinb(n15868), .dout(n16121));
  jnot g16044(.din(n15873), .dout(n16122));
  jand g16045(.dina(n15766), .dinb(n16117), .dout(n16123));
  jor  g16046(.dina(n16123), .dinb(n16122), .dout(n16124));
  jxor g16047(.dina(n16033), .dinb(n16124), .dout(n16125));
  jxor g16048(.dina(n16042), .dinb(n16125), .dout(n16126));
  jor  g16049(.dina(n16126), .dinb(n16121), .dout(n16127));
  jand g16050(.dina(n16127), .dinb(n16113), .dout(n16128));
  jnot g16051(.din(n16023), .dout(n16129));
  jor  g16052(.dina(n16031), .dinb(n16129), .dout(n16130));
  jor  g16053(.dina(n16032), .dinb(n15875), .dout(n16131));
  jand g16054(.dina(n16131), .dinb(n16130), .dout(n16132));
  jnot g16055(.din(n16013), .dout(n16133));
  jor  g16056(.dina(n16021), .dinb(n16133), .dout(n16134));
  jor  g16057(.dina(n16022), .dinb(n15879), .dout(n16135));
  jand g16058(.dina(n16135), .dinb(n16134), .dout(n16136));
  jor  g16059(.dina(n16011), .dinb(n16003), .dout(n16137));
  jnot g16060(.din(n16137), .dout(n16138));
  jand g16061(.dina(n16012), .dinb(n15883), .dout(n16139));
  jor  g16062(.dina(n16139), .dinb(n16138), .dout(n16140));
  jor  g16063(.dina(n16000), .dinb(n15992), .dout(n16141));
  jand g16064(.dina(n16001), .dinb(n15888), .dout(n16142));
  jnot g16065(.din(n16142), .dout(n16143));
  jand g16066(.dina(n16143), .dinb(n16141), .dout(n16144));
  jnot g16067(.din(n16144), .dout(n16145));
  jor  g16068(.dina(n15989), .dinb(n15981), .dout(n16146));
  jand g16069(.dina(n15990), .dinb(n15893), .dout(n16147));
  jnot g16070(.din(n16147), .dout(n16148));
  jand g16071(.dina(n16148), .dinb(n16146), .dout(n16149));
  jnot g16072(.din(n16149), .dout(n16150));
  jor  g16073(.dina(n15978), .dinb(n15970), .dout(n16151));
  jand g16074(.dina(n15979), .dinb(n15898), .dout(n16152));
  jnot g16075(.din(n16152), .dout(n16153));
  jand g16076(.dina(n16153), .dinb(n16151), .dout(n16154));
  jnot g16077(.din(n16154), .dout(n16155));
  jand g16078(.dina(n15967), .dinb(n15959), .dout(n16156));
  jand g16079(.dina(n15968), .dinb(n15903), .dout(n16157));
  jor  g16080(.dina(n16157), .dinb(n16156), .dout(n16158));
  jand g16081(.dina(n15957), .dinb(n15950), .dout(n16159));
  jand g16082(.dina(n15958), .dinb(n15906), .dout(n16160));
  jor  g16083(.dina(n16160), .dinb(n16159), .dout(n16161));
  jand g16084(.dina(n7259), .dinb(n1465), .dout(n16162));
  jand g16085(.dina(n1579), .dinb(n685), .dout(n16163));
  jand g16086(.dina(n16163), .dinb(n16162), .dout(n16164));
  jand g16087(.dina(n3834), .dinb(n2605), .dout(n16165));
  jand g16088(.dina(n16165), .dinb(n16164), .dout(n16166));
  jand g16089(.dina(n1227), .dinb(n541), .dout(n16167));
  jand g16090(.dina(n16167), .dinb(n1971), .dout(n16168));
  jand g16091(.dina(n16168), .dinb(n7496), .dout(n16169));
  jand g16092(.dina(n16169), .dinb(n8402), .dout(n16170));
  jand g16093(.dina(n16170), .dinb(n326), .dout(n16171));
  jand g16094(.dina(n16171), .dinb(n16166), .dout(n16172));
  jand g16095(.dina(n1017), .dinb(n701), .dout(n16173));
  jand g16096(.dina(n16173), .dinb(n622), .dout(n16174));
  jand g16097(.dina(n1589), .dinb(n1366), .dout(n16175));
  jand g16098(.dina(n1713), .dinb(n428), .dout(n16176));
  jand g16099(.dina(n16176), .dinb(n1317), .dout(n16177));
  jand g16100(.dina(n16177), .dinb(n16175), .dout(n16178));
  jand g16101(.dina(n16178), .dinb(n13177), .dout(n16179));
  jand g16102(.dina(n16179), .dinb(n16174), .dout(n16180));
  jand g16103(.dina(n16180), .dinb(n1286), .dout(n16181));
  jand g16104(.dina(n14219), .dinb(n8134), .dout(n16182));
  jand g16105(.dina(n16182), .dinb(n16181), .dout(n16183));
  jand g16106(.dina(n16183), .dinb(n16172), .dout(n16184));
  jand g16107(.dina(n7254), .dinb(n714), .dout(n16185));
  jand g16108(.dina(n8602), .dinb(n7105), .dout(n16186));
  jand g16109(.dina(n16186), .dinb(n1473), .dout(n16187));
  jand g16110(.dina(n16187), .dinb(n16185), .dout(n16188));
  jand g16111(.dina(n3978), .dinb(n563), .dout(n16189));
  jand g16112(.dina(n7499), .dinb(n1169), .dout(n16190));
  jand g16113(.dina(n16190), .dinb(n2023), .dout(n16191));
  jand g16114(.dina(n16191), .dinb(n16189), .dout(n16192));
  jand g16115(.dina(n16192), .dinb(n16188), .dout(n16193));
  jand g16116(.dina(n886), .dinb(n1903), .dout(n16194));
  jand g16117(.dina(n16194), .dinb(n13420), .dout(n16195));
  jand g16118(.dina(n16195), .dinb(n1824), .dout(n16196));
  jand g16119(.dina(n16196), .dinb(n7247), .dout(n16197));
  jand g16120(.dina(n16197), .dinb(n16193), .dout(n16198));
  jand g16121(.dina(n1228), .dinb(n1432), .dout(n16199));
  jand g16122(.dina(n16199), .dinb(n716), .dout(n16200));
  jand g16123(.dina(n16200), .dinb(n908), .dout(n16201));
  jand g16124(.dina(n16201), .dinb(n4675), .dout(n16202));
  jand g16125(.dina(n16202), .dinb(n463), .dout(n16203));
  jand g16126(.dina(n16203), .dinb(n7831), .dout(n16204));
  jand g16127(.dina(n11394), .dinb(n3329), .dout(n16205));
  jand g16128(.dina(n16205), .dinb(n13157), .dout(n16206));
  jand g16129(.dina(n3396), .dinb(n586), .dout(n16207));
  jand g16130(.dina(n16207), .dinb(n16206), .dout(n16208));
  jand g16131(.dina(n16208), .dinb(n3737), .dout(n16209));
  jand g16132(.dina(n16209), .dinb(n13186), .dout(n16210));
  jand g16133(.dina(n16210), .dinb(n16204), .dout(n16211));
  jand g16134(.dina(n16211), .dinb(n16198), .dout(n16212));
  jand g16135(.dina(n16212), .dinb(n16184), .dout(n16213));
  jnot g16136(.din(n16213), .dout(n16214));
  jand g16137(.dina(n8950), .dinb(n5076), .dout(n16215));
  jand g16138(.dina(n8723), .dinb(n5084), .dout(n16216));
  jand g16139(.dina(n8268), .dinb(n6050), .dout(n16217));
  jand g16140(.dina(n8740), .dinb(n5082), .dout(n16218));
  jor  g16141(.dina(n16218), .dinb(n16217), .dout(n16219));
  jor  g16142(.dina(n16219), .dinb(n16216), .dout(n16220));
  jor  g16143(.dina(n16220), .dinb(n16215), .dout(n16221));
  jxor g16144(.dina(n16221), .dinb(n16214), .dout(n16222));
  jxor g16145(.dina(n16222), .dinb(n16161), .dout(n16223));
  jnot g16146(.din(n16223), .dout(n16224));
  jand g16147(.dina(n9898), .dinb(n2936), .dout(n16225));
  jand g16148(.dina(n9250), .dinb(n2940), .dout(n16226));
  jand g16149(.dina(n9656), .dinb(n2943), .dout(n16227));
  jor  g16150(.dina(n16227), .dinb(n16226), .dout(n16228));
  jand g16151(.dina(n8936), .dinb(n3684), .dout(n16229));
  jor  g16152(.dina(n16229), .dinb(n16228), .dout(n16230));
  jor  g16153(.dina(n16230), .dinb(n16225), .dout(n16231));
  jxor g16154(.dina(n16231), .dinb(n93), .dout(n16232));
  jxor g16155(.dina(n16232), .dinb(n16224), .dout(n16233));
  jxor g16156(.dina(n16233), .dinb(n16158), .dout(n16234));
  jnot g16157(.din(n16234), .dout(n16235));
  jand g16158(.dina(n10307), .dinb(n71), .dout(n16236));
  jand g16159(.dina(n10305), .dinb(n796), .dout(n16237));
  jand g16160(.dina(n9872), .dinb(n731), .dout(n16238));
  jand g16161(.dina(n9655), .dinb(n1806), .dout(n16239));
  jor  g16162(.dina(n16239), .dinb(n16238), .dout(n16240));
  jor  g16163(.dina(n16240), .dinb(n16237), .dout(n16241));
  jor  g16164(.dina(n16241), .dinb(n16236), .dout(n16242));
  jxor g16165(.dina(n16242), .dinb(n77), .dout(n16243));
  jxor g16166(.dina(n16243), .dinb(n16235), .dout(n16244));
  jxor g16167(.dina(n16244), .dinb(n16155), .dout(n16245));
  jnot g16168(.din(n16245), .dout(n16246));
  jand g16169(.dina(n10838), .dinb(n806), .dout(n16247));
  jand g16170(.dina(n10836), .dinb(n1620), .dout(n16248));
  jand g16171(.dina(n10640), .dinb(n1612), .dout(n16249));
  jand g16172(.dina(n10647), .dinb(n1644), .dout(n16250));
  jor  g16173(.dina(n16250), .dinb(n16249), .dout(n16251));
  jor  g16174(.dina(n16251), .dinb(n16248), .dout(n16252));
  jor  g16175(.dina(n16252), .dinb(n16247), .dout(n16253));
  jxor g16176(.dina(n16253), .dinb(n65), .dout(n16254));
  jxor g16177(.dina(n16254), .dinb(n16246), .dout(n16255));
  jxor g16178(.dina(n16255), .dinb(n16150), .dout(n16256));
  jnot g16179(.din(n16256), .dout(n16257));
  jand g16180(.dina(n11812), .dinb(n1819), .dout(n16258));
  jand g16181(.dina(n11647), .dinb(n2180), .dout(n16259));
  jand g16182(.dina(n11646), .dinb(n2243), .dout(n16260));
  jor  g16183(.dina(n16260), .dinb(n16259), .dout(n16261));
  jand g16184(.dina(n11306), .dinb(n2185), .dout(n16262));
  jor  g16185(.dina(n16262), .dinb(n16261), .dout(n16263));
  jor  g16186(.dina(n16263), .dinb(n16258), .dout(n16264));
  jxor g16187(.dina(n16264), .dinb(n2196), .dout(n16265));
  jxor g16188(.dina(n16265), .dinb(n16257), .dout(n16266));
  jxor g16189(.dina(n16266), .dinb(n16145), .dout(n16267));
  jand g16190(.dina(n12696), .dinb(n2743), .dout(n16268));
  jand g16191(.dina(n12547), .dinb(n2752), .dout(n16269));
  jand g16192(.dina(n12282), .dinb(n2748), .dout(n16270));
  jand g16193(.dina(n11798), .dinb(n2757), .dout(n16271));
  jor  g16194(.dina(n16271), .dinb(n16270), .dout(n16272));
  jor  g16195(.dina(n16272), .dinb(n16269), .dout(n16273));
  jor  g16196(.dina(n16273), .dinb(n16268), .dout(n16274));
  jxor g16197(.dina(n16274), .dinb(\a[17] ), .dout(n16275));
  jxor g16198(.dina(n16275), .dinb(n16267), .dout(n16276));
  jxor g16199(.dina(n16276), .dinb(n16140), .dout(n16277));
  jand g16200(.dina(n13250), .dinb(n3423), .dout(n16278));
  jand g16201(.dina(n12669), .dinb(n3428), .dout(n16279));
  jand g16202(.dina(n13248), .dinb(n3569), .dout(n16280));
  jor  g16203(.dina(n16280), .dinb(n16279), .dout(n16281));
  jand g16204(.dina(n12536), .dinb(n3210), .dout(n16282));
  jor  g16205(.dina(n16282), .dinb(n16281), .dout(n16283));
  jor  g16206(.dina(n16283), .dinb(n16278), .dout(n16284));
  jxor g16207(.dina(n16284), .dinb(n3473), .dout(n16285));
  jxor g16208(.dina(n16285), .dinb(n16277), .dout(n16286));
  jxor g16209(.dina(n16286), .dinb(n16136), .dout(n16287));
  jand g16210(.dina(n13616), .dinb(n4022), .dout(n16288));
  jand g16211(.dina(n13469), .dinb(n4027), .dout(n16289));
  jand g16212(.dina(n13614), .dinb(n4220), .dout(n16290));
  jor  g16213(.dina(n16290), .dinb(n16289), .dout(n16291));
  jand g16214(.dina(n13478), .dinb(n3870), .dout(n16292));
  jor  g16215(.dina(n16292), .dinb(n16291), .dout(n16293));
  jor  g16216(.dina(n16293), .dinb(n16288), .dout(n16294));
  jxor g16217(.dina(n16294), .dinb(n4050), .dout(n16295));
  jxor g16218(.dina(n16295), .dinb(n16287), .dout(n16296));
  jnot g16219(.din(n16296), .dout(n16297));
  jxor g16220(.dina(n16297), .dinb(n16132), .dout(n16298));
  jand g16221(.dina(n14562), .dinb(n4691), .dout(n16299));
  jand g16222(.dina(n14448), .dinb(n4696), .dout(n16300));
  jand g16223(.dina(n14447), .dinb(n4941), .dout(n16301));
  jor  g16224(.dina(n16301), .dinb(n16300), .dout(n16302));
  jand g16225(.dina(n14249), .dinb(n4701), .dout(n16303));
  jor  g16226(.dina(n16303), .dinb(n16302), .dout(n16304));
  jor  g16227(.dina(n16304), .dinb(n16299), .dout(n16305));
  jxor g16228(.dina(n16305), .dinb(n4713), .dout(n16306));
  jxor g16229(.dina(n16306), .dinb(n16298), .dout(n16307));
  jxor g16230(.dina(n16307), .dinb(n16128), .dout(n16308));
  jand g16231(.dina(n15569), .dinb(n5280), .dout(n16309));
  jand g16232(.dina(n15315), .dinb(n5531), .dout(n16310));
  jand g16233(.dina(n15567), .dinb(n5814), .dout(n16311));
  jor  g16234(.dina(n16311), .dinb(n16310), .dout(n16312));
  jand g16235(.dina(n14549), .dinb(n5536), .dout(n16313));
  jor  g16236(.dina(n16313), .dinb(n16312), .dout(n16314));
  jor  g16237(.dina(n16314), .dinb(n16309), .dout(n16315));
  jxor g16238(.dina(n16315), .dinb(n5277), .dout(n16316));
  jxor g16239(.dina(n16316), .dinb(n16308), .dout(n16317));
  jxor g16240(.dina(n16317), .dinb(n16112), .dout(n16318));
  jand g16241(.dina(n16082), .dinb(n15829), .dout(n16319));
  jand g16242(.dina(n16083), .dinb(n16057), .dout(n16320));
  jor  g16243(.dina(n16320), .dinb(n16319), .dout(n16321));
  jand g16244(.dina(n16071), .dinb(n16061), .dout(n16322));
  jand g16245(.dina(n15566), .dinb(n15518), .dout(n16323));
  jor  g16246(.dina(n16323), .dinb(n15817), .dout(n16324));
  jand g16247(.dina(n16324), .dinb(n15815), .dout(n16325));
  jor  g16248(.dina(n16325), .dinb(n16078), .dout(n16326));
  jand g16249(.dina(n16326), .dinb(n16076), .dout(n16327));
  jor  g16250(.dina(n16327), .dinb(n16322), .dout(n16328));
  jand g16251(.dina(n6449), .dinb(n6175), .dout(n16329));
  jand g16252(.dina(n1036), .dinb(n843), .dout(n16330));
  jand g16253(.dina(n16330), .dinb(n7671), .dout(n16331));
  jand g16254(.dina(n16331), .dinb(n7661), .dout(n16332));
  jand g16255(.dina(n16332), .dinb(n16329), .dout(n16333));
  jand g16256(.dina(n16333), .dinb(n7275), .dout(n16334));
  jxor g16257(.dina(n16334), .dinb(n15811), .dout(n16335));
  jnot g16258(.din(n16335), .dout(n16336));
  jand g16259(.dina(n16070), .dinb(n15811), .dout(n16339));
  jxor g16260(.dina(n16339), .dinb(n16336), .dout(n16342));
  jxor g16261(.dina(n16342), .dinb(n16328), .dout(n16343));
  jxor g16262(.dina(n16343), .dinb(n16082), .dout(n16344));
  jxor g16263(.dina(n16344), .dinb(n16321), .dout(n16345));
  jand g16264(.dina(n16345), .dinb(n6495), .dout(n16346));
  jand g16265(.dina(n16343), .dinb(n6503), .dout(n16347));
  jand g16266(.dina(n16082), .dinb(n6506), .dout(n16348));
  jand g16267(.dina(n15829), .dinb(n6500), .dout(n16349));
  jor  g16268(.dina(n16349), .dinb(n16348), .dout(n16350));
  jor  g16269(.dina(n16350), .dinb(n16347), .dout(n16351));
  jor  g16270(.dina(n16351), .dinb(n16346), .dout(n16352));
  jxor g16271(.dina(n16352), .dinb(n6219), .dout(n16353));
  jxor g16272(.dina(n16353), .dinb(n16318), .dout(n16354));
  jxor g16273(.dina(n16354), .dinb(n16109), .dout(n16355));
  jnot g16274(.din(n16094), .dout(n16356));
  jand g16275(.dina(n15840), .dinb(n15595), .dout(n16357));
  jor  g16276(.dina(n16357), .dinb(n16356), .dout(n16358));
  jxor g16277(.dina(n16092), .dinb(n16054), .dout(n16359));
  jxor g16278(.dina(n16359), .dinb(n16358), .dout(n16360));
  jand g16279(.dina(n16360), .dinb(n16355), .dout(n16361));
  jand g16280(.dina(n16360), .dinb(n15841), .dout(n16362));
  jand g16281(.dina(n15841), .dinb(n15579), .dout(n16363));
  jand g16282(.dina(n15847), .dinb(n15842), .dout(n16364));
  jor  g16283(.dina(n16364), .dinb(n16363), .dout(n16365));
  jxor g16284(.dina(n16360), .dinb(n15841), .dout(n16366));
  jand g16285(.dina(n16366), .dinb(n16365), .dout(n16367));
  jor  g16286(.dina(n16367), .dinb(n16362), .dout(n16368));
  jxor g16287(.dina(n16360), .dinb(n16355), .dout(n16369));
  jand g16288(.dina(n16369), .dinb(n16368), .dout(n16370));
  jor  g16289(.dina(n16370), .dinb(n16361), .dout(n16371));
  jnot g16290(.din(n16318), .dout(n16372));
  jor  g16291(.dina(n16353), .dinb(n16372), .dout(n16373));
  jor  g16292(.dina(n16354), .dinb(n16109), .dout(n16374));
  jand g16293(.dina(n16374), .dinb(n16373), .dout(n16375));
  jor  g16294(.dina(n16316), .dinb(n16308), .dout(n16376));
  jnot g16295(.din(n16376), .dout(n16377));
  jand g16296(.dina(n16317), .dinb(n16112), .dout(n16378));
  jor  g16297(.dina(n16378), .dinb(n16377), .dout(n16379));
  jor  g16298(.dina(n16306), .dinb(n16298), .dout(n16380));
  jnot g16299(.din(n16130), .dout(n16381));
  jand g16300(.dina(n16033), .dinb(n16124), .dout(n16382));
  jor  g16301(.dina(n16382), .dinb(n16381), .dout(n16383));
  jxor g16302(.dina(n16297), .dinb(n16383), .dout(n16384));
  jxor g16303(.dina(n16306), .dinb(n16384), .dout(n16385));
  jor  g16304(.dina(n16385), .dinb(n16128), .dout(n16386));
  jand g16305(.dina(n16386), .dinb(n16380), .dout(n16387));
  jnot g16306(.din(n16287), .dout(n16388));
  jor  g16307(.dina(n16295), .dinb(n16388), .dout(n16389));
  jor  g16308(.dina(n16296), .dinb(n16132), .dout(n16390));
  jand g16309(.dina(n16390), .dinb(n16389), .dout(n16391));
  jnot g16310(.din(n16277), .dout(n16392));
  jor  g16311(.dina(n16285), .dinb(n16392), .dout(n16393));
  jor  g16312(.dina(n16286), .dinb(n16136), .dout(n16394));
  jand g16313(.dina(n16394), .dinb(n16393), .dout(n16395));
  jand g16314(.dina(n16275), .dinb(n16267), .dout(n16396));
  jand g16315(.dina(n16276), .dinb(n16140), .dout(n16397));
  jor  g16316(.dina(n16397), .dinb(n16396), .dout(n16398));
  jor  g16317(.dina(n16265), .dinb(n16257), .dout(n16399));
  jand g16318(.dina(n16266), .dinb(n16145), .dout(n16400));
  jnot g16319(.din(n16400), .dout(n16401));
  jand g16320(.dina(n16401), .dinb(n16399), .dout(n16402));
  jnot g16321(.din(n16402), .dout(n16403));
  jor  g16322(.dina(n16254), .dinb(n16246), .dout(n16404));
  jand g16323(.dina(n16255), .dinb(n16150), .dout(n16405));
  jnot g16324(.din(n16405), .dout(n16406));
  jand g16325(.dina(n16406), .dinb(n16404), .dout(n16407));
  jnot g16326(.din(n16407), .dout(n16408));
  jor  g16327(.dina(n16243), .dinb(n16235), .dout(n16409));
  jand g16328(.dina(n16244), .dinb(n16155), .dout(n16410));
  jnot g16329(.din(n16410), .dout(n16411));
  jand g16330(.dina(n16411), .dinb(n16409), .dout(n16412));
  jnot g16331(.din(n16412), .dout(n16413));
  jor  g16332(.dina(n16232), .dinb(n16224), .dout(n16414));
  jand g16333(.dina(n16233), .dinb(n16158), .dout(n16415));
  jnot g16334(.din(n16415), .dout(n16416));
  jand g16335(.dina(n16416), .dinb(n16414), .dout(n16417));
  jnot g16336(.din(n16417), .dout(n16418));
  jand g16337(.dina(n16221), .dinb(n16214), .dout(n16419));
  jand g16338(.dina(n16222), .dinb(n16161), .dout(n16420));
  jor  g16339(.dina(n16420), .dinb(n16419), .dout(n16421));
  jand g16340(.dina(n2530), .dinb(n916), .dout(n16422));
  jand g16341(.dina(n16422), .dinb(n3829), .dout(n16423));
  jand g16342(.dina(n16423), .dinb(n14049), .dout(n16424));
  jand g16343(.dina(n7105), .dinb(n1090), .dout(n16425));
  jand g16344(.dina(n16425), .dinb(n981), .dout(n16426));
  jand g16345(.dina(n16426), .dinb(n456), .dout(n16427));
  jand g16346(.dina(n16427), .dinb(n16424), .dout(n16428));
  jand g16347(.dina(n2588), .dinb(n82), .dout(n16429));
  jand g16348(.dina(n1470), .dinb(n695), .dout(n16430));
  jand g16349(.dina(n16430), .dinb(n3092), .dout(n16431));
  jand g16350(.dina(n16431), .dinb(n16429), .dout(n16432));
  jand g16351(.dina(n16432), .dinb(n6349), .dout(n16433));
  jand g16352(.dina(n16433), .dinb(n16428), .dout(n16434));
  jand g16353(.dina(n16434), .dinb(n13164), .dout(n16435));
  jand g16354(.dina(n16435), .dinb(n13529), .dout(n16436));
  jnot g16355(.din(n16436), .dout(n16437));
  jand g16356(.dina(n8938), .dinb(n5076), .dout(n16438));
  jand g16357(.dina(n8936), .dinb(n5084), .dout(n16439));
  jand g16358(.dina(n8740), .dinb(n6050), .dout(n16440));
  jand g16359(.dina(n8723), .dinb(n5082), .dout(n16441));
  jor  g16360(.dina(n16441), .dinb(n16440), .dout(n16442));
  jor  g16361(.dina(n16442), .dinb(n16439), .dout(n16443));
  jor  g16362(.dina(n16443), .dinb(n16438), .dout(n16444));
  jxor g16363(.dina(n16444), .dinb(n16437), .dout(n16445));
  jxor g16364(.dina(n16445), .dinb(n16421), .dout(n16446));
  jnot g16365(.din(n16446), .dout(n16447));
  jand g16366(.dina(n9886), .dinb(n2936), .dout(n16448));
  jand g16367(.dina(n9655), .dinb(n2943), .dout(n16449));
  jand g16368(.dina(n9656), .dinb(n2940), .dout(n16450));
  jand g16369(.dina(n9250), .dinb(n3684), .dout(n16451));
  jor  g16370(.dina(n16451), .dinb(n16450), .dout(n16452));
  jor  g16371(.dina(n16452), .dinb(n16449), .dout(n16453));
  jor  g16372(.dina(n16453), .dinb(n16448), .dout(n16454));
  jxor g16373(.dina(n16454), .dinb(n93), .dout(n16455));
  jxor g16374(.dina(n16455), .dinb(n16447), .dout(n16456));
  jxor g16375(.dina(n16456), .dinb(n16418), .dout(n16457));
  jnot g16376(.din(n16457), .dout(n16458));
  jand g16377(.dina(n10862), .dinb(n71), .dout(n16459));
  jand g16378(.dina(n10647), .dinb(n796), .dout(n16460));
  jand g16379(.dina(n10305), .dinb(n731), .dout(n16461));
  jand g16380(.dina(n9872), .dinb(n1806), .dout(n16462));
  jor  g16381(.dina(n16462), .dinb(n16461), .dout(n16463));
  jor  g16382(.dina(n16463), .dinb(n16460), .dout(n16464));
  jor  g16383(.dina(n16464), .dinb(n16459), .dout(n16465));
  jxor g16384(.dina(n16465), .dinb(n77), .dout(n16466));
  jxor g16385(.dina(n16466), .dinb(n16458), .dout(n16467));
  jxor g16386(.dina(n16467), .dinb(n16413), .dout(n16468));
  jand g16387(.dina(n11308), .dinb(n806), .dout(n16469));
  jand g16388(.dina(n11306), .dinb(n1620), .dout(n16470));
  jand g16389(.dina(n10836), .dinb(n1612), .dout(n16471));
  jand g16390(.dina(n10640), .dinb(n1644), .dout(n16472));
  jor  g16391(.dina(n16472), .dinb(n16471), .dout(n16473));
  jor  g16392(.dina(n16473), .dinb(n16470), .dout(n16474));
  jor  g16393(.dina(n16474), .dinb(n16469), .dout(n16475));
  jxor g16394(.dina(n16475), .dinb(\a[23] ), .dout(n16476));
  jxor g16395(.dina(n16476), .dinb(n16468), .dout(n16477));
  jxor g16396(.dina(n16477), .dinb(n16408), .dout(n16478));
  jnot g16397(.din(n16478), .dout(n16479));
  jand g16398(.dina(n11800), .dinb(n1819), .dout(n16480));
  jand g16399(.dina(n11646), .dinb(n2180), .dout(n16481));
  jand g16400(.dina(n11798), .dinb(n2243), .dout(n16482));
  jor  g16401(.dina(n16482), .dinb(n16481), .dout(n16483));
  jand g16402(.dina(n11647), .dinb(n2185), .dout(n16484));
  jor  g16403(.dina(n16484), .dinb(n16483), .dout(n16485));
  jor  g16404(.dina(n16485), .dinb(n16480), .dout(n16486));
  jxor g16405(.dina(n16486), .dinb(n2196), .dout(n16487));
  jxor g16406(.dina(n16487), .dinb(n16479), .dout(n16488));
  jxor g16407(.dina(n16488), .dinb(n16403), .dout(n16489));
  jand g16408(.dina(n12684), .dinb(n2743), .dout(n16490));
  jand g16409(.dina(n12536), .dinb(n2752), .dout(n16491));
  jand g16410(.dina(n12547), .dinb(n2748), .dout(n16492));
  jand g16411(.dina(n12282), .dinb(n2757), .dout(n16493));
  jor  g16412(.dina(n16493), .dinb(n16492), .dout(n16494));
  jor  g16413(.dina(n16494), .dinb(n16491), .dout(n16495));
  jor  g16414(.dina(n16495), .dinb(n16490), .dout(n16496));
  jxor g16415(.dina(n16496), .dinb(n2441), .dout(n16497));
  jxor g16416(.dina(n16497), .dinb(n16489), .dout(n16498));
  jxor g16417(.dina(n16498), .dinb(n16398), .dout(n16499));
  jand g16418(.dina(n13639), .dinb(n3423), .dout(n16500));
  jand g16419(.dina(n13478), .dinb(n3569), .dout(n16501));
  jand g16420(.dina(n13248), .dinb(n3428), .dout(n16502));
  jand g16421(.dina(n12669), .dinb(n3210), .dout(n16503));
  jor  g16422(.dina(n16503), .dinb(n16502), .dout(n16504));
  jor  g16423(.dina(n16504), .dinb(n16501), .dout(n16505));
  jor  g16424(.dina(n16505), .dinb(n16500), .dout(n16506));
  jxor g16425(.dina(n16506), .dinb(n3473), .dout(n16507));
  jxor g16426(.dina(n16507), .dinb(n16499), .dout(n16508));
  jnot g16427(.din(n16508), .dout(n16509));
  jxor g16428(.dina(n16509), .dinb(n16395), .dout(n16510));
  jand g16429(.dina(n14251), .dinb(n4022), .dout(n16511));
  jand g16430(.dina(n13614), .dinb(n4027), .dout(n16512));
  jand g16431(.dina(n14249), .dinb(n4220), .dout(n16513));
  jor  g16432(.dina(n16513), .dinb(n16512), .dout(n16514));
  jand g16433(.dina(n13469), .dinb(n3870), .dout(n16515));
  jor  g16434(.dina(n16515), .dinb(n16514), .dout(n16516));
  jor  g16435(.dina(n16516), .dinb(n16511), .dout(n16517));
  jxor g16436(.dina(n16517), .dinb(n4050), .dout(n16518));
  jxor g16437(.dina(n16518), .dinb(n16510), .dout(n16519));
  jnot g16438(.din(n16519), .dout(n16520));
  jxor g16439(.dina(n16520), .dinb(n16391), .dout(n16521));
  jand g16440(.dina(n14551), .dinb(n4691), .dout(n16522));
  jand g16441(.dina(n14447), .dinb(n4696), .dout(n16523));
  jand g16442(.dina(n14549), .dinb(n4941), .dout(n16524));
  jor  g16443(.dina(n16524), .dinb(n16523), .dout(n16525));
  jand g16444(.dina(n14448), .dinb(n4701), .dout(n16526));
  jor  g16445(.dina(n16526), .dinb(n16525), .dout(n16527));
  jor  g16446(.dina(n16527), .dinb(n16522), .dout(n16528));
  jxor g16447(.dina(n16528), .dinb(n4713), .dout(n16529));
  jxor g16448(.dina(n16529), .dinb(n16521), .dout(n16530));
  jxor g16449(.dina(n16530), .dinb(n16387), .dout(n16531));
  jand g16450(.dina(n15831), .dinb(n5280), .dout(n16532));
  jand g16451(.dina(n15829), .dinb(n5814), .dout(n16533));
  jand g16452(.dina(n15567), .dinb(n5531), .dout(n16534));
  jand g16453(.dina(n15315), .dinb(n5536), .dout(n16535));
  jor  g16454(.dina(n16535), .dinb(n16534), .dout(n16536));
  jor  g16455(.dina(n16536), .dinb(n16533), .dout(n16537));
  jor  g16456(.dina(n16537), .dinb(n16532), .dout(n16538));
  jxor g16457(.dina(n16538), .dinb(n5277), .dout(n16539));
  jxor g16458(.dina(n16539), .dinb(n16531), .dout(n16540));
  jxor g16459(.dina(n16540), .dinb(n16379), .dout(n16541));
  jand g16460(.dina(n16343), .dinb(n16082), .dout(n16542));
  jand g16461(.dina(n16344), .dinb(n16321), .dout(n16543));
  jor  g16462(.dina(n16543), .dinb(n16542), .dout(n16544));
  jnot g16463(.din(n16339), .dout(n16546));
  jnot g16464(.din(n16322), .dout(n16547));
  jor  g16465(.dina(n16081), .dinb(n16077), .dout(n16548));
  jand g16466(.dina(n16548), .dinb(n16547), .dout(n16549));
  jnot g16467(.din(n16342), .dout(n16550));
  jor  g16468(.dina(n16550), .dinb(n16549), .dout(n16551));
  jand g16469(.dina(n16551), .dinb(n16546), .dout(n16552));
  jand g16470(.dina(n16334), .dinb(n15811), .dout(n16553));
  jand g16471(.dina(n3336), .dinb(n1713), .dout(n16554));
  jand g16472(.dina(n668), .dinb(n1701), .dout(n16555));
  jand g16473(.dina(n16555), .dinb(n1591), .dout(n16556));
  jand g16474(.dina(n16556), .dinb(n16554), .dout(n16557));
  jand g16475(.dina(n16557), .dinb(n472), .dout(n16558));
  jand g16476(.dina(n2526), .dinb(n1596), .dout(n16559));
  jand g16477(.dina(n16559), .dinb(n1832), .dout(n16560));
  jand g16478(.dina(n16560), .dinb(n16558), .dout(n16561));
  jand g16479(.dina(n1569), .dinb(n817), .dout(n16562));
  jand g16480(.dina(n16562), .dinb(n100), .dout(n16563));
  jand g16481(.dina(n1470), .dinb(n1213), .dout(n16564));
  jand g16482(.dina(n16564), .dinb(n551), .dout(n16565));
  jand g16483(.dina(n1270), .dinb(n493), .dout(n16566));
  jand g16484(.dina(n16566), .dinb(n3108), .dout(n16567));
  jand g16485(.dina(n16567), .dinb(n16565), .dout(n16568));
  jand g16486(.dina(n16568), .dinb(n16563), .dout(n16569));
  jand g16487(.dina(n16569), .dinb(n1339), .dout(n16570));
  jand g16488(.dina(n16570), .dinb(n16561), .dout(n16571));
  jand g16489(.dina(n16571), .dinb(n3402), .dout(n16572));
  jand g16490(.dina(n16572), .dinb(n14291), .dout(n16573));
  jand g16491(.dina(n14323), .dinb(n7670), .dout(n16589));
  jand g16492(.dina(n16589), .dinb(n24501), .dout(n16590));
  jxor g16493(.dina(n16590), .dinb(n16553), .dout(n16591));
  jxor g16494(.dina(n16591), .dinb(n16552), .dout(n16592));
  jxor g16495(.dina(n16592), .dinb(n16343), .dout(n16593));
  jxor g16496(.dina(n16593), .dinb(n16544), .dout(n16594));
  jand g16497(.dina(n16594), .dinb(n6495), .dout(n16595));
  jand g16498(.dina(n16592), .dinb(n6503), .dout(n16596));
  jand g16499(.dina(n16343), .dinb(n6506), .dout(n16597));
  jand g16500(.dina(n16082), .dinb(n6500), .dout(n16598));
  jor  g16501(.dina(n16598), .dinb(n16597), .dout(n16599));
  jor  g16502(.dina(n16599), .dinb(n16596), .dout(n16600));
  jor  g16503(.dina(n16600), .dinb(n16595), .dout(n16601));
  jxor g16504(.dina(n16601), .dinb(n6219), .dout(n16602));
  jxor g16505(.dina(n16602), .dinb(n16541), .dout(n16603));
  jxor g16506(.dina(n16603), .dinb(n16375), .dout(n16604));
  jxor g16507(.dina(n16604), .dinb(n16355), .dout(n16605));
  jxor g16508(.dina(n16605), .dinb(n16371), .dout(n16606));
  jand g16509(.dina(n16606), .dinb(n806), .dout(n16607));
  jand g16510(.dina(n16355), .dinb(n1612), .dout(n16608));
  jand g16511(.dina(n16604), .dinb(n1620), .dout(n16609));
  jor  g16512(.dina(n16609), .dinb(n16608), .dout(n16610));
  jand g16513(.dina(n16360), .dinb(n1644), .dout(n16611));
  jor  g16514(.dina(n16611), .dinb(n16610), .dout(n16612));
  jor  g16515(.dina(n16612), .dinb(n16607), .dout(n16613));
  jxor g16516(.dina(n16613), .dinb(n65), .dout(n16614));
  jor  g16517(.dina(n16614), .dinb(n15858), .dout(n16615));
  jxor g16518(.dina(n16369), .dinb(n16368), .dout(n16616));
  jand g16519(.dina(n16616), .dinb(n806), .dout(n16617));
  jand g16520(.dina(n16360), .dinb(n1612), .dout(n16618));
  jand g16521(.dina(n16355), .dinb(n1620), .dout(n16619));
  jor  g16522(.dina(n16619), .dinb(n16618), .dout(n16620));
  jand g16523(.dina(n15841), .dinb(n1644), .dout(n16621));
  jor  g16524(.dina(n16621), .dinb(n16620), .dout(n16622));
  jor  g16525(.dina(n16622), .dinb(n16617), .dout(n16623));
  jxor g16526(.dina(n16623), .dinb(n65), .dout(n16624));
  jnot g16527(.din(n16624), .dout(n16625));
  jor  g16528(.dina(n15339), .dinb(n77), .dout(n16626));
  jxor g16529(.dina(n16626), .dinb(n15588), .dout(n16627));
  jand g16530(.dina(n16627), .dinb(n16625), .dout(n16628));
  jand g16531(.dina(n15336), .dinb(\a[26] ), .dout(n16629));
  jxor g16532(.dina(n16629), .dinb(n15334), .dout(n16630));
  jnot g16533(.din(n16630), .dout(n16631));
  jxor g16534(.dina(n16366), .dinb(n16365), .dout(n16632));
  jand g16535(.dina(n16632), .dinb(n806), .dout(n16633));
  jand g16536(.dina(n15841), .dinb(n1612), .dout(n16634));
  jand g16537(.dina(n16360), .dinb(n1620), .dout(n16635));
  jor  g16538(.dina(n16635), .dinb(n16634), .dout(n16636));
  jand g16539(.dina(n15579), .dinb(n1644), .dout(n16637));
  jor  g16540(.dina(n16637), .dinb(n16636), .dout(n16638));
  jor  g16541(.dina(n16638), .dinb(n16633), .dout(n16639));
  jxor g16542(.dina(n16639), .dinb(n65), .dout(n16640));
  jor  g16543(.dina(n16640), .dinb(n16631), .dout(n16641));
  jand g16544(.dina(n15329), .dinb(n806), .dout(n16642));
  jand g16545(.dina(n15020), .dinb(n1612), .dout(n16643));
  jand g16546(.dina(n15327), .dinb(n1620), .dout(n16644));
  jor  g16547(.dina(n16644), .dinb(n16643), .dout(n16645));
  jor  g16548(.dina(n16645), .dinb(n16642), .dout(n16646));
  jnot g16549(.din(n16646), .dout(n16647));
  jand g16550(.dina(n15020), .dinb(n804), .dout(n16648));
  jnot g16551(.din(n16648), .dout(n16649));
  jand g16552(.dina(n16649), .dinb(\a[23] ), .dout(n16650));
  jand g16553(.dina(n16650), .dinb(n16647), .dout(n16651));
  jand g16554(.dina(n15580), .dinb(n806), .dout(n16652));
  jand g16555(.dina(n15327), .dinb(n1612), .dout(n16653));
  jor  g16556(.dina(n16653), .dinb(n16652), .dout(n16654));
  jand g16557(.dina(n15579), .dinb(n1620), .dout(n16655));
  jand g16558(.dina(n15020), .dinb(n1644), .dout(n16656));
  jor  g16559(.dina(n16656), .dinb(n16655), .dout(n16657));
  jor  g16560(.dina(n16657), .dinb(n16654), .dout(n16658));
  jnot g16561(.din(n16658), .dout(n16659));
  jand g16562(.dina(n16659), .dinb(n16651), .dout(n16660));
  jand g16563(.dina(n16660), .dinb(n15336), .dout(n16661));
  jnot g16564(.din(n16661), .dout(n16662));
  jxor g16565(.dina(n16660), .dinb(n15336), .dout(n16663));
  jnot g16566(.din(n16663), .dout(n16664));
  jand g16567(.dina(n15848), .dinb(n806), .dout(n16665));
  jand g16568(.dina(n15579), .dinb(n1612), .dout(n16666));
  jand g16569(.dina(n15841), .dinb(n1620), .dout(n16667));
  jor  g16570(.dina(n16667), .dinb(n16666), .dout(n16668));
  jand g16571(.dina(n15327), .dinb(n1644), .dout(n16669));
  jor  g16572(.dina(n16669), .dinb(n16668), .dout(n16670));
  jor  g16573(.dina(n16670), .dinb(n16665), .dout(n16671));
  jxor g16574(.dina(n16671), .dinb(n65), .dout(n16672));
  jor  g16575(.dina(n16672), .dinb(n16664), .dout(n16673));
  jand g16576(.dina(n16673), .dinb(n16662), .dout(n16674));
  jnot g16577(.din(n16674), .dout(n16675));
  jxor g16578(.dina(n16640), .dinb(n16631), .dout(n16676));
  jand g16579(.dina(n16676), .dinb(n16675), .dout(n16677));
  jnot g16580(.din(n16677), .dout(n16678));
  jand g16581(.dina(n16678), .dinb(n16641), .dout(n16679));
  jnot g16582(.din(n16679), .dout(n16680));
  jxor g16583(.dina(n16627), .dinb(n16625), .dout(n16681));
  jand g16584(.dina(n16681), .dinb(n16680), .dout(n16682));
  jor  g16585(.dina(n16682), .dinb(n16628), .dout(n16683));
  jxor g16586(.dina(n16614), .dinb(n15858), .dout(n16684));
  jand g16587(.dina(n16684), .dinb(n16683), .dout(n16685));
  jnot g16588(.din(n16685), .dout(n16686));
  jand g16589(.dina(n16686), .dinb(n16615), .dout(n16687));
  jnot g16590(.din(n16687), .dout(n16688));
  jand g16591(.dina(n15589), .dinb(n15021), .dout(n16689));
  jnot g16592(.din(n16689), .dout(n16690));
  jor  g16593(.dina(n15856), .dinb(n15591), .dout(n16691));
  jand g16594(.dina(n16691), .dinb(n16690), .dout(n16692));
  jnot g16595(.din(n16692), .dout(n16693));
  jand g16596(.dina(n15329), .dinb(n2936), .dout(n16694));
  jand g16597(.dina(n15020), .dinb(n2940), .dout(n16695));
  jand g16598(.dina(n15327), .dinb(n2943), .dout(n16696));
  jor  g16599(.dina(n16696), .dinb(n16695), .dout(n16697));
  jor  g16600(.dina(n16697), .dinb(n16694), .dout(n16698));
  jnot g16601(.din(n15021), .dout(n16699));
  jor  g16602(.dina(n16699), .dinb(n93), .dout(n16700));
  jxor g16603(.dina(n16700), .dinb(n16698), .dout(n16701));
  jand g16604(.dina(n16632), .dinb(n71), .dout(n16702));
  jand g16605(.dina(n15841), .dinb(n731), .dout(n16703));
  jand g16606(.dina(n16360), .dinb(n796), .dout(n16704));
  jor  g16607(.dina(n16704), .dinb(n16703), .dout(n16705));
  jand g16608(.dina(n15579), .dinb(n1806), .dout(n16706));
  jor  g16609(.dina(n16706), .dinb(n16705), .dout(n16707));
  jor  g16610(.dina(n16707), .dinb(n16702), .dout(n16708));
  jxor g16611(.dina(n16708), .dinb(n77), .dout(n16709));
  jxor g16612(.dina(n16709), .dinb(n16701), .dout(n16710));
  jxor g16613(.dina(n16710), .dinb(n16693), .dout(n16711));
  jnot g16614(.din(n16711), .dout(n16712));
  jand g16615(.dina(n16604), .dinb(n16355), .dout(n16713));
  jand g16616(.dina(n16605), .dinb(n16371), .dout(n16714));
  jor  g16617(.dina(n16714), .dinb(n16713), .dout(n16715));
  jnot g16618(.din(n16541), .dout(n16716));
  jor  g16619(.dina(n16602), .dinb(n16716), .dout(n16717));
  jor  g16620(.dina(n16603), .dinb(n16375), .dout(n16718));
  jand g16621(.dina(n16718), .dinb(n16717), .dout(n16719));
  jor  g16622(.dina(n16539), .dinb(n16531), .dout(n16720));
  jnot g16623(.din(n16110), .dout(n16721));
  jxor g16624(.dina(n16043), .dinb(n16121), .dout(n16722));
  jxor g16625(.dina(n16052), .dinb(n16722), .dout(n16723));
  jor  g16626(.dina(n16723), .dinb(n15867), .dout(n16724));
  jand g16627(.dina(n16724), .dinb(n16721), .dout(n16725));
  jnot g16628(.din(n16113), .dout(n16726));
  jand g16629(.dina(n16043), .dinb(n15871), .dout(n16727));
  jor  g16630(.dina(n16727), .dinb(n16726), .dout(n16728));
  jxor g16631(.dina(n16307), .dinb(n16728), .dout(n16729));
  jxor g16632(.dina(n16316), .dinb(n16729), .dout(n16730));
  jor  g16633(.dina(n16730), .dinb(n16725), .dout(n16731));
  jand g16634(.dina(n16731), .dinb(n16376), .dout(n16732));
  jnot g16635(.din(n16380), .dout(n16733));
  jand g16636(.dina(n16307), .dinb(n16728), .dout(n16734));
  jor  g16637(.dina(n16734), .dinb(n16733), .dout(n16735));
  jxor g16638(.dina(n16530), .dinb(n16735), .dout(n16736));
  jxor g16639(.dina(n16539), .dinb(n16736), .dout(n16737));
  jor  g16640(.dina(n16737), .dinb(n16732), .dout(n16738));
  jand g16641(.dina(n16738), .dinb(n16720), .dout(n16739));
  jor  g16642(.dina(n16529), .dinb(n16521), .dout(n16740));
  jnot g16643(.din(n16740), .dout(n16741));
  jand g16644(.dina(n16530), .dinb(n16735), .dout(n16742));
  jor  g16645(.dina(n16742), .dinb(n16741), .dout(n16743));
  jnot g16646(.din(n16510), .dout(n16744));
  jor  g16647(.dina(n16518), .dinb(n16744), .dout(n16745));
  jor  g16648(.dina(n16519), .dinb(n16391), .dout(n16746));
  jand g16649(.dina(n16746), .dinb(n16745), .dout(n16747));
  jor  g16650(.dina(n16507), .dinb(n16499), .dout(n16748));
  jor  g16651(.dina(n16509), .dinb(n16395), .dout(n16749));
  jand g16652(.dina(n16749), .dinb(n16748), .dout(n16750));
  jnot g16653(.din(n16489), .dout(n16751));
  jor  g16654(.dina(n16497), .dinb(n16751), .dout(n16752));
  jnot g16655(.din(n16498), .dout(n16753));
  jand g16656(.dina(n16753), .dinb(n16398), .dout(n16754));
  jnot g16657(.din(n16754), .dout(n16755));
  jand g16658(.dina(n16755), .dinb(n16752), .dout(n16756));
  jor  g16659(.dina(n16487), .dinb(n16479), .dout(n16757));
  jnot g16660(.din(n16757), .dout(n16758));
  jand g16661(.dina(n16488), .dinb(n16403), .dout(n16759));
  jor  g16662(.dina(n16759), .dinb(n16758), .dout(n16760));
  jand g16663(.dina(n16476), .dinb(n16468), .dout(n16761));
  jand g16664(.dina(n16477), .dinb(n16408), .dout(n16762));
  jor  g16665(.dina(n16762), .dinb(n16761), .dout(n16763));
  jor  g16666(.dina(n16466), .dinb(n16458), .dout(n16764));
  jand g16667(.dina(n16467), .dinb(n16413), .dout(n16765));
  jnot g16668(.din(n16765), .dout(n16766));
  jand g16669(.dina(n16766), .dinb(n16764), .dout(n16767));
  jnot g16670(.din(n16767), .dout(n16768));
  jor  g16671(.dina(n16455), .dinb(n16447), .dout(n16769));
  jand g16672(.dina(n16456), .dinb(n16418), .dout(n16770));
  jnot g16673(.din(n16770), .dout(n16771));
  jand g16674(.dina(n16771), .dinb(n16769), .dout(n16772));
  jnot g16675(.din(n16772), .dout(n16773));
  jand g16676(.dina(n16444), .dinb(n16437), .dout(n16774));
  jand g16677(.dina(n16445), .dinb(n16421), .dout(n16775));
  jor  g16678(.dina(n16775), .dinb(n16774), .dout(n16776));
  jand g16679(.dina(n3149), .dinb(n1471), .dout(n16777));
  jand g16680(.dina(n10739), .dinb(n1700), .dout(n16778));
  jand g16681(.dina(n16778), .dinb(n2024), .dout(n16779));
  jand g16682(.dina(n16779), .dinb(n8143), .dout(n16780));
  jand g16683(.dina(n16780), .dinb(n16777), .dout(n16781));
  jand g16684(.dina(n1565), .dinb(n696), .dout(n16782));
  jand g16685(.dina(n16782), .dinb(n716), .dout(n16783));
  jand g16686(.dina(n2477), .dinb(n1824), .dout(n16784));
  jand g16687(.dina(n983), .dinb(n472), .dout(n16785));
  jand g16688(.dina(n553), .dinb(n964), .dout(n16786));
  jand g16689(.dina(n16786), .dinb(n16785), .dout(n16787));
  jand g16690(.dina(n16787), .dinb(n1016), .dout(n16788));
  jand g16691(.dina(n16788), .dinb(n16784), .dout(n16789));
  jand g16692(.dina(n13551), .dinb(n560), .dout(n16790));
  jand g16693(.dina(n16790), .dinb(n16789), .dout(n16791));
  jand g16694(.dina(n16791), .dinb(n16783), .dout(n16792));
  jand g16695(.dina(n16792), .dinb(n16781), .dout(n16793));
  jand g16696(.dina(n3364), .dinb(n685), .dout(n16794));
  jand g16697(.dina(n16794), .dinb(n114), .dout(n16795));
  jand g16698(.dina(n16795), .dinb(n1096), .dout(n16796));
  jand g16699(.dina(n16796), .dinb(n3116), .dout(n16797));
  jand g16700(.dina(n16797), .dinb(n16793), .dout(n16798));
  jand g16701(.dina(n3026), .dinb(n2483), .dout(n16799));
  jand g16702(.dina(n16799), .dinb(n1055), .dout(n16800));
  jand g16703(.dina(n16800), .dinb(n11224), .dout(n16801));
  jand g16704(.dina(n3214), .dinb(n3190), .dout(n16802));
  jand g16705(.dina(n16802), .dinb(n16801), .dout(n16803));
  jand g16706(.dina(n16803), .dinb(n16798), .dout(n16804));
  jand g16707(.dina(n1162), .dinb(n917), .dout(n16805));
  jand g16708(.dina(n1846), .dinb(n175), .dout(n16806));
  jand g16709(.dina(n16806), .dinb(n16805), .dout(n16807));
  jand g16710(.dina(n16807), .dinb(n7244), .dout(n16808));
  jand g16711(.dina(n3092), .dinb(n1273), .dout(n16809));
  jand g16712(.dina(n16809), .dinb(n1443), .dout(n16810));
  jand g16713(.dina(n16810), .dinb(n16808), .dout(n16811));
  jand g16714(.dina(n16811), .dinb(n16804), .dout(n16812));
  jnot g16715(.din(n16812), .dout(n16813));
  jand g16716(.dina(n9252), .dinb(n5076), .dout(n16814));
  jand g16717(.dina(n9250), .dinb(n5084), .dout(n16815));
  jand g16718(.dina(n8723), .dinb(n6050), .dout(n16816));
  jand g16719(.dina(n8936), .dinb(n5082), .dout(n16817));
  jor  g16720(.dina(n16817), .dinb(n16816), .dout(n16818));
  jor  g16721(.dina(n16818), .dinb(n16815), .dout(n16819));
  jor  g16722(.dina(n16819), .dinb(n16814), .dout(n16820));
  jxor g16723(.dina(n16820), .dinb(n16813), .dout(n16821));
  jxor g16724(.dina(n16821), .dinb(n16776), .dout(n16822));
  jnot g16725(.din(n16822), .dout(n16823));
  jand g16726(.dina(n9874), .dinb(n2936), .dout(n16824));
  jand g16727(.dina(n9655), .dinb(n2940), .dout(n16825));
  jand g16728(.dina(n9872), .dinb(n2943), .dout(n16826));
  jor  g16729(.dina(n16826), .dinb(n16825), .dout(n16827));
  jand g16730(.dina(n9656), .dinb(n3684), .dout(n16828));
  jor  g16731(.dina(n16828), .dinb(n16827), .dout(n16829));
  jor  g16732(.dina(n16829), .dinb(n16824), .dout(n16830));
  jxor g16733(.dina(n16830), .dinb(n93), .dout(n16831));
  jxor g16734(.dina(n16831), .dinb(n16823), .dout(n16832));
  jxor g16735(.dina(n16832), .dinb(n16773), .dout(n16833));
  jnot g16736(.din(n16833), .dout(n16834));
  jand g16737(.dina(n10850), .dinb(n71), .dout(n16835));
  jand g16738(.dina(n10640), .dinb(n796), .dout(n16836));
  jand g16739(.dina(n10647), .dinb(n731), .dout(n16837));
  jand g16740(.dina(n10305), .dinb(n1806), .dout(n16838));
  jor  g16741(.dina(n16838), .dinb(n16837), .dout(n16839));
  jor  g16742(.dina(n16839), .dinb(n16836), .dout(n16840));
  jor  g16743(.dina(n16840), .dinb(n16835), .dout(n16841));
  jxor g16744(.dina(n16841), .dinb(n77), .dout(n16842));
  jxor g16745(.dina(n16842), .dinb(n16834), .dout(n16843));
  jxor g16746(.dina(n16843), .dinb(n16768), .dout(n16844));
  jnot g16747(.din(n16844), .dout(n16845));
  jand g16748(.dina(n11824), .dinb(n806), .dout(n16846));
  jand g16749(.dina(n11647), .dinb(n1620), .dout(n16847));
  jand g16750(.dina(n11306), .dinb(n1612), .dout(n16848));
  jand g16751(.dina(n10836), .dinb(n1644), .dout(n16849));
  jor  g16752(.dina(n16849), .dinb(n16848), .dout(n16850));
  jor  g16753(.dina(n16850), .dinb(n16847), .dout(n16851));
  jor  g16754(.dina(n16851), .dinb(n16846), .dout(n16852));
  jxor g16755(.dina(n16852), .dinb(n65), .dout(n16853));
  jxor g16756(.dina(n16853), .dinb(n16845), .dout(n16854));
  jxor g16757(.dina(n16854), .dinb(n16763), .dout(n16855));
  jnot g16758(.din(n16855), .dout(n16856));
  jand g16759(.dina(n12284), .dinb(n1819), .dout(n16857));
  jand g16760(.dina(n11798), .dinb(n2180), .dout(n16858));
  jand g16761(.dina(n12282), .dinb(n2243), .dout(n16859));
  jor  g16762(.dina(n16859), .dinb(n16858), .dout(n16860));
  jand g16763(.dina(n11646), .dinb(n2185), .dout(n16861));
  jor  g16764(.dina(n16861), .dinb(n16860), .dout(n16862));
  jor  g16765(.dina(n16862), .dinb(n16857), .dout(n16863));
  jxor g16766(.dina(n16863), .dinb(n2196), .dout(n16864));
  jxor g16767(.dina(n16864), .dinb(n16856), .dout(n16865));
  jxor g16768(.dina(n16865), .dinb(n16760), .dout(n16866));
  jand g16769(.dina(n12671), .dinb(n2743), .dout(n16867));
  jand g16770(.dina(n12669), .dinb(n2752), .dout(n16868));
  jand g16771(.dina(n12536), .dinb(n2748), .dout(n16869));
  jand g16772(.dina(n12547), .dinb(n2757), .dout(n16870));
  jor  g16773(.dina(n16870), .dinb(n16869), .dout(n16871));
  jor  g16774(.dina(n16871), .dinb(n16868), .dout(n16872));
  jor  g16775(.dina(n16872), .dinb(n16867), .dout(n16873));
  jxor g16776(.dina(n16873), .dinb(n2441), .dout(n16874));
  jxor g16777(.dina(n16874), .dinb(n16866), .dout(n16875));
  jxor g16778(.dina(n16875), .dinb(n16756), .dout(n16876));
  jnot g16779(.din(n16876), .dout(n16877));
  jand g16780(.dina(n13627), .dinb(n3423), .dout(n16878));
  jand g16781(.dina(n13478), .dinb(n3428), .dout(n16879));
  jand g16782(.dina(n13469), .dinb(n3569), .dout(n16880));
  jor  g16783(.dina(n16880), .dinb(n16879), .dout(n16881));
  jand g16784(.dina(n13248), .dinb(n3210), .dout(n16882));
  jor  g16785(.dina(n16882), .dinb(n16881), .dout(n16883));
  jor  g16786(.dina(n16883), .dinb(n16878), .dout(n16884));
  jxor g16787(.dina(n16884), .dinb(n3473), .dout(n16885));
  jxor g16788(.dina(n16885), .dinb(n16877), .dout(n16886));
  jnot g16789(.din(n16886), .dout(n16887));
  jxor g16790(.dina(n16887), .dinb(n16750), .dout(n16888));
  jand g16791(.dina(n14579), .dinb(n4022), .dout(n16889));
  jand g16792(.dina(n14448), .dinb(n4220), .dout(n16890));
  jand g16793(.dina(n14249), .dinb(n4027), .dout(n16891));
  jand g16794(.dina(n13614), .dinb(n3870), .dout(n16892));
  jor  g16795(.dina(n16892), .dinb(n16891), .dout(n16893));
  jor  g16796(.dina(n16893), .dinb(n16890), .dout(n16894));
  jor  g16797(.dina(n16894), .dinb(n16889), .dout(n16895));
  jxor g16798(.dina(n16895), .dinb(n4050), .dout(n16896));
  jxor g16799(.dina(n16896), .dinb(n16888), .dout(n16897));
  jnot g16800(.din(n16897), .dout(n16898));
  jxor g16801(.dina(n16898), .dinb(n16747), .dout(n16899));
  jand g16802(.dina(n15317), .dinb(n4691), .dout(n16900));
  jand g16803(.dina(n14549), .dinb(n4696), .dout(n16901));
  jand g16804(.dina(n15315), .dinb(n4941), .dout(n16902));
  jor  g16805(.dina(n16902), .dinb(n16901), .dout(n16903));
  jand g16806(.dina(n14447), .dinb(n4701), .dout(n16904));
  jor  g16807(.dina(n16904), .dinb(n16903), .dout(n16905));
  jor  g16808(.dina(n16905), .dinb(n16900), .dout(n16906));
  jxor g16809(.dina(n16906), .dinb(n4713), .dout(n16907));
  jxor g16810(.dina(n16907), .dinb(n16899), .dout(n16908));
  jxor g16811(.dina(n16908), .dinb(n16743), .dout(n16909));
  jand g16812(.dina(n16084), .dinb(n5280), .dout(n16910));
  jand g16813(.dina(n15829), .dinb(n5531), .dout(n16911));
  jand g16814(.dina(n16082), .dinb(n5814), .dout(n16912));
  jor  g16815(.dina(n16912), .dinb(n16911), .dout(n16913));
  jand g16816(.dina(n15567), .dinb(n5536), .dout(n16914));
  jor  g16817(.dina(n16914), .dinb(n16913), .dout(n16915));
  jor  g16818(.dina(n16915), .dinb(n16910), .dout(n16916));
  jxor g16819(.dina(n16916), .dinb(n5277), .dout(n16917));
  jxor g16820(.dina(n16917), .dinb(n16909), .dout(n16918));
  jxor g16821(.dina(n16918), .dinb(n16739), .dout(n16919));
  jand g16822(.dina(n16592), .dinb(n16343), .dout(n16920));
  jand g16823(.dina(n16593), .dinb(n16544), .dout(n16921));
  jor  g16824(.dina(n16921), .dinb(n16920), .dout(n16922));
  jor  g16825(.dina(n16591), .dinb(n16552), .dout(n16924));
  jand g16826(.dina(n16590), .dinb(n16553), .dout(n16925));
  jand g16827(.dina(n16925), .dinb(n16552), .dout(n16926));
  jnot g16828(.din(n16926), .dout(n16927));
  jand g16829(.dina(n16927), .dinb(n16924), .dout(n16928));
  jxor g16830(.dina(n16928), .dinb(n16592), .dout(n16929));
  jxor g16831(.dina(n16929), .dinb(n16922), .dout(n16930));
  jand g16832(.dina(n16930), .dinb(n6495), .dout(n16931));
  jand g16833(.dina(n16592), .dinb(n6506), .dout(n16932));
  jand g16834(.dina(n16928), .dinb(n6503), .dout(n16933));
  jor  g16835(.dina(n16933), .dinb(n16932), .dout(n16934));
  jand g16836(.dina(n16343), .dinb(n6500), .dout(n16935));
  jor  g16837(.dina(n16935), .dinb(n16934), .dout(n16936));
  jor  g16838(.dina(n16936), .dinb(n16931), .dout(n16937));
  jxor g16839(.dina(n16937), .dinb(n6219), .dout(n16938));
  jxor g16840(.dina(n16938), .dinb(n16919), .dout(n16939));
  jxor g16841(.dina(n16939), .dinb(n16719), .dout(n16940));
  jxor g16842(.dina(n16940), .dinb(n16604), .dout(n16941));
  jxor g16843(.dina(n16941), .dinb(n16715), .dout(n16942));
  jand g16844(.dina(n16942), .dinb(n806), .dout(n16943));
  jand g16845(.dina(n16940), .dinb(n1620), .dout(n16944));
  jand g16846(.dina(n16355), .dinb(n1644), .dout(n16945));
  jand g16847(.dina(n16604), .dinb(n1612), .dout(n16946));
  jor  g16848(.dina(n16946), .dinb(n16945), .dout(n16947));
  jor  g16849(.dina(n16947), .dinb(n16944), .dout(n16948));
  jor  g16850(.dina(n16948), .dinb(n16943), .dout(n16949));
  jxor g16851(.dina(n16949), .dinb(n65), .dout(n16950));
  jxor g16852(.dina(n16950), .dinb(n16712), .dout(n16951));
  jxor g16853(.dina(n16951), .dinb(n16688), .dout(n16952));
  jnot g16854(.din(n16952), .dout(n16953));
  jor  g16855(.dina(n16907), .dinb(n16899), .dout(n16954));
  jnot g16856(.din(n16954), .dout(n16955));
  jand g16857(.dina(n16908), .dinb(n16743), .dout(n16956));
  jor  g16858(.dina(n16956), .dinb(n16955), .dout(n16957));
  jnot g16859(.din(n16888), .dout(n16958));
  jor  g16860(.dina(n16896), .dinb(n16958), .dout(n16959));
  jor  g16861(.dina(n16897), .dinb(n16747), .dout(n16960));
  jand g16862(.dina(n16960), .dinb(n16959), .dout(n16961));
  jor  g16863(.dina(n16885), .dinb(n16877), .dout(n16962));
  jor  g16864(.dina(n16887), .dinb(n16750), .dout(n16963));
  jand g16865(.dina(n16963), .dinb(n16962), .dout(n16964));
  jnot g16866(.din(n16866), .dout(n16965));
  jor  g16867(.dina(n16874), .dinb(n16965), .dout(n16966));
  jor  g16868(.dina(n16875), .dinb(n16756), .dout(n16967));
  jand g16869(.dina(n16967), .dinb(n16966), .dout(n16968));
  jor  g16870(.dina(n16864), .dinb(n16856), .dout(n16969));
  jnot g16871(.din(n16969), .dout(n16970));
  jand g16872(.dina(n16865), .dinb(n16760), .dout(n16971));
  jor  g16873(.dina(n16971), .dinb(n16970), .dout(n16972));
  jor  g16874(.dina(n16853), .dinb(n16845), .dout(n16973));
  jand g16875(.dina(n16854), .dinb(n16763), .dout(n16974));
  jnot g16876(.din(n16974), .dout(n16975));
  jand g16877(.dina(n16975), .dinb(n16973), .dout(n16976));
  jnot g16878(.din(n16976), .dout(n16977));
  jor  g16879(.dina(n16842), .dinb(n16834), .dout(n16978));
  jand g16880(.dina(n16843), .dinb(n16768), .dout(n16979));
  jnot g16881(.din(n16979), .dout(n16980));
  jand g16882(.dina(n16980), .dinb(n16978), .dout(n16981));
  jnot g16883(.din(n16981), .dout(n16982));
  jor  g16884(.dina(n16831), .dinb(n16823), .dout(n16983));
  jand g16885(.dina(n16832), .dinb(n16773), .dout(n16984));
  jnot g16886(.din(n16984), .dout(n16985));
  jand g16887(.dina(n16985), .dinb(n16983), .dout(n16986));
  jnot g16888(.din(n16986), .dout(n16987));
  jand g16889(.dina(n16820), .dinb(n16813), .dout(n16988));
  jand g16890(.dina(n16821), .dinb(n16776), .dout(n16989));
  jor  g16891(.dina(n16989), .dinb(n16988), .dout(n16990));
  jand g16892(.dina(n456), .dinb(n510), .dout(n16991));
  jand g16893(.dina(n978), .dinb(n1270), .dout(n16992));
  jand g16894(.dina(n16992), .dinb(n16991), .dout(n16993));
  jand g16895(.dina(n1559), .dinb(n584), .dout(n16994));
  jand g16896(.dina(n16994), .dinb(n16993), .dout(n16995));
  jand g16897(.dina(n5379), .dinb(n818), .dout(n16996));
  jand g16898(.dina(n16996), .dinb(n13313), .dout(n16997));
  jand g16899(.dina(n16997), .dinb(n2077), .dout(n16998));
  jand g16900(.dina(n16998), .dinb(n16995), .dout(n16999));
  jand g16901(.dina(n16999), .dinb(n9140), .dout(n17000));
  jand g16902(.dina(n17000), .dinb(n2707), .dout(n17001));
  jand g16903(.dina(n4532), .dinb(n3996), .dout(n17002));
  jand g16904(.dina(n17002), .dinb(n1509), .dout(n17003));
  jand g16905(.dina(n17003), .dinb(n14484), .dout(n17004));
  jand g16906(.dina(n17004), .dinb(n5193), .dout(n17005));
  jand g16907(.dina(n17005), .dinb(n17001), .dout(n17006));
  jnot g16908(.din(n17006), .dout(n17007));
  jand g16909(.dina(n9898), .dinb(n5076), .dout(n17008));
  jand g16910(.dina(n9656), .dinb(n5084), .dout(n17009));
  jand g16911(.dina(n8936), .dinb(n6050), .dout(n17010));
  jand g16912(.dina(n9250), .dinb(n5082), .dout(n17011));
  jor  g16913(.dina(n17011), .dinb(n17010), .dout(n17012));
  jor  g16914(.dina(n17012), .dinb(n17009), .dout(n17013));
  jor  g16915(.dina(n17013), .dinb(n17008), .dout(n17014));
  jxor g16916(.dina(n17014), .dinb(n17007), .dout(n17015));
  jxor g16917(.dina(n17015), .dinb(n16990), .dout(n17016));
  jnot g16918(.din(n17016), .dout(n17017));
  jand g16919(.dina(n10307), .dinb(n2936), .dout(n17018));
  jand g16920(.dina(n10305), .dinb(n2943), .dout(n17019));
  jand g16921(.dina(n9872), .dinb(n2940), .dout(n17020));
  jand g16922(.dina(n9655), .dinb(n3684), .dout(n17021));
  jor  g16923(.dina(n17021), .dinb(n17020), .dout(n17022));
  jor  g16924(.dina(n17022), .dinb(n17019), .dout(n17023));
  jor  g16925(.dina(n17023), .dinb(n17018), .dout(n17024));
  jxor g16926(.dina(n17024), .dinb(n93), .dout(n17025));
  jxor g16927(.dina(n17025), .dinb(n17017), .dout(n17026));
  jxor g16928(.dina(n17026), .dinb(n16987), .dout(n17027));
  jnot g16929(.din(n17027), .dout(n17028));
  jand g16930(.dina(n10838), .dinb(n71), .dout(n17029));
  jand g16931(.dina(n10836), .dinb(n796), .dout(n17030));
  jand g16932(.dina(n10640), .dinb(n731), .dout(n17031));
  jand g16933(.dina(n10647), .dinb(n1806), .dout(n17032));
  jor  g16934(.dina(n17032), .dinb(n17031), .dout(n17033));
  jor  g16935(.dina(n17033), .dinb(n17030), .dout(n17034));
  jor  g16936(.dina(n17034), .dinb(n17029), .dout(n17035));
  jxor g16937(.dina(n17035), .dinb(n77), .dout(n17036));
  jxor g16938(.dina(n17036), .dinb(n17028), .dout(n17037));
  jxor g16939(.dina(n17037), .dinb(n16982), .dout(n17038));
  jnot g16940(.din(n17038), .dout(n17039));
  jand g16941(.dina(n11812), .dinb(n806), .dout(n17040));
  jand g16942(.dina(n11647), .dinb(n1612), .dout(n17041));
  jand g16943(.dina(n11646), .dinb(n1620), .dout(n17042));
  jor  g16944(.dina(n17042), .dinb(n17041), .dout(n17043));
  jand g16945(.dina(n11306), .dinb(n1644), .dout(n17044));
  jor  g16946(.dina(n17044), .dinb(n17043), .dout(n17045));
  jor  g16947(.dina(n17045), .dinb(n17040), .dout(n17046));
  jxor g16948(.dina(n17046), .dinb(n65), .dout(n17047));
  jxor g16949(.dina(n17047), .dinb(n17039), .dout(n17048));
  jxor g16950(.dina(n17048), .dinb(n16977), .dout(n17049));
  jnot g16951(.din(n17049), .dout(n17050));
  jand g16952(.dina(n12696), .dinb(n1819), .dout(n17051));
  jand g16953(.dina(n12547), .dinb(n2243), .dout(n17052));
  jand g16954(.dina(n12282), .dinb(n2180), .dout(n17053));
  jand g16955(.dina(n11798), .dinb(n2185), .dout(n17054));
  jor  g16956(.dina(n17054), .dinb(n17053), .dout(n17055));
  jor  g16957(.dina(n17055), .dinb(n17052), .dout(n17056));
  jor  g16958(.dina(n17056), .dinb(n17051), .dout(n17057));
  jxor g16959(.dina(n17057), .dinb(n2196), .dout(n17058));
  jxor g16960(.dina(n17058), .dinb(n17050), .dout(n17059));
  jxor g16961(.dina(n17059), .dinb(n16972), .dout(n17060));
  jand g16962(.dina(n13250), .dinb(n2743), .dout(n17061));
  jand g16963(.dina(n13248), .dinb(n2752), .dout(n17062));
  jand g16964(.dina(n12669), .dinb(n2748), .dout(n17063));
  jand g16965(.dina(n12536), .dinb(n2757), .dout(n17064));
  jor  g16966(.dina(n17064), .dinb(n17063), .dout(n17065));
  jor  g16967(.dina(n17065), .dinb(n17062), .dout(n17066));
  jor  g16968(.dina(n17066), .dinb(n17061), .dout(n17067));
  jxor g16969(.dina(n17067), .dinb(n2441), .dout(n17068));
  jxor g16970(.dina(n17068), .dinb(n17060), .dout(n17069));
  jxor g16971(.dina(n17069), .dinb(n16968), .dout(n17070));
  jnot g16972(.din(n17070), .dout(n17071));
  jand g16973(.dina(n13616), .dinb(n3423), .dout(n17072));
  jand g16974(.dina(n13469), .dinb(n3428), .dout(n17073));
  jand g16975(.dina(n13614), .dinb(n3569), .dout(n17074));
  jor  g16976(.dina(n17074), .dinb(n17073), .dout(n17075));
  jand g16977(.dina(n13478), .dinb(n3210), .dout(n17076));
  jor  g16978(.dina(n17076), .dinb(n17075), .dout(n17077));
  jor  g16979(.dina(n17077), .dinb(n17072), .dout(n17078));
  jxor g16980(.dina(n17078), .dinb(n3473), .dout(n17079));
  jxor g16981(.dina(n17079), .dinb(n17071), .dout(n17080));
  jnot g16982(.din(n17080), .dout(n17081));
  jxor g16983(.dina(n17081), .dinb(n16964), .dout(n17082));
  jand g16984(.dina(n14562), .dinb(n4022), .dout(n17083));
  jand g16985(.dina(n14448), .dinb(n4027), .dout(n17084));
  jand g16986(.dina(n14447), .dinb(n4220), .dout(n17085));
  jor  g16987(.dina(n17085), .dinb(n17084), .dout(n17086));
  jand g16988(.dina(n14249), .dinb(n3870), .dout(n17087));
  jor  g16989(.dina(n17087), .dinb(n17086), .dout(n17088));
  jor  g16990(.dina(n17088), .dinb(n17083), .dout(n17089));
  jxor g16991(.dina(n17089), .dinb(n4050), .dout(n17090));
  jxor g16992(.dina(n17090), .dinb(n17082), .dout(n17091));
  jnot g16993(.din(n17091), .dout(n17092));
  jxor g16994(.dina(n17092), .dinb(n16961), .dout(n17093));
  jand g16995(.dina(n15569), .dinb(n4691), .dout(n17094));
  jand g16996(.dina(n15315), .dinb(n4696), .dout(n17095));
  jand g16997(.dina(n15567), .dinb(n4941), .dout(n17096));
  jor  g16998(.dina(n17096), .dinb(n17095), .dout(n17097));
  jand g16999(.dina(n14549), .dinb(n4701), .dout(n17098));
  jor  g17000(.dina(n17098), .dinb(n17097), .dout(n17099));
  jor  g17001(.dina(n17099), .dinb(n17094), .dout(n17100));
  jxor g17002(.dina(n17100), .dinb(n4713), .dout(n17101));
  jxor g17003(.dina(n17101), .dinb(n17093), .dout(n17102));
  jxor g17004(.dina(n17102), .dinb(n16957), .dout(n17103));
  jnot g17005(.din(n17103), .dout(n17104));
  jand g17006(.dina(n16345), .dinb(n5280), .dout(n17105));
  jand g17007(.dina(n16082), .dinb(n5531), .dout(n17106));
  jand g17008(.dina(n16343), .dinb(n5814), .dout(n17107));
  jor  g17009(.dina(n17107), .dinb(n17106), .dout(n17108));
  jand g17010(.dina(n15829), .dinb(n5536), .dout(n17109));
  jor  g17011(.dina(n17109), .dinb(n17108), .dout(n17110));
  jor  g17012(.dina(n17110), .dinb(n17105), .dout(n17111));
  jxor g17013(.dina(n17111), .dinb(n5277), .dout(n17112));
  jor  g17014(.dina(n17112), .dinb(n17104), .dout(n17113));
  jxor g17015(.dina(n16897), .dinb(n16747), .dout(n17114));
  jxor g17016(.dina(n16907), .dinb(n17114), .dout(n17115));
  jxor g17017(.dina(n17115), .dinb(n16743), .dout(n17116));
  jor  g17018(.dina(n16917), .dinb(n17116), .dout(n17117));
  jor  g17019(.dina(n16918), .dinb(n16739), .dout(n17118));
  jand g17020(.dina(n17118), .dinb(n17117), .dout(n17119));
  jxor g17021(.dina(n17112), .dinb(n17103), .dout(n17120));
  jor  g17022(.dina(n17120), .dinb(n17119), .dout(n17121));
  jand g17023(.dina(n17121), .dinb(n17113), .dout(n17122));
  jor  g17024(.dina(n17101), .dinb(n17093), .dout(n17123));
  jnot g17025(.din(n17123), .dout(n17124));
  jand g17026(.dina(n17102), .dinb(n16957), .dout(n17125));
  jor  g17027(.dina(n17125), .dinb(n17124), .dout(n17126));
  jnot g17028(.din(n17082), .dout(n17127));
  jor  g17029(.dina(n17090), .dinb(n17127), .dout(n17128));
  jor  g17030(.dina(n17091), .dinb(n16961), .dout(n17129));
  jand g17031(.dina(n17129), .dinb(n17128), .dout(n17130));
  jor  g17032(.dina(n17079), .dinb(n17071), .dout(n17131));
  jor  g17033(.dina(n17081), .dinb(n16964), .dout(n17132));
  jand g17034(.dina(n17132), .dinb(n17131), .dout(n17133));
  jnot g17035(.din(n17060), .dout(n17134));
  jor  g17036(.dina(n17068), .dinb(n17134), .dout(n17135));
  jor  g17037(.dina(n17069), .dinb(n16968), .dout(n17136));
  jand g17038(.dina(n17136), .dinb(n17135), .dout(n17137));
  jor  g17039(.dina(n17058), .dinb(n17050), .dout(n17138));
  jnot g17040(.din(n17138), .dout(n17139));
  jand g17041(.dina(n17059), .dinb(n16972), .dout(n17140));
  jor  g17042(.dina(n17140), .dinb(n17139), .dout(n17141));
  jor  g17043(.dina(n17047), .dinb(n17039), .dout(n17142));
  jand g17044(.dina(n17048), .dinb(n16977), .dout(n17143));
  jnot g17045(.din(n17143), .dout(n17144));
  jand g17046(.dina(n17144), .dinb(n17142), .dout(n17145));
  jnot g17047(.din(n17145), .dout(n17146));
  jor  g17048(.dina(n17036), .dinb(n17028), .dout(n17147));
  jand g17049(.dina(n17037), .dinb(n16982), .dout(n17148));
  jnot g17050(.din(n17148), .dout(n17149));
  jand g17051(.dina(n17149), .dinb(n17147), .dout(n17150));
  jnot g17052(.din(n17150), .dout(n17151));
  jor  g17053(.dina(n17025), .dinb(n17017), .dout(n17152));
  jand g17054(.dina(n17026), .dinb(n16987), .dout(n17153));
  jnot g17055(.din(n17153), .dout(n17154));
  jand g17056(.dina(n17154), .dinb(n17152), .dout(n17155));
  jnot g17057(.din(n17155), .dout(n17156));
  jand g17058(.dina(n17014), .dinb(n17007), .dout(n17157));
  jand g17059(.dina(n17015), .dinb(n16990), .dout(n17158));
  jor  g17060(.dina(n17158), .dinb(n17157), .dout(n17159));
  jand g17061(.dina(n1968), .dinb(n499), .dout(n17160));
  jand g17062(.dina(n17160), .dinb(n1312), .dout(n17161));
  jand g17063(.dina(n17161), .dinb(n5298), .dout(n17162));
  jand g17064(.dina(n676), .dinb(n501), .dout(n17163));
  jand g17065(.dina(n17163), .dinb(n17162), .dout(n17164));
  jand g17066(.dina(n14327), .dinb(n2100), .dout(n17165));
  jand g17067(.dina(n700), .dinb(n991), .dout(n17166));
  jand g17068(.dina(n1721), .dinb(n2148), .dout(n17167));
  jand g17069(.dina(n17167), .dinb(n17166), .dout(n17168));
  jand g17070(.dina(n17168), .dinb(n17165), .dout(n17169));
  jand g17071(.dina(n10699), .dinb(n108), .dout(n17170));
  jand g17072(.dina(n1495), .dinb(n472), .dout(n17171));
  jand g17073(.dina(n1867), .dinb(n921), .dout(n17172));
  jand g17074(.dina(n17172), .dinb(n17171), .dout(n17173));
  jand g17075(.dina(n17173), .dinb(n17170), .dout(n17174));
  jand g17076(.dina(n1753), .dinb(n1732), .dout(n17175));
  jand g17077(.dina(n17175), .dinb(n13171), .dout(n17176));
  jand g17078(.dina(n17176), .dinb(n17174), .dout(n17177));
  jand g17079(.dina(n17177), .dinb(n17169), .dout(n17178));
  jand g17080(.dina(n1915), .dinb(n1837), .dout(n17179));
  jand g17081(.dina(n17179), .dinb(n431), .dout(n17180));
  jand g17082(.dina(n17180), .dinb(n17178), .dout(n17181));
  jand g17083(.dina(n17181), .dinb(n4649), .dout(n17182));
  jand g17084(.dina(n17182), .dinb(n11381), .dout(n17183));
  jand g17085(.dina(n17183), .dinb(n17164), .dout(n17184));
  jnot g17086(.din(n17184), .dout(n17185));
  jand g17087(.dina(n9886), .dinb(n5076), .dout(n17186));
  jand g17088(.dina(n9655), .dinb(n5084), .dout(n17187));
  jand g17089(.dina(n9250), .dinb(n6050), .dout(n17188));
  jand g17090(.dina(n9656), .dinb(n5082), .dout(n17189));
  jor  g17091(.dina(n17189), .dinb(n17188), .dout(n17190));
  jor  g17092(.dina(n17190), .dinb(n17187), .dout(n17191));
  jor  g17093(.dina(n17191), .dinb(n17186), .dout(n17192));
  jxor g17094(.dina(n17192), .dinb(n17185), .dout(n17193));
  jxor g17095(.dina(n17193), .dinb(n17159), .dout(n17194));
  jnot g17096(.din(n17194), .dout(n17195));
  jand g17097(.dina(n10862), .dinb(n2936), .dout(n17196));
  jand g17098(.dina(n10647), .dinb(n2943), .dout(n17197));
  jand g17099(.dina(n10305), .dinb(n2940), .dout(n17198));
  jand g17100(.dina(n9872), .dinb(n3684), .dout(n17199));
  jor  g17101(.dina(n17199), .dinb(n17198), .dout(n17200));
  jor  g17102(.dina(n17200), .dinb(n17197), .dout(n17201));
  jor  g17103(.dina(n17201), .dinb(n17196), .dout(n17202));
  jxor g17104(.dina(n17202), .dinb(n93), .dout(n17203));
  jxor g17105(.dina(n17203), .dinb(n17195), .dout(n17204));
  jxor g17106(.dina(n17204), .dinb(n17156), .dout(n17205));
  jnot g17107(.din(n17205), .dout(n17206));
  jand g17108(.dina(n11308), .dinb(n71), .dout(n17207));
  jand g17109(.dina(n10836), .dinb(n731), .dout(n17208));
  jand g17110(.dina(n11306), .dinb(n796), .dout(n17209));
  jor  g17111(.dina(n17209), .dinb(n17208), .dout(n17210));
  jand g17112(.dina(n10640), .dinb(n1806), .dout(n17211));
  jor  g17113(.dina(n17211), .dinb(n17210), .dout(n17212));
  jor  g17114(.dina(n17212), .dinb(n17207), .dout(n17213));
  jxor g17115(.dina(n17213), .dinb(n77), .dout(n17214));
  jxor g17116(.dina(n17214), .dinb(n17206), .dout(n17215));
  jxor g17117(.dina(n17215), .dinb(n17151), .dout(n17216));
  jnot g17118(.din(n17216), .dout(n17217));
  jand g17119(.dina(n11800), .dinb(n806), .dout(n17218));
  jand g17120(.dina(n11646), .dinb(n1612), .dout(n17219));
  jand g17121(.dina(n11798), .dinb(n1620), .dout(n17220));
  jor  g17122(.dina(n17220), .dinb(n17219), .dout(n17221));
  jand g17123(.dina(n11647), .dinb(n1644), .dout(n17222));
  jor  g17124(.dina(n17222), .dinb(n17221), .dout(n17223));
  jor  g17125(.dina(n17223), .dinb(n17218), .dout(n17224));
  jxor g17126(.dina(n17224), .dinb(n65), .dout(n17225));
  jxor g17127(.dina(n17225), .dinb(n17217), .dout(n17226));
  jxor g17128(.dina(n17226), .dinb(n17146), .dout(n17227));
  jnot g17129(.din(n17227), .dout(n17228));
  jand g17130(.dina(n12684), .dinb(n1819), .dout(n17229));
  jand g17131(.dina(n12547), .dinb(n2180), .dout(n17230));
  jand g17132(.dina(n12536), .dinb(n2243), .dout(n17231));
  jor  g17133(.dina(n17231), .dinb(n17230), .dout(n17232));
  jand g17134(.dina(n12282), .dinb(n2185), .dout(n17233));
  jor  g17135(.dina(n17233), .dinb(n17232), .dout(n17234));
  jor  g17136(.dina(n17234), .dinb(n17229), .dout(n17235));
  jxor g17137(.dina(n17235), .dinb(n2196), .dout(n17236));
  jxor g17138(.dina(n17236), .dinb(n17228), .dout(n17237));
  jxor g17139(.dina(n17237), .dinb(n17141), .dout(n17238));
  jand g17140(.dina(n13639), .dinb(n2743), .dout(n17239));
  jand g17141(.dina(n13478), .dinb(n2752), .dout(n17240));
  jand g17142(.dina(n13248), .dinb(n2748), .dout(n17241));
  jand g17143(.dina(n12669), .dinb(n2757), .dout(n17242));
  jor  g17144(.dina(n17242), .dinb(n17241), .dout(n17243));
  jor  g17145(.dina(n17243), .dinb(n17240), .dout(n17244));
  jor  g17146(.dina(n17244), .dinb(n17239), .dout(n17245));
  jxor g17147(.dina(n17245), .dinb(\a[17] ), .dout(n17246));
  jxor g17148(.dina(n17246), .dinb(n17238), .dout(n17247));
  jxor g17149(.dina(n17247), .dinb(n17137), .dout(n17248));
  jand g17150(.dina(n14251), .dinb(n3423), .dout(n17249));
  jand g17151(.dina(n13614), .dinb(n3428), .dout(n17250));
  jand g17152(.dina(n14249), .dinb(n3569), .dout(n17251));
  jor  g17153(.dina(n17251), .dinb(n17250), .dout(n17252));
  jand g17154(.dina(n13469), .dinb(n3210), .dout(n17253));
  jor  g17155(.dina(n17253), .dinb(n17252), .dout(n17254));
  jor  g17156(.dina(n17254), .dinb(n17249), .dout(n17255));
  jxor g17157(.dina(n17255), .dinb(n3473), .dout(n17256));
  jxor g17158(.dina(n17256), .dinb(n17248), .dout(n17257));
  jxor g17159(.dina(n17257), .dinb(n17133), .dout(n17258));
  jand g17160(.dina(n14551), .dinb(n4022), .dout(n17259));
  jand g17161(.dina(n14549), .dinb(n4220), .dout(n17260));
  jand g17162(.dina(n14447), .dinb(n4027), .dout(n17261));
  jand g17163(.dina(n14448), .dinb(n3870), .dout(n17262));
  jor  g17164(.dina(n17262), .dinb(n17261), .dout(n17263));
  jor  g17165(.dina(n17263), .dinb(n17260), .dout(n17264));
  jor  g17166(.dina(n17264), .dinb(n17259), .dout(n17265));
  jxor g17167(.dina(n17265), .dinb(n4050), .dout(n17266));
  jxor g17168(.dina(n17266), .dinb(n17258), .dout(n17267));
  jxor g17169(.dina(n17267), .dinb(n17130), .dout(n17268));
  jand g17170(.dina(n15831), .dinb(n4691), .dout(n17269));
  jand g17171(.dina(n15567), .dinb(n4696), .dout(n17270));
  jand g17172(.dina(n15829), .dinb(n4941), .dout(n17271));
  jor  g17173(.dina(n17271), .dinb(n17270), .dout(n17272));
  jand g17174(.dina(n15315), .dinb(n4701), .dout(n17273));
  jor  g17175(.dina(n17273), .dinb(n17272), .dout(n17274));
  jor  g17176(.dina(n17274), .dinb(n17269), .dout(n17275));
  jxor g17177(.dina(n17275), .dinb(n4713), .dout(n17276));
  jxor g17178(.dina(n17276), .dinb(n17268), .dout(n17277));
  jxor g17179(.dina(n17277), .dinb(n17126), .dout(n17278));
  jand g17180(.dina(n16594), .dinb(n5280), .dout(n17279));
  jand g17181(.dina(n16343), .dinb(n5531), .dout(n17280));
  jand g17182(.dina(n16592), .dinb(n5814), .dout(n17281));
  jor  g17183(.dina(n17281), .dinb(n17280), .dout(n17282));
  jand g17184(.dina(n16082), .dinb(n5536), .dout(n17283));
  jor  g17185(.dina(n17283), .dinb(n17282), .dout(n17284));
  jor  g17186(.dina(n17284), .dinb(n17279), .dout(n17285));
  jxor g17187(.dina(n17285), .dinb(n5277), .dout(n17286));
  jxor g17188(.dina(n17286), .dinb(n17278), .dout(n17287));
  jnot g17189(.din(n16928), .dout(n17288));
  jnot g17190(.din(n16592), .dout(n17289));
  jnot g17191(.din(n16922), .dout(n17291));
  jnot g17192(.din(n16929), .dout(n17292));
  jor  g17193(.dina(n17292), .dinb(n17291), .dout(n17293));
  jand g17194(.dina(n17293), .dinb(n17289), .dout(n17294));
  jor  g17195(.dina(n17294), .dinb(n16927), .dout(n17295));
  jand g17196(.dina(n17295), .dinb(n17288), .dout(n17296));
  jor  g17197(.dina(n17296), .dinb(n6496), .dout(n17297));
  jand g17198(.dina(n16342), .dinb(n16328), .dout(n17298));
  jor  g17199(.dina(n17298), .dinb(n16339), .dout(n17299));
  jnot g17200(.din(n16591), .dout(n17300));
  jand g17201(.dina(n17300), .dinb(n17299), .dout(n17301));
  jor  g17202(.dina(n6499), .dinb(n6495), .dout(n17303));
  jand g17203(.dina(n17303), .dinb(n6501), .dout(n17304));
  jor  g17204(.dina(n17304), .dinb(n17301), .dout(n17305));
  jand g17205(.dina(n17305), .dinb(n17297), .dout(n17306));
  jxor g17206(.dina(n17306), .dinb(\a[2] ), .dout(n17307));
  jxor g17207(.dina(n17307), .dinb(n17287), .dout(n17308));
  jxor g17208(.dina(n17308), .dinb(n17122), .dout(n17309));
  jxor g17209(.dina(n17120), .dinb(n17119), .dout(n17310));
  jnot g17210(.din(n17310), .dout(n17311));
  jxor g17211(.dina(n17294), .dinb(n16927), .dout(n17312));
  jand g17212(.dina(n17312), .dinb(n6495), .dout(n17313));
  jand g17213(.dina(n16928), .dinb(n6506), .dout(n17314));
  jand g17214(.dina(n16592), .dinb(n6500), .dout(n17315));
  jand g17215(.dina(n16924), .dinb(n6503), .dout(n17316));
  jor  g17216(.dina(n17316), .dinb(n17315), .dout(n17317));
  jor  g17217(.dina(n17317), .dinb(n17314), .dout(n17318));
  jor  g17218(.dina(n17318), .dinb(n17313), .dout(n17319));
  jxor g17219(.dina(n17319), .dinb(n6219), .dout(n17320));
  jor  g17220(.dina(n17320), .dinb(n17311), .dout(n17321));
  jnot g17221(.din(n16919), .dout(n17322));
  jor  g17222(.dina(n16938), .dinb(n17322), .dout(n17323));
  jor  g17223(.dina(n16939), .dinb(n16719), .dout(n17324));
  jand g17224(.dina(n17324), .dinb(n17323), .dout(n17325));
  jxor g17225(.dina(n17320), .dinb(n17310), .dout(n17326));
  jor  g17226(.dina(n17326), .dinb(n17325), .dout(n17327));
  jand g17227(.dina(n17327), .dinb(n17321), .dout(n17328));
  jxor g17228(.dina(n17328), .dinb(n17309), .dout(n17329));
  jxor g17229(.dina(n17326), .dinb(n17325), .dout(n17330));
  jand g17230(.dina(n17330), .dinb(n17329), .dout(n17331));
  jand g17231(.dina(n17330), .dinb(n16940), .dout(n17332));
  jand g17232(.dina(n16940), .dinb(n16604), .dout(n17333));
  jand g17233(.dina(n16941), .dinb(n16715), .dout(n17334));
  jor  g17234(.dina(n17334), .dinb(n17333), .dout(n17335));
  jxor g17235(.dina(n17330), .dinb(n16940), .dout(n17336));
  jand g17236(.dina(n17336), .dinb(n17335), .dout(n17337));
  jor  g17237(.dina(n17337), .dinb(n17332), .dout(n17338));
  jxor g17238(.dina(n17330), .dinb(n17329), .dout(n17339));
  jand g17239(.dina(n17339), .dinb(n17338), .dout(n17340));
  jor  g17240(.dina(n17340), .dinb(n17331), .dout(n17341));
  jnot g17241(.din(n17278), .dout(n17342));
  jor  g17242(.dina(n17286), .dinb(n17342), .dout(n17343));
  jor  g17243(.dina(n17307), .dinb(n17287), .dout(n17344));
  jand g17244(.dina(n17344), .dinb(n17343), .dout(n17345));
  jor  g17245(.dina(n17276), .dinb(n17268), .dout(n17346));
  jand g17246(.dina(n17277), .dinb(n17126), .dout(n17347));
  jnot g17247(.din(n17347), .dout(n17348));
  jand g17248(.dina(n17348), .dinb(n17346), .dout(n17349));
  jor  g17249(.dina(n17266), .dinb(n17258), .dout(n17350));
  jnot g17250(.din(n17267), .dout(n17351));
  jor  g17251(.dina(n17351), .dinb(n17130), .dout(n17352));
  jand g17252(.dina(n17352), .dinb(n17350), .dout(n17353));
  jor  g17253(.dina(n17256), .dinb(n17248), .dout(n17354));
  jnot g17254(.din(n17257), .dout(n17355));
  jor  g17255(.dina(n17355), .dinb(n17133), .dout(n17356));
  jand g17256(.dina(n17356), .dinb(n17354), .dout(n17357));
  jand g17257(.dina(n17246), .dinb(n17238), .dout(n17358));
  jnot g17258(.din(n17358), .dout(n17359));
  jnot g17259(.din(n17247), .dout(n17360));
  jor  g17260(.dina(n17360), .dinb(n17137), .dout(n17361));
  jand g17261(.dina(n17361), .dinb(n17359), .dout(n17362));
  jor  g17262(.dina(n17236), .dinb(n17228), .dout(n17363));
  jand g17263(.dina(n17237), .dinb(n17141), .dout(n17364));
  jnot g17264(.din(n17364), .dout(n17365));
  jand g17265(.dina(n17365), .dinb(n17363), .dout(n17366));
  jor  g17266(.dina(n17225), .dinb(n17217), .dout(n17367));
  jand g17267(.dina(n17226), .dinb(n17146), .dout(n17368));
  jnot g17268(.din(n17368), .dout(n17369));
  jand g17269(.dina(n17369), .dinb(n17367), .dout(n17370));
  jor  g17270(.dina(n17214), .dinb(n17206), .dout(n17371));
  jand g17271(.dina(n17215), .dinb(n17151), .dout(n17372));
  jnot g17272(.din(n17372), .dout(n17373));
  jand g17273(.dina(n17373), .dinb(n17371), .dout(n17374));
  jor  g17274(.dina(n17203), .dinb(n17195), .dout(n17375));
  jand g17275(.dina(n17204), .dinb(n17156), .dout(n17376));
  jnot g17276(.din(n17376), .dout(n17377));
  jand g17277(.dina(n17377), .dinb(n17375), .dout(n17378));
  jand g17278(.dina(n17192), .dinb(n17185), .dout(n17379));
  jand g17279(.dina(n17193), .dinb(n17159), .dout(n17380));
  jor  g17280(.dina(n17380), .dinb(n17379), .dout(n17381));
  jand g17281(.dina(n9874), .dinb(n5076), .dout(n17382));
  jand g17282(.dina(n9872), .dinb(n5084), .dout(n17383));
  jand g17283(.dina(n9655), .dinb(n5082), .dout(n17384));
  jand g17284(.dina(n9656), .dinb(n6050), .dout(n17385));
  jor  g17285(.dina(n17385), .dinb(n17384), .dout(n17386));
  jor  g17286(.dina(n17386), .dinb(n17383), .dout(n17387));
  jor  g17287(.dina(n17387), .dinb(n17382), .dout(n17388));
  jand g17288(.dina(n1437), .dinb(n92), .dout(n17389));
  jand g17289(.dina(n17389), .dinb(n6368), .dout(n17390));
  jand g17290(.dina(n17390), .dinb(n5171), .dout(n17391));
  jand g17291(.dina(n3264), .dinb(n453), .dout(n17392));
  jand g17292(.dina(n17392), .dinb(n17391), .dout(n17393));
  jand g17293(.dina(n1426), .dinb(n532), .dout(n17394));
  jand g17294(.dina(n17394), .dinb(n630), .dout(n17395));
  jand g17295(.dina(n3136), .dinb(n1040), .dout(n17396));
  jand g17296(.dina(n17396), .dinb(n17395), .dout(n17397));
  jand g17297(.dina(n1713), .dinb(n895), .dout(n17398));
  jand g17298(.dina(n17398), .dinb(n1832), .dout(n17399));
  jand g17299(.dina(n17399), .dinb(n674), .dout(n17400));
  jand g17300(.dina(n17400), .dinb(n17397), .dout(n17401));
  jand g17301(.dina(n17401), .dinb(n2547), .dout(n17402));
  jand g17302(.dina(n17402), .dinb(n17393), .dout(n17403));
  jand g17303(.dina(n1374), .dinb(n1326), .dout(n17404));
  jand g17304(.dina(n17404), .dinb(n2406), .dout(n17405));
  jand g17305(.dina(n15135), .dinb(n3194), .dout(n17406));
  jand g17306(.dina(n17406), .dinb(n17405), .dout(n17407));
  jand g17307(.dina(n17407), .dinb(n17403), .dout(n17408));
  jand g17308(.dina(n1583), .dinb(n1708), .dout(n17409));
  jand g17309(.dina(n17409), .dinb(n619), .dout(n17410));
  jand g17310(.dina(n1731), .dinb(n461), .dout(n17411));
  jand g17311(.dina(n988), .dinb(n1088), .dout(n17412));
  jand g17312(.dina(n17412), .dinb(n17411), .dout(n17413));
  jand g17313(.dina(n17413), .dinb(n17410), .dout(n17414));
  jand g17314(.dina(n15104), .dinb(n3338), .dout(n17415));
  jand g17315(.dina(n17415), .dinb(n17414), .dout(n17416));
  jand g17316(.dina(n17416), .dinb(n17408), .dout(n17417));
  jand g17317(.dina(n17417), .dinb(n16798), .dout(n17418));
  jor  g17318(.dina(n16924), .dinb(n6219), .dout(n17419));
  jor  g17319(.dina(n6499), .dinb(\a[2] ), .dout(n17420));
  jor  g17320(.dina(n17420), .dinb(n17301), .dout(n17421));
  jand g17321(.dina(n17421), .dinb(n17419), .dout(n17422));
  jxor g17322(.dina(n17422), .dinb(n17418), .dout(n17423));
  jxor g17323(.dina(n17423), .dinb(n17388), .dout(n17424));
  jxor g17324(.dina(n17424), .dinb(n17381), .dout(n17425));
  jnot g17325(.din(n10850), .dout(n17426));
  jor  g17326(.dina(n17426), .dinb(n4343), .dout(n17427));
  jnot g17327(.din(n10647), .dout(n17428));
  jor  g17328(.dina(n17428), .dinb(n4346), .dout(n17429));
  jor  g17329(.dina(n14955), .dinb(n4348), .dout(n17430));
  jand g17330(.dina(n17430), .dinb(n17429), .dout(n17431));
  jor  g17331(.dina(n14771), .dinb(n3683), .dout(n17432));
  jand g17332(.dina(n17432), .dinb(n17431), .dout(n17433));
  jand g17333(.dina(n17433), .dinb(n17427), .dout(n17434));
  jxor g17334(.dina(n17434), .dinb(\a[29] ), .dout(n17435));
  jnot g17335(.din(n17435), .dout(n17436));
  jxor g17336(.dina(n17436), .dinb(n17425), .dout(n17437));
  jxor g17337(.dina(n17437), .dinb(n17378), .dout(n17438));
  jand g17338(.dina(n11824), .dinb(n71), .dout(n17439));
  jand g17339(.dina(n11647), .dinb(n796), .dout(n17440));
  jand g17340(.dina(n11306), .dinb(n731), .dout(n17441));
  jand g17341(.dina(n10836), .dinb(n1806), .dout(n17442));
  jor  g17342(.dina(n17442), .dinb(n17441), .dout(n17443));
  jor  g17343(.dina(n17443), .dinb(n17440), .dout(n17444));
  jor  g17344(.dina(n17444), .dinb(n17439), .dout(n17445));
  jxor g17345(.dina(n17445), .dinb(n77), .dout(n17446));
  jxor g17346(.dina(n17446), .dinb(n17438), .dout(n17447));
  jxor g17347(.dina(n17447), .dinb(n17374), .dout(n17448));
  jand g17348(.dina(n12284), .dinb(n806), .dout(n17449));
  jand g17349(.dina(n11798), .dinb(n1612), .dout(n17450));
  jand g17350(.dina(n12282), .dinb(n1620), .dout(n17451));
  jor  g17351(.dina(n17451), .dinb(n17450), .dout(n17452));
  jand g17352(.dina(n11646), .dinb(n1644), .dout(n17453));
  jor  g17353(.dina(n17453), .dinb(n17452), .dout(n17454));
  jor  g17354(.dina(n17454), .dinb(n17449), .dout(n17455));
  jxor g17355(.dina(n17455), .dinb(n65), .dout(n17456));
  jxor g17356(.dina(n17456), .dinb(n17448), .dout(n17457));
  jxor g17357(.dina(n17457), .dinb(n17370), .dout(n17458));
  jand g17358(.dina(n12671), .dinb(n1819), .dout(n17459));
  jand g17359(.dina(n12669), .dinb(n2243), .dout(n17460));
  jand g17360(.dina(n12536), .dinb(n2180), .dout(n17461));
  jand g17361(.dina(n12547), .dinb(n2185), .dout(n17462));
  jor  g17362(.dina(n17462), .dinb(n17461), .dout(n17463));
  jor  g17363(.dina(n17463), .dinb(n17460), .dout(n17464));
  jor  g17364(.dina(n17464), .dinb(n17459), .dout(n17465));
  jxor g17365(.dina(n17465), .dinb(n2196), .dout(n17466));
  jxor g17366(.dina(n17466), .dinb(n17458), .dout(n17467));
  jxor g17367(.dina(n17467), .dinb(n17366), .dout(n17468));
  jnot g17368(.din(n13627), .dout(n17469));
  jor  g17369(.dina(n17469), .dinb(n2744), .dout(n17470));
  jor  g17370(.dina(n14988), .dinb(n2753), .dout(n17471));
  jor  g17371(.dina(n14990), .dinb(n2749), .dout(n17472));
  jnot g17372(.din(n13248), .dout(n17473));
  jor  g17373(.dina(n17473), .dinb(n2758), .dout(n17474));
  jand g17374(.dina(n17474), .dinb(n17472), .dout(n17475));
  jand g17375(.dina(n17475), .dinb(n17471), .dout(n17476));
  jand g17376(.dina(n17476), .dinb(n17470), .dout(n17477));
  jxor g17377(.dina(n17477), .dinb(\a[17] ), .dout(n17478));
  jxor g17378(.dina(n17478), .dinb(n17468), .dout(n17479));
  jxor g17379(.dina(n17479), .dinb(n17362), .dout(n17480));
  jor  g17380(.dina(n14580), .dinb(n3424), .dout(n17481));
  jor  g17381(.dina(n14567), .dinb(n3426), .dout(n17482));
  jor  g17382(.dina(n14569), .dinb(n3429), .dout(n17483));
  jor  g17383(.dina(n14584), .dinb(n3211), .dout(n17484));
  jand g17384(.dina(n17484), .dinb(n17483), .dout(n17485));
  jand g17385(.dina(n17485), .dinb(n17482), .dout(n17486));
  jand g17386(.dina(n17486), .dinb(n17481), .dout(n17487));
  jxor g17387(.dina(n17487), .dinb(\a[14] ), .dout(n17488));
  jxor g17388(.dina(n17488), .dinb(n17480), .dout(n17489));
  jxor g17389(.dina(n17489), .dinb(n17357), .dout(n17490));
  jnot g17390(.din(n15317), .dout(n17491));
  jor  g17391(.dina(n17491), .dinb(n4023), .dout(n17492));
  jnot g17392(.din(n14549), .dout(n17493));
  jor  g17393(.dina(n17493), .dinb(n4028), .dout(n17494));
  jnot g17394(.din(n15315), .dout(n17495));
  jor  g17395(.dina(n17495), .dinb(n4025), .dout(n17496));
  jand g17396(.dina(n17496), .dinb(n17494), .dout(n17497));
  jor  g17397(.dina(n14565), .dinb(n3871), .dout(n17498));
  jand g17398(.dina(n17498), .dinb(n17497), .dout(n17499));
  jand g17399(.dina(n17499), .dinb(n17492), .dout(n17500));
  jxor g17400(.dina(n17500), .dinb(\a[11] ), .dout(n17501));
  jxor g17401(.dina(n17501), .dinb(n17490), .dout(n17502));
  jxor g17402(.dina(n17502), .dinb(n17353), .dout(n17503));
  jnot g17403(.din(n16084), .dout(n17504));
  jor  g17404(.dina(n17504), .dinb(n4692), .dout(n17505));
  jnot g17405(.din(n15829), .dout(n17506));
  jor  g17406(.dina(n17506), .dinb(n4697), .dout(n17507));
  jnot g17407(.din(n16082), .dout(n17508));
  jor  g17408(.dina(n17508), .dinb(n4705), .dout(n17509));
  jand g17409(.dina(n17509), .dinb(n17507), .dout(n17510));
  jnot g17410(.din(n15567), .dout(n17511));
  jor  g17411(.dina(n17511), .dinb(n4702), .dout(n17512));
  jand g17412(.dina(n17512), .dinb(n17510), .dout(n17513));
  jand g17413(.dina(n17513), .dinb(n17505), .dout(n17514));
  jxor g17414(.dina(n17514), .dinb(\a[8] ), .dout(n17515));
  jxor g17415(.dina(n17515), .dinb(n17503), .dout(n17516));
  jxor g17416(.dina(n17516), .dinb(n17349), .dout(n17517));
  jnot g17417(.din(n16930), .dout(n17518));
  jor  g17418(.dina(n17518), .dinb(n5281), .dout(n17519));
  jor  g17419(.dina(n17289), .dinb(n5532), .dout(n17520));
  jor  g17420(.dina(n17288), .dinb(n5539), .dout(n17521));
  jand g17421(.dina(n17521), .dinb(n17520), .dout(n17522));
  jnot g17422(.din(n16343), .dout(n17523));
  jor  g17423(.dina(n17523), .dinb(n5537), .dout(n17524));
  jand g17424(.dina(n17524), .dinb(n17522), .dout(n17525));
  jand g17425(.dina(n17525), .dinb(n17519), .dout(n17526));
  jxor g17426(.dina(n17526), .dinb(\a[5] ), .dout(n17527));
  jxor g17427(.dina(n17527), .dinb(n17517), .dout(n17528));
  jxor g17428(.dina(n17528), .dinb(n17345), .dout(n17529));
  jnot g17429(.din(n17122), .dout(n17530));
  jand g17430(.dina(n17308), .dinb(n17530), .dout(n17531));
  jnot g17431(.din(n17531), .dout(n17532));
  jor  g17432(.dina(n17328), .dinb(n17309), .dout(n17533));
  jand g17433(.dina(n17533), .dinb(n17532), .dout(n17534));
  jxor g17434(.dina(n17534), .dinb(n17529), .dout(n17535));
  jxor g17435(.dina(n17535), .dinb(n17329), .dout(n17536));
  jxor g17436(.dina(n17536), .dinb(n17341), .dout(n17537));
  jand g17437(.dina(n17537), .dinb(n1819), .dout(n17538));
  jand g17438(.dina(n17535), .dinb(n2243), .dout(n17539));
  jand g17439(.dina(n17329), .dinb(n2180), .dout(n17540));
  jand g17440(.dina(n17330), .dinb(n2185), .dout(n17541));
  jor  g17441(.dina(n17541), .dinb(n17540), .dout(n17542));
  jor  g17442(.dina(n17542), .dinb(n17539), .dout(n17543));
  jor  g17443(.dina(n17543), .dinb(n17538), .dout(n17544));
  jxor g17444(.dina(n17544), .dinb(n2196), .dout(n17545));
  jor  g17445(.dina(n17545), .dinb(n16953), .dout(n17546));
  jxor g17446(.dina(n16684), .dinb(n16683), .dout(n17547));
  jnot g17447(.din(n17547), .dout(n17548));
  jxor g17448(.dina(n17339), .dinb(n17338), .dout(n17549));
  jand g17449(.dina(n17549), .dinb(n1819), .dout(n17550));
  jand g17450(.dina(n17329), .dinb(n2243), .dout(n17551));
  jand g17451(.dina(n17330), .dinb(n2180), .dout(n17552));
  jand g17452(.dina(n16940), .dinb(n2185), .dout(n17553));
  jor  g17453(.dina(n17553), .dinb(n17552), .dout(n17554));
  jor  g17454(.dina(n17554), .dinb(n17551), .dout(n17555));
  jor  g17455(.dina(n17555), .dinb(n17550), .dout(n17556));
  jxor g17456(.dina(n17556), .dinb(n2196), .dout(n17557));
  jor  g17457(.dina(n17557), .dinb(n17548), .dout(n17558));
  jxor g17458(.dina(n16681), .dinb(n16680), .dout(n17559));
  jnot g17459(.din(n17559), .dout(n17560));
  jxor g17460(.dina(n17336), .dinb(n17335), .dout(n17561));
  jand g17461(.dina(n17561), .dinb(n1819), .dout(n17562));
  jand g17462(.dina(n16940), .dinb(n2180), .dout(n17563));
  jand g17463(.dina(n17330), .dinb(n2243), .dout(n17564));
  jor  g17464(.dina(n17564), .dinb(n17563), .dout(n17565));
  jand g17465(.dina(n16604), .dinb(n2185), .dout(n17566));
  jor  g17466(.dina(n17566), .dinb(n17565), .dout(n17567));
  jor  g17467(.dina(n17567), .dinb(n17562), .dout(n17568));
  jxor g17468(.dina(n17568), .dinb(n2196), .dout(n17569));
  jor  g17469(.dina(n17569), .dinb(n17560), .dout(n17570));
  jxor g17470(.dina(n16676), .dinb(n16675), .dout(n17571));
  jnot g17471(.din(n17571), .dout(n17572));
  jand g17472(.dina(n16942), .dinb(n1819), .dout(n17573));
  jand g17473(.dina(n16604), .dinb(n2180), .dout(n17574));
  jand g17474(.dina(n16940), .dinb(n2243), .dout(n17575));
  jor  g17475(.dina(n17575), .dinb(n17574), .dout(n17576));
  jand g17476(.dina(n16355), .dinb(n2185), .dout(n17577));
  jor  g17477(.dina(n17577), .dinb(n17576), .dout(n17578));
  jor  g17478(.dina(n17578), .dinb(n17573), .dout(n17579));
  jxor g17479(.dina(n17579), .dinb(n2196), .dout(n17580));
  jor  g17480(.dina(n17580), .dinb(n17572), .dout(n17581));
  jxor g17481(.dina(n16672), .dinb(n16664), .dout(n17582));
  jnot g17482(.din(n17582), .dout(n17583));
  jand g17483(.dina(n16606), .dinb(n1819), .dout(n17584));
  jand g17484(.dina(n16355), .dinb(n2180), .dout(n17585));
  jand g17485(.dina(n16604), .dinb(n2243), .dout(n17586));
  jor  g17486(.dina(n17586), .dinb(n17585), .dout(n17587));
  jand g17487(.dina(n16360), .dinb(n2185), .dout(n17588));
  jor  g17488(.dina(n17588), .dinb(n17587), .dout(n17589));
  jor  g17489(.dina(n17589), .dinb(n17584), .dout(n17590));
  jxor g17490(.dina(n17590), .dinb(n2196), .dout(n17591));
  jor  g17491(.dina(n17591), .dinb(n17583), .dout(n17592));
  jand g17492(.dina(n16616), .dinb(n1819), .dout(n17593));
  jand g17493(.dina(n16355), .dinb(n2243), .dout(n17594));
  jand g17494(.dina(n16360), .dinb(n2180), .dout(n17595));
  jand g17495(.dina(n15841), .dinb(n2185), .dout(n17596));
  jor  g17496(.dina(n17596), .dinb(n17595), .dout(n17597));
  jor  g17497(.dina(n17597), .dinb(n17594), .dout(n17598));
  jor  g17498(.dina(n17598), .dinb(n17593), .dout(n17599));
  jxor g17499(.dina(n17599), .dinb(n2196), .dout(n17600));
  jnot g17500(.din(n17600), .dout(n17601));
  jor  g17501(.dina(n16651), .dinb(n65), .dout(n17602));
  jxor g17502(.dina(n17602), .dinb(n16659), .dout(n17603));
  jand g17503(.dina(n17603), .dinb(n17601), .dout(n17604));
  jand g17504(.dina(n16648), .dinb(\a[23] ), .dout(n17605));
  jxor g17505(.dina(n17605), .dinb(n16646), .dout(n17606));
  jnot g17506(.din(n17606), .dout(n17607));
  jand g17507(.dina(n16632), .dinb(n1819), .dout(n17608));
  jand g17508(.dina(n15841), .dinb(n2180), .dout(n17609));
  jand g17509(.dina(n16360), .dinb(n2243), .dout(n17610));
  jor  g17510(.dina(n17610), .dinb(n17609), .dout(n17611));
  jand g17511(.dina(n15579), .dinb(n2185), .dout(n17612));
  jor  g17512(.dina(n17612), .dinb(n17611), .dout(n17613));
  jor  g17513(.dina(n17613), .dinb(n17608), .dout(n17614));
  jxor g17514(.dina(n17614), .dinb(n2196), .dout(n17615));
  jor  g17515(.dina(n17615), .dinb(n17607), .dout(n17616));
  jand g17516(.dina(n15329), .dinb(n1819), .dout(n17617));
  jand g17517(.dina(n15020), .dinb(n2180), .dout(n17618));
  jand g17518(.dina(n15327), .dinb(n2243), .dout(n17619));
  jor  g17519(.dina(n17619), .dinb(n17618), .dout(n17620));
  jor  g17520(.dina(n17620), .dinb(n17617), .dout(n17621));
  jnot g17521(.din(n17621), .dout(n17622));
  jand g17522(.dina(n15020), .dinb(n1817), .dout(n17623));
  jnot g17523(.din(n17623), .dout(n17624));
  jand g17524(.dina(n17624), .dinb(\a[20] ), .dout(n17625));
  jand g17525(.dina(n17625), .dinb(n17622), .dout(n17626));
  jand g17526(.dina(n15580), .dinb(n1819), .dout(n17627));
  jand g17527(.dina(n15327), .dinb(n2180), .dout(n17628));
  jor  g17528(.dina(n17628), .dinb(n17627), .dout(n17629));
  jand g17529(.dina(n15579), .dinb(n2243), .dout(n17630));
  jand g17530(.dina(n15020), .dinb(n2185), .dout(n17631));
  jor  g17531(.dina(n17631), .dinb(n17630), .dout(n17632));
  jor  g17532(.dina(n17632), .dinb(n17629), .dout(n17633));
  jnot g17533(.din(n17633), .dout(n17634));
  jand g17534(.dina(n17634), .dinb(n17626), .dout(n17635));
  jand g17535(.dina(n17635), .dinb(n16648), .dout(n17636));
  jnot g17536(.din(n17636), .dout(n17637));
  jxor g17537(.dina(n17635), .dinb(n16648), .dout(n17638));
  jnot g17538(.din(n17638), .dout(n17639));
  jand g17539(.dina(n15848), .dinb(n1819), .dout(n17640));
  jand g17540(.dina(n15841), .dinb(n2243), .dout(n17641));
  jand g17541(.dina(n15579), .dinb(n2180), .dout(n17642));
  jand g17542(.dina(n15327), .dinb(n2185), .dout(n17643));
  jor  g17543(.dina(n17643), .dinb(n17642), .dout(n17644));
  jor  g17544(.dina(n17644), .dinb(n17641), .dout(n17645));
  jor  g17545(.dina(n17645), .dinb(n17640), .dout(n17646));
  jxor g17546(.dina(n17646), .dinb(n2196), .dout(n17647));
  jor  g17547(.dina(n17647), .dinb(n17639), .dout(n17648));
  jand g17548(.dina(n17648), .dinb(n17637), .dout(n17649));
  jnot g17549(.din(n17649), .dout(n17650));
  jxor g17550(.dina(n17615), .dinb(n17607), .dout(n17651));
  jand g17551(.dina(n17651), .dinb(n17650), .dout(n17652));
  jnot g17552(.din(n17652), .dout(n17653));
  jand g17553(.dina(n17653), .dinb(n17616), .dout(n17654));
  jnot g17554(.din(n17654), .dout(n17655));
  jxor g17555(.dina(n17603), .dinb(n17601), .dout(n17656));
  jand g17556(.dina(n17656), .dinb(n17655), .dout(n17657));
  jor  g17557(.dina(n17657), .dinb(n17604), .dout(n17658));
  jxor g17558(.dina(n17591), .dinb(n17583), .dout(n17659));
  jand g17559(.dina(n17659), .dinb(n17658), .dout(n17660));
  jnot g17560(.din(n17660), .dout(n17661));
  jand g17561(.dina(n17661), .dinb(n17592), .dout(n17662));
  jnot g17562(.din(n17662), .dout(n17663));
  jxor g17563(.dina(n17580), .dinb(n17572), .dout(n17664));
  jand g17564(.dina(n17664), .dinb(n17663), .dout(n17665));
  jnot g17565(.din(n17665), .dout(n17666));
  jand g17566(.dina(n17666), .dinb(n17581), .dout(n17667));
  jnot g17567(.din(n17667), .dout(n17668));
  jxor g17568(.dina(n17569), .dinb(n17560), .dout(n17669));
  jand g17569(.dina(n17669), .dinb(n17668), .dout(n17670));
  jnot g17570(.din(n17670), .dout(n17671));
  jand g17571(.dina(n17671), .dinb(n17570), .dout(n17672));
  jnot g17572(.din(n17672), .dout(n17673));
  jxor g17573(.dina(n17557), .dinb(n17548), .dout(n17674));
  jand g17574(.dina(n17674), .dinb(n17673), .dout(n17675));
  jnot g17575(.din(n17675), .dout(n17676));
  jand g17576(.dina(n17676), .dinb(n17558), .dout(n17677));
  jnot g17577(.din(n17677), .dout(n17678));
  jxor g17578(.dina(n17545), .dinb(n16953), .dout(n17679));
  jand g17579(.dina(n17679), .dinb(n17678), .dout(n17680));
  jnot g17580(.din(n17680), .dout(n17681));
  jand g17581(.dina(n17681), .dinb(n17546), .dout(n17682));
  jnot g17582(.din(n17682), .dout(n17683));
  jor  g17583(.dina(n16950), .dinb(n16712), .dout(n17684));
  jand g17584(.dina(n16951), .dinb(n16688), .dout(n17685));
  jnot g17585(.din(n17685), .dout(n17686));
  jand g17586(.dina(n17686), .dinb(n17684), .dout(n17687));
  jnot g17587(.din(n17687), .dout(n17688));
  jor  g17588(.dina(n16709), .dinb(n16701), .dout(n17689));
  jand g17589(.dina(n16710), .dinb(n16693), .dout(n17690));
  jnot g17590(.din(n17690), .dout(n17691));
  jand g17591(.dina(n17691), .dinb(n17689), .dout(n17692));
  jnot g17592(.din(n17692), .dout(n17693));
  jand g17593(.dina(n16616), .dinb(n71), .dout(n17694));
  jand g17594(.dina(n16360), .dinb(n731), .dout(n17695));
  jand g17595(.dina(n16355), .dinb(n796), .dout(n17696));
  jor  g17596(.dina(n17696), .dinb(n17695), .dout(n17697));
  jand g17597(.dina(n15841), .dinb(n1806), .dout(n17698));
  jor  g17598(.dina(n17698), .dinb(n17697), .dout(n17699));
  jor  g17599(.dina(n17699), .dinb(n17694), .dout(n17700));
  jxor g17600(.dina(n17700), .dinb(n77), .dout(n17701));
  jnot g17601(.din(n17701), .dout(n17702));
  jand g17602(.dina(n15580), .dinb(n2936), .dout(n17703));
  jand g17603(.dina(n15327), .dinb(n2940), .dout(n17704));
  jand g17604(.dina(n15579), .dinb(n2943), .dout(n17705));
  jor  g17605(.dina(n17705), .dinb(n17704), .dout(n17706));
  jand g17606(.dina(n15020), .dinb(n3684), .dout(n17707));
  jor  g17607(.dina(n17707), .dinb(n17706), .dout(n17708));
  jor  g17608(.dina(n17708), .dinb(n17703), .dout(n17709));
  jor  g17609(.dina(n15021), .dinb(n93), .dout(n17710));
  jor  g17610(.dina(n17710), .dinb(n16698), .dout(n17711));
  jand g17611(.dina(n17711), .dinb(\a[29] ), .dout(n17712));
  jxor g17612(.dina(n17712), .dinb(n17709), .dout(n17713));
  jxor g17613(.dina(n17713), .dinb(n17702), .dout(n17714));
  jxor g17614(.dina(n17714), .dinb(n17693), .dout(n17715));
  jnot g17615(.din(n17715), .dout(n17716));
  jand g17616(.dina(n17561), .dinb(n806), .dout(n17717));
  jand g17617(.dina(n17330), .dinb(n1620), .dout(n17718));
  jand g17618(.dina(n16940), .dinb(n1612), .dout(n17719));
  jand g17619(.dina(n16604), .dinb(n1644), .dout(n17720));
  jor  g17620(.dina(n17720), .dinb(n17719), .dout(n17721));
  jor  g17621(.dina(n17721), .dinb(n17718), .dout(n17722));
  jor  g17622(.dina(n17722), .dinb(n17717), .dout(n17723));
  jxor g17623(.dina(n17723), .dinb(n65), .dout(n17724));
  jxor g17624(.dina(n17724), .dinb(n17716), .dout(n17725));
  jxor g17625(.dina(n17725), .dinb(n17688), .dout(n17726));
  jnot g17626(.din(n17726), .dout(n17727));
  jand g17627(.dina(n17535), .dinb(n17329), .dout(n17728));
  jand g17628(.dina(n17536), .dinb(n17341), .dout(n17729));
  jor  g17629(.dina(n17729), .dinb(n17728), .dout(n17730));
  jnot g17630(.din(n17349), .dout(n17731));
  jand g17631(.dina(n17516), .dinb(n17731), .dout(n17732));
  jnot g17632(.din(n17732), .dout(n17733));
  jor  g17633(.dina(n17527), .dinb(n17517), .dout(n17734));
  jand g17634(.dina(n17734), .dinb(n17733), .dout(n17735));
  jnot g17635(.din(n17353), .dout(n17736));
  jand g17636(.dina(n17502), .dinb(n17736), .dout(n17737));
  jnot g17637(.din(n17737), .dout(n17738));
  jor  g17638(.dina(n17515), .dinb(n17503), .dout(n17739));
  jand g17639(.dina(n17739), .dinb(n17738), .dout(n17740));
  jnot g17640(.din(n17357), .dout(n17741));
  jand g17641(.dina(n17489), .dinb(n17741), .dout(n17742));
  jnot g17642(.din(n17742), .dout(n17743));
  jor  g17643(.dina(n17501), .dinb(n17490), .dout(n17744));
  jand g17644(.dina(n17744), .dinb(n17743), .dout(n17745));
  jnot g17645(.din(n17362), .dout(n17746));
  jand g17646(.dina(n17479), .dinb(n17746), .dout(n17747));
  jnot g17647(.din(n17747), .dout(n17748));
  jor  g17648(.dina(n17488), .dinb(n17480), .dout(n17749));
  jand g17649(.dina(n17749), .dinb(n17748), .dout(n17750));
  jnot g17650(.din(n17467), .dout(n17751));
  jor  g17651(.dina(n17751), .dinb(n17366), .dout(n17752));
  jor  g17652(.dina(n17478), .dinb(n17468), .dout(n17753));
  jand g17653(.dina(n17753), .dinb(n17752), .dout(n17754));
  jnot g17654(.din(n17457), .dout(n17755));
  jor  g17655(.dina(n17755), .dinb(n17370), .dout(n17756));
  jor  g17656(.dina(n17466), .dinb(n17458), .dout(n17757));
  jand g17657(.dina(n17757), .dinb(n17756), .dout(n17758));
  jnot g17658(.din(n17447), .dout(n17759));
  jor  g17659(.dina(n17759), .dinb(n17374), .dout(n17760));
  jor  g17660(.dina(n17456), .dinb(n17448), .dout(n17761));
  jand g17661(.dina(n17761), .dinb(n17760), .dout(n17762));
  jnot g17662(.din(n17437), .dout(n17763));
  jor  g17663(.dina(n17763), .dinb(n17378), .dout(n17764));
  jor  g17664(.dina(n17446), .dinb(n17438), .dout(n17765));
  jand g17665(.dina(n17765), .dinb(n17764), .dout(n17766));
  jand g17666(.dina(n17424), .dinb(n17381), .dout(n17767));
  jand g17667(.dina(n17436), .dinb(n17425), .dout(n17768));
  jor  g17668(.dina(n17768), .dinb(n17767), .dout(n17769));
  jand g17669(.dina(n10307), .dinb(n5076), .dout(n17770));
  jand g17670(.dina(n10305), .dinb(n5084), .dout(n17771));
  jand g17671(.dina(n9872), .dinb(n5082), .dout(n17772));
  jand g17672(.dina(n9655), .dinb(n6050), .dout(n17773));
  jor  g17673(.dina(n17773), .dinb(n17772), .dout(n17774));
  jor  g17674(.dina(n17774), .dinb(n17771), .dout(n17775));
  jor  g17675(.dina(n17775), .dinb(n17770), .dout(n17776));
  jnot g17676(.din(n17418), .dout(n17777));
  jand g17677(.dina(n17301), .dinb(\a[2] ), .dout(n17778));
  jnot g17678(.din(n17420), .dout(n17779));
  jand g17679(.dina(n17779), .dinb(n16924), .dout(n17780));
  jor  g17680(.dina(n17780), .dinb(n17778), .dout(n17781));
  jand g17681(.dina(n17781), .dinb(n17777), .dout(n17782));
  jand g17682(.dina(n17423), .dinb(n17388), .dout(n17783));
  jor  g17683(.dina(n17783), .dinb(n17782), .dout(n17784));
  jand g17684(.dina(n16563), .dinb(n4494), .dout(n17785));
  jand g17685(.dina(n6149), .dinb(n838), .dout(n17786));
  jand g17686(.dina(n4517), .dinb(n2154), .dout(n17787));
  jand g17687(.dina(n17787), .dinb(n1096), .dout(n17788));
  jand g17688(.dina(n17788), .dinb(n10527), .dout(n17789));
  jand g17689(.dina(n17789), .dinb(n17786), .dout(n17790));
  jand g17690(.dina(n632), .dinb(n3185), .dout(n17791));
  jand g17691(.dina(n3328), .dinb(n1846), .dout(n17792));
  jand g17692(.dina(n17792), .dinb(n3989), .dout(n17793));
  jand g17693(.dina(n17793), .dinb(n445), .dout(n17794));
  jand g17694(.dina(n17794), .dinb(n17791), .dout(n17795));
  jand g17695(.dina(n17795), .dinb(n17790), .dout(n17796));
  jand g17696(.dina(n4440), .dinb(n929), .dout(n17797));
  jand g17697(.dina(n17797), .dinb(n9734), .dout(n17798));
  jand g17698(.dina(n5518), .dinb(n827), .dout(n17799));
  jand g17699(.dina(n17799), .dinb(n5367), .dout(n17800));
  jand g17700(.dina(n17800), .dinb(n17798), .dout(n17801));
  jand g17701(.dina(n17801), .dinb(n1196), .dout(n17802));
  jand g17702(.dina(n1270), .dinb(n1226), .dout(n17803));
  jand g17703(.dina(n17803), .dinb(n1160), .dout(n17804));
  jand g17704(.dina(n17804), .dinb(n15104), .dout(n17805));
  jand g17705(.dina(n17805), .dinb(n14310), .dout(n17806));
  jand g17706(.dina(n3066), .dinb(n1913), .dout(n17807));
  jand g17707(.dina(n17807), .dinb(n17806), .dout(n17808));
  jand g17708(.dina(n17808), .dinb(n17802), .dout(n17809));
  jand g17709(.dina(n17809), .dinb(n17796), .dout(n17810));
  jand g17710(.dina(n1532), .dinb(n650), .dout(n17811));
  jand g17711(.dina(n17811), .dinb(n683), .dout(n17812));
  jand g17712(.dina(n17812), .dinb(n3827), .dout(n17813));
  jand g17713(.dina(n2509), .dinb(n2331), .dout(n17814));
  jand g17714(.dina(n17814), .dinb(n17813), .dout(n17815));
  jand g17715(.dina(n1579), .dinb(n542), .dout(n17816));
  jand g17716(.dina(n1903), .dinb(n1378), .dout(n17817));
  jand g17717(.dina(n17817), .dinb(n17816), .dout(n17818));
  jand g17718(.dina(n17818), .dinb(n17815), .dout(n17819));
  jand g17719(.dina(n908), .dinb(n1358), .dout(n17820));
  jand g17720(.dina(n17820), .dinb(n5258), .dout(n17821));
  jand g17721(.dina(n17821), .dinb(n17819), .dout(n17822));
  jand g17722(.dina(n873), .dinb(n893), .dout(n17823));
  jand g17723(.dina(n1306), .dinb(n843), .dout(n17824));
  jand g17724(.dina(n17824), .dinb(n17823), .dout(n17825));
  jand g17725(.dina(n11394), .dinb(n326), .dout(n17826));
  jand g17726(.dina(n17826), .dinb(n17825), .dout(n17827));
  jand g17727(.dina(n17827), .dinb(n17822), .dout(n17828));
  jand g17728(.dina(n17828), .dinb(n17810), .dout(n17829));
  jand g17729(.dina(n17829), .dinb(n17785), .dout(n17830));
  jxor g17730(.dina(n17830), .dinb(n17422), .dout(n17831));
  jxor g17731(.dina(n17831), .dinb(n17784), .dout(n17832));
  jxor g17732(.dina(n17832), .dinb(n17776), .dout(n17833));
  jxor g17733(.dina(n17833), .dinb(n17769), .dout(n17834));
  jand g17734(.dina(n10838), .dinb(n2936), .dout(n17835));
  jand g17735(.dina(n10640), .dinb(n2940), .dout(n17836));
  jand g17736(.dina(n10836), .dinb(n2943), .dout(n17837));
  jor  g17737(.dina(n17837), .dinb(n17836), .dout(n17838));
  jand g17738(.dina(n10647), .dinb(n3684), .dout(n17839));
  jor  g17739(.dina(n17839), .dinb(n17838), .dout(n17840));
  jor  g17740(.dina(n17840), .dinb(n17835), .dout(n17841));
  jxor g17741(.dina(n17841), .dinb(n93), .dout(n17842));
  jxor g17742(.dina(n17842), .dinb(n17834), .dout(n17843));
  jnot g17743(.din(n11812), .dout(n17844));
  jor  g17744(.dina(n17844), .dinb(n2303), .dout(n17845));
  jnot g17745(.din(n11646), .dout(n17846));
  jor  g17746(.dina(n17846), .dinb(n2309), .dout(n17847));
  jor  g17747(.dina(n14951), .dinb(n1805), .dout(n17848));
  jnot g17748(.din(n11647), .dout(n17849));
  jor  g17749(.dina(n17849), .dinb(n2306), .dout(n17850));
  jand g17750(.dina(n17850), .dinb(n17848), .dout(n17851));
  jand g17751(.dina(n17851), .dinb(n17847), .dout(n17852));
  jand g17752(.dina(n17852), .dinb(n17845), .dout(n17853));
  jxor g17753(.dina(n17853), .dinb(\a[26] ), .dout(n17854));
  jxor g17754(.dina(n17854), .dinb(n17843), .dout(n17855));
  jxor g17755(.dina(n17855), .dinb(n17766), .dout(n17856));
  jnot g17756(.din(n12696), .dout(n17857));
  jor  g17757(.dina(n17857), .dinb(n807), .dout(n17858));
  jnot g17758(.din(n12547), .dout(n17859));
  jor  g17759(.dina(n17859), .dinb(n1621), .dout(n17860));
  jnot g17760(.din(n12282), .dout(n17861));
  jor  g17761(.dina(n17861), .dinb(n1613), .dout(n17862));
  jnot g17762(.din(n11798), .dout(n17863));
  jor  g17763(.dina(n17863), .dinb(n1617), .dout(n17864));
  jand g17764(.dina(n17864), .dinb(n17862), .dout(n17865));
  jand g17765(.dina(n17865), .dinb(n17860), .dout(n17866));
  jand g17766(.dina(n17866), .dinb(n17858), .dout(n17867));
  jxor g17767(.dina(n17867), .dinb(\a[23] ), .dout(n17868));
  jxor g17768(.dina(n17868), .dinb(n17856), .dout(n17869));
  jxor g17769(.dina(n17869), .dinb(n17762), .dout(n17870));
  jnot g17770(.din(n13250), .dout(n17871));
  jor  g17771(.dina(n17871), .dinb(n1820), .dout(n17872));
  jor  g17772(.dina(n17473), .dinb(n2189), .dout(n17873));
  jnot g17773(.din(n12669), .dout(n17874));
  jor  g17774(.dina(n17874), .dinb(n2181), .dout(n17875));
  jnot g17775(.din(n12536), .dout(n17876));
  jor  g17776(.dina(n17876), .dinb(n2186), .dout(n17877));
  jand g17777(.dina(n17877), .dinb(n17875), .dout(n17878));
  jand g17778(.dina(n17878), .dinb(n17873), .dout(n17879));
  jand g17779(.dina(n17879), .dinb(n17872), .dout(n17880));
  jxor g17780(.dina(n17880), .dinb(\a[20] ), .dout(n17881));
  jxor g17781(.dina(n17881), .dinb(n17870), .dout(n17882));
  jxor g17782(.dina(n17882), .dinb(n17758), .dout(n17883));
  jor  g17783(.dina(n14985), .dinb(n2744), .dout(n17884));
  jor  g17784(.dina(n14584), .dinb(n2753), .dout(n17885));
  jor  g17785(.dina(n14988), .dinb(n2749), .dout(n17886));
  jor  g17786(.dina(n14990), .dinb(n2758), .dout(n17887));
  jand g17787(.dina(n17887), .dinb(n17886), .dout(n17888));
  jand g17788(.dina(n17888), .dinb(n17885), .dout(n17889));
  jand g17789(.dina(n17889), .dinb(n17884), .dout(n17890));
  jxor g17790(.dina(n17890), .dinb(\a[17] ), .dout(n17891));
  jxor g17791(.dina(n17891), .dinb(n17883), .dout(n17892));
  jxor g17792(.dina(n17892), .dinb(n17754), .dout(n17893));
  jor  g17793(.dina(n14563), .dinb(n3424), .dout(n17894));
  jor  g17794(.dina(n14565), .dinb(n3426), .dout(n17895));
  jor  g17795(.dina(n14567), .dinb(n3429), .dout(n17896));
  jor  g17796(.dina(n14569), .dinb(n3211), .dout(n17897));
  jand g17797(.dina(n17897), .dinb(n17896), .dout(n17898));
  jand g17798(.dina(n17898), .dinb(n17895), .dout(n17899));
  jand g17799(.dina(n17899), .dinb(n17894), .dout(n17900));
  jxor g17800(.dina(n17900), .dinb(\a[14] ), .dout(n17901));
  jxor g17801(.dina(n17901), .dinb(n17893), .dout(n17902));
  jxor g17802(.dina(n17902), .dinb(n17750), .dout(n17903));
  jnot g17803(.din(n15569), .dout(n17904));
  jor  g17804(.dina(n17904), .dinb(n4023), .dout(n17905));
  jor  g17805(.dina(n17511), .dinb(n4025), .dout(n17906));
  jor  g17806(.dina(n17495), .dinb(n4028), .dout(n17907));
  jor  g17807(.dina(n17493), .dinb(n3871), .dout(n17908));
  jand g17808(.dina(n17908), .dinb(n17907), .dout(n17909));
  jand g17809(.dina(n17909), .dinb(n17906), .dout(n17910));
  jand g17810(.dina(n17910), .dinb(n17905), .dout(n17911));
  jxor g17811(.dina(n17911), .dinb(\a[11] ), .dout(n17912));
  jxor g17812(.dina(n17912), .dinb(n17903), .dout(n17913));
  jxor g17813(.dina(n17913), .dinb(n17745), .dout(n17914));
  jnot g17814(.din(n16345), .dout(n17915));
  jor  g17815(.dina(n17915), .dinb(n4692), .dout(n17916));
  jor  g17816(.dina(n17508), .dinb(n4697), .dout(n17917));
  jor  g17817(.dina(n17523), .dinb(n4705), .dout(n17918));
  jand g17818(.dina(n17918), .dinb(n17917), .dout(n17919));
  jor  g17819(.dina(n17506), .dinb(n4702), .dout(n17920));
  jand g17820(.dina(n17920), .dinb(n17919), .dout(n17921));
  jand g17821(.dina(n17921), .dinb(n17916), .dout(n17922));
  jxor g17822(.dina(n17922), .dinb(\a[8] ), .dout(n17923));
  jxor g17823(.dina(n17923), .dinb(n17914), .dout(n17924));
  jxor g17824(.dina(n17924), .dinb(n17740), .dout(n17925));
  jnot g17825(.din(n17312), .dout(n17926));
  jor  g17826(.dina(n17926), .dinb(n5281), .dout(n17927));
  jor  g17827(.dina(n17288), .dinb(n5532), .dout(n17928));
  jor  g17828(.dina(n17289), .dinb(n5537), .dout(n17929));
  jor  g17829(.dina(n17301), .dinb(n5539), .dout(n17930));
  jand g17830(.dina(n17930), .dinb(n17929), .dout(n17931));
  jand g17831(.dina(n17931), .dinb(n17928), .dout(n17932));
  jand g17832(.dina(n17932), .dinb(n17927), .dout(n17933));
  jxor g17833(.dina(n17933), .dinb(\a[5] ), .dout(n17934));
  jxor g17834(.dina(n17934), .dinb(n17925), .dout(n17935));
  jxor g17835(.dina(n17935), .dinb(n17735), .dout(n17936));
  jxor g17836(.dina(n17516), .dinb(n17731), .dout(n17937));
  jxor g17837(.dina(n17527), .dinb(n17937), .dout(n17938));
  jor  g17838(.dina(n17938), .dinb(n17345), .dout(n17939));
  jor  g17839(.dina(n17534), .dinb(n17529), .dout(n17940));
  jand g17840(.dina(n17940), .dinb(n17939), .dout(n17941));
  jxor g17841(.dina(n17941), .dinb(n17936), .dout(n17942));
  jxor g17842(.dina(n17942), .dinb(n17535), .dout(n17943));
  jxor g17843(.dina(n17943), .dinb(n17730), .dout(n17944));
  jand g17844(.dina(n17944), .dinb(n1819), .dout(n17945));
  jand g17845(.dina(n17535), .dinb(n2180), .dout(n17946));
  jand g17846(.dina(n17942), .dinb(n2243), .dout(n17947));
  jor  g17847(.dina(n17947), .dinb(n17946), .dout(n17948));
  jand g17848(.dina(n17329), .dinb(n2185), .dout(n17949));
  jor  g17849(.dina(n17949), .dinb(n17948), .dout(n17950));
  jor  g17850(.dina(n17950), .dinb(n17945), .dout(n17951));
  jxor g17851(.dina(n17951), .dinb(n2196), .dout(n17952));
  jxor g17852(.dina(n17952), .dinb(n17727), .dout(n17953));
  jxor g17853(.dina(n17953), .dinb(n17683), .dout(n17954));
  jnot g17854(.din(n17954), .dout(n17955));
  jnot g17855(.din(n17740), .dout(n17956));
  jand g17856(.dina(n17924), .dinb(n17956), .dout(n17957));
  jnot g17857(.din(n17957), .dout(n17958));
  jor  g17858(.dina(n17934), .dinb(n17925), .dout(n17959));
  jand g17859(.dina(n17959), .dinb(n17958), .dout(n17960));
  jnot g17860(.din(n17745), .dout(n17961));
  jand g17861(.dina(n17913), .dinb(n17961), .dout(n17962));
  jnot g17862(.din(n17962), .dout(n17963));
  jor  g17863(.dina(n17923), .dinb(n17914), .dout(n17964));
  jand g17864(.dina(n17964), .dinb(n17963), .dout(n17965));
  jor  g17865(.dina(n5535), .dinb(n5280), .dout(n17966));
  jxor g17866(.dina(n18201), .dinb(n17965), .dout(n17973));
  jnot g17867(.din(n17750), .dout(n17974));
  jand g17868(.dina(n17902), .dinb(n17974), .dout(n17975));
  jnot g17869(.din(n17975), .dout(n17976));
  jor  g17870(.dina(n17912), .dinb(n17903), .dout(n17977));
  jand g17871(.dina(n17977), .dinb(n17976), .dout(n17978));
  jnot g17872(.din(n17754), .dout(n17979));
  jand g17873(.dina(n17892), .dinb(n17979), .dout(n17980));
  jnot g17874(.din(n17980), .dout(n17981));
  jor  g17875(.dina(n17901), .dinb(n17893), .dout(n17982));
  jand g17876(.dina(n17982), .dinb(n17981), .dout(n17983));
  jnot g17877(.din(n17882), .dout(n17984));
  jor  g17878(.dina(n17984), .dinb(n17758), .dout(n17985));
  jor  g17879(.dina(n17891), .dinb(n17883), .dout(n17986));
  jand g17880(.dina(n17986), .dinb(n17985), .dout(n17987));
  jnot g17881(.din(n17869), .dout(n17988));
  jor  g17882(.dina(n17988), .dinb(n17762), .dout(n17989));
  jor  g17883(.dina(n17881), .dinb(n17870), .dout(n17990));
  jand g17884(.dina(n17990), .dinb(n17989), .dout(n17991));
  jnot g17885(.din(n17855), .dout(n17992));
  jor  g17886(.dina(n17992), .dinb(n17766), .dout(n17993));
  jor  g17887(.dina(n17868), .dinb(n17856), .dout(n17994));
  jand g17888(.dina(n17994), .dinb(n17993), .dout(n17995));
  jnot g17889(.din(n17834), .dout(n17996));
  jor  g17890(.dina(n17842), .dinb(n17996), .dout(n17997));
  jor  g17891(.dina(n17854), .dinb(n17843), .dout(n17998));
  jand g17892(.dina(n17998), .dinb(n17997), .dout(n17999));
  jand g17893(.dina(n17832), .dinb(n17776), .dout(n18000));
  jand g17894(.dina(n17833), .dinb(n17769), .dout(n18001));
  jor  g17895(.dina(n18001), .dinb(n18000), .dout(n18002));
  jand g17896(.dina(n10862), .dinb(n5076), .dout(n18003));
  jand g17897(.dina(n10647), .dinb(n5084), .dout(n18004));
  jand g17898(.dina(n10305), .dinb(n5082), .dout(n18005));
  jand g17899(.dina(n9872), .dinb(n6050), .dout(n18006));
  jor  g17900(.dina(n18006), .dinb(n18005), .dout(n18007));
  jor  g17901(.dina(n18007), .dinb(n18004), .dout(n18008));
  jor  g17902(.dina(n18008), .dinb(n18003), .dout(n18009));
  jnot g17903(.din(n17830), .dout(n18010));
  jand g17904(.dina(n18010), .dinb(n17781), .dout(n18011));
  jand g17905(.dina(n17831), .dinb(n17784), .dout(n18012));
  jor  g17906(.dina(n18012), .dinb(n18011), .dout(n18013));
  jand g17907(.dina(n1515), .dinb(n685), .dout(n18014));
  jand g17908(.dina(n18014), .dinb(n1577), .dout(n18015));
  jand g17909(.dina(n3750), .dinb(n411), .dout(n18016));
  jand g17910(.dina(n18016), .dinb(n2713), .dout(n18017));
  jand g17911(.dina(n18017), .dinb(n3377), .dout(n18018));
  jand g17912(.dina(n18018), .dinb(n18015), .dout(n18019));
  jand g17913(.dina(n18019), .dinb(n9361), .dout(n18020));
  jand g17914(.dina(n510), .dinb(n555), .dout(n18021));
  jand g17915(.dina(n18021), .dinb(n619), .dout(n18022));
  jand g17916(.dina(n18022), .dinb(n2019), .dout(n18023));
  jand g17917(.dina(n18023), .dinb(n1323), .dout(n18024));
  jand g17918(.dina(n820), .dinb(n678), .dout(n18025));
  jand g17919(.dina(n18025), .dinb(n18024), .dout(n18026));
  jand g17920(.dina(n18026), .dinb(n6239), .dout(n18027));
  jand g17921(.dina(n18027), .dinb(n18020), .dout(n18028));
  jand g17922(.dina(n18028), .dinb(n13401), .dout(n18029));
  jxor g17923(.dina(n18029), .dinb(n17422), .dout(n18030));
  jxor g17924(.dina(n18030), .dinb(n18013), .dout(n18031));
  jxor g17925(.dina(n18031), .dinb(n18009), .dout(n18032));
  jxor g17926(.dina(n18032), .dinb(n18002), .dout(n18033));
  jand g17927(.dina(n11308), .dinb(n2936), .dout(n18034));
  jand g17928(.dina(n10836), .dinb(n2940), .dout(n18035));
  jand g17929(.dina(n11306), .dinb(n2943), .dout(n18036));
  jor  g17930(.dina(n18036), .dinb(n18035), .dout(n18037));
  jand g17931(.dina(n10640), .dinb(n3684), .dout(n18038));
  jor  g17932(.dina(n18038), .dinb(n18037), .dout(n18039));
  jor  g17933(.dina(n18039), .dinb(n18034), .dout(n18040));
  jxor g17934(.dina(n18040), .dinb(n93), .dout(n18041));
  jxor g17935(.dina(n18041), .dinb(n18033), .dout(n18042));
  jand g17936(.dina(n11800), .dinb(n71), .dout(n18043));
  jand g17937(.dina(n11646), .dinb(n731), .dout(n18044));
  jand g17938(.dina(n11798), .dinb(n796), .dout(n18045));
  jor  g17939(.dina(n18045), .dinb(n18044), .dout(n18046));
  jand g17940(.dina(n11647), .dinb(n1806), .dout(n18047));
  jor  g17941(.dina(n18047), .dinb(n18046), .dout(n18048));
  jor  g17942(.dina(n18048), .dinb(n18043), .dout(n18049));
  jxor g17943(.dina(n18049), .dinb(n77), .dout(n18050));
  jxor g17944(.dina(n18050), .dinb(n18042), .dout(n18051));
  jxor g17945(.dina(n18051), .dinb(n17999), .dout(n18052));
  jand g17946(.dina(n12684), .dinb(n806), .dout(n18053));
  jand g17947(.dina(n12547), .dinb(n1612), .dout(n18054));
  jand g17948(.dina(n12536), .dinb(n1620), .dout(n18055));
  jor  g17949(.dina(n18055), .dinb(n18054), .dout(n18056));
  jand g17950(.dina(n12282), .dinb(n1644), .dout(n18057));
  jor  g17951(.dina(n18057), .dinb(n18056), .dout(n18058));
  jor  g17952(.dina(n18058), .dinb(n18053), .dout(n18059));
  jxor g17953(.dina(n18059), .dinb(n65), .dout(n18060));
  jxor g17954(.dina(n18060), .dinb(n18052), .dout(n18061));
  jxor g17955(.dina(n18061), .dinb(n17995), .dout(n18062));
  jand g17956(.dina(n13639), .dinb(n1819), .dout(n18063));
  jand g17957(.dina(n13478), .dinb(n2243), .dout(n18064));
  jand g17958(.dina(n13248), .dinb(n2180), .dout(n18065));
  jand g17959(.dina(n12669), .dinb(n2185), .dout(n18066));
  jor  g17960(.dina(n18066), .dinb(n18065), .dout(n18067));
  jor  g17961(.dina(n18067), .dinb(n18064), .dout(n18068));
  jor  g17962(.dina(n18068), .dinb(n18063), .dout(n18069));
  jxor g17963(.dina(n18069), .dinb(n2196), .dout(n18070));
  jxor g17964(.dina(n18070), .dinb(n18062), .dout(n18071));
  jxor g17965(.dina(n18071), .dinb(n17991), .dout(n18072));
  jor  g17966(.dina(n15000), .dinb(n2744), .dout(n18073));
  jor  g17967(.dina(n14569), .dinb(n2753), .dout(n18074));
  jor  g17968(.dina(n14584), .dinb(n2749), .dout(n18075));
  jor  g17969(.dina(n14988), .dinb(n2758), .dout(n18076));
  jand g17970(.dina(n18076), .dinb(n18075), .dout(n18077));
  jand g17971(.dina(n18077), .dinb(n18074), .dout(n18078));
  jand g17972(.dina(n18078), .dinb(n18073), .dout(n18079));
  jxor g17973(.dina(n18079), .dinb(\a[17] ), .dout(n18080));
  jxor g17974(.dina(n18080), .dinb(n18072), .dout(n18081));
  jxor g17975(.dina(n18081), .dinb(n17987), .dout(n18082));
  jnot g17976(.din(n14551), .dout(n18083));
  jor  g17977(.dina(n18083), .dinb(n3424), .dout(n18084));
  jor  g17978(.dina(n14565), .dinb(n3429), .dout(n18085));
  jor  g17979(.dina(n17493), .dinb(n3426), .dout(n18086));
  jand g17980(.dina(n18086), .dinb(n18085), .dout(n18087));
  jor  g17981(.dina(n14567), .dinb(n3211), .dout(n18088));
  jand g17982(.dina(n18088), .dinb(n18087), .dout(n18089));
  jand g17983(.dina(n18089), .dinb(n18084), .dout(n18090));
  jxor g17984(.dina(n18090), .dinb(\a[14] ), .dout(n18091));
  jxor g17985(.dina(n18091), .dinb(n18082), .dout(n18092));
  jxor g17986(.dina(n18092), .dinb(n17983), .dout(n18093));
  jnot g17987(.din(n15831), .dout(n18094));
  jor  g17988(.dina(n18094), .dinb(n4023), .dout(n18095));
  jor  g17989(.dina(n17511), .dinb(n4028), .dout(n18096));
  jor  g17990(.dina(n17506), .dinb(n4025), .dout(n18097));
  jand g17991(.dina(n18097), .dinb(n18096), .dout(n18098));
  jor  g17992(.dina(n17495), .dinb(n3871), .dout(n18099));
  jand g17993(.dina(n18099), .dinb(n18098), .dout(n18100));
  jand g17994(.dina(n18100), .dinb(n18095), .dout(n18101));
  jxor g17995(.dina(n18101), .dinb(\a[11] ), .dout(n18102));
  jxor g17996(.dina(n18102), .dinb(n18093), .dout(n18103));
  jxor g17997(.dina(n18103), .dinb(n17978), .dout(n18104));
  jnot g17998(.din(n16594), .dout(n18105));
  jor  g17999(.dina(n18105), .dinb(n4692), .dout(n18106));
  jor  g18000(.dina(n17523), .dinb(n4697), .dout(n18107));
  jor  g18001(.dina(n17289), .dinb(n4705), .dout(n18108));
  jand g18002(.dina(n18108), .dinb(n18107), .dout(n18109));
  jor  g18003(.dina(n17508), .dinb(n4702), .dout(n18110));
  jand g18004(.dina(n18110), .dinb(n18109), .dout(n18111));
  jand g18005(.dina(n18111), .dinb(n18106), .dout(n18112));
  jxor g18006(.dina(n18112), .dinb(\a[8] ), .dout(n18113));
  jxor g18007(.dina(n18113), .dinb(n18104), .dout(n18114));
  jxor g18008(.dina(n18114), .dinb(n17973), .dout(n18115));
  jnot g18009(.din(n18115), .dout(n18116));
  jor  g18010(.dina(n18116), .dinb(n17960), .dout(n18117));
  jxor g18011(.dina(n18115), .dinb(n17960), .dout(n18118));
  jxor g18012(.dina(n17924), .dinb(n17956), .dout(n18119));
  jxor g18013(.dina(n17934), .dinb(n18119), .dout(n18120));
  jor  g18014(.dina(n18120), .dinb(n17735), .dout(n18121));
  jor  g18015(.dina(n17941), .dinb(n17936), .dout(n18122));
  jand g18016(.dina(n18122), .dinb(n18121), .dout(n18123));
  jor  g18017(.dina(n18123), .dinb(n18118), .dout(n18124));
  jand g18018(.dina(n18124), .dinb(n18117), .dout(n18125));
  jor  g18019(.dina(n18201), .dinb(n17965), .dout(n18126));
  jand g18020(.dina(n18114), .dinb(n17973), .dout(n18127));
  jnot g18021(.din(n18127), .dout(n18128));
  jand g18022(.dina(n18128), .dinb(n18126), .dout(n18129));
  jnot g18023(.din(n17983), .dout(n18130));
  jand g18024(.dina(n18092), .dinb(n18130), .dout(n18131));
  jnot g18025(.din(n18131), .dout(n18132));
  jor  g18026(.dina(n18102), .dinb(n18093), .dout(n18133));
  jand g18027(.dina(n18133), .dinb(n18132), .dout(n18134));
  jnot g18028(.din(n17987), .dout(n18135));
  jand g18029(.dina(n18081), .dinb(n18135), .dout(n18136));
  jnot g18030(.din(n18136), .dout(n18137));
  jor  g18031(.dina(n18091), .dinb(n18082), .dout(n18138));
  jand g18032(.dina(n18138), .dinb(n18137), .dout(n18139));
  jnot g18033(.din(n17991), .dout(n18140));
  jand g18034(.dina(n18071), .dinb(n18140), .dout(n18141));
  jnot g18035(.din(n18141), .dout(n18142));
  jor  g18036(.dina(n18080), .dinb(n18072), .dout(n18143));
  jand g18037(.dina(n18143), .dinb(n18142), .dout(n18144));
  jnot g18038(.din(n18144), .dout(n18145));
  jnot g18039(.din(n18061), .dout(n18146));
  jor  g18040(.dina(n18146), .dinb(n17995), .dout(n18147));
  jor  g18041(.dina(n18070), .dinb(n18062), .dout(n18148));
  jand g18042(.dina(n18148), .dinb(n18147), .dout(n18149));
  jnot g18043(.din(n18051), .dout(n18150));
  jor  g18044(.dina(n18150), .dinb(n17999), .dout(n18151));
  jor  g18045(.dina(n18060), .dinb(n18052), .dout(n18152));
  jand g18046(.dina(n18152), .dinb(n18151), .dout(n18153));
  jnot g18047(.din(n18033), .dout(n18154));
  jor  g18048(.dina(n18041), .dinb(n18154), .dout(n18155));
  jor  g18049(.dina(n18050), .dinb(n18042), .dout(n18156));
  jand g18050(.dina(n18156), .dinb(n18155), .dout(n18157));
  jnot g18051(.din(n18009), .dout(n18158));
  jnot g18052(.din(n18031), .dout(n18159));
  jor  g18053(.dina(n18159), .dinb(n18158), .dout(n18160));
  jnot g18054(.din(n18002), .dout(n18161));
  jnot g18055(.din(n18032), .dout(n18162));
  jor  g18056(.dina(n18162), .dinb(n18161), .dout(n18163));
  jand g18057(.dina(n18163), .dinb(n18160), .dout(n18164));
  jand g18058(.dina(n10850), .dinb(n5076), .dout(n18165));
  jand g18059(.dina(n10640), .dinb(n5084), .dout(n18166));
  jand g18060(.dina(n10647), .dinb(n5082), .dout(n18167));
  jand g18061(.dina(n10305), .dinb(n6050), .dout(n18168));
  jor  g18062(.dina(n18168), .dinb(n18167), .dout(n18169));
  jor  g18063(.dina(n18169), .dinb(n18166), .dout(n18170));
  jor  g18064(.dina(n18170), .dinb(n18165), .dout(n18171));
  jor  g18065(.dina(n18029), .dinb(n17422), .dout(n18172));
  jnot g18066(.din(n18172), .dout(n18173));
  jand g18067(.dina(n18030), .dinb(n18013), .dout(n18174));
  jor  g18068(.dina(n18174), .dinb(n18173), .dout(n18175));
  jand g18069(.dina(n3842), .dinb(n352), .dout(n18176));
  jand g18070(.dina(n558), .dinb(n447), .dout(n18177));
  jand g18071(.dina(n678), .dinb(n1738), .dout(n18178));
  jand g18072(.dina(n18178), .dinb(n1821), .dout(n18179));
  jand g18073(.dina(n18179), .dinb(n18177), .dout(n18180));
  jand g18074(.dina(n411), .dinb(n808), .dout(n18181));
  jand g18075(.dina(n18181), .dinb(n1207), .dout(n18182));
  jand g18076(.dina(n18182), .dinb(n18180), .dout(n18183));
  jand g18077(.dina(n18183), .dinb(n18176), .dout(n18184));
  jand g18078(.dina(n1454), .dinb(n114), .dout(n18185));
  jand g18079(.dina(n18185), .dinb(n9125), .dout(n18186));
  jand g18080(.dina(n1317), .dinb(n172), .dout(n18187));
  jand g18081(.dina(n18187), .dinb(n1088), .dout(n18188));
  jand g18082(.dina(n18188), .dinb(n18186), .dout(n18189));
  jand g18083(.dina(n18189), .dinb(n7502), .dout(n18190));
  jand g18084(.dina(n18190), .dinb(n18184), .dout(n18191));
  jand g18085(.dina(n8820), .dinb(n3322), .dout(n18192));
  jand g18086(.dina(n18192), .dinb(n5378), .dout(n18193));
  jand g18087(.dina(n18193), .dinb(n8622), .dout(n18194));
  jand g18088(.dina(n18194), .dinb(n13548), .dout(n18195));
  jand g18089(.dina(n18195), .dinb(n18191), .dout(n18196));
  jand g18090(.dina(n18196), .dinb(n17810), .dout(n18197));
  jxor g18091(.dina(n18197), .dinb(n17781), .dout(n18198));
  jor  g18092(.dina(n5534), .dinb(n5278), .dout(n18199));
  jand g18093(.dina(n18199), .dinb(n16924), .dout(n18200));
  jxor g18094(.dina(n18200), .dinb(n5277), .dout(n18201));
  jxor g18095(.dina(n18201), .dinb(n18198), .dout(n18202));
  jxor g18096(.dina(n18202), .dinb(n18175), .dout(n18203));
  jxor g18097(.dina(n18203), .dinb(n18171), .dout(n18204));
  jnot g18098(.din(n18204), .dout(n18205));
  jxor g18099(.dina(n18205), .dinb(n18164), .dout(n18206));
  jand g18100(.dina(n11824), .dinb(n2936), .dout(n18207));
  jand g18101(.dina(n11306), .dinb(n2940), .dout(n18208));
  jand g18102(.dina(n11647), .dinb(n2943), .dout(n18209));
  jor  g18103(.dina(n18209), .dinb(n18208), .dout(n18210));
  jand g18104(.dina(n10836), .dinb(n3684), .dout(n18211));
  jor  g18105(.dina(n18211), .dinb(n18210), .dout(n18212));
  jor  g18106(.dina(n18212), .dinb(n18207), .dout(n18213));
  jxor g18107(.dina(n18213), .dinb(n93), .dout(n18214));
  jxor g18108(.dina(n18214), .dinb(n18206), .dout(n18215));
  jand g18109(.dina(n12284), .dinb(n71), .dout(n18216));
  jand g18110(.dina(n11798), .dinb(n731), .dout(n18217));
  jand g18111(.dina(n12282), .dinb(n796), .dout(n18218));
  jor  g18112(.dina(n18218), .dinb(n18217), .dout(n18219));
  jand g18113(.dina(n11646), .dinb(n1806), .dout(n18220));
  jor  g18114(.dina(n18220), .dinb(n18219), .dout(n18221));
  jor  g18115(.dina(n18221), .dinb(n18216), .dout(n18222));
  jxor g18116(.dina(n18222), .dinb(n77), .dout(n18223));
  jxor g18117(.dina(n18223), .dinb(n18215), .dout(n18224));
  jxor g18118(.dina(n18224), .dinb(n18157), .dout(n18225));
  jand g18119(.dina(n12671), .dinb(n806), .dout(n18226));
  jand g18120(.dina(n12536), .dinb(n1612), .dout(n18227));
  jand g18121(.dina(n12669), .dinb(n1620), .dout(n18228));
  jor  g18122(.dina(n18228), .dinb(n18227), .dout(n18229));
  jand g18123(.dina(n12547), .dinb(n1644), .dout(n18230));
  jor  g18124(.dina(n18230), .dinb(n18229), .dout(n18231));
  jor  g18125(.dina(n18231), .dinb(n18226), .dout(n18232));
  jxor g18126(.dina(n18232), .dinb(n65), .dout(n18233));
  jxor g18127(.dina(n18233), .dinb(n18225), .dout(n18234));
  jxor g18128(.dina(n18234), .dinb(n18153), .dout(n18235));
  jand g18129(.dina(n13627), .dinb(n1819), .dout(n18236));
  jand g18130(.dina(n13478), .dinb(n2180), .dout(n18237));
  jand g18131(.dina(n13469), .dinb(n2243), .dout(n18238));
  jor  g18132(.dina(n18238), .dinb(n18237), .dout(n18239));
  jand g18133(.dina(n13248), .dinb(n2185), .dout(n18240));
  jor  g18134(.dina(n18240), .dinb(n18239), .dout(n18241));
  jor  g18135(.dina(n18241), .dinb(n18236), .dout(n18242));
  jxor g18136(.dina(n18242), .dinb(n2196), .dout(n18243));
  jxor g18137(.dina(n18243), .dinb(n18235), .dout(n18244));
  jxor g18138(.dina(n18244), .dinb(n18149), .dout(n18245));
  jand g18139(.dina(n14579), .dinb(n2743), .dout(n18246));
  jand g18140(.dina(n14448), .dinb(n2752), .dout(n18247));
  jand g18141(.dina(n14249), .dinb(n2748), .dout(n18248));
  jand g18142(.dina(n13614), .dinb(n2757), .dout(n18249));
  jor  g18143(.dina(n18249), .dinb(n18248), .dout(n18250));
  jor  g18144(.dina(n18250), .dinb(n18247), .dout(n18251));
  jor  g18145(.dina(n18251), .dinb(n18246), .dout(n18252));
  jxor g18146(.dina(n18252), .dinb(n2441), .dout(n18253));
  jxor g18147(.dina(n18253), .dinb(n18245), .dout(n18254));
  jxor g18148(.dina(n18254), .dinb(n18145), .dout(n18255));
  jand g18149(.dina(n15317), .dinb(n3423), .dout(n18256));
  jand g18150(.dina(n14549), .dinb(n3428), .dout(n18257));
  jand g18151(.dina(n15315), .dinb(n3569), .dout(n18258));
  jor  g18152(.dina(n18258), .dinb(n18257), .dout(n18259));
  jand g18153(.dina(n14447), .dinb(n3210), .dout(n18260));
  jor  g18154(.dina(n18260), .dinb(n18259), .dout(n18261));
  jor  g18155(.dina(n18261), .dinb(n18256), .dout(n18262));
  jxor g18156(.dina(n18262), .dinb(n3473), .dout(n18263));
  jxor g18157(.dina(n18263), .dinb(n18255), .dout(n18264));
  jxor g18158(.dina(n18264), .dinb(n18139), .dout(n18265));
  jor  g18159(.dina(n17504), .dinb(n4023), .dout(n18266));
  jor  g18160(.dina(n17506), .dinb(n4028), .dout(n18267));
  jor  g18161(.dina(n17508), .dinb(n4025), .dout(n18268));
  jand g18162(.dina(n18268), .dinb(n18267), .dout(n18269));
  jor  g18163(.dina(n17511), .dinb(n3871), .dout(n18270));
  jand g18164(.dina(n18270), .dinb(n18269), .dout(n18271));
  jand g18165(.dina(n18271), .dinb(n18266), .dout(n18272));
  jxor g18166(.dina(n18272), .dinb(\a[11] ), .dout(n18273));
  jxor g18167(.dina(n18273), .dinb(n18265), .dout(n18274));
  jxor g18168(.dina(n18274), .dinb(n18134), .dout(n18275));
  jnot g18169(.din(n17978), .dout(n18276));
  jand g18170(.dina(n18103), .dinb(n18276), .dout(n18277));
  jnot g18171(.din(n18277), .dout(n18278));
  jor  g18172(.dina(n18113), .dinb(n18104), .dout(n18279));
  jand g18173(.dina(n18279), .dinb(n18278), .dout(n18280));
  jor  g18174(.dina(n17518), .dinb(n4692), .dout(n18281));
  jor  g18175(.dina(n17289), .dinb(n4697), .dout(n18282));
  jor  g18176(.dina(n17288), .dinb(n4705), .dout(n18283));
  jand g18177(.dina(n18283), .dinb(n18282), .dout(n18284));
  jor  g18178(.dina(n17523), .dinb(n4702), .dout(n18285));
  jand g18179(.dina(n18285), .dinb(n18284), .dout(n18286));
  jand g18180(.dina(n18286), .dinb(n18281), .dout(n18287));
  jxor g18181(.dina(n18287), .dinb(\a[8] ), .dout(n18288));
  jxor g18182(.dina(n18288), .dinb(n18280), .dout(n18289));
  jxor g18183(.dina(n18289), .dinb(n18275), .dout(n18290));
  jxor g18184(.dina(n18290), .dinb(n18129), .dout(n18291));
  jxor g18185(.dina(n18291), .dinb(n18125), .dout(n18292));
  jxor g18186(.dina(n18123), .dinb(n18118), .dout(n18293));
  jand g18187(.dina(n18293), .dinb(n18292), .dout(n18294));
  jand g18188(.dina(n18293), .dinb(n17942), .dout(n18295));
  jand g18189(.dina(n17942), .dinb(n17535), .dout(n18296));
  jand g18190(.dina(n17943), .dinb(n17730), .dout(n18297));
  jor  g18191(.dina(n18297), .dinb(n18296), .dout(n18298));
  jxor g18192(.dina(n18293), .dinb(n17942), .dout(n18299));
  jand g18193(.dina(n18299), .dinb(n18298), .dout(n18300));
  jor  g18194(.dina(n18300), .dinb(n18295), .dout(n18301));
  jxor g18195(.dina(n18293), .dinb(n18292), .dout(n18302));
  jand g18196(.dina(n18302), .dinb(n18301), .dout(n18303));
  jor  g18197(.dina(n18303), .dinb(n18294), .dout(n18304));
  jnot g18198(.din(n18290), .dout(n18305));
  jor  g18199(.dina(n18305), .dinb(n18129), .dout(n18306));
  jor  g18200(.dina(n18291), .dinb(n18125), .dout(n18307));
  jand g18201(.dina(n18307), .dinb(n18306), .dout(n18308));
  jor  g18202(.dina(n18288), .dinb(n18280), .dout(n18309));
  jand g18203(.dina(n18289), .dinb(n18275), .dout(n18310));
  jnot g18204(.din(n18310), .dout(n18311));
  jand g18205(.dina(n18311), .dinb(n18309), .dout(n18312));
  jxor g18206(.dina(n18254), .dinb(n18144), .dout(n18313));
  jxor g18207(.dina(n18263), .dinb(n18313), .dout(n18314));
  jxor g18208(.dina(n18314), .dinb(n18139), .dout(n18315));
  jor  g18209(.dina(n18273), .dinb(n18315), .dout(n18316));
  jor  g18210(.dina(n18274), .dinb(n18134), .dout(n18317));
  jand g18211(.dina(n18317), .dinb(n18316), .dout(n18318));
  jor  g18212(.dina(n18263), .dinb(n18313), .dout(n18319));
  jor  g18213(.dina(n18264), .dinb(n18139), .dout(n18320));
  jand g18214(.dina(n18320), .dinb(n18319), .dout(n18321));
  jor  g18215(.dina(n18253), .dinb(n18245), .dout(n18322));
  jnot g18216(.din(n18322), .dout(n18323));
  jand g18217(.dina(n18254), .dinb(n18145), .dout(n18324));
  jor  g18218(.dina(n18324), .dinb(n18323), .dout(n18325));
  jor  g18219(.dina(n18243), .dinb(n18235), .dout(n18326));
  jxor g18220(.dina(n18204), .dinb(n18164), .dout(n18327));
  jxor g18221(.dina(n18214), .dinb(n18327), .dout(n18328));
  jxor g18222(.dina(n18223), .dinb(n18328), .dout(n18329));
  jxor g18223(.dina(n18329), .dinb(n18157), .dout(n18330));
  jxor g18224(.dina(n18233), .dinb(n18330), .dout(n18331));
  jxor g18225(.dina(n18331), .dinb(n18153), .dout(n18332));
  jxor g18226(.dina(n18243), .dinb(n18332), .dout(n18333));
  jor  g18227(.dina(n18333), .dinb(n18149), .dout(n18334));
  jand g18228(.dina(n18334), .dinb(n18326), .dout(n18335));
  jor  g18229(.dina(n18233), .dinb(n18225), .dout(n18336));
  jor  g18230(.dina(n18331), .dinb(n18153), .dout(n18337));
  jand g18231(.dina(n18337), .dinb(n18336), .dout(n18338));
  jor  g18232(.dina(n18223), .dinb(n18215), .dout(n18339));
  jor  g18233(.dina(n18329), .dinb(n18157), .dout(n18340));
  jand g18234(.dina(n18340), .dinb(n18339), .dout(n18341));
  jor  g18235(.dina(n18205), .dinb(n18164), .dout(n18342));
  jor  g18236(.dina(n18214), .dinb(n18327), .dout(n18343));
  jand g18237(.dina(n18343), .dinb(n18342), .dout(n18344));
  jand g18238(.dina(n18202), .dinb(n18175), .dout(n18345));
  jand g18239(.dina(n18203), .dinb(n18171), .dout(n18346));
  jor  g18240(.dina(n18346), .dinb(n18345), .dout(n18347));
  jand g18241(.dina(n1247), .dinb(n713), .dout(n18348));
  jand g18242(.dina(n18348), .dinb(n12434), .dout(n18349));
  jand g18243(.dina(n1753), .dinb(n907), .dout(n18350));
  jand g18244(.dina(n18350), .dinb(n3750), .dout(n18351));
  jand g18245(.dina(n18351), .dinb(n18349), .dout(n18352));
  jand g18246(.dina(n2586), .dinb(n1461), .dout(n18353));
  jand g18247(.dina(n18353), .dinb(n16195), .dout(n18354));
  jand g18248(.dina(n988), .dinb(n1429), .dout(n18355));
  jand g18249(.dina(n18355), .dinb(n428), .dout(n18356));
  jand g18250(.dina(n632), .dinb(n2148), .dout(n18357));
  jand g18251(.dina(n18357), .dinb(n18356), .dout(n18358));
  jand g18252(.dina(n18358), .dinb(n18354), .dout(n18359));
  jand g18253(.dina(n1707), .dinb(n6441), .dout(n18360));
  jand g18254(.dina(n18360), .dinb(n818), .dout(n18361));
  jand g18255(.dina(n18361), .dinb(n5466), .dout(n18362));
  jand g18256(.dina(n18362), .dinb(n18359), .dout(n18363));
  jand g18257(.dina(n18363), .dinb(n18352), .dout(n18364));
  jand g18258(.dina(n12219), .dinb(n3178), .dout(n18365));
  jand g18259(.dina(n5253), .dinb(n4639), .dout(n18366));
  jand g18260(.dina(n18366), .dinb(n18365), .dout(n18367));
  jand g18261(.dina(n18367), .dinb(n499), .dout(n18368));
  jand g18262(.dina(n981), .dinb(n660), .dout(n18369));
  jand g18263(.dina(n553), .dinb(n991), .dout(n18370));
  jand g18264(.dina(n18370), .dinb(n18369), .dout(n18371));
  jand g18265(.dina(n18371), .dinb(n2663), .dout(n18372));
  jand g18266(.dina(n18372), .dinb(n5978), .dout(n18373));
  jand g18267(.dina(n18373), .dinb(n18368), .dout(n18374));
  jand g18268(.dina(n1365), .dinb(n619), .dout(n18375));
  jand g18269(.dina(n18375), .dinb(n600), .dout(n18376));
  jand g18270(.dina(n18376), .dinb(n1470), .dout(n18377));
  jand g18271(.dina(n6343), .dinb(n1743), .dout(n18378));
  jand g18272(.dina(n680), .dinb(n933), .dout(n18379));
  jand g18273(.dina(n18379), .dinb(n3989), .dout(n18380));
  jand g18274(.dina(n18380), .dinb(n18378), .dout(n18381));
  jand g18275(.dina(n2023), .dinb(n1366), .dout(n18382));
  jand g18276(.dina(n18382), .dinb(n1538), .dout(n18383));
  jand g18277(.dina(n18383), .dinb(n18381), .dout(n18384));
  jand g18278(.dina(n18384), .dinb(n18377), .dout(n18385));
  jand g18279(.dina(n18385), .dinb(n18374), .dout(n18386));
  jand g18280(.dina(n5353), .dinb(n1272), .dout(n18387));
  jand g18281(.dina(n18387), .dinb(n18386), .dout(n18388));
  jand g18282(.dina(n18388), .dinb(n1986), .dout(n18389));
  jand g18283(.dina(n18389), .dinb(n18364), .dout(n18390));
  jnot g18284(.din(n18390), .dout(n18391));
  jor  g18285(.dina(n18197), .dinb(n17781), .dout(n18392));
  jand g18286(.dina(n18201), .dinb(n18198), .dout(n18393));
  jnot g18287(.din(n18393), .dout(n18394));
  jand g18288(.dina(n18394), .dinb(n18392), .dout(n18395));
  jxor g18289(.dina(n18395), .dinb(n18391), .dout(n18396));
  jand g18290(.dina(n10838), .dinb(n5076), .dout(n18397));
  jand g18291(.dina(n10836), .dinb(n5084), .dout(n18398));
  jand g18292(.dina(n10647), .dinb(n6050), .dout(n18399));
  jand g18293(.dina(n10640), .dinb(n5082), .dout(n18400));
  jor  g18294(.dina(n18400), .dinb(n18399), .dout(n18401));
  jor  g18295(.dina(n18401), .dinb(n18398), .dout(n18402));
  jor  g18296(.dina(n18402), .dinb(n18397), .dout(n18403));
  jxor g18297(.dina(n18403), .dinb(n18396), .dout(n18404));
  jxor g18298(.dina(n18404), .dinb(n18347), .dout(n18405));
  jand g18299(.dina(n11812), .dinb(n2936), .dout(n18406));
  jand g18300(.dina(n11646), .dinb(n2943), .dout(n18407));
  jand g18301(.dina(n11647), .dinb(n2940), .dout(n18408));
  jand g18302(.dina(n11306), .dinb(n3684), .dout(n18409));
  jor  g18303(.dina(n18409), .dinb(n18408), .dout(n18410));
  jor  g18304(.dina(n18410), .dinb(n18407), .dout(n18411));
  jor  g18305(.dina(n18411), .dinb(n18406), .dout(n18412));
  jxor g18306(.dina(n18412), .dinb(n93), .dout(n18413));
  jnot g18307(.din(n18413), .dout(n18414));
  jxor g18308(.dina(n18414), .dinb(n18405), .dout(n18415));
  jxor g18309(.dina(n18415), .dinb(n18344), .dout(n18416));
  jand g18310(.dina(n12696), .dinb(n71), .dout(n18417));
  jand g18311(.dina(n12282), .dinb(n731), .dout(n18418));
  jand g18312(.dina(n12547), .dinb(n796), .dout(n18419));
  jor  g18313(.dina(n18419), .dinb(n18418), .dout(n18420));
  jand g18314(.dina(n11798), .dinb(n1806), .dout(n18421));
  jor  g18315(.dina(n18421), .dinb(n18420), .dout(n18422));
  jor  g18316(.dina(n18422), .dinb(n18417), .dout(n18423));
  jxor g18317(.dina(n18423), .dinb(n77), .dout(n18424));
  jxor g18318(.dina(n18424), .dinb(n18416), .dout(n18425));
  jxor g18319(.dina(n18425), .dinb(n18341), .dout(n18426));
  jand g18320(.dina(n13250), .dinb(n806), .dout(n18427));
  jand g18321(.dina(n12669), .dinb(n1612), .dout(n18428));
  jand g18322(.dina(n13248), .dinb(n1620), .dout(n18429));
  jor  g18323(.dina(n18429), .dinb(n18428), .dout(n18430));
  jand g18324(.dina(n12536), .dinb(n1644), .dout(n18431));
  jor  g18325(.dina(n18431), .dinb(n18430), .dout(n18432));
  jor  g18326(.dina(n18432), .dinb(n18427), .dout(n18433));
  jxor g18327(.dina(n18433), .dinb(n65), .dout(n18434));
  jxor g18328(.dina(n18434), .dinb(n18426), .dout(n18435));
  jxor g18329(.dina(n18435), .dinb(n18338), .dout(n18436));
  jand g18330(.dina(n13616), .dinb(n1819), .dout(n18437));
  jand g18331(.dina(n13614), .dinb(n2243), .dout(n18438));
  jand g18332(.dina(n13469), .dinb(n2180), .dout(n18439));
  jand g18333(.dina(n13478), .dinb(n2185), .dout(n18440));
  jor  g18334(.dina(n18440), .dinb(n18439), .dout(n18441));
  jor  g18335(.dina(n18441), .dinb(n18438), .dout(n18442));
  jor  g18336(.dina(n18442), .dinb(n18437), .dout(n18443));
  jxor g18337(.dina(n18443), .dinb(n2196), .dout(n18444));
  jxor g18338(.dina(n18444), .dinb(n18436), .dout(n18445));
  jxor g18339(.dina(n18445), .dinb(n18335), .dout(n18446));
  jand g18340(.dina(n14562), .dinb(n2743), .dout(n18447));
  jand g18341(.dina(n14447), .dinb(n2752), .dout(n18448));
  jand g18342(.dina(n14448), .dinb(n2748), .dout(n18449));
  jand g18343(.dina(n14249), .dinb(n2757), .dout(n18450));
  jor  g18344(.dina(n18450), .dinb(n18449), .dout(n18451));
  jor  g18345(.dina(n18451), .dinb(n18448), .dout(n18452));
  jor  g18346(.dina(n18452), .dinb(n18447), .dout(n18453));
  jxor g18347(.dina(n18453), .dinb(n2441), .dout(n18454));
  jxor g18348(.dina(n18454), .dinb(n18446), .dout(n18455));
  jxor g18349(.dina(n18455), .dinb(n18325), .dout(n18456));
  jnot g18350(.din(n18456), .dout(n18457));
  jor  g18351(.dina(n17904), .dinb(n3424), .dout(n18458));
  jor  g18352(.dina(n17495), .dinb(n3429), .dout(n18459));
  jor  g18353(.dina(n17511), .dinb(n3426), .dout(n18460));
  jand g18354(.dina(n18460), .dinb(n18459), .dout(n18461));
  jor  g18355(.dina(n17493), .dinb(n3211), .dout(n18462));
  jand g18356(.dina(n18462), .dinb(n18461), .dout(n18463));
  jand g18357(.dina(n18463), .dinb(n18458), .dout(n18464));
  jxor g18358(.dina(n18464), .dinb(\a[14] ), .dout(n18465));
  jxor g18359(.dina(n18465), .dinb(n18457), .dout(n18466));
  jxor g18360(.dina(n18466), .dinb(n18321), .dout(n18467));
  jand g18361(.dina(n16345), .dinb(n4022), .dout(n18468));
  jand g18362(.dina(n16082), .dinb(n4027), .dout(n18469));
  jand g18363(.dina(n16343), .dinb(n4220), .dout(n18470));
  jor  g18364(.dina(n18470), .dinb(n18469), .dout(n18471));
  jand g18365(.dina(n15829), .dinb(n3870), .dout(n18472));
  jor  g18366(.dina(n18472), .dinb(n18471), .dout(n18473));
  jor  g18367(.dina(n18473), .dinb(n18468), .dout(n18474));
  jxor g18368(.dina(n18474), .dinb(n4050), .dout(n18475));
  jxor g18369(.dina(n18475), .dinb(n18467), .dout(n18476));
  jxor g18370(.dina(n18476), .dinb(n18318), .dout(n18477));
  jor  g18371(.dina(n17926), .dinb(n4692), .dout(n18478));
  jor  g18372(.dina(n17289), .dinb(n4702), .dout(n18479));
  jand g18373(.dina(n18775), .dinb(n18479), .dout(n18483));
  jand g18374(.dina(n18483), .dinb(n18478), .dout(n18484));
  jxor g18375(.dina(n18484), .dinb(\a[8] ), .dout(n18485));
  jxor g18376(.dina(n18485), .dinb(n18477), .dout(n18486));
  jxor g18377(.dina(n18486), .dinb(n18312), .dout(n18487));
  jxor g18378(.dina(n18487), .dinb(n18308), .dout(n18488));
  jxor g18379(.dina(n18488), .dinb(n18292), .dout(n18489));
  jxor g18380(.dina(n18489), .dinb(n18304), .dout(n18490));
  jand g18381(.dina(n18490), .dinb(n2743), .dout(n18491));
  jand g18382(.dina(n18488), .dinb(n2752), .dout(n18492));
  jand g18383(.dina(n18292), .dinb(n2748), .dout(n18493));
  jand g18384(.dina(n18293), .dinb(n2757), .dout(n18494));
  jor  g18385(.dina(n18494), .dinb(n18493), .dout(n18495));
  jor  g18386(.dina(n18495), .dinb(n18492), .dout(n18496));
  jor  g18387(.dina(n18496), .dinb(n18491), .dout(n18497));
  jxor g18388(.dina(n18497), .dinb(n2441), .dout(n18498));
  jor  g18389(.dina(n18498), .dinb(n17955), .dout(n18499));
  jxor g18390(.dina(n17679), .dinb(n17678), .dout(n18500));
  jnot g18391(.din(n18500), .dout(n18501));
  jxor g18392(.dina(n18302), .dinb(n18301), .dout(n18502));
  jand g18393(.dina(n18502), .dinb(n2743), .dout(n18503));
  jand g18394(.dina(n18292), .dinb(n2752), .dout(n18504));
  jand g18395(.dina(n18293), .dinb(n2748), .dout(n18505));
  jand g18396(.dina(n17942), .dinb(n2757), .dout(n18506));
  jor  g18397(.dina(n18506), .dinb(n18505), .dout(n18507));
  jor  g18398(.dina(n18507), .dinb(n18504), .dout(n18508));
  jor  g18399(.dina(n18508), .dinb(n18503), .dout(n18509));
  jxor g18400(.dina(n18509), .dinb(n2441), .dout(n18510));
  jor  g18401(.dina(n18510), .dinb(n18501), .dout(n18511));
  jxor g18402(.dina(n17674), .dinb(n17673), .dout(n18512));
  jnot g18403(.din(n18512), .dout(n18513));
  jxor g18404(.dina(n18299), .dinb(n18298), .dout(n18514));
  jand g18405(.dina(n18514), .dinb(n2743), .dout(n18515));
  jand g18406(.dina(n18293), .dinb(n2752), .dout(n18516));
  jand g18407(.dina(n17942), .dinb(n2748), .dout(n18517));
  jand g18408(.dina(n17535), .dinb(n2757), .dout(n18518));
  jor  g18409(.dina(n18518), .dinb(n18517), .dout(n18519));
  jor  g18410(.dina(n18519), .dinb(n18516), .dout(n18520));
  jor  g18411(.dina(n18520), .dinb(n18515), .dout(n18521));
  jxor g18412(.dina(n18521), .dinb(n2441), .dout(n18522));
  jor  g18413(.dina(n18522), .dinb(n18513), .dout(n18523));
  jxor g18414(.dina(n17669), .dinb(n17668), .dout(n18524));
  jnot g18415(.din(n18524), .dout(n18525));
  jand g18416(.dina(n17944), .dinb(n2743), .dout(n18526));
  jand g18417(.dina(n17942), .dinb(n2752), .dout(n18527));
  jand g18418(.dina(n17535), .dinb(n2748), .dout(n18528));
  jand g18419(.dina(n17329), .dinb(n2757), .dout(n18529));
  jor  g18420(.dina(n18529), .dinb(n18528), .dout(n18530));
  jor  g18421(.dina(n18530), .dinb(n18527), .dout(n18531));
  jor  g18422(.dina(n18531), .dinb(n18526), .dout(n18532));
  jxor g18423(.dina(n18532), .dinb(n2441), .dout(n18533));
  jor  g18424(.dina(n18533), .dinb(n18525), .dout(n18534));
  jxor g18425(.dina(n17664), .dinb(n17663), .dout(n18535));
  jnot g18426(.din(n18535), .dout(n18536));
  jand g18427(.dina(n17537), .dinb(n2743), .dout(n18537));
  jand g18428(.dina(n17535), .dinb(n2752), .dout(n18538));
  jand g18429(.dina(n17329), .dinb(n2748), .dout(n18539));
  jand g18430(.dina(n17330), .dinb(n2757), .dout(n18540));
  jor  g18431(.dina(n18540), .dinb(n18539), .dout(n18541));
  jor  g18432(.dina(n18541), .dinb(n18538), .dout(n18542));
  jor  g18433(.dina(n18542), .dinb(n18537), .dout(n18543));
  jxor g18434(.dina(n18543), .dinb(n2441), .dout(n18544));
  jor  g18435(.dina(n18544), .dinb(n18536), .dout(n18545));
  jxor g18436(.dina(n17659), .dinb(n17658), .dout(n18546));
  jnot g18437(.din(n18546), .dout(n18547));
  jand g18438(.dina(n17549), .dinb(n2743), .dout(n18548));
  jand g18439(.dina(n17329), .dinb(n2752), .dout(n18549));
  jand g18440(.dina(n17330), .dinb(n2748), .dout(n18550));
  jand g18441(.dina(n16940), .dinb(n2757), .dout(n18551));
  jor  g18442(.dina(n18551), .dinb(n18550), .dout(n18552));
  jor  g18443(.dina(n18552), .dinb(n18549), .dout(n18553));
  jor  g18444(.dina(n18553), .dinb(n18548), .dout(n18554));
  jxor g18445(.dina(n18554), .dinb(n2441), .dout(n18555));
  jor  g18446(.dina(n18555), .dinb(n18547), .dout(n18556));
  jxor g18447(.dina(n17656), .dinb(n17655), .dout(n18557));
  jnot g18448(.din(n18557), .dout(n18558));
  jand g18449(.dina(n17561), .dinb(n2743), .dout(n18559));
  jand g18450(.dina(n16940), .dinb(n2748), .dout(n18560));
  jand g18451(.dina(n17330), .dinb(n2752), .dout(n18561));
  jor  g18452(.dina(n18561), .dinb(n18560), .dout(n18562));
  jand g18453(.dina(n16604), .dinb(n2757), .dout(n18563));
  jor  g18454(.dina(n18563), .dinb(n18562), .dout(n18564));
  jor  g18455(.dina(n18564), .dinb(n18559), .dout(n18565));
  jxor g18456(.dina(n18565), .dinb(n2441), .dout(n18566));
  jor  g18457(.dina(n18566), .dinb(n18558), .dout(n18567));
  jxor g18458(.dina(n17651), .dinb(n17650), .dout(n18568));
  jnot g18459(.din(n18568), .dout(n18569));
  jand g18460(.dina(n16942), .dinb(n2743), .dout(n18570));
  jand g18461(.dina(n16940), .dinb(n2752), .dout(n18571));
  jand g18462(.dina(n16604), .dinb(n2748), .dout(n18572));
  jand g18463(.dina(n16355), .dinb(n2757), .dout(n18573));
  jor  g18464(.dina(n18573), .dinb(n18572), .dout(n18574));
  jor  g18465(.dina(n18574), .dinb(n18571), .dout(n18575));
  jor  g18466(.dina(n18575), .dinb(n18570), .dout(n18576));
  jxor g18467(.dina(n18576), .dinb(n2441), .dout(n18577));
  jor  g18468(.dina(n18577), .dinb(n18569), .dout(n18578));
  jxor g18469(.dina(n17647), .dinb(n17639), .dout(n18579));
  jnot g18470(.din(n18579), .dout(n18580));
  jand g18471(.dina(n16606), .dinb(n2743), .dout(n18581));
  jand g18472(.dina(n16604), .dinb(n2752), .dout(n18582));
  jand g18473(.dina(n16355), .dinb(n2748), .dout(n18583));
  jand g18474(.dina(n16360), .dinb(n2757), .dout(n18584));
  jor  g18475(.dina(n18584), .dinb(n18583), .dout(n18585));
  jor  g18476(.dina(n18585), .dinb(n18582), .dout(n18586));
  jor  g18477(.dina(n18586), .dinb(n18581), .dout(n18587));
  jxor g18478(.dina(n18587), .dinb(n2441), .dout(n18588));
  jor  g18479(.dina(n18588), .dinb(n18580), .dout(n18589));
  jand g18480(.dina(n16616), .dinb(n2743), .dout(n18590));
  jand g18481(.dina(n16355), .dinb(n2752), .dout(n18591));
  jand g18482(.dina(n16360), .dinb(n2748), .dout(n18592));
  jand g18483(.dina(n15841), .dinb(n2757), .dout(n18593));
  jor  g18484(.dina(n18593), .dinb(n18592), .dout(n18594));
  jor  g18485(.dina(n18594), .dinb(n18591), .dout(n18595));
  jor  g18486(.dina(n18595), .dinb(n18590), .dout(n18596));
  jxor g18487(.dina(n18596), .dinb(n2441), .dout(n18597));
  jnot g18488(.din(n18597), .dout(n18598));
  jor  g18489(.dina(n17626), .dinb(n2196), .dout(n18599));
  jxor g18490(.dina(n18599), .dinb(n17634), .dout(n18600));
  jand g18491(.dina(n18600), .dinb(n18598), .dout(n18601));
  jand g18492(.dina(n17623), .dinb(\a[20] ), .dout(n18602));
  jxor g18493(.dina(n18602), .dinb(n17621), .dout(n18603));
  jnot g18494(.din(n18603), .dout(n18604));
  jand g18495(.dina(n16632), .dinb(n2743), .dout(n18605));
  jand g18496(.dina(n15841), .dinb(n2748), .dout(n18606));
  jand g18497(.dina(n16360), .dinb(n2752), .dout(n18607));
  jor  g18498(.dina(n18607), .dinb(n18606), .dout(n18608));
  jand g18499(.dina(n15579), .dinb(n2757), .dout(n18609));
  jor  g18500(.dina(n18609), .dinb(n18608), .dout(n18610));
  jor  g18501(.dina(n18610), .dinb(n18605), .dout(n18611));
  jxor g18502(.dina(n18611), .dinb(n2441), .dout(n18612));
  jor  g18503(.dina(n18612), .dinb(n18604), .dout(n18613));
  jand g18504(.dina(n15329), .dinb(n2743), .dout(n18614));
  jand g18505(.dina(n15020), .dinb(n2748), .dout(n18615));
  jand g18506(.dina(n15327), .dinb(n2752), .dout(n18616));
  jor  g18507(.dina(n18616), .dinb(n18615), .dout(n18617));
  jor  g18508(.dina(n18617), .dinb(n18614), .dout(n18618));
  jnot g18509(.din(n18618), .dout(n18619));
  jand g18510(.dina(n15020), .dinb(n2741), .dout(n18620));
  jnot g18511(.din(n18620), .dout(n18621));
  jand g18512(.dina(n18621), .dinb(\a[17] ), .dout(n18622));
  jand g18513(.dina(n18622), .dinb(n18619), .dout(n18623));
  jand g18514(.dina(n15580), .dinb(n2743), .dout(n18624));
  jand g18515(.dina(n15327), .dinb(n2748), .dout(n18625));
  jor  g18516(.dina(n18625), .dinb(n18624), .dout(n18626));
  jand g18517(.dina(n15579), .dinb(n2752), .dout(n18627));
  jand g18518(.dina(n15020), .dinb(n2757), .dout(n18628));
  jor  g18519(.dina(n18628), .dinb(n18627), .dout(n18629));
  jor  g18520(.dina(n18629), .dinb(n18626), .dout(n18630));
  jnot g18521(.din(n18630), .dout(n18631));
  jand g18522(.dina(n18631), .dinb(n18623), .dout(n18632));
  jand g18523(.dina(n18632), .dinb(n17623), .dout(n18633));
  jnot g18524(.din(n18633), .dout(n18634));
  jxor g18525(.dina(n18632), .dinb(n17623), .dout(n18635));
  jnot g18526(.din(n18635), .dout(n18636));
  jand g18527(.dina(n15848), .dinb(n2743), .dout(n18637));
  jand g18528(.dina(n15841), .dinb(n2752), .dout(n18638));
  jand g18529(.dina(n15579), .dinb(n2748), .dout(n18639));
  jand g18530(.dina(n15327), .dinb(n2757), .dout(n18640));
  jor  g18531(.dina(n18640), .dinb(n18639), .dout(n18641));
  jor  g18532(.dina(n18641), .dinb(n18638), .dout(n18642));
  jor  g18533(.dina(n18642), .dinb(n18637), .dout(n18643));
  jxor g18534(.dina(n18643), .dinb(n2441), .dout(n18644));
  jor  g18535(.dina(n18644), .dinb(n18636), .dout(n18645));
  jand g18536(.dina(n18645), .dinb(n18634), .dout(n18646));
  jnot g18537(.din(n18646), .dout(n18647));
  jxor g18538(.dina(n18612), .dinb(n18604), .dout(n18648));
  jand g18539(.dina(n18648), .dinb(n18647), .dout(n18649));
  jnot g18540(.din(n18649), .dout(n18650));
  jand g18541(.dina(n18650), .dinb(n18613), .dout(n18651));
  jnot g18542(.din(n18651), .dout(n18652));
  jxor g18543(.dina(n18600), .dinb(n18598), .dout(n18653));
  jand g18544(.dina(n18653), .dinb(n18652), .dout(n18654));
  jor  g18545(.dina(n18654), .dinb(n18601), .dout(n18655));
  jxor g18546(.dina(n18588), .dinb(n18580), .dout(n18656));
  jand g18547(.dina(n18656), .dinb(n18655), .dout(n18657));
  jnot g18548(.din(n18657), .dout(n18658));
  jand g18549(.dina(n18658), .dinb(n18589), .dout(n18659));
  jnot g18550(.din(n18659), .dout(n18660));
  jxor g18551(.dina(n18577), .dinb(n18569), .dout(n18661));
  jand g18552(.dina(n18661), .dinb(n18660), .dout(n18662));
  jnot g18553(.din(n18662), .dout(n18663));
  jand g18554(.dina(n18663), .dinb(n18578), .dout(n18664));
  jnot g18555(.din(n18664), .dout(n18665));
  jxor g18556(.dina(n18566), .dinb(n18558), .dout(n18666));
  jand g18557(.dina(n18666), .dinb(n18665), .dout(n18667));
  jnot g18558(.din(n18667), .dout(n18668));
  jand g18559(.dina(n18668), .dinb(n18567), .dout(n18669));
  jnot g18560(.din(n18669), .dout(n18670));
  jxor g18561(.dina(n18555), .dinb(n18547), .dout(n18671));
  jand g18562(.dina(n18671), .dinb(n18670), .dout(n18672));
  jnot g18563(.din(n18672), .dout(n18673));
  jand g18564(.dina(n18673), .dinb(n18556), .dout(n18674));
  jnot g18565(.din(n18674), .dout(n18675));
  jxor g18566(.dina(n18544), .dinb(n18536), .dout(n18676));
  jand g18567(.dina(n18676), .dinb(n18675), .dout(n18677));
  jnot g18568(.din(n18677), .dout(n18678));
  jand g18569(.dina(n18678), .dinb(n18545), .dout(n18679));
  jnot g18570(.din(n18679), .dout(n18680));
  jxor g18571(.dina(n18533), .dinb(n18525), .dout(n18681));
  jand g18572(.dina(n18681), .dinb(n18680), .dout(n18682));
  jnot g18573(.din(n18682), .dout(n18683));
  jand g18574(.dina(n18683), .dinb(n18534), .dout(n18684));
  jnot g18575(.din(n18684), .dout(n18685));
  jxor g18576(.dina(n18522), .dinb(n18513), .dout(n18686));
  jand g18577(.dina(n18686), .dinb(n18685), .dout(n18687));
  jnot g18578(.din(n18687), .dout(n18688));
  jand g18579(.dina(n18688), .dinb(n18523), .dout(n18689));
  jnot g18580(.din(n18689), .dout(n18690));
  jxor g18581(.dina(n18510), .dinb(n18501), .dout(n18691));
  jand g18582(.dina(n18691), .dinb(n18690), .dout(n18692));
  jnot g18583(.din(n18692), .dout(n18693));
  jand g18584(.dina(n18693), .dinb(n18511), .dout(n18694));
  jnot g18585(.din(n18694), .dout(n18695));
  jxor g18586(.dina(n18498), .dinb(n17955), .dout(n18696));
  jand g18587(.dina(n18696), .dinb(n18695), .dout(n18697));
  jnot g18588(.din(n18697), .dout(n18698));
  jand g18589(.dina(n18698), .dinb(n18499), .dout(n18699));
  jnot g18590(.din(n18699), .dout(n18700));
  jor  g18591(.dina(n17952), .dinb(n17727), .dout(n18701));
  jand g18592(.dina(n17953), .dinb(n17683), .dout(n18702));
  jnot g18593(.din(n18702), .dout(n18703));
  jand g18594(.dina(n18703), .dinb(n18701), .dout(n18704));
  jnot g18595(.din(n18704), .dout(n18705));
  jor  g18596(.dina(n17724), .dinb(n17716), .dout(n18706));
  jand g18597(.dina(n17725), .dinb(n17688), .dout(n18707));
  jnot g18598(.din(n18707), .dout(n18708));
  jand g18599(.dina(n18708), .dinb(n18706), .dout(n18709));
  jnot g18600(.din(n18709), .dout(n18710));
  jand g18601(.dina(n17713), .dinb(n17702), .dout(n18711));
  jand g18602(.dina(n17714), .dinb(n17693), .dout(n18712));
  jor  g18603(.dina(n18712), .dinb(n18711), .dout(n18713));
  jor  g18604(.dina(n17711), .dinb(n17709), .dout(n18714));
  jnot g18605(.din(n18714), .dout(n18715));
  jand g18606(.dina(n15020), .dinb(n4338), .dout(n18716));
  jxor g18607(.dina(n18716), .dinb(n18715), .dout(n18717));
  jnot g18608(.din(n18717), .dout(n18718));
  jand g18609(.dina(n15848), .dinb(n2936), .dout(n18719));
  jand g18610(.dina(n15579), .dinb(n2940), .dout(n18720));
  jand g18611(.dina(n15841), .dinb(n2943), .dout(n18721));
  jor  g18612(.dina(n18721), .dinb(n18720), .dout(n18722));
  jand g18613(.dina(n15327), .dinb(n3684), .dout(n18723));
  jor  g18614(.dina(n18723), .dinb(n18722), .dout(n18724));
  jor  g18615(.dina(n18724), .dinb(n18719), .dout(n18725));
  jxor g18616(.dina(n18725), .dinb(n93), .dout(n18726));
  jxor g18617(.dina(n18726), .dinb(n18718), .dout(n18727));
  jnot g18618(.din(n18727), .dout(n18728));
  jand g18619(.dina(n16606), .dinb(n71), .dout(n18729));
  jand g18620(.dina(n16355), .dinb(n731), .dout(n18730));
  jand g18621(.dina(n16604), .dinb(n796), .dout(n18731));
  jor  g18622(.dina(n18731), .dinb(n18730), .dout(n18732));
  jand g18623(.dina(n16360), .dinb(n1806), .dout(n18733));
  jor  g18624(.dina(n18733), .dinb(n18732), .dout(n18734));
  jor  g18625(.dina(n18734), .dinb(n18729), .dout(n18735));
  jxor g18626(.dina(n18735), .dinb(n77), .dout(n18736));
  jxor g18627(.dina(n18736), .dinb(n18728), .dout(n18737));
  jxor g18628(.dina(n18737), .dinb(n18713), .dout(n18738));
  jnot g18629(.din(n18738), .dout(n18739));
  jand g18630(.dina(n17549), .dinb(n806), .dout(n18740));
  jand g18631(.dina(n17329), .dinb(n1620), .dout(n18741));
  jand g18632(.dina(n17330), .dinb(n1612), .dout(n18742));
  jand g18633(.dina(n16940), .dinb(n1644), .dout(n18743));
  jor  g18634(.dina(n18743), .dinb(n18742), .dout(n18744));
  jor  g18635(.dina(n18744), .dinb(n18741), .dout(n18745));
  jor  g18636(.dina(n18745), .dinb(n18740), .dout(n18746));
  jxor g18637(.dina(n18746), .dinb(n65), .dout(n18747));
  jxor g18638(.dina(n18747), .dinb(n18739), .dout(n18748));
  jxor g18639(.dina(n18748), .dinb(n18710), .dout(n18749));
  jnot g18640(.din(n18749), .dout(n18750));
  jand g18641(.dina(n18514), .dinb(n1819), .dout(n18751));
  jand g18642(.dina(n17942), .dinb(n2180), .dout(n18752));
  jand g18643(.dina(n18293), .dinb(n2243), .dout(n18753));
  jor  g18644(.dina(n18753), .dinb(n18752), .dout(n18754));
  jand g18645(.dina(n17535), .dinb(n2185), .dout(n18755));
  jor  g18646(.dina(n18755), .dinb(n18754), .dout(n18756));
  jor  g18647(.dina(n18756), .dinb(n18751), .dout(n18757));
  jxor g18648(.dina(n18757), .dinb(n2196), .dout(n18758));
  jxor g18649(.dina(n18758), .dinb(n18750), .dout(n18759));
  jxor g18650(.dina(n18759), .dinb(n18705), .dout(n18760));
  jnot g18651(.din(n18760), .dout(n18761));
  jand g18652(.dina(n18488), .dinb(n18292), .dout(n18762));
  jand g18653(.dina(n18489), .dinb(n18304), .dout(n18763));
  jor  g18654(.dina(n18763), .dinb(n18762), .dout(n18764));
  jnot g18655(.din(n18318), .dout(n18765));
  jand g18656(.dina(n18476), .dinb(n18765), .dout(n18766));
  jnot g18657(.din(n18766), .dout(n18767));
  jor  g18658(.dina(n18485), .dinb(n18477), .dout(n18768));
  jand g18659(.dina(n18768), .dinb(n18767), .dout(n18769));
  jnot g18660(.din(n18466), .dout(n18770));
  jor  g18661(.dina(n18770), .dinb(n18321), .dout(n18771));
  jor  g18662(.dina(n18475), .dinb(n18467), .dout(n18772));
  jand g18663(.dina(n18772), .dinb(n18771), .dout(n18773));
  jor  g18664(.dina(n4700), .dinb(n4691), .dout(n18774));
  jor  g18665(.dina(n18774), .dinb(n17301), .dout(n18775));
  jxor g18666(.dina(n18994), .dinb(n18773), .dout(n18781));
  jand g18667(.dina(n18455), .dinb(n18325), .dout(n18782));
  jnot g18668(.din(n18782), .dout(n18783));
  jor  g18669(.dina(n18465), .dinb(n18457), .dout(n18784));
  jand g18670(.dina(n18784), .dinb(n18783), .dout(n18785));
  jnot g18671(.din(n18445), .dout(n18786));
  jor  g18672(.dina(n18786), .dinb(n18335), .dout(n18787));
  jor  g18673(.dina(n18454), .dinb(n18446), .dout(n18788));
  jand g18674(.dina(n18788), .dinb(n18787), .dout(n18789));
  jnot g18675(.din(n18789), .dout(n18790));
  jnot g18676(.din(n18435), .dout(n18791));
  jor  g18677(.dina(n18791), .dinb(n18338), .dout(n18792));
  jor  g18678(.dina(n18444), .dinb(n18436), .dout(n18793));
  jand g18679(.dina(n18793), .dinb(n18792), .dout(n18794));
  jnot g18680(.din(n18425), .dout(n18795));
  jor  g18681(.dina(n18795), .dinb(n18341), .dout(n18796));
  jor  g18682(.dina(n18434), .dinb(n18426), .dout(n18797));
  jand g18683(.dina(n18797), .dinb(n18796), .dout(n18798));
  jnot g18684(.din(n18415), .dout(n18799));
  jor  g18685(.dina(n18799), .dinb(n18344), .dout(n18800));
  jor  g18686(.dina(n18424), .dinb(n18416), .dout(n18801));
  jand g18687(.dina(n18801), .dinb(n18800), .dout(n18802));
  jand g18688(.dina(n18404), .dinb(n18347), .dout(n18803));
  jand g18689(.dina(n18414), .dinb(n18405), .dout(n18804));
  jor  g18690(.dina(n18804), .dinb(n18803), .dout(n18805));
  jand g18691(.dina(n11308), .dinb(n5076), .dout(n18806));
  jand g18692(.dina(n11306), .dinb(n5084), .dout(n18807));
  jand g18693(.dina(n10836), .dinb(n5082), .dout(n18808));
  jand g18694(.dina(n10640), .dinb(n6050), .dout(n18809));
  jor  g18695(.dina(n18809), .dinb(n18808), .dout(n18810));
  jor  g18696(.dina(n18810), .dinb(n18807), .dout(n18811));
  jor  g18697(.dina(n18811), .dinb(n18806), .dout(n18812));
  jor  g18698(.dina(n18395), .dinb(n18391), .dout(n18813));
  jand g18699(.dina(n18403), .dinb(n18396), .dout(n18814));
  jnot g18700(.din(n18814), .dout(n18815));
  jand g18701(.dina(n18815), .dinb(n18813), .dout(n18816));
  jnot g18702(.din(n18816), .dout(n18817));
  jand g18703(.dina(n2452), .dinb(n1261), .dout(n18818));
  jand g18704(.dina(n6166), .dinb(n3980), .dout(n18819));
  jand g18705(.dina(n1934), .dinb(n1427), .dout(n18820));
  jand g18706(.dina(n18820), .dinb(n6335), .dout(n18821));
  jand g18707(.dina(n18821), .dinb(n9535), .dout(n18822));
  jand g18708(.dina(n18822), .dinb(n18819), .dout(n18823));
  jand g18709(.dina(n2106), .dinb(n452), .dout(n18824));
  jand g18710(.dina(n18824), .dinb(n1378), .dout(n18825));
  jand g18711(.dina(n9323), .dinb(n7648), .dout(n18826));
  jand g18712(.dina(n18826), .dinb(n499), .dout(n18827));
  jand g18713(.dina(n18827), .dinb(n1162), .dout(n18828));
  jand g18714(.dina(n18828), .dinb(n18825), .dout(n18829));
  jand g18715(.dina(n18829), .dinb(n18823), .dout(n18830));
  jand g18716(.dina(n18830), .dinb(n18818), .dout(n18831));
  jand g18717(.dina(n3011), .dinb(n2507), .dout(n18832));
  jand g18718(.dina(n18832), .dinb(n18831), .dout(n18833));
  jxor g18719(.dina(n18833), .dinb(n18391), .dout(n18834));
  jxor g18720(.dina(n18834), .dinb(n18817), .dout(n18835));
  jxor g18721(.dina(n18835), .dinb(n18812), .dout(n18836));
  jxor g18722(.dina(n18836), .dinb(n18805), .dout(n18837));
  jand g18723(.dina(n11800), .dinb(n2936), .dout(n18838));
  jand g18724(.dina(n11798), .dinb(n2943), .dout(n18839));
  jand g18725(.dina(n11646), .dinb(n2940), .dout(n18840));
  jand g18726(.dina(n11647), .dinb(n3684), .dout(n18841));
  jor  g18727(.dina(n18841), .dinb(n18840), .dout(n18842));
  jor  g18728(.dina(n18842), .dinb(n18839), .dout(n18843));
  jor  g18729(.dina(n18843), .dinb(n18838), .dout(n18844));
  jxor g18730(.dina(n18844), .dinb(n93), .dout(n18845));
  jxor g18731(.dina(n18845), .dinb(n18837), .dout(n18846));
  jand g18732(.dina(n12684), .dinb(n71), .dout(n18847));
  jand g18733(.dina(n12547), .dinb(n731), .dout(n18848));
  jand g18734(.dina(n12536), .dinb(n796), .dout(n18849));
  jor  g18735(.dina(n18849), .dinb(n18848), .dout(n18850));
  jand g18736(.dina(n12282), .dinb(n1806), .dout(n18851));
  jor  g18737(.dina(n18851), .dinb(n18850), .dout(n18852));
  jor  g18738(.dina(n18852), .dinb(n18847), .dout(n18853));
  jxor g18739(.dina(n18853), .dinb(n77), .dout(n18854));
  jxor g18740(.dina(n18854), .dinb(n18846), .dout(n18855));
  jxor g18741(.dina(n18855), .dinb(n18802), .dout(n18856));
  jand g18742(.dina(n13639), .dinb(n806), .dout(n18857));
  jand g18743(.dina(n13478), .dinb(n1620), .dout(n18858));
  jand g18744(.dina(n13248), .dinb(n1612), .dout(n18859));
  jand g18745(.dina(n12669), .dinb(n1644), .dout(n18860));
  jor  g18746(.dina(n18860), .dinb(n18859), .dout(n18861));
  jor  g18747(.dina(n18861), .dinb(n18858), .dout(n18862));
  jor  g18748(.dina(n18862), .dinb(n18857), .dout(n18863));
  jxor g18749(.dina(n18863), .dinb(n65), .dout(n18864));
  jxor g18750(.dina(n18864), .dinb(n18856), .dout(n18865));
  jxor g18751(.dina(n18865), .dinb(n18798), .dout(n18866));
  jand g18752(.dina(n14251), .dinb(n1819), .dout(n18867));
  jand g18753(.dina(n14249), .dinb(n2243), .dout(n18868));
  jand g18754(.dina(n13614), .dinb(n2180), .dout(n18869));
  jand g18755(.dina(n13469), .dinb(n2185), .dout(n18870));
  jor  g18756(.dina(n18870), .dinb(n18869), .dout(n18871));
  jor  g18757(.dina(n18871), .dinb(n18868), .dout(n18872));
  jor  g18758(.dina(n18872), .dinb(n18867), .dout(n18873));
  jxor g18759(.dina(n18873), .dinb(n2196), .dout(n18874));
  jxor g18760(.dina(n18874), .dinb(n18866), .dout(n18875));
  jxor g18761(.dina(n18875), .dinb(n18794), .dout(n18876));
  jand g18762(.dina(n14551), .dinb(n2743), .dout(n18877));
  jand g18763(.dina(n14549), .dinb(n2752), .dout(n18878));
  jand g18764(.dina(n14447), .dinb(n2748), .dout(n18879));
  jand g18765(.dina(n14448), .dinb(n2757), .dout(n18880));
  jor  g18766(.dina(n18880), .dinb(n18879), .dout(n18881));
  jor  g18767(.dina(n18881), .dinb(n18878), .dout(n18882));
  jor  g18768(.dina(n18882), .dinb(n18877), .dout(n18883));
  jxor g18769(.dina(n18883), .dinb(n2441), .dout(n18884));
  jxor g18770(.dina(n18884), .dinb(n18876), .dout(n18885));
  jxor g18771(.dina(n18885), .dinb(n18790), .dout(n18886));
  jnot g18772(.din(n18886), .dout(n18887));
  jand g18773(.dina(n15831), .dinb(n3423), .dout(n18888));
  jand g18774(.dina(n15567), .dinb(n3428), .dout(n18889));
  jand g18775(.dina(n15829), .dinb(n3569), .dout(n18890));
  jor  g18776(.dina(n18890), .dinb(n18889), .dout(n18891));
  jand g18777(.dina(n15315), .dinb(n3210), .dout(n18892));
  jor  g18778(.dina(n18892), .dinb(n18891), .dout(n18893));
  jor  g18779(.dina(n18893), .dinb(n18888), .dout(n18894));
  jxor g18780(.dina(n18894), .dinb(n3473), .dout(n18895));
  jxor g18781(.dina(n18895), .dinb(n18887), .dout(n18896));
  jxor g18782(.dina(n18896), .dinb(n18785), .dout(n18897));
  jand g18783(.dina(n16594), .dinb(n4022), .dout(n18898));
  jand g18784(.dina(n16343), .dinb(n4027), .dout(n18899));
  jand g18785(.dina(n16592), .dinb(n4220), .dout(n18900));
  jor  g18786(.dina(n18900), .dinb(n18899), .dout(n18901));
  jand g18787(.dina(n16082), .dinb(n3870), .dout(n18902));
  jor  g18788(.dina(n18902), .dinb(n18901), .dout(n18903));
  jor  g18789(.dina(n18903), .dinb(n18898), .dout(n18904));
  jxor g18790(.dina(n18904), .dinb(n4050), .dout(n18905));
  jxor g18791(.dina(n18905), .dinb(n18897), .dout(n18906));
  jxor g18792(.dina(n18906), .dinb(n18781), .dout(n18907));
  jxor g18793(.dina(n18907), .dinb(n18769), .dout(n18908));
  jxor g18794(.dina(n18476), .dinb(n18765), .dout(n18909));
  jxor g18795(.dina(n18485), .dinb(n18909), .dout(n18910));
  jor  g18796(.dina(n18910), .dinb(n18312), .dout(n18911));
  jor  g18797(.dina(n18487), .dinb(n18308), .dout(n18912));
  jand g18798(.dina(n18912), .dinb(n18911), .dout(n18913));
  jxor g18799(.dina(n18913), .dinb(n18908), .dout(n18914));
  jxor g18800(.dina(n18914), .dinb(n18488), .dout(n18915));
  jxor g18801(.dina(n18915), .dinb(n18764), .dout(n18916));
  jand g18802(.dina(n18916), .dinb(n2743), .dout(n18917));
  jand g18803(.dina(n18914), .dinb(n2752), .dout(n18918));
  jand g18804(.dina(n18488), .dinb(n2748), .dout(n18919));
  jand g18805(.dina(n18292), .dinb(n2757), .dout(n18920));
  jor  g18806(.dina(n18920), .dinb(n18919), .dout(n18921));
  jor  g18807(.dina(n18921), .dinb(n18918), .dout(n18922));
  jor  g18808(.dina(n18922), .dinb(n18917), .dout(n18923));
  jxor g18809(.dina(n18923), .dinb(n2441), .dout(n18924));
  jxor g18810(.dina(n18924), .dinb(n18761), .dout(n18925));
  jxor g18811(.dina(n18925), .dinb(n18700), .dout(n18926));
  jnot g18812(.din(n18926), .dout(n18927));
  jor  g18813(.dina(n18994), .dinb(n18773), .dout(n18928));
  jand g18814(.dina(n18906), .dinb(n18781), .dout(n18929));
  jnot g18815(.din(n18929), .dout(n18930));
  jand g18816(.dina(n18930), .dinb(n18928), .dout(n18931));
  jand g18817(.dina(n18885), .dinb(n18790), .dout(n18932));
  jnot g18818(.din(n18932), .dout(n18933));
  jor  g18819(.dina(n18895), .dinb(n18887), .dout(n18934));
  jand g18820(.dina(n18934), .dinb(n18933), .dout(n18935));
  jnot g18821(.din(n18794), .dout(n18936));
  jand g18822(.dina(n18875), .dinb(n18936), .dout(n18937));
  jnot g18823(.din(n18937), .dout(n18938));
  jor  g18824(.dina(n18884), .dinb(n18876), .dout(n18939));
  jand g18825(.dina(n18939), .dinb(n18938), .dout(n18940));
  jnot g18826(.din(n18798), .dout(n18941));
  jand g18827(.dina(n18865), .dinb(n18941), .dout(n18942));
  jnot g18828(.din(n18942), .dout(n18943));
  jor  g18829(.dina(n18874), .dinb(n18866), .dout(n18944));
  jand g18830(.dina(n18944), .dinb(n18943), .dout(n18945));
  jnot g18831(.din(n18802), .dout(n18946));
  jand g18832(.dina(n18855), .dinb(n18946), .dout(n18947));
  jnot g18833(.din(n18947), .dout(n18948));
  jor  g18834(.dina(n18864), .dinb(n18856), .dout(n18949));
  jand g18835(.dina(n18949), .dinb(n18948), .dout(n18950));
  jnot g18836(.din(n18837), .dout(n18951));
  jor  g18837(.dina(n18845), .dinb(n18951), .dout(n18952));
  jor  g18838(.dina(n18854), .dinb(n18846), .dout(n18953));
  jand g18839(.dina(n18953), .dinb(n18952), .dout(n18954));
  jand g18840(.dina(n18835), .dinb(n18812), .dout(n18955));
  jand g18841(.dina(n18836), .dinb(n18805), .dout(n18956));
  jor  g18842(.dina(n18956), .dinb(n18955), .dout(n18957));
  jand g18843(.dina(n11824), .dinb(n5076), .dout(n18958));
  jand g18844(.dina(n11647), .dinb(n5084), .dout(n18959));
  jand g18845(.dina(n11306), .dinb(n5082), .dout(n18960));
  jand g18846(.dina(n10836), .dinb(n6050), .dout(n18961));
  jor  g18847(.dina(n18961), .dinb(n18960), .dout(n18962));
  jor  g18848(.dina(n18962), .dinb(n18959), .dout(n18963));
  jor  g18849(.dina(n18963), .dinb(n18958), .dout(n18964));
  jnot g18850(.din(n18964), .dout(n18965));
  jor  g18851(.dina(n18833), .dinb(n18391), .dout(n18966));
  jand g18852(.dina(n18834), .dinb(n18817), .dout(n18967));
  jnot g18853(.din(n18967), .dout(n18968));
  jand g18854(.dina(n18968), .dinb(n18966), .dout(n18969));
  jand g18855(.dina(n1042), .dinb(n492), .dout(n18970));
  jand g18856(.dina(n18970), .dinb(n1846), .dout(n18971));
  jand g18857(.dina(n18971), .dinb(n4661), .dout(n18972));
  jand g18858(.dina(n18972), .dinb(n1213), .dout(n18973));
  jand g18859(.dina(n18973), .dinb(n521), .dout(n18974));
  jand g18860(.dina(n18974), .dinb(n15913), .dout(n18975));
  jand g18861(.dina(n978), .dinb(n1429), .dout(n18976));
  jand g18862(.dina(n18976), .dinb(n1366), .dout(n18977));
  jand g18863(.dina(n1159), .dinb(n325), .dout(n18978));
  jand g18864(.dina(n18978), .dinb(n9540), .dout(n18979));
  jand g18865(.dina(n18979), .dinb(n18977), .dout(n18980));
  jand g18866(.dina(n18980), .dinb(n1751), .dout(n18981));
  jand g18867(.dina(n2715), .dinb(n1957), .dout(n18982));
  jand g18868(.dina(n10400), .dinb(n7086), .dout(n18983));
  jand g18869(.dina(n2409), .dinb(n1432), .dout(n18984));
  jand g18870(.dina(n18984), .dinb(n18983), .dout(n18985));
  jand g18871(.dina(n18985), .dinb(n18982), .dout(n18986));
  jand g18872(.dina(n18986), .dinb(n18981), .dout(n18987));
  jand g18873(.dina(n18987), .dinb(n4004), .dout(n18988));
  jand g18874(.dina(n18988), .dinb(n14401), .dout(n18989));
  jand g18875(.dina(n18989), .dinb(n18975), .dout(n18990));
  jxor g18876(.dina(n18990), .dinb(n18390), .dout(n18991));
  jor  g18877(.dina(n4699), .dinb(n4690), .dout(n18992));
  jand g18878(.dina(n18992), .dinb(n16924), .dout(n18993));
  jxor g18879(.dina(n18993), .dinb(n4713), .dout(n18994));
  jxor g18880(.dina(n18994), .dinb(n18991), .dout(n18995));
  jxor g18881(.dina(n18995), .dinb(n18969), .dout(n18996));
  jxor g18882(.dina(n18996), .dinb(n18965), .dout(n18997));
  jand g18883(.dina(n12284), .dinb(n2936), .dout(n18998));
  jand g18884(.dina(n12282), .dinb(n2943), .dout(n18999));
  jand g18885(.dina(n11798), .dinb(n2940), .dout(n19000));
  jand g18886(.dina(n11646), .dinb(n3684), .dout(n19001));
  jor  g18887(.dina(n19001), .dinb(n19000), .dout(n19002));
  jor  g18888(.dina(n19002), .dinb(n18999), .dout(n19003));
  jor  g18889(.dina(n19003), .dinb(n18998), .dout(n19004));
  jxor g18890(.dina(n19004), .dinb(n93), .dout(n19005));
  jxor g18891(.dina(n19005), .dinb(n18997), .dout(n19006));
  jxor g18892(.dina(n19006), .dinb(n18957), .dout(n19007));
  jand g18893(.dina(n12671), .dinb(n71), .dout(n19008));
  jand g18894(.dina(n12669), .dinb(n796), .dout(n19009));
  jand g18895(.dina(n12536), .dinb(n731), .dout(n19010));
  jand g18896(.dina(n12547), .dinb(n1806), .dout(n19011));
  jor  g18897(.dina(n19011), .dinb(n19010), .dout(n19012));
  jor  g18898(.dina(n19012), .dinb(n19009), .dout(n19013));
  jor  g18899(.dina(n19013), .dinb(n19008), .dout(n19014));
  jxor g18900(.dina(n19014), .dinb(n77), .dout(n19015));
  jxor g18901(.dina(n19015), .dinb(n19007), .dout(n19016));
  jxor g18902(.dina(n19016), .dinb(n18954), .dout(n19017));
  jand g18903(.dina(n13627), .dinb(n806), .dout(n19018));
  jand g18904(.dina(n13478), .dinb(n1612), .dout(n19019));
  jand g18905(.dina(n13469), .dinb(n1620), .dout(n19020));
  jor  g18906(.dina(n19020), .dinb(n19019), .dout(n19021));
  jand g18907(.dina(n13248), .dinb(n1644), .dout(n19022));
  jor  g18908(.dina(n19022), .dinb(n19021), .dout(n19023));
  jor  g18909(.dina(n19023), .dinb(n19018), .dout(n19024));
  jxor g18910(.dina(n19024), .dinb(n65), .dout(n19025));
  jxor g18911(.dina(n19025), .dinb(n19017), .dout(n19026));
  jxor g18912(.dina(n19026), .dinb(n18950), .dout(n19027));
  jand g18913(.dina(n14579), .dinb(n1819), .dout(n19028));
  jand g18914(.dina(n14448), .dinb(n2243), .dout(n19029));
  jand g18915(.dina(n14249), .dinb(n2180), .dout(n19030));
  jand g18916(.dina(n13614), .dinb(n2185), .dout(n19031));
  jor  g18917(.dina(n19031), .dinb(n19030), .dout(n19032));
  jor  g18918(.dina(n19032), .dinb(n19029), .dout(n19033));
  jor  g18919(.dina(n19033), .dinb(n19028), .dout(n19034));
  jxor g18920(.dina(n19034), .dinb(n2196), .dout(n19035));
  jxor g18921(.dina(n19035), .dinb(n19027), .dout(n19036));
  jxor g18922(.dina(n19036), .dinb(n18945), .dout(n19037));
  jand g18923(.dina(n15317), .dinb(n2743), .dout(n19038));
  jand g18924(.dina(n14549), .dinb(n2748), .dout(n19039));
  jand g18925(.dina(n15315), .dinb(n2752), .dout(n19040));
  jor  g18926(.dina(n19040), .dinb(n19039), .dout(n19041));
  jand g18927(.dina(n14447), .dinb(n2757), .dout(n19042));
  jor  g18928(.dina(n19042), .dinb(n19041), .dout(n19043));
  jor  g18929(.dina(n19043), .dinb(n19038), .dout(n19044));
  jxor g18930(.dina(n19044), .dinb(n2441), .dout(n19045));
  jxor g18931(.dina(n19045), .dinb(n19037), .dout(n19046));
  jxor g18932(.dina(n19046), .dinb(n18940), .dout(n19047));
  jand g18933(.dina(n16084), .dinb(n3423), .dout(n19048));
  jand g18934(.dina(n15829), .dinb(n3428), .dout(n19049));
  jand g18935(.dina(n16082), .dinb(n3569), .dout(n19050));
  jor  g18936(.dina(n19050), .dinb(n19049), .dout(n19051));
  jand g18937(.dina(n15567), .dinb(n3210), .dout(n19052));
  jor  g18938(.dina(n19052), .dinb(n19051), .dout(n19053));
  jor  g18939(.dina(n19053), .dinb(n19048), .dout(n19054));
  jxor g18940(.dina(n19054), .dinb(n3473), .dout(n19055));
  jxor g18941(.dina(n19055), .dinb(n19047), .dout(n19056));
  jnot g18942(.din(n19056), .dout(n19057));
  jxor g18943(.dina(n19057), .dinb(n18935), .dout(n19058));
  jnot g18944(.din(n18896), .dout(n19059));
  jor  g18945(.dina(n19059), .dinb(n18785), .dout(n19060));
  jor  g18946(.dina(n18905), .dinb(n18897), .dout(n19061));
  jand g18947(.dina(n19061), .dinb(n19060), .dout(n19062));
  jand g18948(.dina(n16930), .dinb(n4022), .dout(n19063));
  jand g18949(.dina(n16592), .dinb(n4027), .dout(n19064));
  jand g18950(.dina(n16928), .dinb(n4220), .dout(n19065));
  jor  g18951(.dina(n19065), .dinb(n19064), .dout(n19066));
  jand g18952(.dina(n16343), .dinb(n3870), .dout(n19067));
  jor  g18953(.dina(n19067), .dinb(n19066), .dout(n19068));
  jor  g18954(.dina(n19068), .dinb(n19063), .dout(n19069));
  jxor g18955(.dina(n19069), .dinb(n4050), .dout(n19070));
  jxor g18956(.dina(n19070), .dinb(n19062), .dout(n19071));
  jxor g18957(.dina(n19071), .dinb(n19058), .dout(n19072));
  jnot g18958(.din(n19072), .dout(n19073));
  jor  g18959(.dina(n19073), .dinb(n18931), .dout(n19074));
  jnot g18960(.din(n18907), .dout(n19075));
  jor  g18961(.dina(n19075), .dinb(n18769), .dout(n19076));
  jor  g18962(.dina(n18913), .dinb(n18908), .dout(n19077));
  jand g18963(.dina(n19077), .dinb(n19076), .dout(n19078));
  jxor g18964(.dina(n19072), .dinb(n18931), .dout(n19079));
  jor  g18965(.dina(n19079), .dinb(n19078), .dout(n19080));
  jand g18966(.dina(n19080), .dinb(n19074), .dout(n19081));
  jor  g18967(.dina(n19070), .dinb(n19062), .dout(n19082));
  jnot g18968(.din(n19082), .dout(n19083));
  jand g18969(.dina(n19071), .dinb(n19058), .dout(n19084));
  jor  g18970(.dina(n19084), .dinb(n19083), .dout(n19085));
  jor  g18971(.dina(n19055), .dinb(n19047), .dout(n19086));
  jor  g18972(.dina(n19057), .dinb(n18935), .dout(n19087));
  jand g18973(.dina(n19087), .dinb(n19086), .dout(n19088));
  jor  g18974(.dina(n19045), .dinb(n19037), .dout(n19089));
  jnot g18975(.din(n19046), .dout(n19090));
  jor  g18976(.dina(n19090), .dinb(n18940), .dout(n19091));
  jand g18977(.dina(n19091), .dinb(n19089), .dout(n19092));
  jor  g18978(.dina(n19035), .dinb(n19027), .dout(n19093));
  jnot g18979(.din(n19036), .dout(n19094));
  jor  g18980(.dina(n19094), .dinb(n18945), .dout(n19095));
  jand g18981(.dina(n19095), .dinb(n19093), .dout(n19096));
  jor  g18982(.dina(n19025), .dinb(n19017), .dout(n19097));
  jnot g18983(.din(n19026), .dout(n19098));
  jor  g18984(.dina(n19098), .dinb(n18950), .dout(n19099));
  jand g18985(.dina(n19099), .dinb(n19097), .dout(n19100));
  jor  g18986(.dina(n19015), .dinb(n19007), .dout(n19101));
  jnot g18987(.din(n19016), .dout(n19102));
  jor  g18988(.dina(n19102), .dinb(n18954), .dout(n19103));
  jand g18989(.dina(n19103), .dinb(n19101), .dout(n19104));
  jnot g18990(.din(n18997), .dout(n19105));
  jor  g18991(.dina(n19005), .dinb(n19105), .dout(n19106));
  jnot g18992(.din(n18957), .dout(n19107));
  jor  g18993(.dina(n19006), .dinb(n19107), .dout(n19108));
  jand g18994(.dina(n19108), .dinb(n19106), .dout(n19109));
  jnot g18995(.din(n18969), .dout(n19110));
  jand g18996(.dina(n18995), .dinb(n19110), .dout(n19111));
  jnot g18997(.din(n19111), .dout(n19112));
  jor  g18998(.dina(n18996), .dinb(n18965), .dout(n19113));
  jand g18999(.dina(n19113), .dinb(n19112), .dout(n19114));
  jand g19000(.dina(n1716), .dinb(n982), .dout(n19115));
  jand g19001(.dina(n19115), .dinb(n5974), .dout(n19116));
  jand g19002(.dina(n15282), .dinb(n697), .dout(n19117));
  jand g19003(.dina(n19117), .dinb(n3782), .dout(n19118));
  jand g19004(.dina(n19118), .dinb(n17174), .dout(n19119));
  jand g19005(.dina(n19119), .dinb(n19116), .dout(n19120));
  jand g19006(.dina(n19120), .dinb(n1300), .dout(n19121));
  jand g19007(.dina(n1228), .dinb(n1534), .dout(n19122));
  jand g19008(.dina(n19122), .dinb(n964), .dout(n19123));
  jand g19009(.dina(n19123), .dinb(n2615), .dout(n19124));
  jand g19010(.dina(n19124), .dinb(n1245), .dout(n19125));
  jand g19011(.dina(n19125), .dinb(n18184), .dout(n19126));
  jand g19012(.dina(n1162), .dinb(n470), .dout(n19127));
  jand g19013(.dina(n19127), .dinb(n1304), .dout(n19128));
  jand g19014(.dina(n19128), .dinb(n1375), .dout(n19129));
  jand g19015(.dina(n19129), .dinb(n8610), .dout(n19130));
  jand g19016(.dina(n19130), .dinb(n19126), .dout(n19131));
  jand g19017(.dina(n19131), .dinb(n19121), .dout(n19132));
  jnot g19018(.din(n19132), .dout(n19133));
  jor  g19019(.dina(n18990), .dinb(n18390), .dout(n19134));
  jand g19020(.dina(n18994), .dinb(n18991), .dout(n19135));
  jnot g19021(.din(n19135), .dout(n19136));
  jand g19022(.dina(n19136), .dinb(n19134), .dout(n19137));
  jxor g19023(.dina(n19137), .dinb(n19133), .dout(n19138));
  jand g19024(.dina(n11812), .dinb(n5076), .dout(n19139));
  jand g19025(.dina(n11646), .dinb(n5084), .dout(n19140));
  jand g19026(.dina(n11306), .dinb(n6050), .dout(n19141));
  jand g19027(.dina(n11647), .dinb(n5082), .dout(n19142));
  jor  g19028(.dina(n19142), .dinb(n19141), .dout(n19143));
  jor  g19029(.dina(n19143), .dinb(n19140), .dout(n19144));
  jor  g19030(.dina(n19144), .dinb(n19139), .dout(n19145));
  jxor g19031(.dina(n19145), .dinb(n19138), .dout(n19146));
  jxor g19032(.dina(n19146), .dinb(n19114), .dout(n19147));
  jand g19033(.dina(n12696), .dinb(n2936), .dout(n19148));
  jand g19034(.dina(n12282), .dinb(n2940), .dout(n19149));
  jand g19035(.dina(n12547), .dinb(n2943), .dout(n19150));
  jor  g19036(.dina(n19150), .dinb(n19149), .dout(n19151));
  jand g19037(.dina(n11798), .dinb(n3684), .dout(n19152));
  jor  g19038(.dina(n19152), .dinb(n19151), .dout(n19153));
  jor  g19039(.dina(n19153), .dinb(n19148), .dout(n19154));
  jxor g19040(.dina(n19154), .dinb(n93), .dout(n19155));
  jxor g19041(.dina(n19155), .dinb(n19147), .dout(n19156));
  jxor g19042(.dina(n19156), .dinb(n19109), .dout(n19157));
  jand g19043(.dina(n13250), .dinb(n71), .dout(n19158));
  jand g19044(.dina(n13248), .dinb(n796), .dout(n19159));
  jand g19045(.dina(n12669), .dinb(n731), .dout(n19160));
  jand g19046(.dina(n12536), .dinb(n1806), .dout(n19161));
  jor  g19047(.dina(n19161), .dinb(n19160), .dout(n19162));
  jor  g19048(.dina(n19162), .dinb(n19159), .dout(n19163));
  jor  g19049(.dina(n19163), .dinb(n19158), .dout(n19164));
  jxor g19050(.dina(n19164), .dinb(n77), .dout(n19165));
  jxor g19051(.dina(n19165), .dinb(n19157), .dout(n19166));
  jxor g19052(.dina(n19166), .dinb(n19104), .dout(n19167));
  jand g19053(.dina(n13616), .dinb(n806), .dout(n19168));
  jand g19054(.dina(n13469), .dinb(n1612), .dout(n19169));
  jand g19055(.dina(n13614), .dinb(n1620), .dout(n19170));
  jor  g19056(.dina(n19170), .dinb(n19169), .dout(n19171));
  jand g19057(.dina(n13478), .dinb(n1644), .dout(n19172));
  jor  g19058(.dina(n19172), .dinb(n19171), .dout(n19173));
  jor  g19059(.dina(n19173), .dinb(n19168), .dout(n19174));
  jxor g19060(.dina(n19174), .dinb(n65), .dout(n19175));
  jxor g19061(.dina(n19175), .dinb(n19167), .dout(n19176));
  jxor g19062(.dina(n19176), .dinb(n19100), .dout(n19177));
  jand g19063(.dina(n14562), .dinb(n1819), .dout(n19178));
  jand g19064(.dina(n14447), .dinb(n2243), .dout(n19179));
  jand g19065(.dina(n14448), .dinb(n2180), .dout(n19180));
  jand g19066(.dina(n14249), .dinb(n2185), .dout(n19181));
  jor  g19067(.dina(n19181), .dinb(n19180), .dout(n19182));
  jor  g19068(.dina(n19182), .dinb(n19179), .dout(n19183));
  jor  g19069(.dina(n19183), .dinb(n19178), .dout(n19184));
  jxor g19070(.dina(n19184), .dinb(n2196), .dout(n19185));
  jxor g19071(.dina(n19185), .dinb(n19177), .dout(n19186));
  jxor g19072(.dina(n19186), .dinb(n19096), .dout(n19187));
  jand g19073(.dina(n15569), .dinb(n2743), .dout(n19188));
  jand g19074(.dina(n15567), .dinb(n2752), .dout(n19189));
  jand g19075(.dina(n15315), .dinb(n2748), .dout(n19190));
  jand g19076(.dina(n14549), .dinb(n2757), .dout(n19191));
  jor  g19077(.dina(n19191), .dinb(n19190), .dout(n19192));
  jor  g19078(.dina(n19192), .dinb(n19189), .dout(n19193));
  jor  g19079(.dina(n19193), .dinb(n19188), .dout(n19194));
  jxor g19080(.dina(n19194), .dinb(n2441), .dout(n19195));
  jxor g19081(.dina(n19195), .dinb(n19187), .dout(n19196));
  jxor g19082(.dina(n19196), .dinb(n19092), .dout(n19197));
  jand g19083(.dina(n16345), .dinb(n3423), .dout(n19198));
  jand g19084(.dina(n16343), .dinb(n3569), .dout(n19199));
  jand g19085(.dina(n16082), .dinb(n3428), .dout(n19200));
  jand g19086(.dina(n15829), .dinb(n3210), .dout(n19201));
  jor  g19087(.dina(n19201), .dinb(n19200), .dout(n19202));
  jor  g19088(.dina(n19202), .dinb(n19199), .dout(n19203));
  jor  g19089(.dina(n19203), .dinb(n19198), .dout(n19204));
  jxor g19090(.dina(n19204), .dinb(n3473), .dout(n19205));
  jxor g19091(.dina(n19205), .dinb(n19197), .dout(n19206));
  jxor g19092(.dina(n19206), .dinb(n19088), .dout(n19207));
  jand g19093(.dina(n17312), .dinb(n4022), .dout(n19208));
  jand g19094(.dina(n16928), .dinb(n4027), .dout(n19209));
  jand g19095(.dina(n16592), .dinb(n3870), .dout(n19210));
  jand g19096(.dina(n16924), .dinb(n4220), .dout(n19211));
  jor  g19097(.dina(n19211), .dinb(n19210), .dout(n19212));
  jor  g19098(.dina(n19212), .dinb(n19209), .dout(n19213));
  jor  g19099(.dina(n19213), .dinb(n19208), .dout(n19214));
  jxor g19100(.dina(n19214), .dinb(n4050), .dout(n19215));
  jxor g19101(.dina(n19215), .dinb(n19207), .dout(n19216));
  jxor g19102(.dina(n19216), .dinb(n19085), .dout(n19217));
  jnot g19103(.din(n19217), .dout(n19218));
  jxor g19104(.dina(n19218), .dinb(n19081), .dout(n19219));
  jxor g19105(.dina(n19079), .dinb(n19078), .dout(n19220));
  jand g19106(.dina(n19220), .dinb(n19219), .dout(n19221));
  jand g19107(.dina(n19220), .dinb(n18914), .dout(n19222));
  jand g19108(.dina(n18914), .dinb(n18488), .dout(n19223));
  jand g19109(.dina(n18915), .dinb(n18764), .dout(n19224));
  jor  g19110(.dina(n19224), .dinb(n19223), .dout(n19225));
  jxor g19111(.dina(n19220), .dinb(n18914), .dout(n19226));
  jand g19112(.dina(n19226), .dinb(n19225), .dout(n19227));
  jor  g19113(.dina(n19227), .dinb(n19222), .dout(n19228));
  jxor g19114(.dina(n19220), .dinb(n19219), .dout(n19229));
  jand g19115(.dina(n19229), .dinb(n19228), .dout(n19230));
  jor  g19116(.dina(n19230), .dinb(n19221), .dout(n19231));
  jnot g19117(.din(n19088), .dout(n19232));
  jand g19118(.dina(n19206), .dinb(n19232), .dout(n19233));
  jor  g19119(.dina(n19215), .dinb(n19207), .dout(n19234));
  jnot g19120(.din(n19234), .dout(n19235));
  jor  g19121(.dina(n19235), .dinb(n19233), .dout(n19236));
  jnot g19122(.din(n19092), .dout(n19237));
  jand g19123(.dina(n19196), .dinb(n19237), .dout(n19238));
  jnot g19124(.din(n19238), .dout(n19239));
  jor  g19125(.dina(n19205), .dinb(n19197), .dout(n19240));
  jand g19126(.dina(n19240), .dinb(n19239), .dout(n19241));
  jand g19127(.dina(n4028), .dinb(n4025), .dout(n19242));
  jxor g19128(.dina(n19849), .dinb(n19241), .dout(n19249));
  jnot g19129(.din(n19096), .dout(n19250));
  jand g19130(.dina(n19186), .dinb(n19250), .dout(n19251));
  jnot g19131(.din(n19251), .dout(n19252));
  jor  g19132(.dina(n19195), .dinb(n19187), .dout(n19253));
  jand g19133(.dina(n19253), .dinb(n19252), .dout(n19254));
  jnot g19134(.din(n19100), .dout(n19255));
  jand g19135(.dina(n19176), .dinb(n19255), .dout(n19256));
  jnot g19136(.din(n19256), .dout(n19257));
  jor  g19137(.dina(n19185), .dinb(n19177), .dout(n19258));
  jand g19138(.dina(n19258), .dinb(n19257), .dout(n19259));
  jnot g19139(.din(n19104), .dout(n19260));
  jand g19140(.dina(n19166), .dinb(n19260), .dout(n19261));
  jnot g19141(.din(n19261), .dout(n19262));
  jor  g19142(.dina(n19175), .dinb(n19167), .dout(n19263));
  jand g19143(.dina(n19263), .dinb(n19262), .dout(n19264));
  jnot g19144(.din(n19109), .dout(n19265));
  jand g19145(.dina(n19156), .dinb(n19265), .dout(n19266));
  jnot g19146(.din(n19266), .dout(n19267));
  jor  g19147(.dina(n19165), .dinb(n19157), .dout(n19268));
  jand g19148(.dina(n19268), .dinb(n19267), .dout(n19269));
  jnot g19149(.din(n19114), .dout(n19270));
  jand g19150(.dina(n19146), .dinb(n19270), .dout(n19271));
  jnot g19151(.din(n19271), .dout(n19272));
  jor  g19152(.dina(n19155), .dinb(n19147), .dout(n19273));
  jand g19153(.dina(n19273), .dinb(n19272), .dout(n19274));
  jand g19154(.dina(n11800), .dinb(n5076), .dout(n19275));
  jand g19155(.dina(n11798), .dinb(n5084), .dout(n19276));
  jand g19156(.dina(n11646), .dinb(n5082), .dout(n19277));
  jand g19157(.dina(n11647), .dinb(n6050), .dout(n19278));
  jor  g19158(.dina(n19278), .dinb(n19277), .dout(n19279));
  jor  g19159(.dina(n19279), .dinb(n19276), .dout(n19280));
  jor  g19160(.dina(n19280), .dinb(n19275), .dout(n19281));
  jor  g19161(.dina(n19137), .dinb(n19133), .dout(n19282));
  jand g19162(.dina(n19145), .dinb(n19138), .dout(n19283));
  jnot g19163(.din(n19283), .dout(n19284));
  jand g19164(.dina(n19284), .dinb(n19282), .dout(n19285));
  jnot g19165(.din(n19285), .dout(n19286));
  jand g19166(.dina(n3266), .dinb(n1168), .dout(n19287));
  jand g19167(.dina(n691), .dinb(n1226), .dout(n19288));
  jand g19168(.dina(n19288), .dinb(n1289), .dout(n19289));
  jand g19169(.dina(n4641), .dinb(n3897), .dout(n19290));
  jand g19170(.dina(n19290), .dinb(n19289), .dout(n19291));
  jand g19171(.dina(n19291), .dinb(n19287), .dout(n19292));
  jand g19172(.dina(n1753), .dinb(n639), .dout(n19293));
  jand g19173(.dina(n1495), .dinb(n499), .dout(n19294));
  jand g19174(.dina(n19294), .dinb(n562), .dout(n19295));
  jand g19175(.dina(n7242), .dinb(n1961), .dout(n19296));
  jand g19176(.dina(n19296), .dinb(n19295), .dout(n19297));
  jand g19177(.dina(n19297), .dinb(n19293), .dout(n19298));
  jand g19178(.dina(n19298), .dinb(n15671), .dout(n19299));
  jand g19179(.dina(n19299), .dinb(n19292), .dout(n19300));
  jand g19180(.dina(n19300), .dinb(n11720), .dout(n19301));
  jand g19181(.dina(n19301), .dinb(n15108), .dout(n19302));
  jxor g19182(.dina(n19302), .dinb(n19133), .dout(n19303));
  jxor g19183(.dina(n19303), .dinb(n19286), .dout(n19304));
  jxor g19184(.dina(n19304), .dinb(n19281), .dout(n19305));
  jnot g19185(.din(n19305), .dout(n19306));
  jand g19186(.dina(n12684), .dinb(n2936), .dout(n19307));
  jand g19187(.dina(n12547), .dinb(n2940), .dout(n19308));
  jand g19188(.dina(n12536), .dinb(n2943), .dout(n19309));
  jor  g19189(.dina(n19309), .dinb(n19308), .dout(n19310));
  jand g19190(.dina(n12282), .dinb(n3684), .dout(n19311));
  jor  g19191(.dina(n19311), .dinb(n19310), .dout(n19312));
  jor  g19192(.dina(n19312), .dinb(n19307), .dout(n19313));
  jxor g19193(.dina(n19313), .dinb(n93), .dout(n19314));
  jxor g19194(.dina(n19314), .dinb(n19306), .dout(n19315));
  jxor g19195(.dina(n19315), .dinb(n19274), .dout(n19316));
  jand g19196(.dina(n13639), .dinb(n71), .dout(n19317));
  jand g19197(.dina(n13478), .dinb(n796), .dout(n19318));
  jand g19198(.dina(n13248), .dinb(n731), .dout(n19319));
  jand g19199(.dina(n12669), .dinb(n1806), .dout(n19320));
  jor  g19200(.dina(n19320), .dinb(n19319), .dout(n19321));
  jor  g19201(.dina(n19321), .dinb(n19318), .dout(n19322));
  jor  g19202(.dina(n19322), .dinb(n19317), .dout(n19323));
  jxor g19203(.dina(n19323), .dinb(n77), .dout(n19324));
  jxor g19204(.dina(n19324), .dinb(n19316), .dout(n19325));
  jxor g19205(.dina(n19325), .dinb(n19269), .dout(n19326));
  jand g19206(.dina(n14251), .dinb(n806), .dout(n19327));
  jand g19207(.dina(n13614), .dinb(n1612), .dout(n19328));
  jand g19208(.dina(n14249), .dinb(n1620), .dout(n19329));
  jor  g19209(.dina(n19329), .dinb(n19328), .dout(n19330));
  jand g19210(.dina(n13469), .dinb(n1644), .dout(n19331));
  jor  g19211(.dina(n19331), .dinb(n19330), .dout(n19332));
  jor  g19212(.dina(n19332), .dinb(n19327), .dout(n19333));
  jxor g19213(.dina(n19333), .dinb(n65), .dout(n19334));
  jxor g19214(.dina(n19334), .dinb(n19326), .dout(n19335));
  jxor g19215(.dina(n19335), .dinb(n19264), .dout(n19336));
  jand g19216(.dina(n14551), .dinb(n1819), .dout(n19337));
  jand g19217(.dina(n14447), .dinb(n2180), .dout(n19338));
  jand g19218(.dina(n14549), .dinb(n2243), .dout(n19339));
  jor  g19219(.dina(n19339), .dinb(n19338), .dout(n19340));
  jand g19220(.dina(n14448), .dinb(n2185), .dout(n19341));
  jor  g19221(.dina(n19341), .dinb(n19340), .dout(n19342));
  jor  g19222(.dina(n19342), .dinb(n19337), .dout(n19343));
  jxor g19223(.dina(n19343), .dinb(n2196), .dout(n19344));
  jxor g19224(.dina(n19344), .dinb(n19336), .dout(n19345));
  jxor g19225(.dina(n19345), .dinb(n19259), .dout(n19346));
  jand g19226(.dina(n15831), .dinb(n2743), .dout(n19347));
  jand g19227(.dina(n15567), .dinb(n2748), .dout(n19348));
  jand g19228(.dina(n15829), .dinb(n2752), .dout(n19349));
  jor  g19229(.dina(n19349), .dinb(n19348), .dout(n19350));
  jand g19230(.dina(n15315), .dinb(n2757), .dout(n19351));
  jor  g19231(.dina(n19351), .dinb(n19350), .dout(n19352));
  jor  g19232(.dina(n19352), .dinb(n19347), .dout(n19353));
  jxor g19233(.dina(n19353), .dinb(n2441), .dout(n19354));
  jxor g19234(.dina(n19354), .dinb(n19346), .dout(n19355));
  jxor g19235(.dina(n19355), .dinb(n19254), .dout(n19356));
  jand g19236(.dina(n16594), .dinb(n3423), .dout(n19357));
  jand g19237(.dina(n16592), .dinb(n3569), .dout(n19358));
  jand g19238(.dina(n16343), .dinb(n3428), .dout(n19359));
  jand g19239(.dina(n16082), .dinb(n3210), .dout(n19360));
  jor  g19240(.dina(n19360), .dinb(n19359), .dout(n19361));
  jor  g19241(.dina(n19361), .dinb(n19358), .dout(n19362));
  jor  g19242(.dina(n19362), .dinb(n19357), .dout(n19363));
  jxor g19243(.dina(n19363), .dinb(n3473), .dout(n19364));
  jxor g19244(.dina(n19364), .dinb(n19356), .dout(n19365));
  jxor g19245(.dina(n19365), .dinb(n19249), .dout(n19366));
  jxor g19246(.dina(n19366), .dinb(n19236), .dout(n19367));
  jnot g19247(.din(n19367), .dout(n19368));
  jand g19248(.dina(n19216), .dinb(n19085), .dout(n19369));
  jnot g19249(.din(n19369), .dout(n19370));
  jor  g19250(.dina(n19218), .dinb(n19081), .dout(n19371));
  jand g19251(.dina(n19371), .dinb(n19370), .dout(n19372));
  jxor g19252(.dina(n19372), .dinb(n19368), .dout(n19373));
  jxor g19253(.dina(n19373), .dinb(n19219), .dout(n19374));
  jxor g19254(.dina(n19374), .dinb(n19231), .dout(n19375));
  jand g19255(.dina(n19375), .dinb(n3423), .dout(n19376));
  jand g19256(.dina(n19219), .dinb(n3428), .dout(n19377));
  jand g19257(.dina(n19373), .dinb(n3569), .dout(n19378));
  jor  g19258(.dina(n19378), .dinb(n19377), .dout(n19379));
  jand g19259(.dina(n19220), .dinb(n3210), .dout(n19380));
  jor  g19260(.dina(n19380), .dinb(n19379), .dout(n19381));
  jor  g19261(.dina(n19381), .dinb(n19376), .dout(n19382));
  jxor g19262(.dina(n19382), .dinb(n3473), .dout(n19383));
  jor  g19263(.dina(n19383), .dinb(n18927), .dout(n19384));
  jxor g19264(.dina(n18696), .dinb(n18695), .dout(n19385));
  jnot g19265(.din(n19385), .dout(n19386));
  jxor g19266(.dina(n19229), .dinb(n19228), .dout(n19387));
  jand g19267(.dina(n19387), .dinb(n3423), .dout(n19388));
  jand g19268(.dina(n19219), .dinb(n3569), .dout(n19389));
  jand g19269(.dina(n19220), .dinb(n3428), .dout(n19390));
  jand g19270(.dina(n18914), .dinb(n3210), .dout(n19391));
  jor  g19271(.dina(n19391), .dinb(n19390), .dout(n19392));
  jor  g19272(.dina(n19392), .dinb(n19389), .dout(n19393));
  jor  g19273(.dina(n19393), .dinb(n19388), .dout(n19394));
  jxor g19274(.dina(n19394), .dinb(n3473), .dout(n19395));
  jor  g19275(.dina(n19395), .dinb(n19386), .dout(n19396));
  jxor g19276(.dina(n18691), .dinb(n18690), .dout(n19397));
  jnot g19277(.din(n19397), .dout(n19398));
  jxor g19278(.dina(n19226), .dinb(n19225), .dout(n19399));
  jand g19279(.dina(n19399), .dinb(n3423), .dout(n19400));
  jand g19280(.dina(n18914), .dinb(n3428), .dout(n19401));
  jand g19281(.dina(n19220), .dinb(n3569), .dout(n19402));
  jor  g19282(.dina(n19402), .dinb(n19401), .dout(n19403));
  jand g19283(.dina(n18488), .dinb(n3210), .dout(n19404));
  jor  g19284(.dina(n19404), .dinb(n19403), .dout(n19405));
  jor  g19285(.dina(n19405), .dinb(n19400), .dout(n19406));
  jxor g19286(.dina(n19406), .dinb(n3473), .dout(n19407));
  jor  g19287(.dina(n19407), .dinb(n19398), .dout(n19408));
  jxor g19288(.dina(n18686), .dinb(n18685), .dout(n19409));
  jnot g19289(.din(n19409), .dout(n19410));
  jand g19290(.dina(n18916), .dinb(n3423), .dout(n19411));
  jand g19291(.dina(n18914), .dinb(n3569), .dout(n19412));
  jand g19292(.dina(n18488), .dinb(n3428), .dout(n19413));
  jand g19293(.dina(n18292), .dinb(n3210), .dout(n19414));
  jor  g19294(.dina(n19414), .dinb(n19413), .dout(n19415));
  jor  g19295(.dina(n19415), .dinb(n19412), .dout(n19416));
  jor  g19296(.dina(n19416), .dinb(n19411), .dout(n19417));
  jxor g19297(.dina(n19417), .dinb(n3473), .dout(n19418));
  jor  g19298(.dina(n19418), .dinb(n19410), .dout(n19419));
  jxor g19299(.dina(n18681), .dinb(n18680), .dout(n19420));
  jnot g19300(.din(n19420), .dout(n19421));
  jand g19301(.dina(n18490), .dinb(n3423), .dout(n19422));
  jand g19302(.dina(n18292), .dinb(n3428), .dout(n19423));
  jand g19303(.dina(n18488), .dinb(n3569), .dout(n19424));
  jor  g19304(.dina(n19424), .dinb(n19423), .dout(n19425));
  jand g19305(.dina(n18293), .dinb(n3210), .dout(n19426));
  jor  g19306(.dina(n19426), .dinb(n19425), .dout(n19427));
  jor  g19307(.dina(n19427), .dinb(n19422), .dout(n19428));
  jxor g19308(.dina(n19428), .dinb(n3473), .dout(n19429));
  jor  g19309(.dina(n19429), .dinb(n19421), .dout(n19430));
  jxor g19310(.dina(n18676), .dinb(n18675), .dout(n19431));
  jand g19311(.dina(n18502), .dinb(n3423), .dout(n19432));
  jand g19312(.dina(n18292), .dinb(n3569), .dout(n19433));
  jand g19313(.dina(n18293), .dinb(n3428), .dout(n19434));
  jand g19314(.dina(n17942), .dinb(n3210), .dout(n19435));
  jor  g19315(.dina(n19435), .dinb(n19434), .dout(n19436));
  jor  g19316(.dina(n19436), .dinb(n19433), .dout(n19437));
  jor  g19317(.dina(n19437), .dinb(n19432), .dout(n19438));
  jxor g19318(.dina(n19438), .dinb(\a[14] ), .dout(n19439));
  jand g19319(.dina(n19439), .dinb(n19431), .dout(n19440));
  jxor g19320(.dina(n18671), .dinb(n18670), .dout(n19441));
  jnot g19321(.din(n19441), .dout(n19442));
  jand g19322(.dina(n18514), .dinb(n3423), .dout(n19443));
  jand g19323(.dina(n18293), .dinb(n3569), .dout(n19444));
  jand g19324(.dina(n17942), .dinb(n3428), .dout(n19445));
  jand g19325(.dina(n17535), .dinb(n3210), .dout(n19446));
  jor  g19326(.dina(n19446), .dinb(n19445), .dout(n19447));
  jor  g19327(.dina(n19447), .dinb(n19444), .dout(n19448));
  jor  g19328(.dina(n19448), .dinb(n19443), .dout(n19449));
  jxor g19329(.dina(n19449), .dinb(n3473), .dout(n19450));
  jor  g19330(.dina(n19450), .dinb(n19442), .dout(n19451));
  jxor g19331(.dina(n18666), .dinb(n18665), .dout(n19452));
  jnot g19332(.din(n19452), .dout(n19453));
  jand g19333(.dina(n17944), .dinb(n3423), .dout(n19454));
  jand g19334(.dina(n17535), .dinb(n3428), .dout(n19455));
  jand g19335(.dina(n17942), .dinb(n3569), .dout(n19456));
  jor  g19336(.dina(n19456), .dinb(n19455), .dout(n19457));
  jand g19337(.dina(n17329), .dinb(n3210), .dout(n19458));
  jor  g19338(.dina(n19458), .dinb(n19457), .dout(n19459));
  jor  g19339(.dina(n19459), .dinb(n19454), .dout(n19460));
  jxor g19340(.dina(n19460), .dinb(n3473), .dout(n19461));
  jor  g19341(.dina(n19461), .dinb(n19453), .dout(n19462));
  jxor g19342(.dina(n18661), .dinb(n18660), .dout(n19463));
  jnot g19343(.din(n19463), .dout(n19464));
  jand g19344(.dina(n17537), .dinb(n3423), .dout(n19465));
  jand g19345(.dina(n17329), .dinb(n3428), .dout(n19466));
  jand g19346(.dina(n17535), .dinb(n3569), .dout(n19467));
  jor  g19347(.dina(n19467), .dinb(n19466), .dout(n19468));
  jand g19348(.dina(n17330), .dinb(n3210), .dout(n19469));
  jor  g19349(.dina(n19469), .dinb(n19468), .dout(n19470));
  jor  g19350(.dina(n19470), .dinb(n19465), .dout(n19471));
  jxor g19351(.dina(n19471), .dinb(n3473), .dout(n19472));
  jor  g19352(.dina(n19472), .dinb(n19464), .dout(n19473));
  jxor g19353(.dina(n18656), .dinb(n18655), .dout(n19474));
  jnot g19354(.din(n19474), .dout(n19475));
  jand g19355(.dina(n17549), .dinb(n3423), .dout(n19476));
  jand g19356(.dina(n17329), .dinb(n3569), .dout(n19477));
  jand g19357(.dina(n17330), .dinb(n3428), .dout(n19478));
  jand g19358(.dina(n16940), .dinb(n3210), .dout(n19479));
  jor  g19359(.dina(n19479), .dinb(n19478), .dout(n19480));
  jor  g19360(.dina(n19480), .dinb(n19477), .dout(n19481));
  jor  g19361(.dina(n19481), .dinb(n19476), .dout(n19482));
  jxor g19362(.dina(n19482), .dinb(n3473), .dout(n19483));
  jor  g19363(.dina(n19483), .dinb(n19475), .dout(n19484));
  jxor g19364(.dina(n18653), .dinb(n18652), .dout(n19485));
  jnot g19365(.din(n19485), .dout(n19486));
  jand g19366(.dina(n17561), .dinb(n3423), .dout(n19487));
  jand g19367(.dina(n16940), .dinb(n3428), .dout(n19488));
  jand g19368(.dina(n17330), .dinb(n3569), .dout(n19489));
  jor  g19369(.dina(n19489), .dinb(n19488), .dout(n19490));
  jand g19370(.dina(n16604), .dinb(n3210), .dout(n19491));
  jor  g19371(.dina(n19491), .dinb(n19490), .dout(n19492));
  jor  g19372(.dina(n19492), .dinb(n19487), .dout(n19493));
  jxor g19373(.dina(n19493), .dinb(n3473), .dout(n19494));
  jor  g19374(.dina(n19494), .dinb(n19486), .dout(n19495));
  jxor g19375(.dina(n18648), .dinb(n18647), .dout(n19496));
  jnot g19376(.din(n19496), .dout(n19497));
  jand g19377(.dina(n16942), .dinb(n3423), .dout(n19498));
  jand g19378(.dina(n16940), .dinb(n3569), .dout(n19499));
  jand g19379(.dina(n16604), .dinb(n3428), .dout(n19500));
  jand g19380(.dina(n16355), .dinb(n3210), .dout(n19501));
  jor  g19381(.dina(n19501), .dinb(n19500), .dout(n19502));
  jor  g19382(.dina(n19502), .dinb(n19499), .dout(n19503));
  jor  g19383(.dina(n19503), .dinb(n19498), .dout(n19504));
  jxor g19384(.dina(n19504), .dinb(n3473), .dout(n19505));
  jor  g19385(.dina(n19505), .dinb(n19497), .dout(n19506));
  jxor g19386(.dina(n18644), .dinb(n18636), .dout(n19507));
  jnot g19387(.din(n19507), .dout(n19508));
  jand g19388(.dina(n16606), .dinb(n3423), .dout(n19509));
  jand g19389(.dina(n16604), .dinb(n3569), .dout(n19510));
  jand g19390(.dina(n16355), .dinb(n3428), .dout(n19511));
  jand g19391(.dina(n16360), .dinb(n3210), .dout(n19512));
  jor  g19392(.dina(n19512), .dinb(n19511), .dout(n19513));
  jor  g19393(.dina(n19513), .dinb(n19510), .dout(n19514));
  jor  g19394(.dina(n19514), .dinb(n19509), .dout(n19515));
  jxor g19395(.dina(n19515), .dinb(n3473), .dout(n19516));
  jor  g19396(.dina(n19516), .dinb(n19508), .dout(n19517));
  jand g19397(.dina(n16616), .dinb(n3423), .dout(n19518));
  jand g19398(.dina(n16355), .dinb(n3569), .dout(n19519));
  jand g19399(.dina(n16360), .dinb(n3428), .dout(n19520));
  jand g19400(.dina(n15841), .dinb(n3210), .dout(n19521));
  jor  g19401(.dina(n19521), .dinb(n19520), .dout(n19522));
  jor  g19402(.dina(n19522), .dinb(n19519), .dout(n19523));
  jor  g19403(.dina(n19523), .dinb(n19518), .dout(n19524));
  jxor g19404(.dina(n19524), .dinb(n3473), .dout(n19525));
  jnot g19405(.din(n19525), .dout(n19526));
  jor  g19406(.dina(n18623), .dinb(n2441), .dout(n19527));
  jxor g19407(.dina(n19527), .dinb(n18631), .dout(n19528));
  jand g19408(.dina(n19528), .dinb(n19526), .dout(n19529));
  jand g19409(.dina(n18620), .dinb(\a[17] ), .dout(n19530));
  jxor g19410(.dina(n19530), .dinb(n18618), .dout(n19531));
  jnot g19411(.din(n19531), .dout(n19532));
  jand g19412(.dina(n16632), .dinb(n3423), .dout(n19533));
  jand g19413(.dina(n16360), .dinb(n3569), .dout(n19534));
  jand g19414(.dina(n15841), .dinb(n3428), .dout(n19535));
  jand g19415(.dina(n15579), .dinb(n3210), .dout(n19536));
  jor  g19416(.dina(n19536), .dinb(n19535), .dout(n19537));
  jor  g19417(.dina(n19537), .dinb(n19534), .dout(n19538));
  jor  g19418(.dina(n19538), .dinb(n19533), .dout(n19539));
  jxor g19419(.dina(n19539), .dinb(n3473), .dout(n19540));
  jor  g19420(.dina(n19540), .dinb(n19532), .dout(n19541));
  jand g19421(.dina(n15329), .dinb(n3423), .dout(n19542));
  jand g19422(.dina(n15020), .dinb(n3428), .dout(n19543));
  jand g19423(.dina(n15327), .dinb(n3569), .dout(n19544));
  jor  g19424(.dina(n19544), .dinb(n19543), .dout(n19545));
  jor  g19425(.dina(n19545), .dinb(n19542), .dout(n19546));
  jnot g19426(.din(n19546), .dout(n19547));
  jand g19427(.dina(n15020), .dinb(n3205), .dout(n19548));
  jnot g19428(.din(n19548), .dout(n19549));
  jand g19429(.dina(n19549), .dinb(\a[14] ), .dout(n19550));
  jand g19430(.dina(n19550), .dinb(n19547), .dout(n19551));
  jand g19431(.dina(n15580), .dinb(n3423), .dout(n19552));
  jand g19432(.dina(n15327), .dinb(n3428), .dout(n19553));
  jor  g19433(.dina(n19553), .dinb(n19552), .dout(n19554));
  jand g19434(.dina(n15579), .dinb(n3569), .dout(n19555));
  jand g19435(.dina(n15020), .dinb(n3210), .dout(n19556));
  jor  g19436(.dina(n19556), .dinb(n19555), .dout(n19557));
  jor  g19437(.dina(n19557), .dinb(n19554), .dout(n19558));
  jnot g19438(.din(n19558), .dout(n19559));
  jand g19439(.dina(n19559), .dinb(n19551), .dout(n19560));
  jand g19440(.dina(n19560), .dinb(n18620), .dout(n19561));
  jnot g19441(.din(n19561), .dout(n19562));
  jxor g19442(.dina(n19560), .dinb(n18620), .dout(n19563));
  jnot g19443(.din(n19563), .dout(n19564));
  jand g19444(.dina(n15848), .dinb(n3423), .dout(n19565));
  jand g19445(.dina(n15841), .dinb(n3569), .dout(n19566));
  jand g19446(.dina(n15579), .dinb(n3428), .dout(n19567));
  jand g19447(.dina(n15327), .dinb(n3210), .dout(n19568));
  jor  g19448(.dina(n19568), .dinb(n19567), .dout(n19569));
  jor  g19449(.dina(n19569), .dinb(n19566), .dout(n19570));
  jor  g19450(.dina(n19570), .dinb(n19565), .dout(n19571));
  jxor g19451(.dina(n19571), .dinb(n3473), .dout(n19572));
  jor  g19452(.dina(n19572), .dinb(n19564), .dout(n19573));
  jand g19453(.dina(n19573), .dinb(n19562), .dout(n19574));
  jnot g19454(.din(n19574), .dout(n19575));
  jxor g19455(.dina(n19540), .dinb(n19532), .dout(n19576));
  jand g19456(.dina(n19576), .dinb(n19575), .dout(n19577));
  jnot g19457(.din(n19577), .dout(n19578));
  jand g19458(.dina(n19578), .dinb(n19541), .dout(n19579));
  jnot g19459(.din(n19579), .dout(n19580));
  jxor g19460(.dina(n19528), .dinb(n19526), .dout(n19581));
  jand g19461(.dina(n19581), .dinb(n19580), .dout(n19582));
  jor  g19462(.dina(n19582), .dinb(n19529), .dout(n19583));
  jxor g19463(.dina(n19516), .dinb(n19508), .dout(n19584));
  jand g19464(.dina(n19584), .dinb(n19583), .dout(n19585));
  jnot g19465(.din(n19585), .dout(n19586));
  jand g19466(.dina(n19586), .dinb(n19517), .dout(n19587));
  jnot g19467(.din(n19587), .dout(n19588));
  jxor g19468(.dina(n19505), .dinb(n19497), .dout(n19589));
  jand g19469(.dina(n19589), .dinb(n19588), .dout(n19590));
  jnot g19470(.din(n19590), .dout(n19591));
  jand g19471(.dina(n19591), .dinb(n19506), .dout(n19592));
  jnot g19472(.din(n19592), .dout(n19593));
  jxor g19473(.dina(n19494), .dinb(n19486), .dout(n19594));
  jand g19474(.dina(n19594), .dinb(n19593), .dout(n19595));
  jnot g19475(.din(n19595), .dout(n19596));
  jand g19476(.dina(n19596), .dinb(n19495), .dout(n19597));
  jnot g19477(.din(n19597), .dout(n19598));
  jxor g19478(.dina(n19483), .dinb(n19475), .dout(n19599));
  jand g19479(.dina(n19599), .dinb(n19598), .dout(n19600));
  jnot g19480(.din(n19600), .dout(n19601));
  jand g19481(.dina(n19601), .dinb(n19484), .dout(n19602));
  jnot g19482(.din(n19602), .dout(n19603));
  jxor g19483(.dina(n19472), .dinb(n19464), .dout(n19604));
  jand g19484(.dina(n19604), .dinb(n19603), .dout(n19605));
  jnot g19485(.din(n19605), .dout(n19606));
  jand g19486(.dina(n19606), .dinb(n19473), .dout(n19607));
  jnot g19487(.din(n19607), .dout(n19608));
  jxor g19488(.dina(n19461), .dinb(n19453), .dout(n19609));
  jand g19489(.dina(n19609), .dinb(n19608), .dout(n19610));
  jnot g19490(.din(n19610), .dout(n19611));
  jand g19491(.dina(n19611), .dinb(n19462), .dout(n19612));
  jnot g19492(.din(n19612), .dout(n19613));
  jxor g19493(.dina(n19450), .dinb(n19442), .dout(n19614));
  jand g19494(.dina(n19614), .dinb(n19613), .dout(n19615));
  jnot g19495(.din(n19615), .dout(n19616));
  jand g19496(.dina(n19616), .dinb(n19451), .dout(n19617));
  jnot g19497(.din(n19617), .dout(n19618));
  jxor g19498(.dina(n19439), .dinb(n19431), .dout(n19619));
  jand g19499(.dina(n19619), .dinb(n19618), .dout(n19620));
  jor  g19500(.dina(n19620), .dinb(n19440), .dout(n19621));
  jxor g19501(.dina(n19429), .dinb(n19421), .dout(n19622));
  jand g19502(.dina(n19622), .dinb(n19621), .dout(n19623));
  jnot g19503(.din(n19623), .dout(n19624));
  jand g19504(.dina(n19624), .dinb(n19430), .dout(n19625));
  jnot g19505(.din(n19625), .dout(n19626));
  jxor g19506(.dina(n19418), .dinb(n19410), .dout(n19627));
  jand g19507(.dina(n19627), .dinb(n19626), .dout(n19628));
  jnot g19508(.din(n19628), .dout(n19629));
  jand g19509(.dina(n19629), .dinb(n19419), .dout(n19630));
  jnot g19510(.din(n19630), .dout(n19631));
  jxor g19511(.dina(n19407), .dinb(n19398), .dout(n19632));
  jand g19512(.dina(n19632), .dinb(n19631), .dout(n19633));
  jnot g19513(.din(n19633), .dout(n19634));
  jand g19514(.dina(n19634), .dinb(n19408), .dout(n19635));
  jnot g19515(.din(n19635), .dout(n19636));
  jxor g19516(.dina(n19395), .dinb(n19386), .dout(n19637));
  jand g19517(.dina(n19637), .dinb(n19636), .dout(n19638));
  jnot g19518(.din(n19638), .dout(n19639));
  jand g19519(.dina(n19639), .dinb(n19396), .dout(n19640));
  jnot g19520(.din(n19640), .dout(n19641));
  jxor g19521(.dina(n19383), .dinb(n18927), .dout(n19642));
  jand g19522(.dina(n19642), .dinb(n19641), .dout(n19643));
  jnot g19523(.din(n19643), .dout(n19644));
  jand g19524(.dina(n19644), .dinb(n19384), .dout(n19645));
  jnot g19525(.din(n19645), .dout(n19646));
  jor  g19526(.dina(n18924), .dinb(n18761), .dout(n19647));
  jand g19527(.dina(n18925), .dinb(n18700), .dout(n19648));
  jnot g19528(.din(n19648), .dout(n19649));
  jand g19529(.dina(n19649), .dinb(n19647), .dout(n19650));
  jnot g19530(.din(n19650), .dout(n19651));
  jor  g19531(.dina(n18758), .dinb(n18750), .dout(n19652));
  jand g19532(.dina(n18759), .dinb(n18705), .dout(n19653));
  jnot g19533(.din(n19653), .dout(n19654));
  jand g19534(.dina(n19654), .dinb(n19652), .dout(n19655));
  jnot g19535(.din(n19655), .dout(n19656));
  jor  g19536(.dina(n18747), .dinb(n18739), .dout(n19657));
  jand g19537(.dina(n18748), .dinb(n18710), .dout(n19658));
  jnot g19538(.din(n19658), .dout(n19659));
  jand g19539(.dina(n19659), .dinb(n19657), .dout(n19660));
  jnot g19540(.din(n19660), .dout(n19661));
  jor  g19541(.dina(n18736), .dinb(n18728), .dout(n19662));
  jand g19542(.dina(n18737), .dinb(n18713), .dout(n19663));
  jnot g19543(.din(n19663), .dout(n19664));
  jand g19544(.dina(n19664), .dinb(n19662), .dout(n19665));
  jnot g19545(.din(n19665), .dout(n19666));
  jand g19546(.dina(n18716), .dinb(n18715), .dout(n19667));
  jnot g19547(.din(n19667), .dout(n19668));
  jor  g19548(.dina(n18726), .dinb(n18718), .dout(n19669));
  jand g19549(.dina(n19669), .dinb(n19668), .dout(n19670));
  jnot g19550(.din(n19670), .dout(n19671));
  jand g19551(.dina(n1688), .dinb(n2117), .dout(n19672));
  jand g19552(.dina(n2131), .dinb(n492), .dout(n19673));
  jand g19553(.dina(n19673), .dinb(n19672), .dout(n19674));
  jand g19554(.dina(n19674), .dinb(n2342), .dout(n19675));
  jand g19555(.dina(n921), .dinb(n873), .dout(n19676));
  jand g19556(.dina(n19676), .dinb(n1366), .dout(n19677));
  jand g19557(.dina(n19677), .dinb(n621), .dout(n19678));
  jand g19558(.dina(n19678), .dinb(n19675), .dout(n19679));
  jand g19559(.dina(n19679), .dinb(n16211), .dout(n19680));
  jand g19560(.dina(n7658), .dinb(n1697), .dout(n19681));
  jand g19561(.dina(n19681), .dinb(n12218), .dout(n19682));
  jand g19562(.dina(n2500), .dinb(n1308), .dout(n19683));
  jand g19563(.dina(n19683), .dinb(n9545), .dout(n19684));
  jand g19564(.dina(n447), .dinb(n1306), .dout(n19685));
  jand g19565(.dina(n1374), .dinb(n1370), .dout(n19686));
  jand g19566(.dina(n19686), .dinb(n19685), .dout(n19687));
  jand g19567(.dina(n19687), .dinb(n19684), .dout(n19688));
  jand g19568(.dina(n19688), .dinb(n19682), .dout(n19689));
  jand g19569(.dina(n1016), .dinb(n1284), .dout(n19690));
  jand g19570(.dina(n893), .dinb(n168), .dout(n19691));
  jand g19571(.dina(n7516), .dinb(n2693), .dout(n19692));
  jand g19572(.dina(n19692), .dinb(n19691), .dout(n19693));
  jand g19573(.dina(n7649), .dinb(n1476), .dout(n19694));
  jand g19574(.dina(n19694), .dinb(n19693), .dout(n19695));
  jand g19575(.dina(n19695), .dinb(n19690), .dout(n19696));
  jand g19576(.dina(n19696), .dinb(n19689), .dout(n19697));
  jand g19577(.dina(n3750), .dinb(n934), .dout(n19698));
  jand g19578(.dina(n1987), .dinb(n1561), .dout(n19699));
  jand g19579(.dina(n19699), .dinb(n5327), .dout(n19700));
  jand g19580(.dina(n931), .dinb(n925), .dout(n19701));
  jand g19581(.dina(n19701), .dinb(n662), .dout(n19702));
  jand g19582(.dina(n19702), .dinb(n19700), .dout(n19703));
  jand g19583(.dina(n9559), .dinb(n1968), .dout(n19704));
  jand g19584(.dina(n2357), .dinb(n639), .dout(n19705));
  jand g19585(.dina(n19705), .dinb(n19704), .dout(n19706));
  jand g19586(.dina(n19706), .dinb(n19703), .dout(n19707));
  jand g19587(.dina(n19707), .dinb(n19698), .dout(n19708));
  jand g19588(.dina(n15658), .dinb(n3136), .dout(n19709));
  jand g19589(.dina(n19709), .dinb(n3762), .dout(n19710));
  jand g19590(.dina(n19710), .dinb(n4464), .dout(n19711));
  jand g19591(.dina(n19711), .dinb(n19708), .dout(n19712));
  jand g19592(.dina(n19712), .dinb(n19697), .dout(n19713));
  jand g19593(.dina(n19713), .dinb(n19680), .dout(n19714));
  jnot g19594(.din(n19714), .dout(n19715));
  jand g19595(.dina(n15329), .dinb(n5076), .dout(n19716));
  jand g19596(.dina(n15327), .dinb(n5084), .dout(n19717));
  jand g19597(.dina(n15020), .dinb(n5082), .dout(n19718));
  jor  g19598(.dina(n19718), .dinb(n19717), .dout(n19719));
  jor  g19599(.dina(n19719), .dinb(n19716), .dout(n19720));
  jxor g19600(.dina(n19720), .dinb(n19715), .dout(n19721));
  jnot g19601(.din(n19721), .dout(n19722));
  jand g19602(.dina(n16632), .dinb(n2936), .dout(n19723));
  jand g19603(.dina(n16360), .dinb(n2943), .dout(n19724));
  jand g19604(.dina(n15579), .dinb(n3684), .dout(n19725));
  jand g19605(.dina(n15841), .dinb(n2940), .dout(n19726));
  jor  g19606(.dina(n19726), .dinb(n19725), .dout(n19727));
  jor  g19607(.dina(n19727), .dinb(n19724), .dout(n19728));
  jor  g19608(.dina(n19728), .dinb(n19723), .dout(n19729));
  jxor g19609(.dina(n19729), .dinb(n93), .dout(n19730));
  jxor g19610(.dina(n19730), .dinb(n19722), .dout(n19731));
  jxor g19611(.dina(n19731), .dinb(n19671), .dout(n19732));
  jnot g19612(.din(n19732), .dout(n19733));
  jand g19613(.dina(n16942), .dinb(n71), .dout(n19734));
  jand g19614(.dina(n16604), .dinb(n731), .dout(n19735));
  jand g19615(.dina(n16940), .dinb(n796), .dout(n19736));
  jor  g19616(.dina(n19736), .dinb(n19735), .dout(n19737));
  jand g19617(.dina(n16355), .dinb(n1806), .dout(n19738));
  jor  g19618(.dina(n19738), .dinb(n19737), .dout(n19739));
  jor  g19619(.dina(n19739), .dinb(n19734), .dout(n19740));
  jxor g19620(.dina(n19740), .dinb(n77), .dout(n19741));
  jxor g19621(.dina(n19741), .dinb(n19733), .dout(n19742));
  jxor g19622(.dina(n19742), .dinb(n19666), .dout(n19743));
  jnot g19623(.din(n19743), .dout(n19744));
  jand g19624(.dina(n17537), .dinb(n806), .dout(n19745));
  jand g19625(.dina(n17329), .dinb(n1612), .dout(n19746));
  jand g19626(.dina(n17535), .dinb(n1620), .dout(n19747));
  jor  g19627(.dina(n19747), .dinb(n19746), .dout(n19748));
  jand g19628(.dina(n17330), .dinb(n1644), .dout(n19749));
  jor  g19629(.dina(n19749), .dinb(n19748), .dout(n19750));
  jor  g19630(.dina(n19750), .dinb(n19745), .dout(n19751));
  jxor g19631(.dina(n19751), .dinb(n65), .dout(n19752));
  jxor g19632(.dina(n19752), .dinb(n19744), .dout(n19753));
  jxor g19633(.dina(n19753), .dinb(n19661), .dout(n19754));
  jnot g19634(.din(n19754), .dout(n19755));
  jand g19635(.dina(n18502), .dinb(n1819), .dout(n19756));
  jand g19636(.dina(n18292), .dinb(n2243), .dout(n19757));
  jand g19637(.dina(n18293), .dinb(n2180), .dout(n19758));
  jand g19638(.dina(n17942), .dinb(n2185), .dout(n19759));
  jor  g19639(.dina(n19759), .dinb(n19758), .dout(n19760));
  jor  g19640(.dina(n19760), .dinb(n19757), .dout(n19761));
  jor  g19641(.dina(n19761), .dinb(n19756), .dout(n19762));
  jxor g19642(.dina(n19762), .dinb(n2196), .dout(n19763));
  jxor g19643(.dina(n19763), .dinb(n19755), .dout(n19764));
  jxor g19644(.dina(n19764), .dinb(n19656), .dout(n19765));
  jand g19645(.dina(n19399), .dinb(n2743), .dout(n19766));
  jand g19646(.dina(n19220), .dinb(n2752), .dout(n19767));
  jand g19647(.dina(n18914), .dinb(n2748), .dout(n19768));
  jand g19648(.dina(n18488), .dinb(n2757), .dout(n19769));
  jor  g19649(.dina(n19769), .dinb(n19768), .dout(n19770));
  jor  g19650(.dina(n19770), .dinb(n19767), .dout(n19771));
  jor  g19651(.dina(n19771), .dinb(n19766), .dout(n19772));
  jxor g19652(.dina(n19772), .dinb(\a[17] ), .dout(n19773));
  jxor g19653(.dina(n19773), .dinb(n19765), .dout(n19774));
  jxor g19654(.dina(n19774), .dinb(n19651), .dout(n19775));
  jnot g19655(.din(n19775), .dout(n19776));
  jand g19656(.dina(n19373), .dinb(n19219), .dout(n19777));
  jand g19657(.dina(n19374), .dinb(n19231), .dout(n19778));
  jor  g19658(.dina(n19778), .dinb(n19777), .dout(n19779));
  jand g19659(.dina(n19366), .dinb(n19236), .dout(n19780));
  jnot g19660(.din(n19780), .dout(n19781));
  jor  g19661(.dina(n19372), .dinb(n19368), .dout(n19782));
  jand g19662(.dina(n19782), .dinb(n19781), .dout(n19783));
  jor  g19663(.dina(n19849), .dinb(n19241), .dout(n19784));
  jnot g19664(.din(n19784), .dout(n19785));
  jand g19665(.dina(n19365), .dinb(n19249), .dout(n19786));
  jor  g19666(.dina(n19786), .dinb(n19785), .dout(n19787));
  jnot g19667(.din(n19259), .dout(n19788));
  jand g19668(.dina(n19345), .dinb(n19788), .dout(n19789));
  jnot g19669(.din(n19789), .dout(n19790));
  jor  g19670(.dina(n19354), .dinb(n19346), .dout(n19791));
  jand g19671(.dina(n19791), .dinb(n19790), .dout(n19792));
  jnot g19672(.din(n19264), .dout(n19793));
  jand g19673(.dina(n19335), .dinb(n19793), .dout(n19794));
  jnot g19674(.din(n19794), .dout(n19795));
  jor  g19675(.dina(n19344), .dinb(n19336), .dout(n19796));
  jand g19676(.dina(n19796), .dinb(n19795), .dout(n19797));
  jnot g19677(.din(n19269), .dout(n19798));
  jand g19678(.dina(n19325), .dinb(n19798), .dout(n19799));
  jnot g19679(.din(n19799), .dout(n19800));
  jor  g19680(.dina(n19334), .dinb(n19326), .dout(n19801));
  jand g19681(.dina(n19801), .dinb(n19800), .dout(n19802));
  jnot g19682(.din(n19274), .dout(n19803));
  jand g19683(.dina(n19315), .dinb(n19803), .dout(n19804));
  jnot g19684(.din(n19804), .dout(n19805));
  jor  g19685(.dina(n19324), .dinb(n19316), .dout(n19806));
  jand g19686(.dina(n19806), .dinb(n19805), .dout(n19807));
  jnot g19687(.din(n19807), .dout(n19808));
  jand g19688(.dina(n19304), .dinb(n19281), .dout(n19809));
  jnot g19689(.din(n19809), .dout(n19810));
  jor  g19690(.dina(n19314), .dinb(n19306), .dout(n19811));
  jand g19691(.dina(n19811), .dinb(n19810), .dout(n19812));
  jnot g19692(.din(n19812), .dout(n19813));
  jor  g19693(.dina(n19302), .dinb(n19133), .dout(n19814));
  jand g19694(.dina(n19303), .dinb(n19286), .dout(n19815));
  jnot g19695(.din(n19815), .dout(n19816));
  jand g19696(.dina(n19816), .dinb(n19814), .dout(n19817));
  jnot g19697(.din(n19817), .dout(n19818));
  jand g19698(.dina(n12284), .dinb(n5076), .dout(n19819));
  jand g19699(.dina(n12282), .dinb(n5084), .dout(n19820));
  jand g19700(.dina(n11798), .dinb(n5082), .dout(n19821));
  jand g19701(.dina(n11646), .dinb(n6050), .dout(n19822));
  jor  g19702(.dina(n19822), .dinb(n19821), .dout(n19823));
  jor  g19703(.dina(n19823), .dinb(n19820), .dout(n19824));
  jor  g19704(.dina(n19824), .dinb(n19819), .dout(n19825));
  jand g19705(.dina(n9761), .dinb(n3960), .dout(n19826));
  jand g19706(.dina(n521), .dinb(n469), .dout(n19827));
  jand g19707(.dina(n19827), .dinb(n1431), .dout(n19828));
  jand g19708(.dina(n2352), .dinb(n496), .dout(n19829));
  jand g19709(.dina(n19829), .dinb(n19828), .dout(n19830));
  jand g19710(.dina(n19830), .dinb(n5492), .dout(n19831));
  jand g19711(.dina(n630), .dinb(n713), .dout(n19832));
  jand g19712(.dina(n19832), .dinb(n1827), .dout(n19833));
  jand g19713(.dina(n19833), .dinb(n3880), .dout(n19834));
  jand g19714(.dina(n19834), .dinb(n993), .dout(n19835));
  jand g19715(.dina(n1096), .dinb(n130), .dout(n19836));
  jand g19716(.dina(n19836), .dinb(n2044), .dout(n19837));
  jand g19717(.dina(n11224), .dinb(n4531), .dout(n19838));
  jand g19718(.dina(n19838), .dinb(n19837), .dout(n19839));
  jand g19719(.dina(n19839), .dinb(n19835), .dout(n19840));
  jand g19720(.dina(n19840), .dinb(n19831), .dout(n19841));
  jand g19721(.dina(n19841), .dinb(n19826), .dout(n19842));
  jand g19722(.dina(n6323), .dinb(n5382), .dout(n19843));
  jand g19723(.dina(n19843), .dinb(n19842), .dout(n19844));
  jxor g19724(.dina(n19844), .dinb(n19132), .dout(n19845));
  jnot g19725(.din(n3869), .dout(n19846));
  jor  g19726(.dina(n19846), .dinb(n3864), .dout(n19847));
  jand g19727(.dina(n19847), .dinb(n16924), .dout(n19848));
  jxor g19728(.dina(n19848), .dinb(n4050), .dout(n19849));
  jxor g19729(.dina(n19849), .dinb(n19845), .dout(n19850));
  jxor g19730(.dina(n19850), .dinb(n19825), .dout(n19851));
  jxor g19731(.dina(n19851), .dinb(n19818), .dout(n19852));
  jxor g19732(.dina(n19852), .dinb(n19813), .dout(n19853));
  jnot g19733(.din(n19853), .dout(n19854));
  jand g19734(.dina(n12671), .dinb(n2936), .dout(n19855));
  jand g19735(.dina(n12536), .dinb(n2940), .dout(n19856));
  jand g19736(.dina(n12669), .dinb(n2943), .dout(n19857));
  jor  g19737(.dina(n19857), .dinb(n19856), .dout(n19858));
  jand g19738(.dina(n12547), .dinb(n3684), .dout(n19859));
  jor  g19739(.dina(n19859), .dinb(n19858), .dout(n19860));
  jor  g19740(.dina(n19860), .dinb(n19855), .dout(n19861));
  jxor g19741(.dina(n19861), .dinb(n93), .dout(n19862));
  jxor g19742(.dina(n19862), .dinb(n19854), .dout(n19863));
  jnot g19743(.din(n19863), .dout(n19864));
  jand g19744(.dina(n13627), .dinb(n71), .dout(n19865));
  jand g19745(.dina(n13478), .dinb(n731), .dout(n19866));
  jand g19746(.dina(n13469), .dinb(n796), .dout(n19867));
  jor  g19747(.dina(n19867), .dinb(n19866), .dout(n19868));
  jand g19748(.dina(n13248), .dinb(n1806), .dout(n19869));
  jor  g19749(.dina(n19869), .dinb(n19868), .dout(n19870));
  jor  g19750(.dina(n19870), .dinb(n19865), .dout(n19871));
  jxor g19751(.dina(n19871), .dinb(n77), .dout(n19872));
  jxor g19752(.dina(n19872), .dinb(n19864), .dout(n19873));
  jxor g19753(.dina(n19873), .dinb(n19808), .dout(n19874));
  jand g19754(.dina(n14579), .dinb(n806), .dout(n19875));
  jand g19755(.dina(n14448), .dinb(n1620), .dout(n19876));
  jand g19756(.dina(n14249), .dinb(n1612), .dout(n19877));
  jand g19757(.dina(n13614), .dinb(n1644), .dout(n19878));
  jor  g19758(.dina(n19878), .dinb(n19877), .dout(n19879));
  jor  g19759(.dina(n19879), .dinb(n19876), .dout(n19880));
  jor  g19760(.dina(n19880), .dinb(n19875), .dout(n19881));
  jxor g19761(.dina(n19881), .dinb(n65), .dout(n19882));
  jxor g19762(.dina(n19882), .dinb(n19874), .dout(n19883));
  jxor g19763(.dina(n19883), .dinb(n19802), .dout(n19884));
  jand g19764(.dina(n15317), .dinb(n1819), .dout(n19885));
  jand g19765(.dina(n15315), .dinb(n2243), .dout(n19886));
  jand g19766(.dina(n14549), .dinb(n2180), .dout(n19887));
  jand g19767(.dina(n14447), .dinb(n2185), .dout(n19888));
  jor  g19768(.dina(n19888), .dinb(n19887), .dout(n19889));
  jor  g19769(.dina(n19889), .dinb(n19886), .dout(n19890));
  jor  g19770(.dina(n19890), .dinb(n19885), .dout(n19891));
  jxor g19771(.dina(n19891), .dinb(n2196), .dout(n19892));
  jxor g19772(.dina(n19892), .dinb(n19884), .dout(n19893));
  jxor g19773(.dina(n19893), .dinb(n19797), .dout(n19894));
  jand g19774(.dina(n16084), .dinb(n2743), .dout(n19895));
  jand g19775(.dina(n15829), .dinb(n2748), .dout(n19896));
  jand g19776(.dina(n16082), .dinb(n2752), .dout(n19897));
  jor  g19777(.dina(n19897), .dinb(n19896), .dout(n19898));
  jand g19778(.dina(n15567), .dinb(n2757), .dout(n19899));
  jor  g19779(.dina(n19899), .dinb(n19898), .dout(n19900));
  jor  g19780(.dina(n19900), .dinb(n19895), .dout(n19901));
  jxor g19781(.dina(n19901), .dinb(n2441), .dout(n19902));
  jxor g19782(.dina(n19902), .dinb(n19894), .dout(n19903));
  jxor g19783(.dina(n19903), .dinb(n19792), .dout(n19904));
  jnot g19784(.din(n19254), .dout(n19905));
  jand g19785(.dina(n19355), .dinb(n19905), .dout(n19906));
  jnot g19786(.din(n19906), .dout(n19907));
  jor  g19787(.dina(n19364), .dinb(n19356), .dout(n19908));
  jand g19788(.dina(n19908), .dinb(n19907), .dout(n19909));
  jand g19789(.dina(n16930), .dinb(n3423), .dout(n19910));
  jand g19790(.dina(n16592), .dinb(n3428), .dout(n19911));
  jand g19791(.dina(n16928), .dinb(n3569), .dout(n19912));
  jor  g19792(.dina(n19912), .dinb(n19911), .dout(n19913));
  jand g19793(.dina(n16343), .dinb(n3210), .dout(n19914));
  jor  g19794(.dina(n19914), .dinb(n19913), .dout(n19915));
  jor  g19795(.dina(n19915), .dinb(n19910), .dout(n19916));
  jxor g19796(.dina(n19916), .dinb(n3473), .dout(n19917));
  jxor g19797(.dina(n19917), .dinb(n19909), .dout(n19918));
  jxor g19798(.dina(n19918), .dinb(n19904), .dout(n19919));
  jxor g19799(.dina(n19919), .dinb(n19787), .dout(n19920));
  jnot g19800(.din(n19920), .dout(n19921));
  jxor g19801(.dina(n19921), .dinb(n19783), .dout(n19922));
  jxor g19802(.dina(n19922), .dinb(n19373), .dout(n19923));
  jxor g19803(.dina(n19923), .dinb(n19779), .dout(n19924));
  jand g19804(.dina(n19924), .dinb(n3423), .dout(n19925));
  jand g19805(.dina(n19922), .dinb(n3569), .dout(n19926));
  jand g19806(.dina(n19373), .dinb(n3428), .dout(n19927));
  jand g19807(.dina(n19219), .dinb(n3210), .dout(n19928));
  jor  g19808(.dina(n19928), .dinb(n19927), .dout(n19929));
  jor  g19809(.dina(n19929), .dinb(n19926), .dout(n19930));
  jor  g19810(.dina(n19930), .dinb(n19925), .dout(n19931));
  jxor g19811(.dina(n19931), .dinb(n3473), .dout(n19932));
  jxor g19812(.dina(n19932), .dinb(n19776), .dout(n19933));
  jxor g19813(.dina(n19933), .dinb(n19646), .dout(n19934));
  jnot g19814(.din(n19894), .dout(n19935));
  jor  g19815(.dina(n19902), .dinb(n19935), .dout(n19936));
  jor  g19816(.dina(n19903), .dinb(n19792), .dout(n19937));
  jand g19817(.dina(n19937), .dinb(n19936), .dout(n19938));
  jnot g19818(.din(n19938), .dout(n19939));
  jnot g19819(.din(n19884), .dout(n19940));
  jor  g19820(.dina(n19892), .dinb(n19940), .dout(n19941));
  jor  g19821(.dina(n19893), .dinb(n19797), .dout(n19942));
  jand g19822(.dina(n19942), .dinb(n19941), .dout(n19943));
  jnot g19823(.din(n19874), .dout(n19944));
  jor  g19824(.dina(n19882), .dinb(n19944), .dout(n19945));
  jor  g19825(.dina(n19883), .dinb(n19802), .dout(n19946));
  jand g19826(.dina(n19946), .dinb(n19945), .dout(n19947));
  jor  g19827(.dina(n19872), .dinb(n19864), .dout(n19948));
  jand g19828(.dina(n19873), .dinb(n19808), .dout(n19949));
  jnot g19829(.din(n19949), .dout(n19950));
  jand g19830(.dina(n19950), .dinb(n19948), .dout(n19951));
  jand g19831(.dina(n19852), .dinb(n19813), .dout(n19952));
  jnot g19832(.din(n19952), .dout(n19953));
  jor  g19833(.dina(n19862), .dinb(n19854), .dout(n19954));
  jand g19834(.dina(n19954), .dinb(n19953), .dout(n19955));
  jnot g19835(.din(n19955), .dout(n19956));
  jand g19836(.dina(n19850), .dinb(n19825), .dout(n19957));
  jand g19837(.dina(n19851), .dinb(n19818), .dout(n19958));
  jor  g19838(.dina(n19958), .dinb(n19957), .dout(n19959));
  jand g19839(.dina(n10705), .dinb(n1453), .dout(n19960));
  jand g19840(.dina(n19960), .dinb(n2124), .dout(n19961));
  jand g19841(.dina(n4530), .dinb(n132), .dout(n19962));
  jand g19842(.dina(n19962), .dinb(n2023), .dout(n19963));
  jand g19843(.dina(n19963), .dinb(n713), .dout(n19964));
  jand g19844(.dina(n19964), .dinb(n3998), .dout(n19965));
  jand g19845(.dina(n6443), .dinb(n1212), .dout(n19966));
  jand g19846(.dina(n19966), .dinb(n3217), .dout(n19967));
  jand g19847(.dina(n1360), .dinb(n699), .dout(n19968));
  jand g19848(.dina(n19968), .dinb(n10141), .dout(n19969));
  jand g19849(.dina(n19969), .dinb(n19967), .dout(n19970));
  jand g19850(.dina(n19970), .dinb(n593), .dout(n19971));
  jand g19851(.dina(n19971), .dinb(n19965), .dout(n19972));
  jand g19852(.dina(n19972), .dinb(n5498), .dout(n19973));
  jand g19853(.dina(n19973), .dinb(n19961), .dout(n19974));
  jnot g19854(.din(n19974), .dout(n19975));
  jor  g19855(.dina(n19844), .dinb(n19132), .dout(n19976));
  jand g19856(.dina(n19849), .dinb(n19845), .dout(n19977));
  jnot g19857(.din(n19977), .dout(n19978));
  jand g19858(.dina(n19978), .dinb(n19976), .dout(n19979));
  jxor g19859(.dina(n19979), .dinb(n19975), .dout(n19980));
  jand g19860(.dina(n12696), .dinb(n5076), .dout(n19981));
  jand g19861(.dina(n12547), .dinb(n5084), .dout(n19982));
  jand g19862(.dina(n11798), .dinb(n6050), .dout(n19983));
  jand g19863(.dina(n12282), .dinb(n5082), .dout(n19984));
  jor  g19864(.dina(n19984), .dinb(n19983), .dout(n19985));
  jor  g19865(.dina(n19985), .dinb(n19982), .dout(n19986));
  jor  g19866(.dina(n19986), .dinb(n19981), .dout(n19987));
  jxor g19867(.dina(n19987), .dinb(n19980), .dout(n19988));
  jxor g19868(.dina(n19988), .dinb(n19959), .dout(n19989));
  jnot g19869(.din(n19989), .dout(n19990));
  jand g19870(.dina(n13250), .dinb(n2936), .dout(n19991));
  jand g19871(.dina(n12669), .dinb(n2940), .dout(n19992));
  jand g19872(.dina(n13248), .dinb(n2943), .dout(n19993));
  jor  g19873(.dina(n19993), .dinb(n19992), .dout(n19994));
  jand g19874(.dina(n12536), .dinb(n3684), .dout(n19995));
  jor  g19875(.dina(n19995), .dinb(n19994), .dout(n19996));
  jor  g19876(.dina(n19996), .dinb(n19991), .dout(n19997));
  jxor g19877(.dina(n19997), .dinb(n93), .dout(n19998));
  jxor g19878(.dina(n19998), .dinb(n19990), .dout(n19999));
  jxor g19879(.dina(n19999), .dinb(n19956), .dout(n20000));
  jnot g19880(.din(n20000), .dout(n20001));
  jand g19881(.dina(n13616), .dinb(n71), .dout(n20002));
  jand g19882(.dina(n13614), .dinb(n796), .dout(n20003));
  jand g19883(.dina(n13469), .dinb(n731), .dout(n20004));
  jand g19884(.dina(n13478), .dinb(n1806), .dout(n20005));
  jor  g19885(.dina(n20005), .dinb(n20004), .dout(n20006));
  jor  g19886(.dina(n20006), .dinb(n20003), .dout(n20007));
  jor  g19887(.dina(n20007), .dinb(n20002), .dout(n20008));
  jxor g19888(.dina(n20008), .dinb(n77), .dout(n20009));
  jxor g19889(.dina(n20009), .dinb(n20001), .dout(n20010));
  jxor g19890(.dina(n20010), .dinb(n19951), .dout(n20011));
  jand g19891(.dina(n14562), .dinb(n806), .dout(n20012));
  jand g19892(.dina(n14448), .dinb(n1612), .dout(n20013));
  jand g19893(.dina(n14447), .dinb(n1620), .dout(n20014));
  jor  g19894(.dina(n20014), .dinb(n20013), .dout(n20015));
  jand g19895(.dina(n14249), .dinb(n1644), .dout(n20016));
  jor  g19896(.dina(n20016), .dinb(n20015), .dout(n20017));
  jor  g19897(.dina(n20017), .dinb(n20012), .dout(n20018));
  jxor g19898(.dina(n20018), .dinb(n65), .dout(n20019));
  jxor g19899(.dina(n20019), .dinb(n20011), .dout(n20020));
  jxor g19900(.dina(n20020), .dinb(n19947), .dout(n20021));
  jand g19901(.dina(n15569), .dinb(n1819), .dout(n20022));
  jand g19902(.dina(n15315), .dinb(n2180), .dout(n20023));
  jand g19903(.dina(n15567), .dinb(n2243), .dout(n20024));
  jor  g19904(.dina(n20024), .dinb(n20023), .dout(n20025));
  jand g19905(.dina(n14549), .dinb(n2185), .dout(n20026));
  jor  g19906(.dina(n20026), .dinb(n20025), .dout(n20027));
  jor  g19907(.dina(n20027), .dinb(n20022), .dout(n20028));
  jxor g19908(.dina(n20028), .dinb(n2196), .dout(n20029));
  jxor g19909(.dina(n20029), .dinb(n20021), .dout(n20030));
  jxor g19910(.dina(n20030), .dinb(n19943), .dout(n20031));
  jand g19911(.dina(n16345), .dinb(n2743), .dout(n20032));
  jand g19912(.dina(n16343), .dinb(n2752), .dout(n20033));
  jand g19913(.dina(n16082), .dinb(n2748), .dout(n20034));
  jand g19914(.dina(n15829), .dinb(n2757), .dout(n20035));
  jor  g19915(.dina(n20035), .dinb(n20034), .dout(n20036));
  jor  g19916(.dina(n20036), .dinb(n20033), .dout(n20037));
  jor  g19917(.dina(n20037), .dinb(n20032), .dout(n20038));
  jxor g19918(.dina(n20038), .dinb(n2441), .dout(n20039));
  jxor g19919(.dina(n20039), .dinb(n20031), .dout(n20040));
  jand g19920(.dina(n20040), .dinb(n19939), .dout(n20041));
  jnot g19921(.din(n20041), .dout(n20042));
  jxor g19922(.dina(n20040), .dinb(n19938), .dout(n20043));
  jand g19923(.dina(n17312), .dinb(n3423), .dout(n20044));
  jand g19924(.dina(n16592), .dinb(n3210), .dout(n20045));
  jor  g19925(.dina(n3428), .dinb(n3569), .dout(n20047));
  jand g19926(.dina(n20047), .dinb(n16924), .dout(n20048));
  jor  g19927(.dina(n20048), .dinb(n20045), .dout(n20049));
  jor  g19928(.dina(n20049), .dinb(n20044), .dout(n20050));
  jxor g19929(.dina(n20050), .dinb(n3473), .dout(n20051));
  jor  g19930(.dina(n20051), .dinb(n20043), .dout(n20052));
  jand g19931(.dina(n20052), .dinb(n20042), .dout(n20053));
  jnot g19932(.din(n20053), .dout(n20054));
  jnot g19933(.din(n19943), .dout(n20055));
  jand g19934(.dina(n20030), .dinb(n20055), .dout(n20056));
  jnot g19935(.din(n20056), .dout(n20057));
  jor  g19936(.dina(n20039), .dinb(n20031), .dout(n20058));
  jand g19937(.dina(n20058), .dinb(n20057), .dout(n20059));
  jand g19938(.dina(n3429), .dinb(n3426), .dout(n20060));
  jxor g19939(.dina(n20280), .dinb(n20059), .dout(n20067));
  jnot g19940(.din(n19947), .dout(n20068));
  jand g19941(.dina(n20020), .dinb(n20068), .dout(n20069));
  jnot g19942(.din(n20069), .dout(n20070));
  jor  g19943(.dina(n20029), .dinb(n20021), .dout(n20071));
  jand g19944(.dina(n20071), .dinb(n20070), .dout(n20072));
  jnot g19945(.din(n20072), .dout(n20073));
  jnot g19946(.din(n19951), .dout(n20074));
  jand g19947(.dina(n20010), .dinb(n20074), .dout(n20075));
  jnot g19948(.din(n20075), .dout(n20076));
  jor  g19949(.dina(n20019), .dinb(n20011), .dout(n20077));
  jand g19950(.dina(n20077), .dinb(n20076), .dout(n20078));
  jand g19951(.dina(n19999), .dinb(n19956), .dout(n20079));
  jnot g19952(.din(n20079), .dout(n20080));
  jor  g19953(.dina(n20009), .dinb(n20001), .dout(n20081));
  jand g19954(.dina(n20081), .dinb(n20080), .dout(n20082));
  jnot g19955(.din(n20082), .dout(n20083));
  jor  g19956(.dina(n19979), .dinb(n19975), .dout(n20084));
  jand g19957(.dina(n19987), .dinb(n19980), .dout(n20085));
  jnot g19958(.din(n20085), .dout(n20086));
  jand g19959(.dina(n20086), .dinb(n20084), .dout(n20087));
  jnot g19960(.din(n20087), .dout(n20088));
  jand g19961(.dina(n12684), .dinb(n5076), .dout(n20089));
  jand g19962(.dina(n12536), .dinb(n5084), .dout(n20090));
  jand g19963(.dina(n12547), .dinb(n5082), .dout(n20091));
  jand g19964(.dina(n12282), .dinb(n6050), .dout(n20092));
  jor  g19965(.dina(n20092), .dinb(n20091), .dout(n20093));
  jor  g19966(.dina(n20093), .dinb(n20090), .dout(n20094));
  jor  g19967(.dina(n20094), .dinb(n20089), .dout(n20095));
  jand g19968(.dina(n16205), .dinb(n563), .dout(n20096));
  jand g19969(.dina(n20096), .dinb(n13411), .dout(n20097));
  jand g19970(.dina(n20097), .dinb(n16180), .dout(n20098));
  jand g19971(.dina(n20098), .dinb(n1959), .dout(n20099));
  jand g19972(.dina(n20099), .dinb(n2356), .dout(n20100));
  jand g19973(.dina(n4448), .dinb(n1273), .dout(n20101));
  jand g19974(.dina(n20101), .dinb(n4639), .dout(n20102));
  jand g19975(.dina(n20102), .dinb(n325), .dout(n20103));
  jand g19976(.dina(n19693), .dinb(n3949), .dout(n20104));
  jand g19977(.dina(n481), .dinb(n351), .dout(n20105));
  jand g19978(.dina(n20105), .dinb(n1753), .dout(n20106));
  jand g19979(.dina(n20106), .dinb(n9359), .dout(n20107));
  jand g19980(.dina(n20107), .dinb(n4577), .dout(n20108));
  jand g19981(.dina(n2698), .dinb(n514), .dout(n20109));
  jand g19982(.dina(n20109), .dinb(n3897), .dout(n20110));
  jand g19983(.dina(n1716), .dinb(n881), .dout(n20111));
  jand g19984(.dina(n20111), .dinb(n5512), .dout(n20112));
  jand g19985(.dina(n20112), .dinb(n20110), .dout(n20113));
  jand g19986(.dina(n20113), .dinb(n20108), .dout(n20114));
  jand g19987(.dina(n20114), .dinb(n20104), .dout(n20115));
  jand g19988(.dina(n1706), .dinb(n808), .dout(n20116));
  jand g19989(.dina(n680), .dinb(n503), .dout(n20117));
  jand g19990(.dina(n1453), .dinb(n650), .dout(n20118));
  jand g19991(.dina(n20118), .dinb(n1167), .dout(n20119));
  jand g19992(.dina(n20119), .dinb(n20117), .dout(n20120));
  jand g19993(.dina(n20120), .dinb(n20116), .dout(n20121));
  jand g19994(.dina(n20121), .dinb(n20115), .dout(n20122));
  jand g19995(.dina(n20122), .dinb(n20103), .dout(n20123));
  jand g19996(.dina(n20123), .dinb(n20100), .dout(n20124));
  jxor g19997(.dina(n20124), .dinb(n19975), .dout(n20125));
  jxor g19998(.dina(n20125), .dinb(n20095), .dout(n20126));
  jxor g19999(.dina(n20126), .dinb(n20088), .dout(n20127));
  jnot g20000(.din(n20127), .dout(n20128));
  jand g20001(.dina(n19988), .dinb(n19959), .dout(n20129));
  jnot g20002(.din(n20129), .dout(n20130));
  jor  g20003(.dina(n19998), .dinb(n19990), .dout(n20131));
  jand g20004(.dina(n20131), .dinb(n20130), .dout(n20132));
  jxor g20005(.dina(n20132), .dinb(n20128), .dout(n20133));
  jnot g20006(.din(n20133), .dout(n20134));
  jand g20007(.dina(n13639), .dinb(n2936), .dout(n20135));
  jand g20008(.dina(n13248), .dinb(n2940), .dout(n20136));
  jand g20009(.dina(n13478), .dinb(n2943), .dout(n20137));
  jor  g20010(.dina(n20137), .dinb(n20136), .dout(n20138));
  jand g20011(.dina(n12669), .dinb(n3684), .dout(n20139));
  jor  g20012(.dina(n20139), .dinb(n20138), .dout(n20140));
  jor  g20013(.dina(n20140), .dinb(n20135), .dout(n20141));
  jxor g20014(.dina(n20141), .dinb(n93), .dout(n20142));
  jxor g20015(.dina(n20142), .dinb(n20134), .dout(n20143));
  jnot g20016(.din(n20143), .dout(n20144));
  jand g20017(.dina(n14251), .dinb(n71), .dout(n20145));
  jand g20018(.dina(n14249), .dinb(n796), .dout(n20146));
  jand g20019(.dina(n13614), .dinb(n731), .dout(n20147));
  jand g20020(.dina(n13469), .dinb(n1806), .dout(n20148));
  jor  g20021(.dina(n20148), .dinb(n20147), .dout(n20149));
  jor  g20022(.dina(n20149), .dinb(n20146), .dout(n20150));
  jor  g20023(.dina(n20150), .dinb(n20145), .dout(n20151));
  jxor g20024(.dina(n20151), .dinb(n77), .dout(n20152));
  jxor g20025(.dina(n20152), .dinb(n20144), .dout(n20153));
  jxor g20026(.dina(n20153), .dinb(n20083), .dout(n20154));
  jnot g20027(.din(n20154), .dout(n20155));
  jand g20028(.dina(n14551), .dinb(n806), .dout(n20156));
  jand g20029(.dina(n14549), .dinb(n1620), .dout(n20157));
  jand g20030(.dina(n14447), .dinb(n1612), .dout(n20158));
  jand g20031(.dina(n14448), .dinb(n1644), .dout(n20159));
  jor  g20032(.dina(n20159), .dinb(n20158), .dout(n20160));
  jor  g20033(.dina(n20160), .dinb(n20157), .dout(n20161));
  jor  g20034(.dina(n20161), .dinb(n20156), .dout(n20162));
  jxor g20035(.dina(n20162), .dinb(n65), .dout(n20163));
  jxor g20036(.dina(n20163), .dinb(n20155), .dout(n20164));
  jxor g20037(.dina(n20164), .dinb(n20078), .dout(n20165));
  jand g20038(.dina(n15831), .dinb(n1819), .dout(n20166));
  jand g20039(.dina(n15567), .dinb(n2180), .dout(n20167));
  jand g20040(.dina(n15829), .dinb(n2243), .dout(n20168));
  jor  g20041(.dina(n20168), .dinb(n20167), .dout(n20169));
  jand g20042(.dina(n15315), .dinb(n2185), .dout(n20170));
  jor  g20043(.dina(n20170), .dinb(n20169), .dout(n20171));
  jor  g20044(.dina(n20171), .dinb(n20166), .dout(n20172));
  jxor g20045(.dina(n20172), .dinb(n2196), .dout(n20173));
  jxor g20046(.dina(n20173), .dinb(n20165), .dout(n20174));
  jxor g20047(.dina(n20174), .dinb(n20073), .dout(n20175));
  jnot g20048(.din(n20175), .dout(n20176));
  jand g20049(.dina(n16594), .dinb(n2743), .dout(n20177));
  jand g20050(.dina(n16592), .dinb(n2752), .dout(n20178));
  jand g20051(.dina(n16343), .dinb(n2748), .dout(n20179));
  jand g20052(.dina(n16082), .dinb(n2757), .dout(n20180));
  jor  g20053(.dina(n20180), .dinb(n20179), .dout(n20181));
  jor  g20054(.dina(n20181), .dinb(n20178), .dout(n20182));
  jor  g20055(.dina(n20182), .dinb(n20177), .dout(n20183));
  jxor g20056(.dina(n20183), .dinb(n2441), .dout(n20184));
  jxor g20057(.dina(n20184), .dinb(n20176), .dout(n20185));
  jxor g20058(.dina(n20185), .dinb(n20067), .dout(n20186));
  jxor g20059(.dina(n20186), .dinb(n20054), .dout(n20187));
  jnot g20060(.din(n20187), .dout(n20188));
  jor  g20061(.dina(n19917), .dinb(n19909), .dout(n20189));
  jnot g20062(.din(n20189), .dout(n20190));
  jand g20063(.dina(n19918), .dinb(n19904), .dout(n20191));
  jor  g20064(.dina(n20191), .dinb(n20190), .dout(n20192));
  jxor g20065(.dina(n20051), .dinb(n20043), .dout(n20193));
  jand g20066(.dina(n20193), .dinb(n20192), .dout(n20194));
  jnot g20067(.din(n20194), .dout(n20195));
  jand g20068(.dina(n19919), .dinb(n19787), .dout(n20196));
  jnot g20069(.din(n20196), .dout(n20197));
  jor  g20070(.dina(n19921), .dinb(n19783), .dout(n20198));
  jand g20071(.dina(n20198), .dinb(n20197), .dout(n20199));
  jxor g20072(.dina(n20193), .dinb(n20192), .dout(n20200));
  jnot g20073(.din(n20200), .dout(n20201));
  jor  g20074(.dina(n20201), .dinb(n20199), .dout(n20202));
  jand g20075(.dina(n20202), .dinb(n20195), .dout(n20203));
  jxor g20076(.dina(n20203), .dinb(n20188), .dout(n20204));
  jxor g20077(.dina(n20201), .dinb(n20199), .dout(n20205));
  jand g20078(.dina(n20205), .dinb(n20204), .dout(n20206));
  jand g20079(.dina(n20205), .dinb(n19922), .dout(n20207));
  jand g20080(.dina(n19922), .dinb(n19373), .dout(n20208));
  jand g20081(.dina(n19923), .dinb(n19779), .dout(n20209));
  jor  g20082(.dina(n20209), .dinb(n20208), .dout(n20210));
  jxor g20083(.dina(n20205), .dinb(n19922), .dout(n20211));
  jand g20084(.dina(n20211), .dinb(n20210), .dout(n20212));
  jor  g20085(.dina(n20212), .dinb(n20207), .dout(n20213));
  jxor g20086(.dina(n20205), .dinb(n20204), .dout(n20214));
  jand g20087(.dina(n20214), .dinb(n20213), .dout(n20215));
  jor  g20088(.dina(n20215), .dinb(n20206), .dout(n20216));
  jand g20089(.dina(n20186), .dinb(n20054), .dout(n20217));
  jnot g20090(.din(n20217), .dout(n20218));
  jor  g20091(.dina(n20203), .dinb(n20188), .dout(n20219));
  jand g20092(.dina(n20219), .dinb(n20218), .dout(n20220));
  jor  g20093(.dina(n20280), .dinb(n20059), .dout(n20221));
  jnot g20094(.din(n20221), .dout(n20222));
  jand g20095(.dina(n20185), .dinb(n20067), .dout(n20223));
  jor  g20096(.dina(n20223), .dinb(n20222), .dout(n20224));
  jnot g20097(.din(n20078), .dout(n20225));
  jand g20098(.dina(n20164), .dinb(n20225), .dout(n20226));
  jnot g20099(.din(n20226), .dout(n20227));
  jor  g20100(.dina(n20173), .dinb(n20165), .dout(n20228));
  jand g20101(.dina(n20228), .dinb(n20227), .dout(n20229));
  jnot g20102(.din(n20229), .dout(n20230));
  jand g20103(.dina(n20153), .dinb(n20083), .dout(n20231));
  jnot g20104(.din(n20231), .dout(n20232));
  jor  g20105(.dina(n20163), .dinb(n20155), .dout(n20233));
  jand g20106(.dina(n20233), .dinb(n20232), .dout(n20234));
  jnot g20107(.din(n20234), .dout(n20235));
  jor  g20108(.dina(n20142), .dinb(n20134), .dout(n20236));
  jor  g20109(.dina(n20152), .dinb(n20144), .dout(n20237));
  jand g20110(.dina(n20237), .dinb(n20236), .dout(n20238));
  jnot g20111(.din(n20238), .dout(n20239));
  jand g20112(.dina(n20126), .dinb(n20088), .dout(n20240));
  jnot g20113(.din(n20240), .dout(n20241));
  jor  g20114(.dina(n20132), .dinb(n20128), .dout(n20242));
  jand g20115(.dina(n20242), .dinb(n20241), .dout(n20243));
  jnot g20116(.din(n20243), .dout(n20244));
  jand g20117(.dina(n12671), .dinb(n5076), .dout(n20245));
  jand g20118(.dina(n12669), .dinb(n5084), .dout(n20246));
  jand g20119(.dina(n12536), .dinb(n5082), .dout(n20247));
  jand g20120(.dina(n12547), .dinb(n6050), .dout(n20248));
  jor  g20121(.dina(n20248), .dinb(n20247), .dout(n20249));
  jor  g20122(.dina(n20249), .dinb(n20246), .dout(n20250));
  jor  g20123(.dina(n20250), .dinb(n20245), .dout(n20251));
  jor  g20124(.dina(n20124), .dinb(n19975), .dout(n20252));
  jand g20125(.dina(n20125), .dinb(n20095), .dout(n20253));
  jnot g20126(.din(n20253), .dout(n20254));
  jand g20127(.dina(n20254), .dinb(n20252), .dout(n20255));
  jnot g20128(.din(n20255), .dout(n20256));
  jand g20129(.dina(n13296), .dinb(n5196), .dout(n20257));
  jand g20130(.dina(n20257), .dinb(n2990), .dout(n20258));
  jand g20131(.dina(n20258), .dinb(n714), .dout(n20259));
  jand g20132(.dina(n20259), .dinb(n8377), .dout(n20260));
  jand g20133(.dina(n16167), .dinb(n2152), .dout(n20261));
  jand g20134(.dina(n1053), .dinb(n670), .dout(n20262));
  jand g20135(.dina(n20262), .dinb(n3758), .dout(n20263));
  jand g20136(.dina(n20263), .dinb(n20261), .dout(n20264));
  jand g20137(.dina(n20264), .dinb(n3812), .dout(n20265));
  jand g20138(.dina(n20265), .dinb(n586), .dout(n20266));
  jand g20139(.dina(n20266), .dinb(n839), .dout(n20267));
  jand g20140(.dina(n1577), .dinb(n925), .dout(n20268));
  jand g20141(.dina(n17799), .dinb(n15672), .dout(n20269));
  jand g20142(.dina(n20269), .dinb(n11236), .dout(n20270));
  jand g20143(.dina(n20270), .dinb(n534), .dout(n20271));
  jand g20144(.dina(n20271), .dinb(n20268), .dout(n20272));
  jand g20145(.dina(n20272), .dinb(n20267), .dout(n20273));
  jand g20146(.dina(n20273), .dinb(n3055), .dout(n20274));
  jand g20147(.dina(n20274), .dinb(n20260), .dout(n20275));
  jxor g20148(.dina(n20275), .dinb(n19974), .dout(n20276));
  jnot g20149(.din(n3209), .dout(n20277));
  jor  g20150(.dina(n20277), .dinb(n3204), .dout(n20278));
  jand g20151(.dina(n20278), .dinb(n16924), .dout(n20279));
  jxor g20152(.dina(n20279), .dinb(n3473), .dout(n20280));
  jxor g20153(.dina(n20280), .dinb(n20276), .dout(n20281));
  jxor g20154(.dina(n20281), .dinb(n20256), .dout(n20282));
  jxor g20155(.dina(n20282), .dinb(n20251), .dout(n20283));
  jnot g20156(.din(n20283), .dout(n20284));
  jand g20157(.dina(n13627), .dinb(n2936), .dout(n20285));
  jand g20158(.dina(n13469), .dinb(n2943), .dout(n20286));
  jand g20159(.dina(n13478), .dinb(n2940), .dout(n20287));
  jand g20160(.dina(n13248), .dinb(n3684), .dout(n20288));
  jor  g20161(.dina(n20288), .dinb(n20287), .dout(n20289));
  jor  g20162(.dina(n20289), .dinb(n20286), .dout(n20290));
  jor  g20163(.dina(n20290), .dinb(n20285), .dout(n20291));
  jxor g20164(.dina(n20291), .dinb(n93), .dout(n20292));
  jxor g20165(.dina(n20292), .dinb(n20284), .dout(n20293));
  jxor g20166(.dina(n20293), .dinb(n20244), .dout(n20294));
  jnot g20167(.din(n20294), .dout(n20295));
  jand g20168(.dina(n14579), .dinb(n71), .dout(n20296));
  jand g20169(.dina(n14249), .dinb(n731), .dout(n20297));
  jand g20170(.dina(n14448), .dinb(n796), .dout(n20298));
  jor  g20171(.dina(n20298), .dinb(n20297), .dout(n20299));
  jand g20172(.dina(n13614), .dinb(n1806), .dout(n20300));
  jor  g20173(.dina(n20300), .dinb(n20299), .dout(n20301));
  jor  g20174(.dina(n20301), .dinb(n20296), .dout(n20302));
  jxor g20175(.dina(n20302), .dinb(n77), .dout(n20303));
  jxor g20176(.dina(n20303), .dinb(n20295), .dout(n20304));
  jxor g20177(.dina(n20304), .dinb(n20239), .dout(n20305));
  jnot g20178(.din(n20305), .dout(n20306));
  jand g20179(.dina(n15317), .dinb(n806), .dout(n20307));
  jand g20180(.dina(n15315), .dinb(n1620), .dout(n20308));
  jand g20181(.dina(n14549), .dinb(n1612), .dout(n20309));
  jand g20182(.dina(n14447), .dinb(n1644), .dout(n20310));
  jor  g20183(.dina(n20310), .dinb(n20309), .dout(n20311));
  jor  g20184(.dina(n20311), .dinb(n20308), .dout(n20312));
  jor  g20185(.dina(n20312), .dinb(n20307), .dout(n20313));
  jxor g20186(.dina(n20313), .dinb(n65), .dout(n20314));
  jxor g20187(.dina(n20314), .dinb(n20306), .dout(n20315));
  jxor g20188(.dina(n20315), .dinb(n20235), .dout(n20316));
  jnot g20189(.din(n20316), .dout(n20317));
  jand g20190(.dina(n16084), .dinb(n1819), .dout(n20318));
  jand g20191(.dina(n16082), .dinb(n2243), .dout(n20319));
  jand g20192(.dina(n15829), .dinb(n2180), .dout(n20320));
  jand g20193(.dina(n15567), .dinb(n2185), .dout(n20321));
  jor  g20194(.dina(n20321), .dinb(n20320), .dout(n20322));
  jor  g20195(.dina(n20322), .dinb(n20319), .dout(n20323));
  jor  g20196(.dina(n20323), .dinb(n20318), .dout(n20324));
  jxor g20197(.dina(n20324), .dinb(n2196), .dout(n20325));
  jxor g20198(.dina(n20325), .dinb(n20317), .dout(n20326));
  jxor g20199(.dina(n20326), .dinb(n20230), .dout(n20327));
  jand g20200(.dina(n20174), .dinb(n20073), .dout(n20328));
  jnot g20201(.din(n20328), .dout(n20329));
  jor  g20202(.dina(n20184), .dinb(n20176), .dout(n20330));
  jand g20203(.dina(n20330), .dinb(n20329), .dout(n20331));
  jand g20204(.dina(n16930), .dinb(n2743), .dout(n20332));
  jand g20205(.dina(n16592), .dinb(n2748), .dout(n20333));
  jand g20206(.dina(n16928), .dinb(n2752), .dout(n20334));
  jor  g20207(.dina(n20334), .dinb(n20333), .dout(n20335));
  jand g20208(.dina(n16343), .dinb(n2757), .dout(n20336));
  jor  g20209(.dina(n20336), .dinb(n20335), .dout(n20337));
  jor  g20210(.dina(n20337), .dinb(n20332), .dout(n20338));
  jxor g20211(.dina(n20338), .dinb(n2441), .dout(n20339));
  jxor g20212(.dina(n20339), .dinb(n20331), .dout(n20340));
  jxor g20213(.dina(n20340), .dinb(n20327), .dout(n20341));
  jxor g20214(.dina(n20341), .dinb(n20224), .dout(n20342));
  jnot g20215(.din(n20342), .dout(n20343));
  jxor g20216(.dina(n20343), .dinb(n20220), .dout(n20344));
  jxor g20217(.dina(n20344), .dinb(n20204), .dout(n20345));
  jxor g20218(.dina(n20345), .dinb(n20216), .dout(n20346));
  jand g20219(.dina(n20346), .dinb(n4022), .dout(n20347));
  jand g20220(.dina(n20344), .dinb(n4220), .dout(n20348));
  jand g20221(.dina(n20204), .dinb(n4027), .dout(n20349));
  jand g20222(.dina(n20205), .dinb(n3870), .dout(n20350));
  jor  g20223(.dina(n20350), .dinb(n20349), .dout(n20351));
  jor  g20224(.dina(n20351), .dinb(n20348), .dout(n20352));
  jor  g20225(.dina(n20352), .dinb(n20347), .dout(n20353));
  jxor g20226(.dina(n20353), .dinb(\a[11] ), .dout(n20354));
  jand g20227(.dina(n20354), .dinb(n19934), .dout(n20355));
  jxor g20228(.dina(n19642), .dinb(n19641), .dout(n20356));
  jnot g20229(.din(n20356), .dout(n20357));
  jxor g20230(.dina(n20214), .dinb(n20213), .dout(n20358));
  jand g20231(.dina(n20358), .dinb(n4022), .dout(n20359));
  jand g20232(.dina(n20205), .dinb(n4027), .dout(n20360));
  jand g20233(.dina(n20204), .dinb(n4220), .dout(n20361));
  jor  g20234(.dina(n20361), .dinb(n20360), .dout(n20362));
  jand g20235(.dina(n19922), .dinb(n3870), .dout(n20363));
  jor  g20236(.dina(n20363), .dinb(n20362), .dout(n20364));
  jor  g20237(.dina(n20364), .dinb(n20359), .dout(n20365));
  jxor g20238(.dina(n20365), .dinb(n4050), .dout(n20366));
  jor  g20239(.dina(n20366), .dinb(n20357), .dout(n20367));
  jnot g20240(.din(n20367), .dout(n20368));
  jxor g20241(.dina(n19637), .dinb(n19636), .dout(n20369));
  jnot g20242(.din(n20369), .dout(n20370));
  jxor g20243(.dina(n20211), .dinb(n20210), .dout(n20371));
  jand g20244(.dina(n20371), .dinb(n4022), .dout(n20372));
  jand g20245(.dina(n20205), .dinb(n4220), .dout(n20373));
  jand g20246(.dina(n19922), .dinb(n4027), .dout(n20374));
  jand g20247(.dina(n19373), .dinb(n3870), .dout(n20375));
  jor  g20248(.dina(n20375), .dinb(n20374), .dout(n20376));
  jor  g20249(.dina(n20376), .dinb(n20373), .dout(n20377));
  jor  g20250(.dina(n20377), .dinb(n20372), .dout(n20378));
  jxor g20251(.dina(n20378), .dinb(n4050), .dout(n20379));
  jor  g20252(.dina(n20379), .dinb(n20370), .dout(n20380));
  jnot g20253(.din(n20380), .dout(n20381));
  jxor g20254(.dina(n19632), .dinb(n19631), .dout(n20382));
  jand g20255(.dina(n19924), .dinb(n4022), .dout(n20383));
  jand g20256(.dina(n19922), .dinb(n4220), .dout(n20384));
  jand g20257(.dina(n19373), .dinb(n4027), .dout(n20385));
  jand g20258(.dina(n19219), .dinb(n3870), .dout(n20386));
  jor  g20259(.dina(n20386), .dinb(n20385), .dout(n20387));
  jor  g20260(.dina(n20387), .dinb(n20384), .dout(n20388));
  jor  g20261(.dina(n20388), .dinb(n20383), .dout(n20389));
  jxor g20262(.dina(n20389), .dinb(\a[11] ), .dout(n20390));
  jand g20263(.dina(n20390), .dinb(n20382), .dout(n20391));
  jxor g20264(.dina(n19627), .dinb(n19626), .dout(n20392));
  jnot g20265(.din(n20392), .dout(n20393));
  jand g20266(.dina(n19375), .dinb(n4022), .dout(n20394));
  jand g20267(.dina(n19219), .dinb(n4027), .dout(n20395));
  jand g20268(.dina(n19373), .dinb(n4220), .dout(n20396));
  jor  g20269(.dina(n20396), .dinb(n20395), .dout(n20397));
  jand g20270(.dina(n19220), .dinb(n3870), .dout(n20398));
  jor  g20271(.dina(n20398), .dinb(n20397), .dout(n20399));
  jor  g20272(.dina(n20399), .dinb(n20394), .dout(n20400));
  jxor g20273(.dina(n20400), .dinb(n4050), .dout(n20401));
  jor  g20274(.dina(n20401), .dinb(n20393), .dout(n20402));
  jxor g20275(.dina(n19622), .dinb(n19621), .dout(n20403));
  jnot g20276(.din(n20403), .dout(n20404));
  jand g20277(.dina(n19387), .dinb(n4022), .dout(n20405));
  jand g20278(.dina(n19220), .dinb(n4027), .dout(n20406));
  jand g20279(.dina(n19219), .dinb(n4220), .dout(n20407));
  jor  g20280(.dina(n20407), .dinb(n20406), .dout(n20408));
  jand g20281(.dina(n18914), .dinb(n3870), .dout(n20409));
  jor  g20282(.dina(n20409), .dinb(n20408), .dout(n20410));
  jor  g20283(.dina(n20410), .dinb(n20405), .dout(n20411));
  jxor g20284(.dina(n20411), .dinb(n4050), .dout(n20412));
  jor  g20285(.dina(n20412), .dinb(n20404), .dout(n20413));
  jxor g20286(.dina(n19619), .dinb(n19618), .dout(n20414));
  jnot g20287(.din(n20414), .dout(n20415));
  jand g20288(.dina(n19399), .dinb(n4022), .dout(n20416));
  jand g20289(.dina(n19220), .dinb(n4220), .dout(n20417));
  jand g20290(.dina(n18914), .dinb(n4027), .dout(n20418));
  jand g20291(.dina(n18488), .dinb(n3870), .dout(n20419));
  jor  g20292(.dina(n20419), .dinb(n20418), .dout(n20420));
  jor  g20293(.dina(n20420), .dinb(n20417), .dout(n20421));
  jor  g20294(.dina(n20421), .dinb(n20416), .dout(n20422));
  jxor g20295(.dina(n20422), .dinb(n4050), .dout(n20423));
  jor  g20296(.dina(n20423), .dinb(n20415), .dout(n20424));
  jxor g20297(.dina(n19614), .dinb(n19613), .dout(n20425));
  jnot g20298(.din(n20425), .dout(n20426));
  jand g20299(.dina(n18916), .dinb(n4022), .dout(n20427));
  jand g20300(.dina(n18488), .dinb(n4027), .dout(n20428));
  jand g20301(.dina(n18914), .dinb(n4220), .dout(n20429));
  jor  g20302(.dina(n20429), .dinb(n20428), .dout(n20430));
  jand g20303(.dina(n18292), .dinb(n3870), .dout(n20431));
  jor  g20304(.dina(n20431), .dinb(n20430), .dout(n20432));
  jor  g20305(.dina(n20432), .dinb(n20427), .dout(n20433));
  jxor g20306(.dina(n20433), .dinb(n4050), .dout(n20434));
  jor  g20307(.dina(n20434), .dinb(n20426), .dout(n20435));
  jxor g20308(.dina(n19609), .dinb(n19608), .dout(n20436));
  jnot g20309(.din(n20436), .dout(n20437));
  jand g20310(.dina(n18490), .dinb(n4022), .dout(n20438));
  jand g20311(.dina(n18488), .dinb(n4220), .dout(n20439));
  jand g20312(.dina(n18292), .dinb(n4027), .dout(n20440));
  jand g20313(.dina(n18293), .dinb(n3870), .dout(n20441));
  jor  g20314(.dina(n20441), .dinb(n20440), .dout(n20442));
  jor  g20315(.dina(n20442), .dinb(n20439), .dout(n20443));
  jor  g20316(.dina(n20443), .dinb(n20438), .dout(n20444));
  jxor g20317(.dina(n20444), .dinb(n4050), .dout(n20445));
  jor  g20318(.dina(n20445), .dinb(n20437), .dout(n20446));
  jxor g20319(.dina(n19604), .dinb(n19603), .dout(n20447));
  jnot g20320(.din(n20447), .dout(n20448));
  jand g20321(.dina(n18502), .dinb(n4022), .dout(n20449));
  jand g20322(.dina(n18293), .dinb(n4027), .dout(n20450));
  jand g20323(.dina(n18292), .dinb(n4220), .dout(n20451));
  jor  g20324(.dina(n20451), .dinb(n20450), .dout(n20452));
  jand g20325(.dina(n17942), .dinb(n3870), .dout(n20453));
  jor  g20326(.dina(n20453), .dinb(n20452), .dout(n20454));
  jor  g20327(.dina(n20454), .dinb(n20449), .dout(n20455));
  jxor g20328(.dina(n20455), .dinb(n4050), .dout(n20456));
  jor  g20329(.dina(n20456), .dinb(n20448), .dout(n20457));
  jxor g20330(.dina(n19599), .dinb(n19598), .dout(n20458));
  jnot g20331(.din(n20458), .dout(n20459));
  jand g20332(.dina(n18514), .dinb(n4022), .dout(n20460));
  jand g20333(.dina(n17942), .dinb(n4027), .dout(n20461));
  jand g20334(.dina(n18293), .dinb(n4220), .dout(n20462));
  jor  g20335(.dina(n20462), .dinb(n20461), .dout(n20463));
  jand g20336(.dina(n17535), .dinb(n3870), .dout(n20464));
  jor  g20337(.dina(n20464), .dinb(n20463), .dout(n20465));
  jor  g20338(.dina(n20465), .dinb(n20460), .dout(n20466));
  jxor g20339(.dina(n20466), .dinb(n4050), .dout(n20467));
  jor  g20340(.dina(n20467), .dinb(n20459), .dout(n20468));
  jxor g20341(.dina(n19594), .dinb(n19593), .dout(n20469));
  jnot g20342(.din(n20469), .dout(n20470));
  jand g20343(.dina(n17944), .dinb(n4022), .dout(n20471));
  jand g20344(.dina(n17942), .dinb(n4220), .dout(n20472));
  jand g20345(.dina(n17535), .dinb(n4027), .dout(n20473));
  jand g20346(.dina(n17329), .dinb(n3870), .dout(n20474));
  jor  g20347(.dina(n20474), .dinb(n20473), .dout(n20475));
  jor  g20348(.dina(n20475), .dinb(n20472), .dout(n20476));
  jor  g20349(.dina(n20476), .dinb(n20471), .dout(n20477));
  jxor g20350(.dina(n20477), .dinb(n4050), .dout(n20478));
  jor  g20351(.dina(n20478), .dinb(n20470), .dout(n20479));
  jxor g20352(.dina(n19589), .dinb(n19588), .dout(n20480));
  jnot g20353(.din(n20480), .dout(n20481));
  jand g20354(.dina(n17537), .dinb(n4022), .dout(n20482));
  jand g20355(.dina(n17329), .dinb(n4027), .dout(n20483));
  jand g20356(.dina(n17535), .dinb(n4220), .dout(n20484));
  jor  g20357(.dina(n20484), .dinb(n20483), .dout(n20485));
  jand g20358(.dina(n17330), .dinb(n3870), .dout(n20486));
  jor  g20359(.dina(n20486), .dinb(n20485), .dout(n20487));
  jor  g20360(.dina(n20487), .dinb(n20482), .dout(n20488));
  jxor g20361(.dina(n20488), .dinb(n4050), .dout(n20489));
  jor  g20362(.dina(n20489), .dinb(n20481), .dout(n20490));
  jxor g20363(.dina(n19584), .dinb(n19583), .dout(n20491));
  jnot g20364(.din(n20491), .dout(n20492));
  jand g20365(.dina(n17549), .dinb(n4022), .dout(n20493));
  jand g20366(.dina(n17329), .dinb(n4220), .dout(n20494));
  jand g20367(.dina(n17330), .dinb(n4027), .dout(n20495));
  jand g20368(.dina(n16940), .dinb(n3870), .dout(n20496));
  jor  g20369(.dina(n20496), .dinb(n20495), .dout(n20497));
  jor  g20370(.dina(n20497), .dinb(n20494), .dout(n20498));
  jor  g20371(.dina(n20498), .dinb(n20493), .dout(n20499));
  jxor g20372(.dina(n20499), .dinb(n4050), .dout(n20500));
  jor  g20373(.dina(n20500), .dinb(n20492), .dout(n20501));
  jxor g20374(.dina(n19581), .dinb(n19580), .dout(n20502));
  jnot g20375(.din(n20502), .dout(n20503));
  jand g20376(.dina(n17561), .dinb(n4022), .dout(n20504));
  jand g20377(.dina(n16940), .dinb(n4027), .dout(n20505));
  jand g20378(.dina(n17330), .dinb(n4220), .dout(n20506));
  jor  g20379(.dina(n20506), .dinb(n20505), .dout(n20507));
  jand g20380(.dina(n16604), .dinb(n3870), .dout(n20508));
  jor  g20381(.dina(n20508), .dinb(n20507), .dout(n20509));
  jor  g20382(.dina(n20509), .dinb(n20504), .dout(n20510));
  jxor g20383(.dina(n20510), .dinb(n4050), .dout(n20511));
  jor  g20384(.dina(n20511), .dinb(n20503), .dout(n20512));
  jxor g20385(.dina(n19576), .dinb(n19575), .dout(n20513));
  jnot g20386(.din(n20513), .dout(n20514));
  jand g20387(.dina(n16942), .dinb(n4022), .dout(n20515));
  jand g20388(.dina(n16604), .dinb(n4027), .dout(n20516));
  jand g20389(.dina(n16940), .dinb(n4220), .dout(n20517));
  jor  g20390(.dina(n20517), .dinb(n20516), .dout(n20518));
  jand g20391(.dina(n16355), .dinb(n3870), .dout(n20519));
  jor  g20392(.dina(n20519), .dinb(n20518), .dout(n20520));
  jor  g20393(.dina(n20520), .dinb(n20515), .dout(n20521));
  jxor g20394(.dina(n20521), .dinb(n4050), .dout(n20522));
  jor  g20395(.dina(n20522), .dinb(n20514), .dout(n20523));
  jxor g20396(.dina(n19572), .dinb(n19564), .dout(n20524));
  jnot g20397(.din(n20524), .dout(n20525));
  jand g20398(.dina(n16606), .dinb(n4022), .dout(n20526));
  jand g20399(.dina(n16355), .dinb(n4027), .dout(n20527));
  jand g20400(.dina(n16604), .dinb(n4220), .dout(n20528));
  jor  g20401(.dina(n20528), .dinb(n20527), .dout(n20529));
  jand g20402(.dina(n16360), .dinb(n3870), .dout(n20530));
  jor  g20403(.dina(n20530), .dinb(n20529), .dout(n20531));
  jor  g20404(.dina(n20531), .dinb(n20526), .dout(n20532));
  jxor g20405(.dina(n20532), .dinb(n4050), .dout(n20533));
  jor  g20406(.dina(n20533), .dinb(n20525), .dout(n20534));
  jand g20407(.dina(n16616), .dinb(n4022), .dout(n20535));
  jand g20408(.dina(n16360), .dinb(n4027), .dout(n20536));
  jand g20409(.dina(n16355), .dinb(n4220), .dout(n20537));
  jor  g20410(.dina(n20537), .dinb(n20536), .dout(n20538));
  jand g20411(.dina(n15841), .dinb(n3870), .dout(n20539));
  jor  g20412(.dina(n20539), .dinb(n20538), .dout(n20540));
  jor  g20413(.dina(n20540), .dinb(n20535), .dout(n20541));
  jxor g20414(.dina(n20541), .dinb(n4050), .dout(n20542));
  jnot g20415(.din(n20542), .dout(n20543));
  jor  g20416(.dina(n19551), .dinb(n3473), .dout(n20544));
  jxor g20417(.dina(n20544), .dinb(n19559), .dout(n20545));
  jand g20418(.dina(n20545), .dinb(n20543), .dout(n20546));
  jand g20419(.dina(n19548), .dinb(\a[14] ), .dout(n20547));
  jxor g20420(.dina(n20547), .dinb(n19546), .dout(n20548));
  jnot g20421(.din(n20548), .dout(n20549));
  jand g20422(.dina(n16632), .dinb(n4022), .dout(n20550));
  jand g20423(.dina(n15841), .dinb(n4027), .dout(n20551));
  jand g20424(.dina(n16360), .dinb(n4220), .dout(n20552));
  jor  g20425(.dina(n20552), .dinb(n20551), .dout(n20553));
  jand g20426(.dina(n15579), .dinb(n3870), .dout(n20554));
  jor  g20427(.dina(n20554), .dinb(n20553), .dout(n20555));
  jor  g20428(.dina(n20555), .dinb(n20550), .dout(n20556));
  jxor g20429(.dina(n20556), .dinb(n4050), .dout(n20557));
  jor  g20430(.dina(n20557), .dinb(n20549), .dout(n20558));
  jand g20431(.dina(n15329), .dinb(n4022), .dout(n20559));
  jand g20432(.dina(n15020), .dinb(n4027), .dout(n20560));
  jand g20433(.dina(n15327), .dinb(n4220), .dout(n20561));
  jor  g20434(.dina(n20561), .dinb(n20560), .dout(n20562));
  jor  g20435(.dina(n20562), .dinb(n20559), .dout(n20563));
  jnot g20436(.din(n20563), .dout(n20564));
  jand g20437(.dina(n15020), .dinb(n3865), .dout(n20565));
  jnot g20438(.din(n20565), .dout(n20566));
  jand g20439(.dina(n20566), .dinb(\a[11] ), .dout(n20567));
  jand g20440(.dina(n20567), .dinb(n20564), .dout(n20568));
  jand g20441(.dina(n15580), .dinb(n4022), .dout(n20569));
  jand g20442(.dina(n15327), .dinb(n4027), .dout(n20570));
  jand g20443(.dina(n15579), .dinb(n4220), .dout(n20571));
  jor  g20444(.dina(n20571), .dinb(n20570), .dout(n20572));
  jand g20445(.dina(n15020), .dinb(n3870), .dout(n20573));
  jor  g20446(.dina(n20573), .dinb(n20572), .dout(n20574));
  jor  g20447(.dina(n20574), .dinb(n20569), .dout(n20575));
  jnot g20448(.din(n20575), .dout(n20576));
  jand g20449(.dina(n20576), .dinb(n20568), .dout(n20577));
  jand g20450(.dina(n20577), .dinb(n19548), .dout(n20578));
  jnot g20451(.din(n20578), .dout(n20579));
  jxor g20452(.dina(n20577), .dinb(n19548), .dout(n20580));
  jnot g20453(.din(n20580), .dout(n20581));
  jand g20454(.dina(n15848), .dinb(n4022), .dout(n20582));
  jand g20455(.dina(n15841), .dinb(n4220), .dout(n20583));
  jand g20456(.dina(n15579), .dinb(n4027), .dout(n20584));
  jand g20457(.dina(n15327), .dinb(n3870), .dout(n20585));
  jor  g20458(.dina(n20585), .dinb(n20584), .dout(n20586));
  jor  g20459(.dina(n20586), .dinb(n20583), .dout(n20587));
  jor  g20460(.dina(n20587), .dinb(n20582), .dout(n20588));
  jxor g20461(.dina(n20588), .dinb(n4050), .dout(n20589));
  jor  g20462(.dina(n20589), .dinb(n20581), .dout(n20590));
  jand g20463(.dina(n20590), .dinb(n20579), .dout(n20591));
  jnot g20464(.din(n20591), .dout(n20592));
  jxor g20465(.dina(n20557), .dinb(n20549), .dout(n20593));
  jand g20466(.dina(n20593), .dinb(n20592), .dout(n20594));
  jnot g20467(.din(n20594), .dout(n20595));
  jand g20468(.dina(n20595), .dinb(n20558), .dout(n20596));
  jnot g20469(.din(n20596), .dout(n20597));
  jxor g20470(.dina(n20545), .dinb(n20543), .dout(n20598));
  jand g20471(.dina(n20598), .dinb(n20597), .dout(n20599));
  jor  g20472(.dina(n20599), .dinb(n20546), .dout(n20600));
  jxor g20473(.dina(n20533), .dinb(n20525), .dout(n20601));
  jand g20474(.dina(n20601), .dinb(n20600), .dout(n20602));
  jnot g20475(.din(n20602), .dout(n20603));
  jand g20476(.dina(n20603), .dinb(n20534), .dout(n20604));
  jnot g20477(.din(n20604), .dout(n20605));
  jxor g20478(.dina(n20522), .dinb(n20514), .dout(n20606));
  jand g20479(.dina(n20606), .dinb(n20605), .dout(n20607));
  jnot g20480(.din(n20607), .dout(n20608));
  jand g20481(.dina(n20608), .dinb(n20523), .dout(n20609));
  jnot g20482(.din(n20609), .dout(n20610));
  jxor g20483(.dina(n20511), .dinb(n20503), .dout(n20611));
  jand g20484(.dina(n20611), .dinb(n20610), .dout(n20612));
  jnot g20485(.din(n20612), .dout(n20613));
  jand g20486(.dina(n20613), .dinb(n20512), .dout(n20614));
  jnot g20487(.din(n20614), .dout(n20615));
  jxor g20488(.dina(n20500), .dinb(n20492), .dout(n20616));
  jand g20489(.dina(n20616), .dinb(n20615), .dout(n20617));
  jnot g20490(.din(n20617), .dout(n20618));
  jand g20491(.dina(n20618), .dinb(n20501), .dout(n20619));
  jnot g20492(.din(n20619), .dout(n20620));
  jxor g20493(.dina(n20489), .dinb(n20481), .dout(n20621));
  jand g20494(.dina(n20621), .dinb(n20620), .dout(n20622));
  jnot g20495(.din(n20622), .dout(n20623));
  jand g20496(.dina(n20623), .dinb(n20490), .dout(n20624));
  jnot g20497(.din(n20624), .dout(n20625));
  jxor g20498(.dina(n20478), .dinb(n20470), .dout(n20626));
  jand g20499(.dina(n20626), .dinb(n20625), .dout(n20627));
  jnot g20500(.din(n20627), .dout(n20628));
  jand g20501(.dina(n20628), .dinb(n20479), .dout(n20629));
  jnot g20502(.din(n20629), .dout(n20630));
  jxor g20503(.dina(n20467), .dinb(n20459), .dout(n20631));
  jand g20504(.dina(n20631), .dinb(n20630), .dout(n20632));
  jnot g20505(.din(n20632), .dout(n20633));
  jand g20506(.dina(n20633), .dinb(n20468), .dout(n20634));
  jnot g20507(.din(n20634), .dout(n20635));
  jxor g20508(.dina(n20456), .dinb(n20448), .dout(n20636));
  jand g20509(.dina(n20636), .dinb(n20635), .dout(n20637));
  jnot g20510(.din(n20637), .dout(n20638));
  jand g20511(.dina(n20638), .dinb(n20457), .dout(n20639));
  jnot g20512(.din(n20639), .dout(n20640));
  jxor g20513(.dina(n20445), .dinb(n20437), .dout(n20641));
  jand g20514(.dina(n20641), .dinb(n20640), .dout(n20642));
  jnot g20515(.din(n20642), .dout(n20643));
  jand g20516(.dina(n20643), .dinb(n20446), .dout(n20644));
  jnot g20517(.din(n20644), .dout(n20645));
  jxor g20518(.dina(n20434), .dinb(n20426), .dout(n20646));
  jand g20519(.dina(n20646), .dinb(n20645), .dout(n20647));
  jnot g20520(.din(n20647), .dout(n20648));
  jand g20521(.dina(n20648), .dinb(n20435), .dout(n20649));
  jxor g20522(.dina(n20423), .dinb(n20415), .dout(n20650));
  jnot g20523(.din(n20650), .dout(n20651));
  jor  g20524(.dina(n20651), .dinb(n20649), .dout(n20652));
  jand g20525(.dina(n20652), .dinb(n20424), .dout(n20653));
  jxor g20526(.dina(n20412), .dinb(n20404), .dout(n20654));
  jnot g20527(.din(n20654), .dout(n20655));
  jor  g20528(.dina(n20655), .dinb(n20653), .dout(n20656));
  jand g20529(.dina(n20656), .dinb(n20413), .dout(n20657));
  jxor g20530(.dina(n20401), .dinb(n20393), .dout(n20658));
  jnot g20531(.din(n20658), .dout(n20659));
  jor  g20532(.dina(n20659), .dinb(n20657), .dout(n20660));
  jand g20533(.dina(n20660), .dinb(n20402), .dout(n20661));
  jnot g20534(.din(n20661), .dout(n20662));
  jxor g20535(.dina(n20390), .dinb(n20382), .dout(n20663));
  jand g20536(.dina(n20663), .dinb(n20662), .dout(n20664));
  jor  g20537(.dina(n20664), .dinb(n20391), .dout(n20665));
  jxor g20538(.dina(n20379), .dinb(n20370), .dout(n20666));
  jand g20539(.dina(n20666), .dinb(n20665), .dout(n20667));
  jor  g20540(.dina(n20667), .dinb(n20381), .dout(n20668));
  jxor g20541(.dina(n20366), .dinb(n20357), .dout(n20669));
  jand g20542(.dina(n20669), .dinb(n20668), .dout(n20670));
  jor  g20543(.dina(n20670), .dinb(n20368), .dout(n20671));
  jxor g20544(.dina(n20354), .dinb(n19934), .dout(n20672));
  jand g20545(.dina(n20672), .dinb(n20671), .dout(n20673));
  jor  g20546(.dina(n20673), .dinb(n20355), .dout(n20674));
  jor  g20547(.dina(n19932), .dinb(n19776), .dout(n20675));
  jnot g20548(.din(n20675), .dout(n20676));
  jand g20549(.dina(n19933), .dinb(n19646), .dout(n20677));
  jor  g20550(.dina(n20677), .dinb(n20676), .dout(n20678));
  jand g20551(.dina(n19773), .dinb(n19765), .dout(n20679));
  jand g20552(.dina(n19774), .dinb(n19651), .dout(n20680));
  jor  g20553(.dina(n20680), .dinb(n20679), .dout(n20681));
  jor  g20554(.dina(n19763), .dinb(n19755), .dout(n20682));
  jand g20555(.dina(n19764), .dinb(n19656), .dout(n20683));
  jnot g20556(.din(n20683), .dout(n20684));
  jand g20557(.dina(n20684), .dinb(n20682), .dout(n20685));
  jnot g20558(.din(n20685), .dout(n20686));
  jor  g20559(.dina(n19752), .dinb(n19744), .dout(n20687));
  jand g20560(.dina(n19753), .dinb(n19661), .dout(n20688));
  jnot g20561(.din(n20688), .dout(n20689));
  jand g20562(.dina(n20689), .dinb(n20687), .dout(n20690));
  jnot g20563(.din(n20690), .dout(n20691));
  jor  g20564(.dina(n19741), .dinb(n19733), .dout(n20692));
  jand g20565(.dina(n19742), .dinb(n19666), .dout(n20693));
  jnot g20566(.din(n20693), .dout(n20694));
  jand g20567(.dina(n20694), .dinb(n20692), .dout(n20695));
  jnot g20568(.din(n20695), .dout(n20696));
  jor  g20569(.dina(n19730), .dinb(n19722), .dout(n20697));
  jand g20570(.dina(n19731), .dinb(n19671), .dout(n20698));
  jnot g20571(.din(n20698), .dout(n20699));
  jand g20572(.dina(n20699), .dinb(n20697), .dout(n20700));
  jnot g20573(.din(n20700), .dout(n20701));
  jand g20574(.dina(n15580), .dinb(n5076), .dout(n20702));
  jand g20575(.dina(n15327), .dinb(n5082), .dout(n20703));
  jor  g20576(.dina(n20703), .dinb(n20702), .dout(n20704));
  jand g20577(.dina(n15579), .dinb(n5084), .dout(n20705));
  jand g20578(.dina(n15020), .dinb(n6050), .dout(n20706));
  jor  g20579(.dina(n20706), .dinb(n20705), .dout(n20707));
  jor  g20580(.dina(n20707), .dinb(n20704), .dout(n20708));
  jand g20581(.dina(n19720), .dinb(n19715), .dout(n20709));
  jnot g20582(.din(n20709), .dout(n20710));
  jand g20583(.dina(n12597), .dinb(n4460), .dout(n20711));
  jand g20584(.dina(n13538), .dinb(n1890), .dout(n20712));
  jand g20585(.dina(n20712), .dinb(n20711), .dout(n20713));
  jand g20586(.dina(n16211), .dinb(n1971), .dout(n20714));
  jand g20587(.dina(n20714), .dinb(n20713), .dout(n20715));
  jand g20588(.dina(n950), .dinb(n532), .dout(n20716));
  jand g20589(.dina(n20716), .dinb(n1559), .dout(n20717));
  jand g20590(.dina(n964), .dinb(n653), .dout(n20718));
  jand g20591(.dina(n20718), .dinb(n6443), .dout(n20719));
  jand g20592(.dina(n17823), .dinb(n2587), .dout(n20720));
  jand g20593(.dina(n20720), .dinb(n20719), .dout(n20721));
  jand g20594(.dina(n20721), .dinb(n20717), .dout(n20722));
  jand g20595(.dina(n2023), .dinb(n925), .dout(n20723));
  jand g20596(.dina(n20723), .dinb(n1426), .dout(n20724));
  jand g20597(.dina(n7789), .dinb(n641), .dout(n20725));
  jand g20598(.dina(n20725), .dinb(n20724), .dout(n20726));
  jand g20599(.dina(n20726), .dinb(n20722), .dout(n20727));
  jand g20600(.dina(n20727), .dinb(n7823), .dout(n20728));
  jand g20601(.dina(n20728), .dinb(n4440), .dout(n20729));
  jand g20602(.dina(n20729), .dinb(n20715), .dout(n20730));
  jxor g20603(.dina(n20730), .dinb(n20710), .dout(n20731));
  jxor g20604(.dina(n20731), .dinb(n20708), .dout(n20732));
  jnot g20605(.din(n20732), .dout(n20733));
  jand g20606(.dina(n16616), .dinb(n2936), .dout(n20734));
  jand g20607(.dina(n16360), .dinb(n2940), .dout(n20735));
  jand g20608(.dina(n16355), .dinb(n2943), .dout(n20736));
  jor  g20609(.dina(n20736), .dinb(n20735), .dout(n20737));
  jand g20610(.dina(n15841), .dinb(n3684), .dout(n20738));
  jor  g20611(.dina(n20738), .dinb(n20737), .dout(n20739));
  jor  g20612(.dina(n20739), .dinb(n20734), .dout(n20740));
  jxor g20613(.dina(n20740), .dinb(n93), .dout(n20741));
  jxor g20614(.dina(n20741), .dinb(n20733), .dout(n20742));
  jxor g20615(.dina(n20742), .dinb(n20701), .dout(n20743));
  jnot g20616(.din(n20743), .dout(n20744));
  jand g20617(.dina(n17561), .dinb(n71), .dout(n20745));
  jand g20618(.dina(n16940), .dinb(n731), .dout(n20746));
  jand g20619(.dina(n17330), .dinb(n796), .dout(n20747));
  jor  g20620(.dina(n20747), .dinb(n20746), .dout(n20748));
  jand g20621(.dina(n16604), .dinb(n1806), .dout(n20749));
  jor  g20622(.dina(n20749), .dinb(n20748), .dout(n20750));
  jor  g20623(.dina(n20750), .dinb(n20745), .dout(n20751));
  jxor g20624(.dina(n20751), .dinb(n77), .dout(n20752));
  jxor g20625(.dina(n20752), .dinb(n20744), .dout(n20753));
  jxor g20626(.dina(n20753), .dinb(n20696), .dout(n20754));
  jnot g20627(.din(n20754), .dout(n20755));
  jand g20628(.dina(n17944), .dinb(n806), .dout(n20756));
  jand g20629(.dina(n17535), .dinb(n1612), .dout(n20757));
  jand g20630(.dina(n17942), .dinb(n1620), .dout(n20758));
  jor  g20631(.dina(n20758), .dinb(n20757), .dout(n20759));
  jand g20632(.dina(n17329), .dinb(n1644), .dout(n20760));
  jor  g20633(.dina(n20760), .dinb(n20759), .dout(n20761));
  jor  g20634(.dina(n20761), .dinb(n20756), .dout(n20762));
  jxor g20635(.dina(n20762), .dinb(n65), .dout(n20763));
  jxor g20636(.dina(n20763), .dinb(n20755), .dout(n20764));
  jxor g20637(.dina(n20764), .dinb(n20691), .dout(n20765));
  jnot g20638(.din(n20765), .dout(n20766));
  jand g20639(.dina(n18490), .dinb(n1819), .dout(n20767));
  jand g20640(.dina(n18488), .dinb(n2243), .dout(n20768));
  jand g20641(.dina(n18292), .dinb(n2180), .dout(n20769));
  jand g20642(.dina(n18293), .dinb(n2185), .dout(n20770));
  jor  g20643(.dina(n20770), .dinb(n20769), .dout(n20771));
  jor  g20644(.dina(n20771), .dinb(n20768), .dout(n20772));
  jor  g20645(.dina(n20772), .dinb(n20767), .dout(n20773));
  jxor g20646(.dina(n20773), .dinb(n2196), .dout(n20774));
  jxor g20647(.dina(n20774), .dinb(n20766), .dout(n20775));
  jxor g20648(.dina(n20775), .dinb(n20686), .dout(n20776));
  jnot g20649(.din(n20776), .dout(n20777));
  jand g20650(.dina(n19387), .dinb(n2743), .dout(n20778));
  jand g20651(.dina(n19219), .dinb(n2752), .dout(n20779));
  jand g20652(.dina(n19220), .dinb(n2748), .dout(n20780));
  jand g20653(.dina(n18914), .dinb(n2757), .dout(n20781));
  jor  g20654(.dina(n20781), .dinb(n20780), .dout(n20782));
  jor  g20655(.dina(n20782), .dinb(n20779), .dout(n20783));
  jor  g20656(.dina(n20783), .dinb(n20778), .dout(n20784));
  jxor g20657(.dina(n20784), .dinb(n2441), .dout(n20785));
  jxor g20658(.dina(n20785), .dinb(n20777), .dout(n20786));
  jxor g20659(.dina(n20786), .dinb(n20681), .dout(n20787));
  jnot g20660(.din(n20787), .dout(n20788));
  jand g20661(.dina(n20371), .dinb(n3423), .dout(n20789));
  jand g20662(.dina(n19922), .dinb(n3428), .dout(n20790));
  jand g20663(.dina(n20205), .dinb(n3569), .dout(n20791));
  jor  g20664(.dina(n20791), .dinb(n20790), .dout(n20792));
  jand g20665(.dina(n19373), .dinb(n3210), .dout(n20793));
  jor  g20666(.dina(n20793), .dinb(n20792), .dout(n20794));
  jor  g20667(.dina(n20794), .dinb(n20789), .dout(n20795));
  jxor g20668(.dina(n20795), .dinb(n3473), .dout(n20796));
  jxor g20669(.dina(n20796), .dinb(n20788), .dout(n20797));
  jxor g20670(.dina(n20797), .dinb(n20678), .dout(n20798));
  jand g20671(.dina(n20344), .dinb(n20204), .dout(n20799));
  jand g20672(.dina(n20345), .dinb(n20216), .dout(n20800));
  jor  g20673(.dina(n20800), .dinb(n20799), .dout(n20801));
  jand g20674(.dina(n20341), .dinb(n20224), .dout(n20802));
  jnot g20675(.din(n20802), .dout(n20803));
  jor  g20676(.dina(n20343), .dinb(n20220), .dout(n20804));
  jand g20677(.dina(n20804), .dinb(n20803), .dout(n20805));
  jor  g20678(.dina(n20339), .dinb(n20331), .dout(n20806));
  jnot g20679(.din(n20806), .dout(n20807));
  jand g20680(.dina(n20340), .dinb(n20327), .dout(n20808));
  jor  g20681(.dina(n20808), .dinb(n20807), .dout(n20809));
  jor  g20682(.dina(n20325), .dinb(n20317), .dout(n20810));
  jand g20683(.dina(n20326), .dinb(n20230), .dout(n20811));
  jnot g20684(.din(n20811), .dout(n20812));
  jand g20685(.dina(n20812), .dinb(n20810), .dout(n20813));
  jor  g20686(.dina(n20314), .dinb(n20306), .dout(n20814));
  jand g20687(.dina(n20315), .dinb(n20235), .dout(n20815));
  jnot g20688(.din(n20815), .dout(n20816));
  jand g20689(.dina(n20816), .dinb(n20814), .dout(n20817));
  jnot g20690(.din(n20817), .dout(n20818));
  jor  g20691(.dina(n20303), .dinb(n20295), .dout(n20819));
  jand g20692(.dina(n20304), .dinb(n20239), .dout(n20820));
  jnot g20693(.din(n20820), .dout(n20821));
  jand g20694(.dina(n20821), .dinb(n20819), .dout(n20822));
  jnot g20695(.din(n20822), .dout(n20823));
  jor  g20696(.dina(n20292), .dinb(n20284), .dout(n20824));
  jand g20697(.dina(n20293), .dinb(n20244), .dout(n20825));
  jnot g20698(.din(n20825), .dout(n20826));
  jand g20699(.dina(n20826), .dinb(n20824), .dout(n20827));
  jnot g20700(.din(n20827), .dout(n20828));
  jand g20701(.dina(n20281), .dinb(n20256), .dout(n20829));
  jand g20702(.dina(n20282), .dinb(n20251), .dout(n20830));
  jor  g20703(.dina(n20830), .dinb(n20829), .dout(n20831));
  jand g20704(.dina(n9756), .dinb(n1378), .dout(n20832));
  jand g20705(.dina(n20832), .dinb(n534), .dout(n20833));
  jand g20706(.dina(n20833), .dinb(n9129), .dout(n20834));
  jand g20707(.dina(n1465), .dinb(n1375), .dout(n20835));
  jand g20708(.dina(n20835), .dinb(n20834), .dout(n20836));
  jnot g20709(.din(n889), .dout(n20837));
  jand g20710(.dina(n881), .dinb(n440), .dout(n20838));
  jand g20711(.dina(n20838), .dinb(n1212), .dout(n20839));
  jand g20712(.dina(n1731), .dinb(n114), .dout(n20840));
  jand g20713(.dina(n20840), .dinb(n1205), .dout(n20841));
  jand g20714(.dina(n20841), .dinb(n20839), .dout(n20842));
  jand g20715(.dina(n20842), .dinb(n20837), .dout(n20843));
  jand g20716(.dina(n3758), .dinb(n452), .dout(n20844));
  jand g20717(.dina(n20844), .dinb(n17823), .dout(n20845));
  jand g20718(.dina(n20845), .dinb(n553), .dout(n20846));
  jand g20719(.dina(n20846), .dinb(n20843), .dout(n20847));
  jand g20720(.dina(n20847), .dinb(n11192), .dout(n20848));
  jand g20721(.dina(n20848), .dinb(n20836), .dout(n20849));
  jand g20722(.dina(n1096), .dinb(n673), .dout(n20850));
  jand g20723(.dina(n20850), .dinb(n20849), .dout(n20851));
  jand g20724(.dina(n1226), .dinb(n653), .dout(n20852));
  jand g20725(.dina(n693), .dinb(n600), .dout(n20853));
  jand g20726(.dina(n20853), .dinb(n20852), .dout(n20854));
  jand g20727(.dina(n20854), .dinb(n1898), .dout(n20855));
  jand g20728(.dina(n20855), .dinb(n9373), .dout(n20856));
  jand g20729(.dina(n1190), .dinb(n499), .dout(n20857));
  jand g20730(.dina(n833), .dinb(n908), .dout(n20858));
  jand g20731(.dina(n20858), .dinb(n6270), .dout(n20859));
  jand g20732(.dina(n1289), .dinb(n179), .dout(n20860));
  jand g20733(.dina(n20860), .dinb(n20859), .dout(n20861));
  jand g20734(.dina(n1524), .dinb(n641), .dout(n20862));
  jand g20735(.dina(n20862), .dinb(n549), .dout(n20863));
  jand g20736(.dina(n20863), .dinb(n20861), .dout(n20864));
  jand g20737(.dina(n20864), .dinb(n20857), .dout(n20865));
  jand g20738(.dina(n3276), .dinb(n3136), .dout(n20866));
  jand g20739(.dina(n1168), .dinb(n504), .dout(n20867));
  jand g20740(.dina(n20867), .dinb(n20866), .dout(n20868));
  jand g20741(.dina(n703), .dinb(n1233), .dout(n20869));
  jand g20742(.dina(n20869), .dinb(n869), .dout(n20870));
  jand g20743(.dina(n20870), .dinb(n2650), .dout(n20871));
  jand g20744(.dina(n20871), .dinb(n20868), .dout(n20872));
  jand g20745(.dina(n20872), .dinb(n20865), .dout(n20873));
  jand g20746(.dina(n20873), .dinb(n20856), .dout(n20874));
  jand g20747(.dina(n20874), .dinb(n1341), .dout(n20875));
  jand g20748(.dina(n20875), .dinb(n20851), .dout(n20876));
  jnot g20749(.din(n20876), .dout(n20877));
  jor  g20750(.dina(n20275), .dinb(n19974), .dout(n20878));
  jand g20751(.dina(n20280), .dinb(n20276), .dout(n20879));
  jnot g20752(.din(n20879), .dout(n20880));
  jand g20753(.dina(n20880), .dinb(n20878), .dout(n20881));
  jxor g20754(.dina(n20881), .dinb(n20877), .dout(n20882));
  jand g20755(.dina(n13250), .dinb(n5076), .dout(n20883));
  jand g20756(.dina(n13248), .dinb(n5084), .dout(n20884));
  jand g20757(.dina(n12536), .dinb(n6050), .dout(n20885));
  jand g20758(.dina(n12669), .dinb(n5082), .dout(n20886));
  jor  g20759(.dina(n20886), .dinb(n20885), .dout(n20887));
  jor  g20760(.dina(n20887), .dinb(n20884), .dout(n20888));
  jor  g20761(.dina(n20888), .dinb(n20883), .dout(n20889));
  jxor g20762(.dina(n20889), .dinb(n20882), .dout(n20890));
  jxor g20763(.dina(n20890), .dinb(n20831), .dout(n20891));
  jnot g20764(.din(n20891), .dout(n20892));
  jand g20765(.dina(n13616), .dinb(n2936), .dout(n20893));
  jand g20766(.dina(n13469), .dinb(n2940), .dout(n20894));
  jand g20767(.dina(n13614), .dinb(n2943), .dout(n20895));
  jor  g20768(.dina(n20895), .dinb(n20894), .dout(n20896));
  jand g20769(.dina(n13478), .dinb(n3684), .dout(n20897));
  jor  g20770(.dina(n20897), .dinb(n20896), .dout(n20898));
  jor  g20771(.dina(n20898), .dinb(n20893), .dout(n20899));
  jxor g20772(.dina(n20899), .dinb(n93), .dout(n20900));
  jxor g20773(.dina(n20900), .dinb(n20892), .dout(n20901));
  jxor g20774(.dina(n20901), .dinb(n20828), .dout(n20902));
  jnot g20775(.din(n20902), .dout(n20903));
  jand g20776(.dina(n14562), .dinb(n71), .dout(n20904));
  jand g20777(.dina(n14447), .dinb(n796), .dout(n20905));
  jand g20778(.dina(n14448), .dinb(n731), .dout(n20906));
  jand g20779(.dina(n14249), .dinb(n1806), .dout(n20907));
  jor  g20780(.dina(n20907), .dinb(n20906), .dout(n20908));
  jor  g20781(.dina(n20908), .dinb(n20905), .dout(n20909));
  jor  g20782(.dina(n20909), .dinb(n20904), .dout(n20910));
  jxor g20783(.dina(n20910), .dinb(n77), .dout(n20911));
  jxor g20784(.dina(n20911), .dinb(n20903), .dout(n20912));
  jxor g20785(.dina(n20912), .dinb(n20823), .dout(n20913));
  jnot g20786(.din(n20913), .dout(n20914));
  jand g20787(.dina(n15569), .dinb(n806), .dout(n20915));
  jand g20788(.dina(n15567), .dinb(n1620), .dout(n20916));
  jand g20789(.dina(n15315), .dinb(n1612), .dout(n20917));
  jand g20790(.dina(n14549), .dinb(n1644), .dout(n20918));
  jor  g20791(.dina(n20918), .dinb(n20917), .dout(n20919));
  jor  g20792(.dina(n20919), .dinb(n20916), .dout(n20920));
  jor  g20793(.dina(n20920), .dinb(n20915), .dout(n20921));
  jxor g20794(.dina(n20921), .dinb(n65), .dout(n20922));
  jxor g20795(.dina(n20922), .dinb(n20914), .dout(n20923));
  jxor g20796(.dina(n20923), .dinb(n20818), .dout(n20924));
  jnot g20797(.din(n20924), .dout(n20925));
  jand g20798(.dina(n16345), .dinb(n1819), .dout(n20926));
  jand g20799(.dina(n16082), .dinb(n2180), .dout(n20927));
  jand g20800(.dina(n16343), .dinb(n2243), .dout(n20928));
  jor  g20801(.dina(n20928), .dinb(n20927), .dout(n20929));
  jand g20802(.dina(n15829), .dinb(n2185), .dout(n20930));
  jor  g20803(.dina(n20930), .dinb(n20929), .dout(n20931));
  jor  g20804(.dina(n20931), .dinb(n20926), .dout(n20932));
  jxor g20805(.dina(n20932), .dinb(n2196), .dout(n20933));
  jxor g20806(.dina(n20933), .dinb(n20925), .dout(n20934));
  jxor g20807(.dina(n20934), .dinb(n20813), .dout(n20935));
  jand g20808(.dina(n17312), .dinb(n2743), .dout(n20936));
  jand g20809(.dina(n16928), .dinb(n2748), .dout(n20937));
  jand g20810(.dina(n16592), .dinb(n2757), .dout(n20938));
  jand g20811(.dina(n16924), .dinb(n2752), .dout(n20939));
  jor  g20812(.dina(n20939), .dinb(n20938), .dout(n20940));
  jor  g20813(.dina(n20940), .dinb(n20937), .dout(n20941));
  jor  g20814(.dina(n20941), .dinb(n20936), .dout(n20942));
  jxor g20815(.dina(n20942), .dinb(n2441), .dout(n20943));
  jxor g20816(.dina(n20943), .dinb(n20935), .dout(n20944));
  jxor g20817(.dina(n20944), .dinb(n20809), .dout(n20945));
  jnot g20818(.din(n20945), .dout(n20946));
  jxor g20819(.dina(n20946), .dinb(n20805), .dout(n20947));
  jxor g20820(.dina(n20947), .dinb(n20344), .dout(n20948));
  jxor g20821(.dina(n20948), .dinb(n20801), .dout(n20949));
  jand g20822(.dina(n20949), .dinb(n4022), .dout(n20950));
  jand g20823(.dina(n20344), .dinb(n4027), .dout(n20951));
  jand g20824(.dina(n20947), .dinb(n4220), .dout(n20952));
  jor  g20825(.dina(n20952), .dinb(n20951), .dout(n20953));
  jand g20826(.dina(n20204), .dinb(n3870), .dout(n20954));
  jor  g20827(.dina(n20954), .dinb(n20953), .dout(n20955));
  jor  g20828(.dina(n20955), .dinb(n20950), .dout(n20956));
  jxor g20829(.dina(n20956), .dinb(n4050), .dout(n20957));
  jxor g20830(.dina(n20957), .dinb(n20798), .dout(n20958));
  jxor g20831(.dina(n20958), .dinb(n20674), .dout(n20959));
  jnot g20832(.din(n20813), .dout(n20960));
  jand g20833(.dina(n20934), .dinb(n20960), .dout(n20961));
  jor  g20834(.dina(n20943), .dinb(n20935), .dout(n20962));
  jnot g20835(.din(n20962), .dout(n20963));
  jor  g20836(.dina(n20963), .dinb(n20961), .dout(n20964));
  jand g20837(.dina(n20923), .dinb(n20818), .dout(n20965));
  jnot g20838(.din(n20965), .dout(n20966));
  jor  g20839(.dina(n20933), .dinb(n20925), .dout(n20967));
  jand g20840(.dina(n20967), .dinb(n20966), .dout(n20968));
  jand g20841(.dina(n2753), .dinb(n2749), .dout(n20969));
  jor  g20842(.dina(n20969), .dinb(n17301), .dout(n20970));
  jor  g20843(.dina(n17296), .dinb(n2744), .dout(n20971));
  jor  g20844(.dina(n17288), .dinb(n2758), .dout(n20972));
  jand g20845(.dina(n20972), .dinb(n20971), .dout(n20973));
  jand g20846(.dina(n20973), .dinb(n20970), .dout(n20974));
  jxor g20847(.dina(n20974), .dinb(\a[17] ), .dout(n20975));
  jxor g20848(.dina(n20975), .dinb(n20968), .dout(n20976));
  jand g20849(.dina(n20912), .dinb(n20823), .dout(n20977));
  jnot g20850(.din(n20977), .dout(n20978));
  jor  g20851(.dina(n20922), .dinb(n20914), .dout(n20979));
  jand g20852(.dina(n20979), .dinb(n20978), .dout(n20980));
  jnot g20853(.din(n20980), .dout(n20981));
  jand g20854(.dina(n20901), .dinb(n20828), .dout(n20982));
  jnot g20855(.din(n20982), .dout(n20983));
  jor  g20856(.dina(n20911), .dinb(n20903), .dout(n20984));
  jand g20857(.dina(n20984), .dinb(n20983), .dout(n20985));
  jnot g20858(.din(n20985), .dout(n20986));
  jand g20859(.dina(n20890), .dinb(n20831), .dout(n20987));
  jnot g20860(.din(n20987), .dout(n20988));
  jor  g20861(.dina(n20900), .dinb(n20892), .dout(n20989));
  jand g20862(.dina(n20989), .dinb(n20988), .dout(n20990));
  jnot g20863(.din(n20990), .dout(n20991));
  jand g20864(.dina(n13639), .dinb(n5076), .dout(n20992));
  jand g20865(.dina(n13478), .dinb(n5084), .dout(n20993));
  jand g20866(.dina(n13248), .dinb(n5082), .dout(n20994));
  jand g20867(.dina(n12669), .dinb(n6050), .dout(n20995));
  jor  g20868(.dina(n20995), .dinb(n20994), .dout(n20996));
  jor  g20869(.dina(n20996), .dinb(n20993), .dout(n20997));
  jor  g20870(.dina(n20997), .dinb(n20992), .dout(n20998));
  jor  g20871(.dina(n20881), .dinb(n20877), .dout(n20999));
  jand g20872(.dina(n20889), .dinb(n20882), .dout(n21000));
  jnot g20873(.din(n21000), .dout(n21001));
  jand g20874(.dina(n21001), .dinb(n20999), .dout(n21002));
  jnot g20875(.din(n21002), .dout(n21003));
  jand g20876(.dina(n1571), .dinb(n450), .dout(n21004));
  jand g20877(.dina(n325), .dinb(n1288), .dout(n21005));
  jand g20878(.dina(n21005), .dinb(n8580), .dout(n21006));
  jand g20879(.dina(n21006), .dinb(n2094), .dout(n21007));
  jand g20880(.dina(n21007), .dinb(n1462), .dout(n21008));
  jand g20881(.dina(n21008), .dinb(n21004), .dout(n21009));
  jand g20882(.dina(n21009), .dinb(n10152), .dout(n21010));
  jand g20883(.dina(n21010), .dinb(n2007), .dout(n21011));
  jand g20884(.dina(n1936), .dinb(n621), .dout(n21012));
  jand g20885(.dina(n15656), .dinb(n2511), .dout(n21013));
  jand g20886(.dina(n21013), .dinb(n21012), .dout(n21014));
  jand g20887(.dina(n3007), .dinb(n1559), .dout(n21015));
  jand g20888(.dina(n21015), .dinb(n1310), .dout(n21016));
  jand g20889(.dina(n21016), .dinb(n21014), .dout(n21017));
  jand g20890(.dina(n537), .dinb(n1344), .dout(n21018));
  jand g20891(.dina(n1713), .dinb(n929), .dout(n21019));
  jand g20892(.dina(n21019), .dinb(n21018), .dout(n21020));
  jand g20893(.dina(n1506), .dinb(n871), .dout(n21021));
  jand g20894(.dina(n21021), .dinb(n1374), .dout(n21022));
  jand g20895(.dina(n21022), .dinb(n21020), .dout(n21023));
  jand g20896(.dina(n21023), .dinb(n697), .dout(n21024));
  jand g20897(.dina(n21024), .dinb(n21017), .dout(n21025));
  jand g20898(.dina(n21025), .dinb(n12465), .dout(n21026));
  jand g20899(.dina(n21026), .dinb(n21011), .dout(n21027));
  jxor g20900(.dina(n21027), .dinb(n20877), .dout(n21028));
  jxor g20901(.dina(n21028), .dinb(n21003), .dout(n21029));
  jxor g20902(.dina(n21029), .dinb(n20998), .dout(n21030));
  jnot g20903(.din(n21030), .dout(n21031));
  jand g20904(.dina(n14251), .dinb(n2936), .dout(n21032));
  jand g20905(.dina(n14249), .dinb(n2943), .dout(n21033));
  jand g20906(.dina(n13614), .dinb(n2940), .dout(n21034));
  jand g20907(.dina(n13469), .dinb(n3684), .dout(n21035));
  jor  g20908(.dina(n21035), .dinb(n21034), .dout(n21036));
  jor  g20909(.dina(n21036), .dinb(n21033), .dout(n21037));
  jor  g20910(.dina(n21037), .dinb(n21032), .dout(n21038));
  jxor g20911(.dina(n21038), .dinb(n93), .dout(n21039));
  jxor g20912(.dina(n21039), .dinb(n21031), .dout(n21040));
  jxor g20913(.dina(n21040), .dinb(n20991), .dout(n21041));
  jnot g20914(.din(n21041), .dout(n21042));
  jand g20915(.dina(n14551), .dinb(n71), .dout(n21043));
  jand g20916(.dina(n14447), .dinb(n731), .dout(n21044));
  jand g20917(.dina(n14549), .dinb(n796), .dout(n21045));
  jor  g20918(.dina(n21045), .dinb(n21044), .dout(n21046));
  jand g20919(.dina(n14448), .dinb(n1806), .dout(n21047));
  jor  g20920(.dina(n21047), .dinb(n21046), .dout(n21048));
  jor  g20921(.dina(n21048), .dinb(n21043), .dout(n21049));
  jxor g20922(.dina(n21049), .dinb(n77), .dout(n21050));
  jxor g20923(.dina(n21050), .dinb(n21042), .dout(n21051));
  jxor g20924(.dina(n21051), .dinb(n20986), .dout(n21052));
  jnot g20925(.din(n21052), .dout(n21053));
  jand g20926(.dina(n15831), .dinb(n806), .dout(n21054));
  jand g20927(.dina(n15567), .dinb(n1612), .dout(n21055));
  jand g20928(.dina(n15829), .dinb(n1620), .dout(n21056));
  jor  g20929(.dina(n21056), .dinb(n21055), .dout(n21057));
  jand g20930(.dina(n15315), .dinb(n1644), .dout(n21058));
  jor  g20931(.dina(n21058), .dinb(n21057), .dout(n21059));
  jor  g20932(.dina(n21059), .dinb(n21054), .dout(n21060));
  jxor g20933(.dina(n21060), .dinb(n65), .dout(n21061));
  jxor g20934(.dina(n21061), .dinb(n21053), .dout(n21062));
  jxor g20935(.dina(n21062), .dinb(n20981), .dout(n21063));
  jnot g20936(.din(n21063), .dout(n21064));
  jand g20937(.dina(n16594), .dinb(n1819), .dout(n21065));
  jand g20938(.dina(n16592), .dinb(n2243), .dout(n21066));
  jand g20939(.dina(n16343), .dinb(n2180), .dout(n21067));
  jand g20940(.dina(n16082), .dinb(n2185), .dout(n21068));
  jor  g20941(.dina(n21068), .dinb(n21067), .dout(n21069));
  jor  g20942(.dina(n21069), .dinb(n21066), .dout(n21070));
  jor  g20943(.dina(n21070), .dinb(n21065), .dout(n21071));
  jxor g20944(.dina(n21071), .dinb(n2196), .dout(n21072));
  jxor g20945(.dina(n21072), .dinb(n21064), .dout(n21073));
  jxor g20946(.dina(n21073), .dinb(n20976), .dout(n21074));
  jand g20947(.dina(n21074), .dinb(n20964), .dout(n21075));
  jnot g20948(.din(n21075), .dout(n21076));
  jxor g20949(.dina(n21074), .dinb(n20964), .dout(n21077));
  jnot g20950(.din(n21077), .dout(n21078));
  jand g20951(.dina(n20944), .dinb(n20809), .dout(n21079));
  jnot g20952(.din(n21079), .dout(n21080));
  jor  g20953(.dina(n20946), .dinb(n20805), .dout(n21081));
  jand g20954(.dina(n21081), .dinb(n21080), .dout(n21082));
  jor  g20955(.dina(n21082), .dinb(n21078), .dout(n21083));
  jand g20956(.dina(n21083), .dinb(n21076), .dout(n21084));
  jor  g20957(.dina(n20975), .dinb(n20968), .dout(n21085));
  jand g20958(.dina(n21073), .dinb(n20976), .dout(n21086));
  jnot g20959(.din(n21086), .dout(n21087));
  jand g20960(.dina(n21087), .dinb(n21085), .dout(n21088));
  jnot g20961(.din(n21088), .dout(n21089));
  jand g20962(.dina(n21051), .dinb(n20986), .dout(n21090));
  jnot g20963(.din(n21090), .dout(n21091));
  jor  g20964(.dina(n21061), .dinb(n21053), .dout(n21092));
  jand g20965(.dina(n21092), .dinb(n21091), .dout(n21093));
  jnot g20966(.din(n21093), .dout(n21094));
  jand g20967(.dina(n21040), .dinb(n20991), .dout(n21095));
  jnot g20968(.din(n21095), .dout(n21096));
  jor  g20969(.dina(n21050), .dinb(n21042), .dout(n21097));
  jand g20970(.dina(n21097), .dinb(n21096), .dout(n21098));
  jnot g20971(.din(n21098), .dout(n21099));
  jand g20972(.dina(n21029), .dinb(n20998), .dout(n21100));
  jnot g20973(.din(n21100), .dout(n21101));
  jor  g20974(.dina(n21039), .dinb(n21031), .dout(n21102));
  jand g20975(.dina(n21102), .dinb(n21101), .dout(n21103));
  jnot g20976(.din(n21103), .dout(n21104));
  jand g20977(.dina(n21027), .dinb(n20877), .dout(n21105));
  jand g20978(.dina(n21028), .dinb(n21003), .dout(n21106));
  jor  g20979(.dina(n21106), .dinb(n21105), .dout(n21107));
  jand g20980(.dina(n13627), .dinb(n5076), .dout(n21108));
  jand g20981(.dina(n13469), .dinb(n5084), .dout(n21109));
  jand g20982(.dina(n13478), .dinb(n5082), .dout(n21110));
  jand g20983(.dina(n13248), .dinb(n6050), .dout(n21111));
  jor  g20984(.dina(n21111), .dinb(n21110), .dout(n21112));
  jor  g20985(.dina(n21112), .dinb(n21109), .dout(n21113));
  jor  g20986(.dina(n21113), .dinb(n21108), .dout(n21114));
  jand g20987(.dina(n11381), .dinb(n137), .dout(n21115));
  jand g20988(.dina(n10388), .dinb(n686), .dout(n21116));
  jand g20989(.dina(n1219), .dinb(n1437), .dout(n21117));
  jand g20990(.dina(n21117), .dinb(n3238), .dout(n21118));
  jand g20991(.dina(n21118), .dinb(n1532), .dout(n21119));
  jand g20992(.dina(n13403), .dinb(n5379), .dout(n21120));
  jand g20993(.dina(n21120), .dinb(n838), .dout(n21121));
  jand g20994(.dina(n21121), .dinb(n21119), .dout(n21122));
  jand g20995(.dina(n21122), .dinb(n21116), .dout(n21123));
  jand g20996(.dina(n1744), .dinb(n1304), .dout(n21124));
  jand g20997(.dina(n21124), .dinb(n2148), .dout(n21125));
  jand g20998(.dina(n3276), .dinb(n326), .dout(n21126));
  jand g20999(.dina(n7518), .dinb(n1763), .dout(n21127));
  jand g21000(.dina(n21127), .dinb(n21126), .dout(n21128));
  jand g21001(.dina(n21128), .dinb(n21125), .dout(n21129));
  jand g21002(.dina(n21129), .dinb(n21123), .dout(n21130));
  jand g21003(.dina(n21130), .dinb(n15280), .dout(n21131));
  jand g21004(.dina(n18376), .dinb(n1522), .dout(n21132));
  jand g21005(.dina(n1203), .dinb(n933), .dout(n21133));
  jand g21006(.dina(n21133), .dinb(n1288), .dout(n21134));
  jand g21007(.dina(n21134), .dinb(n469), .dout(n21135));
  jand g21008(.dina(n21135), .dinb(n21132), .dout(n21136));
  jand g21009(.dina(n21136), .dinb(n1183), .dout(n21137));
  jand g21010(.dina(n21137), .dinb(n1453), .dout(n21138));
  jand g21011(.dina(n21138), .dinb(n21131), .dout(n21139));
  jand g21012(.dina(n21139), .dinb(n21115), .dout(n21140));
  jxor g21013(.dina(n21140), .dinb(n21027), .dout(n21141));
  jand g21014(.dina(n2756), .dinb(n2751), .dout(n21142));
  jor  g21015(.dina(n21142), .dinb(n17301), .dout(n21143));
  jxor g21016(.dina(n21143), .dinb(\a[17] ), .dout(n21144));
  jxor g21017(.dina(n21144), .dinb(n21141), .dout(n21145));
  jxor g21018(.dina(n21145), .dinb(n21114), .dout(n21146));
  jxor g21019(.dina(n21146), .dinb(n21107), .dout(n21147));
  jxor g21020(.dina(n21147), .dinb(n21104), .dout(n21148));
  jnot g21021(.din(n21148), .dout(n21149));
  jand g21022(.dina(n14579), .dinb(n2936), .dout(n21150));
  jand g21023(.dina(n14249), .dinb(n2940), .dout(n21151));
  jand g21024(.dina(n14448), .dinb(n2943), .dout(n21152));
  jor  g21025(.dina(n21152), .dinb(n21151), .dout(n21153));
  jand g21026(.dina(n13614), .dinb(n3684), .dout(n21154));
  jor  g21027(.dina(n21154), .dinb(n21153), .dout(n21155));
  jor  g21028(.dina(n21155), .dinb(n21150), .dout(n21156));
  jxor g21029(.dina(n21156), .dinb(n93), .dout(n21157));
  jxor g21030(.dina(n21157), .dinb(n21149), .dout(n21158));
  jnot g21031(.din(n21158), .dout(n21159));
  jand g21032(.dina(n15317), .dinb(n71), .dout(n21160));
  jand g21033(.dina(n14549), .dinb(n731), .dout(n21161));
  jand g21034(.dina(n15315), .dinb(n796), .dout(n21162));
  jor  g21035(.dina(n21162), .dinb(n21161), .dout(n21163));
  jand g21036(.dina(n14447), .dinb(n1806), .dout(n21164));
  jor  g21037(.dina(n21164), .dinb(n21163), .dout(n21165));
  jor  g21038(.dina(n21165), .dinb(n21160), .dout(n21166));
  jxor g21039(.dina(n21166), .dinb(n77), .dout(n21167));
  jxor g21040(.dina(n21167), .dinb(n21159), .dout(n21168));
  jxor g21041(.dina(n21168), .dinb(n21099), .dout(n21169));
  jnot g21042(.din(n21169), .dout(n21170));
  jand g21043(.dina(n16084), .dinb(n806), .dout(n21171));
  jand g21044(.dina(n15829), .dinb(n1612), .dout(n21172));
  jand g21045(.dina(n16082), .dinb(n1620), .dout(n21173));
  jor  g21046(.dina(n21173), .dinb(n21172), .dout(n21174));
  jand g21047(.dina(n15567), .dinb(n1644), .dout(n21175));
  jor  g21048(.dina(n21175), .dinb(n21174), .dout(n21176));
  jor  g21049(.dina(n21176), .dinb(n21171), .dout(n21177));
  jxor g21050(.dina(n21177), .dinb(n65), .dout(n21178));
  jxor g21051(.dina(n21178), .dinb(n21170), .dout(n21179));
  jxor g21052(.dina(n21179), .dinb(n21094), .dout(n21180));
  jand g21053(.dina(n21062), .dinb(n20981), .dout(n21181));
  jnot g21054(.din(n21181), .dout(n21182));
  jor  g21055(.dina(n21072), .dinb(n21064), .dout(n21183));
  jand g21056(.dina(n21183), .dinb(n21182), .dout(n21184));
  jand g21057(.dina(n16930), .dinb(n1819), .dout(n21185));
  jand g21058(.dina(n16592), .dinb(n2180), .dout(n21186));
  jand g21059(.dina(n16928), .dinb(n2243), .dout(n21187));
  jor  g21060(.dina(n21187), .dinb(n21186), .dout(n21188));
  jand g21061(.dina(n16343), .dinb(n2185), .dout(n21189));
  jor  g21062(.dina(n21189), .dinb(n21188), .dout(n21190));
  jor  g21063(.dina(n21190), .dinb(n21185), .dout(n21191));
  jxor g21064(.dina(n21191), .dinb(n2196), .dout(n21192));
  jxor g21065(.dina(n21192), .dinb(n21184), .dout(n21193));
  jxor g21066(.dina(n21193), .dinb(n21180), .dout(n21194));
  jxor g21067(.dina(n21194), .dinb(n21089), .dout(n21195));
  jnot g21068(.din(n21195), .dout(n21196));
  jxor g21069(.dina(n21196), .dinb(n21084), .dout(n21197));
  jxor g21070(.dina(n21082), .dinb(n21078), .dout(n21198));
  jand g21071(.dina(n21198), .dinb(n21197), .dout(n21199));
  jand g21072(.dina(n21198), .dinb(n20947), .dout(n21200));
  jand g21073(.dina(n20947), .dinb(n20344), .dout(n21201));
  jand g21074(.dina(n20948), .dinb(n20801), .dout(n21202));
  jor  g21075(.dina(n21202), .dinb(n21201), .dout(n21203));
  jxor g21076(.dina(n21198), .dinb(n20947), .dout(n21204));
  jand g21077(.dina(n21204), .dinb(n21203), .dout(n21205));
  jor  g21078(.dina(n21205), .dinb(n21200), .dout(n21206));
  jxor g21079(.dina(n21198), .dinb(n21197), .dout(n21207));
  jand g21080(.dina(n21207), .dinb(n21206), .dout(n21208));
  jor  g21081(.dina(n21208), .dinb(n21199), .dout(n21209));
  jand g21082(.dina(n21194), .dinb(n21089), .dout(n21210));
  jnot g21083(.din(n21210), .dout(n21211));
  jor  g21084(.dina(n21196), .dinb(n21084), .dout(n21212));
  jand g21085(.dina(n21212), .dinb(n21211), .dout(n21213));
  jor  g21086(.dina(n21192), .dinb(n21184), .dout(n21214));
  jand g21087(.dina(n21193), .dinb(n21180), .dout(n21215));
  jnot g21088(.din(n21215), .dout(n21216));
  jand g21089(.dina(n21216), .dinb(n21214), .dout(n21217));
  jnot g21090(.din(n21217), .dout(n21218));
  jor  g21091(.dina(n21178), .dinb(n21170), .dout(n21219));
  jand g21092(.dina(n21179), .dinb(n21094), .dout(n21220));
  jnot g21093(.din(n21220), .dout(n21221));
  jand g21094(.dina(n21221), .dinb(n21219), .dout(n21222));
  jnot g21095(.din(n21222), .dout(n21223));
  jor  g21096(.dina(n21167), .dinb(n21159), .dout(n21224));
  jand g21097(.dina(n21168), .dinb(n21099), .dout(n21225));
  jnot g21098(.din(n21225), .dout(n21226));
  jand g21099(.dina(n21226), .dinb(n21224), .dout(n21227));
  jnot g21100(.din(n21227), .dout(n21228));
  jand g21101(.dina(n21147), .dinb(n21104), .dout(n21229));
  jnot g21102(.din(n21229), .dout(n21230));
  jor  g21103(.dina(n21157), .dinb(n21149), .dout(n21231));
  jand g21104(.dina(n21231), .dinb(n21230), .dout(n21232));
  jnot g21105(.din(n21232), .dout(n21233));
  jand g21106(.dina(n21145), .dinb(n21114), .dout(n21234));
  jand g21107(.dina(n21146), .dinb(n21107), .dout(n21235));
  jor  g21108(.dina(n21235), .dinb(n21234), .dout(n21236));
  jand g21109(.dina(n654), .dinb(n1283), .dout(n21237));
  jand g21110(.dina(n21237), .dinb(n1317), .dout(n21238));
  jand g21111(.dina(n5408), .dinb(n699), .dout(n21239));
  jand g21112(.dina(n21239), .dinb(n1326), .dout(n21240));
  jand g21113(.dina(n21240), .dinb(n21238), .dout(n21241));
  jand g21114(.dina(n1522), .dinb(n1559), .dout(n21242));
  jand g21115(.dina(n21242), .dinb(n3779), .dout(n21243));
  jand g21116(.dina(n21243), .dinb(n270), .dout(n21244));
  jand g21117(.dina(n1721), .dinb(n622), .dout(n21245));
  jand g21118(.dina(n21245), .dinb(n21244), .dout(n21246));
  jand g21119(.dina(n8355), .dinb(n1328), .dout(n21247));
  jand g21120(.dina(n21247), .dinb(n21246), .dout(n21248));
  jand g21121(.dina(n7088), .dinb(n583), .dout(n21249));
  jand g21122(.dina(n908), .dinb(n1316), .dout(n21250));
  jand g21123(.dina(n21250), .dinb(n2394), .dout(n21251));
  jand g21124(.dina(n21251), .dinb(n21249), .dout(n21252));
  jand g21125(.dina(n4617), .dinb(n1453), .dout(n21253));
  jand g21126(.dina(n21253), .dinb(n1272), .dout(n21254));
  jand g21127(.dina(n21254), .dinb(n21252), .dout(n21255));
  jand g21128(.dina(n10398), .dinb(n1855), .dout(n21256));
  jand g21129(.dina(n21256), .dinb(n21255), .dout(n21257));
  jand g21130(.dina(n21257), .dinb(n21248), .dout(n21258));
  jand g21131(.dina(n21258), .dinb(n21241), .dout(n21259));
  jand g21132(.dina(n1971), .dinb(n954), .dout(n21260));
  jand g21133(.dina(n21260), .dinb(n11224), .dout(n21261));
  jand g21134(.dina(n510), .dinb(n1351), .dout(n21262));
  jand g21135(.dina(n826), .dinb(n557), .dout(n21263));
  jand g21136(.dina(n21263), .dinb(n21262), .dout(n21264));
  jand g21137(.dina(n1903), .dinb(n452), .dout(n21265));
  jand g21138(.dina(n428), .dinb(n676), .dout(n21266));
  jand g21139(.dina(n21266), .dinb(n21265), .dout(n21267));
  jand g21140(.dina(n21267), .dinb(n21264), .dout(n21268));
  jand g21141(.dina(n21268), .dinb(n549), .dout(n21269));
  jand g21142(.dina(n2386), .dinb(n989), .dout(n21270));
  jand g21143(.dina(n645), .dinb(n1701), .dout(n21271));
  jand g21144(.dina(n21271), .dinb(n1471), .dout(n21272));
  jand g21145(.dina(n21272), .dinb(n664), .dout(n21273));
  jand g21146(.dina(n21273), .dinb(n21270), .dout(n21274));
  jand g21147(.dina(n21274), .dinb(n21269), .dout(n21275));
  jand g21148(.dina(n21275), .dinb(n21123), .dout(n21276));
  jand g21149(.dina(n21276), .dinb(n21261), .dout(n21277));
  jand g21150(.dina(n21277), .dinb(n21259), .dout(n21278));
  jand g21151(.dina(n21278), .dinb(n1202), .dout(n21279));
  jnot g21152(.din(n21279), .dout(n21280));
  jor  g21153(.dina(n21140), .dinb(n21027), .dout(n21281));
  jand g21154(.dina(n21144), .dinb(n21141), .dout(n21282));
  jnot g21155(.din(n21282), .dout(n21283));
  jand g21156(.dina(n21283), .dinb(n21281), .dout(n21284));
  jxor g21157(.dina(n21284), .dinb(n21280), .dout(n21285));
  jand g21158(.dina(n13616), .dinb(n5076), .dout(n21286));
  jand g21159(.dina(n13614), .dinb(n5084), .dout(n21287));
  jand g21160(.dina(n13478), .dinb(n6050), .dout(n21288));
  jand g21161(.dina(n13469), .dinb(n5082), .dout(n21289));
  jor  g21162(.dina(n21289), .dinb(n21288), .dout(n21290));
  jor  g21163(.dina(n21290), .dinb(n21287), .dout(n21291));
  jor  g21164(.dina(n21291), .dinb(n21286), .dout(n21292));
  jxor g21165(.dina(n21292), .dinb(n21285), .dout(n21293));
  jxor g21166(.dina(n21293), .dinb(n21236), .dout(n21294));
  jnot g21167(.din(n21294), .dout(n21295));
  jand g21168(.dina(n14562), .dinb(n2936), .dout(n21296));
  jand g21169(.dina(n14448), .dinb(n2940), .dout(n21297));
  jand g21170(.dina(n14447), .dinb(n2943), .dout(n21298));
  jor  g21171(.dina(n21298), .dinb(n21297), .dout(n21299));
  jand g21172(.dina(n14249), .dinb(n3684), .dout(n21300));
  jor  g21173(.dina(n21300), .dinb(n21299), .dout(n21301));
  jor  g21174(.dina(n21301), .dinb(n21296), .dout(n21302));
  jxor g21175(.dina(n21302), .dinb(n93), .dout(n21303));
  jxor g21176(.dina(n21303), .dinb(n21295), .dout(n21304));
  jxor g21177(.dina(n21304), .dinb(n21233), .dout(n21305));
  jnot g21178(.din(n21305), .dout(n21306));
  jand g21179(.dina(n15569), .dinb(n71), .dout(n21307));
  jand g21180(.dina(n15567), .dinb(n796), .dout(n21308));
  jand g21181(.dina(n15315), .dinb(n731), .dout(n21309));
  jand g21182(.dina(n14549), .dinb(n1806), .dout(n21310));
  jor  g21183(.dina(n21310), .dinb(n21309), .dout(n21311));
  jor  g21184(.dina(n21311), .dinb(n21308), .dout(n21312));
  jor  g21185(.dina(n21312), .dinb(n21307), .dout(n21313));
  jxor g21186(.dina(n21313), .dinb(n77), .dout(n21314));
  jxor g21187(.dina(n21314), .dinb(n21306), .dout(n21315));
  jxor g21188(.dina(n21315), .dinb(n21228), .dout(n21316));
  jnot g21189(.din(n21316), .dout(n21317));
  jand g21190(.dina(n16345), .dinb(n806), .dout(n21318));
  jand g21191(.dina(n16082), .dinb(n1612), .dout(n21319));
  jand g21192(.dina(n16343), .dinb(n1620), .dout(n21320));
  jor  g21193(.dina(n21320), .dinb(n21319), .dout(n21321));
  jand g21194(.dina(n15829), .dinb(n1644), .dout(n21322));
  jor  g21195(.dina(n21322), .dinb(n21321), .dout(n21323));
  jor  g21196(.dina(n21323), .dinb(n21318), .dout(n21324));
  jxor g21197(.dina(n21324), .dinb(n65), .dout(n21325));
  jxor g21198(.dina(n21325), .dinb(n21317), .dout(n21326));
  jxor g21199(.dina(n21326), .dinb(n21223), .dout(n21327));
  jnot g21200(.din(n21327), .dout(n21328));
  jand g21201(.dina(n17312), .dinb(n1819), .dout(n21329));
  jand g21202(.dina(n16928), .dinb(n2180), .dout(n21330));
  jand g21203(.dina(n16924), .dinb(n2243), .dout(n21331));
  jand g21204(.dina(n16592), .dinb(n2185), .dout(n21332));
  jor  g21205(.dina(n21332), .dinb(n21331), .dout(n21333));
  jor  g21206(.dina(n21333), .dinb(n21330), .dout(n21334));
  jor  g21207(.dina(n21334), .dinb(n21329), .dout(n21335));
  jxor g21208(.dina(n21335), .dinb(n2196), .dout(n21336));
  jxor g21209(.dina(n21336), .dinb(n21328), .dout(n21337));
  jxor g21210(.dina(n21337), .dinb(n21218), .dout(n21338));
  jnot g21211(.din(n21338), .dout(n21339));
  jxor g21212(.dina(n21339), .dinb(n21213), .dout(n21340));
  jxor g21213(.dina(n21340), .dinb(n21197), .dout(n21341));
  jxor g21214(.dina(n21341), .dinb(n21209), .dout(n21342));
  jand g21215(.dina(n21342), .dinb(n4691), .dout(n21343));
  jand g21216(.dina(n21340), .dinb(n4941), .dout(n21344));
  jand g21217(.dina(n21197), .dinb(n4696), .dout(n21345));
  jand g21218(.dina(n21198), .dinb(n4701), .dout(n21346));
  jor  g21219(.dina(n21346), .dinb(n21345), .dout(n21347));
  jor  g21220(.dina(n21347), .dinb(n21344), .dout(n21348));
  jor  g21221(.dina(n21348), .dinb(n21343), .dout(n21349));
  jxor g21222(.dina(n21349), .dinb(n4713), .dout(n21350));
  jor  g21223(.dina(n21350), .dinb(n20959), .dout(n21351));
  jnot g21224(.din(n21351), .dout(n21352));
  jxor g21225(.dina(n20672), .dinb(n20671), .dout(n21353));
  jnot g21226(.din(n21353), .dout(n21354));
  jxor g21227(.dina(n21207), .dinb(n21206), .dout(n21355));
  jand g21228(.dina(n21355), .dinb(n4691), .dout(n21356));
  jand g21229(.dina(n21198), .dinb(n4696), .dout(n21357));
  jand g21230(.dina(n21197), .dinb(n4941), .dout(n21358));
  jor  g21231(.dina(n21358), .dinb(n21357), .dout(n21359));
  jand g21232(.dina(n20947), .dinb(n4701), .dout(n21360));
  jor  g21233(.dina(n21360), .dinb(n21359), .dout(n21361));
  jor  g21234(.dina(n21361), .dinb(n21356), .dout(n21362));
  jxor g21235(.dina(n21362), .dinb(n4713), .dout(n21363));
  jor  g21236(.dina(n21363), .dinb(n21354), .dout(n21364));
  jxor g21237(.dina(n20669), .dinb(n20668), .dout(n21365));
  jnot g21238(.din(n21365), .dout(n21366));
  jxor g21239(.dina(n21204), .dinb(n21203), .dout(n21367));
  jand g21240(.dina(n21367), .dinb(n4691), .dout(n21368));
  jand g21241(.dina(n20947), .dinb(n4696), .dout(n21369));
  jand g21242(.dina(n21198), .dinb(n4941), .dout(n21370));
  jor  g21243(.dina(n21370), .dinb(n21369), .dout(n21371));
  jand g21244(.dina(n20344), .dinb(n4701), .dout(n21372));
  jor  g21245(.dina(n21372), .dinb(n21371), .dout(n21373));
  jor  g21246(.dina(n21373), .dinb(n21368), .dout(n21374));
  jxor g21247(.dina(n21374), .dinb(n4713), .dout(n21375));
  jor  g21248(.dina(n21375), .dinb(n21366), .dout(n21376));
  jxor g21249(.dina(n20666), .dinb(n20665), .dout(n21377));
  jnot g21250(.din(n21377), .dout(n21378));
  jand g21251(.dina(n20949), .dinb(n4691), .dout(n21379));
  jand g21252(.dina(n20344), .dinb(n4696), .dout(n21380));
  jand g21253(.dina(n20947), .dinb(n4941), .dout(n21381));
  jor  g21254(.dina(n21381), .dinb(n21380), .dout(n21382));
  jand g21255(.dina(n20204), .dinb(n4701), .dout(n21383));
  jor  g21256(.dina(n21383), .dinb(n21382), .dout(n21384));
  jor  g21257(.dina(n21384), .dinb(n21379), .dout(n21385));
  jxor g21258(.dina(n21385), .dinb(n4713), .dout(n21386));
  jor  g21259(.dina(n21386), .dinb(n21378), .dout(n21387));
  jxor g21260(.dina(n20663), .dinb(n20661), .dout(n21388));
  jand g21261(.dina(n20346), .dinb(n4691), .dout(n21389));
  jand g21262(.dina(n20344), .dinb(n4941), .dout(n21390));
  jand g21263(.dina(n20204), .dinb(n4696), .dout(n21391));
  jand g21264(.dina(n20205), .dinb(n4701), .dout(n21392));
  jor  g21265(.dina(n21392), .dinb(n21391), .dout(n21393));
  jor  g21266(.dina(n21393), .dinb(n21390), .dout(n21394));
  jor  g21267(.dina(n21394), .dinb(n21389), .dout(n21395));
  jxor g21268(.dina(n21395), .dinb(n4713), .dout(n21396));
  jor  g21269(.dina(n21396), .dinb(n21388), .dout(n21397));
  jxor g21270(.dina(n20659), .dinb(n20657), .dout(n21398));
  jnot g21271(.din(n21398), .dout(n21399));
  jand g21272(.dina(n20358), .dinb(n4691), .dout(n21400));
  jand g21273(.dina(n20205), .dinb(n4696), .dout(n21401));
  jand g21274(.dina(n20204), .dinb(n4941), .dout(n21402));
  jor  g21275(.dina(n21402), .dinb(n21401), .dout(n21403));
  jand g21276(.dina(n19922), .dinb(n4701), .dout(n21404));
  jor  g21277(.dina(n21404), .dinb(n21403), .dout(n21405));
  jor  g21278(.dina(n21405), .dinb(n21400), .dout(n21406));
  jxor g21279(.dina(n21406), .dinb(n4713), .dout(n21407));
  jor  g21280(.dina(n21407), .dinb(n21399), .dout(n21408));
  jxor g21281(.dina(n20655), .dinb(n20653), .dout(n21409));
  jnot g21282(.din(n21409), .dout(n21410));
  jand g21283(.dina(n20371), .dinb(n4691), .dout(n21411));
  jand g21284(.dina(n19922), .dinb(n4696), .dout(n21412));
  jand g21285(.dina(n20205), .dinb(n4941), .dout(n21413));
  jor  g21286(.dina(n21413), .dinb(n21412), .dout(n21414));
  jand g21287(.dina(n19373), .dinb(n4701), .dout(n21415));
  jor  g21288(.dina(n21415), .dinb(n21414), .dout(n21416));
  jor  g21289(.dina(n21416), .dinb(n21411), .dout(n21417));
  jxor g21290(.dina(n21417), .dinb(n4713), .dout(n21418));
  jor  g21291(.dina(n21418), .dinb(n21410), .dout(n21419));
  jxor g21292(.dina(n20651), .dinb(n20649), .dout(n21420));
  jnot g21293(.din(n21420), .dout(n21421));
  jand g21294(.dina(n19924), .dinb(n4691), .dout(n21422));
  jand g21295(.dina(n19922), .dinb(n4941), .dout(n21423));
  jand g21296(.dina(n19373), .dinb(n4696), .dout(n21424));
  jand g21297(.dina(n19219), .dinb(n4701), .dout(n21425));
  jor  g21298(.dina(n21425), .dinb(n21424), .dout(n21426));
  jor  g21299(.dina(n21426), .dinb(n21423), .dout(n21427));
  jor  g21300(.dina(n21427), .dinb(n21422), .dout(n21428));
  jxor g21301(.dina(n21428), .dinb(n4713), .dout(n21429));
  jor  g21302(.dina(n21429), .dinb(n21421), .dout(n21430));
  jxor g21303(.dina(n20646), .dinb(n20645), .dout(n21431));
  jnot g21304(.din(n21431), .dout(n21432));
  jand g21305(.dina(n19375), .dinb(n4691), .dout(n21433));
  jand g21306(.dina(n19219), .dinb(n4696), .dout(n21434));
  jand g21307(.dina(n19373), .dinb(n4941), .dout(n21435));
  jor  g21308(.dina(n21435), .dinb(n21434), .dout(n21436));
  jand g21309(.dina(n19220), .dinb(n4701), .dout(n21437));
  jor  g21310(.dina(n21437), .dinb(n21436), .dout(n21438));
  jor  g21311(.dina(n21438), .dinb(n21433), .dout(n21439));
  jxor g21312(.dina(n21439), .dinb(n4713), .dout(n21440));
  jor  g21313(.dina(n21440), .dinb(n21432), .dout(n21441));
  jxor g21314(.dina(n20641), .dinb(n20640), .dout(n21442));
  jnot g21315(.din(n21442), .dout(n21443));
  jand g21316(.dina(n19387), .dinb(n4691), .dout(n21444));
  jand g21317(.dina(n19219), .dinb(n4941), .dout(n21445));
  jand g21318(.dina(n19220), .dinb(n4696), .dout(n21446));
  jand g21319(.dina(n18914), .dinb(n4701), .dout(n21447));
  jor  g21320(.dina(n21447), .dinb(n21446), .dout(n21448));
  jor  g21321(.dina(n21448), .dinb(n21445), .dout(n21449));
  jor  g21322(.dina(n21449), .dinb(n21444), .dout(n21450));
  jxor g21323(.dina(n21450), .dinb(n4713), .dout(n21451));
  jor  g21324(.dina(n21451), .dinb(n21443), .dout(n21452));
  jxor g21325(.dina(n20636), .dinb(n20635), .dout(n21453));
  jnot g21326(.din(n21453), .dout(n21454));
  jand g21327(.dina(n19399), .dinb(n4691), .dout(n21455));
  jand g21328(.dina(n19220), .dinb(n4941), .dout(n21456));
  jand g21329(.dina(n18914), .dinb(n4696), .dout(n21457));
  jand g21330(.dina(n18488), .dinb(n4701), .dout(n21458));
  jor  g21331(.dina(n21458), .dinb(n21457), .dout(n21459));
  jor  g21332(.dina(n21459), .dinb(n21456), .dout(n21460));
  jor  g21333(.dina(n21460), .dinb(n21455), .dout(n21461));
  jxor g21334(.dina(n21461), .dinb(n4713), .dout(n21462));
  jor  g21335(.dina(n21462), .dinb(n21454), .dout(n21463));
  jxor g21336(.dina(n20631), .dinb(n20630), .dout(n21464));
  jnot g21337(.din(n21464), .dout(n21465));
  jand g21338(.dina(n18916), .dinb(n4691), .dout(n21466));
  jand g21339(.dina(n18488), .dinb(n4696), .dout(n21467));
  jand g21340(.dina(n18914), .dinb(n4941), .dout(n21468));
  jor  g21341(.dina(n21468), .dinb(n21467), .dout(n21469));
  jand g21342(.dina(n18292), .dinb(n4701), .dout(n21470));
  jor  g21343(.dina(n21470), .dinb(n21469), .dout(n21471));
  jor  g21344(.dina(n21471), .dinb(n21466), .dout(n21472));
  jxor g21345(.dina(n21472), .dinb(n4713), .dout(n21473));
  jor  g21346(.dina(n21473), .dinb(n21465), .dout(n21474));
  jxor g21347(.dina(n20626), .dinb(n20625), .dout(n21475));
  jnot g21348(.din(n21475), .dout(n21476));
  jand g21349(.dina(n18490), .dinb(n4691), .dout(n21477));
  jand g21350(.dina(n18488), .dinb(n4941), .dout(n21478));
  jand g21351(.dina(n18292), .dinb(n4696), .dout(n21479));
  jand g21352(.dina(n18293), .dinb(n4701), .dout(n21480));
  jor  g21353(.dina(n21480), .dinb(n21479), .dout(n21481));
  jor  g21354(.dina(n21481), .dinb(n21478), .dout(n21482));
  jor  g21355(.dina(n21482), .dinb(n21477), .dout(n21483));
  jxor g21356(.dina(n21483), .dinb(n4713), .dout(n21484));
  jor  g21357(.dina(n21484), .dinb(n21476), .dout(n21485));
  jxor g21358(.dina(n20621), .dinb(n20620), .dout(n21486));
  jnot g21359(.din(n21486), .dout(n21487));
  jand g21360(.dina(n18502), .dinb(n4691), .dout(n21488));
  jand g21361(.dina(n18293), .dinb(n4696), .dout(n21489));
  jand g21362(.dina(n18292), .dinb(n4941), .dout(n21490));
  jor  g21363(.dina(n21490), .dinb(n21489), .dout(n21491));
  jand g21364(.dina(n17942), .dinb(n4701), .dout(n21492));
  jor  g21365(.dina(n21492), .dinb(n21491), .dout(n21493));
  jor  g21366(.dina(n21493), .dinb(n21488), .dout(n21494));
  jxor g21367(.dina(n21494), .dinb(n4713), .dout(n21495));
  jor  g21368(.dina(n21495), .dinb(n21487), .dout(n21496));
  jxor g21369(.dina(n20616), .dinb(n20615), .dout(n21497));
  jnot g21370(.din(n21497), .dout(n21498));
  jand g21371(.dina(n18514), .dinb(n4691), .dout(n21499));
  jand g21372(.dina(n18293), .dinb(n4941), .dout(n21500));
  jand g21373(.dina(n17942), .dinb(n4696), .dout(n21501));
  jand g21374(.dina(n17535), .dinb(n4701), .dout(n21502));
  jor  g21375(.dina(n21502), .dinb(n21501), .dout(n21503));
  jor  g21376(.dina(n21503), .dinb(n21500), .dout(n21504));
  jor  g21377(.dina(n21504), .dinb(n21499), .dout(n21505));
  jxor g21378(.dina(n21505), .dinb(n4713), .dout(n21506));
  jor  g21379(.dina(n21506), .dinb(n21498), .dout(n21507));
  jxor g21380(.dina(n20611), .dinb(n20610), .dout(n21508));
  jnot g21381(.din(n21508), .dout(n21509));
  jand g21382(.dina(n17944), .dinb(n4691), .dout(n21510));
  jand g21383(.dina(n17942), .dinb(n4941), .dout(n21511));
  jand g21384(.dina(n17535), .dinb(n4696), .dout(n21512));
  jand g21385(.dina(n17329), .dinb(n4701), .dout(n21513));
  jor  g21386(.dina(n21513), .dinb(n21512), .dout(n21514));
  jor  g21387(.dina(n21514), .dinb(n21511), .dout(n21515));
  jor  g21388(.dina(n21515), .dinb(n21510), .dout(n21516));
  jxor g21389(.dina(n21516), .dinb(n4713), .dout(n21517));
  jor  g21390(.dina(n21517), .dinb(n21509), .dout(n21518));
  jxor g21391(.dina(n20606), .dinb(n20605), .dout(n21519));
  jnot g21392(.din(n21519), .dout(n21520));
  jand g21393(.dina(n17537), .dinb(n4691), .dout(n21521));
  jand g21394(.dina(n17535), .dinb(n4941), .dout(n21522));
  jand g21395(.dina(n17329), .dinb(n4696), .dout(n21523));
  jand g21396(.dina(n17330), .dinb(n4701), .dout(n21524));
  jor  g21397(.dina(n21524), .dinb(n21523), .dout(n21525));
  jor  g21398(.dina(n21525), .dinb(n21522), .dout(n21526));
  jor  g21399(.dina(n21526), .dinb(n21521), .dout(n21527));
  jxor g21400(.dina(n21527), .dinb(n4713), .dout(n21528));
  jor  g21401(.dina(n21528), .dinb(n21520), .dout(n21529));
  jxor g21402(.dina(n20601), .dinb(n20600), .dout(n21530));
  jnot g21403(.din(n21530), .dout(n21531));
  jand g21404(.dina(n17549), .dinb(n4691), .dout(n21532));
  jand g21405(.dina(n17329), .dinb(n4941), .dout(n21533));
  jand g21406(.dina(n17330), .dinb(n4696), .dout(n21534));
  jand g21407(.dina(n16940), .dinb(n4701), .dout(n21535));
  jor  g21408(.dina(n21535), .dinb(n21534), .dout(n21536));
  jor  g21409(.dina(n21536), .dinb(n21533), .dout(n21537));
  jor  g21410(.dina(n21537), .dinb(n21532), .dout(n21538));
  jxor g21411(.dina(n21538), .dinb(n4713), .dout(n21539));
  jor  g21412(.dina(n21539), .dinb(n21531), .dout(n21540));
  jxor g21413(.dina(n20598), .dinb(n20597), .dout(n21541));
  jnot g21414(.din(n21541), .dout(n21542));
  jand g21415(.dina(n17561), .dinb(n4691), .dout(n21543));
  jand g21416(.dina(n16940), .dinb(n4696), .dout(n21544));
  jand g21417(.dina(n17330), .dinb(n4941), .dout(n21545));
  jor  g21418(.dina(n21545), .dinb(n21544), .dout(n21546));
  jand g21419(.dina(n16604), .dinb(n4701), .dout(n21547));
  jor  g21420(.dina(n21547), .dinb(n21546), .dout(n21548));
  jor  g21421(.dina(n21548), .dinb(n21543), .dout(n21549));
  jxor g21422(.dina(n21549), .dinb(n4713), .dout(n21550));
  jor  g21423(.dina(n21550), .dinb(n21542), .dout(n21551));
  jxor g21424(.dina(n20593), .dinb(n20592), .dout(n21552));
  jnot g21425(.din(n21552), .dout(n21553));
  jand g21426(.dina(n16942), .dinb(n4691), .dout(n21554));
  jand g21427(.dina(n16940), .dinb(n4941), .dout(n21555));
  jand g21428(.dina(n16355), .dinb(n4701), .dout(n21556));
  jand g21429(.dina(n16604), .dinb(n4696), .dout(n21557));
  jor  g21430(.dina(n21557), .dinb(n21556), .dout(n21558));
  jor  g21431(.dina(n21558), .dinb(n21555), .dout(n21559));
  jor  g21432(.dina(n21559), .dinb(n21554), .dout(n21560));
  jxor g21433(.dina(n21560), .dinb(n4713), .dout(n21561));
  jor  g21434(.dina(n21561), .dinb(n21553), .dout(n21562));
  jxor g21435(.dina(n20589), .dinb(n20581), .dout(n21563));
  jnot g21436(.din(n21563), .dout(n21564));
  jand g21437(.dina(n16606), .dinb(n4691), .dout(n21565));
  jand g21438(.dina(n16355), .dinb(n4696), .dout(n21566));
  jand g21439(.dina(n16604), .dinb(n4941), .dout(n21567));
  jor  g21440(.dina(n21567), .dinb(n21566), .dout(n21568));
  jand g21441(.dina(n16360), .dinb(n4701), .dout(n21569));
  jor  g21442(.dina(n21569), .dinb(n21568), .dout(n21570));
  jor  g21443(.dina(n21570), .dinb(n21565), .dout(n21571));
  jxor g21444(.dina(n21571), .dinb(n4713), .dout(n21572));
  jor  g21445(.dina(n21572), .dinb(n21564), .dout(n21573));
  jand g21446(.dina(n16616), .dinb(n4691), .dout(n21574));
  jand g21447(.dina(n16360), .dinb(n4696), .dout(n21575));
  jand g21448(.dina(n16355), .dinb(n4941), .dout(n21576));
  jor  g21449(.dina(n21576), .dinb(n21575), .dout(n21577));
  jand g21450(.dina(n15841), .dinb(n4701), .dout(n21578));
  jor  g21451(.dina(n21578), .dinb(n21577), .dout(n21579));
  jor  g21452(.dina(n21579), .dinb(n21574), .dout(n21580));
  jxor g21453(.dina(n21580), .dinb(n4713), .dout(n21581));
  jnot g21454(.din(n21581), .dout(n21582));
  jor  g21455(.dina(n20568), .dinb(n4050), .dout(n21583));
  jxor g21456(.dina(n21583), .dinb(n20576), .dout(n21584));
  jand g21457(.dina(n21584), .dinb(n21582), .dout(n21585));
  jand g21458(.dina(n20565), .dinb(\a[11] ), .dout(n21586));
  jxor g21459(.dina(n21586), .dinb(n20563), .dout(n21587));
  jnot g21460(.din(n21587), .dout(n21588));
  jand g21461(.dina(n16632), .dinb(n4691), .dout(n21589));
  jand g21462(.dina(n15841), .dinb(n4696), .dout(n21590));
  jand g21463(.dina(n16360), .dinb(n4941), .dout(n21591));
  jor  g21464(.dina(n21591), .dinb(n21590), .dout(n21592));
  jand g21465(.dina(n15579), .dinb(n4701), .dout(n21593));
  jor  g21466(.dina(n21593), .dinb(n21592), .dout(n21594));
  jor  g21467(.dina(n21594), .dinb(n21589), .dout(n21595));
  jxor g21468(.dina(n21595), .dinb(n4713), .dout(n21596));
  jor  g21469(.dina(n21596), .dinb(n21588), .dout(n21597));
  jand g21470(.dina(n15329), .dinb(n4691), .dout(n21598));
  jand g21471(.dina(n15327), .dinb(n4941), .dout(n21599));
  jand g21472(.dina(n15020), .dinb(n4696), .dout(n21600));
  jor  g21473(.dina(n21600), .dinb(n21599), .dout(n21601));
  jor  g21474(.dina(n21601), .dinb(n21598), .dout(n21602));
  jnot g21475(.din(n21602), .dout(n21603));
  jand g21476(.dina(n15020), .dinb(n4689), .dout(n21604));
  jnot g21477(.din(n21604), .dout(n21605));
  jand g21478(.dina(n21605), .dinb(\a[8] ), .dout(n21606));
  jand g21479(.dina(n21606), .dinb(n21603), .dout(n21607));
  jand g21480(.dina(n15580), .dinb(n4691), .dout(n21608));
  jand g21481(.dina(n15327), .dinb(n4696), .dout(n21609));
  jor  g21482(.dina(n21609), .dinb(n21608), .dout(n21610));
  jand g21483(.dina(n15579), .dinb(n4941), .dout(n21611));
  jand g21484(.dina(n15020), .dinb(n4701), .dout(n21612));
  jor  g21485(.dina(n21612), .dinb(n21611), .dout(n21613));
  jor  g21486(.dina(n21613), .dinb(n21610), .dout(n21614));
  jnot g21487(.din(n21614), .dout(n21615));
  jand g21488(.dina(n21615), .dinb(n21607), .dout(n21616));
  jand g21489(.dina(n21616), .dinb(n20565), .dout(n21617));
  jnot g21490(.din(n21617), .dout(n21618));
  jxor g21491(.dina(n21616), .dinb(n20565), .dout(n21619));
  jnot g21492(.din(n21619), .dout(n21620));
  jand g21493(.dina(n15848), .dinb(n4691), .dout(n21621));
  jand g21494(.dina(n15841), .dinb(n4941), .dout(n21622));
  jand g21495(.dina(n15579), .dinb(n4696), .dout(n21623));
  jand g21496(.dina(n15327), .dinb(n4701), .dout(n21624));
  jor  g21497(.dina(n21624), .dinb(n21623), .dout(n21625));
  jor  g21498(.dina(n21625), .dinb(n21622), .dout(n21626));
  jor  g21499(.dina(n21626), .dinb(n21621), .dout(n21627));
  jxor g21500(.dina(n21627), .dinb(n4713), .dout(n21628));
  jor  g21501(.dina(n21628), .dinb(n21620), .dout(n21629));
  jand g21502(.dina(n21629), .dinb(n21618), .dout(n21630));
  jnot g21503(.din(n21630), .dout(n21631));
  jxor g21504(.dina(n21596), .dinb(n21588), .dout(n21632));
  jand g21505(.dina(n21632), .dinb(n21631), .dout(n21633));
  jnot g21506(.din(n21633), .dout(n21634));
  jand g21507(.dina(n21634), .dinb(n21597), .dout(n21635));
  jnot g21508(.din(n21635), .dout(n21636));
  jxor g21509(.dina(n21584), .dinb(n21582), .dout(n21637));
  jand g21510(.dina(n21637), .dinb(n21636), .dout(n21638));
  jor  g21511(.dina(n21638), .dinb(n21585), .dout(n21639));
  jxor g21512(.dina(n21572), .dinb(n21564), .dout(n21640));
  jand g21513(.dina(n21640), .dinb(n21639), .dout(n21641));
  jnot g21514(.din(n21641), .dout(n21642));
  jand g21515(.dina(n21642), .dinb(n21573), .dout(n21643));
  jnot g21516(.din(n21643), .dout(n21644));
  jxor g21517(.dina(n21561), .dinb(n21553), .dout(n21645));
  jand g21518(.dina(n21645), .dinb(n21644), .dout(n21646));
  jnot g21519(.din(n21646), .dout(n21647));
  jand g21520(.dina(n21647), .dinb(n21562), .dout(n21648));
  jnot g21521(.din(n21648), .dout(n21649));
  jxor g21522(.dina(n21550), .dinb(n21542), .dout(n21650));
  jand g21523(.dina(n21650), .dinb(n21649), .dout(n21651));
  jnot g21524(.din(n21651), .dout(n21652));
  jand g21525(.dina(n21652), .dinb(n21551), .dout(n21653));
  jnot g21526(.din(n21653), .dout(n21654));
  jxor g21527(.dina(n21539), .dinb(n21531), .dout(n21655));
  jand g21528(.dina(n21655), .dinb(n21654), .dout(n21656));
  jnot g21529(.din(n21656), .dout(n21657));
  jand g21530(.dina(n21657), .dinb(n21540), .dout(n21658));
  jnot g21531(.din(n21658), .dout(n21659));
  jxor g21532(.dina(n21528), .dinb(n21520), .dout(n21660));
  jand g21533(.dina(n21660), .dinb(n21659), .dout(n21661));
  jnot g21534(.din(n21661), .dout(n21662));
  jand g21535(.dina(n21662), .dinb(n21529), .dout(n21663));
  jnot g21536(.din(n21663), .dout(n21664));
  jxor g21537(.dina(n21517), .dinb(n21509), .dout(n21665));
  jand g21538(.dina(n21665), .dinb(n21664), .dout(n21666));
  jnot g21539(.din(n21666), .dout(n21667));
  jand g21540(.dina(n21667), .dinb(n21518), .dout(n21668));
  jnot g21541(.din(n21668), .dout(n21669));
  jxor g21542(.dina(n21506), .dinb(n21498), .dout(n21670));
  jand g21543(.dina(n21670), .dinb(n21669), .dout(n21671));
  jnot g21544(.din(n21671), .dout(n21672));
  jand g21545(.dina(n21672), .dinb(n21507), .dout(n21673));
  jnot g21546(.din(n21673), .dout(n21674));
  jxor g21547(.dina(n21495), .dinb(n21487), .dout(n21675));
  jand g21548(.dina(n21675), .dinb(n21674), .dout(n21676));
  jnot g21549(.din(n21676), .dout(n21677));
  jand g21550(.dina(n21677), .dinb(n21496), .dout(n21678));
  jxor g21551(.dina(n21484), .dinb(n21476), .dout(n21679));
  jnot g21552(.din(n21679), .dout(n21680));
  jor  g21553(.dina(n21680), .dinb(n21678), .dout(n21681));
  jand g21554(.dina(n21681), .dinb(n21485), .dout(n21682));
  jxor g21555(.dina(n21473), .dinb(n21465), .dout(n21683));
  jnot g21556(.din(n21683), .dout(n21684));
  jor  g21557(.dina(n21684), .dinb(n21682), .dout(n21685));
  jand g21558(.dina(n21685), .dinb(n21474), .dout(n21686));
  jxor g21559(.dina(n21462), .dinb(n21454), .dout(n21687));
  jnot g21560(.din(n21687), .dout(n21688));
  jor  g21561(.dina(n21688), .dinb(n21686), .dout(n21689));
  jand g21562(.dina(n21689), .dinb(n21463), .dout(n21690));
  jxor g21563(.dina(n21451), .dinb(n21443), .dout(n21691));
  jnot g21564(.din(n21691), .dout(n21692));
  jor  g21565(.dina(n21692), .dinb(n21690), .dout(n21693));
  jand g21566(.dina(n21693), .dinb(n21452), .dout(n21694));
  jxor g21567(.dina(n21440), .dinb(n21432), .dout(n21695));
  jnot g21568(.din(n21695), .dout(n21696));
  jor  g21569(.dina(n21696), .dinb(n21694), .dout(n21697));
  jand g21570(.dina(n21697), .dinb(n21441), .dout(n21698));
  jxor g21571(.dina(n21429), .dinb(n21420), .dout(n21699));
  jor  g21572(.dina(n21699), .dinb(n21698), .dout(n21700));
  jand g21573(.dina(n21700), .dinb(n21430), .dout(n21701));
  jxor g21574(.dina(n21418), .dinb(n21409), .dout(n21702));
  jor  g21575(.dina(n21702), .dinb(n21701), .dout(n21703));
  jand g21576(.dina(n21703), .dinb(n21419), .dout(n21704));
  jxor g21577(.dina(n21407), .dinb(n21398), .dout(n21705));
  jor  g21578(.dina(n21705), .dinb(n21704), .dout(n21706));
  jand g21579(.dina(n21706), .dinb(n21408), .dout(n21707));
  jxor g21580(.dina(n21396), .dinb(n21388), .dout(n21708));
  jnot g21581(.din(n21708), .dout(n21709));
  jor  g21582(.dina(n21709), .dinb(n21707), .dout(n21710));
  jand g21583(.dina(n21710), .dinb(n21397), .dout(n21711));
  jxor g21584(.dina(n21386), .dinb(n21377), .dout(n21712));
  jor  g21585(.dina(n21712), .dinb(n21711), .dout(n21713));
  jand g21586(.dina(n21713), .dinb(n21387), .dout(n21714));
  jxor g21587(.dina(n21375), .dinb(n21365), .dout(n21715));
  jor  g21588(.dina(n21715), .dinb(n21714), .dout(n21716));
  jand g21589(.dina(n21716), .dinb(n21376), .dout(n21717));
  jxor g21590(.dina(n21363), .dinb(n21353), .dout(n21718));
  jor  g21591(.dina(n21718), .dinb(n21717), .dout(n21719));
  jand g21592(.dina(n21719), .dinb(n21364), .dout(n21720));
  jnot g21593(.din(n21720), .dout(n21721));
  jxor g21594(.dina(n21350), .dinb(n20959), .dout(n21722));
  jand g21595(.dina(n21722), .dinb(n21721), .dout(n21723));
  jor  g21596(.dina(n21723), .dinb(n21352), .dout(n21724));
  jnot g21597(.din(n20798), .dout(n21725));
  jor  g21598(.dina(n20957), .dinb(n21725), .dout(n21726));
  jnot g21599(.din(n21726), .dout(n21727));
  jnot g21600(.din(n20958), .dout(n21728));
  jand g21601(.dina(n21728), .dinb(n20674), .dout(n21729));
  jor  g21602(.dina(n21729), .dinb(n21727), .dout(n21730));
  jor  g21603(.dina(n20796), .dinb(n20788), .dout(n21731));
  jnot g21604(.din(n21731), .dout(n21732));
  jand g21605(.dina(n20797), .dinb(n20678), .dout(n21733));
  jor  g21606(.dina(n21733), .dinb(n21732), .dout(n21734));
  jor  g21607(.dina(n20785), .dinb(n20777), .dout(n21735));
  jand g21608(.dina(n20786), .dinb(n20681), .dout(n21736));
  jnot g21609(.din(n21736), .dout(n21737));
  jand g21610(.dina(n21737), .dinb(n21735), .dout(n21738));
  jnot g21611(.din(n21738), .dout(n21739));
  jor  g21612(.dina(n20774), .dinb(n20766), .dout(n21740));
  jand g21613(.dina(n20775), .dinb(n20686), .dout(n21741));
  jnot g21614(.din(n21741), .dout(n21742));
  jand g21615(.dina(n21742), .dinb(n21740), .dout(n21743));
  jnot g21616(.din(n21743), .dout(n21744));
  jor  g21617(.dina(n20763), .dinb(n20755), .dout(n21745));
  jand g21618(.dina(n20764), .dinb(n20691), .dout(n21746));
  jnot g21619(.din(n21746), .dout(n21747));
  jand g21620(.dina(n21747), .dinb(n21745), .dout(n21748));
  jnot g21621(.din(n21748), .dout(n21749));
  jor  g21622(.dina(n20752), .dinb(n20744), .dout(n21750));
  jand g21623(.dina(n20753), .dinb(n20696), .dout(n21751));
  jnot g21624(.din(n21751), .dout(n21752));
  jand g21625(.dina(n21752), .dinb(n21750), .dout(n21753));
  jnot g21626(.din(n21753), .dout(n21754));
  jor  g21627(.dina(n20741), .dinb(n20733), .dout(n21755));
  jand g21628(.dina(n20742), .dinb(n20701), .dout(n21756));
  jnot g21629(.din(n21756), .dout(n21757));
  jand g21630(.dina(n21757), .dinb(n21755), .dout(n21758));
  jnot g21631(.din(n21758), .dout(n21759));
  jor  g21632(.dina(n20730), .dinb(n20710), .dout(n21760));
  jand g21633(.dina(n20731), .dinb(n20708), .dout(n21761));
  jnot g21634(.din(n21761), .dout(n21762));
  jand g21635(.dina(n21762), .dinb(n21760), .dout(n21763));
  jnot g21636(.din(n21763), .dout(n21764));
  jand g21637(.dina(n10202), .dinb(n3228), .dout(n21765));
  jand g21638(.dina(n1915), .dinb(n1225), .dout(n21766));
  jand g21639(.dina(n21766), .dinb(n1569), .dout(n21767));
  jand g21640(.dina(n1852), .dinb(n136), .dout(n21768));
  jand g21641(.dina(n895), .dinb(n662), .dout(n21769));
  jand g21642(.dina(n21769), .dinb(n21768), .dout(n21770));
  jand g21643(.dina(n21770), .dinb(n21767), .dout(n21771));
  jand g21644(.dina(n6335), .dinb(n2024), .dout(n21772));
  jand g21645(.dina(n21772), .dinb(n266), .dout(n21773));
  jand g21646(.dina(n21773), .dinb(n1088), .dout(n21774));
  jand g21647(.dina(n21774), .dinb(n21771), .dout(n21775));
  jand g21648(.dina(n21775), .dinb(n10194), .dout(n21776));
  jand g21649(.dina(n20117), .dinb(n1276), .dout(n21777));
  jand g21650(.dina(n21777), .dinb(n5396), .dout(n21778));
  jand g21651(.dina(n21778), .dinb(n21776), .dout(n21779));
  jand g21652(.dina(n21779), .dinb(n21765), .dout(n21780));
  jand g21653(.dina(n4553), .dinb(n2473), .dout(n21781));
  jand g21654(.dina(n21781), .dinb(n21780), .dout(n21782));
  jnot g21655(.din(n21782), .dout(n21783));
  jand g21656(.dina(n15848), .dinb(n5076), .dout(n21784));
  jand g21657(.dina(n15841), .dinb(n5084), .dout(n21785));
  jand g21658(.dina(n15327), .dinb(n6050), .dout(n21786));
  jand g21659(.dina(n15579), .dinb(n5082), .dout(n21787));
  jor  g21660(.dina(n21787), .dinb(n21786), .dout(n21788));
  jor  g21661(.dina(n21788), .dinb(n21785), .dout(n21789));
  jor  g21662(.dina(n21789), .dinb(n21784), .dout(n21790));
  jxor g21663(.dina(n21790), .dinb(n21783), .dout(n21791));
  jxor g21664(.dina(n21791), .dinb(n21764), .dout(n21792));
  jnot g21665(.din(n21792), .dout(n21793));
  jand g21666(.dina(n16606), .dinb(n2936), .dout(n21794));
  jand g21667(.dina(n16604), .dinb(n2943), .dout(n21795));
  jand g21668(.dina(n16355), .dinb(n2940), .dout(n21796));
  jand g21669(.dina(n16360), .dinb(n3684), .dout(n21797));
  jor  g21670(.dina(n21797), .dinb(n21796), .dout(n21798));
  jor  g21671(.dina(n21798), .dinb(n21795), .dout(n21799));
  jor  g21672(.dina(n21799), .dinb(n21794), .dout(n21800));
  jxor g21673(.dina(n21800), .dinb(n93), .dout(n21801));
  jxor g21674(.dina(n21801), .dinb(n21793), .dout(n21802));
  jxor g21675(.dina(n21802), .dinb(n21759), .dout(n21803));
  jnot g21676(.din(n21803), .dout(n21804));
  jand g21677(.dina(n17549), .dinb(n71), .dout(n21805));
  jand g21678(.dina(n17329), .dinb(n796), .dout(n21806));
  jand g21679(.dina(n17330), .dinb(n731), .dout(n21807));
  jand g21680(.dina(n16940), .dinb(n1806), .dout(n21808));
  jor  g21681(.dina(n21808), .dinb(n21807), .dout(n21809));
  jor  g21682(.dina(n21809), .dinb(n21806), .dout(n21810));
  jor  g21683(.dina(n21810), .dinb(n21805), .dout(n21811));
  jxor g21684(.dina(n21811), .dinb(n77), .dout(n21812));
  jxor g21685(.dina(n21812), .dinb(n21804), .dout(n21813));
  jxor g21686(.dina(n21813), .dinb(n21754), .dout(n21814));
  jnot g21687(.din(n21814), .dout(n21815));
  jand g21688(.dina(n18514), .dinb(n806), .dout(n21816));
  jand g21689(.dina(n18293), .dinb(n1620), .dout(n21817));
  jand g21690(.dina(n17942), .dinb(n1612), .dout(n21818));
  jand g21691(.dina(n17535), .dinb(n1644), .dout(n21819));
  jor  g21692(.dina(n21819), .dinb(n21818), .dout(n21820));
  jor  g21693(.dina(n21820), .dinb(n21817), .dout(n21821));
  jor  g21694(.dina(n21821), .dinb(n21816), .dout(n21822));
  jxor g21695(.dina(n21822), .dinb(n65), .dout(n21823));
  jxor g21696(.dina(n21823), .dinb(n21815), .dout(n21824));
  jxor g21697(.dina(n21824), .dinb(n21749), .dout(n21825));
  jnot g21698(.din(n21825), .dout(n21826));
  jand g21699(.dina(n18916), .dinb(n1819), .dout(n21827));
  jand g21700(.dina(n18914), .dinb(n2243), .dout(n21828));
  jand g21701(.dina(n18488), .dinb(n2180), .dout(n21829));
  jand g21702(.dina(n18292), .dinb(n2185), .dout(n21830));
  jor  g21703(.dina(n21830), .dinb(n21829), .dout(n21831));
  jor  g21704(.dina(n21831), .dinb(n21828), .dout(n21832));
  jor  g21705(.dina(n21832), .dinb(n21827), .dout(n21833));
  jxor g21706(.dina(n21833), .dinb(n2196), .dout(n21834));
  jxor g21707(.dina(n21834), .dinb(n21826), .dout(n21835));
  jxor g21708(.dina(n21835), .dinb(n21744), .dout(n21836));
  jnot g21709(.din(n21836), .dout(n21837));
  jand g21710(.dina(n19375), .dinb(n2743), .dout(n21838));
  jand g21711(.dina(n19373), .dinb(n2752), .dout(n21839));
  jand g21712(.dina(n19219), .dinb(n2748), .dout(n21840));
  jand g21713(.dina(n19220), .dinb(n2757), .dout(n21841));
  jor  g21714(.dina(n21841), .dinb(n21840), .dout(n21842));
  jor  g21715(.dina(n21842), .dinb(n21839), .dout(n21843));
  jor  g21716(.dina(n21843), .dinb(n21838), .dout(n21844));
  jxor g21717(.dina(n21844), .dinb(n2441), .dout(n21845));
  jxor g21718(.dina(n21845), .dinb(n21837), .dout(n21846));
  jxor g21719(.dina(n21846), .dinb(n21739), .dout(n21847));
  jnot g21720(.din(n21847), .dout(n21848));
  jand g21721(.dina(n20358), .dinb(n3423), .dout(n21849));
  jand g21722(.dina(n20204), .dinb(n3569), .dout(n21850));
  jand g21723(.dina(n20205), .dinb(n3428), .dout(n21851));
  jand g21724(.dina(n19922), .dinb(n3210), .dout(n21852));
  jor  g21725(.dina(n21852), .dinb(n21851), .dout(n21853));
  jor  g21726(.dina(n21853), .dinb(n21850), .dout(n21854));
  jor  g21727(.dina(n21854), .dinb(n21849), .dout(n21855));
  jxor g21728(.dina(n21855), .dinb(n3473), .dout(n21856));
  jxor g21729(.dina(n21856), .dinb(n21848), .dout(n21857));
  jxor g21730(.dina(n21857), .dinb(n21734), .dout(n21858));
  jand g21731(.dina(n21367), .dinb(n4022), .dout(n21859));
  jand g21732(.dina(n21198), .dinb(n4220), .dout(n21860));
  jand g21733(.dina(n20947), .dinb(n4027), .dout(n21861));
  jand g21734(.dina(n20344), .dinb(n3870), .dout(n21862));
  jor  g21735(.dina(n21862), .dinb(n21861), .dout(n21863));
  jor  g21736(.dina(n21863), .dinb(n21860), .dout(n21864));
  jor  g21737(.dina(n21864), .dinb(n21859), .dout(n21865));
  jxor g21738(.dina(n21865), .dinb(n4050), .dout(n21866));
  jxor g21739(.dina(n21866), .dinb(n21858), .dout(n21867));
  jnot g21740(.din(n21867), .dout(n21868));
  jxor g21741(.dina(n21868), .dinb(n21730), .dout(n21869));
  jand g21742(.dina(n21340), .dinb(n21197), .dout(n21870));
  jand g21743(.dina(n21341), .dinb(n21209), .dout(n21871));
  jor  g21744(.dina(n21871), .dinb(n21870), .dout(n21872));
  jand g21745(.dina(n21326), .dinb(n21223), .dout(n21873));
  jnot g21746(.din(n21873), .dout(n21874));
  jor  g21747(.dina(n21336), .dinb(n21328), .dout(n21875));
  jand g21748(.dina(n21875), .dinb(n21874), .dout(n21876));
  jnot g21749(.din(n21876), .dout(n21877));
  jand g21750(.dina(n21315), .dinb(n21228), .dout(n21878));
  jnot g21751(.din(n21878), .dout(n21879));
  jor  g21752(.dina(n21325), .dinb(n21317), .dout(n21880));
  jand g21753(.dina(n21880), .dinb(n21879), .dout(n21881));
  jor  g21754(.dina(n2184), .dinb(n1819), .dout(n21882));
  jxor g21755(.dina(n22046), .dinb(n21881), .dout(n21889));
  jand g21756(.dina(n21304), .dinb(n21233), .dout(n21890));
  jnot g21757(.din(n21890), .dout(n21891));
  jor  g21758(.dina(n21314), .dinb(n21306), .dout(n21892));
  jand g21759(.dina(n21892), .dinb(n21891), .dout(n21893));
  jnot g21760(.din(n21893), .dout(n21894));
  jor  g21761(.dina(n21284), .dinb(n21280), .dout(n21895));
  jand g21762(.dina(n21292), .dinb(n21285), .dout(n21896));
  jnot g21763(.din(n21896), .dout(n21897));
  jand g21764(.dina(n21897), .dinb(n21895), .dout(n21898));
  jnot g21765(.din(n21898), .dout(n21899));
  jand g21766(.dina(n14251), .dinb(n5076), .dout(n21900));
  jand g21767(.dina(n14249), .dinb(n5084), .dout(n21901));
  jand g21768(.dina(n13614), .dinb(n5082), .dout(n21902));
  jand g21769(.dina(n13469), .dinb(n6050), .dout(n21903));
  jor  g21770(.dina(n21903), .dinb(n21902), .dout(n21904));
  jor  g21771(.dina(n21904), .dinb(n21901), .dout(n21905));
  jor  g21772(.dina(n21905), .dinb(n21900), .dout(n21906));
  jand g21773(.dina(n499), .dinb(n699), .dout(n21907));
  jand g21774(.dina(n21907), .dinb(n11242), .dout(n21908));
  jand g21775(.dina(n1227), .dinb(n270), .dout(n21909));
  jand g21776(.dina(n21909), .dinb(n6441), .dout(n21910));
  jand g21777(.dina(n21910), .dinb(n21908), .dout(n21911));
  jand g21778(.dina(n3322), .dinb(n965), .dout(n21912));
  jand g21779(.dina(n21912), .dinb(n1465), .dout(n21913));
  jand g21780(.dina(n21913), .dinb(n3915), .dout(n21914));
  jand g21781(.dina(n21914), .dinb(n21911), .dout(n21915));
  jand g21782(.dina(n1162), .dinb(n1218), .dout(n21916));
  jand g21783(.dina(n21916), .dinb(n1822), .dout(n21917));
  jand g21784(.dina(n21917), .dinb(n4562), .dout(n21918));
  jand g21785(.dina(n9731), .dinb(n7104), .dout(n21919));
  jand g21786(.dina(n21919), .dinb(n21918), .dout(n21920));
  jand g21787(.dina(n7242), .dinb(n1283), .dout(n21921));
  jand g21788(.dina(n21921), .dinb(n21920), .dout(n21922));
  jand g21789(.dina(n21922), .dinb(n21915), .dout(n21923));
  jand g21790(.dina(n21923), .dinb(n2520), .dout(n21924));
  jand g21791(.dina(n17403), .dinb(n7792), .dout(n21925));
  jand g21792(.dina(n21925), .dinb(n21924), .dout(n21926));
  jxor g21793(.dina(n21926), .dinb(n21280), .dout(n21927));
  jxor g21794(.dina(n21927), .dinb(n21906), .dout(n21928));
  jxor g21795(.dina(n21928), .dinb(n21899), .dout(n21929));
  jnot g21796(.din(n21929), .dout(n21930));
  jand g21797(.dina(n21293), .dinb(n21236), .dout(n21931));
  jnot g21798(.din(n21931), .dout(n21932));
  jor  g21799(.dina(n21303), .dinb(n21295), .dout(n21933));
  jand g21800(.dina(n21933), .dinb(n21932), .dout(n21934));
  jxor g21801(.dina(n21934), .dinb(n21930), .dout(n21935));
  jnot g21802(.din(n21935), .dout(n21936));
  jand g21803(.dina(n14551), .dinb(n2936), .dout(n21937));
  jand g21804(.dina(n14447), .dinb(n2940), .dout(n21938));
  jand g21805(.dina(n14549), .dinb(n2943), .dout(n21939));
  jor  g21806(.dina(n21939), .dinb(n21938), .dout(n21940));
  jand g21807(.dina(n14448), .dinb(n3684), .dout(n21941));
  jor  g21808(.dina(n21941), .dinb(n21940), .dout(n21942));
  jor  g21809(.dina(n21942), .dinb(n21937), .dout(n21943));
  jxor g21810(.dina(n21943), .dinb(n93), .dout(n21944));
  jxor g21811(.dina(n21944), .dinb(n21936), .dout(n21945));
  jnot g21812(.din(n21945), .dout(n21946));
  jand g21813(.dina(n15831), .dinb(n71), .dout(n21947));
  jand g21814(.dina(n15829), .dinb(n796), .dout(n21948));
  jand g21815(.dina(n15567), .dinb(n731), .dout(n21949));
  jand g21816(.dina(n15315), .dinb(n1806), .dout(n21950));
  jor  g21817(.dina(n21950), .dinb(n21949), .dout(n21951));
  jor  g21818(.dina(n21951), .dinb(n21948), .dout(n21952));
  jor  g21819(.dina(n21952), .dinb(n21947), .dout(n21953));
  jxor g21820(.dina(n21953), .dinb(n77), .dout(n21954));
  jxor g21821(.dina(n21954), .dinb(n21946), .dout(n21955));
  jxor g21822(.dina(n21955), .dinb(n21894), .dout(n21956));
  jnot g21823(.din(n21956), .dout(n21957));
  jand g21824(.dina(n16594), .dinb(n806), .dout(n21958));
  jand g21825(.dina(n16592), .dinb(n1620), .dout(n21959));
  jand g21826(.dina(n16343), .dinb(n1612), .dout(n21960));
  jand g21827(.dina(n16082), .dinb(n1644), .dout(n21961));
  jor  g21828(.dina(n21961), .dinb(n21960), .dout(n21962));
  jor  g21829(.dina(n21962), .dinb(n21959), .dout(n21963));
  jor  g21830(.dina(n21963), .dinb(n21958), .dout(n21964));
  jxor g21831(.dina(n21964), .dinb(n65), .dout(n21965));
  jxor g21832(.dina(n21965), .dinb(n21957), .dout(n21966));
  jxor g21833(.dina(n21966), .dinb(n21889), .dout(n21967));
  jxor g21834(.dina(n21967), .dinb(n21877), .dout(n21968));
  jnot g21835(.din(n21968), .dout(n21969));
  jand g21836(.dina(n21337), .dinb(n21218), .dout(n21970));
  jnot g21837(.din(n21970), .dout(n21971));
  jor  g21838(.dina(n21339), .dinb(n21213), .dout(n21972));
  jand g21839(.dina(n21972), .dinb(n21971), .dout(n21973));
  jxor g21840(.dina(n21973), .dinb(n21969), .dout(n21974));
  jxor g21841(.dina(n21974), .dinb(n21340), .dout(n21975));
  jxor g21842(.dina(n21975), .dinb(n21872), .dout(n21976));
  jand g21843(.dina(n21976), .dinb(n4691), .dout(n21977));
  jand g21844(.dina(n21974), .dinb(n4941), .dout(n21978));
  jand g21845(.dina(n21340), .dinb(n4696), .dout(n21979));
  jand g21846(.dina(n21197), .dinb(n4701), .dout(n21980));
  jor  g21847(.dina(n21980), .dinb(n21979), .dout(n21981));
  jor  g21848(.dina(n21981), .dinb(n21978), .dout(n21982));
  jor  g21849(.dina(n21982), .dinb(n21977), .dout(n21983));
  jxor g21850(.dina(n21983), .dinb(n4713), .dout(n21984));
  jxor g21851(.dina(n21984), .dinb(n21869), .dout(n21985));
  jnot g21852(.din(n21985), .dout(n21986));
  jxor g21853(.dina(n21986), .dinb(n21724), .dout(n21987));
  jnot g21854(.din(n21987), .dout(n21988));
  jor  g21855(.dina(n22046), .dinb(n21881), .dout(n21989));
  jand g21856(.dina(n21966), .dinb(n21889), .dout(n21990));
  jnot g21857(.din(n21990), .dout(n21991));
  jand g21858(.dina(n21991), .dinb(n21989), .dout(n21992));
  jnot g21859(.din(n21992), .dout(n21993));
  jor  g21860(.dina(n21944), .dinb(n21936), .dout(n21994));
  jor  g21861(.dina(n21954), .dinb(n21946), .dout(n21995));
  jand g21862(.dina(n21995), .dinb(n21994), .dout(n21996));
  jnot g21863(.din(n21996), .dout(n21997));
  jand g21864(.dina(n21928), .dinb(n21899), .dout(n21998));
  jnot g21865(.din(n21998), .dout(n21999));
  jor  g21866(.dina(n21934), .dinb(n21930), .dout(n22000));
  jand g21867(.dina(n22000), .dinb(n21999), .dout(n22001));
  jnot g21868(.din(n22001), .dout(n22002));
  jand g21869(.dina(n14579), .dinb(n5076), .dout(n22003));
  jand g21870(.dina(n14448), .dinb(n5084), .dout(n22004));
  jand g21871(.dina(n14249), .dinb(n5082), .dout(n22005));
  jand g21872(.dina(n13614), .dinb(n6050), .dout(n22006));
  jor  g21873(.dina(n22006), .dinb(n22005), .dout(n22007));
  jor  g21874(.dina(n22007), .dinb(n22004), .dout(n22008));
  jor  g21875(.dina(n22008), .dinb(n22003), .dout(n22009));
  jor  g21876(.dina(n21926), .dinb(n21280), .dout(n22010));
  jand g21877(.dina(n21927), .dinb(n21906), .dout(n22011));
  jnot g21878(.din(n22011), .dout(n22012));
  jand g21879(.dina(n22012), .dinb(n22010), .dout(n22013));
  jnot g21880(.din(n22013), .dout(n22014));
  jnot g21881(.din(n1029), .dout(n22015));
  jand g21882(.dina(n2713), .dinb(n2052), .dout(n22016));
  jand g21883(.dina(n22016), .dinb(n22015), .dout(n22017));
  jand g21884(.dina(n1367), .dinb(n1233), .dout(n22018));
  jand g21885(.dina(n534), .dinb(n1226), .dout(n22019));
  jand g21886(.dina(n22019), .dinb(n2020), .dout(n22020));
  jand g21887(.dina(n22020), .dinb(n22018), .dout(n22021));
  jand g21888(.dina(n10413), .dinb(n4440), .dout(n22022));
  jand g21889(.dina(n22022), .dinb(n480), .dout(n22023));
  jand g21890(.dina(n22023), .dinb(n22021), .dout(n22024));
  jand g21891(.dina(n22024), .dinb(n22017), .dout(n22025));
  jand g21892(.dina(n6366), .dinb(n1525), .dout(n22026));
  jand g21893(.dina(n22026), .dinb(n3811), .dout(n22027));
  jand g21894(.dina(n22027), .dinb(n22025), .dout(n22028));
  jand g21895(.dina(n10530), .dinb(n683), .dout(n22029));
  jand g21896(.dina(n22029), .dinb(n11538), .dout(n22030));
  jand g21897(.dina(n22030), .dinb(n1562), .dout(n22031));
  jand g21898(.dina(n22031), .dinb(n22028), .dout(n22032));
  jand g21899(.dina(n582), .dinb(n175), .dout(n22033));
  jand g21900(.dina(n18187), .dinb(n4639), .dout(n22034));
  jand g21901(.dina(n22034), .dinb(n22033), .dout(n22035));
  jand g21902(.dina(n3198), .dinb(n7503), .dout(n22036));
  jand g21903(.dina(n22036), .dinb(n4588), .dout(n22037));
  jand g21904(.dina(n22037), .dinb(n22035), .dout(n22038));
  jand g21905(.dina(n22038), .dinb(n1357), .dout(n22039));
  jand g21906(.dina(n22039), .dinb(n4439), .dout(n22040));
  jand g21907(.dina(n22040), .dinb(n22032), .dout(n22041));
  jand g21908(.dina(n22041), .dinb(n3129), .dout(n22042));
  jxor g21909(.dina(n22042), .dinb(n21279), .dout(n22043));
  jand g21910(.dina(n2186), .dinb(n2184), .dout(n22044));
  jor  g21911(.dina(n22044), .dinb(n17301), .dout(n22045));
  jxor g21912(.dina(n22045), .dinb(\a[20] ), .dout(n22046));
  jxor g21913(.dina(n22046), .dinb(n22043), .dout(n22047));
  jxor g21914(.dina(n22047), .dinb(n22014), .dout(n22048));
  jxor g21915(.dina(n22048), .dinb(n22009), .dout(n22049));
  jxor g21916(.dina(n22049), .dinb(n22002), .dout(n22050));
  jnot g21917(.din(n22050), .dout(n22051));
  jand g21918(.dina(n15317), .dinb(n2936), .dout(n22052));
  jand g21919(.dina(n15315), .dinb(n2943), .dout(n22053));
  jand g21920(.dina(n14549), .dinb(n2940), .dout(n22054));
  jand g21921(.dina(n14447), .dinb(n3684), .dout(n22055));
  jor  g21922(.dina(n22055), .dinb(n22054), .dout(n22056));
  jor  g21923(.dina(n22056), .dinb(n22053), .dout(n22057));
  jor  g21924(.dina(n22057), .dinb(n22052), .dout(n22058));
  jxor g21925(.dina(n22058), .dinb(n93), .dout(n22059));
  jxor g21926(.dina(n22059), .dinb(n22051), .dout(n22060));
  jnot g21927(.din(n22060), .dout(n22061));
  jand g21928(.dina(n16084), .dinb(n71), .dout(n22062));
  jand g21929(.dina(n15829), .dinb(n731), .dout(n22063));
  jand g21930(.dina(n16082), .dinb(n796), .dout(n22064));
  jor  g21931(.dina(n22064), .dinb(n22063), .dout(n22065));
  jand g21932(.dina(n15567), .dinb(n1806), .dout(n22066));
  jor  g21933(.dina(n22066), .dinb(n22065), .dout(n22067));
  jor  g21934(.dina(n22067), .dinb(n22062), .dout(n22068));
  jxor g21935(.dina(n22068), .dinb(n77), .dout(n22069));
  jxor g21936(.dina(n22069), .dinb(n22061), .dout(n22070));
  jxor g21937(.dina(n22070), .dinb(n21997), .dout(n22071));
  jand g21938(.dina(n21955), .dinb(n21894), .dout(n22072));
  jnot g21939(.din(n22072), .dout(n22073));
  jor  g21940(.dina(n21965), .dinb(n21957), .dout(n22074));
  jand g21941(.dina(n22074), .dinb(n22073), .dout(n22075));
  jand g21942(.dina(n16930), .dinb(n806), .dout(n22076));
  jand g21943(.dina(n16592), .dinb(n1612), .dout(n22077));
  jand g21944(.dina(n16928), .dinb(n1620), .dout(n22078));
  jor  g21945(.dina(n22078), .dinb(n22077), .dout(n22079));
  jand g21946(.dina(n16343), .dinb(n1644), .dout(n22080));
  jor  g21947(.dina(n22080), .dinb(n22079), .dout(n22081));
  jor  g21948(.dina(n22081), .dinb(n22076), .dout(n22082));
  jxor g21949(.dina(n22082), .dinb(n65), .dout(n22083));
  jxor g21950(.dina(n22083), .dinb(n22075), .dout(n22084));
  jxor g21951(.dina(n22084), .dinb(n22071), .dout(n22085));
  jand g21952(.dina(n22085), .dinb(n21993), .dout(n22086));
  jnot g21953(.din(n22086), .dout(n22087));
  jand g21954(.dina(n21967), .dinb(n21877), .dout(n22088));
  jnot g21955(.din(n22088), .dout(n22089));
  jor  g21956(.dina(n21973), .dinb(n21969), .dout(n22090));
  jand g21957(.dina(n22090), .dinb(n22089), .dout(n22091));
  jxor g21958(.dina(n22085), .dinb(n21993), .dout(n22092));
  jnot g21959(.din(n22092), .dout(n22093));
  jor  g21960(.dina(n22093), .dinb(n22091), .dout(n22094));
  jand g21961(.dina(n22094), .dinb(n22087), .dout(n22095));
  jor  g21962(.dina(n22083), .dinb(n22075), .dout(n22096));
  jand g21963(.dina(n22084), .dinb(n22071), .dout(n22097));
  jnot g21964(.din(n22097), .dout(n22098));
  jand g21965(.dina(n22098), .dinb(n22096), .dout(n22099));
  jnot g21966(.din(n22099), .dout(n22100));
  jor  g21967(.dina(n22069), .dinb(n22061), .dout(n22101));
  jand g21968(.dina(n22070), .dinb(n21997), .dout(n22102));
  jnot g21969(.din(n22102), .dout(n22103));
  jand g21970(.dina(n22103), .dinb(n22101), .dout(n22104));
  jnot g21971(.din(n22104), .dout(n22105));
  jand g21972(.dina(n22049), .dinb(n22002), .dout(n22106));
  jnot g21973(.din(n22106), .dout(n22107));
  jor  g21974(.dina(n22059), .dinb(n22051), .dout(n22108));
  jand g21975(.dina(n22108), .dinb(n22107), .dout(n22109));
  jnot g21976(.din(n22109), .dout(n22110));
  jand g21977(.dina(n22047), .dinb(n22014), .dout(n22111));
  jand g21978(.dina(n22048), .dinb(n22009), .dout(n22112));
  jor  g21979(.dina(n22112), .dinb(n22111), .dout(n22113));
  jnot g21980(.din(n16573), .dout(n22114));
  jor  g21981(.dina(n22042), .dinb(n21279), .dout(n22115));
  jand g21982(.dina(n22046), .dinb(n22043), .dout(n22116));
  jnot g21983(.din(n22116), .dout(n22117));
  jand g21984(.dina(n22117), .dinb(n22115), .dout(n22118));
  jxor g21985(.dina(n22118), .dinb(n22114), .dout(n22119));
  jand g21986(.dina(n14562), .dinb(n5076), .dout(n22120));
  jand g21987(.dina(n14447), .dinb(n5084), .dout(n22121));
  jand g21988(.dina(n14249), .dinb(n6050), .dout(n22122));
  jand g21989(.dina(n14448), .dinb(n5082), .dout(n22123));
  jor  g21990(.dina(n22123), .dinb(n22122), .dout(n22124));
  jor  g21991(.dina(n22124), .dinb(n22121), .dout(n22125));
  jor  g21992(.dina(n22125), .dinb(n22120), .dout(n22126));
  jxor g21993(.dina(n22126), .dinb(n22119), .dout(n22127));
  jxor g21994(.dina(n22127), .dinb(n22113), .dout(n22128));
  jnot g21995(.din(n22128), .dout(n22129));
  jand g21996(.dina(n15569), .dinb(n2936), .dout(n22130));
  jand g21997(.dina(n15315), .dinb(n2940), .dout(n22131));
  jand g21998(.dina(n15567), .dinb(n2943), .dout(n22132));
  jor  g21999(.dina(n22132), .dinb(n22131), .dout(n22133));
  jand g22000(.dina(n14549), .dinb(n3684), .dout(n22134));
  jor  g22001(.dina(n22134), .dinb(n22133), .dout(n22135));
  jor  g22002(.dina(n22135), .dinb(n22130), .dout(n22136));
  jxor g22003(.dina(n22136), .dinb(n93), .dout(n22137));
  jxor g22004(.dina(n22137), .dinb(n22129), .dout(n22138));
  jxor g22005(.dina(n22138), .dinb(n22110), .dout(n22139));
  jnot g22006(.din(n22139), .dout(n22140));
  jand g22007(.dina(n16345), .dinb(n71), .dout(n22141));
  jand g22008(.dina(n16082), .dinb(n731), .dout(n22142));
  jand g22009(.dina(n16343), .dinb(n796), .dout(n22143));
  jor  g22010(.dina(n22143), .dinb(n22142), .dout(n22144));
  jand g22011(.dina(n15829), .dinb(n1806), .dout(n22145));
  jor  g22012(.dina(n22145), .dinb(n22144), .dout(n22146));
  jor  g22013(.dina(n22146), .dinb(n22141), .dout(n22147));
  jxor g22014(.dina(n22147), .dinb(n77), .dout(n22148));
  jxor g22015(.dina(n22148), .dinb(n22140), .dout(n22149));
  jxor g22016(.dina(n22149), .dinb(n22105), .dout(n22150));
  jnot g22017(.din(n22150), .dout(n22151));
  jand g22018(.dina(n17312), .dinb(n806), .dout(n22152));
  jand g22019(.dina(n16928), .dinb(n1612), .dout(n22153));
  jand g22020(.dina(n16592), .dinb(n1644), .dout(n22154));
  jand g22021(.dina(n16924), .dinb(n1620), .dout(n22155));
  jor  g22022(.dina(n22155), .dinb(n22154), .dout(n22156));
  jor  g22023(.dina(n22156), .dinb(n22153), .dout(n22157));
  jor  g22024(.dina(n22157), .dinb(n22152), .dout(n22158));
  jxor g22025(.dina(n22158), .dinb(n65), .dout(n22159));
  jxor g22026(.dina(n22159), .dinb(n22151), .dout(n22160));
  jxor g22027(.dina(n22160), .dinb(n22100), .dout(n22161));
  jnot g22028(.din(n22161), .dout(n22162));
  jxor g22029(.dina(n22162), .dinb(n22095), .dout(n22163));
  jxor g22030(.dina(n22093), .dinb(n22091), .dout(n22164));
  jand g22031(.dina(n22164), .dinb(n22163), .dout(n22165));
  jand g22032(.dina(n22164), .dinb(n21974), .dout(n22166));
  jand g22033(.dina(n21974), .dinb(n21340), .dout(n22167));
  jand g22034(.dina(n21975), .dinb(n21872), .dout(n22168));
  jor  g22035(.dina(n22168), .dinb(n22167), .dout(n22169));
  jxor g22036(.dina(n22164), .dinb(n21974), .dout(n22170));
  jand g22037(.dina(n22170), .dinb(n22169), .dout(n22171));
  jor  g22038(.dina(n22171), .dinb(n22166), .dout(n22172));
  jxor g22039(.dina(n22164), .dinb(n22163), .dout(n22173));
  jand g22040(.dina(n22173), .dinb(n22172), .dout(n22174));
  jor  g22041(.dina(n22174), .dinb(n22165), .dout(n22175));
  jand g22042(.dina(n22149), .dinb(n22105), .dout(n22176));
  jnot g22043(.din(n22176), .dout(n22177));
  jor  g22044(.dina(n22159), .dinb(n22151), .dout(n22178));
  jand g22045(.dina(n22178), .dinb(n22177), .dout(n22179));
  jnot g22046(.din(n22179), .dout(n22180));
  jand g22047(.dina(n22138), .dinb(n22110), .dout(n22181));
  jnot g22048(.din(n22181), .dout(n22182));
  jor  g22049(.dina(n22148), .dinb(n22140), .dout(n22183));
  jand g22050(.dina(n22183), .dinb(n22182), .dout(n22184));
  jand g22051(.dina(n1621), .dinb(n1613), .dout(n22185));
  jxor g22052(.dina(n22912), .dinb(n22184), .dout(n22192));
  jand g22053(.dina(n22127), .dinb(n22113), .dout(n22193));
  jnot g22054(.din(n22193), .dout(n22194));
  jor  g22055(.dina(n22137), .dinb(n22129), .dout(n22195));
  jand g22056(.dina(n22195), .dinb(n22194), .dout(n22196));
  jnot g22057(.din(n22196), .dout(n22197));
  jand g22058(.dina(n14551), .dinb(n5076), .dout(n22198));
  jand g22059(.dina(n14549), .dinb(n5084), .dout(n22199));
  jand g22060(.dina(n14447), .dinb(n5082), .dout(n22200));
  jand g22061(.dina(n14448), .dinb(n6050), .dout(n22201));
  jor  g22062(.dina(n22201), .dinb(n22200), .dout(n22202));
  jor  g22063(.dina(n22202), .dinb(n22199), .dout(n22203));
  jor  g22064(.dina(n22203), .dinb(n22198), .dout(n22204));
  jor  g22065(.dina(n22118), .dinb(n22114), .dout(n22205));
  jand g22066(.dina(n22126), .dinb(n22119), .dout(n22206));
  jnot g22067(.din(n22206), .dout(n22207));
  jand g22068(.dina(n22207), .dinb(n22205), .dout(n22208));
  jnot g22069(.din(n22208), .dout(n22209));
  jand g22070(.dina(n6439), .dinb(n178), .dout(n22210));
  jand g22071(.dina(n22210), .dinb(n588), .dout(n22211));
  jand g22072(.dina(n22211), .dinb(n1552), .dout(n22212));
  jand g22073(.dina(n22212), .dinb(n21258), .dout(n22213));
  jand g22074(.dina(n13536), .dinb(n6317), .dout(n22214));
  jand g22075(.dina(n1698), .dinb(n1713), .dout(n22215));
  jand g22076(.dina(n22215), .dinb(n1580), .dout(n22216));
  jand g22077(.dina(n22216), .dinb(n22214), .dout(n22217));
  jand g22078(.dina(n3827), .dinb(n630), .dout(n22218));
  jand g22079(.dina(n22218), .dinb(n13541), .dout(n22219));
  jand g22080(.dina(n22219), .dinb(n11358), .dout(n22220));
  jand g22081(.dina(n6151), .dinb(n1017), .dout(n22221));
  jand g22082(.dina(n713), .dinb(n1430), .dout(n22222));
  jand g22083(.dina(n22222), .dinb(n1236), .dout(n22223));
  jand g22084(.dina(n22223), .dinb(n22221), .dout(n22224));
  jand g22085(.dina(n6280), .dinb(n680), .dout(n22225));
  jand g22086(.dina(n22225), .dinb(n22224), .dout(n22226));
  jand g22087(.dina(n22226), .dinb(n22220), .dout(n22227));
  jand g22088(.dina(n1731), .dinb(n1188), .dout(n22228));
  jand g22089(.dina(n22228), .dinb(n9747), .dout(n22229));
  jand g22090(.dina(n22229), .dinb(n22227), .dout(n22230));
  jand g22091(.dina(n22230), .dinb(n22217), .dout(n22231));
  jand g22092(.dina(n22231), .dinb(n11215), .dout(n22232));
  jand g22093(.dina(n22232), .dinb(n22213), .dout(n22233));
  jxor g22094(.dina(n22233), .dinb(n22114), .dout(n22234));
  jxor g22095(.dina(n22234), .dinb(n22209), .dout(n22235));
  jxor g22096(.dina(n22235), .dinb(n22204), .dout(n22236));
  jnot g22097(.din(n22236), .dout(n22237));
  jand g22098(.dina(n15831), .dinb(n2936), .dout(n22238));
  jand g22099(.dina(n15567), .dinb(n2940), .dout(n22239));
  jand g22100(.dina(n15829), .dinb(n2943), .dout(n22240));
  jor  g22101(.dina(n22240), .dinb(n22239), .dout(n22241));
  jand g22102(.dina(n15315), .dinb(n3684), .dout(n22242));
  jor  g22103(.dina(n22242), .dinb(n22241), .dout(n22243));
  jor  g22104(.dina(n22243), .dinb(n22238), .dout(n22244));
  jxor g22105(.dina(n22244), .dinb(n93), .dout(n22245));
  jxor g22106(.dina(n22245), .dinb(n22237), .dout(n22246));
  jxor g22107(.dina(n22246), .dinb(n22197), .dout(n22247));
  jnot g22108(.din(n22247), .dout(n22248));
  jand g22109(.dina(n16594), .dinb(n71), .dout(n22249));
  jand g22110(.dina(n16592), .dinb(n796), .dout(n22250));
  jand g22111(.dina(n16343), .dinb(n731), .dout(n22251));
  jand g22112(.dina(n16082), .dinb(n1806), .dout(n22252));
  jor  g22113(.dina(n22252), .dinb(n22251), .dout(n22253));
  jor  g22114(.dina(n22253), .dinb(n22250), .dout(n22254));
  jor  g22115(.dina(n22254), .dinb(n22249), .dout(n22255));
  jxor g22116(.dina(n22255), .dinb(n77), .dout(n22256));
  jxor g22117(.dina(n22256), .dinb(n22248), .dout(n22257));
  jxor g22118(.dina(n22257), .dinb(n22192), .dout(n22258));
  jxor g22119(.dina(n22258), .dinb(n22180), .dout(n22259));
  jnot g22120(.din(n22259), .dout(n22260));
  jand g22121(.dina(n22160), .dinb(n22100), .dout(n22261));
  jnot g22122(.din(n22261), .dout(n22262));
  jor  g22123(.dina(n22162), .dinb(n22095), .dout(n22263));
  jand g22124(.dina(n22263), .dinb(n22262), .dout(n22264));
  jxor g22125(.dina(n22264), .dinb(n22260), .dout(n22265));
  jxor g22126(.dina(n22265), .dinb(n22163), .dout(n22266));
  jxor g22127(.dina(n22266), .dinb(n22175), .dout(n22267));
  jand g22128(.dina(n22267), .dinb(n5280), .dout(n22268));
  jand g22129(.dina(n22265), .dinb(n5814), .dout(n22269));
  jand g22130(.dina(n22163), .dinb(n5531), .dout(n22270));
  jand g22131(.dina(n22164), .dinb(n5536), .dout(n22271));
  jor  g22132(.dina(n22271), .dinb(n22270), .dout(n22272));
  jor  g22133(.dina(n22272), .dinb(n22269), .dout(n22273));
  jor  g22134(.dina(n22273), .dinb(n22268), .dout(n22274));
  jxor g22135(.dina(n22274), .dinb(n5277), .dout(n22275));
  jor  g22136(.dina(n22275), .dinb(n21988), .dout(n22276));
  jxor g22137(.dina(n21722), .dinb(n21720), .dout(n22277));
  jnot g22138(.din(n22277), .dout(n22278));
  jxor g22139(.dina(n22173), .dinb(n22172), .dout(n22279));
  jand g22140(.dina(n22279), .dinb(n5280), .dout(n22280));
  jand g22141(.dina(n22163), .dinb(n5814), .dout(n22281));
  jand g22142(.dina(n22164), .dinb(n5531), .dout(n22282));
  jand g22143(.dina(n21974), .dinb(n5536), .dout(n22283));
  jor  g22144(.dina(n22283), .dinb(n22282), .dout(n22284));
  jor  g22145(.dina(n22284), .dinb(n22281), .dout(n22285));
  jor  g22146(.dina(n22285), .dinb(n22280), .dout(n22286));
  jxor g22147(.dina(n22286), .dinb(\a[5] ), .dout(n22287));
  jand g22148(.dina(n22287), .dinb(n22278), .dout(n22288));
  jnot g22149(.din(n22288), .dout(n22289));
  jxor g22150(.dina(n21718), .dinb(n21717), .dout(n22290));
  jxor g22151(.dina(n22170), .dinb(n22169), .dout(n22291));
  jand g22152(.dina(n22291), .dinb(n5280), .dout(n22292));
  jand g22153(.dina(n22164), .dinb(n5814), .dout(n22293));
  jand g22154(.dina(n21974), .dinb(n5531), .dout(n22294));
  jand g22155(.dina(n21340), .dinb(n5536), .dout(n22295));
  jor  g22156(.dina(n22295), .dinb(n22294), .dout(n22296));
  jor  g22157(.dina(n22296), .dinb(n22293), .dout(n22297));
  jor  g22158(.dina(n22297), .dinb(n22292), .dout(n22298));
  jxor g22159(.dina(n22298), .dinb(\a[5] ), .dout(n22299));
  jand g22160(.dina(n22299), .dinb(n22290), .dout(n22300));
  jnot g22161(.din(n22300), .dout(n22301));
  jxor g22162(.dina(n21715), .dinb(n21714), .dout(n22302));
  jnot g22163(.din(n22302), .dout(n22303));
  jand g22164(.dina(n21976), .dinb(n5280), .dout(n22304));
  jand g22165(.dina(n21340), .dinb(n5531), .dout(n22305));
  jand g22166(.dina(n21974), .dinb(n5814), .dout(n22306));
  jor  g22167(.dina(n22306), .dinb(n22305), .dout(n22307));
  jand g22168(.dina(n21197), .dinb(n5536), .dout(n22308));
  jor  g22169(.dina(n22308), .dinb(n22307), .dout(n22309));
  jor  g22170(.dina(n22309), .dinb(n22304), .dout(n22310));
  jxor g22171(.dina(n22310), .dinb(n5277), .dout(n22311));
  jor  g22172(.dina(n22311), .dinb(n22303), .dout(n22312));
  jxor g22173(.dina(n21712), .dinb(n21711), .dout(n22313));
  jnot g22174(.din(n22313), .dout(n22314));
  jand g22175(.dina(n21342), .dinb(n5280), .dout(n22315));
  jand g22176(.dina(n21340), .dinb(n5814), .dout(n22316));
  jand g22177(.dina(n21197), .dinb(n5531), .dout(n22317));
  jand g22178(.dina(n21198), .dinb(n5536), .dout(n22318));
  jor  g22179(.dina(n22318), .dinb(n22317), .dout(n22319));
  jor  g22180(.dina(n22319), .dinb(n22316), .dout(n22320));
  jor  g22181(.dina(n22320), .dinb(n22315), .dout(n22321));
  jxor g22182(.dina(n22321), .dinb(n5277), .dout(n22322));
  jor  g22183(.dina(n22322), .dinb(n22314), .dout(n22323));
  jxor g22184(.dina(n21708), .dinb(n21707), .dout(n22324));
  jand g22185(.dina(n21355), .dinb(n5280), .dout(n22325));
  jand g22186(.dina(n21198), .dinb(n5531), .dout(n22326));
  jand g22187(.dina(n21197), .dinb(n5814), .dout(n22327));
  jor  g22188(.dina(n22327), .dinb(n22326), .dout(n22328));
  jand g22189(.dina(n20947), .dinb(n5536), .dout(n22329));
  jor  g22190(.dina(n22329), .dinb(n22328), .dout(n22330));
  jor  g22191(.dina(n22330), .dinb(n22325), .dout(n22331));
  jxor g22192(.dina(n22331), .dinb(n5277), .dout(n22332));
  jor  g22193(.dina(n22332), .dinb(n22324), .dout(n22333));
  jnot g22194(.din(n22333), .dout(n22334));
  jnot g22195(.din(n21705), .dout(n22335));
  jxor g22196(.dina(n22335), .dinb(n21704), .dout(n22336));
  jand g22197(.dina(n21367), .dinb(n5280), .dout(n22337));
  jand g22198(.dina(n20947), .dinb(n5531), .dout(n22338));
  jand g22199(.dina(n21198), .dinb(n5814), .dout(n22339));
  jor  g22200(.dina(n22339), .dinb(n22338), .dout(n22340));
  jand g22201(.dina(n20344), .dinb(n5536), .dout(n22341));
  jor  g22202(.dina(n22341), .dinb(n22340), .dout(n22342));
  jor  g22203(.dina(n22342), .dinb(n22337), .dout(n22343));
  jxor g22204(.dina(n22343), .dinb(n5277), .dout(n22344));
  jor  g22205(.dina(n22344), .dinb(n22336), .dout(n22345));
  jnot g22206(.din(n22345), .dout(n22346));
  jnot g22207(.din(n21702), .dout(n22347));
  jxor g22208(.dina(n22347), .dinb(n21701), .dout(n22348));
  jand g22209(.dina(n20949), .dinb(n5280), .dout(n22349));
  jand g22210(.dina(n20344), .dinb(n5531), .dout(n22350));
  jand g22211(.dina(n20947), .dinb(n5814), .dout(n22351));
  jor  g22212(.dina(n22351), .dinb(n22350), .dout(n22352));
  jand g22213(.dina(n20204), .dinb(n5536), .dout(n22353));
  jor  g22214(.dina(n22353), .dinb(n22352), .dout(n22354));
  jor  g22215(.dina(n22354), .dinb(n22349), .dout(n22355));
  jxor g22216(.dina(n22355), .dinb(n5277), .dout(n22356));
  jor  g22217(.dina(n22356), .dinb(n22348), .dout(n22357));
  jnot g22218(.din(n22357), .dout(n22358));
  jnot g22219(.din(n21699), .dout(n22359));
  jxor g22220(.dina(n22359), .dinb(n21698), .dout(n22360));
  jand g22221(.dina(n20346), .dinb(n5280), .dout(n22361));
  jand g22222(.dina(n20344), .dinb(n5814), .dout(n22362));
  jand g22223(.dina(n20204), .dinb(n5531), .dout(n22363));
  jand g22224(.dina(n20205), .dinb(n5536), .dout(n22364));
  jor  g22225(.dina(n22364), .dinb(n22363), .dout(n22365));
  jor  g22226(.dina(n22365), .dinb(n22362), .dout(n22366));
  jor  g22227(.dina(n22366), .dinb(n22361), .dout(n22367));
  jxor g22228(.dina(n22367), .dinb(n5277), .dout(n22368));
  jor  g22229(.dina(n22368), .dinb(n22360), .dout(n22369));
  jnot g22230(.din(n22369), .dout(n22370));
  jxor g22231(.dina(n21695), .dinb(n21694), .dout(n22371));
  jand g22232(.dina(n20358), .dinb(n5280), .dout(n22372));
  jand g22233(.dina(n20205), .dinb(n5531), .dout(n22373));
  jand g22234(.dina(n20204), .dinb(n5814), .dout(n22374));
  jor  g22235(.dina(n22374), .dinb(n22373), .dout(n22375));
  jand g22236(.dina(n19922), .dinb(n5536), .dout(n22376));
  jor  g22237(.dina(n22376), .dinb(n22375), .dout(n22377));
  jor  g22238(.dina(n22377), .dinb(n22372), .dout(n22378));
  jxor g22239(.dina(n22378), .dinb(n5277), .dout(n22379));
  jor  g22240(.dina(n22379), .dinb(n22371), .dout(n22380));
  jnot g22241(.din(n22380), .dout(n22381));
  jxor g22242(.dina(n21692), .dinb(n21690), .dout(n22382));
  jnot g22243(.din(n22382), .dout(n22383));
  jand g22244(.dina(n20371), .dinb(n5280), .dout(n22384));
  jand g22245(.dina(n19922), .dinb(n5531), .dout(n22385));
  jand g22246(.dina(n20205), .dinb(n5814), .dout(n22386));
  jor  g22247(.dina(n22386), .dinb(n22385), .dout(n22387));
  jand g22248(.dina(n19373), .dinb(n5536), .dout(n22388));
  jor  g22249(.dina(n22388), .dinb(n22387), .dout(n22389));
  jor  g22250(.dina(n22389), .dinb(n22384), .dout(n22390));
  jxor g22251(.dina(n22390), .dinb(n5277), .dout(n22391));
  jor  g22252(.dina(n22391), .dinb(n22383), .dout(n22392));
  jnot g22253(.din(n22392), .dout(n22393));
  jxor g22254(.dina(n21688), .dinb(n21686), .dout(n22394));
  jnot g22255(.din(n22394), .dout(n22395));
  jand g22256(.dina(n19924), .dinb(n5280), .dout(n22396));
  jand g22257(.dina(n19373), .dinb(n5531), .dout(n22397));
  jand g22258(.dina(n19922), .dinb(n5814), .dout(n22398));
  jor  g22259(.dina(n22398), .dinb(n22397), .dout(n22399));
  jand g22260(.dina(n19219), .dinb(n5536), .dout(n22400));
  jor  g22261(.dina(n22400), .dinb(n22399), .dout(n22401));
  jor  g22262(.dina(n22401), .dinb(n22396), .dout(n22402));
  jxor g22263(.dina(n22402), .dinb(n5277), .dout(n22403));
  jor  g22264(.dina(n22403), .dinb(n22395), .dout(n22404));
  jnot g22265(.din(n22404), .dout(n22405));
  jxor g22266(.dina(n21684), .dinb(n21682), .dout(n22406));
  jand g22267(.dina(n19375), .dinb(n5280), .dout(n22407));
  jand g22268(.dina(n19373), .dinb(n5814), .dout(n22408));
  jand g22269(.dina(n19219), .dinb(n5531), .dout(n22409));
  jand g22270(.dina(n19220), .dinb(n5536), .dout(n22410));
  jor  g22271(.dina(n22410), .dinb(n22409), .dout(n22411));
  jor  g22272(.dina(n22411), .dinb(n22408), .dout(n22412));
  jor  g22273(.dina(n22412), .dinb(n22407), .dout(n22413));
  jxor g22274(.dina(n22413), .dinb(\a[5] ), .dout(n22414));
  jand g22275(.dina(n22414), .dinb(n22406), .dout(n22415));
  jxor g22276(.dina(n21680), .dinb(n21678), .dout(n22416));
  jnot g22277(.din(n22416), .dout(n22417));
  jand g22278(.dina(n19387), .dinb(n5280), .dout(n22418));
  jand g22279(.dina(n19220), .dinb(n5531), .dout(n22419));
  jand g22280(.dina(n19219), .dinb(n5814), .dout(n22420));
  jor  g22281(.dina(n22420), .dinb(n22419), .dout(n22421));
  jand g22282(.dina(n18914), .dinb(n5536), .dout(n22422));
  jor  g22283(.dina(n22422), .dinb(n22421), .dout(n22423));
  jor  g22284(.dina(n22423), .dinb(n22418), .dout(n22424));
  jxor g22285(.dina(n22424), .dinb(n5277), .dout(n22425));
  jor  g22286(.dina(n22425), .dinb(n22417), .dout(n22426));
  jnot g22287(.din(n22426), .dout(n22427));
  jxor g22288(.dina(n21675), .dinb(n21674), .dout(n22428));
  jnot g22289(.din(n22428), .dout(n22429));
  jand g22290(.dina(n19399), .dinb(n5280), .dout(n22430));
  jand g22291(.dina(n19220), .dinb(n5814), .dout(n22431));
  jand g22292(.dina(n18914), .dinb(n5531), .dout(n22432));
  jand g22293(.dina(n18488), .dinb(n5536), .dout(n22433));
  jor  g22294(.dina(n22433), .dinb(n22432), .dout(n22434));
  jor  g22295(.dina(n22434), .dinb(n22431), .dout(n22435));
  jor  g22296(.dina(n22435), .dinb(n22430), .dout(n22436));
  jxor g22297(.dina(n22436), .dinb(n5277), .dout(n22437));
  jor  g22298(.dina(n22437), .dinb(n22429), .dout(n22438));
  jnot g22299(.din(n22438), .dout(n22439));
  jxor g22300(.dina(n21670), .dinb(n21669), .dout(n22440));
  jnot g22301(.din(n22440), .dout(n22441));
  jand g22302(.dina(n18916), .dinb(n5280), .dout(n22442));
  jand g22303(.dina(n18488), .dinb(n5531), .dout(n22443));
  jand g22304(.dina(n18914), .dinb(n5814), .dout(n22444));
  jor  g22305(.dina(n22444), .dinb(n22443), .dout(n22445));
  jand g22306(.dina(n18292), .dinb(n5536), .dout(n22446));
  jor  g22307(.dina(n22446), .dinb(n22445), .dout(n22447));
  jor  g22308(.dina(n22447), .dinb(n22442), .dout(n22448));
  jxor g22309(.dina(n22448), .dinb(n5277), .dout(n22449));
  jor  g22310(.dina(n22449), .dinb(n22441), .dout(n22450));
  jnot g22311(.din(n22450), .dout(n22451));
  jxor g22312(.dina(n21665), .dinb(n21664), .dout(n22452));
  jnot g22313(.din(n22452), .dout(n22453));
  jand g22314(.dina(n18490), .dinb(n5280), .dout(n22454));
  jand g22315(.dina(n18488), .dinb(n5814), .dout(n22455));
  jand g22316(.dina(n18292), .dinb(n5531), .dout(n22456));
  jand g22317(.dina(n18293), .dinb(n5536), .dout(n22457));
  jor  g22318(.dina(n22457), .dinb(n22456), .dout(n22458));
  jor  g22319(.dina(n22458), .dinb(n22455), .dout(n22459));
  jor  g22320(.dina(n22459), .dinb(n22454), .dout(n22460));
  jxor g22321(.dina(n22460), .dinb(n5277), .dout(n22461));
  jor  g22322(.dina(n22461), .dinb(n22453), .dout(n22462));
  jnot g22323(.din(n22462), .dout(n22463));
  jxor g22324(.dina(n21660), .dinb(n21659), .dout(n22464));
  jnot g22325(.din(n22464), .dout(n22465));
  jand g22326(.dina(n18502), .dinb(n5280), .dout(n22466));
  jand g22327(.dina(n18293), .dinb(n5531), .dout(n22467));
  jand g22328(.dina(n18292), .dinb(n5814), .dout(n22468));
  jor  g22329(.dina(n22468), .dinb(n22467), .dout(n22469));
  jand g22330(.dina(n17942), .dinb(n5536), .dout(n22470));
  jor  g22331(.dina(n22470), .dinb(n22469), .dout(n22471));
  jor  g22332(.dina(n22471), .dinb(n22466), .dout(n22472));
  jxor g22333(.dina(n22472), .dinb(n5277), .dout(n22473));
  jor  g22334(.dina(n22473), .dinb(n22465), .dout(n22474));
  jnot g22335(.din(n22474), .dout(n22475));
  jxor g22336(.dina(n21655), .dinb(n21654), .dout(n22476));
  jnot g22337(.din(n22476), .dout(n22477));
  jand g22338(.dina(n18514), .dinb(n5280), .dout(n22478));
  jand g22339(.dina(n17942), .dinb(n5531), .dout(n22479));
  jand g22340(.dina(n18293), .dinb(n5814), .dout(n22480));
  jor  g22341(.dina(n22480), .dinb(n22479), .dout(n22481));
  jand g22342(.dina(n17535), .dinb(n5536), .dout(n22482));
  jor  g22343(.dina(n22482), .dinb(n22481), .dout(n22483));
  jor  g22344(.dina(n22483), .dinb(n22478), .dout(n22484));
  jxor g22345(.dina(n22484), .dinb(n5277), .dout(n22485));
  jor  g22346(.dina(n22485), .dinb(n22477), .dout(n22486));
  jnot g22347(.din(n22486), .dout(n22487));
  jxor g22348(.dina(n21650), .dinb(n21649), .dout(n22488));
  jnot g22349(.din(n22488), .dout(n22489));
  jand g22350(.dina(n17944), .dinb(n5280), .dout(n22490));
  jand g22351(.dina(n17942), .dinb(n5814), .dout(n22491));
  jand g22352(.dina(n17535), .dinb(n5531), .dout(n22492));
  jand g22353(.dina(n17329), .dinb(n5536), .dout(n22493));
  jor  g22354(.dina(n22493), .dinb(n22492), .dout(n22494));
  jor  g22355(.dina(n22494), .dinb(n22491), .dout(n22495));
  jor  g22356(.dina(n22495), .dinb(n22490), .dout(n22496));
  jxor g22357(.dina(n22496), .dinb(n5277), .dout(n22497));
  jor  g22358(.dina(n22497), .dinb(n22489), .dout(n22498));
  jxor g22359(.dina(n21645), .dinb(n21644), .dout(n22499));
  jnot g22360(.din(n22499), .dout(n22500));
  jand g22361(.dina(n17537), .dinb(n5280), .dout(n22501));
  jand g22362(.dina(n17329), .dinb(n5531), .dout(n22502));
  jand g22363(.dina(n17535), .dinb(n5814), .dout(n22503));
  jor  g22364(.dina(n22503), .dinb(n22502), .dout(n22504));
  jand g22365(.dina(n17330), .dinb(n5536), .dout(n22505));
  jor  g22366(.dina(n22505), .dinb(n22504), .dout(n22506));
  jor  g22367(.dina(n22506), .dinb(n22501), .dout(n22507));
  jxor g22368(.dina(n22507), .dinb(n5277), .dout(n22508));
  jor  g22369(.dina(n22508), .dinb(n22500), .dout(n22509));
  jxor g22370(.dina(n21640), .dinb(n21639), .dout(n22510));
  jnot g22371(.din(n22510), .dout(n22511));
  jand g22372(.dina(n17549), .dinb(n5280), .dout(n22512));
  jand g22373(.dina(n17329), .dinb(n5814), .dout(n22513));
  jand g22374(.dina(n17330), .dinb(n5531), .dout(n22514));
  jand g22375(.dina(n16940), .dinb(n5536), .dout(n22515));
  jor  g22376(.dina(n22515), .dinb(n22514), .dout(n22516));
  jor  g22377(.dina(n22516), .dinb(n22513), .dout(n22517));
  jor  g22378(.dina(n22517), .dinb(n22512), .dout(n22518));
  jxor g22379(.dina(n22518), .dinb(n5277), .dout(n22519));
  jor  g22380(.dina(n22519), .dinb(n22511), .dout(n22520));
  jxor g22381(.dina(n21637), .dinb(n21636), .dout(n22521));
  jnot g22382(.din(n22521), .dout(n22522));
  jand g22383(.dina(n17561), .dinb(n5280), .dout(n22523));
  jand g22384(.dina(n17330), .dinb(n5814), .dout(n22524));
  jand g22385(.dina(n16940), .dinb(n5531), .dout(n22525));
  jand g22386(.dina(n16604), .dinb(n5536), .dout(n22526));
  jor  g22387(.dina(n22526), .dinb(n22525), .dout(n22527));
  jor  g22388(.dina(n22527), .dinb(n22524), .dout(n22528));
  jor  g22389(.dina(n22528), .dinb(n22523), .dout(n22529));
  jxor g22390(.dina(n22529), .dinb(n5277), .dout(n22530));
  jor  g22391(.dina(n22530), .dinb(n22522), .dout(n22531));
  jxor g22392(.dina(n21632), .dinb(n21631), .dout(n22532));
  jnot g22393(.din(n22532), .dout(n22533));
  jand g22394(.dina(n16942), .dinb(n5280), .dout(n22534));
  jand g22395(.dina(n16940), .dinb(n5814), .dout(n22535));
  jand g22396(.dina(n16604), .dinb(n5531), .dout(n22536));
  jand g22397(.dina(n16355), .dinb(n5536), .dout(n22537));
  jor  g22398(.dina(n22537), .dinb(n22536), .dout(n22538));
  jor  g22399(.dina(n22538), .dinb(n22535), .dout(n22539));
  jor  g22400(.dina(n22539), .dinb(n22534), .dout(n22540));
  jxor g22401(.dina(n22540), .dinb(n5277), .dout(n22541));
  jor  g22402(.dina(n22541), .dinb(n22533), .dout(n22542));
  jxor g22403(.dina(n21628), .dinb(n21620), .dout(n22543));
  jnot g22404(.din(n22543), .dout(n22544));
  jand g22405(.dina(n16606), .dinb(n5280), .dout(n22545));
  jand g22406(.dina(n16355), .dinb(n5531), .dout(n22546));
  jand g22407(.dina(n16604), .dinb(n5814), .dout(n22547));
  jor  g22408(.dina(n22547), .dinb(n22546), .dout(n22548));
  jand g22409(.dina(n16360), .dinb(n5536), .dout(n22549));
  jor  g22410(.dina(n22549), .dinb(n22548), .dout(n22550));
  jor  g22411(.dina(n22550), .dinb(n22545), .dout(n22551));
  jxor g22412(.dina(n22551), .dinb(n5277), .dout(n22552));
  jor  g22413(.dina(n22552), .dinb(n22544), .dout(n22553));
  jand g22414(.dina(n16616), .dinb(n5280), .dout(n22554));
  jand g22415(.dina(n16355), .dinb(n5814), .dout(n22555));
  jand g22416(.dina(n16360), .dinb(n5531), .dout(n22556));
  jand g22417(.dina(n15841), .dinb(n5536), .dout(n22557));
  jor  g22418(.dina(n22557), .dinb(n22556), .dout(n22558));
  jor  g22419(.dina(n22558), .dinb(n22555), .dout(n22559));
  jor  g22420(.dina(n22559), .dinb(n22554), .dout(n22560));
  jxor g22421(.dina(n22560), .dinb(n5277), .dout(n22561));
  jnot g22422(.din(n22561), .dout(n22562));
  jor  g22423(.dina(n21607), .dinb(n4713), .dout(n22563));
  jxor g22424(.dina(n22563), .dinb(n21615), .dout(n22564));
  jand g22425(.dina(n22564), .dinb(n22562), .dout(n22565));
  jand g22426(.dina(n21604), .dinb(\a[8] ), .dout(n22566));
  jxor g22427(.dina(n22566), .dinb(n21602), .dout(n22567));
  jnot g22428(.din(n22567), .dout(n22568));
  jand g22429(.dina(n16632), .dinb(n5280), .dout(n22569));
  jand g22430(.dina(n15841), .dinb(n5531), .dout(n22570));
  jand g22431(.dina(n16360), .dinb(n5814), .dout(n22571));
  jor  g22432(.dina(n22571), .dinb(n22570), .dout(n22572));
  jand g22433(.dina(n15579), .dinb(n5536), .dout(n22573));
  jor  g22434(.dina(n22573), .dinb(n22572), .dout(n22574));
  jor  g22435(.dina(n22574), .dinb(n22569), .dout(n22575));
  jxor g22436(.dina(n22575), .dinb(n5277), .dout(n22576));
  jor  g22437(.dina(n22576), .dinb(n22568), .dout(n22577));
  jand g22438(.dina(n15329), .dinb(n5280), .dout(n22578));
  jand g22439(.dina(n15020), .dinb(n5531), .dout(n22579));
  jand g22440(.dina(n15327), .dinb(n5814), .dout(n22580));
  jor  g22441(.dina(n22580), .dinb(n22579), .dout(n22581));
  jor  g22442(.dina(n22581), .dinb(n22578), .dout(n22582));
  jnot g22443(.din(n22582), .dout(n22583));
  jand g22444(.dina(n15020), .dinb(n5279), .dout(n22584));
  jnot g22445(.din(n22584), .dout(n22585));
  jand g22446(.dina(n22585), .dinb(\a[5] ), .dout(n22586));
  jand g22447(.dina(n22586), .dinb(n22583), .dout(n22587));
  jand g22448(.dina(n15580), .dinb(n5280), .dout(n22588));
  jand g22449(.dina(n15327), .dinb(n5531), .dout(n22589));
  jand g22450(.dina(n15579), .dinb(n5814), .dout(n22590));
  jor  g22451(.dina(n22590), .dinb(n22589), .dout(n22591));
  jand g22452(.dina(n15020), .dinb(n5536), .dout(n22592));
  jor  g22453(.dina(n22592), .dinb(n22591), .dout(n22593));
  jor  g22454(.dina(n22593), .dinb(n22588), .dout(n22594));
  jnot g22455(.din(n22594), .dout(n22595));
  jand g22456(.dina(n22595), .dinb(n22587), .dout(n22596));
  jand g22457(.dina(n22596), .dinb(n21604), .dout(n22597));
  jnot g22458(.din(n22597), .dout(n22598));
  jxor g22459(.dina(n22596), .dinb(n21604), .dout(n22599));
  jnot g22460(.din(n22599), .dout(n22600));
  jand g22461(.dina(n15848), .dinb(n5280), .dout(n22601));
  jand g22462(.dina(n15579), .dinb(n5531), .dout(n22602));
  jand g22463(.dina(n15841), .dinb(n5814), .dout(n22603));
  jor  g22464(.dina(n22603), .dinb(n22602), .dout(n22604));
  jand g22465(.dina(n15327), .dinb(n5536), .dout(n22605));
  jor  g22466(.dina(n22605), .dinb(n22604), .dout(n22606));
  jor  g22467(.dina(n22606), .dinb(n22601), .dout(n22607));
  jxor g22468(.dina(n22607), .dinb(n5277), .dout(n22608));
  jor  g22469(.dina(n22608), .dinb(n22600), .dout(n22609));
  jand g22470(.dina(n22609), .dinb(n22598), .dout(n22610));
  jnot g22471(.din(n22610), .dout(n22611));
  jxor g22472(.dina(n22576), .dinb(n22568), .dout(n22612));
  jand g22473(.dina(n22612), .dinb(n22611), .dout(n22613));
  jnot g22474(.din(n22613), .dout(n22614));
  jand g22475(.dina(n22614), .dinb(n22577), .dout(n22615));
  jnot g22476(.din(n22615), .dout(n22616));
  jxor g22477(.dina(n22564), .dinb(n22562), .dout(n22617));
  jand g22478(.dina(n22617), .dinb(n22616), .dout(n22618));
  jor  g22479(.dina(n22618), .dinb(n22565), .dout(n22619));
  jxor g22480(.dina(n22552), .dinb(n22544), .dout(n22620));
  jand g22481(.dina(n22620), .dinb(n22619), .dout(n22621));
  jnot g22482(.din(n22621), .dout(n22622));
  jand g22483(.dina(n22622), .dinb(n22553), .dout(n22623));
  jnot g22484(.din(n22623), .dout(n22624));
  jxor g22485(.dina(n22541), .dinb(n22533), .dout(n22625));
  jand g22486(.dina(n22625), .dinb(n22624), .dout(n22626));
  jnot g22487(.din(n22626), .dout(n22627));
  jand g22488(.dina(n22627), .dinb(n22542), .dout(n22628));
  jnot g22489(.din(n22628), .dout(n22629));
  jxor g22490(.dina(n22530), .dinb(n22522), .dout(n22630));
  jand g22491(.dina(n22630), .dinb(n22629), .dout(n22631));
  jnot g22492(.din(n22631), .dout(n22632));
  jand g22493(.dina(n22632), .dinb(n22531), .dout(n22633));
  jnot g22494(.din(n22633), .dout(n22634));
  jxor g22495(.dina(n22519), .dinb(n22511), .dout(n22635));
  jand g22496(.dina(n22635), .dinb(n22634), .dout(n22636));
  jnot g22497(.din(n22636), .dout(n22637));
  jand g22498(.dina(n22637), .dinb(n22520), .dout(n22638));
  jnot g22499(.din(n22638), .dout(n22639));
  jxor g22500(.dina(n22508), .dinb(n22500), .dout(n22640));
  jand g22501(.dina(n22640), .dinb(n22639), .dout(n22641));
  jnot g22502(.din(n22641), .dout(n22642));
  jand g22503(.dina(n22642), .dinb(n22509), .dout(n22643));
  jnot g22504(.din(n22643), .dout(n22644));
  jxor g22505(.dina(n22497), .dinb(n22489), .dout(n22645));
  jand g22506(.dina(n22645), .dinb(n22644), .dout(n22646));
  jnot g22507(.din(n22646), .dout(n22647));
  jand g22508(.dina(n22647), .dinb(n22498), .dout(n22648));
  jnot g22509(.din(n22648), .dout(n22649));
  jxor g22510(.dina(n22485), .dinb(n22477), .dout(n22650));
  jand g22511(.dina(n22650), .dinb(n22649), .dout(n22651));
  jor  g22512(.dina(n22651), .dinb(n22487), .dout(n22652));
  jxor g22513(.dina(n22473), .dinb(n22465), .dout(n22653));
  jand g22514(.dina(n22653), .dinb(n22652), .dout(n22654));
  jor  g22515(.dina(n22654), .dinb(n22475), .dout(n22655));
  jxor g22516(.dina(n22461), .dinb(n22453), .dout(n22656));
  jand g22517(.dina(n22656), .dinb(n22655), .dout(n22657));
  jor  g22518(.dina(n22657), .dinb(n22463), .dout(n22658));
  jxor g22519(.dina(n22449), .dinb(n22441), .dout(n22659));
  jand g22520(.dina(n22659), .dinb(n22658), .dout(n22660));
  jor  g22521(.dina(n22660), .dinb(n22451), .dout(n22661));
  jxor g22522(.dina(n22437), .dinb(n22429), .dout(n22662));
  jand g22523(.dina(n22662), .dinb(n22661), .dout(n22663));
  jor  g22524(.dina(n22663), .dinb(n22439), .dout(n22664));
  jxor g22525(.dina(n22425), .dinb(n22417), .dout(n22665));
  jand g22526(.dina(n22665), .dinb(n22664), .dout(n22666));
  jor  g22527(.dina(n22666), .dinb(n22427), .dout(n22667));
  jxor g22528(.dina(n22414), .dinb(n22406), .dout(n22668));
  jand g22529(.dina(n22668), .dinb(n22667), .dout(n22669));
  jor  g22530(.dina(n22669), .dinb(n22415), .dout(n22670));
  jxor g22531(.dina(n22403), .dinb(n22395), .dout(n22671));
  jand g22532(.dina(n22671), .dinb(n22670), .dout(n22672));
  jor  g22533(.dina(n22672), .dinb(n22405), .dout(n22673));
  jxor g22534(.dina(n22391), .dinb(n22383), .dout(n22674));
  jand g22535(.dina(n22674), .dinb(n22673), .dout(n22675));
  jor  g22536(.dina(n22675), .dinb(n22393), .dout(n22676));
  jxor g22537(.dina(n22379), .dinb(n22371), .dout(n22677));
  jand g22538(.dina(n22677), .dinb(n22676), .dout(n22678));
  jor  g22539(.dina(n22678), .dinb(n22381), .dout(n22679));
  jxor g22540(.dina(n22368), .dinb(n22360), .dout(n22680));
  jand g22541(.dina(n22680), .dinb(n22679), .dout(n22681));
  jor  g22542(.dina(n22681), .dinb(n22370), .dout(n22682));
  jxor g22543(.dina(n22356), .dinb(n22348), .dout(n22683));
  jand g22544(.dina(n22683), .dinb(n22682), .dout(n22684));
  jor  g22545(.dina(n22684), .dinb(n22358), .dout(n22685));
  jxor g22546(.dina(n22344), .dinb(n22336), .dout(n22686));
  jand g22547(.dina(n22686), .dinb(n22685), .dout(n22687));
  jor  g22548(.dina(n22687), .dinb(n22346), .dout(n22688));
  jxor g22549(.dina(n22332), .dinb(n22324), .dout(n22689));
  jand g22550(.dina(n22689), .dinb(n22688), .dout(n22690));
  jor  g22551(.dina(n22690), .dinb(n22334), .dout(n22691));
  jnot g22552(.din(n22691), .dout(n22692));
  jxor g22553(.dina(n22322), .dinb(n22313), .dout(n22693));
  jor  g22554(.dina(n22693), .dinb(n22692), .dout(n22694));
  jand g22555(.dina(n22694), .dinb(n22323), .dout(n22695));
  jxor g22556(.dina(n22311), .dinb(n22302), .dout(n22696));
  jor  g22557(.dina(n22696), .dinb(n22695), .dout(n22697));
  jand g22558(.dina(n22697), .dinb(n22312), .dout(n22698));
  jxor g22559(.dina(n22299), .dinb(n22290), .dout(n22699));
  jnot g22560(.din(n22699), .dout(n22700));
  jor  g22561(.dina(n22700), .dinb(n22698), .dout(n22701));
  jand g22562(.dina(n22701), .dinb(n22301), .dout(n22702));
  jxor g22563(.dina(n22287), .dinb(n22277), .dout(n22703));
  jor  g22564(.dina(n22703), .dinb(n22702), .dout(n22704));
  jand g22565(.dina(n22704), .dinb(n22289), .dout(n22705));
  jxor g22566(.dina(n22275), .dinb(n21987), .dout(n22706));
  jor  g22567(.dina(n22706), .dinb(n22705), .dout(n22707));
  jand g22568(.dina(n22707), .dinb(n22276), .dout(n22708));
  jnot g22569(.din(n21869), .dout(n22709));
  jor  g22570(.dina(n21984), .dinb(n22709), .dout(n22710));
  jnot g22571(.din(n22710), .dout(n22711));
  jand g22572(.dina(n21986), .dinb(n21724), .dout(n22712));
  jor  g22573(.dina(n22712), .dinb(n22711), .dout(n22713));
  jnot g22574(.din(n21858), .dout(n22714));
  jor  g22575(.dina(n21866), .dinb(n22714), .dout(n22715));
  jnot g22576(.din(n22715), .dout(n22716));
  jand g22577(.dina(n21868), .dinb(n21730), .dout(n22717));
  jor  g22578(.dina(n22717), .dinb(n22716), .dout(n22718));
  jor  g22579(.dina(n21856), .dinb(n21848), .dout(n22719));
  jnot g22580(.din(n22719), .dout(n22720));
  jand g22581(.dina(n21857), .dinb(n21734), .dout(n22721));
  jor  g22582(.dina(n22721), .dinb(n22720), .dout(n22722));
  jor  g22583(.dina(n21845), .dinb(n21837), .dout(n22723));
  jand g22584(.dina(n21846), .dinb(n21739), .dout(n22724));
  jnot g22585(.din(n22724), .dout(n22725));
  jand g22586(.dina(n22725), .dinb(n22723), .dout(n22726));
  jnot g22587(.din(n22726), .dout(n22727));
  jor  g22588(.dina(n21834), .dinb(n21826), .dout(n22728));
  jand g22589(.dina(n21835), .dinb(n21744), .dout(n22729));
  jnot g22590(.din(n22729), .dout(n22730));
  jand g22591(.dina(n22730), .dinb(n22728), .dout(n22731));
  jnot g22592(.din(n22731), .dout(n22732));
  jor  g22593(.dina(n21823), .dinb(n21815), .dout(n22733));
  jand g22594(.dina(n21824), .dinb(n21749), .dout(n22734));
  jnot g22595(.din(n22734), .dout(n22735));
  jand g22596(.dina(n22735), .dinb(n22733), .dout(n22736));
  jnot g22597(.din(n22736), .dout(n22737));
  jor  g22598(.dina(n21812), .dinb(n21804), .dout(n22738));
  jand g22599(.dina(n21813), .dinb(n21754), .dout(n22739));
  jnot g22600(.din(n22739), .dout(n22740));
  jand g22601(.dina(n22740), .dinb(n22738), .dout(n22741));
  jnot g22602(.din(n22741), .dout(n22742));
  jor  g22603(.dina(n21801), .dinb(n21793), .dout(n22743));
  jand g22604(.dina(n21802), .dinb(n21759), .dout(n22744));
  jnot g22605(.din(n22744), .dout(n22745));
  jand g22606(.dina(n22745), .dinb(n22743), .dout(n22746));
  jnot g22607(.din(n22746), .dout(n22747));
  jand g22608(.dina(n21790), .dinb(n21783), .dout(n22748));
  jand g22609(.dina(n21791), .dinb(n21764), .dout(n22749));
  jor  g22610(.dina(n22749), .dinb(n22748), .dout(n22750));
  jand g22611(.dina(n7512), .dinb(n4678), .dout(n22751));
  jand g22612(.dina(n22751), .dinb(n21268), .dout(n22752));
  jand g22613(.dina(n22752), .dinb(n3238), .dout(n22753));
  jand g22614(.dina(n901), .dinb(n871), .dout(n22754));
  jand g22615(.dina(n22754), .dinb(n1366), .dout(n22755));
  jand g22616(.dina(n895), .dinb(n472), .dout(n22756));
  jand g22617(.dina(n22756), .dinb(n1324), .dout(n22757));
  jand g22618(.dina(n22757), .dinb(n22755), .dout(n22758));
  jand g22619(.dina(n9763), .dinb(n329), .dout(n22759));
  jand g22620(.dina(n22759), .dinb(n22758), .dout(n22760));
  jand g22621(.dina(n22760), .dinb(n21248), .dout(n22761));
  jand g22622(.dina(n22761), .dinb(n22753), .dout(n22762));
  jand g22623(.dina(n22762), .dinb(n22227), .dout(n22763));
  jand g22624(.dina(n22763), .dinb(n15927), .dout(n22764));
  jnot g22625(.din(n22764), .dout(n22765));
  jand g22626(.dina(n16632), .dinb(n5076), .dout(n22766));
  jand g22627(.dina(n16360), .dinb(n5084), .dout(n22767));
  jand g22628(.dina(n15841), .dinb(n5082), .dout(n22768));
  jand g22629(.dina(n15579), .dinb(n6050), .dout(n22769));
  jor  g22630(.dina(n22769), .dinb(n22768), .dout(n22770));
  jor  g22631(.dina(n22770), .dinb(n22767), .dout(n22771));
  jor  g22632(.dina(n22771), .dinb(n22766), .dout(n22772));
  jxor g22633(.dina(n22772), .dinb(n22765), .dout(n22773));
  jxor g22634(.dina(n22773), .dinb(n22750), .dout(n22774));
  jnot g22635(.din(n22774), .dout(n22775));
  jand g22636(.dina(n16942), .dinb(n2936), .dout(n22776));
  jand g22637(.dina(n16940), .dinb(n2943), .dout(n22777));
  jand g22638(.dina(n16604), .dinb(n2940), .dout(n22778));
  jand g22639(.dina(n16355), .dinb(n3684), .dout(n22779));
  jor  g22640(.dina(n22779), .dinb(n22778), .dout(n22780));
  jor  g22641(.dina(n22780), .dinb(n22777), .dout(n22781));
  jor  g22642(.dina(n22781), .dinb(n22776), .dout(n22782));
  jxor g22643(.dina(n22782), .dinb(n93), .dout(n22783));
  jxor g22644(.dina(n22783), .dinb(n22775), .dout(n22784));
  jxor g22645(.dina(n22784), .dinb(n22747), .dout(n22785));
  jnot g22646(.din(n22785), .dout(n22786));
  jand g22647(.dina(n17537), .dinb(n71), .dout(n22787));
  jand g22648(.dina(n17535), .dinb(n796), .dout(n22788));
  jand g22649(.dina(n17329), .dinb(n731), .dout(n22789));
  jand g22650(.dina(n17330), .dinb(n1806), .dout(n22790));
  jor  g22651(.dina(n22790), .dinb(n22789), .dout(n22791));
  jor  g22652(.dina(n22791), .dinb(n22788), .dout(n22792));
  jor  g22653(.dina(n22792), .dinb(n22787), .dout(n22793));
  jxor g22654(.dina(n22793), .dinb(n77), .dout(n22794));
  jxor g22655(.dina(n22794), .dinb(n22786), .dout(n22795));
  jxor g22656(.dina(n22795), .dinb(n22742), .dout(n22796));
  jand g22657(.dina(n18502), .dinb(n806), .dout(n22797));
  jand g22658(.dina(n18292), .dinb(n1620), .dout(n22798));
  jand g22659(.dina(n18293), .dinb(n1612), .dout(n22799));
  jand g22660(.dina(n17942), .dinb(n1644), .dout(n22800));
  jor  g22661(.dina(n22800), .dinb(n22799), .dout(n22801));
  jor  g22662(.dina(n22801), .dinb(n22798), .dout(n22802));
  jor  g22663(.dina(n22802), .dinb(n22797), .dout(n22803));
  jxor g22664(.dina(n22803), .dinb(\a[23] ), .dout(n22804));
  jxor g22665(.dina(n22804), .dinb(n22796), .dout(n22805));
  jxor g22666(.dina(n22805), .dinb(n22737), .dout(n22806));
  jnot g22667(.din(n22806), .dout(n22807));
  jand g22668(.dina(n19399), .dinb(n1819), .dout(n22808));
  jand g22669(.dina(n19220), .dinb(n2243), .dout(n22809));
  jand g22670(.dina(n18914), .dinb(n2180), .dout(n22810));
  jand g22671(.dina(n18488), .dinb(n2185), .dout(n22811));
  jor  g22672(.dina(n22811), .dinb(n22810), .dout(n22812));
  jor  g22673(.dina(n22812), .dinb(n22809), .dout(n22813));
  jor  g22674(.dina(n22813), .dinb(n22808), .dout(n22814));
  jxor g22675(.dina(n22814), .dinb(n2196), .dout(n22815));
  jxor g22676(.dina(n22815), .dinb(n22807), .dout(n22816));
  jxor g22677(.dina(n22816), .dinb(n22732), .dout(n22817));
  jand g22678(.dina(n19924), .dinb(n2743), .dout(n22818));
  jand g22679(.dina(n19922), .dinb(n2752), .dout(n22819));
  jand g22680(.dina(n19373), .dinb(n2748), .dout(n22820));
  jand g22681(.dina(n19219), .dinb(n2757), .dout(n22821));
  jor  g22682(.dina(n22821), .dinb(n22820), .dout(n22822));
  jor  g22683(.dina(n22822), .dinb(n22819), .dout(n22823));
  jor  g22684(.dina(n22823), .dinb(n22818), .dout(n22824));
  jxor g22685(.dina(n22824), .dinb(\a[17] ), .dout(n22825));
  jxor g22686(.dina(n22825), .dinb(n22817), .dout(n22826));
  jxor g22687(.dina(n22826), .dinb(n22727), .dout(n22827));
  jnot g22688(.din(n22827), .dout(n22828));
  jand g22689(.dina(n20346), .dinb(n3423), .dout(n22829));
  jand g22690(.dina(n20204), .dinb(n3428), .dout(n22830));
  jand g22691(.dina(n20344), .dinb(n3569), .dout(n22831));
  jor  g22692(.dina(n22831), .dinb(n22830), .dout(n22832));
  jand g22693(.dina(n20205), .dinb(n3210), .dout(n22833));
  jor  g22694(.dina(n22833), .dinb(n22832), .dout(n22834));
  jor  g22695(.dina(n22834), .dinb(n22829), .dout(n22835));
  jxor g22696(.dina(n22835), .dinb(n3473), .dout(n22836));
  jxor g22697(.dina(n22836), .dinb(n22828), .dout(n22837));
  jxor g22698(.dina(n22837), .dinb(n22722), .dout(n22838));
  jand g22699(.dina(n21355), .dinb(n4022), .dout(n22839));
  jand g22700(.dina(n21198), .dinb(n4027), .dout(n22840));
  jand g22701(.dina(n21197), .dinb(n4220), .dout(n22841));
  jor  g22702(.dina(n22841), .dinb(n22840), .dout(n22842));
  jand g22703(.dina(n20947), .dinb(n3870), .dout(n22843));
  jor  g22704(.dina(n22843), .dinb(n22842), .dout(n22844));
  jor  g22705(.dina(n22844), .dinb(n22839), .dout(n22845));
  jxor g22706(.dina(n22845), .dinb(n4050), .dout(n22846));
  jxor g22707(.dina(n22846), .dinb(n22838), .dout(n22847));
  jnot g22708(.din(n22847), .dout(n22848));
  jxor g22709(.dina(n22848), .dinb(n22718), .dout(n22849));
  jand g22710(.dina(n22291), .dinb(n4691), .dout(n22850));
  jand g22711(.dina(n22164), .dinb(n4941), .dout(n22851));
  jand g22712(.dina(n21974), .dinb(n4696), .dout(n22852));
  jand g22713(.dina(n21340), .dinb(n4701), .dout(n22853));
  jor  g22714(.dina(n22853), .dinb(n22852), .dout(n22854));
  jor  g22715(.dina(n22854), .dinb(n22851), .dout(n22855));
  jor  g22716(.dina(n22855), .dinb(n22850), .dout(n22856));
  jxor g22717(.dina(n22856), .dinb(n4713), .dout(n22857));
  jxor g22718(.dina(n22857), .dinb(n22849), .dout(n22858));
  jnot g22719(.din(n22858), .dout(n22859));
  jxor g22720(.dina(n22859), .dinb(n22713), .dout(n22860));
  jand g22721(.dina(n22265), .dinb(n22163), .dout(n22861));
  jand g22722(.dina(n22266), .dinb(n22175), .dout(n22862));
  jor  g22723(.dina(n22862), .dinb(n22861), .dout(n22863));
  jand g22724(.dina(n22258), .dinb(n22180), .dout(n22864));
  jnot g22725(.din(n22864), .dout(n22865));
  jor  g22726(.dina(n22264), .dinb(n22260), .dout(n22866));
  jand g22727(.dina(n22866), .dinb(n22865), .dout(n22867));
  jor  g22728(.dina(n22912), .dinb(n22184), .dout(n22868));
  jand g22729(.dina(n22257), .dinb(n22192), .dout(n22869));
  jnot g22730(.din(n22869), .dout(n22870));
  jand g22731(.dina(n22870), .dinb(n22868), .dout(n22871));
  jnot g22732(.din(n22871), .dout(n22872));
  jand g22733(.dina(n22246), .dinb(n22197), .dout(n22873));
  jnot g22734(.din(n22873), .dout(n22874));
  jor  g22735(.dina(n22256), .dinb(n22248), .dout(n22875));
  jand g22736(.dina(n22875), .dinb(n22874), .dout(n22876));
  jand g22737(.dina(n16930), .dinb(n71), .dout(n22877));
  jand g22738(.dina(n16592), .dinb(n731), .dout(n22878));
  jand g22739(.dina(n16928), .dinb(n796), .dout(n22879));
  jor  g22740(.dina(n22879), .dinb(n22878), .dout(n22880));
  jand g22741(.dina(n16343), .dinb(n1806), .dout(n22881));
  jor  g22742(.dina(n22881), .dinb(n22880), .dout(n22882));
  jor  g22743(.dina(n22882), .dinb(n22877), .dout(n22883));
  jxor g22744(.dina(n22883), .dinb(n77), .dout(n22884));
  jxor g22745(.dina(n22884), .dinb(n22876), .dout(n22885));
  jand g22746(.dina(n22235), .dinb(n22204), .dout(n22886));
  jnot g22747(.din(n22886), .dout(n22887));
  jor  g22748(.dina(n22245), .dinb(n22237), .dout(n22888));
  jand g22749(.dina(n22888), .dinb(n22887), .dout(n22889));
  jnot g22750(.din(n22889), .dout(n22890));
  jand g22751(.dina(n22233), .dinb(n22114), .dout(n22891));
  jand g22752(.dina(n22234), .dinb(n22209), .dout(n22892));
  jor  g22753(.dina(n22892), .dinb(n22891), .dout(n22893));
  jand g22754(.dina(n15122), .dinb(n3762), .dout(n22894));
  jand g22755(.dina(n22894), .dinb(n6335), .dout(n22895));
  jand g22756(.dina(n22895), .dinb(n20849), .dout(n22896));
  jand g22757(.dina(n2385), .dinb(n1713), .dout(n22897));
  jand g22758(.dina(n2148), .dinb(n1449), .dout(n22898));
  jand g22759(.dina(n22898), .dinb(n511), .dout(n22899));
  jand g22760(.dina(n22899), .dinb(n22897), .dout(n22900));
  jand g22761(.dina(n22900), .dinb(n7498), .dout(n22901));
  jand g22762(.dina(n8106), .dinb(n6231), .dout(n22902));
  jand g22763(.dina(n22902), .dinb(n22901), .dout(n22903));
  jand g22764(.dina(n22903), .dinb(n11418), .dout(n22904));
  jand g22765(.dina(n18385), .dinb(n13313), .dout(n22905));
  jand g22766(.dina(n22905), .dinb(n22904), .dout(n22906));
  jand g22767(.dina(n22906), .dinb(n839), .dout(n22907));
  jand g22768(.dina(n22907), .dinb(n22896), .dout(n22908));
  jxor g22769(.dina(n22908), .dinb(n22233), .dout(n22909));
  jor  g22770(.dina(n1616), .dinb(n805), .dout(n22910));
  jand g22771(.dina(n22910), .dinb(n16924), .dout(n22911));
  jxor g22772(.dina(n22911), .dinb(n65), .dout(n22912));
  jxor g22773(.dina(n22912), .dinb(n22909), .dout(n22913));
  jxor g22774(.dina(n22913), .dinb(n22893), .dout(n22914));
  jand g22775(.dina(n15317), .dinb(n5076), .dout(n22915));
  jand g22776(.dina(n15315), .dinb(n5084), .dout(n22916));
  jand g22777(.dina(n14549), .dinb(n5082), .dout(n22917));
  jand g22778(.dina(n14447), .dinb(n6050), .dout(n22918));
  jor  g22779(.dina(n22918), .dinb(n22917), .dout(n22919));
  jor  g22780(.dina(n22919), .dinb(n22916), .dout(n22920));
  jor  g22781(.dina(n22920), .dinb(n22915), .dout(n22921));
  jxor g22782(.dina(n22921), .dinb(n22914), .dout(n22922));
  jxor g22783(.dina(n22922), .dinb(n22890), .dout(n22923));
  jnot g22784(.din(n22923), .dout(n22924));
  jand g22785(.dina(n16084), .dinb(n2936), .dout(n22925));
  jand g22786(.dina(n16082), .dinb(n2943), .dout(n22926));
  jand g22787(.dina(n15829), .dinb(n2940), .dout(n22927));
  jand g22788(.dina(n15567), .dinb(n3684), .dout(n22928));
  jor  g22789(.dina(n22928), .dinb(n22927), .dout(n22929));
  jor  g22790(.dina(n22929), .dinb(n22926), .dout(n22930));
  jor  g22791(.dina(n22930), .dinb(n22925), .dout(n22931));
  jxor g22792(.dina(n22931), .dinb(n93), .dout(n22932));
  jxor g22793(.dina(n22932), .dinb(n22924), .dout(n22933));
  jxor g22794(.dina(n22933), .dinb(n22885), .dout(n22934));
  jxor g22795(.dina(n22934), .dinb(n22872), .dout(n22935));
  jnot g22796(.din(n22935), .dout(n22936));
  jxor g22797(.dina(n22936), .dinb(n22867), .dout(n22937));
  jxor g22798(.dina(n22937), .dinb(n22265), .dout(n22938));
  jxor g22799(.dina(n22938), .dinb(n22863), .dout(n22939));
  jand g22800(.dina(n22939), .dinb(n5280), .dout(n22940));
  jand g22801(.dina(n22937), .dinb(n5814), .dout(n22941));
  jand g22802(.dina(n22265), .dinb(n5531), .dout(n22942));
  jand g22803(.dina(n22163), .dinb(n5536), .dout(n22943));
  jor  g22804(.dina(n22943), .dinb(n22942), .dout(n22944));
  jor  g22805(.dina(n22944), .dinb(n22941), .dout(n22945));
  jor  g22806(.dina(n22945), .dinb(n22940), .dout(n22946));
  jxor g22807(.dina(n22946), .dinb(n5277), .dout(n22947));
  jxor g22808(.dina(n22947), .dinb(n22860), .dout(n22948));
  jnot g22809(.din(n22948), .dout(n22949));
  jxor g22810(.dina(n22949), .dinb(n22708), .dout(n22950));
  jor  g22811(.dina(n22884), .dinb(n22876), .dout(n22951));
  jand g22812(.dina(n22933), .dinb(n22885), .dout(n22952));
  jnot g22813(.din(n22952), .dout(n22953));
  jand g22814(.dina(n22953), .dinb(n22951), .dout(n22954));
  jnot g22815(.din(n22954), .dout(n22955));
  jand g22816(.dina(n22922), .dinb(n22890), .dout(n22956));
  jnot g22817(.din(n22956), .dout(n22957));
  jor  g22818(.dina(n22932), .dinb(n22924), .dout(n22958));
  jand g22819(.dina(n22958), .dinb(n22957), .dout(n22959));
  jnot g22820(.din(n22959), .dout(n22960));
  jand g22821(.dina(n22913), .dinb(n22893), .dout(n22961));
  jand g22822(.dina(n22921), .dinb(n22914), .dout(n22962));
  jor  g22823(.dina(n22962), .dinb(n22961), .dout(n22963));
  jor  g22824(.dina(n22908), .dinb(n22233), .dout(n22964));
  jand g22825(.dina(n22912), .dinb(n22909), .dout(n22965));
  jnot g22826(.din(n22965), .dout(n22966));
  jand g22827(.dina(n22966), .dinb(n22964), .dout(n22967));
  jand g22828(.dina(n7085), .dinb(n716), .dout(n22968));
  jand g22829(.dina(n7289), .dinb(n839), .dout(n22969));
  jand g22830(.dina(n22969), .dinb(n6440), .dout(n22970));
  jand g22831(.dina(n22970), .dinb(n884), .dout(n22971));
  jand g22832(.dina(n22971), .dinb(n22968), .dout(n22972));
  jand g22833(.dina(n22972), .dinb(n15536), .dout(n22973));
  jand g22834(.dina(n22973), .dinb(n3782), .dout(n22974));
  jand g22835(.dina(n3900), .dinb(n2716), .dout(n22975));
  jand g22836(.dina(n22975), .dinb(n3852), .dout(n22976));
  jand g22837(.dina(n22976), .dinb(n1370), .dout(n22977));
  jand g22838(.dina(n22977), .dinb(n6289), .dout(n22978));
  jand g22839(.dina(n22978), .dinb(n831), .dout(n22979));
  jand g22840(.dina(n22979), .dinb(n22974), .dout(n22980));
  jand g22841(.dina(n22980), .dinb(n6353), .dout(n22981));
  jnot g22842(.din(n22981), .dout(n22982));
  jxor g22843(.dina(n22982), .dinb(n22967), .dout(n22983));
  jand g22844(.dina(n15569), .dinb(n5076), .dout(n22984));
  jand g22845(.dina(n15567), .dinb(n5084), .dout(n22985));
  jand g22846(.dina(n14549), .dinb(n6050), .dout(n22986));
  jand g22847(.dina(n15315), .dinb(n5082), .dout(n22987));
  jor  g22848(.dina(n22987), .dinb(n22986), .dout(n22988));
  jor  g22849(.dina(n22988), .dinb(n22985), .dout(n22989));
  jor  g22850(.dina(n22989), .dinb(n22984), .dout(n22990));
  jxor g22851(.dina(n22990), .dinb(n22983), .dout(n22991));
  jxor g22852(.dina(n22991), .dinb(n22963), .dout(n22992));
  jnot g22853(.din(n22992), .dout(n22993));
  jand g22854(.dina(n16345), .dinb(n2936), .dout(n22994));
  jand g22855(.dina(n16082), .dinb(n2940), .dout(n22995));
  jand g22856(.dina(n16343), .dinb(n2943), .dout(n22996));
  jor  g22857(.dina(n22996), .dinb(n22995), .dout(n22997));
  jand g22858(.dina(n15829), .dinb(n3684), .dout(n22998));
  jor  g22859(.dina(n22998), .dinb(n22997), .dout(n22999));
  jor  g22860(.dina(n22999), .dinb(n22994), .dout(n23000));
  jxor g22861(.dina(n23000), .dinb(n93), .dout(n23001));
  jxor g22862(.dina(n23001), .dinb(n22993), .dout(n23002));
  jxor g22863(.dina(n23002), .dinb(n22960), .dout(n23003));
  jnot g22864(.din(n23003), .dout(n23004));
  jand g22865(.dina(n17312), .dinb(n71), .dout(n23005));
  jand g22866(.dina(n16928), .dinb(n731), .dout(n23006));
  jand g22867(.dina(n16592), .dinb(n1806), .dout(n23007));
  jand g22868(.dina(n16924), .dinb(n796), .dout(n23008));
  jor  g22869(.dina(n23008), .dinb(n23007), .dout(n23009));
  jor  g22870(.dina(n23009), .dinb(n23006), .dout(n23010));
  jor  g22871(.dina(n23010), .dinb(n23005), .dout(n23011));
  jxor g22872(.dina(n23011), .dinb(n77), .dout(n23012));
  jxor g22873(.dina(n23012), .dinb(n23004), .dout(n23013));
  jand g22874(.dina(n23013), .dinb(n22955), .dout(n23014));
  jnot g22875(.din(n23014), .dout(n23015));
  jand g22876(.dina(n22934), .dinb(n22872), .dout(n23016));
  jnot g22877(.din(n23016), .dout(n23017));
  jor  g22878(.dina(n22936), .dinb(n22867), .dout(n23018));
  jand g22879(.dina(n23018), .dinb(n23017), .dout(n23019));
  jxor g22880(.dina(n23013), .dinb(n22955), .dout(n23020));
  jnot g22881(.din(n23020), .dout(n23021));
  jor  g22882(.dina(n23021), .dinb(n23019), .dout(n23022));
  jand g22883(.dina(n23022), .dinb(n23015), .dout(n23023));
  jand g22884(.dina(n23002), .dinb(n22960), .dout(n23024));
  jnot g22885(.din(n23024), .dout(n23025));
  jor  g22886(.dina(n23012), .dinb(n23004), .dout(n23026));
  jand g22887(.dina(n23026), .dinb(n23025), .dout(n23027));
  jnot g22888(.din(n23027), .dout(n23028));
  jnot g22889(.din(n22967), .dout(n23029));
  jand g22890(.dina(n22981), .dinb(n23029), .dout(n23030));
  jand g22891(.dina(n22990), .dinb(n22983), .dout(n23031));
  jor  g22892(.dina(n23031), .dinb(n23030), .dout(n23032));
  jand g22893(.dina(n15831), .dinb(n5076), .dout(n23033));
  jand g22894(.dina(n15829), .dinb(n5084), .dout(n23034));
  jand g22895(.dina(n15567), .dinb(n5082), .dout(n23035));
  jand g22896(.dina(n15315), .dinb(n6050), .dout(n23036));
  jor  g22897(.dina(n23036), .dinb(n23035), .dout(n23037));
  jor  g22898(.dina(n23037), .dinb(n23034), .dout(n23038));
  jor  g22899(.dina(n23038), .dinb(n23033), .dout(n23039));
  jand g22900(.dina(n1560), .dinb(n1309), .dout(n23040));
  jand g22901(.dina(n23040), .dinb(n7292), .dout(n23041));
  jand g22902(.dina(n9768), .dinb(n542), .dout(n23042));
  jand g22903(.dina(n23042), .dinb(n1427), .dout(n23043));
  jand g22904(.dina(n23043), .dinb(n3170), .dout(n23044));
  jand g22905(.dina(n23044), .dinb(n23041), .dout(n23045));
  jand g22906(.dina(n5223), .dinb(n1189), .dout(n23046));
  jand g22907(.dina(n23046), .dinb(n15536), .dout(n23047));
  jand g22908(.dina(n23047), .dinb(n4449), .dout(n23048));
  jand g22909(.dina(n23048), .dinb(n23045), .dout(n23049));
  jand g22910(.dina(n23049), .dinb(n6268), .dout(n23050));
  jxor g22911(.dina(n23050), .dinb(n22982), .dout(n23051));
  jxor g22912(.dina(n23051), .dinb(n23039), .dout(n23052));
  jxor g22913(.dina(n23052), .dinb(n23032), .dout(n23053));
  jnot g22914(.din(n23053), .dout(n23054));
  jand g22915(.dina(n22991), .dinb(n22963), .dout(n23055));
  jnot g22916(.din(n23055), .dout(n23056));
  jor  g22917(.dina(n23001), .dinb(n22993), .dout(n23057));
  jand g22918(.dina(n23057), .dinb(n23056), .dout(n23058));
  jxor g22919(.dina(n23058), .dinb(n23054), .dout(n23059));
  jand g22920(.dina(n2309), .dinb(n2306), .dout(n23060));
  jand g22921(.dina(n16594), .dinb(n2936), .dout(n23067));
  jand g22922(.dina(n16343), .dinb(n2940), .dout(n23068));
  jand g22923(.dina(n16592), .dinb(n2943), .dout(n23069));
  jor  g22924(.dina(n23069), .dinb(n23068), .dout(n23070));
  jand g22925(.dina(n16082), .dinb(n3684), .dout(n23071));
  jor  g22926(.dina(n23071), .dinb(n23070), .dout(n23072));
  jor  g22927(.dina(n23072), .dinb(n23067), .dout(n23073));
  jxor g22928(.dina(n23073), .dinb(n93), .dout(n23074));
  jxor g22929(.dina(n23074), .dinb(n23115), .dout(n23075));
  jxor g22930(.dina(n23075), .dinb(n23059), .dout(n23076));
  jxor g22931(.dina(n23076), .dinb(n23028), .dout(n23077));
  jnot g22932(.din(n23077), .dout(n23078));
  jxor g22933(.dina(n23078), .dinb(n23023), .dout(n23079));
  jxor g22934(.dina(n23021), .dinb(n23019), .dout(n23080));
  jand g22935(.dina(n23080), .dinb(n23079), .dout(n23081));
  jand g22936(.dina(n23080), .dinb(n22937), .dout(n23082));
  jand g22937(.dina(n22937), .dinb(n22265), .dout(n23083));
  jand g22938(.dina(n22938), .dinb(n22863), .dout(n23084));
  jor  g22939(.dina(n23084), .dinb(n23083), .dout(n23085));
  jxor g22940(.dina(n23080), .dinb(n22937), .dout(n23086));
  jand g22941(.dina(n23086), .dinb(n23085), .dout(n23087));
  jor  g22942(.dina(n23087), .dinb(n23082), .dout(n23088));
  jxor g22943(.dina(n23080), .dinb(n23079), .dout(n23089));
  jand g22944(.dina(n23089), .dinb(n23088), .dout(n23090));
  jor  g22945(.dina(n23090), .dinb(n23081), .dout(n23091));
  jand g22946(.dina(n23076), .dinb(n23028), .dout(n23092));
  jnot g22947(.din(n23092), .dout(n23093));
  jor  g22948(.dina(n23078), .dinb(n23023), .dout(n23094));
  jand g22949(.dina(n23094), .dinb(n23093), .dout(n23095));
  jand g22950(.dina(n23052), .dinb(n23032), .dout(n23096));
  jnot g22951(.din(n23096), .dout(n23097));
  jor  g22952(.dina(n23058), .dinb(n23054), .dout(n23098));
  jand g22953(.dina(n23098), .dinb(n23097), .dout(n23099));
  jnot g22954(.din(n23099), .dout(n23100));
  jor  g22955(.dina(n23050), .dinb(n22982), .dout(n23101));
  jand g22956(.dina(n23051), .dinb(n23039), .dout(n23102));
  jnot g22957(.din(n23102), .dout(n23103));
  jand g22958(.dina(n23103), .dinb(n23101), .dout(n23104));
  jnot g22959(.din(n23104), .dout(n23105));
  jand g22960(.dina(n7975), .dinb(n7664), .dout(n23106));
  jand g22961(.dina(n583), .dinb(n843), .dout(n23107));
  jand g22962(.dina(n23107), .dinb(n23106), .dout(n23108));
  jand g22963(.dina(n7266), .dinb(n1291), .dout(n23109));
  jand g22964(.dina(n23109), .dinb(n7285), .dout(n23110));
  jand g22965(.dina(n23110), .dinb(n23108), .dout(n23111));
  jxor g22966(.dina(n23111), .dinb(n22981), .dout(n23112));
  jand g22967(.dina(n451), .dinb(n408), .dout(n23113));
  jand g22968(.dina(n23113), .dinb(n16924), .dout(n23114));
  jxor g22969(.dina(n23114), .dinb(n77), .dout(n23115));
  jxor g22970(.dina(n23115), .dinb(n23112), .dout(n23116));
  jxor g22971(.dina(n23116), .dinb(n23105), .dout(n23117));
  jand g22972(.dina(n16084), .dinb(n5076), .dout(n23118));
  jand g22973(.dina(n16082), .dinb(n5084), .dout(n23119));
  jand g22974(.dina(n15829), .dinb(n5082), .dout(n23120));
  jand g22975(.dina(n15567), .dinb(n6050), .dout(n23121));
  jor  g22976(.dina(n23121), .dinb(n23120), .dout(n23122));
  jor  g22977(.dina(n23122), .dinb(n23119), .dout(n23123));
  jor  g22978(.dina(n23123), .dinb(n23118), .dout(n23124));
  jxor g22979(.dina(n23124), .dinb(n23117), .dout(n23125));
  jnot g22980(.din(n23125), .dout(n23126));
  jand g22981(.dina(n16930), .dinb(n2936), .dout(n23127));
  jand g22982(.dina(n16592), .dinb(n2940), .dout(n23128));
  jand g22983(.dina(n16928), .dinb(n2943), .dout(n23129));
  jor  g22984(.dina(n23129), .dinb(n23128), .dout(n23130));
  jand g22985(.dina(n16343), .dinb(n3684), .dout(n23131));
  jor  g22986(.dina(n23131), .dinb(n23130), .dout(n23132));
  jor  g22987(.dina(n23132), .dinb(n23127), .dout(n23133));
  jxor g22988(.dina(n23133), .dinb(n93), .dout(n23134));
  jxor g22989(.dina(n23134), .dinb(n23126), .dout(n23135));
  jxor g22990(.dina(n23135), .dinb(n23100), .dout(n23136));
  jnot g22991(.din(n23136), .dout(n23137));
  jor  g22992(.dina(n23074), .dinb(n23115), .dout(n23138));
  jand g22993(.dina(n23075), .dinb(n23059), .dout(n23139));
  jnot g22994(.din(n23139), .dout(n23140));
  jand g22995(.dina(n23140), .dinb(n23138), .dout(n23141));
  jxor g22996(.dina(n23141), .dinb(n23137), .dout(n23142));
  jnot g22997(.din(n23142), .dout(n23143));
  jxor g22998(.dina(n23143), .dinb(n23095), .dout(n23144));
  jxor g22999(.dina(n23144), .dinb(n23079), .dout(n23145));
  jxor g23000(.dina(n23145), .dinb(n23091), .dout(n23146));
  jand g23001(.dina(n23146), .dinb(n6495), .dout(n23147));
  jand g23002(.dina(n23144), .dinb(n6503), .dout(n23148));
  jand g23003(.dina(n23079), .dinb(n6506), .dout(n23149));
  jand g23004(.dina(n23080), .dinb(n6500), .dout(n23150));
  jor  g23005(.dina(n23150), .dinb(n23149), .dout(n23151));
  jor  g23006(.dina(n23151), .dinb(n23148), .dout(n23152));
  jor  g23007(.dina(n23152), .dinb(n23147), .dout(n23153));
  jxor g23008(.dina(n23153), .dinb(n6219), .dout(n23154));
  jor  g23009(.dina(n23154), .dinb(n22950), .dout(n23155));
  jnot g23010(.din(n23155), .dout(n23156));
  jxor g23011(.dina(n23154), .dinb(n22950), .dout(n23157));
  jxor g23012(.dina(n22706), .dinb(n22705), .dout(n23158));
  jxor g23013(.dina(n23089), .dinb(n23088), .dout(n23159));
  jand g23014(.dina(n23159), .dinb(n6495), .dout(n23160));
  jand g23015(.dina(n23079), .dinb(n6503), .dout(n23161));
  jand g23016(.dina(n23080), .dinb(n6506), .dout(n23162));
  jand g23017(.dina(n22937), .dinb(n6500), .dout(n23163));
  jor  g23018(.dina(n23163), .dinb(n23162), .dout(n23164));
  jor  g23019(.dina(n23164), .dinb(n23161), .dout(n23165));
  jor  g23020(.dina(n23165), .dinb(n23160), .dout(n23166));
  jxor g23021(.dina(n23166), .dinb(n6219), .dout(n23167));
  jnot g23022(.din(n23167), .dout(n23168));
  jand g23023(.dina(n23168), .dinb(n23158), .dout(n23169));
  jor  g23024(.dina(n23168), .dinb(n23158), .dout(n23170));
  jxor g23025(.dina(n22703), .dinb(n22702), .dout(n23171));
  jxor g23026(.dina(n23086), .dinb(n23085), .dout(n23172));
  jand g23027(.dina(n23172), .dinb(n6495), .dout(n23173));
  jand g23028(.dina(n23080), .dinb(n6503), .dout(n23174));
  jand g23029(.dina(n22937), .dinb(n6506), .dout(n23175));
  jand g23030(.dina(n22265), .dinb(n6500), .dout(n23176));
  jor  g23031(.dina(n23176), .dinb(n23175), .dout(n23177));
  jor  g23032(.dina(n23177), .dinb(n23174), .dout(n23178));
  jor  g23033(.dina(n23178), .dinb(n23173), .dout(n23179));
  jxor g23034(.dina(n23179), .dinb(n6219), .dout(n23180));
  jnot g23035(.din(n23180), .dout(n23181));
  jand g23036(.dina(n23181), .dinb(n23171), .dout(n23182));
  jor  g23037(.dina(n23181), .dinb(n23171), .dout(n23183));
  jxor g23038(.dina(n22700), .dinb(n22698), .dout(n23184));
  jand g23039(.dina(n22939), .dinb(n6495), .dout(n23185));
  jand g23040(.dina(n22937), .dinb(n6503), .dout(n23186));
  jand g23041(.dina(n22265), .dinb(n6506), .dout(n23187));
  jand g23042(.dina(n22163), .dinb(n6500), .dout(n23188));
  jor  g23043(.dina(n23188), .dinb(n23187), .dout(n23189));
  jor  g23044(.dina(n23189), .dinb(n23186), .dout(n23190));
  jor  g23045(.dina(n23190), .dinb(n23185), .dout(n23191));
  jxor g23046(.dina(n23191), .dinb(n6219), .dout(n23192));
  jnot g23047(.din(n23192), .dout(n23193));
  jand g23048(.dina(n23193), .dinb(n23184), .dout(n23194));
  jor  g23049(.dina(n23193), .dinb(n23184), .dout(n23195));
  jxor g23050(.dina(n22696), .dinb(n22695), .dout(n23196));
  jand g23051(.dina(n22267), .dinb(n6495), .dout(n23197));
  jand g23052(.dina(n22265), .dinb(n6503), .dout(n23198));
  jand g23053(.dina(n22163), .dinb(n6506), .dout(n23199));
  jand g23054(.dina(n22164), .dinb(n6500), .dout(n23200));
  jor  g23055(.dina(n23200), .dinb(n23199), .dout(n23201));
  jor  g23056(.dina(n23201), .dinb(n23198), .dout(n23202));
  jor  g23057(.dina(n23202), .dinb(n23197), .dout(n23203));
  jxor g23058(.dina(n23203), .dinb(\a[2] ), .dout(n23204));
  jand g23059(.dina(n23204), .dinb(n23196), .dout(n23205));
  jor  g23060(.dina(n23204), .dinb(n23196), .dout(n23206));
  jxor g23061(.dina(n22693), .dinb(n22692), .dout(n23207));
  jand g23062(.dina(n22279), .dinb(n6495), .dout(n23208));
  jand g23063(.dina(n22163), .dinb(n6503), .dout(n23209));
  jand g23064(.dina(n22164), .dinb(n6506), .dout(n23210));
  jand g23065(.dina(n21974), .dinb(n6500), .dout(n23211));
  jor  g23066(.dina(n23211), .dinb(n23210), .dout(n23212));
  jor  g23067(.dina(n23212), .dinb(n23209), .dout(n23213));
  jor  g23068(.dina(n23213), .dinb(n23208), .dout(n23214));
  jxor g23069(.dina(n23214), .dinb(\a[2] ), .dout(n23215));
  jand g23070(.dina(n23215), .dinb(n23207), .dout(n23216));
  jor  g23071(.dina(n23215), .dinb(n23207), .dout(n23217));
  jxor g23072(.dina(n22686), .dinb(n22685), .dout(n23218));
  jnot g23073(.din(n23218), .dout(n23219));
  jnot g23074(.din(n21976), .dout(n23220));
  jor  g23075(.dina(n23220), .dinb(n6496), .dout(n23221));
  jnot g23076(.din(n21974), .dout(n23222));
  jor  g23077(.dina(n23222), .dinb(n6504), .dout(n23223));
  jnot g23078(.din(n21340), .dout(n23224));
  jor  g23079(.dina(n23224), .dinb(n6507), .dout(n23225));
  jnot g23080(.din(n21197), .dout(n23226));
  jor  g23081(.dina(n23226), .dinb(n6501), .dout(n23227));
  jand g23082(.dina(n23227), .dinb(n23225), .dout(n23228));
  jand g23083(.dina(n23228), .dinb(n23223), .dout(n23229));
  jand g23084(.dina(n23229), .dinb(n23221), .dout(n23230));
  jxor g23085(.dina(n23230), .dinb(\a[2] ), .dout(n23231));
  jand g23086(.dina(n23231), .dinb(n23219), .dout(n23232));
  jnot g23087(.din(n23232), .dout(n23233));
  jxor g23088(.dina(n22689), .dinb(n22688), .dout(n23234));
  jand g23089(.dina(n22291), .dinb(n6495), .dout(n23235));
  jand g23090(.dina(n22164), .dinb(n6503), .dout(n23236));
  jand g23091(.dina(n21974), .dinb(n6506), .dout(n23237));
  jand g23092(.dina(n21340), .dinb(n6500), .dout(n23238));
  jor  g23093(.dina(n23238), .dinb(n23237), .dout(n23239));
  jor  g23094(.dina(n23239), .dinb(n23236), .dout(n23240));
  jor  g23095(.dina(n23240), .dinb(n23235), .dout(n23241));
  jxor g23096(.dina(n23241), .dinb(\a[2] ), .dout(n23242));
  jor  g23097(.dina(n23242), .dinb(n23234), .dout(n23243));
  jnot g23098(.din(n23231), .dout(n23244));
  jand g23099(.dina(n23244), .dinb(n23218), .dout(n23245));
  jxor g23100(.dina(n22683), .dinb(n22682), .dout(n23246));
  jnot g23101(.din(n23246), .dout(n23247));
  jnot g23102(.din(n21342), .dout(n23248));
  jor  g23103(.dina(n23248), .dinb(n6496), .dout(n23249));
  jor  g23104(.dina(n23224), .dinb(n6504), .dout(n23250));
  jor  g23105(.dina(n23226), .dinb(n6507), .dout(n23251));
  jnot g23106(.din(n21198), .dout(n23252));
  jor  g23107(.dina(n23252), .dinb(n6501), .dout(n23253));
  jand g23108(.dina(n23253), .dinb(n23251), .dout(n23254));
  jand g23109(.dina(n23254), .dinb(n23250), .dout(n23255));
  jand g23110(.dina(n23255), .dinb(n23249), .dout(n23256));
  jxor g23111(.dina(n23256), .dinb(\a[2] ), .dout(n23257));
  jand g23112(.dina(n23257), .dinb(n23247), .dout(n23258));
  jnot g23113(.din(n23258), .dout(n23259));
  jnot g23114(.din(n23257), .dout(n23260));
  jand g23115(.dina(n23260), .dinb(n23246), .dout(n23261));
  jxor g23116(.dina(n22680), .dinb(n22679), .dout(n23262));
  jnot g23117(.din(n23262), .dout(n23263));
  jnot g23118(.din(n21355), .dout(n23264));
  jor  g23119(.dina(n23264), .dinb(n6496), .dout(n23265));
  jor  g23120(.dina(n23226), .dinb(n6504), .dout(n23266));
  jor  g23121(.dina(n23252), .dinb(n6507), .dout(n23267));
  jnot g23122(.din(n20947), .dout(n23268));
  jor  g23123(.dina(n23268), .dinb(n6501), .dout(n23269));
  jand g23124(.dina(n23269), .dinb(n23267), .dout(n23270));
  jand g23125(.dina(n23270), .dinb(n23266), .dout(n23271));
  jand g23126(.dina(n23271), .dinb(n23265), .dout(n23272));
  jxor g23127(.dina(n23272), .dinb(\a[2] ), .dout(n23273));
  jand g23128(.dina(n23273), .dinb(n23263), .dout(n23274));
  jnot g23129(.din(n23274), .dout(n23275));
  jnot g23130(.din(n23273), .dout(n23276));
  jand g23131(.dina(n23276), .dinb(n23262), .dout(n23277));
  jxor g23132(.dina(n22677), .dinb(n22676), .dout(n23278));
  jand g23133(.dina(n21367), .dinb(n6495), .dout(n23279));
  jand g23134(.dina(n21198), .dinb(n6503), .dout(n23280));
  jand g23135(.dina(n20947), .dinb(n6506), .dout(n23281));
  jand g23136(.dina(n20344), .dinb(n6500), .dout(n23282));
  jor  g23137(.dina(n23282), .dinb(n23281), .dout(n23283));
  jor  g23138(.dina(n23283), .dinb(n23280), .dout(n23284));
  jor  g23139(.dina(n23284), .dinb(n23279), .dout(n23285));
  jxor g23140(.dina(n23285), .dinb(\a[2] ), .dout(n23286));
  jand g23141(.dina(n23286), .dinb(n23278), .dout(n23287));
  jor  g23142(.dina(n23286), .dinb(n23278), .dout(n23288));
  jxor g23143(.dina(n22674), .dinb(n22673), .dout(n23289));
  jand g23144(.dina(n20949), .dinb(n6495), .dout(n23290));
  jand g23145(.dina(n20947), .dinb(n6503), .dout(n23291));
  jand g23146(.dina(n20344), .dinb(n6506), .dout(n23292));
  jand g23147(.dina(n20204), .dinb(n6500), .dout(n23293));
  jor  g23148(.dina(n23293), .dinb(n23292), .dout(n23294));
  jor  g23149(.dina(n23294), .dinb(n23291), .dout(n23295));
  jor  g23150(.dina(n23295), .dinb(n23290), .dout(n23296));
  jxor g23151(.dina(n23296), .dinb(\a[2] ), .dout(n23297));
  jand g23152(.dina(n23297), .dinb(n23289), .dout(n23298));
  jxor g23153(.dina(n22671), .dinb(n22670), .dout(n23299));
  jxor g23154(.dina(n22668), .dinb(n22667), .dout(n23300));
  jand g23155(.dina(n20358), .dinb(n6495), .dout(n23301));
  jand g23156(.dina(n20204), .dinb(n6503), .dout(n23302));
  jand g23157(.dina(n20205), .dinb(n6506), .dout(n23303));
  jand g23158(.dina(n19922), .dinb(n6500), .dout(n23304));
  jor  g23159(.dina(n23304), .dinb(n23303), .dout(n23305));
  jor  g23160(.dina(n23305), .dinb(n23302), .dout(n23306));
  jor  g23161(.dina(n23306), .dinb(n23301), .dout(n23307));
  jxor g23162(.dina(n23307), .dinb(n6219), .dout(n23308));
  jnot g23163(.din(n23308), .dout(n23309));
  jand g23164(.dina(n23309), .dinb(n23300), .dout(n23310));
  jxor g23165(.dina(n22665), .dinb(n22664), .dout(n23311));
  jxor g23166(.dina(n22662), .dinb(n22661), .dout(n23312));
  jand g23167(.dina(n19924), .dinb(n6495), .dout(n23313));
  jand g23168(.dina(n19922), .dinb(n6503), .dout(n23314));
  jand g23169(.dina(n19373), .dinb(n6506), .dout(n23315));
  jand g23170(.dina(n19219), .dinb(n6500), .dout(n23316));
  jor  g23171(.dina(n23316), .dinb(n23315), .dout(n23317));
  jor  g23172(.dina(n23317), .dinb(n23314), .dout(n23318));
  jor  g23173(.dina(n23318), .dinb(n23313), .dout(n23319));
  jxor g23174(.dina(n23319), .dinb(\a[2] ), .dout(n23320));
  jand g23175(.dina(n23320), .dinb(n23312), .dout(n23321));
  jor  g23176(.dina(n23320), .dinb(n23312), .dout(n23322));
  jxor g23177(.dina(n22659), .dinb(n22658), .dout(n23323));
  jand g23178(.dina(n19375), .dinb(n6495), .dout(n23324));
  jand g23179(.dina(n19373), .dinb(n6503), .dout(n23325));
  jand g23180(.dina(n19219), .dinb(n6506), .dout(n23326));
  jand g23181(.dina(n19220), .dinb(n6500), .dout(n23327));
  jor  g23182(.dina(n23327), .dinb(n23326), .dout(n23328));
  jor  g23183(.dina(n23328), .dinb(n23325), .dout(n23329));
  jor  g23184(.dina(n23329), .dinb(n23324), .dout(n23330));
  jxor g23185(.dina(n23330), .dinb(\a[2] ), .dout(n23331));
  jand g23186(.dina(n23331), .dinb(n23323), .dout(n23332));
  jor  g23187(.dina(n23331), .dinb(n23323), .dout(n23333));
  jxor g23188(.dina(n22656), .dinb(n22655), .dout(n23334));
  jand g23189(.dina(n19387), .dinb(n6495), .dout(n23335));
  jand g23190(.dina(n19219), .dinb(n6503), .dout(n23336));
  jand g23191(.dina(n19220), .dinb(n6506), .dout(n23337));
  jand g23192(.dina(n18914), .dinb(n6500), .dout(n23338));
  jor  g23193(.dina(n23338), .dinb(n23337), .dout(n23339));
  jor  g23194(.dina(n23339), .dinb(n23336), .dout(n23340));
  jor  g23195(.dina(n23340), .dinb(n23335), .dout(n23341));
  jxor g23196(.dina(n23341), .dinb(\a[2] ), .dout(n23342));
  jand g23197(.dina(n23342), .dinb(n23334), .dout(n23343));
  jor  g23198(.dina(n23342), .dinb(n23334), .dout(n23344));
  jxor g23199(.dina(n22653), .dinb(n22652), .dout(n23345));
  jand g23200(.dina(n19399), .dinb(n6495), .dout(n23346));
  jand g23201(.dina(n19220), .dinb(n6503), .dout(n23347));
  jand g23202(.dina(n18914), .dinb(n6506), .dout(n23348));
  jand g23203(.dina(n18488), .dinb(n6500), .dout(n23349));
  jor  g23204(.dina(n23349), .dinb(n23348), .dout(n23350));
  jor  g23205(.dina(n23350), .dinb(n23347), .dout(n23351));
  jor  g23206(.dina(n23351), .dinb(n23346), .dout(n23352));
  jxor g23207(.dina(n23352), .dinb(n6219), .dout(n23353));
  jnot g23208(.din(n23353), .dout(n23354));
  jand g23209(.dina(n23354), .dinb(n23345), .dout(n23355));
  jor  g23210(.dina(n23354), .dinb(n23345), .dout(n23356));
  jxor g23211(.dina(n22650), .dinb(n22649), .dout(n23357));
  jand g23212(.dina(n18916), .dinb(n6495), .dout(n23358));
  jand g23213(.dina(n18914), .dinb(n6503), .dout(n23359));
  jand g23214(.dina(n18488), .dinb(n6506), .dout(n23360));
  jand g23215(.dina(n18292), .dinb(n6500), .dout(n23361));
  jor  g23216(.dina(n23361), .dinb(n23360), .dout(n23362));
  jor  g23217(.dina(n23362), .dinb(n23359), .dout(n23363));
  jor  g23218(.dina(n23363), .dinb(n23358), .dout(n23364));
  jxor g23219(.dina(n23364), .dinb(n6219), .dout(n23365));
  jnot g23220(.din(n23365), .dout(n23366));
  jand g23221(.dina(n23366), .dinb(n23357), .dout(n23367));
  jor  g23222(.dina(n23366), .dinb(n23357), .dout(n23368));
  jxor g23223(.dina(n22645), .dinb(n22644), .dout(n23369));
  jand g23224(.dina(n18490), .dinb(n6495), .dout(n23370));
  jand g23225(.dina(n18488), .dinb(n6503), .dout(n23371));
  jand g23226(.dina(n18292), .dinb(n6506), .dout(n23372));
  jand g23227(.dina(n18293), .dinb(n6500), .dout(n23373));
  jor  g23228(.dina(n23373), .dinb(n23372), .dout(n23374));
  jor  g23229(.dina(n23374), .dinb(n23371), .dout(n23375));
  jor  g23230(.dina(n23375), .dinb(n23370), .dout(n23376));
  jxor g23231(.dina(n23376), .dinb(\a[2] ), .dout(n23377));
  jand g23232(.dina(n23377), .dinb(n23369), .dout(n23378));
  jxor g23233(.dina(n22640), .dinb(n22639), .dout(n23379));
  jnot g23234(.din(n23379), .dout(n23380));
  jnot g23235(.din(n18502), .dout(n23381));
  jor  g23236(.dina(n23381), .dinb(n6496), .dout(n23382));
  jnot g23237(.din(n18292), .dout(n23383));
  jor  g23238(.dina(n23383), .dinb(n6504), .dout(n23384));
  jnot g23239(.din(n18293), .dout(n23385));
  jor  g23240(.dina(n23385), .dinb(n6507), .dout(n23386));
  jnot g23241(.din(n17942), .dout(n23387));
  jor  g23242(.dina(n23387), .dinb(n6501), .dout(n23388));
  jand g23243(.dina(n23388), .dinb(n23386), .dout(n23389));
  jand g23244(.dina(n23389), .dinb(n23384), .dout(n23390));
  jand g23245(.dina(n23390), .dinb(n23382), .dout(n23391));
  jxor g23246(.dina(n23391), .dinb(n6219), .dout(n23392));
  jnot g23247(.din(n23392), .dout(n23393));
  jand g23248(.dina(n23393), .dinb(n23380), .dout(n23394));
  jnot g23249(.din(n23394), .dout(n23395));
  jxor g23250(.dina(n22630), .dinb(n22629), .dout(n23396));
  jxor g23251(.dina(n22625), .dinb(n22624), .dout(n23397));
  jnot g23252(.din(n23397), .dout(n23398));
  jxor g23253(.dina(n22620), .dinb(n22619), .dout(n23399));
  jand g23254(.dina(n17549), .dinb(n6495), .dout(n23400));
  jand g23255(.dina(n17329), .dinb(n6503), .dout(n23401));
  jand g23256(.dina(n17330), .dinb(n6506), .dout(n23402));
  jand g23257(.dina(n16940), .dinb(n6500), .dout(n23403));
  jor  g23258(.dina(n23403), .dinb(n23402), .dout(n23404));
  jor  g23259(.dina(n23404), .dinb(n23401), .dout(n23405));
  jor  g23260(.dina(n23405), .dinb(n23400), .dout(n23406));
  jxor g23261(.dina(n23406), .dinb(n6219), .dout(n23407));
  jnot g23262(.din(n23407), .dout(n23408));
  jand g23263(.dina(n23408), .dinb(n23399), .dout(n23409));
  jor  g23264(.dina(n23408), .dinb(n23399), .dout(n23410));
  jxor g23265(.dina(n22617), .dinb(n22616), .dout(n23411));
  jnot g23266(.din(n23411), .dout(n23412));
  jand g23267(.dina(n17561), .dinb(n6495), .dout(n23413));
  jand g23268(.dina(n17330), .dinb(n6503), .dout(n23414));
  jand g23269(.dina(n16940), .dinb(n6506), .dout(n23415));
  jand g23270(.dina(n16604), .dinb(n6500), .dout(n23416));
  jor  g23271(.dina(n23416), .dinb(n23415), .dout(n23417));
  jor  g23272(.dina(n23417), .dinb(n23414), .dout(n23418));
  jor  g23273(.dina(n23418), .dinb(n23413), .dout(n23419));
  jxor g23274(.dina(n23419), .dinb(n6219), .dout(n23420));
  jand g23275(.dina(n23420), .dinb(n23412), .dout(n23421));
  jor  g23276(.dina(n23420), .dinb(n23412), .dout(n23422));
  jxor g23277(.dina(n22612), .dinb(n22611), .dout(n23423));
  jnot g23278(.din(n23423), .dout(n23424));
  jnot g23279(.din(n16942), .dout(n23425));
  jor  g23280(.dina(n23425), .dinb(n6496), .dout(n23426));
  jnot g23281(.din(n16940), .dout(n23427));
  jor  g23282(.dina(n23427), .dinb(n6504), .dout(n23428));
  jnot g23283(.din(n16604), .dout(n23429));
  jor  g23284(.dina(n23429), .dinb(n6507), .dout(n23430));
  jnot g23285(.din(n16355), .dout(n23431));
  jor  g23286(.dina(n23431), .dinb(n6501), .dout(n23432));
  jand g23287(.dina(n23432), .dinb(n23430), .dout(n23433));
  jand g23288(.dina(n23433), .dinb(n23428), .dout(n23434));
  jand g23289(.dina(n23434), .dinb(n23426), .dout(n23435));
  jxor g23290(.dina(n23435), .dinb(n6219), .dout(n23436));
  jnot g23291(.din(n23436), .dout(n23437));
  jand g23292(.dina(n23437), .dinb(n23424), .dout(n23438));
  jand g23293(.dina(n23436), .dinb(n23423), .dout(n23439));
  jnot g23294(.din(n23439), .dout(n23440));
  jxor g23295(.dina(n22608), .dinb(n22600), .dout(n23441));
  jnot g23296(.din(n23441), .dout(n23442));
  jand g23297(.dina(n16606), .dinb(n6495), .dout(n23443));
  jand g23298(.dina(n16604), .dinb(n6503), .dout(n23444));
  jand g23299(.dina(n16355), .dinb(n6506), .dout(n23445));
  jand g23300(.dina(n16360), .dinb(n6500), .dout(n23446));
  jor  g23301(.dina(n23446), .dinb(n23445), .dout(n23447));
  jor  g23302(.dina(n23447), .dinb(n23444), .dout(n23448));
  jor  g23303(.dina(n23448), .dinb(n23443), .dout(n23449));
  jxor g23304(.dina(n23449), .dinb(n6219), .dout(n23450));
  jand g23305(.dina(n23450), .dinb(n23442), .dout(n23451));
  jor  g23306(.dina(n23450), .dinb(n23442), .dout(n23452));
  jor  g23307(.dina(n22587), .dinb(n5277), .dout(n23453));
  jxor g23308(.dina(n23453), .dinb(n22595), .dout(n23454));
  jand g23309(.dina(n16616), .dinb(n6495), .dout(n23455));
  jand g23310(.dina(n16355), .dinb(n6503), .dout(n23456));
  jand g23311(.dina(n16360), .dinb(n6506), .dout(n23457));
  jand g23312(.dina(n15841), .dinb(n6500), .dout(n23458));
  jor  g23313(.dina(n23458), .dinb(n23457), .dout(n23459));
  jor  g23314(.dina(n23459), .dinb(n23456), .dout(n23460));
  jor  g23315(.dina(n23460), .dinb(n23455), .dout(n23461));
  jxor g23316(.dina(n23461), .dinb(\a[2] ), .dout(n23462));
  jand g23317(.dina(n23462), .dinb(n23454), .dout(n23463));
  jand g23318(.dina(n15579), .dinb(n6503), .dout(n23464));
  jnot g23319(.din(n23464), .dout(n23465));
  jand g23320(.dina(n15843), .dinb(n15020), .dout(n23466));
  jnot g23321(.din(n23466), .dout(n23467));
  jnot g23322(.din(n15340), .dout(n23468));
  jand g23323(.dina(n15844), .dinb(n23468), .dout(n23469));
  jand g23324(.dina(n23469), .dinb(n23467), .dout(n23470));
  jor  g23325(.dina(n23470), .dinb(n6861), .dout(n23471));
  jand g23326(.dina(n15022), .dinb(\a[2] ), .dout(n23472));
  jand g23327(.dina(n15327), .dinb(n6856), .dout(n23473));
  jnot g23328(.din(n23473), .dout(n23474));
  jand g23329(.dina(n23474), .dinb(n23472), .dout(n23475));
  jand g23330(.dina(n23475), .dinb(n23471), .dout(n23476));
  jand g23331(.dina(n23476), .dinb(n23465), .dout(n23477));
  jor  g23332(.dina(n23477), .dinb(n22584), .dout(n23479));
  jand g23333(.dina(n15848), .dinb(n6495), .dout(n23480));
  jand g23334(.dina(n15841), .dinb(n6503), .dout(n23481));
  jand g23335(.dina(n15579), .dinb(n6506), .dout(n23482));
  jand g23336(.dina(n15327), .dinb(n6500), .dout(n23483));
  jor  g23337(.dina(n23483), .dinb(n23482), .dout(n23484));
  jor  g23338(.dina(n23484), .dinb(n23481), .dout(n23485));
  jor  g23339(.dina(n23485), .dinb(n23480), .dout(n23486));
  jxor g23340(.dina(n23486), .dinb(n6219), .dout(n23487));
  jnot g23341(.din(n23487), .dout(n23488));
  jand g23342(.dina(n23488), .dinb(n23479), .dout(n23489));
  jand g23343(.dina(n16632), .dinb(n6495), .dout(n23491));
  jand g23344(.dina(n16360), .dinb(n6503), .dout(n23492));
  jand g23345(.dina(n15841), .dinb(n6506), .dout(n23493));
  jand g23346(.dina(n15579), .dinb(n6500), .dout(n23494));
  jor  g23347(.dina(n23494), .dinb(n23493), .dout(n23495));
  jor  g23348(.dina(n23495), .dinb(n23492), .dout(n23496));
  jor  g23349(.dina(n23496), .dinb(n23491), .dout(n23497));
  jxor g23350(.dina(n23497), .dinb(n6219), .dout(n23498));
  jnot g23351(.din(n23498), .dout(n23499));
  jand g23352(.dina(n23499), .dinb(n23489), .dout(n23500));
  jor  g23353(.dina(n23499), .dinb(n23489), .dout(n23501));
  jand g23354(.dina(n22584), .dinb(\a[5] ), .dout(n23502));
  jxor g23355(.dina(n23502), .dinb(n22582), .dout(n23503));
  jand g23356(.dina(n23503), .dinb(n23501), .dout(n23504));
  jor  g23357(.dina(n23504), .dinb(n23500), .dout(n23505));
  jor  g23358(.dina(n23462), .dinb(n23454), .dout(n23506));
  jand g23359(.dina(n23506), .dinb(n23505), .dout(n23507));
  jor  g23360(.dina(n23507), .dinb(n23463), .dout(n23508));
  jnot g23361(.din(n23508), .dout(n23509));
  jand g23362(.dina(n23509), .dinb(n23452), .dout(n23510));
  jor  g23363(.dina(n23510), .dinb(n23451), .dout(n23511));
  jand g23364(.dina(n23511), .dinb(n23440), .dout(n23512));
  jor  g23365(.dina(n23512), .dinb(n23438), .dout(n23513));
  jand g23366(.dina(n23513), .dinb(n23422), .dout(n23514));
  jor  g23367(.dina(n23514), .dinb(n23421), .dout(n23515));
  jnot g23368(.din(n23515), .dout(n23516));
  jand g23369(.dina(n23516), .dinb(n23410), .dout(n23517));
  jor  g23370(.dina(n23517), .dinb(n23409), .dout(n23518));
  jnot g23371(.din(n23518), .dout(n23519));
  jand g23372(.dina(n23519), .dinb(n23398), .dout(n23520));
  jand g23373(.dina(n23518), .dinb(n23397), .dout(n23521));
  jnot g23374(.din(n23521), .dout(n23522));
  jand g23375(.dina(n17537), .dinb(n6495), .dout(n23523));
  jand g23376(.dina(n17535), .dinb(n6503), .dout(n23524));
  jand g23377(.dina(n17329), .dinb(n6506), .dout(n23525));
  jand g23378(.dina(n17330), .dinb(n6500), .dout(n23526));
  jor  g23379(.dina(n23526), .dinb(n23525), .dout(n23527));
  jor  g23380(.dina(n23527), .dinb(n23524), .dout(n23528));
  jor  g23381(.dina(n23528), .dinb(n23523), .dout(n23529));
  jxor g23382(.dina(n23529), .dinb(n6219), .dout(n23530));
  jand g23383(.dina(n23530), .dinb(n23522), .dout(n23531));
  jor  g23384(.dina(n23531), .dinb(n23520), .dout(n23532));
  jnot g23385(.din(n23532), .dout(n23533));
  jand g23386(.dina(n23533), .dinb(n23396), .dout(n23534));
  jand g23387(.dina(n17944), .dinb(n6495), .dout(n23535));
  jand g23388(.dina(n17942), .dinb(n6503), .dout(n23536));
  jand g23389(.dina(n17535), .dinb(n6506), .dout(n23537));
  jand g23390(.dina(n17329), .dinb(n6500), .dout(n23538));
  jor  g23391(.dina(n23538), .dinb(n23537), .dout(n23539));
  jor  g23392(.dina(n23539), .dinb(n23536), .dout(n23540));
  jor  g23393(.dina(n23540), .dinb(n23535), .dout(n23541));
  jxor g23394(.dina(n23541), .dinb(\a[2] ), .dout(n23542));
  jor  g23395(.dina(n23542), .dinb(n23534), .dout(n23543));
  jor  g23396(.dina(n23533), .dinb(n23396), .dout(n23544));
  jxor g23397(.dina(n22635), .dinb(n22634), .dout(n23545));
  jnot g23398(.din(n23545), .dout(n23546));
  jnot g23399(.din(n18514), .dout(n23547));
  jor  g23400(.dina(n23547), .dinb(n6496), .dout(n23548));
  jor  g23401(.dina(n23385), .dinb(n6504), .dout(n23549));
  jor  g23402(.dina(n23387), .dinb(n6507), .dout(n23550));
  jnot g23403(.din(n17535), .dout(n23551));
  jor  g23404(.dina(n23551), .dinb(n6501), .dout(n23552));
  jand g23405(.dina(n23552), .dinb(n23550), .dout(n23553));
  jand g23406(.dina(n23553), .dinb(n23549), .dout(n23554));
  jand g23407(.dina(n23554), .dinb(n23548), .dout(n23555));
  jxor g23408(.dina(n23555), .dinb(n6219), .dout(n23556));
  jnot g23409(.din(n23556), .dout(n23557));
  jand g23410(.dina(n23557), .dinb(n23546), .dout(n23558));
  jnot g23411(.din(n23558), .dout(n23559));
  jand g23412(.dina(n23559), .dinb(n23544), .dout(n23560));
  jand g23413(.dina(n23560), .dinb(n23543), .dout(n23561));
  jand g23414(.dina(n23556), .dinb(n23545), .dout(n23562));
  jor  g23415(.dina(n23562), .dinb(n23561), .dout(n23563));
  jand g23416(.dina(n23392), .dinb(n23379), .dout(n23564));
  jor  g23417(.dina(n23564), .dinb(n23563), .dout(n23565));
  jand g23418(.dina(n23565), .dinb(n23395), .dout(n23566));
  jor  g23419(.dina(n23377), .dinb(n23369), .dout(n23567));
  jand g23420(.dina(n23567), .dinb(n23566), .dout(n23568));
  jor  g23421(.dina(n23568), .dinb(n23378), .dout(n23569));
  jand g23422(.dina(n23569), .dinb(n23368), .dout(n23570));
  jor  g23423(.dina(n23570), .dinb(n23367), .dout(n23571));
  jand g23424(.dina(n23571), .dinb(n23356), .dout(n23572));
  jor  g23425(.dina(n23572), .dinb(n23355), .dout(n23573));
  jand g23426(.dina(n23573), .dinb(n23344), .dout(n23574));
  jor  g23427(.dina(n23574), .dinb(n23343), .dout(n23575));
  jand g23428(.dina(n23575), .dinb(n23333), .dout(n23576));
  jor  g23429(.dina(n23576), .dinb(n23332), .dout(n23577));
  jand g23430(.dina(n23577), .dinb(n23322), .dout(n23578));
  jor  g23431(.dina(n23578), .dinb(n23321), .dout(n23579));
  jand g23432(.dina(n23579), .dinb(n23311), .dout(n23580));
  jand g23433(.dina(n20371), .dinb(n6495), .dout(n23581));
  jand g23434(.dina(n20205), .dinb(n6503), .dout(n23582));
  jand g23435(.dina(n19922), .dinb(n6506), .dout(n23583));
  jand g23436(.dina(n19373), .dinb(n6500), .dout(n23584));
  jor  g23437(.dina(n23584), .dinb(n23583), .dout(n23585));
  jor  g23438(.dina(n23585), .dinb(n23582), .dout(n23586));
  jor  g23439(.dina(n23586), .dinb(n23581), .dout(n23587));
  jxor g23440(.dina(n23587), .dinb(n6219), .dout(n23588));
  jnot g23441(.din(n23588), .dout(n23589));
  jor  g23442(.dina(n23589), .dinb(n23580), .dout(n23590));
  jor  g23443(.dina(n23579), .dinb(n23311), .dout(n23591));
  jor  g23444(.dina(n23309), .dinb(n23300), .dout(n23592));
  jand g23445(.dina(n23592), .dinb(n23591), .dout(n23593));
  jand g23446(.dina(n23593), .dinb(n23590), .dout(n23594));
  jor  g23447(.dina(n23594), .dinb(n23310), .dout(n23595));
  jand g23448(.dina(n23595), .dinb(n23299), .dout(n23596));
  jand g23449(.dina(n20346), .dinb(n6495), .dout(n23597));
  jand g23450(.dina(n20344), .dinb(n6503), .dout(n23598));
  jand g23451(.dina(n20204), .dinb(n6506), .dout(n23599));
  jand g23452(.dina(n20205), .dinb(n6500), .dout(n23600));
  jor  g23453(.dina(n23600), .dinb(n23599), .dout(n23601));
  jor  g23454(.dina(n23601), .dinb(n23598), .dout(n23602));
  jor  g23455(.dina(n23602), .dinb(n23597), .dout(n23603));
  jxor g23456(.dina(n23603), .dinb(n6219), .dout(n23604));
  jnot g23457(.din(n23604), .dout(n23605));
  jor  g23458(.dina(n23605), .dinb(n23596), .dout(n23606));
  jor  g23459(.dina(n23297), .dinb(n23289), .dout(n23607));
  jor  g23460(.dina(n23595), .dinb(n23299), .dout(n23608));
  jand g23461(.dina(n23608), .dinb(n23607), .dout(n23609));
  jand g23462(.dina(n23609), .dinb(n23606), .dout(n23610));
  jor  g23463(.dina(n23610), .dinb(n23298), .dout(n23611));
  jand g23464(.dina(n23611), .dinb(n23288), .dout(n23612));
  jor  g23465(.dina(n23612), .dinb(n23287), .dout(n23613));
  jor  g23466(.dina(n23613), .dinb(n23277), .dout(n23614));
  jand g23467(.dina(n23614), .dinb(n23275), .dout(n23615));
  jor  g23468(.dina(n23615), .dinb(n23261), .dout(n23616));
  jand g23469(.dina(n23616), .dinb(n23259), .dout(n23617));
  jor  g23470(.dina(n23617), .dinb(n23245), .dout(n23618));
  jand g23471(.dina(n23618), .dinb(n23243), .dout(n23619));
  jand g23472(.dina(n23619), .dinb(n23233), .dout(n23620));
  jand g23473(.dina(n23242), .dinb(n23234), .dout(n23621));
  jor  g23474(.dina(n23621), .dinb(n23620), .dout(n23622));
  jand g23475(.dina(n23622), .dinb(n23217), .dout(n23623));
  jor  g23476(.dina(n23623), .dinb(n23216), .dout(n23624));
  jand g23477(.dina(n23624), .dinb(n23206), .dout(n23625));
  jor  g23478(.dina(n23625), .dinb(n23205), .dout(n23626));
  jand g23479(.dina(n23626), .dinb(n23195), .dout(n23627));
  jor  g23480(.dina(n23627), .dinb(n23194), .dout(n23628));
  jand g23481(.dina(n23628), .dinb(n23183), .dout(n23629));
  jor  g23482(.dina(n23629), .dinb(n23182), .dout(n23630));
  jand g23483(.dina(n23630), .dinb(n23170), .dout(n23631));
  jor  g23484(.dina(n23631), .dinb(n23169), .dout(n23632));
  jand g23485(.dina(n23632), .dinb(n23157), .dout(n23633));
  jor  g23486(.dina(n23633), .dinb(n23156), .dout(n23634));
  jnot g23487(.din(n22860), .dout(n23635));
  jor  g23488(.dina(n22947), .dinb(n23635), .dout(n23636));
  jor  g23489(.dina(n22948), .dinb(n22708), .dout(n23637));
  jand g23490(.dina(n23637), .dinb(n23636), .dout(n23638));
  jnot g23491(.din(n22849), .dout(n23639));
  jor  g23492(.dina(n22857), .dinb(n23639), .dout(n23640));
  jnot g23493(.din(n21724), .dout(n23641));
  jor  g23494(.dina(n21985), .dinb(n23641), .dout(n23642));
  jand g23495(.dina(n23642), .dinb(n22710), .dout(n23643));
  jor  g23496(.dina(n22858), .dinb(n23643), .dout(n23644));
  jand g23497(.dina(n23644), .dinb(n23640), .dout(n23645));
  jnot g23498(.din(n22838), .dout(n23646));
  jor  g23499(.dina(n22846), .dinb(n23646), .dout(n23647));
  jnot g23500(.din(n23647), .dout(n23648));
  jand g23501(.dina(n22848), .dinb(n22718), .dout(n23649));
  jor  g23502(.dina(n23649), .dinb(n23648), .dout(n23650));
  jor  g23503(.dina(n22836), .dinb(n22828), .dout(n23651));
  jnot g23504(.din(n23651), .dout(n23652));
  jand g23505(.dina(n22837), .dinb(n22722), .dout(n23653));
  jor  g23506(.dina(n23653), .dinb(n23652), .dout(n23654));
  jand g23507(.dina(n22825), .dinb(n22817), .dout(n23655));
  jand g23508(.dina(n22826), .dinb(n22727), .dout(n23656));
  jor  g23509(.dina(n23656), .dinb(n23655), .dout(n23657));
  jor  g23510(.dina(n22815), .dinb(n22807), .dout(n23658));
  jand g23511(.dina(n22816), .dinb(n22732), .dout(n23659));
  jnot g23512(.din(n23659), .dout(n23660));
  jand g23513(.dina(n23660), .dinb(n23658), .dout(n23661));
  jnot g23514(.din(n23661), .dout(n23662));
  jand g23515(.dina(n22804), .dinb(n22796), .dout(n23663));
  jand g23516(.dina(n22805), .dinb(n22737), .dout(n23664));
  jor  g23517(.dina(n23664), .dinb(n23663), .dout(n23665));
  jor  g23518(.dina(n22794), .dinb(n22786), .dout(n23666));
  jand g23519(.dina(n22795), .dinb(n22742), .dout(n23667));
  jnot g23520(.din(n23667), .dout(n23668));
  jand g23521(.dina(n23668), .dinb(n23666), .dout(n23669));
  jnot g23522(.din(n23669), .dout(n23670));
  jor  g23523(.dina(n22783), .dinb(n22775), .dout(n23671));
  jand g23524(.dina(n22784), .dinb(n22747), .dout(n23672));
  jnot g23525(.din(n23672), .dout(n23673));
  jand g23526(.dina(n23673), .dinb(n23671), .dout(n23674));
  jnot g23527(.din(n23674), .dout(n23675));
  jand g23528(.dina(n22772), .dinb(n22765), .dout(n23676));
  jand g23529(.dina(n22773), .dinb(n22750), .dout(n23677));
  jor  g23530(.dina(n23677), .dinb(n23676), .dout(n23678));
  jand g23531(.dina(n2127), .dinb(n510), .dout(n23679));
  jand g23532(.dina(n23679), .dinb(n11398), .dout(n23680));
  jand g23533(.dina(n23680), .dinb(n1843), .dout(n23681));
  jand g23534(.dina(n1782), .dinb(n496), .dout(n23682));
  jand g23535(.dina(n13544), .dinb(n557), .dout(n23683));
  jand g23536(.dina(n23683), .dinb(n23682), .dout(n23684));
  jand g23537(.dina(n1772), .dinb(n1213), .dout(n23685));
  jand g23538(.dina(n1915), .dinb(n1326), .dout(n23686));
  jand g23539(.dina(n23686), .dinb(n23685), .dout(n23687));
  jand g23540(.dina(n23687), .dinb(n23684), .dout(n23688));
  jand g23541(.dina(n23688), .dinb(n21023), .dout(n23689));
  jand g23542(.dina(n23689), .dinb(n23681), .dout(n23690));
  jand g23543(.dina(n23690), .dinb(n13202), .dout(n23691));
  jand g23544(.dina(n20851), .dinb(n11240), .dout(n23692));
  jand g23545(.dina(n23692), .dinb(n23691), .dout(n23693));
  jnot g23546(.din(n23693), .dout(n23694));
  jand g23547(.dina(n16616), .dinb(n5076), .dout(n23695));
  jand g23548(.dina(n16355), .dinb(n5084), .dout(n23696));
  jand g23549(.dina(n15841), .dinb(n6050), .dout(n23697));
  jand g23550(.dina(n16360), .dinb(n5082), .dout(n23698));
  jor  g23551(.dina(n23698), .dinb(n23697), .dout(n23699));
  jor  g23552(.dina(n23699), .dinb(n23696), .dout(n23700));
  jor  g23553(.dina(n23700), .dinb(n23695), .dout(n23701));
  jxor g23554(.dina(n23701), .dinb(n23694), .dout(n23702));
  jxor g23555(.dina(n23702), .dinb(n23678), .dout(n23703));
  jnot g23556(.din(n23703), .dout(n23704));
  jand g23557(.dina(n17561), .dinb(n2936), .dout(n23705));
  jand g23558(.dina(n16940), .dinb(n2940), .dout(n23706));
  jand g23559(.dina(n17330), .dinb(n2943), .dout(n23707));
  jor  g23560(.dina(n23707), .dinb(n23706), .dout(n23708));
  jand g23561(.dina(n16604), .dinb(n3684), .dout(n23709));
  jor  g23562(.dina(n23709), .dinb(n23708), .dout(n23710));
  jor  g23563(.dina(n23710), .dinb(n23705), .dout(n23711));
  jxor g23564(.dina(n23711), .dinb(n93), .dout(n23712));
  jxor g23565(.dina(n23712), .dinb(n23704), .dout(n23713));
  jxor g23566(.dina(n23713), .dinb(n23675), .dout(n23714));
  jnot g23567(.din(n23714), .dout(n23715));
  jand g23568(.dina(n17944), .dinb(n71), .dout(n23716));
  jand g23569(.dina(n17942), .dinb(n796), .dout(n23717));
  jand g23570(.dina(n17535), .dinb(n731), .dout(n23718));
  jand g23571(.dina(n17329), .dinb(n1806), .dout(n23719));
  jor  g23572(.dina(n23719), .dinb(n23718), .dout(n23720));
  jor  g23573(.dina(n23720), .dinb(n23717), .dout(n23721));
  jor  g23574(.dina(n23721), .dinb(n23716), .dout(n23722));
  jxor g23575(.dina(n23722), .dinb(n77), .dout(n23723));
  jxor g23576(.dina(n23723), .dinb(n23715), .dout(n23724));
  jxor g23577(.dina(n23724), .dinb(n23670), .dout(n23725));
  jnot g23578(.din(n23725), .dout(n23726));
  jand g23579(.dina(n18490), .dinb(n806), .dout(n23727));
  jand g23580(.dina(n18488), .dinb(n1620), .dout(n23728));
  jand g23581(.dina(n18292), .dinb(n1612), .dout(n23729));
  jand g23582(.dina(n18293), .dinb(n1644), .dout(n23730));
  jor  g23583(.dina(n23730), .dinb(n23729), .dout(n23731));
  jor  g23584(.dina(n23731), .dinb(n23728), .dout(n23732));
  jor  g23585(.dina(n23732), .dinb(n23727), .dout(n23733));
  jxor g23586(.dina(n23733), .dinb(n65), .dout(n23734));
  jxor g23587(.dina(n23734), .dinb(n23726), .dout(n23735));
  jxor g23588(.dina(n23735), .dinb(n23665), .dout(n23736));
  jnot g23589(.din(n23736), .dout(n23737));
  jand g23590(.dina(n19387), .dinb(n1819), .dout(n23738));
  jand g23591(.dina(n19220), .dinb(n2180), .dout(n23739));
  jand g23592(.dina(n19219), .dinb(n2243), .dout(n23740));
  jor  g23593(.dina(n23740), .dinb(n23739), .dout(n23741));
  jand g23594(.dina(n18914), .dinb(n2185), .dout(n23742));
  jor  g23595(.dina(n23742), .dinb(n23741), .dout(n23743));
  jor  g23596(.dina(n23743), .dinb(n23738), .dout(n23744));
  jxor g23597(.dina(n23744), .dinb(n2196), .dout(n23745));
  jxor g23598(.dina(n23745), .dinb(n23737), .dout(n23746));
  jxor g23599(.dina(n23746), .dinb(n23662), .dout(n23747));
  jand g23600(.dina(n20371), .dinb(n2743), .dout(n23748));
  jand g23601(.dina(n20205), .dinb(n2752), .dout(n23749));
  jand g23602(.dina(n19922), .dinb(n2748), .dout(n23750));
  jand g23603(.dina(n19373), .dinb(n2757), .dout(n23751));
  jor  g23604(.dina(n23751), .dinb(n23750), .dout(n23752));
  jor  g23605(.dina(n23752), .dinb(n23749), .dout(n23753));
  jor  g23606(.dina(n23753), .dinb(n23748), .dout(n23754));
  jxor g23607(.dina(n23754), .dinb(\a[17] ), .dout(n23755));
  jxor g23608(.dina(n23755), .dinb(n23747), .dout(n23756));
  jxor g23609(.dina(n23756), .dinb(n23657), .dout(n23757));
  jnot g23610(.din(n23757), .dout(n23758));
  jand g23611(.dina(n20949), .dinb(n3423), .dout(n23759));
  jand g23612(.dina(n20344), .dinb(n3428), .dout(n23760));
  jand g23613(.dina(n20947), .dinb(n3569), .dout(n23761));
  jor  g23614(.dina(n23761), .dinb(n23760), .dout(n23762));
  jand g23615(.dina(n20204), .dinb(n3210), .dout(n23763));
  jor  g23616(.dina(n23763), .dinb(n23762), .dout(n23764));
  jor  g23617(.dina(n23764), .dinb(n23759), .dout(n23765));
  jxor g23618(.dina(n23765), .dinb(n3473), .dout(n23766));
  jxor g23619(.dina(n23766), .dinb(n23758), .dout(n23767));
  jxor g23620(.dina(n23767), .dinb(n23654), .dout(n23768));
  jand g23621(.dina(n21342), .dinb(n4022), .dout(n23769));
  jand g23622(.dina(n21340), .dinb(n4220), .dout(n23770));
  jand g23623(.dina(n21197), .dinb(n4027), .dout(n23771));
  jand g23624(.dina(n21198), .dinb(n3870), .dout(n23772));
  jor  g23625(.dina(n23772), .dinb(n23771), .dout(n23773));
  jor  g23626(.dina(n23773), .dinb(n23770), .dout(n23774));
  jor  g23627(.dina(n23774), .dinb(n23769), .dout(n23775));
  jxor g23628(.dina(n23775), .dinb(\a[11] ), .dout(n23776));
  jxor g23629(.dina(n23776), .dinb(n23768), .dout(n23777));
  jxor g23630(.dina(n23777), .dinb(n23650), .dout(n23778));
  jand g23631(.dina(n22279), .dinb(n4691), .dout(n23779));
  jand g23632(.dina(n22163), .dinb(n4941), .dout(n23780));
  jand g23633(.dina(n22164), .dinb(n4696), .dout(n23781));
  jand g23634(.dina(n21974), .dinb(n4701), .dout(n23782));
  jor  g23635(.dina(n23782), .dinb(n23781), .dout(n23783));
  jor  g23636(.dina(n23783), .dinb(n23780), .dout(n23784));
  jor  g23637(.dina(n23784), .dinb(n23779), .dout(n23785));
  jxor g23638(.dina(n23785), .dinb(n4713), .dout(n23786));
  jxor g23639(.dina(n23786), .dinb(n23778), .dout(n23787));
  jnot g23640(.din(n23787), .dout(n23788));
  jxor g23641(.dina(n23788), .dinb(n23645), .dout(n23789));
  jand g23642(.dina(n23172), .dinb(n5280), .dout(n23790));
  jand g23643(.dina(n23080), .dinb(n5814), .dout(n23791));
  jand g23644(.dina(n22937), .dinb(n5531), .dout(n23792));
  jand g23645(.dina(n22265), .dinb(n5536), .dout(n23793));
  jor  g23646(.dina(n23793), .dinb(n23792), .dout(n23794));
  jor  g23647(.dina(n23794), .dinb(n23791), .dout(n23795));
  jor  g23648(.dina(n23795), .dinb(n23790), .dout(n23796));
  jxor g23649(.dina(n23796), .dinb(\a[5] ), .dout(n23797));
  jxor g23650(.dina(n23797), .dinb(n23789), .dout(n23798));
  jnot g23651(.din(n23798), .dout(n23799));
  jxor g23652(.dina(n23799), .dinb(n23638), .dout(n23800));
  jand g23653(.dina(n23144), .dinb(n23079), .dout(n23801));
  jand g23654(.dina(n23145), .dinb(n23091), .dout(n23802));
  jor  g23655(.dina(n23802), .dinb(n23801), .dout(n23803));
  jor  g23656(.dina(n23141), .dinb(n23137), .dout(n23804));
  jor  g23657(.dina(n23143), .dinb(n23095), .dout(n23805));
  jand g23658(.dina(n23805), .dinb(n23804), .dout(n23806));
  jor  g23659(.dina(n23134), .dinb(n23126), .dout(n23807));
  jand g23660(.dina(n23135), .dinb(n23100), .dout(n23808));
  jnot g23661(.din(n23808), .dout(n23809));
  jand g23662(.dina(n23809), .dinb(n23807), .dout(n23810));
  jnot g23663(.din(n23810), .dout(n23811));
  jand g23664(.dina(n23116), .dinb(n23105), .dout(n23812));
  jand g23665(.dina(n23124), .dinb(n23117), .dout(n23813));
  jor  g23666(.dina(n23813), .dinb(n23812), .dout(n23814));
  jand g23667(.dina(n16345), .dinb(n5076), .dout(n23815));
  jand g23668(.dina(n16343), .dinb(n5084), .dout(n23816));
  jand g23669(.dina(n16082), .dinb(n5082), .dout(n23817));
  jor  g23670(.dina(n23121), .dinb(n23817), .dout(n23819));
  jor  g23671(.dina(n23819), .dinb(n23816), .dout(n23820));
  jor  g23672(.dina(n23820), .dinb(n23815), .dout(n23821));
  jor  g23673(.dina(n23111), .dinb(n22981), .dout(n23822));
  jand g23674(.dina(n23115), .dinb(n23112), .dout(n23823));
  jnot g23675(.din(n23823), .dout(n23824));
  jand g23676(.dina(n23824), .dinb(n23822), .dout(n23825));
  jand g23677(.dina(n7996), .dinb(n843), .dout(n23826));
  jand g23678(.dina(n23826), .dinb(n7235), .dout(n23827));
  jand g23679(.dina(n23827), .dinb(n23106), .dout(n23828));
  jnot g23680(.din(n23828), .dout(n23829));
  jxor g23681(.dina(n23829), .dinb(n23825), .dout(n23830));
  jxor g23682(.dina(n23830), .dinb(n23821), .dout(n23831));
  jxor g23683(.dina(n23831), .dinb(n23814), .dout(n23832));
  jnot g23684(.din(n23832), .dout(n23833));
  jxor g23685(.dina(n24287), .dinb(n23833), .dout(n23842));
  jxor g23686(.dina(n23842), .dinb(n23811), .dout(n23843));
  jnot g23687(.din(n23843), .dout(n23844));
  jxor g23688(.dina(n23844), .dinb(n23806), .dout(n23845));
  jxor g23689(.dina(n23845), .dinb(n23144), .dout(n23846));
  jxor g23690(.dina(n23846), .dinb(n23803), .dout(n23847));
  jand g23691(.dina(n23847), .dinb(n6495), .dout(n23848));
  jand g23692(.dina(n23845), .dinb(n6503), .dout(n23849));
  jand g23693(.dina(n23144), .dinb(n6506), .dout(n23850));
  jand g23694(.dina(n23079), .dinb(n6500), .dout(n23851));
  jor  g23695(.dina(n23851), .dinb(n23850), .dout(n23852));
  jor  g23696(.dina(n23852), .dinb(n23849), .dout(n23853));
  jor  g23697(.dina(n23853), .dinb(n23848), .dout(n23854));
  jxor g23698(.dina(n23854), .dinb(n6219), .dout(n23855));
  jxor g23699(.dina(n23855), .dinb(n23800), .dout(n23856));
  jxor g23700(.dina(n23856), .dinb(n23634), .dout(n23857));
  jxor g23701(.dina(n23632), .dinb(n23157), .dout(n23858));
  jxor g23702(.dina(n23858), .dinb(n23857), .dout(\result[0] ));
  jand g23703(.dina(n23858), .dinb(n23857), .dout(n23860));
  jor  g23704(.dina(n23855), .dinb(n23800), .dout(n23861));
  jnot g23705(.din(n23861), .dout(n23862));
  jand g23706(.dina(n23856), .dinb(n23634), .dout(n23863));
  jor  g23707(.dina(n23863), .dinb(n23862), .dout(n23864));
  jnot g23708(.din(n23640), .dout(n23865));
  jand g23709(.dina(n22859), .dinb(n22713), .dout(n23866));
  jor  g23710(.dina(n23866), .dinb(n23865), .dout(n23867));
  jxor g23711(.dina(n23788), .dinb(n23867), .dout(n23868));
  jand g23712(.dina(n23797), .dinb(n23868), .dout(n23869));
  jnot g23713(.din(n23869), .dout(n23870));
  jor  g23714(.dina(n23798), .dinb(n23638), .dout(n23871));
  jand g23715(.dina(n23871), .dinb(n23870), .dout(n23872));
  jnot g23716(.din(n23778), .dout(n23873));
  jor  g23717(.dina(n23786), .dinb(n23873), .dout(n23874));
  jnot g23718(.din(n23874), .dout(n23875));
  jand g23719(.dina(n23788), .dinb(n23867), .dout(n23876));
  jor  g23720(.dina(n23876), .dinb(n23875), .dout(n23877));
  jand g23721(.dina(n23776), .dinb(n23768), .dout(n23878));
  jand g23722(.dina(n23777), .dinb(n23650), .dout(n23879));
  jor  g23723(.dina(n23879), .dinb(n23878), .dout(n23880));
  jor  g23724(.dina(n23766), .dinb(n23758), .dout(n23881));
  jnot g23725(.din(n23881), .dout(n23882));
  jand g23726(.dina(n23767), .dinb(n23654), .dout(n23883));
  jor  g23727(.dina(n23883), .dinb(n23882), .dout(n23884));
  jand g23728(.dina(n23755), .dinb(n23747), .dout(n23885));
  jand g23729(.dina(n23756), .dinb(n23657), .dout(n23886));
  jor  g23730(.dina(n23886), .dinb(n23885), .dout(n23887));
  jor  g23731(.dina(n23745), .dinb(n23737), .dout(n23888));
  jand g23732(.dina(n23746), .dinb(n23662), .dout(n23889));
  jnot g23733(.din(n23889), .dout(n23890));
  jand g23734(.dina(n23890), .dinb(n23888), .dout(n23891));
  jnot g23735(.din(n23891), .dout(n23892));
  jor  g23736(.dina(n23734), .dinb(n23726), .dout(n23893));
  jand g23737(.dina(n23735), .dinb(n23665), .dout(n23894));
  jnot g23738(.din(n23894), .dout(n23895));
  jand g23739(.dina(n23895), .dinb(n23893), .dout(n23896));
  jnot g23740(.din(n23896), .dout(n23897));
  jor  g23741(.dina(n23723), .dinb(n23715), .dout(n23898));
  jand g23742(.dina(n23724), .dinb(n23670), .dout(n23899));
  jnot g23743(.din(n23899), .dout(n23900));
  jand g23744(.dina(n23900), .dinb(n23898), .dout(n23901));
  jnot g23745(.din(n23901), .dout(n23902));
  jor  g23746(.dina(n23712), .dinb(n23704), .dout(n23903));
  jand g23747(.dina(n23713), .dinb(n23675), .dout(n23904));
  jnot g23748(.din(n23904), .dout(n23905));
  jand g23749(.dina(n23905), .dinb(n23903), .dout(n23906));
  jnot g23750(.din(n23906), .dout(n23907));
  jand g23751(.dina(n23701), .dinb(n23694), .dout(n23908));
  jand g23752(.dina(n23702), .dinb(n23678), .dout(n23909));
  jor  g23753(.dina(n23909), .dinb(n23908), .dout(n23910));
  jand g23754(.dina(n18374), .dinb(n1761), .dout(n23911));
  jand g23755(.dina(n1326), .dinb(n175), .dout(n23912));
  jand g23756(.dina(n6151), .dinb(n3276), .dout(n23913));
  jand g23757(.dina(n23913), .dinb(n23912), .dout(n23914));
  jand g23758(.dina(n697), .dinb(n1260), .dout(n23915));
  jand g23759(.dina(n23915), .dinb(n3173), .dout(n23916));
  jand g23760(.dina(n23916), .dinb(n23914), .dout(n23917));
  jand g23761(.dina(n7795), .dinb(n3329), .dout(n23918));
  jand g23762(.dina(n23918), .dinb(n23917), .dout(n23919));
  jand g23763(.dina(n3045), .dinb(n1695), .dout(n23920));
  jand g23764(.dina(n664), .dinb(n495), .dout(n23921));
  jand g23765(.dina(n23921), .dinb(n5463), .dout(n23922));
  jand g23766(.dina(n23922), .dinb(n23920), .dout(n23923));
  jand g23767(.dina(n23923), .dinb(n23919), .dout(n23924));
  jand g23768(.dina(n23924), .dinb(n23911), .dout(n23925));
  jand g23769(.dina(n6005), .dinb(n5347), .dout(n23926));
  jand g23770(.dina(n23926), .dinb(n23925), .dout(n23927));
  jnot g23771(.din(n23927), .dout(n23928));
  jand g23772(.dina(n16606), .dinb(n5076), .dout(n23929));
  jand g23773(.dina(n16604), .dinb(n5084), .dout(n23930));
  jand g23774(.dina(n16360), .dinb(n6050), .dout(n23931));
  jand g23775(.dina(n16355), .dinb(n5082), .dout(n23932));
  jor  g23776(.dina(n23932), .dinb(n23931), .dout(n23933));
  jor  g23777(.dina(n23933), .dinb(n23930), .dout(n23934));
  jor  g23778(.dina(n23934), .dinb(n23929), .dout(n23935));
  jxor g23779(.dina(n23935), .dinb(n23928), .dout(n23936));
  jxor g23780(.dina(n23936), .dinb(n23910), .dout(n23937));
  jnot g23781(.din(n23937), .dout(n23938));
  jand g23782(.dina(n17549), .dinb(n2936), .dout(n23939));
  jand g23783(.dina(n17329), .dinb(n2943), .dout(n23940));
  jand g23784(.dina(n17330), .dinb(n2940), .dout(n23941));
  jand g23785(.dina(n16940), .dinb(n3684), .dout(n23942));
  jor  g23786(.dina(n23942), .dinb(n23941), .dout(n23943));
  jor  g23787(.dina(n23943), .dinb(n23940), .dout(n23944));
  jor  g23788(.dina(n23944), .dinb(n23939), .dout(n23945));
  jxor g23789(.dina(n23945), .dinb(n93), .dout(n23946));
  jxor g23790(.dina(n23946), .dinb(n23938), .dout(n23947));
  jxor g23791(.dina(n23947), .dinb(n23907), .dout(n23948));
  jnot g23792(.din(n23948), .dout(n23949));
  jand g23793(.dina(n18514), .dinb(n71), .dout(n23950));
  jand g23794(.dina(n18293), .dinb(n796), .dout(n23951));
  jand g23795(.dina(n17942), .dinb(n731), .dout(n23952));
  jand g23796(.dina(n17535), .dinb(n1806), .dout(n23953));
  jor  g23797(.dina(n23953), .dinb(n23952), .dout(n23954));
  jor  g23798(.dina(n23954), .dinb(n23951), .dout(n23955));
  jor  g23799(.dina(n23955), .dinb(n23950), .dout(n23956));
  jxor g23800(.dina(n23956), .dinb(n77), .dout(n23957));
  jxor g23801(.dina(n23957), .dinb(n23949), .dout(n23958));
  jxor g23802(.dina(n23958), .dinb(n23902), .dout(n23959));
  jnot g23803(.din(n23959), .dout(n23960));
  jand g23804(.dina(n18916), .dinb(n806), .dout(n23961));
  jand g23805(.dina(n18914), .dinb(n1620), .dout(n23962));
  jand g23806(.dina(n18488), .dinb(n1612), .dout(n23963));
  jand g23807(.dina(n18292), .dinb(n1644), .dout(n23964));
  jor  g23808(.dina(n23964), .dinb(n23963), .dout(n23965));
  jor  g23809(.dina(n23965), .dinb(n23962), .dout(n23966));
  jor  g23810(.dina(n23966), .dinb(n23961), .dout(n23967));
  jxor g23811(.dina(n23967), .dinb(n65), .dout(n23968));
  jxor g23812(.dina(n23968), .dinb(n23960), .dout(n23969));
  jxor g23813(.dina(n23969), .dinb(n23897), .dout(n23970));
  jnot g23814(.din(n23970), .dout(n23971));
  jand g23815(.dina(n19375), .dinb(n1819), .dout(n23972));
  jand g23816(.dina(n19373), .dinb(n2243), .dout(n23973));
  jand g23817(.dina(n19219), .dinb(n2180), .dout(n23974));
  jand g23818(.dina(n19220), .dinb(n2185), .dout(n23975));
  jor  g23819(.dina(n23975), .dinb(n23974), .dout(n23976));
  jor  g23820(.dina(n23976), .dinb(n23973), .dout(n23977));
  jor  g23821(.dina(n23977), .dinb(n23972), .dout(n23978));
  jxor g23822(.dina(n23978), .dinb(n2196), .dout(n23979));
  jxor g23823(.dina(n23979), .dinb(n23971), .dout(n23980));
  jxor g23824(.dina(n23980), .dinb(n23892), .dout(n23981));
  jnot g23825(.din(n23981), .dout(n23982));
  jand g23826(.dina(n20358), .dinb(n2743), .dout(n23983));
  jand g23827(.dina(n20204), .dinb(n2752), .dout(n23984));
  jand g23828(.dina(n20205), .dinb(n2748), .dout(n23985));
  jand g23829(.dina(n19922), .dinb(n2757), .dout(n23986));
  jor  g23830(.dina(n23986), .dinb(n23985), .dout(n23987));
  jor  g23831(.dina(n23987), .dinb(n23984), .dout(n23988));
  jor  g23832(.dina(n23988), .dinb(n23983), .dout(n23989));
  jxor g23833(.dina(n23989), .dinb(n2441), .dout(n23990));
  jxor g23834(.dina(n23990), .dinb(n23982), .dout(n23991));
  jxor g23835(.dina(n23991), .dinb(n23887), .dout(n23992));
  jnot g23836(.din(n23992), .dout(n23993));
  jand g23837(.dina(n21367), .dinb(n3423), .dout(n23994));
  jand g23838(.dina(n21198), .dinb(n3569), .dout(n23995));
  jand g23839(.dina(n20947), .dinb(n3428), .dout(n23996));
  jand g23840(.dina(n20344), .dinb(n3210), .dout(n23997));
  jor  g23841(.dina(n23997), .dinb(n23996), .dout(n23998));
  jor  g23842(.dina(n23998), .dinb(n23995), .dout(n23999));
  jor  g23843(.dina(n23999), .dinb(n23994), .dout(n24000));
  jxor g23844(.dina(n24000), .dinb(n3473), .dout(n24001));
  jxor g23845(.dina(n24001), .dinb(n23993), .dout(n24002));
  jxor g23846(.dina(n24002), .dinb(n23884), .dout(n24003));
  jand g23847(.dina(n21976), .dinb(n4022), .dout(n24004));
  jand g23848(.dina(n21974), .dinb(n4220), .dout(n24005));
  jand g23849(.dina(n21340), .dinb(n4027), .dout(n24006));
  jand g23850(.dina(n21197), .dinb(n3870), .dout(n24007));
  jor  g23851(.dina(n24007), .dinb(n24006), .dout(n24008));
  jor  g23852(.dina(n24008), .dinb(n24005), .dout(n24009));
  jor  g23853(.dina(n24009), .dinb(n24004), .dout(n24010));
  jxor g23854(.dina(n24010), .dinb(n4050), .dout(n24011));
  jxor g23855(.dina(n24011), .dinb(n24003), .dout(n24012));
  jnot g23856(.din(n24012), .dout(n24013));
  jxor g23857(.dina(n24013), .dinb(n23880), .dout(n24014));
  jand g23858(.dina(n22267), .dinb(n4691), .dout(n24015));
  jand g23859(.dina(n22163), .dinb(n4696), .dout(n24016));
  jand g23860(.dina(n22265), .dinb(n4941), .dout(n24017));
  jor  g23861(.dina(n24017), .dinb(n24016), .dout(n24018));
  jand g23862(.dina(n22164), .dinb(n4701), .dout(n24019));
  jor  g23863(.dina(n24019), .dinb(n24018), .dout(n24020));
  jor  g23864(.dina(n24020), .dinb(n24015), .dout(n24021));
  jxor g23865(.dina(n24021), .dinb(n4713), .dout(n24022));
  jxor g23866(.dina(n24022), .dinb(n24014), .dout(n24023));
  jnot g23867(.din(n24023), .dout(n24024));
  jxor g23868(.dina(n24024), .dinb(n23877), .dout(n24025));
  jand g23869(.dina(n23159), .dinb(n5280), .dout(n24026));
  jand g23870(.dina(n23079), .dinb(n5814), .dout(n24027));
  jand g23871(.dina(n23080), .dinb(n5531), .dout(n24028));
  jand g23872(.dina(n22937), .dinb(n5536), .dout(n24029));
  jor  g23873(.dina(n24029), .dinb(n24028), .dout(n24030));
  jor  g23874(.dina(n24030), .dinb(n24027), .dout(n24031));
  jor  g23875(.dina(n24031), .dinb(n24026), .dout(n24032));
  jxor g23876(.dina(n24032), .dinb(n5277), .dout(n24033));
  jxor g23877(.dina(n24033), .dinb(n24025), .dout(n24034));
  jnot g23878(.din(n24034), .dout(n24035));
  jxor g23879(.dina(n24035), .dinb(n23872), .dout(n24036));
  jand g23880(.dina(n23845), .dinb(n23144), .dout(n24037));
  jand g23881(.dina(n23846), .dinb(n23803), .dout(n24038));
  jor  g23882(.dina(n24038), .dinb(n24037), .dout(n24039));
  jand g23883(.dina(n23842), .dinb(n23811), .dout(n24040));
  jnot g23884(.din(n24040), .dout(n24041));
  jor  g23885(.dina(n23844), .dinb(n23806), .dout(n24042));
  jand g23886(.dina(n24042), .dinb(n24041), .dout(n24043));
  jand g23887(.dina(n23831), .dinb(n23814), .dout(n24044));
  jnot g23888(.din(n24044), .dout(n24045));
  jor  g23889(.dina(n24287), .dinb(n23833), .dout(n24046));
  jand g23890(.dina(n24046), .dinb(n24045), .dout(n24047));
  jnot g23891(.din(n24047), .dout(n24048));
  jand g23892(.dina(n16594), .dinb(n5076), .dout(n24049));
  jand g23893(.dina(n16592), .dinb(n5084), .dout(n24050));
  jand g23894(.dina(n16343), .dinb(n5082), .dout(n24051));
  jand g23895(.dina(n16082), .dinb(n6050), .dout(n24052));
  jor  g23896(.dina(n24052), .dinb(n24051), .dout(n24053));
  jor  g23897(.dina(n24053), .dinb(n24050), .dout(n24054));
  jor  g23898(.dina(n24054), .dinb(n24049), .dout(n24055));
  jnot g23899(.din(n24055), .dout(n24056));
  jxor g23900(.dina(n24287), .dinb(n24056), .dout(n24064));
  jnot g23901(.din(n23825), .dout(n24065));
  jand g23902(.dina(n23828), .dinb(n24065), .dout(n24066));
  jand g23903(.dina(n23830), .dinb(n23821), .dout(n24067));
  jor  g23904(.dina(n24067), .dinb(n24066), .dout(n24068));
  jand g23905(.dina(n7998), .dinb(n7647), .dout(n24069));
  jxor g23906(.dina(n24069), .dinb(n23829), .dout(n24070));
  jxor g23907(.dina(n24070), .dinb(n24068), .dout(n24071));
  jxor g23908(.dina(n24071), .dinb(n24064), .dout(n24072));
  jxor g23909(.dina(n24072), .dinb(n24048), .dout(n24073));
  jnot g23910(.din(n24073), .dout(n24074));
  jxor g23911(.dina(n24074), .dinb(n24043), .dout(n24075));
  jxor g23912(.dina(n24075), .dinb(n23845), .dout(n24076));
  jxor g23913(.dina(n24076), .dinb(n24039), .dout(n24077));
  jand g23914(.dina(n24077), .dinb(n6495), .dout(n24078));
  jand g23915(.dina(n24075), .dinb(n6503), .dout(n24079));
  jand g23916(.dina(n23845), .dinb(n6506), .dout(n24080));
  jand g23917(.dina(n23144), .dinb(n6500), .dout(n24081));
  jor  g23918(.dina(n24081), .dinb(n24080), .dout(n24082));
  jor  g23919(.dina(n24082), .dinb(n24079), .dout(n24083));
  jor  g23920(.dina(n24083), .dinb(n24078), .dout(n24084));
  jxor g23921(.dina(n24084), .dinb(n6219), .dout(n24085));
  jxor g23922(.dina(n24085), .dinb(n24036), .dout(n24086));
  jxor g23923(.dina(n24086), .dinb(n23864), .dout(n24087));
  jxor g23924(.dina(n24087), .dinb(n23860), .dout(\result[1] ));
  jand g23925(.dina(n24087), .dinb(n23860), .dout(n24089));
  jor  g23926(.dina(n24085), .dinb(n24036), .dout(n24090));
  jnot g23927(.din(n24090), .dout(n24091));
  jand g23928(.dina(n24086), .dinb(n23864), .dout(n24092));
  jor  g23929(.dina(n24092), .dinb(n24091), .dout(n24093));
  jnot g23930(.din(n24025), .dout(n24094));
  jor  g23931(.dina(n24033), .dinb(n24094), .dout(n24095));
  jor  g23932(.dina(n24034), .dinb(n23872), .dout(n24096));
  jand g23933(.dina(n24096), .dinb(n24095), .dout(n24097));
  jnot g23934(.din(n24014), .dout(n24098));
  jor  g23935(.dina(n24022), .dinb(n24098), .dout(n24099));
  jnot g23936(.din(n24099), .dout(n24100));
  jand g23937(.dina(n24024), .dinb(n23877), .dout(n24101));
  jor  g23938(.dina(n24101), .dinb(n24100), .dout(n24102));
  jnot g23939(.din(n24003), .dout(n24103));
  jor  g23940(.dina(n24011), .dinb(n24103), .dout(n24104));
  jnot g23941(.din(n24104), .dout(n24105));
  jand g23942(.dina(n24013), .dinb(n23880), .dout(n24106));
  jor  g23943(.dina(n24106), .dinb(n24105), .dout(n24107));
  jor  g23944(.dina(n24001), .dinb(n23993), .dout(n24108));
  jnot g23945(.din(n24108), .dout(n24109));
  jand g23946(.dina(n24002), .dinb(n23884), .dout(n24110));
  jor  g23947(.dina(n24110), .dinb(n24109), .dout(n24111));
  jor  g23948(.dina(n23990), .dinb(n23982), .dout(n24112));
  jand g23949(.dina(n23991), .dinb(n23887), .dout(n24113));
  jnot g23950(.din(n24113), .dout(n24114));
  jand g23951(.dina(n24114), .dinb(n24112), .dout(n24115));
  jnot g23952(.din(n24115), .dout(n24116));
  jor  g23953(.dina(n23979), .dinb(n23971), .dout(n24117));
  jand g23954(.dina(n23980), .dinb(n23892), .dout(n24118));
  jnot g23955(.din(n24118), .dout(n24119));
  jand g23956(.dina(n24119), .dinb(n24117), .dout(n24120));
  jnot g23957(.din(n24120), .dout(n24121));
  jor  g23958(.dina(n23968), .dinb(n23960), .dout(n24122));
  jand g23959(.dina(n23969), .dinb(n23897), .dout(n24123));
  jnot g23960(.din(n24123), .dout(n24124));
  jand g23961(.dina(n24124), .dinb(n24122), .dout(n24125));
  jnot g23962(.din(n24125), .dout(n24126));
  jor  g23963(.dina(n23957), .dinb(n23949), .dout(n24127));
  jand g23964(.dina(n23958), .dinb(n23902), .dout(n24128));
  jnot g23965(.din(n24128), .dout(n24129));
  jand g23966(.dina(n24129), .dinb(n24127), .dout(n24130));
  jnot g23967(.din(n24130), .dout(n24131));
  jor  g23968(.dina(n23946), .dinb(n23938), .dout(n24132));
  jand g23969(.dina(n23947), .dinb(n23907), .dout(n24133));
  jnot g23970(.din(n24133), .dout(n24134));
  jand g23971(.dina(n24134), .dinb(n24132), .dout(n24135));
  jnot g23972(.din(n24135), .dout(n24136));
  jand g23973(.dina(n23935), .dinb(n23928), .dout(n24137));
  jand g23974(.dina(n23936), .dinb(n23910), .dout(n24138));
  jor  g23975(.dina(n24138), .dinb(n24137), .dout(n24139));
  jand g23976(.dina(n3762), .dinb(n3176), .dout(n24140));
  jand g23977(.dina(n24140), .dinb(n1485), .dout(n24141));
  jand g23978(.dina(n3397), .dinb(n447), .dout(n24142));
  jand g23979(.dina(n24142), .dinb(n1324), .dout(n24143));
  jand g23980(.dina(n24143), .dinb(n24141), .dout(n24144));
  jand g23981(.dina(n461), .dinb(n450), .dout(n24145));
  jand g23982(.dina(n24145), .dinb(n7666), .dout(n24146));
  jand g23983(.dina(n24146), .dinb(n17799), .dout(n24147));
  jand g23984(.dina(n24147), .dinb(n7096), .dout(n24148));
  jand g23985(.dina(n24148), .dinb(n24144), .dout(n24149));
  jand g23986(.dina(n24149), .dinb(n3006), .dout(n24150));
  jand g23987(.dina(n24150), .dinb(n2594), .dout(n24151));
  jand g23988(.dina(n18977), .dinb(n1230), .dout(n24152));
  jand g23989(.dina(n24152), .dinb(n9729), .dout(n24153));
  jand g23990(.dina(n24153), .dinb(n13191), .dout(n24154));
  jand g23991(.dina(n24154), .dinb(n24151), .dout(n24155));
  jnot g23992(.din(n24155), .dout(n24156));
  jand g23993(.dina(n16942), .dinb(n5076), .dout(n24157));
  jand g23994(.dina(n16940), .dinb(n5084), .dout(n24158));
  jand g23995(.dina(n16355), .dinb(n6050), .dout(n24159));
  jand g23996(.dina(n16604), .dinb(n5082), .dout(n24160));
  jor  g23997(.dina(n24160), .dinb(n24159), .dout(n24161));
  jor  g23998(.dina(n24161), .dinb(n24158), .dout(n24162));
  jor  g23999(.dina(n24162), .dinb(n24157), .dout(n24163));
  jxor g24000(.dina(n24163), .dinb(n24156), .dout(n24164));
  jxor g24001(.dina(n24164), .dinb(n24139), .dout(n24165));
  jnot g24002(.din(n24165), .dout(n24166));
  jand g24003(.dina(n17537), .dinb(n2936), .dout(n24167));
  jand g24004(.dina(n17535), .dinb(n2943), .dout(n24168));
  jand g24005(.dina(n17329), .dinb(n2940), .dout(n24169));
  jand g24006(.dina(n17330), .dinb(n3684), .dout(n24170));
  jor  g24007(.dina(n24170), .dinb(n24169), .dout(n24171));
  jor  g24008(.dina(n24171), .dinb(n24168), .dout(n24172));
  jor  g24009(.dina(n24172), .dinb(n24167), .dout(n24173));
  jxor g24010(.dina(n24173), .dinb(n93), .dout(n24174));
  jxor g24011(.dina(n24174), .dinb(n24166), .dout(n24175));
  jxor g24012(.dina(n24175), .dinb(n24136), .dout(n24176));
  jnot g24013(.din(n24176), .dout(n24177));
  jand g24014(.dina(n18502), .dinb(n71), .dout(n24178));
  jand g24015(.dina(n18293), .dinb(n731), .dout(n24179));
  jand g24016(.dina(n18292), .dinb(n796), .dout(n24180));
  jor  g24017(.dina(n24180), .dinb(n24179), .dout(n24181));
  jand g24018(.dina(n17942), .dinb(n1806), .dout(n24182));
  jor  g24019(.dina(n24182), .dinb(n24181), .dout(n24183));
  jor  g24020(.dina(n24183), .dinb(n24178), .dout(n24184));
  jxor g24021(.dina(n24184), .dinb(n77), .dout(n24185));
  jxor g24022(.dina(n24185), .dinb(n24177), .dout(n24186));
  jxor g24023(.dina(n24186), .dinb(n24131), .dout(n24187));
  jnot g24024(.din(n24187), .dout(n24188));
  jand g24025(.dina(n19399), .dinb(n806), .dout(n24189));
  jand g24026(.dina(n18914), .dinb(n1612), .dout(n24190));
  jand g24027(.dina(n19220), .dinb(n1620), .dout(n24191));
  jor  g24028(.dina(n24191), .dinb(n24190), .dout(n24192));
  jand g24029(.dina(n18488), .dinb(n1644), .dout(n24193));
  jor  g24030(.dina(n24193), .dinb(n24192), .dout(n24194));
  jor  g24031(.dina(n24194), .dinb(n24189), .dout(n24195));
  jxor g24032(.dina(n24195), .dinb(n65), .dout(n24196));
  jxor g24033(.dina(n24196), .dinb(n24188), .dout(n24197));
  jxor g24034(.dina(n24197), .dinb(n24126), .dout(n24198));
  jnot g24035(.din(n24198), .dout(n24199));
  jand g24036(.dina(n19924), .dinb(n1819), .dout(n24200));
  jand g24037(.dina(n19922), .dinb(n2243), .dout(n24201));
  jand g24038(.dina(n19373), .dinb(n2180), .dout(n24202));
  jand g24039(.dina(n19219), .dinb(n2185), .dout(n24203));
  jor  g24040(.dina(n24203), .dinb(n24202), .dout(n24204));
  jor  g24041(.dina(n24204), .dinb(n24201), .dout(n24205));
  jor  g24042(.dina(n24205), .dinb(n24200), .dout(n24206));
  jxor g24043(.dina(n24206), .dinb(n2196), .dout(n24207));
  jxor g24044(.dina(n24207), .dinb(n24199), .dout(n24208));
  jxor g24045(.dina(n24208), .dinb(n24121), .dout(n24209));
  jnot g24046(.din(n24209), .dout(n24210));
  jand g24047(.dina(n20346), .dinb(n2743), .dout(n24211));
  jand g24048(.dina(n20344), .dinb(n2752), .dout(n24212));
  jand g24049(.dina(n20204), .dinb(n2748), .dout(n24213));
  jand g24050(.dina(n20205), .dinb(n2757), .dout(n24214));
  jor  g24051(.dina(n24214), .dinb(n24213), .dout(n24215));
  jor  g24052(.dina(n24215), .dinb(n24212), .dout(n24216));
  jor  g24053(.dina(n24216), .dinb(n24211), .dout(n24217));
  jxor g24054(.dina(n24217), .dinb(n2441), .dout(n24218));
  jxor g24055(.dina(n24218), .dinb(n24210), .dout(n24219));
  jxor g24056(.dina(n24219), .dinb(n24116), .dout(n24220));
  jnot g24057(.din(n24220), .dout(n24221));
  jand g24058(.dina(n21355), .dinb(n3423), .dout(n24222));
  jand g24059(.dina(n21197), .dinb(n3569), .dout(n24223));
  jand g24060(.dina(n21198), .dinb(n3428), .dout(n24224));
  jand g24061(.dina(n20947), .dinb(n3210), .dout(n24225));
  jor  g24062(.dina(n24225), .dinb(n24224), .dout(n24226));
  jor  g24063(.dina(n24226), .dinb(n24223), .dout(n24227));
  jor  g24064(.dina(n24227), .dinb(n24222), .dout(n24228));
  jxor g24065(.dina(n24228), .dinb(n3473), .dout(n24229));
  jxor g24066(.dina(n24229), .dinb(n24221), .dout(n24230));
  jxor g24067(.dina(n24230), .dinb(n24111), .dout(n24231));
  jand g24068(.dina(n22291), .dinb(n4022), .dout(n24232));
  jand g24069(.dina(n22164), .dinb(n4220), .dout(n24233));
  jand g24070(.dina(n21974), .dinb(n4027), .dout(n24234));
  jand g24071(.dina(n21340), .dinb(n3870), .dout(n24235));
  jor  g24072(.dina(n24235), .dinb(n24234), .dout(n24236));
  jor  g24073(.dina(n24236), .dinb(n24233), .dout(n24237));
  jor  g24074(.dina(n24237), .dinb(n24232), .dout(n24238));
  jxor g24075(.dina(n24238), .dinb(n4050), .dout(n24239));
  jxor g24076(.dina(n24239), .dinb(n24231), .dout(n24240));
  jnot g24077(.din(n24240), .dout(n24241));
  jxor g24078(.dina(n24241), .dinb(n24107), .dout(n24242));
  jand g24079(.dina(n22939), .dinb(n4691), .dout(n24243));
  jand g24080(.dina(n22265), .dinb(n4696), .dout(n24244));
  jand g24081(.dina(n22937), .dinb(n4941), .dout(n24245));
  jor  g24082(.dina(n24245), .dinb(n24244), .dout(n24246));
  jand g24083(.dina(n22163), .dinb(n4701), .dout(n24247));
  jor  g24084(.dina(n24247), .dinb(n24246), .dout(n24248));
  jor  g24085(.dina(n24248), .dinb(n24243), .dout(n24249));
  jxor g24086(.dina(n24249), .dinb(n4713), .dout(n24250));
  jxor g24087(.dina(n24250), .dinb(n24242), .dout(n24251));
  jnot g24088(.din(n24251), .dout(n24252));
  jxor g24089(.dina(n24252), .dinb(n24102), .dout(n24253));
  jand g24090(.dina(n23146), .dinb(n5280), .dout(n24254));
  jand g24091(.dina(n23079), .dinb(n5531), .dout(n24255));
  jand g24092(.dina(n23144), .dinb(n5814), .dout(n24256));
  jor  g24093(.dina(n24256), .dinb(n24255), .dout(n24257));
  jand g24094(.dina(n23080), .dinb(n5536), .dout(n24258));
  jor  g24095(.dina(n24258), .dinb(n24257), .dout(n24259));
  jor  g24096(.dina(n24259), .dinb(n24254), .dout(n24260));
  jxor g24097(.dina(n24260), .dinb(n5277), .dout(n24261));
  jxor g24098(.dina(n24261), .dinb(n24253), .dout(n24262));
  jnot g24099(.din(n24262), .dout(n24263));
  jxor g24100(.dina(n24263), .dinb(n24097), .dout(n24264));
  jnot g24101(.din(n23845), .dout(n24265));
  jnot g24102(.din(n24075), .dout(n24266));
  jor  g24103(.dina(n24266), .dinb(n24265), .dout(n24267));
  jnot g24104(.din(n24039), .dout(n24268));
  jnot g24105(.din(n24076), .dout(n24269));
  jor  g24106(.dina(n24269), .dinb(n24268), .dout(n24270));
  jand g24107(.dina(n24270), .dinb(n24267), .dout(n24271));
  jand g24108(.dina(n24072), .dinb(n24048), .dout(n24272));
  jnot g24109(.din(n24272), .dout(n24273));
  jor  g24110(.dina(n24074), .dinb(n24043), .dout(n24274));
  jand g24111(.dina(n24274), .dinb(n24273), .dout(n24275));
  jor  g24112(.dina(n24287), .dinb(n24056), .dout(n24276));
  jand g24113(.dina(n24071), .dinb(n24064), .dout(n24277));
  jnot g24114(.din(n24277), .dout(n24278));
  jand g24115(.dina(n24278), .dinb(n24276), .dout(n24279));
  jnot g24116(.din(n24279), .dout(n24280));
  jand g24117(.dina(n24069), .dinb(n23829), .dout(n24281));
  jand g24118(.dina(n24070), .dinb(n24068), .dout(n24282));
  jor  g24119(.dina(n24282), .dinb(n24281), .dout(n24283));
  jxor g24120(.dina(n24069), .dinb(n24501), .dout(n24284));
  jor  g24121(.dina(n3682), .dinb(n2935), .dout(n24285));
  jand g24122(.dina(n24285), .dinb(n16924), .dout(n24286));
  jxor g24123(.dina(n24286), .dinb(n93), .dout(n24287));
  jxor g24124(.dina(n24287), .dinb(n24284), .dout(n24288));
  jand g24125(.dina(n16930), .dinb(n5076), .dout(n24289));
  jand g24126(.dina(n16592), .dinb(n5082), .dout(n24290));
  jand g24127(.dina(n16928), .dinb(n5084), .dout(n24291));
  jor  g24128(.dina(n6050), .dinb(n24291), .dout(n24293));
  jor  g24129(.dina(n24293), .dinb(n24290), .dout(n24294));
  jor  g24130(.dina(n24294), .dinb(n24289), .dout(n24295));
  jxor g24131(.dina(n24295), .dinb(n24288), .dout(n24296));
  jxor g24132(.dina(n24296), .dinb(n24283), .dout(n24297));
  jxor g24133(.dina(n24297), .dinb(n24280), .dout(n24298));
  jnot g24134(.din(n24298), .dout(n24299));
  jxor g24135(.dina(n24299), .dinb(n24275), .dout(n24300));
  jxor g24136(.dina(n24300), .dinb(n24075), .dout(n24301));
  jxor g24137(.dina(n24301), .dinb(n24271), .dout(n24302));
  jor  g24138(.dina(n24302), .dinb(n6496), .dout(n24303));
  jnot g24139(.din(n24300), .dout(n24304));
  jor  g24140(.dina(n24304), .dinb(n6504), .dout(n24305));
  jor  g24141(.dina(n24266), .dinb(n6507), .dout(n24306));
  jor  g24142(.dina(n24265), .dinb(n6501), .dout(n24307));
  jand g24143(.dina(n24307), .dinb(n24306), .dout(n24308));
  jand g24144(.dina(n24308), .dinb(n24305), .dout(n24309));
  jand g24145(.dina(n24309), .dinb(n24303), .dout(n24310));
  jxor g24146(.dina(n24310), .dinb(\a[2] ), .dout(n24311));
  jxor g24147(.dina(n24311), .dinb(n24264), .dout(n24312));
  jxor g24148(.dina(n24312), .dinb(n24093), .dout(n24313));
  jxor g24149(.dina(n24313), .dinb(n24089), .dout(\result[2] ));
  jand g24150(.dina(n24313), .dinb(n24089), .dout(n24315));
  jor  g24151(.dina(n24311), .dinb(n24264), .dout(n24316));
  jnot g24152(.din(n24316), .dout(n24317));
  jand g24153(.dina(n24312), .dinb(n24093), .dout(n24318));
  jor  g24154(.dina(n24318), .dinb(n24317), .dout(n24319));
  jnot g24155(.din(n24253), .dout(n24320));
  jor  g24156(.dina(n24261), .dinb(n24320), .dout(n24321));
  jor  g24157(.dina(n24262), .dinb(n24097), .dout(n24322));
  jand g24158(.dina(n24322), .dinb(n24321), .dout(n24323));
  jnot g24159(.din(n24242), .dout(n24324));
  jor  g24160(.dina(n24250), .dinb(n24324), .dout(n24325));
  jnot g24161(.din(n24325), .dout(n24326));
  jand g24162(.dina(n24252), .dinb(n24102), .dout(n24327));
  jor  g24163(.dina(n24327), .dinb(n24326), .dout(n24328));
  jnot g24164(.din(n24231), .dout(n24329));
  jor  g24165(.dina(n24239), .dinb(n24329), .dout(n24330));
  jand g24166(.dina(n24241), .dinb(n24107), .dout(n24331));
  jnot g24167(.din(n24331), .dout(n24332));
  jand g24168(.dina(n24332), .dinb(n24330), .dout(n24333));
  jor  g24169(.dina(n24229), .dinb(n24221), .dout(n24334));
  jnot g24170(.din(n24334), .dout(n24335));
  jand g24171(.dina(n24230), .dinb(n24111), .dout(n24336));
  jor  g24172(.dina(n24336), .dinb(n24335), .dout(n24337));
  jor  g24173(.dina(n24218), .dinb(n24210), .dout(n24338));
  jand g24174(.dina(n24219), .dinb(n24116), .dout(n24339));
  jnot g24175(.din(n24339), .dout(n24340));
  jand g24176(.dina(n24340), .dinb(n24338), .dout(n24341));
  jnot g24177(.din(n24341), .dout(n24342));
  jor  g24178(.dina(n24207), .dinb(n24199), .dout(n24343));
  jand g24179(.dina(n24208), .dinb(n24121), .dout(n24344));
  jnot g24180(.din(n24344), .dout(n24345));
  jand g24181(.dina(n24345), .dinb(n24343), .dout(n24346));
  jnot g24182(.din(n24346), .dout(n24347));
  jor  g24183(.dina(n24196), .dinb(n24188), .dout(n24348));
  jand g24184(.dina(n24197), .dinb(n24126), .dout(n24349));
  jnot g24185(.din(n24349), .dout(n24350));
  jand g24186(.dina(n24350), .dinb(n24348), .dout(n24351));
  jnot g24187(.din(n24351), .dout(n24352));
  jor  g24188(.dina(n24185), .dinb(n24177), .dout(n24353));
  jand g24189(.dina(n24186), .dinb(n24131), .dout(n24354));
  jnot g24190(.din(n24354), .dout(n24355));
  jand g24191(.dina(n24355), .dinb(n24353), .dout(n24356));
  jnot g24192(.din(n24356), .dout(n24357));
  jor  g24193(.dina(n24174), .dinb(n24166), .dout(n24358));
  jand g24194(.dina(n24175), .dinb(n24136), .dout(n24359));
  jnot g24195(.din(n24359), .dout(n24360));
  jand g24196(.dina(n24360), .dinb(n24358), .dout(n24361));
  jnot g24197(.din(n24361), .dout(n24362));
  jand g24198(.dina(n24163), .dinb(n24156), .dout(n24363));
  jand g24199(.dina(n24164), .dinb(n24139), .dout(n24364));
  jor  g24200(.dina(n24364), .dinb(n24363), .dout(n24365));
  jand g24201(.dina(n1462), .dinb(n1438), .dout(n24366));
  jand g24202(.dina(n24366), .dinb(n5351), .dout(n24367));
  jand g24203(.dina(n24367), .dinb(n704), .dout(n24368));
  jand g24204(.dina(n1851), .dinb(n1485), .dout(n24369));
  jand g24205(.dina(n24369), .dinb(n1207), .dout(n24370));
  jand g24206(.dina(n24370), .dinb(n2993), .dout(n24371));
  jand g24207(.dina(n24371), .dinb(n24368), .dout(n24372));
  jand g24208(.dina(n3146), .dinb(n121), .dout(n24373));
  jand g24209(.dina(n24373), .dinb(n11401), .dout(n24374));
  jand g24210(.dina(n24374), .dinb(n3175), .dout(n24375));
  jand g24211(.dina(n24375), .dinb(n24372), .dout(n24376));
  jand g24212(.dina(n17169), .dinb(n1939), .dout(n24377));
  jand g24213(.dina(n24377), .dinb(n24376), .dout(n24378));
  jand g24214(.dina(n24378), .dinb(n7099), .dout(n24379));
  jand g24215(.dina(n24379), .dinb(n6028), .dout(n24380));
  jnot g24216(.din(n24380), .dout(n24381));
  jand g24217(.dina(n17561), .dinb(n5076), .dout(n24382));
  jand g24218(.dina(n17330), .dinb(n5084), .dout(n24383));
  jand g24219(.dina(n16604), .dinb(n6050), .dout(n24384));
  jand g24220(.dina(n16940), .dinb(n5082), .dout(n24385));
  jor  g24221(.dina(n24385), .dinb(n24384), .dout(n24386));
  jor  g24222(.dina(n24386), .dinb(n24383), .dout(n24387));
  jor  g24223(.dina(n24387), .dinb(n24382), .dout(n24388));
  jxor g24224(.dina(n24388), .dinb(n24381), .dout(n24389));
  jxor g24225(.dina(n24389), .dinb(n24365), .dout(n24390));
  jnot g24226(.din(n24390), .dout(n24391));
  jand g24227(.dina(n17944), .dinb(n2936), .dout(n24392));
  jand g24228(.dina(n17942), .dinb(n2943), .dout(n24393));
  jand g24229(.dina(n17535), .dinb(n2940), .dout(n24394));
  jand g24230(.dina(n17329), .dinb(n3684), .dout(n24395));
  jor  g24231(.dina(n24395), .dinb(n24394), .dout(n24396));
  jor  g24232(.dina(n24396), .dinb(n24393), .dout(n24397));
  jor  g24233(.dina(n24397), .dinb(n24392), .dout(n24398));
  jxor g24234(.dina(n24398), .dinb(n93), .dout(n24399));
  jxor g24235(.dina(n24399), .dinb(n24391), .dout(n24400));
  jxor g24236(.dina(n24400), .dinb(n24362), .dout(n24401));
  jnot g24237(.din(n24401), .dout(n24402));
  jand g24238(.dina(n18490), .dinb(n71), .dout(n24403));
  jand g24239(.dina(n18488), .dinb(n796), .dout(n24404));
  jand g24240(.dina(n18292), .dinb(n731), .dout(n24405));
  jand g24241(.dina(n18293), .dinb(n1806), .dout(n24406));
  jor  g24242(.dina(n24406), .dinb(n24405), .dout(n24407));
  jor  g24243(.dina(n24407), .dinb(n24404), .dout(n24408));
  jor  g24244(.dina(n24408), .dinb(n24403), .dout(n24409));
  jxor g24245(.dina(n24409), .dinb(n77), .dout(n24410));
  jxor g24246(.dina(n24410), .dinb(n24402), .dout(n24411));
  jxor g24247(.dina(n24411), .dinb(n24357), .dout(n24412));
  jnot g24248(.din(n24412), .dout(n24413));
  jand g24249(.dina(n19387), .dinb(n806), .dout(n24414));
  jand g24250(.dina(n19220), .dinb(n1612), .dout(n24415));
  jand g24251(.dina(n19219), .dinb(n1620), .dout(n24416));
  jor  g24252(.dina(n24416), .dinb(n24415), .dout(n24417));
  jand g24253(.dina(n18914), .dinb(n1644), .dout(n24418));
  jor  g24254(.dina(n24418), .dinb(n24417), .dout(n24419));
  jor  g24255(.dina(n24419), .dinb(n24414), .dout(n24420));
  jxor g24256(.dina(n24420), .dinb(n65), .dout(n24421));
  jxor g24257(.dina(n24421), .dinb(n24413), .dout(n24422));
  jxor g24258(.dina(n24422), .dinb(n24352), .dout(n24423));
  jnot g24259(.din(n24423), .dout(n24424));
  jand g24260(.dina(n20371), .dinb(n1819), .dout(n24425));
  jand g24261(.dina(n20205), .dinb(n2243), .dout(n24426));
  jand g24262(.dina(n19922), .dinb(n2180), .dout(n24427));
  jand g24263(.dina(n19373), .dinb(n2185), .dout(n24428));
  jor  g24264(.dina(n24428), .dinb(n24427), .dout(n24429));
  jor  g24265(.dina(n24429), .dinb(n24426), .dout(n24430));
  jor  g24266(.dina(n24430), .dinb(n24425), .dout(n24431));
  jxor g24267(.dina(n24431), .dinb(n2196), .dout(n24432));
  jxor g24268(.dina(n24432), .dinb(n24424), .dout(n24433));
  jxor g24269(.dina(n24433), .dinb(n24347), .dout(n24434));
  jand g24270(.dina(n20949), .dinb(n2743), .dout(n24435));
  jand g24271(.dina(n20947), .dinb(n2752), .dout(n24436));
  jand g24272(.dina(n20344), .dinb(n2748), .dout(n24437));
  jand g24273(.dina(n20204), .dinb(n2757), .dout(n24438));
  jor  g24274(.dina(n24438), .dinb(n24437), .dout(n24439));
  jor  g24275(.dina(n24439), .dinb(n24436), .dout(n24440));
  jor  g24276(.dina(n24440), .dinb(n24435), .dout(n24441));
  jxor g24277(.dina(n24441), .dinb(\a[17] ), .dout(n24442));
  jxor g24278(.dina(n24442), .dinb(n24434), .dout(n24443));
  jxor g24279(.dina(n24443), .dinb(n24342), .dout(n24444));
  jand g24280(.dina(n21342), .dinb(n3423), .dout(n24445));
  jand g24281(.dina(n21340), .dinb(n3569), .dout(n24446));
  jand g24282(.dina(n21197), .dinb(n3428), .dout(n24447));
  jand g24283(.dina(n21198), .dinb(n3210), .dout(n24448));
  jor  g24284(.dina(n24448), .dinb(n24447), .dout(n24449));
  jor  g24285(.dina(n24449), .dinb(n24446), .dout(n24450));
  jor  g24286(.dina(n24450), .dinb(n24445), .dout(n24451));
  jxor g24287(.dina(n24451), .dinb(n3473), .dout(n24452));
  jxor g24288(.dina(n24452), .dinb(n24444), .dout(n24453));
  jxor g24289(.dina(n24453), .dinb(n24337), .dout(n24454));
  jand g24290(.dina(n22279), .dinb(n4022), .dout(n24455));
  jand g24291(.dina(n22164), .dinb(n4027), .dout(n24456));
  jand g24292(.dina(n22163), .dinb(n4220), .dout(n24457));
  jor  g24293(.dina(n24457), .dinb(n24456), .dout(n24458));
  jand g24294(.dina(n21974), .dinb(n3870), .dout(n24459));
  jor  g24295(.dina(n24459), .dinb(n24458), .dout(n24460));
  jor  g24296(.dina(n24460), .dinb(n24455), .dout(n24461));
  jxor g24297(.dina(n24461), .dinb(n4050), .dout(n24462));
  jxor g24298(.dina(n24462), .dinb(n24454), .dout(n24463));
  jxor g24299(.dina(n24463), .dinb(n24333), .dout(n24464));
  jand g24300(.dina(n23172), .dinb(n4691), .dout(n24465));
  jand g24301(.dina(n23080), .dinb(n4941), .dout(n24466));
  jand g24302(.dina(n22937), .dinb(n4696), .dout(n24467));
  jand g24303(.dina(n22265), .dinb(n4701), .dout(n24468));
  jor  g24304(.dina(n24468), .dinb(n24467), .dout(n24469));
  jor  g24305(.dina(n24469), .dinb(n24466), .dout(n24470));
  jor  g24306(.dina(n24470), .dinb(n24465), .dout(n24471));
  jxor g24307(.dina(n24471), .dinb(n4713), .dout(n24472));
  jxor g24308(.dina(n24472), .dinb(n24464), .dout(n24473));
  jxor g24309(.dina(n24473), .dinb(n24328), .dout(n24474));
  jand g24310(.dina(n23847), .dinb(n5280), .dout(n24475));
  jand g24311(.dina(n23845), .dinb(n5814), .dout(n24476));
  jand g24312(.dina(n23144), .dinb(n5531), .dout(n24477));
  jand g24313(.dina(n23079), .dinb(n5536), .dout(n24478));
  jor  g24314(.dina(n24478), .dinb(n24477), .dout(n24479));
  jor  g24315(.dina(n24479), .dinb(n24476), .dout(n24480));
  jor  g24316(.dina(n24480), .dinb(n24475), .dout(n24481));
  jxor g24317(.dina(n24481), .dinb(\a[5] ), .dout(n24482));
  jnot g24318(.din(n24482), .dout(n24483));
  jxor g24319(.dina(n24483), .dinb(n24474), .dout(n24484));
  jnot g24320(.din(n24484), .dout(n24485));
  jxor g24321(.dina(n24485), .dinb(n24323), .dout(n24486));
  jor  g24322(.dina(n24304), .dinb(n24266), .dout(n24487));
  jnot g24323(.din(n24301), .dout(n24488));
  jor  g24324(.dina(n24488), .dinb(n24271), .dout(n24489));
  jand g24325(.dina(n24489), .dinb(n24487), .dout(n24490));
  jand g24326(.dina(n24295), .dinb(n24288), .dout(n24491));
  jand g24327(.dina(n24296), .dinb(n24283), .dout(n24492));
  jor  g24328(.dina(n24492), .dinb(n24491), .dout(n24493));
  jand g24329(.dina(n17312), .dinb(n5076), .dout(n24494));
  jand g24330(.dina(n16924), .dinb(n5084), .dout(n24496));
  jand g24331(.dina(n16928), .dinb(n5082), .dout(n24497));
  jor  g24332(.dina(n24497), .dinb(n24496), .dout(n24498));
  jor  g24333(.dina(n24498), .dinb(n6050), .dout(n24499));
  jor  g24334(.dina(n24499), .dinb(n24494), .dout(n24500));
  jnot g24335(.din(n7677), .dout(n24501));
  jand g24336(.dina(n24287), .dinb(n24284), .dout(n24503));
  jnot g24337(.din(n24503), .dout(n24504));
  jand g24338(.dina(n24504), .dinb(n24069), .dout(n24505));
  jxor g24339(.dina(n24505), .dinb(n24501), .dout(n24506));
  jxor g24340(.dina(n24506), .dinb(n24500), .dout(n24507));
  jxor g24341(.dina(n24507), .dinb(n24493), .dout(n24508));
  jnot g24342(.din(n24508), .dout(n24509));
  jand g24343(.dina(n24297), .dinb(n24280), .dout(n24510));
  jnot g24344(.din(n24510), .dout(n24511));
  jor  g24345(.dina(n24299), .dinb(n24275), .dout(n24512));
  jand g24346(.dina(n24512), .dinb(n24511), .dout(n24513));
  jxor g24347(.dina(n24513), .dinb(n24509), .dout(n24514));
  jxor g24348(.dina(n24514), .dinb(n24300), .dout(n24515));
  jxor g24349(.dina(n24515), .dinb(n24490), .dout(n24516));
  jor  g24350(.dina(n24516), .dinb(n6496), .dout(n24517));
  jnot g24351(.din(n24514), .dout(n24518));
  jor  g24352(.dina(n24518), .dinb(n6504), .dout(n24519));
  jor  g24353(.dina(n24304), .dinb(n6507), .dout(n24520));
  jor  g24354(.dina(n24266), .dinb(n6501), .dout(n24521));
  jand g24355(.dina(n24521), .dinb(n24520), .dout(n24522));
  jand g24356(.dina(n24522), .dinb(n24519), .dout(n24523));
  jand g24357(.dina(n24523), .dinb(n24517), .dout(n24524));
  jxor g24358(.dina(n24524), .dinb(\a[2] ), .dout(n24525));
  jxor g24359(.dina(n24525), .dinb(n24486), .dout(n24526));
  jxor g24360(.dina(n24526), .dinb(n24319), .dout(n24527));
  jxor g24361(.dina(n24527), .dinb(n24315), .dout(\result[3] ));
  jand g24362(.dina(n24527), .dinb(n24315), .dout(n24529));
  jor  g24363(.dina(n24525), .dinb(n24486), .dout(n24530));
  jnot g24364(.din(n24530), .dout(n24531));
  jand g24365(.dina(n24526), .dinb(n24319), .dout(n24532));
  jor  g24366(.dina(n24532), .dinb(n24531), .dout(n24533));
  jand g24367(.dina(n24482), .dinb(n24474), .dout(n24534));
  jnot g24368(.din(n24534), .dout(n24535));
  jor  g24369(.dina(n24484), .dinb(n24323), .dout(n24536));
  jand g24370(.dina(n24536), .dinb(n24535), .dout(n24537));
  jor  g24371(.dina(n24472), .dinb(n24464), .dout(n24538));
  jnot g24372(.din(n24538), .dout(n24539));
  jand g24373(.dina(n24473), .dinb(n24328), .dout(n24540));
  jor  g24374(.dina(n24540), .dinb(n24539), .dout(n24541));
  jor  g24375(.dina(n24462), .dinb(n24454), .dout(n24542));
  jnot g24376(.din(n24463), .dout(n24543));
  jor  g24377(.dina(n24543), .dinb(n24333), .dout(n24544));
  jand g24378(.dina(n24544), .dinb(n24542), .dout(n24545));
  jnot g24379(.din(n24444), .dout(n24546));
  jor  g24380(.dina(n24452), .dinb(n24546), .dout(n24547));
  jnot g24381(.din(n24547), .dout(n24548));
  jnot g24382(.din(n24453), .dout(n24549));
  jand g24383(.dina(n24549), .dinb(n24337), .dout(n24550));
  jor  g24384(.dina(n24550), .dinb(n24548), .dout(n24551));
  jand g24385(.dina(n24442), .dinb(n24434), .dout(n24552));
  jand g24386(.dina(n24443), .dinb(n24342), .dout(n24553));
  jor  g24387(.dina(n24553), .dinb(n24552), .dout(n24554));
  jor  g24388(.dina(n24432), .dinb(n24424), .dout(n24555));
  jand g24389(.dina(n24433), .dinb(n24347), .dout(n24556));
  jnot g24390(.din(n24556), .dout(n24557));
  jand g24391(.dina(n24557), .dinb(n24555), .dout(n24558));
  jnot g24392(.din(n24558), .dout(n24559));
  jor  g24393(.dina(n24421), .dinb(n24413), .dout(n24560));
  jand g24394(.dina(n24422), .dinb(n24352), .dout(n24561));
  jnot g24395(.din(n24561), .dout(n24562));
  jand g24396(.dina(n24562), .dinb(n24560), .dout(n24563));
  jnot g24397(.din(n24563), .dout(n24564));
  jor  g24398(.dina(n24410), .dinb(n24402), .dout(n24565));
  jand g24399(.dina(n24411), .dinb(n24357), .dout(n24566));
  jnot g24400(.din(n24566), .dout(n24567));
  jand g24401(.dina(n24567), .dinb(n24565), .dout(n24568));
  jnot g24402(.din(n24568), .dout(n24569));
  jor  g24403(.dina(n24399), .dinb(n24391), .dout(n24570));
  jand g24404(.dina(n24400), .dinb(n24362), .dout(n24571));
  jnot g24405(.din(n24571), .dout(n24572));
  jand g24406(.dina(n24572), .dinb(n24570), .dout(n24573));
  jnot g24407(.din(n24573), .dout(n24574));
  jand g24408(.dina(n24388), .dinb(n24381), .dout(n24575));
  jand g24409(.dina(n24389), .dinb(n24365), .dout(n24576));
  jor  g24410(.dina(n24576), .dinb(n24575), .dout(n24577));
  jand g24411(.dina(n1042), .dinb(n664), .dout(n24578));
  jand g24412(.dina(n24578), .dinb(n1891), .dout(n24579));
  jand g24413(.dina(n24579), .dinb(n2409), .dout(n24580));
  jand g24414(.dina(n5180), .dinb(n1358), .dout(n24581));
  jand g24415(.dina(n24581), .dinb(n2560), .dout(n24582));
  jand g24416(.dina(n24582), .dinb(n24580), .dout(n24583));
  jand g24417(.dina(n3806), .dinb(n2394), .dout(n24584));
  jand g24418(.dina(n4422), .dinb(n3880), .dout(n24585));
  jand g24419(.dina(n24585), .dinb(n24584), .dout(n24586));
  jand g24420(.dina(n3118), .dinb(n1212), .dout(n24587));
  jand g24421(.dina(n6269), .dinb(n3978), .dout(n24588));
  jand g24422(.dina(n24588), .dinb(n24587), .dout(n24589));
  jand g24423(.dina(n24589), .dinb(n24586), .dout(n24590));
  jand g24424(.dina(n24590), .dinb(n24583), .dout(n24591));
  jand g24425(.dina(n24591), .dinb(n12443), .dout(n24592));
  jand g24426(.dina(n3771), .dinb(n130), .dout(n24593));
  jand g24427(.dina(n24593), .dinb(n23913), .dout(n24594));
  jand g24428(.dina(n8843), .dinb(n1934), .dout(n24595));
  jand g24429(.dina(n24595), .dinb(n24594), .dout(n24596));
  jand g24430(.dina(n886), .dinb(n1583), .dout(n24597));
  jand g24431(.dina(n24597), .dinb(n511), .dout(n24598));
  jand g24432(.dina(n24598), .dinb(n521), .dout(n24599));
  jand g24433(.dina(n24599), .dinb(n447), .dout(n24600));
  jand g24434(.dina(n24600), .dinb(n24596), .dout(n24601));
  jand g24435(.dina(n24601), .dinb(n9330), .dout(n24602));
  jand g24436(.dina(n24602), .dinb(n24592), .dout(n24603));
  jnot g24437(.din(n24603), .dout(n24604));
  jand g24438(.dina(n17549), .dinb(n5076), .dout(n24605));
  jand g24439(.dina(n17329), .dinb(n5084), .dout(n24606));
  jand g24440(.dina(n16940), .dinb(n6050), .dout(n24607));
  jand g24441(.dina(n17330), .dinb(n5082), .dout(n24608));
  jor  g24442(.dina(n24608), .dinb(n24607), .dout(n24609));
  jor  g24443(.dina(n24609), .dinb(n24606), .dout(n24610));
  jor  g24444(.dina(n24610), .dinb(n24605), .dout(n24611));
  jxor g24445(.dina(n24611), .dinb(n24604), .dout(n24612));
  jxor g24446(.dina(n24612), .dinb(n24577), .dout(n24613));
  jnot g24447(.din(n24613), .dout(n24614));
  jand g24448(.dina(n18514), .dinb(n2936), .dout(n24615));
  jand g24449(.dina(n17942), .dinb(n2940), .dout(n24616));
  jand g24450(.dina(n18293), .dinb(n2943), .dout(n24617));
  jor  g24451(.dina(n24617), .dinb(n24616), .dout(n24618));
  jand g24452(.dina(n17535), .dinb(n3684), .dout(n24619));
  jor  g24453(.dina(n24619), .dinb(n24618), .dout(n24620));
  jor  g24454(.dina(n24620), .dinb(n24615), .dout(n24621));
  jxor g24455(.dina(n24621), .dinb(n93), .dout(n24622));
  jxor g24456(.dina(n24622), .dinb(n24614), .dout(n24623));
  jxor g24457(.dina(n24623), .dinb(n24574), .dout(n24624));
  jnot g24458(.din(n24624), .dout(n24625));
  jand g24459(.dina(n18916), .dinb(n71), .dout(n24626));
  jand g24460(.dina(n18488), .dinb(n731), .dout(n24627));
  jand g24461(.dina(n18914), .dinb(n796), .dout(n24628));
  jor  g24462(.dina(n24628), .dinb(n24627), .dout(n24629));
  jand g24463(.dina(n18292), .dinb(n1806), .dout(n24630));
  jor  g24464(.dina(n24630), .dinb(n24629), .dout(n24631));
  jor  g24465(.dina(n24631), .dinb(n24626), .dout(n24632));
  jxor g24466(.dina(n24632), .dinb(n77), .dout(n24633));
  jxor g24467(.dina(n24633), .dinb(n24625), .dout(n24634));
  jxor g24468(.dina(n24634), .dinb(n24569), .dout(n24635));
  jnot g24469(.din(n24635), .dout(n24636));
  jand g24470(.dina(n19375), .dinb(n806), .dout(n24637));
  jand g24471(.dina(n19219), .dinb(n1612), .dout(n24638));
  jand g24472(.dina(n19373), .dinb(n1620), .dout(n24639));
  jor  g24473(.dina(n24639), .dinb(n24638), .dout(n24640));
  jand g24474(.dina(n19220), .dinb(n1644), .dout(n24641));
  jor  g24475(.dina(n24641), .dinb(n24640), .dout(n24642));
  jor  g24476(.dina(n24642), .dinb(n24637), .dout(n24643));
  jxor g24477(.dina(n24643), .dinb(n65), .dout(n24644));
  jxor g24478(.dina(n24644), .dinb(n24636), .dout(n24645));
  jxor g24479(.dina(n24645), .dinb(n24564), .dout(n24646));
  jnot g24480(.din(n24646), .dout(n24647));
  jand g24481(.dina(n20358), .dinb(n1819), .dout(n24648));
  jand g24482(.dina(n20204), .dinb(n2243), .dout(n24649));
  jand g24483(.dina(n20205), .dinb(n2180), .dout(n24650));
  jand g24484(.dina(n19922), .dinb(n2185), .dout(n24651));
  jor  g24485(.dina(n24651), .dinb(n24650), .dout(n24652));
  jor  g24486(.dina(n24652), .dinb(n24649), .dout(n24653));
  jor  g24487(.dina(n24653), .dinb(n24648), .dout(n24654));
  jxor g24488(.dina(n24654), .dinb(n2196), .dout(n24655));
  jxor g24489(.dina(n24655), .dinb(n24647), .dout(n24656));
  jxor g24490(.dina(n24656), .dinb(n24559), .dout(n24657));
  jand g24491(.dina(n21367), .dinb(n2743), .dout(n24658));
  jand g24492(.dina(n21198), .dinb(n2752), .dout(n24659));
  jand g24493(.dina(n20947), .dinb(n2748), .dout(n24660));
  jand g24494(.dina(n20344), .dinb(n2757), .dout(n24661));
  jor  g24495(.dina(n24661), .dinb(n24660), .dout(n24662));
  jor  g24496(.dina(n24662), .dinb(n24659), .dout(n24663));
  jor  g24497(.dina(n24663), .dinb(n24658), .dout(n24664));
  jxor g24498(.dina(n24664), .dinb(\a[17] ), .dout(n24665));
  jxor g24499(.dina(n24665), .dinb(n24657), .dout(n24666));
  jxor g24500(.dina(n24666), .dinb(n24554), .dout(n24667));
  jand g24501(.dina(n21976), .dinb(n3423), .dout(n24668));
  jand g24502(.dina(n21974), .dinb(n3569), .dout(n24669));
  jand g24503(.dina(n21340), .dinb(n3428), .dout(n24670));
  jand g24504(.dina(n21197), .dinb(n3210), .dout(n24671));
  jor  g24505(.dina(n24671), .dinb(n24670), .dout(n24672));
  jor  g24506(.dina(n24672), .dinb(n24669), .dout(n24673));
  jor  g24507(.dina(n24673), .dinb(n24668), .dout(n24674));
  jxor g24508(.dina(n24674), .dinb(n3473), .dout(n24675));
  jxor g24509(.dina(n24675), .dinb(n24667), .dout(n24676));
  jnot g24510(.din(n24676), .dout(n24677));
  jxor g24511(.dina(n24677), .dinb(n24551), .dout(n24678));
  jand g24512(.dina(n22267), .dinb(n4022), .dout(n24679));
  jand g24513(.dina(n22265), .dinb(n4220), .dout(n24680));
  jand g24514(.dina(n22163), .dinb(n4027), .dout(n24681));
  jand g24515(.dina(n22164), .dinb(n3870), .dout(n24682));
  jor  g24516(.dina(n24682), .dinb(n24681), .dout(n24683));
  jor  g24517(.dina(n24683), .dinb(n24680), .dout(n24684));
  jor  g24518(.dina(n24684), .dinb(n24679), .dout(n24685));
  jxor g24519(.dina(n24685), .dinb(n4050), .dout(n24686));
  jxor g24520(.dina(n24686), .dinb(n24678), .dout(n24687));
  jnot g24521(.din(n24687), .dout(n24688));
  jxor g24522(.dina(n24688), .dinb(n24545), .dout(n24689));
  jand g24523(.dina(n23159), .dinb(n4691), .dout(n24690));
  jand g24524(.dina(n23080), .dinb(n4696), .dout(n24691));
  jand g24525(.dina(n23079), .dinb(n4941), .dout(n24692));
  jor  g24526(.dina(n24692), .dinb(n24691), .dout(n24693));
  jand g24527(.dina(n22937), .dinb(n4701), .dout(n24694));
  jor  g24528(.dina(n24694), .dinb(n24693), .dout(n24695));
  jor  g24529(.dina(n24695), .dinb(n24690), .dout(n24696));
  jxor g24530(.dina(n24696), .dinb(n4713), .dout(n24697));
  jxor g24531(.dina(n24697), .dinb(n24689), .dout(n24698));
  jxor g24532(.dina(n24698), .dinb(n24541), .dout(n24699));
  jand g24533(.dina(n24077), .dinb(n5280), .dout(n24700));
  jand g24534(.dina(n23845), .dinb(n5531), .dout(n24701));
  jand g24535(.dina(n24075), .dinb(n5814), .dout(n24702));
  jor  g24536(.dina(n24702), .dinb(n24701), .dout(n24703));
  jand g24537(.dina(n23144), .dinb(n5536), .dout(n24704));
  jor  g24538(.dina(n24704), .dinb(n24703), .dout(n24705));
  jor  g24539(.dina(n24705), .dinb(n24700), .dout(n24706));
  jxor g24540(.dina(n24706), .dinb(n5277), .dout(n24707));
  jxor g24541(.dina(n24707), .dinb(n24699), .dout(n24708));
  jnot g24542(.din(n24708), .dout(n24709));
  jxor g24543(.dina(n24709), .dinb(n24537), .dout(n24710));
  jor  g24544(.dina(n24518), .dinb(n24304), .dout(n24711));
  jnot g24545(.din(n24515), .dout(n24712));
  jor  g24546(.dina(n24712), .dinb(n24490), .dout(n24713));
  jand g24547(.dina(n24713), .dinb(n24711), .dout(n24714));
  jor  g24548(.dina(n17296), .dinb(n7061), .dout(n24715));
  jnot g24549(.din(n6050), .dout(n24716));
  jand g24550(.dina(n142), .dinb(n5078), .dout(n24718));
  jor  g24551(.dina(n24718), .dinb(n17301), .dout(n24719));
  jor  g24552(.dina(n24719), .dinb(n5080), .dout(n24720));
  jand g24553(.dina(n24720), .dinb(n24716), .dout(n24721));
  jand g24554(.dina(n24721), .dinb(n24715), .dout(n24722));
  jxor g24555(.dina(n24722), .dinb(n7677), .dout(n24723));
  jand g24556(.dina(n24506), .dinb(n24500), .dout(n24725));
  jnot g24557(.din(n24725), .dout(n24726));
  jand g24558(.dina(n24726), .dinb(n24505), .dout(n24727));
  jxor g24559(.dina(n24727), .dinb(n24723), .dout(n24728));
  jnot g24560(.din(n24728), .dout(n24729));
  jand g24561(.dina(n24507), .dinb(n24493), .dout(n24730));
  jnot g24562(.din(n24730), .dout(n24731));
  jor  g24563(.dina(n24513), .dinb(n24509), .dout(n24732));
  jand g24564(.dina(n24732), .dinb(n24731), .dout(n24733));
  jxor g24565(.dina(n24733), .dinb(n24729), .dout(n24734));
  jxor g24566(.dina(n24734), .dinb(n24514), .dout(n24735));
  jxor g24567(.dina(n24735), .dinb(n24714), .dout(n24736));
  jor  g24568(.dina(n24736), .dinb(n6496), .dout(n24737));
  jnot g24569(.din(n24734), .dout(n24738));
  jor  g24570(.dina(n24738), .dinb(n6504), .dout(n24739));
  jor  g24571(.dina(n24518), .dinb(n6507), .dout(n24740));
  jor  g24572(.dina(n24304), .dinb(n6501), .dout(n24741));
  jand g24573(.dina(n24741), .dinb(n24740), .dout(n24742));
  jand g24574(.dina(n24742), .dinb(n24739), .dout(n24743));
  jand g24575(.dina(n24743), .dinb(n24737), .dout(n24744));
  jxor g24576(.dina(n24744), .dinb(\a[2] ), .dout(n24745));
  jxor g24577(.dina(n24745), .dinb(n24710), .dout(n24746));
  jxor g24578(.dina(n24746), .dinb(n24533), .dout(n24747));
  jxor g24579(.dina(n24747), .dinb(n24529), .dout(\result[4] ));
  jand g24580(.dina(n24747), .dinb(n24529), .dout(n24749));
  jor  g24581(.dina(n24745), .dinb(n24710), .dout(n24750));
  jnot g24582(.din(n24750), .dout(n24751));
  jand g24583(.dina(n24746), .dinb(n24533), .dout(n24752));
  jor  g24584(.dina(n24752), .dinb(n24751), .dout(n24753));
  jnot g24585(.din(n24699), .dout(n24754));
  jor  g24586(.dina(n24707), .dinb(n24754), .dout(n24755));
  jor  g24587(.dina(n24708), .dinb(n24537), .dout(n24756));
  jand g24588(.dina(n24756), .dinb(n24755), .dout(n24757));
  jnot g24589(.din(n24757), .dout(n24758));
  jor  g24590(.dina(n24697), .dinb(n24689), .dout(n24759));
  jnot g24591(.din(n24759), .dout(n24760));
  jand g24592(.dina(n24698), .dinb(n24541), .dout(n24761));
  jor  g24593(.dina(n24761), .dinb(n24760), .dout(n24762));
  jnot g24594(.din(n24678), .dout(n24763));
  jor  g24595(.dina(n24686), .dinb(n24763), .dout(n24764));
  jor  g24596(.dina(n24687), .dinb(n24545), .dout(n24765));
  jand g24597(.dina(n24765), .dinb(n24764), .dout(n24766));
  jnot g24598(.din(n24667), .dout(n24767));
  jor  g24599(.dina(n24675), .dinb(n24767), .dout(n24768));
  jnot g24600(.din(n24768), .dout(n24769));
  jand g24601(.dina(n24677), .dinb(n24551), .dout(n24770));
  jor  g24602(.dina(n24770), .dinb(n24769), .dout(n24771));
  jand g24603(.dina(n24665), .dinb(n24657), .dout(n24772));
  jand g24604(.dina(n24666), .dinb(n24554), .dout(n24773));
  jor  g24605(.dina(n24773), .dinb(n24772), .dout(n24774));
  jor  g24606(.dina(n24655), .dinb(n24647), .dout(n24775));
  jand g24607(.dina(n24656), .dinb(n24559), .dout(n24776));
  jnot g24608(.din(n24776), .dout(n24777));
  jand g24609(.dina(n24777), .dinb(n24775), .dout(n24778));
  jnot g24610(.din(n24778), .dout(n24779));
  jor  g24611(.dina(n24644), .dinb(n24636), .dout(n24780));
  jand g24612(.dina(n24645), .dinb(n24564), .dout(n24781));
  jnot g24613(.din(n24781), .dout(n24782));
  jand g24614(.dina(n24782), .dinb(n24780), .dout(n24783));
  jnot g24615(.din(n24783), .dout(n24784));
  jor  g24616(.dina(n24633), .dinb(n24625), .dout(n24785));
  jand g24617(.dina(n24634), .dinb(n24569), .dout(n24786));
  jnot g24618(.din(n24786), .dout(n24787));
  jand g24619(.dina(n24787), .dinb(n24785), .dout(n24788));
  jnot g24620(.din(n24788), .dout(n24789));
  jor  g24621(.dina(n24622), .dinb(n24614), .dout(n24790));
  jand g24622(.dina(n24623), .dinb(n24574), .dout(n24791));
  jnot g24623(.din(n24791), .dout(n24792));
  jand g24624(.dina(n24792), .dinb(n24790), .dout(n24793));
  jnot g24625(.din(n24793), .dout(n24794));
  jand g24626(.dina(n24611), .dinb(n24604), .dout(n24795));
  jand g24627(.dina(n24612), .dinb(n24577), .dout(n24796));
  jor  g24628(.dina(n24796), .dinb(n24795), .dout(n24797));
  jand g24629(.dina(n1515), .dinb(n270), .dout(n24798));
  jand g24630(.dina(n24798), .dinb(n583), .dout(n24799));
  jand g24631(.dina(n24799), .dinb(n654), .dout(n24800));
  jand g24632(.dina(n24800), .dinb(n6198), .dout(n24801));
  jand g24633(.dina(n24801), .dinb(n13521), .dout(n24802));
  jand g24634(.dina(n6019), .dinb(n1246), .dout(n24803));
  jand g24635(.dina(n1167), .dinb(n1213), .dout(n24804));
  jand g24636(.dina(n24804), .dinb(n24803), .dout(n24805));
  jand g24637(.dina(n24805), .dinb(n5232), .dout(n24806));
  jand g24638(.dina(n24806), .dinb(n24802), .dout(n24807));
  jand g24639(.dina(n4448), .dinb(n1961), .dout(n24808));
  jand g24640(.dina(n13394), .dinb(n4675), .dout(n24809));
  jand g24641(.dina(n24809), .dinb(n24808), .dout(n24810));
  jand g24642(.dina(n24810), .dinb(n24807), .dout(n24811));
  jand g24643(.dina(n24811), .dinb(n15679), .dout(n24812));
  jand g24644(.dina(n24812), .dinb(n10159), .dout(n24813));
  jnot g24645(.din(n24813), .dout(n24814));
  jand g24646(.dina(n17537), .dinb(n5076), .dout(n24815));
  jand g24647(.dina(n17535), .dinb(n5084), .dout(n24816));
  jand g24648(.dina(n17330), .dinb(n6050), .dout(n24817));
  jand g24649(.dina(n17329), .dinb(n5082), .dout(n24818));
  jor  g24650(.dina(n24818), .dinb(n24817), .dout(n24819));
  jor  g24651(.dina(n24819), .dinb(n24816), .dout(n24820));
  jor  g24652(.dina(n24820), .dinb(n24815), .dout(n24821));
  jxor g24653(.dina(n24821), .dinb(n24814), .dout(n24822));
  jxor g24654(.dina(n24822), .dinb(n24797), .dout(n24823));
  jnot g24655(.din(n24823), .dout(n24824));
  jand g24656(.dina(n18502), .dinb(n2936), .dout(n24825));
  jand g24657(.dina(n18293), .dinb(n2940), .dout(n24826));
  jand g24658(.dina(n18292), .dinb(n2943), .dout(n24827));
  jor  g24659(.dina(n24827), .dinb(n24826), .dout(n24828));
  jand g24660(.dina(n17942), .dinb(n3684), .dout(n24829));
  jor  g24661(.dina(n24829), .dinb(n24828), .dout(n24830));
  jor  g24662(.dina(n24830), .dinb(n24825), .dout(n24831));
  jxor g24663(.dina(n24831), .dinb(n93), .dout(n24832));
  jxor g24664(.dina(n24832), .dinb(n24824), .dout(n24833));
  jxor g24665(.dina(n24833), .dinb(n24794), .dout(n24834));
  jnot g24666(.din(n24834), .dout(n24835));
  jand g24667(.dina(n19399), .dinb(n71), .dout(n24836));
  jand g24668(.dina(n19220), .dinb(n796), .dout(n24837));
  jand g24669(.dina(n18914), .dinb(n731), .dout(n24838));
  jand g24670(.dina(n18488), .dinb(n1806), .dout(n24839));
  jor  g24671(.dina(n24839), .dinb(n24838), .dout(n24840));
  jor  g24672(.dina(n24840), .dinb(n24837), .dout(n24841));
  jor  g24673(.dina(n24841), .dinb(n24836), .dout(n24842));
  jxor g24674(.dina(n24842), .dinb(n77), .dout(n24843));
  jxor g24675(.dina(n24843), .dinb(n24835), .dout(n24844));
  jxor g24676(.dina(n24844), .dinb(n24789), .dout(n24845));
  jnot g24677(.din(n24845), .dout(n24846));
  jand g24678(.dina(n19924), .dinb(n806), .dout(n24847));
  jand g24679(.dina(n19373), .dinb(n1612), .dout(n24848));
  jand g24680(.dina(n19922), .dinb(n1620), .dout(n24849));
  jor  g24681(.dina(n24849), .dinb(n24848), .dout(n24850));
  jand g24682(.dina(n19219), .dinb(n1644), .dout(n24851));
  jor  g24683(.dina(n24851), .dinb(n24850), .dout(n24852));
  jor  g24684(.dina(n24852), .dinb(n24847), .dout(n24853));
  jxor g24685(.dina(n24853), .dinb(n65), .dout(n24854));
  jxor g24686(.dina(n24854), .dinb(n24846), .dout(n24855));
  jxor g24687(.dina(n24855), .dinb(n24784), .dout(n24856));
  jnot g24688(.din(n24856), .dout(n24857));
  jand g24689(.dina(n20346), .dinb(n1819), .dout(n24858));
  jand g24690(.dina(n20344), .dinb(n2243), .dout(n24859));
  jand g24691(.dina(n20204), .dinb(n2180), .dout(n24860));
  jand g24692(.dina(n20205), .dinb(n2185), .dout(n24861));
  jor  g24693(.dina(n24861), .dinb(n24860), .dout(n24862));
  jor  g24694(.dina(n24862), .dinb(n24859), .dout(n24863));
  jor  g24695(.dina(n24863), .dinb(n24858), .dout(n24864));
  jxor g24696(.dina(n24864), .dinb(n2196), .dout(n24865));
  jxor g24697(.dina(n24865), .dinb(n24857), .dout(n24866));
  jxor g24698(.dina(n24866), .dinb(n24779), .dout(n24867));
  jand g24699(.dina(n21355), .dinb(n2743), .dout(n24868));
  jand g24700(.dina(n21197), .dinb(n2752), .dout(n24869));
  jand g24701(.dina(n21198), .dinb(n2748), .dout(n24870));
  jand g24702(.dina(n20947), .dinb(n2757), .dout(n24871));
  jor  g24703(.dina(n24871), .dinb(n24870), .dout(n24872));
  jor  g24704(.dina(n24872), .dinb(n24869), .dout(n24873));
  jor  g24705(.dina(n24873), .dinb(n24868), .dout(n24874));
  jxor g24706(.dina(n24874), .dinb(n2441), .dout(n24875));
  jxor g24707(.dina(n24875), .dinb(n24867), .dout(n24876));
  jxor g24708(.dina(n24876), .dinb(n24774), .dout(n24877));
  jand g24709(.dina(n22291), .dinb(n3423), .dout(n24878));
  jand g24710(.dina(n22164), .dinb(n3569), .dout(n24879));
  jand g24711(.dina(n21974), .dinb(n3428), .dout(n24880));
  jand g24712(.dina(n21340), .dinb(n3210), .dout(n24881));
  jor  g24713(.dina(n24881), .dinb(n24880), .dout(n24882));
  jor  g24714(.dina(n24882), .dinb(n24879), .dout(n24883));
  jor  g24715(.dina(n24883), .dinb(n24878), .dout(n24884));
  jxor g24716(.dina(n24884), .dinb(n3473), .dout(n24885));
  jxor g24717(.dina(n24885), .dinb(n24877), .dout(n24886));
  jxor g24718(.dina(n24886), .dinb(n24771), .dout(n24887));
  jnot g24719(.din(n24887), .dout(n24888));
  jand g24720(.dina(n22939), .dinb(n4022), .dout(n24889));
  jand g24721(.dina(n22265), .dinb(n4027), .dout(n24890));
  jand g24722(.dina(n22937), .dinb(n4220), .dout(n24891));
  jor  g24723(.dina(n24891), .dinb(n24890), .dout(n24892));
  jand g24724(.dina(n22163), .dinb(n3870), .dout(n24893));
  jor  g24725(.dina(n24893), .dinb(n24892), .dout(n24894));
  jor  g24726(.dina(n24894), .dinb(n24889), .dout(n24895));
  jxor g24727(.dina(n24895), .dinb(n4050), .dout(n24896));
  jxor g24728(.dina(n24896), .dinb(n24888), .dout(n24897));
  jxor g24729(.dina(n24897), .dinb(n24766), .dout(n24898));
  jand g24730(.dina(n23146), .dinb(n4691), .dout(n24899));
  jand g24731(.dina(n23144), .dinb(n4941), .dout(n24900));
  jand g24732(.dina(n23079), .dinb(n4696), .dout(n24901));
  jand g24733(.dina(n23080), .dinb(n4701), .dout(n24902));
  jor  g24734(.dina(n24902), .dinb(n24901), .dout(n24903));
  jor  g24735(.dina(n24903), .dinb(n24900), .dout(n24904));
  jor  g24736(.dina(n24904), .dinb(n24899), .dout(n24905));
  jxor g24737(.dina(n24905), .dinb(n4713), .dout(n24906));
  jxor g24738(.dina(n24906), .dinb(n24898), .dout(n24907));
  jnot g24739(.din(n24907), .dout(n24908));
  jxor g24740(.dina(n24908), .dinb(n24762), .dout(n24909));
  jor  g24741(.dina(n24302), .dinb(n5281), .dout(n24910));
  jor  g24742(.dina(n24266), .dinb(n5532), .dout(n24911));
  jor  g24743(.dina(n24304), .dinb(n5539), .dout(n24912));
  jand g24744(.dina(n24912), .dinb(n24911), .dout(n24913));
  jor  g24745(.dina(n24265), .dinb(n5537), .dout(n24914));
  jand g24746(.dina(n24914), .dinb(n24913), .dout(n24915));
  jand g24747(.dina(n24915), .dinb(n24910), .dout(n24916));
  jxor g24748(.dina(n24916), .dinb(\a[5] ), .dout(n24917));
  jxor g24749(.dina(n24917), .dinb(n24909), .dout(n24918));
  jxor g24750(.dina(n24918), .dinb(n24758), .dout(n24919));
  jor  g24751(.dina(n24738), .dinb(n24518), .dout(n24920));
  jnot g24752(.din(n24735), .dout(n24921));
  jor  g24753(.dina(n24921), .dinb(n24714), .dout(n24922));
  jand g24754(.dina(n24922), .dinb(n24920), .dout(n24923));
  jor  g24755(.dina(n24727), .dinb(n24723), .dout(n24924));
  jor  g24756(.dina(n24733), .dinb(n24729), .dout(n24925));
  jand g24757(.dina(n24925), .dinb(n24924), .dout(n24926));
  jand g24758(.dina(n24722), .dinb(n7677), .dout(n24927));
  jxor g24759(.dina(n24927), .dinb(n24719), .dout(n24928));
  jnot g24760(.din(n24928), .dout(n24929));
  jxor g24761(.dina(n24929), .dinb(n24926), .dout(n24930));
  jxor g24762(.dina(n24930), .dinb(n24738), .dout(n24931));
  jxor g24763(.dina(n24931), .dinb(n24923), .dout(n24932));
  jor  g24764(.dina(n24932), .dinb(n6496), .dout(n24933));
  jor  g24765(.dina(n24930), .dinb(n6504), .dout(n24934));
  jor  g24766(.dina(n24738), .dinb(n6507), .dout(n24935));
  jor  g24767(.dina(n24518), .dinb(n6501), .dout(n24936));
  jand g24768(.dina(n24936), .dinb(n24935), .dout(n24937));
  jand g24769(.dina(n24937), .dinb(n24934), .dout(n24938));
  jand g24770(.dina(n24938), .dinb(n24933), .dout(n24939));
  jxor g24771(.dina(n24939), .dinb(\a[2] ), .dout(n24940));
  jnot g24772(.din(n24940), .dout(n24941));
  jxor g24773(.dina(n24941), .dinb(n24919), .dout(n24942));
  jxor g24774(.dina(n24942), .dinb(n24753), .dout(n24943));
  jxor g24775(.dina(n24943), .dinb(n24749), .dout(\result[5] ));
  jand g24776(.dina(n24943), .dinb(n24749), .dout(n24945));
  jor  g24777(.dina(n24917), .dinb(n24909), .dout(n24946));
  jnot g24778(.din(n24946), .dout(n24947));
  jand g24779(.dina(n24918), .dinb(n24758), .dout(n24948));
  jor  g24780(.dina(n24948), .dinb(n24947), .dout(n24949));
  jor  g24781(.dina(n24906), .dinb(n24898), .dout(n24950));
  jnot g24782(.din(n24950), .dout(n24951));
  jand g24783(.dina(n24907), .dinb(n24762), .dout(n24952));
  jor  g24784(.dina(n24952), .dinb(n24951), .dout(n24953));
  jor  g24785(.dina(n24896), .dinb(n24888), .dout(n24954));
  jnot g24786(.din(n24897), .dout(n24955));
  jor  g24787(.dina(n24955), .dinb(n24766), .dout(n24956));
  jand g24788(.dina(n24956), .dinb(n24954), .dout(n24957));
  jor  g24789(.dina(n24885), .dinb(n24877), .dout(n24958));
  jnot g24790(.din(n24958), .dout(n24959));
  jand g24791(.dina(n24886), .dinb(n24771), .dout(n24960));
  jor  g24792(.dina(n24960), .dinb(n24959), .dout(n24961));
  jnot g24793(.din(n24867), .dout(n24962));
  jor  g24794(.dina(n24875), .dinb(n24962), .dout(n24963));
  jnot g24795(.din(n24774), .dout(n24964));
  jor  g24796(.dina(n24876), .dinb(n24964), .dout(n24965));
  jand g24797(.dina(n24965), .dinb(n24963), .dout(n24966));
  jor  g24798(.dina(n24865), .dinb(n24857), .dout(n24967));
  jnot g24799(.din(n24967), .dout(n24968));
  jand g24800(.dina(n24866), .dinb(n24779), .dout(n24969));
  jor  g24801(.dina(n24969), .dinb(n24968), .dout(n24970));
  jor  g24802(.dina(n24854), .dinb(n24846), .dout(n24971));
  jand g24803(.dina(n24855), .dinb(n24784), .dout(n24972));
  jnot g24804(.din(n24972), .dout(n24973));
  jand g24805(.dina(n24973), .dinb(n24971), .dout(n24974));
  jnot g24806(.din(n24974), .dout(n24975));
  jor  g24807(.dina(n24843), .dinb(n24835), .dout(n24976));
  jand g24808(.dina(n24844), .dinb(n24789), .dout(n24977));
  jnot g24809(.din(n24977), .dout(n24978));
  jand g24810(.dina(n24978), .dinb(n24976), .dout(n24979));
  jnot g24811(.din(n24979), .dout(n24980));
  jor  g24812(.dina(n24832), .dinb(n24824), .dout(n24981));
  jand g24813(.dina(n24833), .dinb(n24794), .dout(n24982));
  jnot g24814(.din(n24982), .dout(n24983));
  jand g24815(.dina(n24983), .dinb(n24981), .dout(n24984));
  jnot g24816(.din(n24984), .dout(n24985));
  jand g24817(.dina(n24821), .dinb(n24814), .dout(n24986));
  jand g24818(.dina(n24822), .dinb(n24797), .dout(n24987));
  jor  g24819(.dina(n24987), .dinb(n24986), .dout(n24988));
  jand g24820(.dina(n24367), .dinb(n18980), .dout(n24989));
  jand g24821(.dina(n1987), .dinb(n1915), .dout(n24990));
  jand g24822(.dina(n24990), .dinb(n2620), .dout(n24991));
  jand g24823(.dina(n24991), .dinb(n24989), .dout(n24992));
  jand g24824(.dina(n10390), .dinb(n6269), .dout(n24993));
  jand g24825(.dina(n1378), .dinb(n638), .dout(n24994));
  jand g24826(.dina(n24994), .dinb(n172), .dout(n24995));
  jand g24827(.dina(n24995), .dinb(n24993), .dout(n24996));
  jand g24828(.dina(n3182), .dinb(n1772), .dout(n24997));
  jand g24829(.dina(n24997), .dinb(n4423), .dout(n24998));
  jand g24830(.dina(n24998), .dinb(n411), .dout(n24999));
  jand g24831(.dina(n24999), .dinb(n24996), .dout(n25000));
  jand g24832(.dina(n25000), .dinb(n24992), .dout(n25001));
  jand g24833(.dina(n25001), .dinb(n17796), .dout(n25002));
  jand g24834(.dina(n6228), .dinb(n1872), .dout(n25003));
  jand g24835(.dina(n3108), .dinb(n1208), .dout(n25004));
  jand g24836(.dina(n25004), .dinb(n10375), .dout(n25005));
  jand g24837(.dina(n25005), .dinb(n25003), .dout(n25006));
  jand g24838(.dina(n25006), .dinb(n1761), .dout(n25007));
  jand g24839(.dina(n25007), .dinb(n10416), .dout(n25008));
  jand g24840(.dina(n25008), .dinb(n25002), .dout(n25009));
  jnot g24841(.din(n25009), .dout(n25010));
  jand g24842(.dina(n17944), .dinb(n5076), .dout(n25011));
  jand g24843(.dina(n17942), .dinb(n5084), .dout(n25012));
  jand g24844(.dina(n17329), .dinb(n6050), .dout(n25013));
  jand g24845(.dina(n17535), .dinb(n5082), .dout(n25014));
  jor  g24846(.dina(n25014), .dinb(n25013), .dout(n25015));
  jor  g24847(.dina(n25015), .dinb(n25012), .dout(n25016));
  jor  g24848(.dina(n25016), .dinb(n25011), .dout(n25017));
  jxor g24849(.dina(n25017), .dinb(n25010), .dout(n25018));
  jxor g24850(.dina(n25018), .dinb(n24988), .dout(n25019));
  jnot g24851(.din(n25019), .dout(n25020));
  jand g24852(.dina(n18490), .dinb(n2936), .dout(n25021));
  jand g24853(.dina(n18488), .dinb(n2943), .dout(n25022));
  jand g24854(.dina(n18292), .dinb(n2940), .dout(n25023));
  jand g24855(.dina(n18293), .dinb(n3684), .dout(n25024));
  jor  g24856(.dina(n25024), .dinb(n25023), .dout(n25025));
  jor  g24857(.dina(n25025), .dinb(n25022), .dout(n25026));
  jor  g24858(.dina(n25026), .dinb(n25021), .dout(n25027));
  jxor g24859(.dina(n25027), .dinb(n93), .dout(n25028));
  jxor g24860(.dina(n25028), .dinb(n25020), .dout(n25029));
  jxor g24861(.dina(n25029), .dinb(n24985), .dout(n25030));
  jnot g24862(.din(n25030), .dout(n25031));
  jand g24863(.dina(n19387), .dinb(n71), .dout(n25032));
  jand g24864(.dina(n19219), .dinb(n796), .dout(n25033));
  jand g24865(.dina(n19220), .dinb(n731), .dout(n25034));
  jand g24866(.dina(n18914), .dinb(n1806), .dout(n25035));
  jor  g24867(.dina(n25035), .dinb(n25034), .dout(n25036));
  jor  g24868(.dina(n25036), .dinb(n25033), .dout(n25037));
  jor  g24869(.dina(n25037), .dinb(n25032), .dout(n25038));
  jxor g24870(.dina(n25038), .dinb(n77), .dout(n25039));
  jxor g24871(.dina(n25039), .dinb(n25031), .dout(n25040));
  jxor g24872(.dina(n25040), .dinb(n24980), .dout(n25041));
  jnot g24873(.din(n25041), .dout(n25042));
  jand g24874(.dina(n20371), .dinb(n806), .dout(n25043));
  jand g24875(.dina(n20205), .dinb(n1620), .dout(n25044));
  jand g24876(.dina(n19922), .dinb(n1612), .dout(n25045));
  jand g24877(.dina(n19373), .dinb(n1644), .dout(n25046));
  jor  g24878(.dina(n25046), .dinb(n25045), .dout(n25047));
  jor  g24879(.dina(n25047), .dinb(n25044), .dout(n25048));
  jor  g24880(.dina(n25048), .dinb(n25043), .dout(n25049));
  jxor g24881(.dina(n25049), .dinb(n65), .dout(n25050));
  jxor g24882(.dina(n25050), .dinb(n25042), .dout(n25051));
  jxor g24883(.dina(n25051), .dinb(n24975), .dout(n25052));
  jnot g24884(.din(n25052), .dout(n25053));
  jand g24885(.dina(n20949), .dinb(n1819), .dout(n25054));
  jand g24886(.dina(n20344), .dinb(n2180), .dout(n25055));
  jand g24887(.dina(n20947), .dinb(n2243), .dout(n25056));
  jor  g24888(.dina(n25056), .dinb(n25055), .dout(n25057));
  jand g24889(.dina(n20204), .dinb(n2185), .dout(n25058));
  jor  g24890(.dina(n25058), .dinb(n25057), .dout(n25059));
  jor  g24891(.dina(n25059), .dinb(n25054), .dout(n25060));
  jxor g24892(.dina(n25060), .dinb(n2196), .dout(n25061));
  jxor g24893(.dina(n25061), .dinb(n25053), .dout(n25062));
  jxor g24894(.dina(n25062), .dinb(n24970), .dout(n25063));
  jand g24895(.dina(n21342), .dinb(n2743), .dout(n25064));
  jand g24896(.dina(n21340), .dinb(n2752), .dout(n25065));
  jand g24897(.dina(n21197), .dinb(n2748), .dout(n25066));
  jand g24898(.dina(n21198), .dinb(n2757), .dout(n25067));
  jor  g24899(.dina(n25067), .dinb(n25066), .dout(n25068));
  jor  g24900(.dina(n25068), .dinb(n25065), .dout(n25069));
  jor  g24901(.dina(n25069), .dinb(n25064), .dout(n25070));
  jxor g24902(.dina(n25070), .dinb(\a[17] ), .dout(n25071));
  jxor g24903(.dina(n25071), .dinb(n25063), .dout(n25072));
  jxor g24904(.dina(n25072), .dinb(n24966), .dout(n25073));
  jand g24905(.dina(n22279), .dinb(n3423), .dout(n25074));
  jand g24906(.dina(n22164), .dinb(n3428), .dout(n25075));
  jand g24907(.dina(n22163), .dinb(n3569), .dout(n25076));
  jor  g24908(.dina(n25076), .dinb(n25075), .dout(n25077));
  jand g24909(.dina(n21974), .dinb(n3210), .dout(n25078));
  jor  g24910(.dina(n25078), .dinb(n25077), .dout(n25079));
  jor  g24911(.dina(n25079), .dinb(n25074), .dout(n25080));
  jxor g24912(.dina(n25080), .dinb(n3473), .dout(n25081));
  jxor g24913(.dina(n25081), .dinb(n25073), .dout(n25082));
  jxor g24914(.dina(n25082), .dinb(n24961), .dout(n25083));
  jand g24915(.dina(n23172), .dinb(n4022), .dout(n25084));
  jand g24916(.dina(n23080), .dinb(n4220), .dout(n25085));
  jand g24917(.dina(n22937), .dinb(n4027), .dout(n25086));
  jand g24918(.dina(n22265), .dinb(n3870), .dout(n25087));
  jor  g24919(.dina(n25087), .dinb(n25086), .dout(n25088));
  jor  g24920(.dina(n25088), .dinb(n25085), .dout(n25089));
  jor  g24921(.dina(n25089), .dinb(n25084), .dout(n25090));
  jxor g24922(.dina(n25090), .dinb(\a[11] ), .dout(n25091));
  jxor g24923(.dina(n25091), .dinb(n25083), .dout(n25092));
  jxor g24924(.dina(n25092), .dinb(n24957), .dout(n25093));
  jand g24925(.dina(n23847), .dinb(n4691), .dout(n25094));
  jand g24926(.dina(n23144), .dinb(n4696), .dout(n25095));
  jand g24927(.dina(n23845), .dinb(n4941), .dout(n25096));
  jor  g24928(.dina(n25096), .dinb(n25095), .dout(n25097));
  jand g24929(.dina(n23079), .dinb(n4701), .dout(n25098));
  jor  g24930(.dina(n25098), .dinb(n25097), .dout(n25099));
  jor  g24931(.dina(n25099), .dinb(n25094), .dout(n25100));
  jxor g24932(.dina(n25100), .dinb(n4713), .dout(n25101));
  jxor g24933(.dina(n25101), .dinb(n25093), .dout(n25102));
  jxor g24934(.dina(n25102), .dinb(n24953), .dout(n25103));
  jor  g24935(.dina(n24516), .dinb(n5281), .dout(n25104));
  jor  g24936(.dina(n24304), .dinb(n5532), .dout(n25105));
  jor  g24937(.dina(n24518), .dinb(n5539), .dout(n25106));
  jand g24938(.dina(n25106), .dinb(n25105), .dout(n25107));
  jor  g24939(.dina(n24266), .dinb(n5537), .dout(n25108));
  jand g24940(.dina(n25108), .dinb(n25107), .dout(n25109));
  jand g24941(.dina(n25109), .dinb(n25104), .dout(n25110));
  jxor g24942(.dina(n25110), .dinb(\a[5] ), .dout(n25111));
  jxor g24943(.dina(n25111), .dinb(n25103), .dout(n25112));
  jor  g24944(.dina(n24930), .dinb(n24738), .dout(n25113));
  jnot g24945(.din(n24931), .dout(n25114));
  jor  g24946(.dina(n25114), .dinb(n24923), .dout(n25115));
  jand g24947(.dina(n25115), .dinb(n25113), .dout(n25116));
  jor  g24948(.dina(n25116), .dinb(n6496), .dout(n25117));
  jor  g24949(.dina(n24930), .dinb(n17303), .dout(n25118));
  jor  g24950(.dina(n24738), .dinb(n6501), .dout(n25119));
  jand g24951(.dina(n25119), .dinb(n25118), .dout(n25120));
  jand g24952(.dina(n25120), .dinb(n25117), .dout(n25121));
  jxor g24953(.dina(n25121), .dinb(\a[2] ), .dout(n25122));
  jxor g24954(.dina(n25122), .dinb(n25112), .dout(n25123));
  jxor g24955(.dina(n25123), .dinb(n24949), .dout(n25124));
  jand g24956(.dina(n24941), .dinb(n24919), .dout(n25125));
  jand g24957(.dina(n24942), .dinb(n24753), .dout(n25126));
  jor  g24958(.dina(n25126), .dinb(n25125), .dout(n25127));
  jxor g24959(.dina(n25127), .dinb(n25124), .dout(n25128));
  jxor g24960(.dina(n25128), .dinb(n24945), .dout(\result[6] ));
  jand g24961(.dina(n25128), .dinb(n24945), .dout(n25130));
  jnot g24962(.din(n25103), .dout(n25131));
  jor  g24963(.dina(n25111), .dinb(n25131), .dout(n25132));
  jor  g24964(.dina(n25122), .dinb(n25112), .dout(n25133));
  jand g24965(.dina(n25133), .dinb(n25132), .dout(n25134));
  jnot g24966(.din(n25134), .dout(n25135));
  jor  g24967(.dina(n25101), .dinb(n25093), .dout(n25136));
  jand g24968(.dina(n25102), .dinb(n24953), .dout(n25137));
  jnot g24969(.din(n25137), .dout(n25138));
  jand g24970(.dina(n25138), .dinb(n25136), .dout(n25139));
  jnot g24971(.din(n25139), .dout(n25140));
  jand g24972(.dina(n25091), .dinb(n25083), .dout(n25141));
  jnot g24973(.din(n25141), .dout(n25142));
  jnot g24974(.din(n25092), .dout(n25143));
  jor  g24975(.dina(n25143), .dinb(n24957), .dout(n25144));
  jand g24976(.dina(n25144), .dinb(n25142), .dout(n25145));
  jor  g24977(.dina(n25081), .dinb(n25073), .dout(n25146));
  jand g24978(.dina(n25082), .dinb(n24961), .dout(n25147));
  jnot g24979(.din(n25147), .dout(n25148));
  jand g24980(.dina(n25148), .dinb(n25146), .dout(n25149));
  jand g24981(.dina(n25071), .dinb(n25063), .dout(n25150));
  jnot g24982(.din(n25150), .dout(n25151));
  jnot g24983(.din(n25072), .dout(n25152));
  jor  g24984(.dina(n25152), .dinb(n24966), .dout(n25153));
  jand g24985(.dina(n25153), .dinb(n25151), .dout(n25154));
  jor  g24986(.dina(n25061), .dinb(n25053), .dout(n25155));
  jand g24987(.dina(n25062), .dinb(n24970), .dout(n25156));
  jnot g24988(.din(n25156), .dout(n25157));
  jand g24989(.dina(n25157), .dinb(n25155), .dout(n25158));
  jor  g24990(.dina(n25050), .dinb(n25042), .dout(n25159));
  jand g24991(.dina(n25051), .dinb(n24975), .dout(n25160));
  jnot g24992(.din(n25160), .dout(n25161));
  jand g24993(.dina(n25161), .dinb(n25159), .dout(n25162));
  jor  g24994(.dina(n25039), .dinb(n25031), .dout(n25163));
  jand g24995(.dina(n25040), .dinb(n24980), .dout(n25164));
  jnot g24996(.din(n25164), .dout(n25165));
  jand g24997(.dina(n25165), .dinb(n25163), .dout(n25166));
  jor  g24998(.dina(n25028), .dinb(n25020), .dout(n25167));
  jand g24999(.dina(n25029), .dinb(n24985), .dout(n25168));
  jnot g25000(.din(n25168), .dout(n25169));
  jand g25001(.dina(n25169), .dinb(n25167), .dout(n25170));
  jand g25002(.dina(n25017), .dinb(n25010), .dout(n25171));
  jand g25003(.dina(n25018), .dinb(n24988), .dout(n25172));
  jor  g25004(.dina(n25172), .dinb(n25171), .dout(n25173));
  jand g25005(.dina(n18514), .dinb(n5076), .dout(n25174));
  jand g25006(.dina(n18293), .dinb(n5084), .dout(n25175));
  jand g25007(.dina(n17942), .dinb(n5082), .dout(n25176));
  jand g25008(.dina(n17535), .dinb(n6050), .dout(n25177));
  jor  g25009(.dina(n25177), .dinb(n25176), .dout(n25178));
  jor  g25010(.dina(n25178), .dinb(n25175), .dout(n25179));
  jor  g25011(.dina(n25179), .dinb(n25174), .dout(n25180));
  jand g25012(.dina(n21241), .dinb(n7272), .dout(n25181));
  jand g25013(.dina(n1713), .dinb(n1053), .dout(n25182));
  jand g25014(.dina(n25182), .dinb(n993), .dout(n25183));
  jand g25015(.dina(n25183), .dinb(n880), .dout(n25184));
  jand g25016(.dina(n25184), .dinb(n630), .dout(n25185));
  jand g25017(.dina(n1376), .dinb(n583), .dout(n25186));
  jand g25018(.dina(n25186), .dinb(n2377), .dout(n25187));
  jand g25019(.dina(n25187), .dinb(n7103), .dout(n25188));
  jand g25020(.dina(n2522), .dinb(n1512), .dout(n25189));
  jand g25021(.dina(n25189), .dinb(n19115), .dout(n25190));
  jand g25022(.dina(n25190), .dinb(n21135), .dout(n25191));
  jand g25023(.dina(n25191), .dinb(n25188), .dout(n25192));
  jand g25024(.dina(n25192), .dinb(n25185), .dout(n25193));
  jand g25025(.dina(n25193), .dinb(n25181), .dout(n25194));
  jand g25026(.dina(n25194), .dinb(n6248), .dout(n25195));
  jand g25027(.dina(n2712), .dinb(n1484), .dout(n25196));
  jand g25028(.dina(n25196), .dinb(n25195), .dout(n25197));
  jnot g25029(.din(n25197), .dout(n25198));
  jxor g25030(.dina(n24928), .dinb(n24926), .dout(n25199));
  jor  g25031(.dina(n25199), .dinb(\a[2] ), .dout(n25200));
  jor  g25032(.dina(n24930), .dinb(n17779), .dout(n25201));
  jand g25033(.dina(n25201), .dinb(n25200), .dout(n25202));
  jxor g25034(.dina(n25202), .dinb(n25198), .dout(n25203));
  jxor g25035(.dina(n25203), .dinb(n25180), .dout(n25204));
  jxor g25036(.dina(n25204), .dinb(n25173), .dout(n25205));
  jnot g25037(.din(n18916), .dout(n25206));
  jor  g25038(.dina(n25206), .dinb(n4343), .dout(n25207));
  jnot g25039(.din(n18488), .dout(n25208));
  jor  g25040(.dina(n25208), .dinb(n4346), .dout(n25209));
  jnot g25041(.din(n18914), .dout(n25210));
  jor  g25042(.dina(n25210), .dinb(n4348), .dout(n25211));
  jand g25043(.dina(n25211), .dinb(n25209), .dout(n25212));
  jor  g25044(.dina(n23383), .dinb(n3683), .dout(n25213));
  jand g25045(.dina(n25213), .dinb(n25212), .dout(n25214));
  jand g25046(.dina(n25214), .dinb(n25207), .dout(n25215));
  jxor g25047(.dina(n25215), .dinb(\a[29] ), .dout(n25216));
  jnot g25048(.din(n25216), .dout(n25217));
  jxor g25049(.dina(n25217), .dinb(n25205), .dout(n25218));
  jxor g25050(.dina(n25218), .dinb(n25170), .dout(n25219));
  jand g25051(.dina(n19375), .dinb(n71), .dout(n25220));
  jand g25052(.dina(n19219), .dinb(n731), .dout(n25221));
  jand g25053(.dina(n19373), .dinb(n796), .dout(n25222));
  jor  g25054(.dina(n25222), .dinb(n25221), .dout(n25223));
  jand g25055(.dina(n19220), .dinb(n1806), .dout(n25224));
  jor  g25056(.dina(n25224), .dinb(n25223), .dout(n25225));
  jor  g25057(.dina(n25225), .dinb(n25220), .dout(n25226));
  jxor g25058(.dina(n25226), .dinb(n77), .dout(n25227));
  jxor g25059(.dina(n25227), .dinb(n25219), .dout(n25228));
  jxor g25060(.dina(n25228), .dinb(n25166), .dout(n25229));
  jand g25061(.dina(n20358), .dinb(n806), .dout(n25230));
  jand g25062(.dina(n20204), .dinb(n1620), .dout(n25231));
  jand g25063(.dina(n20205), .dinb(n1612), .dout(n25232));
  jand g25064(.dina(n19922), .dinb(n1644), .dout(n25233));
  jor  g25065(.dina(n25233), .dinb(n25232), .dout(n25234));
  jor  g25066(.dina(n25234), .dinb(n25231), .dout(n25235));
  jor  g25067(.dina(n25235), .dinb(n25230), .dout(n25236));
  jxor g25068(.dina(n25236), .dinb(n65), .dout(n25237));
  jxor g25069(.dina(n25237), .dinb(n25229), .dout(n25238));
  jxor g25070(.dina(n25238), .dinb(n25162), .dout(n25239));
  jnot g25071(.din(n21367), .dout(n25240));
  jor  g25072(.dina(n25240), .dinb(n1820), .dout(n25241));
  jor  g25073(.dina(n23252), .dinb(n2189), .dout(n25242));
  jor  g25074(.dina(n23268), .dinb(n2181), .dout(n25243));
  jnot g25075(.din(n20344), .dout(n25244));
  jor  g25076(.dina(n25244), .dinb(n2186), .dout(n25245));
  jand g25077(.dina(n25245), .dinb(n25243), .dout(n25246));
  jand g25078(.dina(n25246), .dinb(n25242), .dout(n25247));
  jand g25079(.dina(n25247), .dinb(n25241), .dout(n25248));
  jxor g25080(.dina(n25248), .dinb(\a[20] ), .dout(n25249));
  jxor g25081(.dina(n25249), .dinb(n25239), .dout(n25250));
  jxor g25082(.dina(n25250), .dinb(n25158), .dout(n25251));
  jor  g25083(.dina(n23220), .dinb(n2744), .dout(n25252));
  jor  g25084(.dina(n23222), .dinb(n2753), .dout(n25253));
  jor  g25085(.dina(n23224), .dinb(n2749), .dout(n25254));
  jor  g25086(.dina(n23226), .dinb(n2758), .dout(n25255));
  jand g25087(.dina(n25255), .dinb(n25254), .dout(n25256));
  jand g25088(.dina(n25256), .dinb(n25253), .dout(n25257));
  jand g25089(.dina(n25257), .dinb(n25252), .dout(n25258));
  jxor g25090(.dina(n25258), .dinb(\a[17] ), .dout(n25259));
  jxor g25091(.dina(n25259), .dinb(n25251), .dout(n25260));
  jxor g25092(.dina(n25260), .dinb(n25154), .dout(n25261));
  jand g25093(.dina(n22267), .dinb(n3423), .dout(n25262));
  jand g25094(.dina(n22265), .dinb(n3569), .dout(n25263));
  jand g25095(.dina(n22163), .dinb(n3428), .dout(n25264));
  jand g25096(.dina(n22164), .dinb(n3210), .dout(n25265));
  jor  g25097(.dina(n25265), .dinb(n25264), .dout(n25266));
  jor  g25098(.dina(n25266), .dinb(n25263), .dout(n25267));
  jor  g25099(.dina(n25267), .dinb(n25262), .dout(n25268));
  jxor g25100(.dina(n25268), .dinb(n3473), .dout(n25269));
  jxor g25101(.dina(n25269), .dinb(n25261), .dout(n25270));
  jxor g25102(.dina(n25270), .dinb(n25149), .dout(n25271));
  jnot g25103(.din(n23159), .dout(n25272));
  jor  g25104(.dina(n25272), .dinb(n4023), .dout(n25273));
  jnot g25105(.din(n23079), .dout(n25274));
  jor  g25106(.dina(n25274), .dinb(n4025), .dout(n25275));
  jnot g25107(.din(n23080), .dout(n25276));
  jor  g25108(.dina(n25276), .dinb(n4028), .dout(n25277));
  jnot g25109(.din(n22937), .dout(n25278));
  jor  g25110(.dina(n25278), .dinb(n3871), .dout(n25279));
  jand g25111(.dina(n25279), .dinb(n25277), .dout(n25280));
  jand g25112(.dina(n25280), .dinb(n25275), .dout(n25281));
  jand g25113(.dina(n25281), .dinb(n25273), .dout(n25282));
  jxor g25114(.dina(n25282), .dinb(\a[11] ), .dout(n25283));
  jxor g25115(.dina(n25283), .dinb(n25271), .dout(n25284));
  jxor g25116(.dina(n25284), .dinb(n25145), .dout(n25285));
  jnot g25117(.din(n24077), .dout(n25286));
  jor  g25118(.dina(n25286), .dinb(n4692), .dout(n25287));
  jor  g25119(.dina(n24266), .dinb(n4705), .dout(n25288));
  jor  g25120(.dina(n24265), .dinb(n4697), .dout(n25289));
  jnot g25121(.din(n23144), .dout(n25290));
  jor  g25122(.dina(n25290), .dinb(n4702), .dout(n25291));
  jand g25123(.dina(n25291), .dinb(n25289), .dout(n25292));
  jand g25124(.dina(n25292), .dinb(n25288), .dout(n25293));
  jand g25125(.dina(n25293), .dinb(n25287), .dout(n25294));
  jxor g25126(.dina(n25294), .dinb(\a[8] ), .dout(n25295));
  jxor g25127(.dina(n25295), .dinb(n25285), .dout(n25296));
  jxor g25128(.dina(n25296), .dinb(n25140), .dout(n25297));
  jor  g25129(.dina(n24736), .dinb(n5281), .dout(n25298));
  jor  g25130(.dina(n24738), .dinb(n5539), .dout(n25299));
  jor  g25131(.dina(n24518), .dinb(n5532), .dout(n25300));
  jor  g25132(.dina(n24304), .dinb(n5537), .dout(n25301));
  jand g25133(.dina(n25301), .dinb(n25300), .dout(n25302));
  jand g25134(.dina(n25302), .dinb(n25299), .dout(n25303));
  jand g25135(.dina(n25303), .dinb(n25298), .dout(n25304));
  jxor g25136(.dina(n25304), .dinb(\a[5] ), .dout(n25305));
  jnot g25137(.din(n25305), .dout(n25306));
  jxor g25138(.dina(n25306), .dinb(n25297), .dout(n25307));
  jxor g25139(.dina(n25307), .dinb(n25135), .dout(n25308));
  jand g25140(.dina(n25123), .dinb(n24949), .dout(n25309));
  jand g25141(.dina(n25127), .dinb(n25124), .dout(n25310));
  jor  g25142(.dina(n25310), .dinb(n25309), .dout(n25311));
  jxor g25143(.dina(n25311), .dinb(n25308), .dout(n25312));
  jxor g25144(.dina(n25312), .dinb(n25130), .dout(\result[7] ));
  jand g25145(.dina(n25312), .dinb(n25130), .dout(n25314));
  jand g25146(.dina(n25296), .dinb(n25140), .dout(n25315));
  jand g25147(.dina(n25306), .dinb(n25297), .dout(n25316));
  jor  g25148(.dina(n25316), .dinb(n25315), .dout(n25317));
  jnot g25149(.din(n25145), .dout(n25318));
  jand g25150(.dina(n25284), .dinb(n25318), .dout(n25319));
  jnot g25151(.din(n25319), .dout(n25320));
  jor  g25152(.dina(n25295), .dinb(n25285), .dout(n25321));
  jand g25153(.dina(n25321), .dinb(n25320), .dout(n25322));
  jnot g25154(.din(n25322), .dout(n25323));
  jnot g25155(.din(n25270), .dout(n25324));
  jor  g25156(.dina(n25324), .dinb(n25149), .dout(n25325));
  jor  g25157(.dina(n25283), .dinb(n25271), .dout(n25326));
  jand g25158(.dina(n25326), .dinb(n25325), .dout(n25327));
  jnot g25159(.din(n25260), .dout(n25328));
  jor  g25160(.dina(n25328), .dinb(n25154), .dout(n25329));
  jor  g25161(.dina(n25269), .dinb(n25261), .dout(n25330));
  jand g25162(.dina(n25330), .dinb(n25329), .dout(n25331));
  jnot g25163(.din(n25250), .dout(n25332));
  jor  g25164(.dina(n25332), .dinb(n25158), .dout(n25333));
  jor  g25165(.dina(n25259), .dinb(n25251), .dout(n25334));
  jand g25166(.dina(n25334), .dinb(n25333), .dout(n25335));
  jnot g25167(.din(n25238), .dout(n25336));
  jor  g25168(.dina(n25336), .dinb(n25162), .dout(n25337));
  jor  g25169(.dina(n25249), .dinb(n25239), .dout(n25338));
  jand g25170(.dina(n25338), .dinb(n25337), .dout(n25339));
  jnot g25171(.din(n25228), .dout(n25340));
  jor  g25172(.dina(n25340), .dinb(n25166), .dout(n25341));
  jor  g25173(.dina(n25237), .dinb(n25229), .dout(n25342));
  jand g25174(.dina(n25342), .dinb(n25341), .dout(n25343));
  jnot g25175(.din(n25218), .dout(n25344));
  jor  g25176(.dina(n25344), .dinb(n25170), .dout(n25345));
  jor  g25177(.dina(n25227), .dinb(n25219), .dout(n25346));
  jand g25178(.dina(n25346), .dinb(n25345), .dout(n25347));
  jand g25179(.dina(n25204), .dinb(n25173), .dout(n25348));
  jand g25180(.dina(n25217), .dinb(n25205), .dout(n25349));
  jor  g25181(.dina(n25349), .dinb(n25348), .dout(n25350));
  jand g25182(.dina(n18502), .dinb(n5076), .dout(n25351));
  jand g25183(.dina(n18292), .dinb(n5084), .dout(n25352));
  jand g25184(.dina(n18293), .dinb(n5082), .dout(n25353));
  jand g25185(.dina(n17942), .dinb(n6050), .dout(n25354));
  jor  g25186(.dina(n25354), .dinb(n25353), .dout(n25355));
  jor  g25187(.dina(n25355), .dinb(n25352), .dout(n25356));
  jor  g25188(.dina(n25356), .dinb(n25351), .dout(n25357));
  jand g25189(.dina(n20717), .dinb(n1098), .dout(n25358));
  jand g25190(.dina(n7082), .dinb(n1037), .dout(n25359));
  jand g25191(.dina(n25359), .dinb(n25358), .dout(n25360));
  jand g25192(.dina(n25360), .dinb(n2655), .dout(n25361));
  jand g25193(.dina(n3814), .dinb(n2086), .dout(n25362));
  jand g25194(.dina(n25362), .dinb(n698), .dout(n25363));
  jand g25195(.dina(n25363), .dinb(n25361), .dout(n25364));
  jand g25196(.dina(n5395), .dinb(n4588), .dout(n25365));
  jand g25197(.dina(n9545), .dinb(n622), .dout(n25366));
  jand g25198(.dina(n25366), .dinb(n25365), .dout(n25367));
  jand g25199(.dina(n1767), .dinb(n1485), .dout(n25368));
  jand g25200(.dina(n15119), .dinb(n1247), .dout(n25369));
  jand g25201(.dina(n988), .dinb(n1378), .dout(n25370));
  jand g25202(.dina(n25370), .dinb(n1270), .dout(n25371));
  jand g25203(.dina(n25371), .dinb(n25369), .dout(n25372));
  jand g25204(.dina(n25372), .dinb(n25368), .dout(n25373));
  jand g25205(.dina(n25373), .dinb(n25367), .dout(n25374));
  jand g25206(.dina(n25374), .dinb(n25364), .dout(n25375));
  jand g25207(.dina(n25375), .dinb(n14070), .dout(n25376));
  jand g25208(.dina(n25376), .dinb(n2356), .dout(n25377));
  jnot g25209(.din(n25377), .dout(n25378));
  jxor g25210(.dina(n25378), .dinb(n25202), .dout(n25379));
  jor  g25211(.dina(n25202), .dinb(n25198), .dout(n25380));
  jand g25212(.dina(n25202), .dinb(n25198), .dout(n25381));
  jor  g25213(.dina(n25381), .dinb(n25180), .dout(n25382));
  jand g25214(.dina(n25382), .dinb(n25380), .dout(n25383));
  jxor g25215(.dina(n25383), .dinb(n25379), .dout(n25384));
  jxor g25216(.dina(n25384), .dinb(n25357), .dout(n25385));
  jxor g25217(.dina(n25385), .dinb(n25350), .dout(n25386));
  jand g25218(.dina(n19399), .dinb(n2936), .dout(n25387));
  jand g25219(.dina(n18914), .dinb(n2940), .dout(n25388));
  jand g25220(.dina(n19220), .dinb(n2943), .dout(n25389));
  jor  g25221(.dina(n25389), .dinb(n25388), .dout(n25390));
  jand g25222(.dina(n18488), .dinb(n3684), .dout(n25391));
  jor  g25223(.dina(n25391), .dinb(n25390), .dout(n25392));
  jor  g25224(.dina(n25392), .dinb(n25387), .dout(n25393));
  jxor g25225(.dina(n25393), .dinb(n93), .dout(n25394));
  jxor g25226(.dina(n25394), .dinb(n25386), .dout(n25395));
  jnot g25227(.din(n19924), .dout(n25396));
  jor  g25228(.dina(n25396), .dinb(n2303), .dout(n25397));
  jnot g25229(.din(n19922), .dout(n25398));
  jor  g25230(.dina(n25398), .dinb(n2309), .dout(n25399));
  jnot g25231(.din(n19373), .dout(n25400));
  jor  g25232(.dina(n25400), .dinb(n2306), .dout(n25401));
  jnot g25233(.din(n19219), .dout(n25402));
  jor  g25234(.dina(n25402), .dinb(n1805), .dout(n25403));
  jand g25235(.dina(n25403), .dinb(n25401), .dout(n25404));
  jand g25236(.dina(n25404), .dinb(n25399), .dout(n25405));
  jand g25237(.dina(n25405), .dinb(n25397), .dout(n25406));
  jxor g25238(.dina(n25406), .dinb(\a[26] ), .dout(n25407));
  jxor g25239(.dina(n25407), .dinb(n25395), .dout(n25408));
  jxor g25240(.dina(n25408), .dinb(n25347), .dout(n25409));
  jnot g25241(.din(n20346), .dout(n25410));
  jor  g25242(.dina(n25410), .dinb(n807), .dout(n25411));
  jor  g25243(.dina(n25244), .dinb(n1621), .dout(n25412));
  jnot g25244(.din(n20204), .dout(n25413));
  jor  g25245(.dina(n25413), .dinb(n1613), .dout(n25414));
  jnot g25246(.din(n20205), .dout(n25415));
  jor  g25247(.dina(n25415), .dinb(n1617), .dout(n25416));
  jand g25248(.dina(n25416), .dinb(n25414), .dout(n25417));
  jand g25249(.dina(n25417), .dinb(n25412), .dout(n25418));
  jand g25250(.dina(n25418), .dinb(n25411), .dout(n25419));
  jxor g25251(.dina(n25419), .dinb(\a[23] ), .dout(n25420));
  jxor g25252(.dina(n25420), .dinb(n25409), .dout(n25421));
  jxor g25253(.dina(n25421), .dinb(n25343), .dout(n25422));
  jand g25254(.dina(n21355), .dinb(n1819), .dout(n25423));
  jand g25255(.dina(n21198), .dinb(n2180), .dout(n25424));
  jand g25256(.dina(n21197), .dinb(n2243), .dout(n25425));
  jor  g25257(.dina(n25425), .dinb(n25424), .dout(n25426));
  jand g25258(.dina(n20947), .dinb(n2185), .dout(n25427));
  jor  g25259(.dina(n25427), .dinb(n25426), .dout(n25428));
  jor  g25260(.dina(n25428), .dinb(n25423), .dout(n25429));
  jxor g25261(.dina(n25429), .dinb(n2196), .dout(n25430));
  jxor g25262(.dina(n25430), .dinb(n25422), .dout(n25431));
  jxor g25263(.dina(n25431), .dinb(n25339), .dout(n25432));
  jnot g25264(.din(n22291), .dout(n25433));
  jor  g25265(.dina(n25433), .dinb(n2744), .dout(n25434));
  jnot g25266(.din(n22164), .dout(n25435));
  jor  g25267(.dina(n25435), .dinb(n2753), .dout(n25436));
  jor  g25268(.dina(n23222), .dinb(n2749), .dout(n25437));
  jor  g25269(.dina(n23224), .dinb(n2758), .dout(n25438));
  jand g25270(.dina(n25438), .dinb(n25437), .dout(n25439));
  jand g25271(.dina(n25439), .dinb(n25436), .dout(n25440));
  jand g25272(.dina(n25440), .dinb(n25434), .dout(n25441));
  jxor g25273(.dina(n25441), .dinb(\a[17] ), .dout(n25442));
  jxor g25274(.dina(n25442), .dinb(n25432), .dout(n25443));
  jxor g25275(.dina(n25443), .dinb(n25335), .dout(n25444));
  jnot g25276(.din(n22939), .dout(n25445));
  jor  g25277(.dina(n25445), .dinb(n3424), .dout(n25446));
  jnot g25278(.din(n22265), .dout(n25447));
  jor  g25279(.dina(n25447), .dinb(n3429), .dout(n25448));
  jor  g25280(.dina(n25278), .dinb(n3426), .dout(n25449));
  jand g25281(.dina(n25449), .dinb(n25448), .dout(n25450));
  jnot g25282(.din(n22163), .dout(n25451));
  jor  g25283(.dina(n25451), .dinb(n3211), .dout(n25452));
  jand g25284(.dina(n25452), .dinb(n25450), .dout(n25453));
  jand g25285(.dina(n25453), .dinb(n25446), .dout(n25454));
  jxor g25286(.dina(n25454), .dinb(\a[14] ), .dout(n25455));
  jxor g25287(.dina(n25455), .dinb(n25444), .dout(n25456));
  jxor g25288(.dina(n25456), .dinb(n25331), .dout(n25457));
  jnot g25289(.din(n23146), .dout(n25458));
  jor  g25290(.dina(n25458), .dinb(n4023), .dout(n25459));
  jor  g25291(.dina(n25290), .dinb(n4025), .dout(n25460));
  jor  g25292(.dina(n25274), .dinb(n4028), .dout(n25461));
  jor  g25293(.dina(n25276), .dinb(n3871), .dout(n25462));
  jand g25294(.dina(n25462), .dinb(n25461), .dout(n25463));
  jand g25295(.dina(n25463), .dinb(n25460), .dout(n25464));
  jand g25296(.dina(n25464), .dinb(n25459), .dout(n25465));
  jxor g25297(.dina(n25465), .dinb(\a[11] ), .dout(n25466));
  jxor g25298(.dina(n25466), .dinb(n25457), .dout(n25467));
  jxor g25299(.dina(n25467), .dinb(n25327), .dout(n25468));
  jor  g25300(.dina(n24302), .dinb(n4692), .dout(n25469));
  jor  g25301(.dina(n24304), .dinb(n4705), .dout(n25470));
  jor  g25302(.dina(n24265), .dinb(n4702), .dout(n25471));
  jor  g25303(.dina(n24266), .dinb(n4697), .dout(n25472));
  jand g25304(.dina(n25472), .dinb(n25471), .dout(n25473));
  jand g25305(.dina(n25473), .dinb(n25470), .dout(n25474));
  jand g25306(.dina(n25474), .dinb(n25469), .dout(n25475));
  jxor g25307(.dina(n25475), .dinb(\a[8] ), .dout(n25476));
  jxor g25308(.dina(n25476), .dinb(n25468), .dout(n25477));
  jxor g25309(.dina(n25477), .dinb(n25323), .dout(n25478));
  jor  g25310(.dina(n24932), .dinb(n5281), .dout(n25479));
  jor  g25311(.dina(n24930), .dinb(n5539), .dout(n25480));
  jor  g25312(.dina(n24738), .dinb(n5532), .dout(n25481));
  jor  g25313(.dina(n24518), .dinb(n5537), .dout(n25482));
  jand g25314(.dina(n25482), .dinb(n25481), .dout(n25483));
  jand g25315(.dina(n25483), .dinb(n25480), .dout(n25484));
  jand g25316(.dina(n25484), .dinb(n25479), .dout(n25485));
  jxor g25317(.dina(n25485), .dinb(\a[5] ), .dout(n25486));
  jnot g25318(.din(n25486), .dout(n25487));
  jxor g25319(.dina(n25487), .dinb(n25478), .dout(n25488));
  jxor g25320(.dina(n25488), .dinb(n25317), .dout(n25489));
  jand g25321(.dina(n25307), .dinb(n25135), .dout(n25490));
  jand g25322(.dina(n25311), .dinb(n25308), .dout(n25491));
  jor  g25323(.dina(n25491), .dinb(n25490), .dout(n25492));
  jxor g25324(.dina(n25492), .dinb(n25489), .dout(n25493));
  jxor g25325(.dina(n25493), .dinb(n25314), .dout(\result[8] ));
  jand g25326(.dina(n25493), .dinb(n25314), .dout(n25495));
  jand g25327(.dina(n25477), .dinb(n25323), .dout(n25496));
  jand g25328(.dina(n25487), .dinb(n25478), .dout(n25497));
  jor  g25329(.dina(n25497), .dinb(n25496), .dout(n25498));
  jnot g25330(.din(n25327), .dout(n25499));
  jand g25331(.dina(n25467), .dinb(n25499), .dout(n25500));
  jnot g25332(.din(n25500), .dout(n25501));
  jor  g25333(.dina(n25476), .dinb(n25468), .dout(n25502));
  jand g25334(.dina(n25502), .dinb(n25501), .dout(n25503));
  jor  g25335(.dina(n25116), .dinb(n5281), .dout(n25504));
  jor  g25336(.dina(n24930), .dinb(n17966), .dout(n25505));
  jor  g25337(.dina(n24738), .dinb(n5537), .dout(n25506));
  jand g25338(.dina(n25506), .dinb(n25505), .dout(n25507));
  jand g25339(.dina(n25507), .dinb(n25504), .dout(n25508));
  jxor g25340(.dina(n25508), .dinb(\a[5] ), .dout(n25509));
  jxor g25341(.dina(n25509), .dinb(n25503), .dout(n25510));
  jnot g25342(.din(n25456), .dout(n25511));
  jor  g25343(.dina(n25511), .dinb(n25331), .dout(n25512));
  jor  g25344(.dina(n25466), .dinb(n25457), .dout(n25513));
  jand g25345(.dina(n25513), .dinb(n25512), .dout(n25514));
  jnot g25346(.din(n25335), .dout(n25515));
  jand g25347(.dina(n25443), .dinb(n25515), .dout(n25516));
  jnot g25348(.din(n25516), .dout(n25517));
  jor  g25349(.dina(n25455), .dinb(n25444), .dout(n25518));
  jand g25350(.dina(n25518), .dinb(n25517), .dout(n25519));
  jnot g25351(.din(n25339), .dout(n25520));
  jand g25352(.dina(n25431), .dinb(n25520), .dout(n25521));
  jnot g25353(.din(n25521), .dout(n25522));
  jor  g25354(.dina(n25442), .dinb(n25432), .dout(n25523));
  jand g25355(.dina(n25523), .dinb(n25522), .dout(n25524));
  jnot g25356(.din(n25421), .dout(n25525));
  jor  g25357(.dina(n25525), .dinb(n25343), .dout(n25526));
  jor  g25358(.dina(n25430), .dinb(n25422), .dout(n25527));
  jand g25359(.dina(n25527), .dinb(n25526), .dout(n25528));
  jnot g25360(.din(n25408), .dout(n25529));
  jor  g25361(.dina(n25529), .dinb(n25347), .dout(n25530));
  jor  g25362(.dina(n25420), .dinb(n25409), .dout(n25531));
  jand g25363(.dina(n25531), .dinb(n25530), .dout(n25532));
  jnot g25364(.din(n25386), .dout(n25533));
  jor  g25365(.dina(n25394), .dinb(n25533), .dout(n25534));
  jor  g25366(.dina(n25407), .dinb(n25395), .dout(n25535));
  jand g25367(.dina(n25535), .dinb(n25534), .dout(n25536));
  jand g25368(.dina(n25384), .dinb(n25357), .dout(n25537));
  jand g25369(.dina(n25385), .dinb(n25350), .dout(n25538));
  jor  g25370(.dina(n25538), .dinb(n25537), .dout(n25539));
  jand g25371(.dina(n18490), .dinb(n5076), .dout(n25540));
  jand g25372(.dina(n18488), .dinb(n5084), .dout(n25541));
  jand g25373(.dina(n18292), .dinb(n5082), .dout(n25542));
  jand g25374(.dina(n18293), .dinb(n6050), .dout(n25543));
  jor  g25375(.dina(n25543), .dinb(n25542), .dout(n25544));
  jor  g25376(.dina(n25544), .dinb(n25541), .dout(n25545));
  jor  g25377(.dina(n25545), .dinb(n25540), .dout(n25546));
  jand g25378(.dina(n25378), .dinb(n25202), .dout(n25547));
  jand g25379(.dina(n25383), .dinb(n25379), .dout(n25548));
  jor  g25380(.dina(n25548), .dinb(n25547), .dout(n25549));
  jnot g25381(.din(n25202), .dout(n25550));
  jand g25382(.dina(n13405), .dinb(n704), .dout(n25551));
  jand g25383(.dina(n17825), .dinb(n584), .dout(n25552));
  jand g25384(.dina(n25552), .dinb(n25551), .dout(n25553));
  jand g25385(.dina(n3857), .dinb(n1272), .dout(n25554));
  jand g25386(.dina(n1005), .dinb(n1708), .dout(n25555));
  jand g25387(.dina(n1351), .dinb(n1317), .dout(n25556));
  jand g25388(.dina(n25556), .dinb(n25555), .dout(n25557));
  jand g25389(.dina(n25557), .dinb(n586), .dout(n25558));
  jand g25390(.dina(n25558), .dinb(n25554), .dout(n25559));
  jand g25391(.dina(n1514), .dinb(n563), .dout(n25560));
  jand g25392(.dina(n25560), .dinb(n25559), .dout(n25561));
  jand g25393(.dina(n25561), .dinb(n25553), .dout(n25562));
  jand g25394(.dina(n25562), .dinb(n2141), .dout(n25563));
  jand g25395(.dina(n7768), .dinb(n5239), .dout(n25564));
  jand g25396(.dina(n25564), .dinb(n4507), .dout(n25565));
  jand g25397(.dina(n25565), .dinb(n25563), .dout(n25566));
  jxor g25398(.dina(n25566), .dinb(n25550), .dout(n25567));
  jxor g25399(.dina(n25567), .dinb(n25549), .dout(n25568));
  jxor g25400(.dina(n25568), .dinb(n25546), .dout(n25569));
  jxor g25401(.dina(n25569), .dinb(n25539), .dout(n25570));
  jand g25402(.dina(n19387), .dinb(n2936), .dout(n25571));
  jand g25403(.dina(n19219), .dinb(n2943), .dout(n25572));
  jand g25404(.dina(n19220), .dinb(n2940), .dout(n25573));
  jand g25405(.dina(n18914), .dinb(n3684), .dout(n25574));
  jor  g25406(.dina(n25574), .dinb(n25573), .dout(n25575));
  jor  g25407(.dina(n25575), .dinb(n25572), .dout(n25576));
  jor  g25408(.dina(n25576), .dinb(n25571), .dout(n25577));
  jxor g25409(.dina(n25577), .dinb(n93), .dout(n25578));
  jxor g25410(.dina(n25578), .dinb(n25570), .dout(n25579));
  jand g25411(.dina(n20371), .dinb(n71), .dout(n25580));
  jand g25412(.dina(n20205), .dinb(n796), .dout(n25581));
  jand g25413(.dina(n19922), .dinb(n731), .dout(n25582));
  jand g25414(.dina(n19373), .dinb(n1806), .dout(n25583));
  jor  g25415(.dina(n25583), .dinb(n25582), .dout(n25584));
  jor  g25416(.dina(n25584), .dinb(n25581), .dout(n25585));
  jor  g25417(.dina(n25585), .dinb(n25580), .dout(n25586));
  jxor g25418(.dina(n25586), .dinb(n77), .dout(n25587));
  jxor g25419(.dina(n25587), .dinb(n25579), .dout(n25588));
  jxor g25420(.dina(n25588), .dinb(n25536), .dout(n25589));
  jand g25421(.dina(n20949), .dinb(n806), .dout(n25590));
  jand g25422(.dina(n20947), .dinb(n1620), .dout(n25591));
  jand g25423(.dina(n20344), .dinb(n1612), .dout(n25592));
  jand g25424(.dina(n20204), .dinb(n1644), .dout(n25593));
  jor  g25425(.dina(n25593), .dinb(n25592), .dout(n25594));
  jor  g25426(.dina(n25594), .dinb(n25591), .dout(n25595));
  jor  g25427(.dina(n25595), .dinb(n25590), .dout(n25596));
  jxor g25428(.dina(n25596), .dinb(n65), .dout(n25597));
  jxor g25429(.dina(n25597), .dinb(n25589), .dout(n25598));
  jxor g25430(.dina(n25598), .dinb(n25532), .dout(n25599));
  jand g25431(.dina(n21342), .dinb(n1819), .dout(n25600));
  jand g25432(.dina(n21340), .dinb(n2243), .dout(n25601));
  jand g25433(.dina(n21197), .dinb(n2180), .dout(n25602));
  jand g25434(.dina(n21198), .dinb(n2185), .dout(n25603));
  jor  g25435(.dina(n25603), .dinb(n25602), .dout(n25604));
  jor  g25436(.dina(n25604), .dinb(n25601), .dout(n25605));
  jor  g25437(.dina(n25605), .dinb(n25600), .dout(n25606));
  jxor g25438(.dina(n25606), .dinb(n2196), .dout(n25607));
  jxor g25439(.dina(n25607), .dinb(n25599), .dout(n25608));
  jxor g25440(.dina(n25608), .dinb(n25528), .dout(n25609));
  jnot g25441(.din(n22279), .dout(n25610));
  jor  g25442(.dina(n25610), .dinb(n2744), .dout(n25611));
  jor  g25443(.dina(n25451), .dinb(n2753), .dout(n25612));
  jor  g25444(.dina(n25435), .dinb(n2749), .dout(n25613));
  jor  g25445(.dina(n23222), .dinb(n2758), .dout(n25614));
  jand g25446(.dina(n25614), .dinb(n25613), .dout(n25615));
  jand g25447(.dina(n25615), .dinb(n25612), .dout(n25616));
  jand g25448(.dina(n25616), .dinb(n25611), .dout(n25617));
  jxor g25449(.dina(n25617), .dinb(\a[17] ), .dout(n25618));
  jxor g25450(.dina(n25618), .dinb(n25609), .dout(n25619));
  jxor g25451(.dina(n25619), .dinb(n25524), .dout(n25620));
  jand g25452(.dina(n23172), .dinb(n3423), .dout(n25621));
  jand g25453(.dina(n22937), .dinb(n3428), .dout(n25622));
  jand g25454(.dina(n23080), .dinb(n3569), .dout(n25623));
  jor  g25455(.dina(n25623), .dinb(n25622), .dout(n25624));
  jand g25456(.dina(n22265), .dinb(n3210), .dout(n25625));
  jor  g25457(.dina(n25625), .dinb(n25624), .dout(n25626));
  jor  g25458(.dina(n25626), .dinb(n25621), .dout(n25627));
  jxor g25459(.dina(n25627), .dinb(n3473), .dout(n25628));
  jxor g25460(.dina(n25628), .dinb(n25620), .dout(n25629));
  jxor g25461(.dina(n25629), .dinb(n25519), .dout(n25630));
  jnot g25462(.din(n23847), .dout(n25631));
  jor  g25463(.dina(n25631), .dinb(n4023), .dout(n25632));
  jor  g25464(.dina(n24265), .dinb(n4025), .dout(n25633));
  jor  g25465(.dina(n25290), .dinb(n4028), .dout(n25634));
  jor  g25466(.dina(n25274), .dinb(n3871), .dout(n25635));
  jand g25467(.dina(n25635), .dinb(n25634), .dout(n25636));
  jand g25468(.dina(n25636), .dinb(n25633), .dout(n25637));
  jand g25469(.dina(n25637), .dinb(n25632), .dout(n25638));
  jxor g25470(.dina(n25638), .dinb(\a[11] ), .dout(n25639));
  jxor g25471(.dina(n25639), .dinb(n25630), .dout(n25640));
  jxor g25472(.dina(n25640), .dinb(n25514), .dout(n25641));
  jor  g25473(.dina(n24516), .dinb(n4692), .dout(n25642));
  jor  g25474(.dina(n24304), .dinb(n4697), .dout(n25643));
  jor  g25475(.dina(n24518), .dinb(n4705), .dout(n25644));
  jand g25476(.dina(n25644), .dinb(n25643), .dout(n25645));
  jor  g25477(.dina(n24266), .dinb(n4702), .dout(n25646));
  jand g25478(.dina(n25646), .dinb(n25645), .dout(n25647));
  jand g25479(.dina(n25647), .dinb(n25642), .dout(n25648));
  jxor g25480(.dina(n25648), .dinb(\a[8] ), .dout(n25649));
  jxor g25481(.dina(n25649), .dinb(n25641), .dout(n25650));
  jxor g25482(.dina(n25650), .dinb(n25510), .dout(n25651));
  jxor g25483(.dina(n25651), .dinb(n25498), .dout(n25652));
  jand g25484(.dina(n25488), .dinb(n25317), .dout(n25653));
  jand g25485(.dina(n25492), .dinb(n25489), .dout(n25654));
  jor  g25486(.dina(n25654), .dinb(n25653), .dout(n25655));
  jxor g25487(.dina(n25655), .dinb(n25652), .dout(n25656));
  jxor g25488(.dina(n25656), .dinb(n25495), .dout(\result[9] ));
  jand g25489(.dina(n25656), .dinb(n25495), .dout(n25658));
  jand g25490(.dina(n25651), .dinb(n25498), .dout(n25659));
  jand g25491(.dina(n25655), .dinb(n25652), .dout(n25660));
  jor  g25492(.dina(n25660), .dinb(n25659), .dout(n25661));
  jor  g25493(.dina(n25509), .dinb(n25503), .dout(n25662));
  jnot g25494(.din(n25662), .dout(n25663));
  jand g25495(.dina(n25650), .dinb(n25510), .dout(n25664));
  jor  g25496(.dina(n25664), .dinb(n25663), .dout(n25665));
  jnot g25497(.din(n25519), .dout(n25666));
  jand g25498(.dina(n25629), .dinb(n25666), .dout(n25667));
  jnot g25499(.din(n25667), .dout(n25668));
  jor  g25500(.dina(n25639), .dinb(n25630), .dout(n25669));
  jand g25501(.dina(n25669), .dinb(n25668), .dout(n25670));
  jnot g25502(.din(n25670), .dout(n25671));
  jnot g25503(.din(n25608), .dout(n25672));
  jor  g25504(.dina(n25672), .dinb(n25528), .dout(n25673));
  jor  g25505(.dina(n25618), .dinb(n25609), .dout(n25674));
  jand g25506(.dina(n25674), .dinb(n25673), .dout(n25675));
  jnot g25507(.din(n25598), .dout(n25676));
  jor  g25508(.dina(n25676), .dinb(n25532), .dout(n25677));
  jor  g25509(.dina(n25607), .dinb(n25599), .dout(n25678));
  jand g25510(.dina(n25678), .dinb(n25677), .dout(n25679));
  jnot g25511(.din(n25588), .dout(n25680));
  jor  g25512(.dina(n25680), .dinb(n25536), .dout(n25681));
  jor  g25513(.dina(n25597), .dinb(n25589), .dout(n25682));
  jand g25514(.dina(n25682), .dinb(n25681), .dout(n25683));
  jnot g25515(.din(n25570), .dout(n25684));
  jor  g25516(.dina(n25578), .dinb(n25684), .dout(n25685));
  jor  g25517(.dina(n25587), .dinb(n25579), .dout(n25686));
  jand g25518(.dina(n25686), .dinb(n25685), .dout(n25687));
  jnot g25519(.din(n25546), .dout(n25688));
  jnot g25520(.din(n25568), .dout(n25689));
  jor  g25521(.dina(n25689), .dinb(n25688), .dout(n25690));
  jnot g25522(.din(n25539), .dout(n25691));
  jnot g25523(.din(n25569), .dout(n25692));
  jor  g25524(.dina(n25692), .dinb(n25691), .dout(n25693));
  jand g25525(.dina(n25693), .dinb(n25690), .dout(n25694));
  jand g25526(.dina(n18916), .dinb(n5076), .dout(n25695));
  jand g25527(.dina(n18914), .dinb(n5084), .dout(n25696));
  jand g25528(.dina(n18488), .dinb(n5082), .dout(n25697));
  jand g25529(.dina(n18292), .dinb(n6050), .dout(n25698));
  jor  g25530(.dina(n25698), .dinb(n25697), .dout(n25699));
  jor  g25531(.dina(n25699), .dinb(n25696), .dout(n25700));
  jor  g25532(.dina(n25700), .dinb(n25695), .dout(n25701));
  jor  g25533(.dina(n25566), .dinb(n25550), .dout(n25702));
  jnot g25534(.din(n25702), .dout(n25703));
  jand g25535(.dina(n25567), .dinb(n25549), .dout(n25704));
  jor  g25536(.dina(n25704), .dinb(n25703), .dout(n25705));
  jand g25537(.dina(n20264), .dinb(n641), .dout(n25706));
  jand g25538(.dina(n562), .dinb(n542), .dout(n25707));
  jand g25539(.dina(n25707), .dinb(n6439), .dout(n25708));
  jand g25540(.dina(n25708), .dinb(n1477), .dout(n25709));
  jand g25541(.dina(n25709), .dinb(n514), .dout(n25710));
  jand g25542(.dina(n25710), .dinb(n25706), .dout(n25711));
  jand g25543(.dina(n3996), .dinb(n1735), .dout(n25712));
  jand g25544(.dina(n25712), .dinb(n9132), .dout(n25713));
  jand g25545(.dina(n8370), .dinb(n3405), .dout(n25714));
  jand g25546(.dina(n25714), .dinb(n25713), .dout(n25715));
  jand g25547(.dina(n25715), .dinb(n1891), .dout(n25716));
  jand g25548(.dina(n25716), .dinb(n25711), .dout(n25717));
  jand g25549(.dina(n19707), .dinb(n13320), .dout(n25718));
  jand g25550(.dina(n25718), .dinb(n25717), .dout(n25719));
  jand g25551(.dina(n25719), .dinb(n3013), .dout(n25720));
  jxor g25552(.dina(n25720), .dinb(n25202), .dout(n25721));
  jand g25553(.dina(n25199), .dinb(n18199), .dout(n25722));
  jxor g25554(.dina(n25722), .dinb(n5277), .dout(n25723));
  jxor g25555(.dina(n25723), .dinb(n25721), .dout(n25724));
  jxor g25556(.dina(n25724), .dinb(n25705), .dout(n25725));
  jxor g25557(.dina(n25725), .dinb(n25701), .dout(n25726));
  jnot g25558(.din(n25726), .dout(n25727));
  jxor g25559(.dina(n25727), .dinb(n25694), .dout(n25728));
  jand g25560(.dina(n19375), .dinb(n2936), .dout(n25729));
  jand g25561(.dina(n19219), .dinb(n2940), .dout(n25730));
  jand g25562(.dina(n19373), .dinb(n2943), .dout(n25731));
  jor  g25563(.dina(n25731), .dinb(n25730), .dout(n25732));
  jand g25564(.dina(n19220), .dinb(n3684), .dout(n25733));
  jor  g25565(.dina(n25733), .dinb(n25732), .dout(n25734));
  jor  g25566(.dina(n25734), .dinb(n25729), .dout(n25735));
  jxor g25567(.dina(n25735), .dinb(n93), .dout(n25736));
  jxor g25568(.dina(n25736), .dinb(n25728), .dout(n25737));
  jand g25569(.dina(n20358), .dinb(n71), .dout(n25738));
  jand g25570(.dina(n20204), .dinb(n796), .dout(n25739));
  jand g25571(.dina(n20205), .dinb(n731), .dout(n25740));
  jand g25572(.dina(n19922), .dinb(n1806), .dout(n25741));
  jor  g25573(.dina(n25741), .dinb(n25740), .dout(n25742));
  jor  g25574(.dina(n25742), .dinb(n25739), .dout(n25743));
  jor  g25575(.dina(n25743), .dinb(n25738), .dout(n25744));
  jxor g25576(.dina(n25744), .dinb(n77), .dout(n25745));
  jxor g25577(.dina(n25745), .dinb(n25737), .dout(n25746));
  jxor g25578(.dina(n25746), .dinb(n25687), .dout(n25747));
  jand g25579(.dina(n21367), .dinb(n806), .dout(n25748));
  jand g25580(.dina(n20947), .dinb(n1612), .dout(n25749));
  jand g25581(.dina(n21198), .dinb(n1620), .dout(n25750));
  jor  g25582(.dina(n25750), .dinb(n25749), .dout(n25751));
  jand g25583(.dina(n20344), .dinb(n1644), .dout(n25752));
  jor  g25584(.dina(n25752), .dinb(n25751), .dout(n25753));
  jor  g25585(.dina(n25753), .dinb(n25748), .dout(n25754));
  jxor g25586(.dina(n25754), .dinb(n65), .dout(n25755));
  jxor g25587(.dina(n25755), .dinb(n25747), .dout(n25756));
  jxor g25588(.dina(n25756), .dinb(n25683), .dout(n25757));
  jand g25589(.dina(n21976), .dinb(n1819), .dout(n25758));
  jand g25590(.dina(n21974), .dinb(n2243), .dout(n25759));
  jand g25591(.dina(n21340), .dinb(n2180), .dout(n25760));
  jand g25592(.dina(n21197), .dinb(n2185), .dout(n25761));
  jor  g25593(.dina(n25761), .dinb(n25760), .dout(n25762));
  jor  g25594(.dina(n25762), .dinb(n25759), .dout(n25763));
  jor  g25595(.dina(n25763), .dinb(n25758), .dout(n25764));
  jxor g25596(.dina(n25764), .dinb(n2196), .dout(n25765));
  jxor g25597(.dina(n25765), .dinb(n25757), .dout(n25766));
  jxor g25598(.dina(n25766), .dinb(n25679), .dout(n25767));
  jand g25599(.dina(n22267), .dinb(n2743), .dout(n25768));
  jand g25600(.dina(n22265), .dinb(n2752), .dout(n25769));
  jand g25601(.dina(n22163), .dinb(n2748), .dout(n25770));
  jand g25602(.dina(n22164), .dinb(n2757), .dout(n25771));
  jor  g25603(.dina(n25771), .dinb(n25770), .dout(n25772));
  jor  g25604(.dina(n25772), .dinb(n25769), .dout(n25773));
  jor  g25605(.dina(n25773), .dinb(n25768), .dout(n25774));
  jxor g25606(.dina(n25774), .dinb(n2441), .dout(n25775));
  jxor g25607(.dina(n25775), .dinb(n25767), .dout(n25776));
  jxor g25608(.dina(n25776), .dinb(n25675), .dout(n25777));
  jnot g25609(.din(n25619), .dout(n25778));
  jor  g25610(.dina(n25778), .dinb(n25524), .dout(n25779));
  jor  g25611(.dina(n25628), .dinb(n25620), .dout(n25780));
  jand g25612(.dina(n25780), .dinb(n25779), .dout(n25781));
  jor  g25613(.dina(n25272), .dinb(n3424), .dout(n25782));
  jor  g25614(.dina(n25276), .dinb(n3429), .dout(n25783));
  jor  g25615(.dina(n25274), .dinb(n3426), .dout(n25784));
  jand g25616(.dina(n25784), .dinb(n25783), .dout(n25785));
  jor  g25617(.dina(n25278), .dinb(n3211), .dout(n25786));
  jand g25618(.dina(n25786), .dinb(n25785), .dout(n25787));
  jand g25619(.dina(n25787), .dinb(n25782), .dout(n25788));
  jxor g25620(.dina(n25788), .dinb(\a[14] ), .dout(n25789));
  jxor g25621(.dina(n25789), .dinb(n25781), .dout(n25790));
  jxor g25622(.dina(n25790), .dinb(n25777), .dout(n25791));
  jor  g25623(.dina(n25286), .dinb(n4023), .dout(n25792));
  jor  g25624(.dina(n24266), .dinb(n4025), .dout(n25793));
  jor  g25625(.dina(n24265), .dinb(n4028), .dout(n25794));
  jor  g25626(.dina(n25290), .dinb(n3871), .dout(n25795));
  jand g25627(.dina(n25795), .dinb(n25794), .dout(n25796));
  jand g25628(.dina(n25796), .dinb(n25793), .dout(n25797));
  jand g25629(.dina(n25797), .dinb(n25792), .dout(n25798));
  jxor g25630(.dina(n25798), .dinb(\a[11] ), .dout(n25799));
  jxor g25631(.dina(n25799), .dinb(n25791), .dout(n25800));
  jxor g25632(.dina(n25800), .dinb(n25671), .dout(n25801));
  jnot g25633(.din(n25514), .dout(n25802));
  jand g25634(.dina(n25640), .dinb(n25802), .dout(n25803));
  jnot g25635(.din(n25803), .dout(n25804));
  jor  g25636(.dina(n25649), .dinb(n25641), .dout(n25805));
  jand g25637(.dina(n25805), .dinb(n25804), .dout(n25806));
  jor  g25638(.dina(n24736), .dinb(n4692), .dout(n25807));
  jor  g25639(.dina(n24738), .dinb(n4705), .dout(n25808));
  jor  g25640(.dina(n24518), .dinb(n4697), .dout(n25809));
  jor  g25641(.dina(n24304), .dinb(n4702), .dout(n25810));
  jand g25642(.dina(n25810), .dinb(n25809), .dout(n25811));
  jand g25643(.dina(n25811), .dinb(n25808), .dout(n25812));
  jand g25644(.dina(n25812), .dinb(n25807), .dout(n25813));
  jxor g25645(.dina(n25813), .dinb(\a[8] ), .dout(n25814));
  jxor g25646(.dina(n25814), .dinb(n25806), .dout(n25815));
  jxor g25647(.dina(n25815), .dinb(n25801), .dout(n25816));
  jxor g25648(.dina(n25816), .dinb(n25665), .dout(n25817));
  jxor g25649(.dina(n25817), .dinb(n25661), .dout(n25818));
  jxor g25650(.dina(n25818), .dinb(n25658), .dout(\result[10] ));
  jand g25651(.dina(n25818), .dinb(n25658), .dout(n25820));
  jand g25652(.dina(n25816), .dinb(n25665), .dout(n25821));
  jand g25653(.dina(n25817), .dinb(n25661), .dout(n25822));
  jor  g25654(.dina(n25822), .dinb(n25821), .dout(n25823));
  jor  g25655(.dina(n25814), .dinb(n25806), .dout(n25824));
  jnot g25656(.din(n25824), .dout(n25825));
  jand g25657(.dina(n25815), .dinb(n25801), .dout(n25826));
  jor  g25658(.dina(n25826), .dinb(n25825), .dout(n25827));
  jnot g25659(.din(n25791), .dout(n25828));
  jnot g25660(.din(n25799), .dout(n25829));
  jand g25661(.dina(n25829), .dinb(n25828), .dout(n25830));
  jand g25662(.dina(n25800), .dinb(n25671), .dout(n25831));
  jor  g25663(.dina(n25831), .dinb(n25830), .dout(n25832));
  jor  g25664(.dina(n25789), .dinb(n25781), .dout(n25833));
  jnot g25665(.din(n25790), .dout(n25834));
  jor  g25666(.dina(n25834), .dinb(n25777), .dout(n25835));
  jand g25667(.dina(n25835), .dinb(n25833), .dout(n25836));
  jor  g25668(.dina(n25775), .dinb(n25767), .dout(n25837));
  jnot g25669(.din(n25837), .dout(n25838));
  jnot g25670(.din(n25675), .dout(n25839));
  jand g25671(.dina(n25776), .dinb(n25839), .dout(n25840));
  jor  g25672(.dina(n25840), .dinb(n25838), .dout(n25841));
  jor  g25673(.dina(n25765), .dinb(n25757), .dout(n25842));
  jxor g25674(.dina(n25726), .dinb(n25694), .dout(n25843));
  jxor g25675(.dina(n25736), .dinb(n25843), .dout(n25844));
  jxor g25676(.dina(n25745), .dinb(n25844), .dout(n25845));
  jxor g25677(.dina(n25845), .dinb(n25687), .dout(n25846));
  jxor g25678(.dina(n25755), .dinb(n25846), .dout(n25847));
  jxor g25679(.dina(n25847), .dinb(n25683), .dout(n25848));
  jxor g25680(.dina(n25765), .dinb(n25848), .dout(n25849));
  jor  g25681(.dina(n25849), .dinb(n25679), .dout(n25850));
  jand g25682(.dina(n25850), .dinb(n25842), .dout(n25851));
  jor  g25683(.dina(n25755), .dinb(n25747), .dout(n25852));
  jor  g25684(.dina(n25847), .dinb(n25683), .dout(n25853));
  jand g25685(.dina(n25853), .dinb(n25852), .dout(n25854));
  jor  g25686(.dina(n25745), .dinb(n25737), .dout(n25855));
  jor  g25687(.dina(n25845), .dinb(n25687), .dout(n25856));
  jand g25688(.dina(n25856), .dinb(n25855), .dout(n25857));
  jor  g25689(.dina(n25727), .dinb(n25694), .dout(n25858));
  jor  g25690(.dina(n25736), .dinb(n25843), .dout(n25859));
  jand g25691(.dina(n25859), .dinb(n25858), .dout(n25860));
  jand g25692(.dina(n25724), .dinb(n25705), .dout(n25861));
  jand g25693(.dina(n25725), .dinb(n25701), .dout(n25862));
  jor  g25694(.dina(n25862), .dinb(n25861), .dout(n25863));
  jand g25695(.dina(n19399), .dinb(n5076), .dout(n25864));
  jand g25696(.dina(n19220), .dinb(n5084), .dout(n25865));
  jand g25697(.dina(n18914), .dinb(n5082), .dout(n25866));
  jand g25698(.dina(n18488), .dinb(n6050), .dout(n25867));
  jor  g25699(.dina(n25867), .dinb(n25866), .dout(n25868));
  jor  g25700(.dina(n25868), .dinb(n25865), .dout(n25869));
  jor  g25701(.dina(n25869), .dinb(n25864), .dout(n25870));
  jand g25702(.dina(n7113), .dinb(n521), .dout(n25871));
  jand g25703(.dina(n8822), .dinb(n2730), .dout(n25872));
  jand g25704(.dina(n25872), .dinb(n25871), .dout(n25873));
  jand g25705(.dina(n1037), .dinb(n1226), .dout(n25874));
  jand g25706(.dina(n3812), .dinb(n1495), .dout(n25875));
  jand g25707(.dina(n25875), .dinb(n25874), .dout(n25876));
  jand g25708(.dina(n25876), .dinb(n1489), .dout(n25877));
  jand g25709(.dina(n25877), .dinb(n25873), .dout(n25878));
  jand g25710(.dina(n4588), .dinb(n3747), .dout(n25879));
  jand g25711(.dina(n5478), .dinb(n2149), .dout(n25880));
  jand g25712(.dina(n25880), .dinb(n25879), .dout(n25881));
  jand g25713(.dina(n25881), .dinb(n25878), .dout(n25882));
  jand g25714(.dina(n1709), .dinb(n481), .dout(n25883));
  jand g25715(.dina(n647), .dinb(n829), .dout(n25884));
  jand g25716(.dina(n25884), .dinb(n1260), .dout(n25885));
  jand g25717(.dina(n25885), .dinb(n25883), .dout(n25886));
  jand g25718(.dina(n886), .dinb(n1213), .dout(n25887));
  jand g25719(.dina(n25887), .dinb(n15651), .dout(n25888));
  jand g25720(.dina(n25888), .dinb(n12439), .dout(n25889));
  jand g25721(.dina(n25889), .dinb(n25886), .dout(n25890));
  jand g25722(.dina(n25890), .dinb(n3784), .dout(n25891));
  jand g25723(.dina(n25891), .dinb(n25882), .dout(n25892));
  jand g25724(.dina(n4674), .dinb(n1868), .dout(n25893));
  jand g25725(.dina(n3329), .dinb(n1877), .dout(n25894));
  jand g25726(.dina(n25894), .dinb(n3161), .dout(n25895));
  jand g25727(.dina(n25895), .dinb(n6033), .dout(n25896));
  jand g25728(.dina(n25896), .dinb(n25893), .dout(n25897));
  jand g25729(.dina(n25897), .dinb(n5228), .dout(n25898));
  jand g25730(.dina(n25898), .dinb(n25892), .dout(n25899));
  jnot g25731(.din(n25899), .dout(n25900));
  jor  g25732(.dina(n25720), .dinb(n25202), .dout(n25901));
  jand g25733(.dina(n25723), .dinb(n25721), .dout(n25902));
  jnot g25734(.din(n25902), .dout(n25903));
  jand g25735(.dina(n25903), .dinb(n25901), .dout(n25904));
  jxor g25736(.dina(n25904), .dinb(n25900), .dout(n25905));
  jxor g25737(.dina(n25905), .dinb(n25870), .dout(n25906));
  jxor g25738(.dina(n25906), .dinb(n25863), .dout(n25907));
  jand g25739(.dina(n19924), .dinb(n2936), .dout(n25908));
  jand g25740(.dina(n19373), .dinb(n2940), .dout(n25909));
  jand g25741(.dina(n19922), .dinb(n2943), .dout(n25910));
  jor  g25742(.dina(n25910), .dinb(n25909), .dout(n25911));
  jand g25743(.dina(n19219), .dinb(n3684), .dout(n25912));
  jor  g25744(.dina(n25912), .dinb(n25911), .dout(n25913));
  jor  g25745(.dina(n25913), .dinb(n25908), .dout(n25914));
  jxor g25746(.dina(n25914), .dinb(n93), .dout(n25915));
  jnot g25747(.din(n25915), .dout(n25916));
  jxor g25748(.dina(n25916), .dinb(n25907), .dout(n25917));
  jxor g25749(.dina(n25917), .dinb(n25860), .dout(n25918));
  jand g25750(.dina(n20346), .dinb(n71), .dout(n25919));
  jand g25751(.dina(n20344), .dinb(n796), .dout(n25920));
  jand g25752(.dina(n20204), .dinb(n731), .dout(n25921));
  jand g25753(.dina(n20205), .dinb(n1806), .dout(n25922));
  jor  g25754(.dina(n25922), .dinb(n25921), .dout(n25923));
  jor  g25755(.dina(n25923), .dinb(n25920), .dout(n25924));
  jor  g25756(.dina(n25924), .dinb(n25919), .dout(n25925));
  jxor g25757(.dina(n25925), .dinb(n77), .dout(n25926));
  jxor g25758(.dina(n25926), .dinb(n25918), .dout(n25927));
  jxor g25759(.dina(n25927), .dinb(n25857), .dout(n25928));
  jand g25760(.dina(n21355), .dinb(n806), .dout(n25929));
  jand g25761(.dina(n21198), .dinb(n1612), .dout(n25930));
  jand g25762(.dina(n21197), .dinb(n1620), .dout(n25931));
  jor  g25763(.dina(n25931), .dinb(n25930), .dout(n25932));
  jand g25764(.dina(n20947), .dinb(n1644), .dout(n25933));
  jor  g25765(.dina(n25933), .dinb(n25932), .dout(n25934));
  jor  g25766(.dina(n25934), .dinb(n25929), .dout(n25935));
  jxor g25767(.dina(n25935), .dinb(n65), .dout(n25936));
  jxor g25768(.dina(n25936), .dinb(n25928), .dout(n25937));
  jxor g25769(.dina(n25937), .dinb(n25854), .dout(n25938));
  jand g25770(.dina(n22291), .dinb(n1819), .dout(n25939));
  jand g25771(.dina(n21974), .dinb(n2180), .dout(n25940));
  jand g25772(.dina(n22164), .dinb(n2243), .dout(n25941));
  jor  g25773(.dina(n25941), .dinb(n25940), .dout(n25942));
  jand g25774(.dina(n21340), .dinb(n2185), .dout(n25943));
  jor  g25775(.dina(n25943), .dinb(n25942), .dout(n25944));
  jor  g25776(.dina(n25944), .dinb(n25939), .dout(n25945));
  jxor g25777(.dina(n25945), .dinb(n2196), .dout(n25946));
  jxor g25778(.dina(n25946), .dinb(n25938), .dout(n25947));
  jxor g25779(.dina(n25947), .dinb(n25851), .dout(n25948));
  jand g25780(.dina(n22939), .dinb(n2743), .dout(n25949));
  jand g25781(.dina(n22937), .dinb(n2752), .dout(n25950));
  jand g25782(.dina(n22265), .dinb(n2748), .dout(n25951));
  jand g25783(.dina(n22163), .dinb(n2757), .dout(n25952));
  jor  g25784(.dina(n25952), .dinb(n25951), .dout(n25953));
  jor  g25785(.dina(n25953), .dinb(n25950), .dout(n25954));
  jor  g25786(.dina(n25954), .dinb(n25949), .dout(n25955));
  jxor g25787(.dina(n25955), .dinb(n2441), .dout(n25956));
  jxor g25788(.dina(n25956), .dinb(n25948), .dout(n25957));
  jxor g25789(.dina(n25957), .dinb(n25841), .dout(n25958));
  jand g25790(.dina(n23146), .dinb(n3423), .dout(n25959));
  jand g25791(.dina(n23079), .dinb(n3428), .dout(n25960));
  jand g25792(.dina(n23144), .dinb(n3569), .dout(n25961));
  jor  g25793(.dina(n25961), .dinb(n25960), .dout(n25962));
  jand g25794(.dina(n23080), .dinb(n3210), .dout(n25963));
  jor  g25795(.dina(n25963), .dinb(n25962), .dout(n25964));
  jor  g25796(.dina(n25964), .dinb(n25959), .dout(n25965));
  jxor g25797(.dina(n25965), .dinb(n3473), .dout(n25966));
  jxor g25798(.dina(n25966), .dinb(n25958), .dout(n25967));
  jxor g25799(.dina(n25967), .dinb(n25836), .dout(n25968));
  jor  g25800(.dina(n24302), .dinb(n4023), .dout(n25969));
  jor  g25801(.dina(n24266), .dinb(n4028), .dout(n25970));
  jor  g25802(.dina(n24304), .dinb(n4025), .dout(n25971));
  jand g25803(.dina(n25971), .dinb(n25970), .dout(n25972));
  jor  g25804(.dina(n24265), .dinb(n3871), .dout(n25973));
  jand g25805(.dina(n25973), .dinb(n25972), .dout(n25974));
  jand g25806(.dina(n25974), .dinb(n25969), .dout(n25975));
  jxor g25807(.dina(n25975), .dinb(\a[11] ), .dout(n25976));
  jnot g25808(.din(n25976), .dout(n25977));
  jxor g25809(.dina(n25977), .dinb(n25968), .dout(n25978));
  jxor g25810(.dina(n25978), .dinb(n25832), .dout(n25979));
  jor  g25811(.dina(n24932), .dinb(n4692), .dout(n25980));
  jor  g25812(.dina(n24738), .dinb(n4697), .dout(n25981));
  jor  g25813(.dina(n24930), .dinb(n4705), .dout(n25982));
  jand g25814(.dina(n25982), .dinb(n25981), .dout(n25983));
  jor  g25815(.dina(n24518), .dinb(n4702), .dout(n25984));
  jand g25816(.dina(n25984), .dinb(n25983), .dout(n25985));
  jand g25817(.dina(n25985), .dinb(n25980), .dout(n25986));
  jxor g25818(.dina(n25986), .dinb(\a[8] ), .dout(n25987));
  jnot g25819(.din(n25987), .dout(n25988));
  jxor g25820(.dina(n25988), .dinb(n25979), .dout(n25989));
  jxor g25821(.dina(n25989), .dinb(n25827), .dout(n25990));
  jxor g25822(.dina(n25990), .dinb(n25823), .dout(n25991));
  jxor g25823(.dina(n25991), .dinb(n25820), .dout(\result[11] ));
  jand g25824(.dina(n25991), .dinb(n25820), .dout(n25993));
  jand g25825(.dina(n25978), .dinb(n25832), .dout(n25994));
  jand g25826(.dina(n25988), .dinb(n25979), .dout(n25995));
  jor  g25827(.dina(n25995), .dinb(n25994), .dout(n25996));
  jor  g25828(.dina(n25967), .dinb(n25836), .dout(n25997));
  jnot g25829(.din(n25997), .dout(n25998));
  jand g25830(.dina(n25977), .dinb(n25968), .dout(n25999));
  jor  g25831(.dina(n25999), .dinb(n25998), .dout(n26000));
  jor  g25832(.dina(n25116), .dinb(n4692), .dout(n26001));
  jor  g25833(.dina(n24930), .dinb(n18774), .dout(n26002));
  jor  g25834(.dina(n24738), .dinb(n4702), .dout(n26003));
  jand g25835(.dina(n26003), .dinb(n26002), .dout(n26004));
  jand g25836(.dina(n26004), .dinb(n26001), .dout(n26005));
  jxor g25837(.dina(n26005), .dinb(\a[8] ), .dout(n26006));
  jnot g25838(.din(n26006), .dout(n26007));
  jxor g25839(.dina(n26007), .dinb(n26000), .dout(n26008));
  jand g25840(.dina(n25957), .dinb(n25841), .dout(n26009));
  jnot g25841(.din(n26009), .dout(n26010));
  jnot g25842(.din(n25958), .dout(n26011));
  jor  g25843(.dina(n25966), .dinb(n26011), .dout(n26012));
  jand g25844(.dina(n26012), .dinb(n26010), .dout(n26013));
  jnot g25845(.din(n25947), .dout(n26014));
  jor  g25846(.dina(n26014), .dinb(n25851), .dout(n26015));
  jor  g25847(.dina(n25956), .dinb(n25948), .dout(n26016));
  jand g25848(.dina(n26016), .dinb(n26015), .dout(n26017));
  jnot g25849(.din(n26017), .dout(n26018));
  jnot g25850(.din(n25937), .dout(n26019));
  jor  g25851(.dina(n26019), .dinb(n25854), .dout(n26020));
  jor  g25852(.dina(n25946), .dinb(n25938), .dout(n26021));
  jand g25853(.dina(n26021), .dinb(n26020), .dout(n26022));
  jnot g25854(.din(n25927), .dout(n26023));
  jor  g25855(.dina(n26023), .dinb(n25857), .dout(n26024));
  jor  g25856(.dina(n25936), .dinb(n25928), .dout(n26025));
  jand g25857(.dina(n26025), .dinb(n26024), .dout(n26026));
  jnot g25858(.din(n25917), .dout(n26027));
  jor  g25859(.dina(n26027), .dinb(n25860), .dout(n26028));
  jor  g25860(.dina(n25926), .dinb(n25918), .dout(n26029));
  jand g25861(.dina(n26029), .dinb(n26028), .dout(n26030));
  jand g25862(.dina(n25906), .dinb(n25863), .dout(n26031));
  jand g25863(.dina(n25916), .dinb(n25907), .dout(n26032));
  jor  g25864(.dina(n26032), .dinb(n26031), .dout(n26033));
  jand g25865(.dina(n19387), .dinb(n5076), .dout(n26034));
  jand g25866(.dina(n19219), .dinb(n5084), .dout(n26035));
  jand g25867(.dina(n19220), .dinb(n5082), .dout(n26036));
  jand g25868(.dina(n18914), .dinb(n6050), .dout(n26037));
  jor  g25869(.dina(n26037), .dinb(n26036), .dout(n26038));
  jor  g25870(.dina(n26038), .dinb(n26035), .dout(n26039));
  jor  g25871(.dina(n26039), .dinb(n26034), .dout(n26040));
  jor  g25872(.dina(n25904), .dinb(n25900), .dout(n26041));
  jand g25873(.dina(n25905), .dinb(n25870), .dout(n26042));
  jnot g25874(.din(n26042), .dout(n26043));
  jand g25875(.dina(n26043), .dinb(n26041), .dout(n26044));
  jnot g25876(.din(n26044), .dout(n26045));
  jand g25877(.dina(n19961), .dinb(n13294), .dout(n26046));
  jand g25878(.dina(n14220), .dinb(n4569), .dout(n26047));
  jand g25879(.dina(n26047), .dinb(n3133), .dout(n26048));
  jand g25880(.dina(n11224), .dinb(n1437), .dout(n26049));
  jand g25881(.dina(n26049), .dinb(n1493), .dout(n26050));
  jand g25882(.dina(n26050), .dinb(n26048), .dout(n26051));
  jand g25883(.dina(n1561), .dinb(n1271), .dout(n26052));
  jand g25884(.dina(n1207), .dinb(n108), .dout(n26053));
  jand g25885(.dina(n26053), .dinb(n1763), .dout(n26054));
  jand g25886(.dina(n26054), .dinb(n26052), .dout(n26055));
  jand g25887(.dina(n26055), .dinb(n4448), .dout(n26056));
  jand g25888(.dina(n26056), .dinb(n26051), .dout(n26057));
  jand g25889(.dina(n26057), .dinb(n8126), .dout(n26058));
  jand g25890(.dina(n26058), .dinb(n553), .dout(n26059));
  jand g25891(.dina(n21120), .dinb(n818), .dout(n26060));
  jand g25892(.dina(n26060), .dinb(n13540), .dout(n26061));
  jand g25893(.dina(n1053), .dinb(n430), .dout(n26062));
  jand g25894(.dina(n26062), .dinb(n920), .dout(n26063));
  jand g25895(.dina(n26063), .dinb(n954), .dout(n26064));
  jand g25896(.dina(n588), .dinb(n1575), .dout(n26065));
  jand g25897(.dina(n1005), .dinb(n1315), .dout(n26066));
  jand g25898(.dina(n886), .dinb(n1310), .dout(n26067));
  jand g25899(.dina(n26067), .dinb(n26066), .dout(n26068));
  jand g25900(.dina(n2148), .dinb(n619), .dout(n26069));
  jand g25901(.dina(n26069), .dinb(n470), .dout(n26070));
  jand g25902(.dina(n26070), .dinb(n26068), .dout(n26071));
  jand g25903(.dina(n26071), .dinb(n26065), .dout(n26072));
  jand g25904(.dina(n26072), .dinb(n532), .dout(n26073));
  jand g25905(.dina(n26073), .dinb(n26064), .dout(n26074));
  jand g25906(.dina(n26074), .dinb(n26061), .dout(n26075));
  jand g25907(.dina(n26075), .dinb(n948), .dout(n26076));
  jand g25908(.dina(n26076), .dinb(n26059), .dout(n26077));
  jand g25909(.dina(n26077), .dinb(n26046), .dout(n26078));
  jxor g25910(.dina(n26078), .dinb(n25900), .dout(n26079));
  jxor g25911(.dina(n26079), .dinb(n26045), .dout(n26080));
  jxor g25912(.dina(n26080), .dinb(n26040), .dout(n26081));
  jxor g25913(.dina(n26081), .dinb(n26033), .dout(n26082));
  jand g25914(.dina(n20371), .dinb(n2936), .dout(n26083));
  jand g25915(.dina(n19922), .dinb(n2940), .dout(n26084));
  jand g25916(.dina(n20205), .dinb(n2943), .dout(n26085));
  jor  g25917(.dina(n26085), .dinb(n26084), .dout(n26086));
  jand g25918(.dina(n19373), .dinb(n3684), .dout(n26087));
  jor  g25919(.dina(n26087), .dinb(n26086), .dout(n26088));
  jor  g25920(.dina(n26088), .dinb(n26083), .dout(n26089));
  jxor g25921(.dina(n26089), .dinb(n93), .dout(n26090));
  jxor g25922(.dina(n26090), .dinb(n26082), .dout(n26091));
  jand g25923(.dina(n20949), .dinb(n71), .dout(n26092));
  jand g25924(.dina(n20947), .dinb(n796), .dout(n26093));
  jand g25925(.dina(n20344), .dinb(n731), .dout(n26094));
  jand g25926(.dina(n20204), .dinb(n1806), .dout(n26095));
  jor  g25927(.dina(n26095), .dinb(n26094), .dout(n26096));
  jor  g25928(.dina(n26096), .dinb(n26093), .dout(n26097));
  jor  g25929(.dina(n26097), .dinb(n26092), .dout(n26098));
  jxor g25930(.dina(n26098), .dinb(n77), .dout(n26099));
  jxor g25931(.dina(n26099), .dinb(n26091), .dout(n26100));
  jxor g25932(.dina(n26100), .dinb(n26030), .dout(n26101));
  jand g25933(.dina(n21342), .dinb(n806), .dout(n26102));
  jand g25934(.dina(n21197), .dinb(n1612), .dout(n26103));
  jand g25935(.dina(n21340), .dinb(n1620), .dout(n26104));
  jor  g25936(.dina(n26104), .dinb(n26103), .dout(n26105));
  jand g25937(.dina(n21198), .dinb(n1644), .dout(n26106));
  jor  g25938(.dina(n26106), .dinb(n26105), .dout(n26107));
  jor  g25939(.dina(n26107), .dinb(n26102), .dout(n26108));
  jxor g25940(.dina(n26108), .dinb(n65), .dout(n26109));
  jxor g25941(.dina(n26109), .dinb(n26101), .dout(n26110));
  jxor g25942(.dina(n26110), .dinb(n26026), .dout(n26111));
  jand g25943(.dina(n22279), .dinb(n1819), .dout(n26112));
  jand g25944(.dina(n22163), .dinb(n2243), .dout(n26113));
  jand g25945(.dina(n22164), .dinb(n2180), .dout(n26114));
  jand g25946(.dina(n21974), .dinb(n2185), .dout(n26115));
  jor  g25947(.dina(n26115), .dinb(n26114), .dout(n26116));
  jor  g25948(.dina(n26116), .dinb(n26113), .dout(n26117));
  jor  g25949(.dina(n26117), .dinb(n26112), .dout(n26118));
  jxor g25950(.dina(n26118), .dinb(n2196), .dout(n26119));
  jxor g25951(.dina(n26119), .dinb(n26111), .dout(n26120));
  jxor g25952(.dina(n26120), .dinb(n26022), .dout(n26121));
  jand g25953(.dina(n23172), .dinb(n2743), .dout(n26122));
  jand g25954(.dina(n23080), .dinb(n2752), .dout(n26123));
  jand g25955(.dina(n22937), .dinb(n2748), .dout(n26124));
  jand g25956(.dina(n22265), .dinb(n2757), .dout(n26125));
  jor  g25957(.dina(n26125), .dinb(n26124), .dout(n26126));
  jor  g25958(.dina(n26126), .dinb(n26123), .dout(n26127));
  jor  g25959(.dina(n26127), .dinb(n26122), .dout(n26128));
  jxor g25960(.dina(n26128), .dinb(n2441), .dout(n26129));
  jxor g25961(.dina(n26129), .dinb(n26121), .dout(n26130));
  jxor g25962(.dina(n26130), .dinb(n26018), .dout(n26131));
  jnot g25963(.din(n26131), .dout(n26132));
  jand g25964(.dina(n23847), .dinb(n3423), .dout(n26133));
  jand g25965(.dina(n23845), .dinb(n3569), .dout(n26134));
  jand g25966(.dina(n23144), .dinb(n3428), .dout(n26135));
  jand g25967(.dina(n23079), .dinb(n3210), .dout(n26136));
  jor  g25968(.dina(n26136), .dinb(n26135), .dout(n26137));
  jor  g25969(.dina(n26137), .dinb(n26134), .dout(n26138));
  jor  g25970(.dina(n26138), .dinb(n26133), .dout(n26139));
  jxor g25971(.dina(n26139), .dinb(n3473), .dout(n26140));
  jxor g25972(.dina(n26140), .dinb(n26132), .dout(n26141));
  jxor g25973(.dina(n26141), .dinb(n26013), .dout(n26142));
  jor  g25974(.dina(n24516), .dinb(n4023), .dout(n26143));
  jor  g25975(.dina(n24304), .dinb(n4028), .dout(n26144));
  jor  g25976(.dina(n24518), .dinb(n4025), .dout(n26145));
  jand g25977(.dina(n26145), .dinb(n26144), .dout(n26146));
  jor  g25978(.dina(n24266), .dinb(n3871), .dout(n26147));
  jand g25979(.dina(n26147), .dinb(n26146), .dout(n26148));
  jand g25980(.dina(n26148), .dinb(n26143), .dout(n26149));
  jxor g25981(.dina(n26149), .dinb(\a[11] ), .dout(n26150));
  jxor g25982(.dina(n26150), .dinb(n26142), .dout(n26151));
  jxor g25983(.dina(n26151), .dinb(n26008), .dout(n26152));
  jxor g25984(.dina(n26152), .dinb(n25996), .dout(n26153));
  jand g25985(.dina(n25989), .dinb(n25827), .dout(n26154));
  jand g25986(.dina(n25990), .dinb(n25823), .dout(n26155));
  jor  g25987(.dina(n26155), .dinb(n26154), .dout(n26156));
  jxor g25988(.dina(n26156), .dinb(n26153), .dout(n26157));
  jxor g25989(.dina(n26157), .dinb(n25993), .dout(\result[12] ));
  jand g25990(.dina(n26157), .dinb(n25993), .dout(n26159));
  jand g25991(.dina(n26152), .dinb(n25996), .dout(n26160));
  jand g25992(.dina(n26156), .dinb(n26153), .dout(n26161));
  jor  g25993(.dina(n26161), .dinb(n26160), .dout(n26162));
  jand g25994(.dina(n26007), .dinb(n26000), .dout(n26163));
  jand g25995(.dina(n26151), .dinb(n26008), .dout(n26164));
  jor  g25996(.dina(n26164), .dinb(n26163), .dout(n26165));
  jand g25997(.dina(n26130), .dinb(n26018), .dout(n26166));
  jnot g25998(.din(n26166), .dout(n26167));
  jor  g25999(.dina(n26140), .dinb(n26132), .dout(n26168));
  jand g26000(.dina(n26168), .dinb(n26167), .dout(n26169));
  jnot g26001(.din(n26026), .dout(n26170));
  jand g26002(.dina(n26110), .dinb(n26170), .dout(n26171));
  jnot g26003(.din(n26171), .dout(n26172));
  jor  g26004(.dina(n26119), .dinb(n26111), .dout(n26173));
  jand g26005(.dina(n26173), .dinb(n26172), .dout(n26174));
  jnot g26006(.din(n26030), .dout(n26175));
  jand g26007(.dina(n26100), .dinb(n26175), .dout(n26176));
  jnot g26008(.din(n26176), .dout(n26177));
  jor  g26009(.dina(n26109), .dinb(n26101), .dout(n26178));
  jand g26010(.dina(n26178), .dinb(n26177), .dout(n26179));
  jnot g26011(.din(n26082), .dout(n26180));
  jor  g26012(.dina(n26090), .dinb(n26180), .dout(n26181));
  jor  g26013(.dina(n26099), .dinb(n26091), .dout(n26182));
  jand g26014(.dina(n26182), .dinb(n26181), .dout(n26183));
  jand g26015(.dina(n26080), .dinb(n26040), .dout(n26184));
  jand g26016(.dina(n26081), .dinb(n26033), .dout(n26185));
  jor  g26017(.dina(n26185), .dinb(n26184), .dout(n26186));
  jor  g26018(.dina(n26078), .dinb(n25900), .dout(n26187));
  jand g26019(.dina(n26079), .dinb(n26045), .dout(n26188));
  jnot g26020(.din(n26188), .dout(n26189));
  jand g26021(.dina(n26189), .dinb(n26187), .dout(n26190));
  jand g26022(.dina(n1541), .dinb(n1427), .dout(n26191));
  jand g26023(.dina(n504), .dinb(n178), .dout(n26192));
  jand g26024(.dina(n26192), .dinb(n3276), .dout(n26193));
  jand g26025(.dina(n26193), .dinb(n26191), .dout(n26194));
  jand g26026(.dina(n5494), .dinb(n3769), .dout(n26195));
  jand g26027(.dina(n2567), .dinb(n1438), .dout(n26196));
  jand g26028(.dina(n26196), .dinb(n26195), .dout(n26197));
  jand g26029(.dina(n3405), .dinb(n1578), .dout(n26198));
  jand g26030(.dina(n26198), .dinb(n20842), .dout(n26199));
  jand g26031(.dina(n26199), .dinb(n26197), .dout(n26200));
  jand g26032(.dina(n26200), .dinb(n26194), .dout(n26201));
  jand g26033(.dina(n26201), .dinb(n2625), .dout(n26202));
  jand g26034(.dina(n5326), .dinb(n724), .dout(n26203));
  jand g26035(.dina(n26203), .dinb(n26202), .dout(n26204));
  jxor g26036(.dina(n26204), .dinb(n25899), .dout(n26205));
  jand g26037(.dina(n25199), .dinb(n18992), .dout(n26206));
  jxor g26038(.dina(n26206), .dinb(n4713), .dout(n26207));
  jxor g26039(.dina(n26207), .dinb(n26205), .dout(n26208));
  jxor g26040(.dina(n26208), .dinb(n26190), .dout(n26209));
  jand g26041(.dina(n19375), .dinb(n5076), .dout(n26210));
  jand g26042(.dina(n19373), .dinb(n5084), .dout(n26211));
  jand g26043(.dina(n19219), .dinb(n5082), .dout(n26212));
  jand g26044(.dina(n19220), .dinb(n6050), .dout(n26213));
  jor  g26045(.dina(n26213), .dinb(n26212), .dout(n26214));
  jor  g26046(.dina(n26214), .dinb(n26211), .dout(n26215));
  jor  g26047(.dina(n26215), .dinb(n26210), .dout(n26216));
  jnot g26048(.din(n26216), .dout(n26217));
  jxor g26049(.dina(n26217), .dinb(n26209), .dout(n26218));
  jand g26050(.dina(n20358), .dinb(n2936), .dout(n26219));
  jand g26051(.dina(n20204), .dinb(n2943), .dout(n26220));
  jand g26052(.dina(n20205), .dinb(n2940), .dout(n26221));
  jand g26053(.dina(n19922), .dinb(n3684), .dout(n26222));
  jor  g26054(.dina(n26222), .dinb(n26221), .dout(n26223));
  jor  g26055(.dina(n26223), .dinb(n26220), .dout(n26224));
  jor  g26056(.dina(n26224), .dinb(n26219), .dout(n26225));
  jxor g26057(.dina(n26225), .dinb(n93), .dout(n26226));
  jxor g26058(.dina(n26226), .dinb(n26218), .dout(n26227));
  jxor g26059(.dina(n26227), .dinb(n26186), .dout(n26228));
  jand g26060(.dina(n21367), .dinb(n71), .dout(n26229));
  jand g26061(.dina(n21198), .dinb(n796), .dout(n26230));
  jand g26062(.dina(n20947), .dinb(n731), .dout(n26231));
  jand g26063(.dina(n20344), .dinb(n1806), .dout(n26232));
  jor  g26064(.dina(n26232), .dinb(n26231), .dout(n26233));
  jor  g26065(.dina(n26233), .dinb(n26230), .dout(n26234));
  jor  g26066(.dina(n26234), .dinb(n26229), .dout(n26235));
  jxor g26067(.dina(n26235), .dinb(n77), .dout(n26236));
  jxor g26068(.dina(n26236), .dinb(n26228), .dout(n26237));
  jxor g26069(.dina(n26237), .dinb(n26183), .dout(n26238));
  jand g26070(.dina(n21976), .dinb(n806), .dout(n26239));
  jand g26071(.dina(n21340), .dinb(n1612), .dout(n26240));
  jand g26072(.dina(n21974), .dinb(n1620), .dout(n26241));
  jor  g26073(.dina(n26241), .dinb(n26240), .dout(n26242));
  jand g26074(.dina(n21197), .dinb(n1644), .dout(n26243));
  jor  g26075(.dina(n26243), .dinb(n26242), .dout(n26244));
  jor  g26076(.dina(n26244), .dinb(n26239), .dout(n26245));
  jxor g26077(.dina(n26245), .dinb(n65), .dout(n26246));
  jxor g26078(.dina(n26246), .dinb(n26238), .dout(n26247));
  jnot g26079(.din(n26247), .dout(n26248));
  jxor g26080(.dina(n26248), .dinb(n26179), .dout(n26249));
  jand g26081(.dina(n22267), .dinb(n1819), .dout(n26250));
  jand g26082(.dina(n22163), .dinb(n2180), .dout(n26251));
  jand g26083(.dina(n22265), .dinb(n2243), .dout(n26252));
  jor  g26084(.dina(n26252), .dinb(n26251), .dout(n26253));
  jand g26085(.dina(n22164), .dinb(n2185), .dout(n26254));
  jor  g26086(.dina(n26254), .dinb(n26253), .dout(n26255));
  jor  g26087(.dina(n26255), .dinb(n26250), .dout(n26256));
  jxor g26088(.dina(n26256), .dinb(n2196), .dout(n26257));
  jxor g26089(.dina(n26257), .dinb(n26249), .dout(n26258));
  jxor g26090(.dina(n26258), .dinb(n26174), .dout(n26259));
  jnot g26091(.din(n26022), .dout(n26260));
  jand g26092(.dina(n26120), .dinb(n26260), .dout(n26261));
  jnot g26093(.din(n26261), .dout(n26262));
  jor  g26094(.dina(n26129), .dinb(n26121), .dout(n26263));
  jand g26095(.dina(n26263), .dinb(n26262), .dout(n26264));
  jor  g26096(.dina(n25272), .dinb(n2744), .dout(n26265));
  jor  g26097(.dina(n25274), .dinb(n2753), .dout(n26266));
  jor  g26098(.dina(n25276), .dinb(n2749), .dout(n26267));
  jor  g26099(.dina(n25278), .dinb(n2758), .dout(n26268));
  jand g26100(.dina(n26268), .dinb(n26267), .dout(n26269));
  jand g26101(.dina(n26269), .dinb(n26266), .dout(n26270));
  jand g26102(.dina(n26270), .dinb(n26265), .dout(n26271));
  jxor g26103(.dina(n26271), .dinb(\a[17] ), .dout(n26272));
  jxor g26104(.dina(n26272), .dinb(n26264), .dout(n26273));
  jxor g26105(.dina(n26273), .dinb(n26259), .dout(n26274));
  jand g26106(.dina(n24077), .dinb(n3423), .dout(n26275));
  jand g26107(.dina(n23845), .dinb(n3428), .dout(n26276));
  jand g26108(.dina(n24075), .dinb(n3569), .dout(n26277));
  jor  g26109(.dina(n26277), .dinb(n26276), .dout(n26278));
  jand g26110(.dina(n23144), .dinb(n3210), .dout(n26279));
  jor  g26111(.dina(n26279), .dinb(n26278), .dout(n26280));
  jor  g26112(.dina(n26280), .dinb(n26275), .dout(n26281));
  jxor g26113(.dina(n26281), .dinb(n3473), .dout(n26282));
  jxor g26114(.dina(n26282), .dinb(n26274), .dout(n26283));
  jxor g26115(.dina(n26283), .dinb(n26169), .dout(n26284));
  jnot g26116(.din(n26141), .dout(n26285));
  jor  g26117(.dina(n26285), .dinb(n26013), .dout(n26286));
  jor  g26118(.dina(n26150), .dinb(n26142), .dout(n26287));
  jand g26119(.dina(n26287), .dinb(n26286), .dout(n26288));
  jor  g26120(.dina(n24736), .dinb(n4023), .dout(n26289));
  jor  g26121(.dina(n24738), .dinb(n4025), .dout(n26290));
  jor  g26122(.dina(n24518), .dinb(n4028), .dout(n26291));
  jor  g26123(.dina(n24304), .dinb(n3871), .dout(n26292));
  jand g26124(.dina(n26292), .dinb(n26291), .dout(n26293));
  jand g26125(.dina(n26293), .dinb(n26290), .dout(n26294));
  jand g26126(.dina(n26294), .dinb(n26289), .dout(n26295));
  jxor g26127(.dina(n26295), .dinb(\a[11] ), .dout(n26296));
  jxor g26128(.dina(n26296), .dinb(n26288), .dout(n26297));
  jxor g26129(.dina(n26297), .dinb(n26284), .dout(n26298));
  jxor g26130(.dina(n26298), .dinb(n26165), .dout(n26299));
  jxor g26131(.dina(n26299), .dinb(n26162), .dout(n26300));
  jxor g26132(.dina(n26300), .dinb(n26159), .dout(\result[13] ));
  jand g26133(.dina(n26300), .dinb(n26159), .dout(n26302));
  jand g26134(.dina(n26298), .dinb(n26165), .dout(n26303));
  jand g26135(.dina(n26299), .dinb(n26162), .dout(n26304));
  jor  g26136(.dina(n26304), .dinb(n26303), .dout(n26305));
  jor  g26137(.dina(n26296), .dinb(n26288), .dout(n26306));
  jnot g26138(.din(n26306), .dout(n26307));
  jand g26139(.dina(n26297), .dinb(n26284), .dout(n26308));
  jor  g26140(.dina(n26308), .dinb(n26307), .dout(n26309));
  jnot g26141(.din(n26274), .dout(n26310));
  jor  g26142(.dina(n26282), .dinb(n26310), .dout(n26311));
  jor  g26143(.dina(n26283), .dinb(n26169), .dout(n26312));
  jand g26144(.dina(n26312), .dinb(n26311), .dout(n26313));
  jor  g26145(.dina(n26272), .dinb(n26264), .dout(n26314));
  jnot g26146(.din(n26259), .dout(n26315));
  jnot g26147(.din(n26273), .dout(n26316));
  jor  g26148(.dina(n26316), .dinb(n26315), .dout(n26317));
  jand g26149(.dina(n26317), .dinb(n26314), .dout(n26318));
  jnot g26150(.din(n26249), .dout(n26319));
  jor  g26151(.dina(n26257), .dinb(n26319), .dout(n26320));
  jor  g26152(.dina(n26258), .dinb(n26174), .dout(n26321));
  jand g26153(.dina(n26321), .dinb(n26320), .dout(n26322));
  jor  g26154(.dina(n26246), .dinb(n26238), .dout(n26323));
  jor  g26155(.dina(n26248), .dinb(n26179), .dout(n26324));
  jand g26156(.dina(n26324), .dinb(n26323), .dout(n26325));
  jor  g26157(.dina(n26236), .dinb(n26228), .dout(n26326));
  jnot g26158(.din(n26237), .dout(n26327));
  jor  g26159(.dina(n26327), .dinb(n26183), .dout(n26328));
  jand g26160(.dina(n26328), .dinb(n26326), .dout(n26329));
  jnot g26161(.din(n26218), .dout(n26330));
  jor  g26162(.dina(n26226), .dinb(n26330), .dout(n26331));
  jnot g26163(.din(n26186), .dout(n26332));
  jor  g26164(.dina(n26227), .dinb(n26332), .dout(n26333));
  jand g26165(.dina(n26333), .dinb(n26331), .dout(n26334));
  jnot g26166(.din(n26190), .dout(n26335));
  jand g26167(.dina(n26208), .dinb(n26335), .dout(n26336));
  jnot g26168(.din(n26336), .dout(n26337));
  jor  g26169(.dina(n26217), .dinb(n26209), .dout(n26338));
  jand g26170(.dina(n26338), .dinb(n26337), .dout(n26339));
  jand g26171(.dina(n19924), .dinb(n5076), .dout(n26340));
  jand g26172(.dina(n19922), .dinb(n5084), .dout(n26341));
  jand g26173(.dina(n19373), .dinb(n5082), .dout(n26342));
  jand g26174(.dina(n19219), .dinb(n6050), .dout(n26343));
  jor  g26175(.dina(n26343), .dinb(n26342), .dout(n26344));
  jor  g26176(.dina(n26344), .dinb(n26341), .dout(n26345));
  jor  g26177(.dina(n26345), .dinb(n26340), .dout(n26346));
  jor  g26178(.dina(n26204), .dinb(n25899), .dout(n26347));
  jand g26179(.dina(n26207), .dinb(n26205), .dout(n26348));
  jnot g26180(.din(n26348), .dout(n26349));
  jand g26181(.dina(n26349), .dinb(n26347), .dout(n26350));
  jand g26182(.dina(n3003), .dinb(n270), .dout(n26351));
  jand g26183(.dina(n26351), .dinb(n16200), .dout(n26352));
  jand g26184(.dina(n8580), .dinb(n519), .dout(n26353));
  jand g26185(.dina(n26353), .dinb(n26352), .dout(n26354));
  jand g26186(.dina(n3380), .dinb(n1708), .dout(n26355));
  jand g26187(.dina(n26355), .dinb(n18357), .dout(n26356));
  jand g26188(.dina(n26356), .dinb(n26354), .dout(n26357));
  jand g26189(.dina(n19835), .dinb(n11386), .dout(n26358));
  jand g26190(.dina(n26358), .dinb(n26357), .dout(n26359));
  jand g26191(.dina(n1731), .dinb(n829), .dout(n26360));
  jand g26192(.dina(n26360), .dinb(n1426), .dout(n26361));
  jand g26193(.dina(n26361), .dinb(n6161), .dout(n26362));
  jand g26194(.dina(n26362), .dinb(n26359), .dout(n26363));
  jand g26195(.dina(n26363), .dinb(n3141), .dout(n26364));
  jnot g26196(.din(n26364), .dout(n26365));
  jxor g26197(.dina(n26365), .dinb(n26350), .dout(n26366));
  jxor g26198(.dina(n26366), .dinb(n26346), .dout(n26367));
  jxor g26199(.dina(n26367), .dinb(n26339), .dout(n26368));
  jand g26200(.dina(n20346), .dinb(n2936), .dout(n26369));
  jand g26201(.dina(n20344), .dinb(n2943), .dout(n26370));
  jand g26202(.dina(n20204), .dinb(n2940), .dout(n26371));
  jand g26203(.dina(n20205), .dinb(n3684), .dout(n26372));
  jor  g26204(.dina(n26372), .dinb(n26371), .dout(n26373));
  jor  g26205(.dina(n26373), .dinb(n26370), .dout(n26374));
  jor  g26206(.dina(n26374), .dinb(n26369), .dout(n26375));
  jxor g26207(.dina(n26375), .dinb(n93), .dout(n26376));
  jxor g26208(.dina(n26376), .dinb(n26368), .dout(n26377));
  jxor g26209(.dina(n26377), .dinb(n26334), .dout(n26378));
  jand g26210(.dina(n21355), .dinb(n71), .dout(n26379));
  jand g26211(.dina(n21197), .dinb(n796), .dout(n26380));
  jand g26212(.dina(n21198), .dinb(n731), .dout(n26381));
  jand g26213(.dina(n20947), .dinb(n1806), .dout(n26382));
  jor  g26214(.dina(n26382), .dinb(n26381), .dout(n26383));
  jor  g26215(.dina(n26383), .dinb(n26380), .dout(n26384));
  jor  g26216(.dina(n26384), .dinb(n26379), .dout(n26385));
  jxor g26217(.dina(n26385), .dinb(n77), .dout(n26386));
  jxor g26218(.dina(n26386), .dinb(n26378), .dout(n26387));
  jxor g26219(.dina(n26387), .dinb(n26329), .dout(n26388));
  jand g26220(.dina(n22291), .dinb(n806), .dout(n26389));
  jand g26221(.dina(n22164), .dinb(n1620), .dout(n26390));
  jand g26222(.dina(n21974), .dinb(n1612), .dout(n26391));
  jand g26223(.dina(n21340), .dinb(n1644), .dout(n26392));
  jor  g26224(.dina(n26392), .dinb(n26391), .dout(n26393));
  jor  g26225(.dina(n26393), .dinb(n26390), .dout(n26394));
  jor  g26226(.dina(n26394), .dinb(n26389), .dout(n26395));
  jxor g26227(.dina(n26395), .dinb(n65), .dout(n26396));
  jxor g26228(.dina(n26396), .dinb(n26388), .dout(n26397));
  jxor g26229(.dina(n26397), .dinb(n26325), .dout(n26398));
  jand g26230(.dina(n22939), .dinb(n1819), .dout(n26399));
  jand g26231(.dina(n22937), .dinb(n2243), .dout(n26400));
  jand g26232(.dina(n22265), .dinb(n2180), .dout(n26401));
  jand g26233(.dina(n22163), .dinb(n2185), .dout(n26402));
  jor  g26234(.dina(n26402), .dinb(n26401), .dout(n26403));
  jor  g26235(.dina(n26403), .dinb(n26400), .dout(n26404));
  jor  g26236(.dina(n26404), .dinb(n26399), .dout(n26405));
  jxor g26237(.dina(n26405), .dinb(n2196), .dout(n26406));
  jxor g26238(.dina(n26406), .dinb(n26398), .dout(n26407));
  jxor g26239(.dina(n26407), .dinb(n26322), .dout(n26408));
  jand g26240(.dina(n23146), .dinb(n2743), .dout(n26409));
  jand g26241(.dina(n23144), .dinb(n2752), .dout(n26410));
  jand g26242(.dina(n23079), .dinb(n2748), .dout(n26411));
  jand g26243(.dina(n23080), .dinb(n2757), .dout(n26412));
  jor  g26244(.dina(n26412), .dinb(n26411), .dout(n26413));
  jor  g26245(.dina(n26413), .dinb(n26410), .dout(n26414));
  jor  g26246(.dina(n26414), .dinb(n26409), .dout(n26415));
  jxor g26247(.dina(n26415), .dinb(n2441), .dout(n26416));
  jxor g26248(.dina(n26416), .dinb(n26408), .dout(n26417));
  jxor g26249(.dina(n26417), .dinb(n26318), .dout(n26418));
  jor  g26250(.dina(n24302), .dinb(n3424), .dout(n26419));
  jor  g26251(.dina(n24304), .dinb(n3426), .dout(n26420));
  jor  g26252(.dina(n24266), .dinb(n3429), .dout(n26421));
  jor  g26253(.dina(n24265), .dinb(n3211), .dout(n26422));
  jand g26254(.dina(n26422), .dinb(n26421), .dout(n26423));
  jand g26255(.dina(n26423), .dinb(n26420), .dout(n26424));
  jand g26256(.dina(n26424), .dinb(n26419), .dout(n26425));
  jxor g26257(.dina(n26425), .dinb(\a[14] ), .dout(n26426));
  jxor g26258(.dina(n26426), .dinb(n26418), .dout(n26427));
  jxor g26259(.dina(n26427), .dinb(n26313), .dout(n26428));
  jor  g26260(.dina(n24932), .dinb(n4023), .dout(n26429));
  jor  g26261(.dina(n24738), .dinb(n4028), .dout(n26430));
  jor  g26262(.dina(n24930), .dinb(n4025), .dout(n26431));
  jand g26263(.dina(n26431), .dinb(n26430), .dout(n26432));
  jor  g26264(.dina(n24518), .dinb(n3871), .dout(n26433));
  jand g26265(.dina(n26433), .dinb(n26432), .dout(n26434));
  jand g26266(.dina(n26434), .dinb(n26429), .dout(n26435));
  jxor g26267(.dina(n26435), .dinb(\a[11] ), .dout(n26436));
  jxor g26268(.dina(n26436), .dinb(n26428), .dout(n26437));
  jxor g26269(.dina(n26437), .dinb(n26309), .dout(n26438));
  jxor g26270(.dina(n26438), .dinb(n26305), .dout(n26439));
  jxor g26271(.dina(n26439), .dinb(n26302), .dout(\result[14] ));
  jand g26272(.dina(n26439), .dinb(n26302), .dout(n26441));
  jnot g26273(.din(n26313), .dout(n26442));
  jand g26274(.dina(n26427), .dinb(n26442), .dout(n26443));
  jor  g26275(.dina(n26436), .dinb(n26428), .dout(n26444));
  jnot g26276(.din(n26444), .dout(n26445));
  jor  g26277(.dina(n26445), .dinb(n26443), .dout(n26446));
  jnot g26278(.din(n26318), .dout(n26447));
  jand g26279(.dina(n26417), .dinb(n26447), .dout(n26448));
  jnot g26280(.din(n26448), .dout(n26449));
  jor  g26281(.dina(n26426), .dinb(n26418), .dout(n26450));
  jand g26282(.dina(n26450), .dinb(n26449), .dout(n26451));
  jor  g26283(.dina(n25116), .dinb(n4023), .dout(n26452));
  jor  g26284(.dina(n24930), .dinb(n19242), .dout(n26453));
  jor  g26285(.dina(n24738), .dinb(n3871), .dout(n26454));
  jand g26286(.dina(n26454), .dinb(n26453), .dout(n26455));
  jand g26287(.dina(n26455), .dinb(n26452), .dout(n26456));
  jxor g26288(.dina(n26456), .dinb(\a[11] ), .dout(n26457));
  jxor g26289(.dina(n26457), .dinb(n26451), .dout(n26458));
  jnot g26290(.din(n26322), .dout(n26459));
  jand g26291(.dina(n26407), .dinb(n26459), .dout(n26460));
  jnot g26292(.din(n26460), .dout(n26461));
  jor  g26293(.dina(n26416), .dinb(n26408), .dout(n26462));
  jand g26294(.dina(n26462), .dinb(n26461), .dout(n26463));
  jnot g26295(.din(n26325), .dout(n26464));
  jand g26296(.dina(n26397), .dinb(n26464), .dout(n26465));
  jnot g26297(.din(n26465), .dout(n26466));
  jor  g26298(.dina(n26406), .dinb(n26398), .dout(n26467));
  jand g26299(.dina(n26467), .dinb(n26466), .dout(n26468));
  jnot g26300(.din(n26329), .dout(n26469));
  jand g26301(.dina(n26387), .dinb(n26469), .dout(n26470));
  jnot g26302(.din(n26470), .dout(n26471));
  jor  g26303(.dina(n26396), .dinb(n26388), .dout(n26472));
  jand g26304(.dina(n26472), .dinb(n26471), .dout(n26473));
  jnot g26305(.din(n26334), .dout(n26474));
  jand g26306(.dina(n26377), .dinb(n26474), .dout(n26475));
  jnot g26307(.din(n26475), .dout(n26476));
  jor  g26308(.dina(n26386), .dinb(n26378), .dout(n26477));
  jand g26309(.dina(n26477), .dinb(n26476), .dout(n26478));
  jnot g26310(.din(n26339), .dout(n26479));
  jand g26311(.dina(n26367), .dinb(n26479), .dout(n26480));
  jnot g26312(.din(n26480), .dout(n26481));
  jor  g26313(.dina(n26376), .dinb(n26368), .dout(n26482));
  jand g26314(.dina(n26482), .dinb(n26481), .dout(n26483));
  jand g26315(.dina(n20371), .dinb(n5076), .dout(n26484));
  jand g26316(.dina(n20205), .dinb(n5084), .dout(n26485));
  jand g26317(.dina(n19922), .dinb(n5082), .dout(n26486));
  jand g26318(.dina(n19373), .dinb(n6050), .dout(n26487));
  jor  g26319(.dina(n26487), .dinb(n26486), .dout(n26488));
  jor  g26320(.dina(n26488), .dinb(n26485), .dout(n26489));
  jor  g26321(.dina(n26489), .dinb(n26484), .dout(n26490));
  jnot g26322(.din(n26350), .dout(n26491));
  jand g26323(.dina(n26364), .dinb(n26491), .dout(n26492));
  jand g26324(.dina(n26366), .dinb(n26346), .dout(n26493));
  jor  g26325(.dina(n26493), .dinb(n26492), .dout(n26494));
  jand g26326(.dina(n25882), .dinb(n2521), .dout(n26495));
  jand g26327(.dina(n26495), .dinb(n10159), .dout(n26496));
  jand g26328(.dina(n5396), .dinb(n2367), .dout(n26497));
  jand g26329(.dina(n2587), .dinb(n1822), .dout(n26498));
  jand g26330(.dina(n26498), .dinb(n26497), .dout(n26499));
  jand g26331(.dina(n26499), .dinb(n110), .dout(n26500));
  jand g26332(.dina(n557), .dinb(n266), .dout(n26501));
  jand g26333(.dina(n589), .dinb(n1160), .dout(n26502));
  jand g26334(.dina(n26502), .dinb(n26501), .dout(n26503));
  jand g26335(.dina(n26503), .dinb(n645), .dout(n26504));
  jand g26336(.dina(n26504), .dinb(n16789), .dout(n26505));
  jand g26337(.dina(n26505), .dinb(n26500), .dout(n26506));
  jand g26338(.dina(n2600), .dinb(n1516), .dout(n26507));
  jand g26339(.dina(n26507), .dinb(n20865), .dout(n26508));
  jand g26340(.dina(n1714), .dinb(n880), .dout(n26509));
  jand g26341(.dina(n26509), .dinb(n26508), .dout(n26510));
  jand g26342(.dina(n26510), .dinb(n26506), .dout(n26511));
  jand g26343(.dina(n26511), .dinb(n26496), .dout(n26512));
  jxor g26344(.dina(n26512), .dinb(n26365), .dout(n26513));
  jxor g26345(.dina(n26513), .dinb(n26494), .dout(n26514));
  jxor g26346(.dina(n26514), .dinb(n26490), .dout(n26515));
  jnot g26347(.din(n26515), .dout(n26516));
  jand g26348(.dina(n20949), .dinb(n2936), .dout(n26517));
  jand g26349(.dina(n20947), .dinb(n2943), .dout(n26518));
  jand g26350(.dina(n20344), .dinb(n2940), .dout(n26519));
  jand g26351(.dina(n20204), .dinb(n3684), .dout(n26520));
  jor  g26352(.dina(n26520), .dinb(n26519), .dout(n26521));
  jor  g26353(.dina(n26521), .dinb(n26518), .dout(n26522));
  jor  g26354(.dina(n26522), .dinb(n26517), .dout(n26523));
  jxor g26355(.dina(n26523), .dinb(n93), .dout(n26524));
  jxor g26356(.dina(n26524), .dinb(n26516), .dout(n26525));
  jxor g26357(.dina(n26525), .dinb(n26483), .dout(n26526));
  jand g26358(.dina(n21342), .dinb(n71), .dout(n26527));
  jand g26359(.dina(n21340), .dinb(n796), .dout(n26528));
  jand g26360(.dina(n21197), .dinb(n731), .dout(n26529));
  jand g26361(.dina(n21198), .dinb(n1806), .dout(n26530));
  jor  g26362(.dina(n26530), .dinb(n26529), .dout(n26531));
  jor  g26363(.dina(n26531), .dinb(n26528), .dout(n26532));
  jor  g26364(.dina(n26532), .dinb(n26527), .dout(n26533));
  jxor g26365(.dina(n26533), .dinb(n77), .dout(n26534));
  jxor g26366(.dina(n26534), .dinb(n26526), .dout(n26535));
  jxor g26367(.dina(n26535), .dinb(n26478), .dout(n26536));
  jand g26368(.dina(n22279), .dinb(n806), .dout(n26537));
  jand g26369(.dina(n22164), .dinb(n1612), .dout(n26538));
  jand g26370(.dina(n22163), .dinb(n1620), .dout(n26539));
  jor  g26371(.dina(n26539), .dinb(n26538), .dout(n26540));
  jand g26372(.dina(n21974), .dinb(n1644), .dout(n26541));
  jor  g26373(.dina(n26541), .dinb(n26540), .dout(n26542));
  jor  g26374(.dina(n26542), .dinb(n26537), .dout(n26543));
  jxor g26375(.dina(n26543), .dinb(n65), .dout(n26544));
  jxor g26376(.dina(n26544), .dinb(n26536), .dout(n26545));
  jxor g26377(.dina(n26545), .dinb(n26473), .dout(n26546));
  jand g26378(.dina(n23172), .dinb(n1819), .dout(n26547));
  jand g26379(.dina(n23080), .dinb(n2243), .dout(n26548));
  jand g26380(.dina(n22937), .dinb(n2180), .dout(n26549));
  jand g26381(.dina(n22265), .dinb(n2185), .dout(n26550));
  jor  g26382(.dina(n26550), .dinb(n26549), .dout(n26551));
  jor  g26383(.dina(n26551), .dinb(n26548), .dout(n26552));
  jor  g26384(.dina(n26552), .dinb(n26547), .dout(n26553));
  jxor g26385(.dina(n26553), .dinb(n2196), .dout(n26554));
  jxor g26386(.dina(n26554), .dinb(n26546), .dout(n26555));
  jxor g26387(.dina(n26555), .dinb(n26468), .dout(n26556));
  jand g26388(.dina(n23847), .dinb(n2743), .dout(n26557));
  jand g26389(.dina(n23845), .dinb(n2752), .dout(n26558));
  jand g26390(.dina(n23144), .dinb(n2748), .dout(n26559));
  jand g26391(.dina(n23079), .dinb(n2757), .dout(n26560));
  jor  g26392(.dina(n26560), .dinb(n26559), .dout(n26561));
  jor  g26393(.dina(n26561), .dinb(n26558), .dout(n26562));
  jor  g26394(.dina(n26562), .dinb(n26557), .dout(n26563));
  jxor g26395(.dina(n26563), .dinb(n2441), .dout(n26564));
  jxor g26396(.dina(n26564), .dinb(n26556), .dout(n26565));
  jxor g26397(.dina(n26565), .dinb(n26463), .dout(n26566));
  jor  g26398(.dina(n24516), .dinb(n3424), .dout(n26567));
  jor  g26399(.dina(n24518), .dinb(n3426), .dout(n26568));
  jor  g26400(.dina(n24304), .dinb(n3429), .dout(n26569));
  jor  g26401(.dina(n24266), .dinb(n3211), .dout(n26570));
  jand g26402(.dina(n26570), .dinb(n26569), .dout(n26571));
  jand g26403(.dina(n26571), .dinb(n26568), .dout(n26572));
  jand g26404(.dina(n26572), .dinb(n26567), .dout(n26573));
  jxor g26405(.dina(n26573), .dinb(\a[14] ), .dout(n26574));
  jxor g26406(.dina(n26574), .dinb(n26566), .dout(n26575));
  jxor g26407(.dina(n26575), .dinb(n26458), .dout(n26576));
  jxor g26408(.dina(n26576), .dinb(n26446), .dout(n26577));
  jand g26409(.dina(n26437), .dinb(n26309), .dout(n26578));
  jand g26410(.dina(n26438), .dinb(n26305), .dout(n26579));
  jor  g26411(.dina(n26579), .dinb(n26578), .dout(n26580));
  jxor g26412(.dina(n26580), .dinb(n26577), .dout(n26581));
  jxor g26413(.dina(n26581), .dinb(n26441), .dout(\result[15] ));
  jand g26414(.dina(n26581), .dinb(n26441), .dout(n26583));
  jand g26415(.dina(n26576), .dinb(n26446), .dout(n26584));
  jand g26416(.dina(n26580), .dinb(n26577), .dout(n26585));
  jor  g26417(.dina(n26585), .dinb(n26584), .dout(n26586));
  jor  g26418(.dina(n26457), .dinb(n26451), .dout(n26587));
  jnot g26419(.din(n26587), .dout(n26588));
  jand g26420(.dina(n26575), .dinb(n26458), .dout(n26589));
  jor  g26421(.dina(n26589), .dinb(n26588), .dout(n26590));
  jnot g26422(.din(n26468), .dout(n26591));
  jand g26423(.dina(n26555), .dinb(n26591), .dout(n26592));
  jnot g26424(.din(n26592), .dout(n26593));
  jor  g26425(.dina(n26564), .dinb(n26556), .dout(n26594));
  jand g26426(.dina(n26594), .dinb(n26593), .dout(n26595));
  jnot g26427(.din(n26478), .dout(n26596));
  jand g26428(.dina(n26535), .dinb(n26596), .dout(n26597));
  jnot g26429(.din(n26597), .dout(n26598));
  jor  g26430(.dina(n26544), .dinb(n26536), .dout(n26599));
  jand g26431(.dina(n26599), .dinb(n26598), .dout(n26600));
  jnot g26432(.din(n26483), .dout(n26601));
  jand g26433(.dina(n26525), .dinb(n26601), .dout(n26602));
  jnot g26434(.din(n26602), .dout(n26603));
  jor  g26435(.dina(n26534), .dinb(n26526), .dout(n26604));
  jand g26436(.dina(n26604), .dinb(n26603), .dout(n26605));
  jnot g26437(.din(n26605), .dout(n26606));
  jand g26438(.dina(n26514), .dinb(n26490), .dout(n26607));
  jnot g26439(.din(n26607), .dout(n26608));
  jor  g26440(.dina(n26524), .dinb(n26516), .dout(n26609));
  jand g26441(.dina(n26609), .dinb(n26608), .dout(n26610));
  jnot g26442(.din(n26610), .dout(n26611));
  jor  g26443(.dina(n26512), .dinb(n26365), .dout(n26612));
  jand g26444(.dina(n26513), .dinb(n26494), .dout(n26613));
  jnot g26445(.din(n26613), .dout(n26614));
  jand g26446(.dina(n26614), .dinb(n26612), .dout(n26615));
  jnot g26447(.din(n26615), .dout(n26616));
  jand g26448(.dina(n2169), .dinb(n114), .dout(n26617));
  jand g26449(.dina(n26617), .dinb(n2092), .dout(n26618));
  jand g26450(.dina(n10379), .dinb(n270), .dout(n26619));
  jand g26451(.dina(n26619), .dinb(n26618), .dout(n26620));
  jand g26452(.dina(n2052), .dinb(n1379), .dout(n26621));
  jand g26453(.dina(n26621), .dinb(n10383), .dout(n26622));
  jand g26454(.dina(n6439), .dinb(n553), .dout(n26623));
  jand g26455(.dina(n26623), .dinb(n874), .dout(n26624));
  jand g26456(.dina(n26624), .dinb(n26622), .dout(n26625));
  jand g26457(.dina(n3150), .dinb(n2020), .dout(n26626));
  jand g26458(.dina(n26626), .dinb(n1098), .dout(n26627));
  jand g26459(.dina(n26627), .dinb(n2586), .dout(n26628));
  jand g26460(.dina(n26628), .dinb(n26625), .dout(n26629));
  jand g26461(.dina(n26629), .dinb(n5461), .dout(n26630));
  jand g26462(.dina(n26630), .dinb(n3757), .dout(n26631));
  jand g26463(.dina(n26631), .dinb(n26620), .dout(n26632));
  jxor g26464(.dina(n26632), .dinb(n26364), .dout(n26633));
  jand g26465(.dina(n25199), .dinb(n19847), .dout(n26634));
  jxor g26466(.dina(n26634), .dinb(n4050), .dout(n26635));
  jxor g26467(.dina(n26635), .dinb(n26633), .dout(n26636));
  jand g26468(.dina(n20358), .dinb(n5076), .dout(n26637));
  jand g26469(.dina(n20204), .dinb(n5084), .dout(n26638));
  jand g26470(.dina(n20205), .dinb(n5082), .dout(n26639));
  jand g26471(.dina(n19922), .dinb(n6050), .dout(n26640));
  jor  g26472(.dina(n26640), .dinb(n26639), .dout(n26641));
  jor  g26473(.dina(n26641), .dinb(n26638), .dout(n26642));
  jor  g26474(.dina(n26642), .dinb(n26637), .dout(n26643));
  jxor g26475(.dina(n26643), .dinb(n26636), .dout(n26644));
  jxor g26476(.dina(n26644), .dinb(n26616), .dout(n26645));
  jxor g26477(.dina(n26645), .dinb(n26611), .dout(n26646));
  jnot g26478(.din(n26646), .dout(n26647));
  jand g26479(.dina(n21367), .dinb(n2936), .dout(n26648));
  jand g26480(.dina(n21198), .dinb(n2943), .dout(n26649));
  jand g26481(.dina(n20947), .dinb(n2940), .dout(n26650));
  jand g26482(.dina(n20344), .dinb(n3684), .dout(n26651));
  jor  g26483(.dina(n26651), .dinb(n26650), .dout(n26652));
  jor  g26484(.dina(n26652), .dinb(n26649), .dout(n26653));
  jor  g26485(.dina(n26653), .dinb(n26648), .dout(n26654));
  jxor g26486(.dina(n26654), .dinb(n93), .dout(n26655));
  jxor g26487(.dina(n26655), .dinb(n26647), .dout(n26656));
  jnot g26488(.din(n26656), .dout(n26657));
  jand g26489(.dina(n21976), .dinb(n71), .dout(n26658));
  jand g26490(.dina(n21974), .dinb(n796), .dout(n26659));
  jand g26491(.dina(n21340), .dinb(n731), .dout(n26660));
  jand g26492(.dina(n21197), .dinb(n1806), .dout(n26661));
  jor  g26493(.dina(n26661), .dinb(n26660), .dout(n26662));
  jor  g26494(.dina(n26662), .dinb(n26659), .dout(n26663));
  jor  g26495(.dina(n26663), .dinb(n26658), .dout(n26664));
  jxor g26496(.dina(n26664), .dinb(n77), .dout(n26665));
  jxor g26497(.dina(n26665), .dinb(n26657), .dout(n26666));
  jxor g26498(.dina(n26666), .dinb(n26606), .dout(n26667));
  jand g26499(.dina(n22267), .dinb(n806), .dout(n26668));
  jand g26500(.dina(n22163), .dinb(n1612), .dout(n26669));
  jand g26501(.dina(n22265), .dinb(n1620), .dout(n26670));
  jor  g26502(.dina(n26670), .dinb(n26669), .dout(n26671));
  jand g26503(.dina(n22164), .dinb(n1644), .dout(n26672));
  jor  g26504(.dina(n26672), .dinb(n26671), .dout(n26673));
  jor  g26505(.dina(n26673), .dinb(n26668), .dout(n26674));
  jxor g26506(.dina(n26674), .dinb(n65), .dout(n26675));
  jxor g26507(.dina(n26675), .dinb(n26667), .dout(n26676));
  jxor g26508(.dina(n26676), .dinb(n26600), .dout(n26677));
  jnot g26509(.din(n26473), .dout(n26678));
  jand g26510(.dina(n26545), .dinb(n26678), .dout(n26679));
  jnot g26511(.din(n26679), .dout(n26680));
  jor  g26512(.dina(n26554), .dinb(n26546), .dout(n26681));
  jand g26513(.dina(n26681), .dinb(n26680), .dout(n26682));
  jand g26514(.dina(n23159), .dinb(n1819), .dout(n26683));
  jand g26515(.dina(n23080), .dinb(n2180), .dout(n26684));
  jand g26516(.dina(n23079), .dinb(n2243), .dout(n26685));
  jor  g26517(.dina(n26685), .dinb(n26684), .dout(n26686));
  jand g26518(.dina(n22937), .dinb(n2185), .dout(n26687));
  jor  g26519(.dina(n26687), .dinb(n26686), .dout(n26688));
  jor  g26520(.dina(n26688), .dinb(n26683), .dout(n26689));
  jxor g26521(.dina(n26689), .dinb(n2196), .dout(n26690));
  jxor g26522(.dina(n26690), .dinb(n26682), .dout(n26691));
  jxor g26523(.dina(n26691), .dinb(n26677), .dout(n26692));
  jand g26524(.dina(n24077), .dinb(n2743), .dout(n26693));
  jand g26525(.dina(n23845), .dinb(n2748), .dout(n26694));
  jand g26526(.dina(n24075), .dinb(n2752), .dout(n26695));
  jor  g26527(.dina(n26695), .dinb(n26694), .dout(n26696));
  jand g26528(.dina(n23144), .dinb(n2757), .dout(n26697));
  jor  g26529(.dina(n26697), .dinb(n26696), .dout(n26698));
  jor  g26530(.dina(n26698), .dinb(n26693), .dout(n26699));
  jxor g26531(.dina(n26699), .dinb(n2441), .dout(n26700));
  jxor g26532(.dina(n26700), .dinb(n26692), .dout(n26701));
  jxor g26533(.dina(n26701), .dinb(n26595), .dout(n26702));
  jnot g26534(.din(n26463), .dout(n26703));
  jand g26535(.dina(n26565), .dinb(n26703), .dout(n26704));
  jnot g26536(.din(n26704), .dout(n26705));
  jor  g26537(.dina(n26574), .dinb(n26566), .dout(n26706));
  jand g26538(.dina(n26706), .dinb(n26705), .dout(n26707));
  jor  g26539(.dina(n24736), .dinb(n3424), .dout(n26708));
  jor  g26540(.dina(n24738), .dinb(n3426), .dout(n26709));
  jor  g26541(.dina(n24518), .dinb(n3429), .dout(n26710));
  jor  g26542(.dina(n24304), .dinb(n3211), .dout(n26711));
  jand g26543(.dina(n26711), .dinb(n26710), .dout(n26712));
  jand g26544(.dina(n26712), .dinb(n26709), .dout(n26713));
  jand g26545(.dina(n26713), .dinb(n26708), .dout(n26714));
  jxor g26546(.dina(n26714), .dinb(\a[14] ), .dout(n26715));
  jxor g26547(.dina(n26715), .dinb(n26707), .dout(n26716));
  jxor g26548(.dina(n26716), .dinb(n26702), .dout(n26717));
  jxor g26549(.dina(n26717), .dinb(n26590), .dout(n26718));
  jxor g26550(.dina(n26718), .dinb(n26586), .dout(n26719));
  jxor g26551(.dina(n26719), .dinb(n26583), .dout(\result[16] ));
  jand g26552(.dina(n26719), .dinb(n26583), .dout(n26721));
  jand g26553(.dina(n26717), .dinb(n26590), .dout(n26722));
  jand g26554(.dina(n26718), .dinb(n26586), .dout(n26723));
  jor  g26555(.dina(n26723), .dinb(n26722), .dout(n26724));
  jor  g26556(.dina(n26715), .dinb(n26707), .dout(n26725));
  jnot g26557(.din(n26725), .dout(n26726));
  jand g26558(.dina(n26716), .dinb(n26702), .dout(n26727));
  jor  g26559(.dina(n26727), .dinb(n26726), .dout(n26728));
  jnot g26560(.din(n26692), .dout(n26729));
  jor  g26561(.dina(n26700), .dinb(n26729), .dout(n26730));
  jor  g26562(.dina(n26701), .dinb(n26595), .dout(n26731));
  jand g26563(.dina(n26731), .dinb(n26730), .dout(n26732));
  jor  g26564(.dina(n26690), .dinb(n26682), .dout(n26733));
  jand g26565(.dina(n26691), .dinb(n26677), .dout(n26734));
  jnot g26566(.din(n26734), .dout(n26735));
  jand g26567(.dina(n26735), .dinb(n26733), .dout(n26736));
  jnot g26568(.din(n26667), .dout(n26737));
  jor  g26569(.dina(n26675), .dinb(n26737), .dout(n26738));
  jor  g26570(.dina(n26676), .dinb(n26600), .dout(n26739));
  jand g26571(.dina(n26739), .dinb(n26738), .dout(n26740));
  jor  g26572(.dina(n26665), .dinb(n26657), .dout(n26741));
  jand g26573(.dina(n26666), .dinb(n26606), .dout(n26742));
  jnot g26574(.din(n26742), .dout(n26743));
  jand g26575(.dina(n26743), .dinb(n26741), .dout(n26744));
  jand g26576(.dina(n26645), .dinb(n26611), .dout(n26745));
  jnot g26577(.din(n26745), .dout(n26746));
  jor  g26578(.dina(n26655), .dinb(n26647), .dout(n26747));
  jand g26579(.dina(n26747), .dinb(n26746), .dout(n26748));
  jnot g26580(.din(n26748), .dout(n26749));
  jand g26581(.dina(n26643), .dinb(n26636), .dout(n26750));
  jand g26582(.dina(n26644), .dinb(n26616), .dout(n26751));
  jor  g26583(.dina(n26751), .dinb(n26750), .dout(n26752));
  jand g26584(.dina(n20346), .dinb(n5076), .dout(n26753));
  jand g26585(.dina(n20344), .dinb(n5084), .dout(n26754));
  jand g26586(.dina(n20204), .dinb(n5082), .dout(n26755));
  jand g26587(.dina(n20205), .dinb(n6050), .dout(n26756));
  jor  g26588(.dina(n26756), .dinb(n26755), .dout(n26757));
  jor  g26589(.dina(n26757), .dinb(n26754), .dout(n26758));
  jor  g26590(.dina(n26758), .dinb(n26753), .dout(n26759));
  jor  g26591(.dina(n26632), .dinb(n26364), .dout(n26760));
  jand g26592(.dina(n26635), .dinb(n26633), .dout(n26761));
  jnot g26593(.din(n26761), .dout(n26762));
  jand g26594(.dina(n26762), .dinb(n26760), .dout(n26763));
  jand g26595(.dina(n934), .dinb(n1393), .dout(n26764));
  jand g26596(.dina(n26764), .dinb(n1687), .dout(n26765));
  jand g26597(.dina(n1327), .dinb(n542), .dout(n26766));
  jand g26598(.dina(n26766), .dinb(n1744), .dout(n26767));
  jand g26599(.dina(n26767), .dinb(n26765), .dout(n26768));
  jand g26600(.dina(n7230), .dinb(n676), .dout(n26769));
  jand g26601(.dina(n26769), .dinb(n3389), .dout(n26770));
  jand g26602(.dina(n21918), .dinb(n5222), .dout(n26771));
  jand g26603(.dina(n26771), .dinb(n26770), .dout(n26772));
  jand g26604(.dina(n26772), .dinb(n26768), .dout(n26773));
  jand g26605(.dina(n26773), .dinb(n24601), .dout(n26774));
  jand g26606(.dina(n25006), .dinb(n22028), .dout(n26775));
  jand g26607(.dina(n26775), .dinb(n16793), .dout(n26776));
  jand g26608(.dina(n26776), .dinb(n26774), .dout(n26777));
  jnot g26609(.din(n26777), .dout(n26778));
  jxor g26610(.dina(n26778), .dinb(n26763), .dout(n26779));
  jxor g26611(.dina(n26779), .dinb(n26759), .dout(n26780));
  jxor g26612(.dina(n26780), .dinb(n26752), .dout(n26781));
  jnot g26613(.din(n26781), .dout(n26782));
  jand g26614(.dina(n21355), .dinb(n2936), .dout(n26783));
  jand g26615(.dina(n21198), .dinb(n2940), .dout(n26784));
  jand g26616(.dina(n21197), .dinb(n2943), .dout(n26785));
  jor  g26617(.dina(n26785), .dinb(n26784), .dout(n26786));
  jand g26618(.dina(n20947), .dinb(n3684), .dout(n26787));
  jor  g26619(.dina(n26787), .dinb(n26786), .dout(n26788));
  jor  g26620(.dina(n26788), .dinb(n26783), .dout(n26789));
  jxor g26621(.dina(n26789), .dinb(n93), .dout(n26790));
  jxor g26622(.dina(n26790), .dinb(n26782), .dout(n26791));
  jxor g26623(.dina(n26791), .dinb(n26749), .dout(n26792));
  jnot g26624(.din(n26792), .dout(n26793));
  jand g26625(.dina(n22291), .dinb(n71), .dout(n26794));
  jand g26626(.dina(n22164), .dinb(n796), .dout(n26795));
  jand g26627(.dina(n21974), .dinb(n731), .dout(n26796));
  jand g26628(.dina(n21340), .dinb(n1806), .dout(n26797));
  jor  g26629(.dina(n26797), .dinb(n26796), .dout(n26798));
  jor  g26630(.dina(n26798), .dinb(n26795), .dout(n26799));
  jor  g26631(.dina(n26799), .dinb(n26794), .dout(n26800));
  jxor g26632(.dina(n26800), .dinb(n77), .dout(n26801));
  jxor g26633(.dina(n26801), .dinb(n26793), .dout(n26802));
  jxor g26634(.dina(n26802), .dinb(n26744), .dout(n26803));
  jand g26635(.dina(n22939), .dinb(n806), .dout(n26804));
  jand g26636(.dina(n22937), .dinb(n1620), .dout(n26805));
  jand g26637(.dina(n22265), .dinb(n1612), .dout(n26806));
  jand g26638(.dina(n22163), .dinb(n1644), .dout(n26807));
  jor  g26639(.dina(n26807), .dinb(n26806), .dout(n26808));
  jor  g26640(.dina(n26808), .dinb(n26805), .dout(n26809));
  jor  g26641(.dina(n26809), .dinb(n26804), .dout(n26810));
  jxor g26642(.dina(n26810), .dinb(n65), .dout(n26811));
  jxor g26643(.dina(n26811), .dinb(n26803), .dout(n26812));
  jxor g26644(.dina(n26812), .dinb(n26740), .dout(n26813));
  jand g26645(.dina(n23146), .dinb(n1819), .dout(n26814));
  jand g26646(.dina(n23079), .dinb(n2180), .dout(n26815));
  jand g26647(.dina(n23144), .dinb(n2243), .dout(n26816));
  jor  g26648(.dina(n26816), .dinb(n26815), .dout(n26817));
  jand g26649(.dina(n23080), .dinb(n2185), .dout(n26818));
  jor  g26650(.dina(n26818), .dinb(n26817), .dout(n26819));
  jor  g26651(.dina(n26819), .dinb(n26814), .dout(n26820));
  jxor g26652(.dina(n26820), .dinb(n2196), .dout(n26821));
  jxor g26653(.dina(n26821), .dinb(n26813), .dout(n26822));
  jxor g26654(.dina(n26822), .dinb(n26736), .dout(n26823));
  jor  g26655(.dina(n24302), .dinb(n2744), .dout(n26824));
  jor  g26656(.dina(n24304), .dinb(n2753), .dout(n26825));
  jor  g26657(.dina(n24266), .dinb(n2749), .dout(n26826));
  jor  g26658(.dina(n24265), .dinb(n2758), .dout(n26827));
  jand g26659(.dina(n26827), .dinb(n26826), .dout(n26828));
  jand g26660(.dina(n26828), .dinb(n26825), .dout(n26829));
  jand g26661(.dina(n26829), .dinb(n26824), .dout(n26830));
  jxor g26662(.dina(n26830), .dinb(\a[17] ), .dout(n26831));
  jxor g26663(.dina(n26831), .dinb(n26823), .dout(n26832));
  jxor g26664(.dina(n26832), .dinb(n26732), .dout(n26833));
  jor  g26665(.dina(n24932), .dinb(n3424), .dout(n26834));
  jor  g26666(.dina(n24738), .dinb(n3429), .dout(n26835));
  jor  g26667(.dina(n24930), .dinb(n3426), .dout(n26836));
  jand g26668(.dina(n26836), .dinb(n26835), .dout(n26837));
  jor  g26669(.dina(n24518), .dinb(n3211), .dout(n26838));
  jand g26670(.dina(n26838), .dinb(n26837), .dout(n26839));
  jand g26671(.dina(n26839), .dinb(n26834), .dout(n26840));
  jxor g26672(.dina(n26840), .dinb(\a[14] ), .dout(n26841));
  jxor g26673(.dina(n26841), .dinb(n26833), .dout(n26842));
  jxor g26674(.dina(n26842), .dinb(n26728), .dout(n26843));
  jxor g26675(.dina(n26843), .dinb(n26724), .dout(n26844));
  jxor g26676(.dina(n26844), .dinb(n26721), .dout(\result[17] ));
  jand g26677(.dina(n26844), .dinb(n26721), .dout(n26846));
  jnot g26678(.din(n26732), .dout(n26847));
  jand g26679(.dina(n26832), .dinb(n26847), .dout(n26848));
  jnot g26680(.din(n26848), .dout(n26849));
  jor  g26681(.dina(n26841), .dinb(n26833), .dout(n26850));
  jand g26682(.dina(n26850), .dinb(n26849), .dout(n26851));
  jnot g26683(.din(n26851), .dout(n26852));
  jnot g26684(.din(n26736), .dout(n26853));
  jand g26685(.dina(n26822), .dinb(n26853), .dout(n26854));
  jnot g26686(.din(n26854), .dout(n26855));
  jor  g26687(.dina(n26831), .dinb(n26823), .dout(n26856));
  jand g26688(.dina(n26856), .dinb(n26855), .dout(n26857));
  jor  g26689(.dina(n25116), .dinb(n3424), .dout(n26858));
  jor  g26690(.dina(n24930), .dinb(n20060), .dout(n26859));
  jor  g26691(.dina(n24738), .dinb(n3211), .dout(n26860));
  jand g26692(.dina(n26860), .dinb(n26859), .dout(n26861));
  jand g26693(.dina(n26861), .dinb(n26858), .dout(n26862));
  jxor g26694(.dina(n26862), .dinb(\a[14] ), .dout(n26863));
  jxor g26695(.dina(n26863), .dinb(n26857), .dout(n26864));
  jnot g26696(.din(n26740), .dout(n26865));
  jand g26697(.dina(n26812), .dinb(n26865), .dout(n26866));
  jnot g26698(.din(n26866), .dout(n26867));
  jor  g26699(.dina(n26821), .dinb(n26813), .dout(n26868));
  jand g26700(.dina(n26868), .dinb(n26867), .dout(n26869));
  jnot g26701(.din(n26869), .dout(n26870));
  jnot g26702(.din(n26744), .dout(n26871));
  jand g26703(.dina(n26802), .dinb(n26871), .dout(n26872));
  jnot g26704(.din(n26872), .dout(n26873));
  jor  g26705(.dina(n26811), .dinb(n26803), .dout(n26874));
  jand g26706(.dina(n26874), .dinb(n26873), .dout(n26875));
  jand g26707(.dina(n26791), .dinb(n26749), .dout(n26876));
  jnot g26708(.din(n26876), .dout(n26877));
  jor  g26709(.dina(n26801), .dinb(n26793), .dout(n26878));
  jand g26710(.dina(n26878), .dinb(n26877), .dout(n26879));
  jnot g26711(.din(n26879), .dout(n26880));
  jnot g26712(.din(n26763), .dout(n26881));
  jand g26713(.dina(n26777), .dinb(n26881), .dout(n26882));
  jand g26714(.dina(n26779), .dinb(n26759), .dout(n26883));
  jor  g26715(.dina(n26883), .dinb(n26882), .dout(n26884));
  jand g26716(.dina(n20949), .dinb(n5076), .dout(n26885));
  jand g26717(.dina(n20947), .dinb(n5084), .dout(n26886));
  jand g26718(.dina(n20344), .dinb(n5082), .dout(n26887));
  jand g26719(.dina(n20204), .dinb(n6050), .dout(n26888));
  jor  g26720(.dina(n26888), .dinb(n26887), .dout(n26889));
  jor  g26721(.dina(n26889), .dinb(n26886), .dout(n26890));
  jor  g26722(.dina(n26890), .dinb(n26885), .dout(n26891));
  jand g26723(.dina(n1237), .dinb(n171), .dout(n26892));
  jand g26724(.dina(n26892), .dinb(n1437), .dout(n26893));
  jand g26725(.dina(n1495), .dinb(n1289), .dout(n26894));
  jand g26726(.dina(n26894), .dinb(n26893), .dout(n26895));
  jand g26727(.dina(n26895), .dinb(n2151), .dout(n26896));
  jand g26728(.dina(n8589), .dinb(n3198), .dout(n26897));
  jand g26729(.dina(n6283), .dinb(n829), .dout(n26898));
  jand g26730(.dina(n26898), .dinb(n1327), .dout(n26899));
  jand g26731(.dina(n26899), .dinb(n26897), .dout(n26900));
  jand g26732(.dina(n26900), .dinb(n26896), .dout(n26901));
  jand g26733(.dina(n26901), .dinb(n1588), .dout(n26902));
  jand g26734(.dina(n26902), .dinb(n12465), .dout(n26903));
  jand g26735(.dina(n15290), .dinb(n6304), .dout(n26904));
  jand g26736(.dina(n14206), .dinb(n7789), .dout(n26905));
  jand g26737(.dina(n26905), .dinb(n26904), .dout(n26906));
  jand g26738(.dina(n26906), .dinb(n26903), .dout(n26907));
  jxor g26739(.dina(n26907), .dinb(n26778), .dout(n26908));
  jxor g26740(.dina(n26908), .dinb(n26891), .dout(n26909));
  jxor g26741(.dina(n26909), .dinb(n26884), .dout(n26910));
  jnot g26742(.din(n26910), .dout(n26911));
  jand g26743(.dina(n26780), .dinb(n26752), .dout(n26912));
  jnot g26744(.din(n26912), .dout(n26913));
  jor  g26745(.dina(n26790), .dinb(n26782), .dout(n26914));
  jand g26746(.dina(n26914), .dinb(n26913), .dout(n26915));
  jxor g26747(.dina(n26915), .dinb(n26911), .dout(n26916));
  jnot g26748(.din(n26916), .dout(n26917));
  jand g26749(.dina(n21342), .dinb(n2936), .dout(n26918));
  jand g26750(.dina(n21197), .dinb(n2940), .dout(n26919));
  jand g26751(.dina(n21340), .dinb(n2943), .dout(n26920));
  jor  g26752(.dina(n26920), .dinb(n26919), .dout(n26921));
  jand g26753(.dina(n21198), .dinb(n3684), .dout(n26922));
  jor  g26754(.dina(n26922), .dinb(n26921), .dout(n26923));
  jor  g26755(.dina(n26923), .dinb(n26918), .dout(n26924));
  jxor g26756(.dina(n26924), .dinb(n93), .dout(n26925));
  jxor g26757(.dina(n26925), .dinb(n26917), .dout(n26926));
  jnot g26758(.din(n26926), .dout(n26927));
  jand g26759(.dina(n22279), .dinb(n71), .dout(n26928));
  jand g26760(.dina(n22163), .dinb(n796), .dout(n26929));
  jand g26761(.dina(n22164), .dinb(n731), .dout(n26930));
  jand g26762(.dina(n21974), .dinb(n1806), .dout(n26931));
  jor  g26763(.dina(n26931), .dinb(n26930), .dout(n26932));
  jor  g26764(.dina(n26932), .dinb(n26929), .dout(n26933));
  jor  g26765(.dina(n26933), .dinb(n26928), .dout(n26934));
  jxor g26766(.dina(n26934), .dinb(n77), .dout(n26935));
  jxor g26767(.dina(n26935), .dinb(n26927), .dout(n26936));
  jxor g26768(.dina(n26936), .dinb(n26880), .dout(n26937));
  jnot g26769(.din(n26937), .dout(n26938));
  jand g26770(.dina(n23172), .dinb(n806), .dout(n26939));
  jand g26771(.dina(n23080), .dinb(n1620), .dout(n26940));
  jand g26772(.dina(n22937), .dinb(n1612), .dout(n26941));
  jand g26773(.dina(n22265), .dinb(n1644), .dout(n26942));
  jor  g26774(.dina(n26942), .dinb(n26941), .dout(n26943));
  jor  g26775(.dina(n26943), .dinb(n26940), .dout(n26944));
  jor  g26776(.dina(n26944), .dinb(n26939), .dout(n26945));
  jxor g26777(.dina(n26945), .dinb(n65), .dout(n26946));
  jxor g26778(.dina(n26946), .dinb(n26938), .dout(n26947));
  jxor g26779(.dina(n26947), .dinb(n26875), .dout(n26948));
  jand g26780(.dina(n23847), .dinb(n1819), .dout(n26949));
  jand g26781(.dina(n23144), .dinb(n2180), .dout(n26950));
  jand g26782(.dina(n23845), .dinb(n2243), .dout(n26951));
  jor  g26783(.dina(n26951), .dinb(n26950), .dout(n26952));
  jand g26784(.dina(n23079), .dinb(n2185), .dout(n26953));
  jor  g26785(.dina(n26953), .dinb(n26952), .dout(n26954));
  jor  g26786(.dina(n26954), .dinb(n26949), .dout(n26955));
  jxor g26787(.dina(n26955), .dinb(n2196), .dout(n26956));
  jxor g26788(.dina(n26956), .dinb(n26948), .dout(n26957));
  jxor g26789(.dina(n26957), .dinb(n26870), .dout(n26958));
  jnot g26790(.din(n26958), .dout(n26959));
  jor  g26791(.dina(n24516), .dinb(n2744), .dout(n26960));
  jor  g26792(.dina(n24518), .dinb(n2753), .dout(n26961));
  jor  g26793(.dina(n24304), .dinb(n2749), .dout(n26962));
  jor  g26794(.dina(n24266), .dinb(n2758), .dout(n26963));
  jand g26795(.dina(n26963), .dinb(n26962), .dout(n26964));
  jand g26796(.dina(n26964), .dinb(n26961), .dout(n26965));
  jand g26797(.dina(n26965), .dinb(n26960), .dout(n26966));
  jxor g26798(.dina(n26966), .dinb(\a[17] ), .dout(n26967));
  jxor g26799(.dina(n26967), .dinb(n26959), .dout(n26968));
  jxor g26800(.dina(n26968), .dinb(n26864), .dout(n26969));
  jxor g26801(.dina(n26969), .dinb(n26852), .dout(n26970));
  jand g26802(.dina(n26842), .dinb(n26728), .dout(n26971));
  jand g26803(.dina(n26843), .dinb(n26724), .dout(n26972));
  jor  g26804(.dina(n26972), .dinb(n26971), .dout(n26973));
  jxor g26805(.dina(n26973), .dinb(n26970), .dout(n26974));
  jxor g26806(.dina(n26974), .dinb(n26846), .dout(\result[18] ));
  jand g26807(.dina(n26974), .dinb(n26846), .dout(n26976));
  jand g26808(.dina(n26969), .dinb(n26852), .dout(n26977));
  jand g26809(.dina(n26973), .dinb(n26970), .dout(n26978));
  jor  g26810(.dina(n26978), .dinb(n26977), .dout(n26979));
  jor  g26811(.dina(n26863), .dinb(n26857), .dout(n26980));
  jnot g26812(.din(n26980), .dout(n26981));
  jand g26813(.dina(n26968), .dinb(n26864), .dout(n26982));
  jor  g26814(.dina(n26982), .dinb(n26981), .dout(n26983));
  jnot g26815(.din(n26875), .dout(n26984));
  jand g26816(.dina(n26947), .dinb(n26984), .dout(n26985));
  jnot g26817(.din(n26985), .dout(n26986));
  jor  g26818(.dina(n26956), .dinb(n26948), .dout(n26987));
  jand g26819(.dina(n26987), .dinb(n26986), .dout(n26988));
  jnot g26820(.din(n26988), .dout(n26989));
  jor  g26821(.dina(n26925), .dinb(n26917), .dout(n26990));
  jor  g26822(.dina(n26935), .dinb(n26927), .dout(n26991));
  jand g26823(.dina(n26991), .dinb(n26990), .dout(n26992));
  jnot g26824(.din(n26992), .dout(n26993));
  jand g26825(.dina(n26909), .dinb(n26884), .dout(n26994));
  jnot g26826(.din(n26994), .dout(n26995));
  jor  g26827(.dina(n26915), .dinb(n26911), .dout(n26996));
  jand g26828(.dina(n26996), .dinb(n26995), .dout(n26997));
  jnot g26829(.din(n26997), .dout(n26998));
  jor  g26830(.dina(n26907), .dinb(n26778), .dout(n26999));
  jand g26831(.dina(n26908), .dinb(n26891), .dout(n27000));
  jnot g26832(.din(n27000), .dout(n27001));
  jand g26833(.dina(n27001), .dinb(n26999), .dout(n27002));
  jnot g26834(.din(n27002), .dout(n27003));
  jand g26835(.dina(n20115), .dinb(n1407), .dout(n27004));
  jand g26836(.dina(n4420), .dinb(n1917), .dout(n27005));
  jand g26837(.dina(n27005), .dinb(n13302), .dout(n27006));
  jand g26838(.dina(n2106), .dinb(n884), .dout(n27007));
  jand g26839(.dina(n2713), .dinb(n454), .dout(n27008));
  jand g26840(.dina(n27008), .dinb(n27007), .dout(n27009));
  jand g26841(.dina(n27009), .dinb(n15099), .dout(n27010));
  jand g26842(.dina(n27010), .dinb(n7079), .dout(n27011));
  jand g26843(.dina(n27011), .dinb(n829), .dout(n27012));
  jand g26844(.dina(n27012), .dinb(n27006), .dout(n27013));
  jand g26845(.dina(n27013), .dinb(n3861), .dout(n27014));
  jand g26846(.dina(n27014), .dinb(n27004), .dout(n27015));
  jxor g26847(.dina(n27015), .dinb(n26777), .dout(n27016));
  jand g26848(.dina(n25199), .dinb(n20278), .dout(n27017));
  jxor g26849(.dina(n27017), .dinb(n3473), .dout(n27018));
  jxor g26850(.dina(n27018), .dinb(n27016), .dout(n27019));
  jxor g26851(.dina(n27019), .dinb(n27003), .dout(n27020));
  jand g26852(.dina(n21367), .dinb(n5076), .dout(n27021));
  jand g26853(.dina(n21198), .dinb(n5084), .dout(n27022));
  jand g26854(.dina(n20947), .dinb(n5082), .dout(n27023));
  jand g26855(.dina(n20344), .dinb(n6050), .dout(n27024));
  jor  g26856(.dina(n27024), .dinb(n27023), .dout(n27025));
  jor  g26857(.dina(n27025), .dinb(n27022), .dout(n27026));
  jor  g26858(.dina(n27026), .dinb(n27021), .dout(n27027));
  jxor g26859(.dina(n27027), .dinb(n27020), .dout(n27028));
  jnot g26860(.din(n27028), .dout(n27029));
  jand g26861(.dina(n21976), .dinb(n2936), .dout(n27030));
  jand g26862(.dina(n21974), .dinb(n2943), .dout(n27031));
  jand g26863(.dina(n21340), .dinb(n2940), .dout(n27032));
  jand g26864(.dina(n21197), .dinb(n3684), .dout(n27033));
  jor  g26865(.dina(n27033), .dinb(n27032), .dout(n27034));
  jor  g26866(.dina(n27034), .dinb(n27031), .dout(n27035));
  jor  g26867(.dina(n27035), .dinb(n27030), .dout(n27036));
  jxor g26868(.dina(n27036), .dinb(n93), .dout(n27037));
  jxor g26869(.dina(n27037), .dinb(n27029), .dout(n27038));
  jxor g26870(.dina(n27038), .dinb(n26998), .dout(n27039));
  jnot g26871(.din(n27039), .dout(n27040));
  jand g26872(.dina(n22267), .dinb(n71), .dout(n27041));
  jand g26873(.dina(n22265), .dinb(n796), .dout(n27042));
  jand g26874(.dina(n22163), .dinb(n731), .dout(n27043));
  jand g26875(.dina(n22164), .dinb(n1806), .dout(n27044));
  jor  g26876(.dina(n27044), .dinb(n27043), .dout(n27045));
  jor  g26877(.dina(n27045), .dinb(n27042), .dout(n27046));
  jor  g26878(.dina(n27046), .dinb(n27041), .dout(n27047));
  jxor g26879(.dina(n27047), .dinb(n77), .dout(n27048));
  jxor g26880(.dina(n27048), .dinb(n27040), .dout(n27049));
  jxor g26881(.dina(n27049), .dinb(n26993), .dout(n27050));
  jand g26882(.dina(n26936), .dinb(n26880), .dout(n27051));
  jnot g26883(.din(n27051), .dout(n27052));
  jor  g26884(.dina(n26946), .dinb(n26938), .dout(n27053));
  jand g26885(.dina(n27053), .dinb(n27052), .dout(n27054));
  jand g26886(.dina(n23159), .dinb(n806), .dout(n27055));
  jand g26887(.dina(n23079), .dinb(n1620), .dout(n27056));
  jand g26888(.dina(n23080), .dinb(n1612), .dout(n27057));
  jand g26889(.dina(n22937), .dinb(n1644), .dout(n27058));
  jor  g26890(.dina(n27058), .dinb(n27057), .dout(n27059));
  jor  g26891(.dina(n27059), .dinb(n27056), .dout(n27060));
  jor  g26892(.dina(n27060), .dinb(n27055), .dout(n27061));
  jxor g26893(.dina(n27061), .dinb(n65), .dout(n27062));
  jxor g26894(.dina(n27062), .dinb(n27054), .dout(n27063));
  jxor g26895(.dina(n27063), .dinb(n27050), .dout(n27064));
  jnot g26896(.din(n27064), .dout(n27065));
  jand g26897(.dina(n24077), .dinb(n1819), .dout(n27066));
  jand g26898(.dina(n24075), .dinb(n2243), .dout(n27067));
  jand g26899(.dina(n23845), .dinb(n2180), .dout(n27068));
  jand g26900(.dina(n23144), .dinb(n2185), .dout(n27069));
  jor  g26901(.dina(n27069), .dinb(n27068), .dout(n27070));
  jor  g26902(.dina(n27070), .dinb(n27067), .dout(n27071));
  jor  g26903(.dina(n27071), .dinb(n27066), .dout(n27072));
  jxor g26904(.dina(n27072), .dinb(n2196), .dout(n27073));
  jxor g26905(.dina(n27073), .dinb(n27065), .dout(n27074));
  jxor g26906(.dina(n27074), .dinb(n26989), .dout(n27075));
  jand g26907(.dina(n26957), .dinb(n26870), .dout(n27076));
  jnot g26908(.din(n27076), .dout(n27077));
  jor  g26909(.dina(n26967), .dinb(n26959), .dout(n27078));
  jand g26910(.dina(n27078), .dinb(n27077), .dout(n27079));
  jor  g26911(.dina(n24736), .dinb(n2744), .dout(n27080));
  jor  g26912(.dina(n24518), .dinb(n2749), .dout(n27081));
  jor  g26913(.dina(n24738), .dinb(n2753), .dout(n27082));
  jand g26914(.dina(n27082), .dinb(n27081), .dout(n27083));
  jor  g26915(.dina(n24304), .dinb(n2758), .dout(n27084));
  jand g26916(.dina(n27084), .dinb(n27083), .dout(n27085));
  jand g26917(.dina(n27085), .dinb(n27080), .dout(n27086));
  jxor g26918(.dina(n27086), .dinb(\a[17] ), .dout(n27087));
  jxor g26919(.dina(n27087), .dinb(n27079), .dout(n27088));
  jxor g26920(.dina(n27088), .dinb(n27075), .dout(n27089));
  jxor g26921(.dina(n27089), .dinb(n26983), .dout(n27090));
  jxor g26922(.dina(n27090), .dinb(n26979), .dout(n27091));
  jxor g26923(.dina(n27091), .dinb(n26976), .dout(\result[19] ));
  jand g26924(.dina(n27091), .dinb(n26976), .dout(n27093));
  jand g26925(.dina(n27089), .dinb(n26983), .dout(n27094));
  jand g26926(.dina(n27090), .dinb(n26979), .dout(n27095));
  jor  g26927(.dina(n27095), .dinb(n27094), .dout(n27096));
  jor  g26928(.dina(n27087), .dinb(n27079), .dout(n27097));
  jnot g26929(.din(n27097), .dout(n27098));
  jand g26930(.dina(n27088), .dinb(n27075), .dout(n27099));
  jor  g26931(.dina(n27099), .dinb(n27098), .dout(n27100));
  jor  g26932(.dina(n27073), .dinb(n27065), .dout(n27101));
  jand g26933(.dina(n27074), .dinb(n26989), .dout(n27102));
  jnot g26934(.din(n27102), .dout(n27103));
  jand g26935(.dina(n27103), .dinb(n27101), .dout(n27104));
  jor  g26936(.dina(n27062), .dinb(n27054), .dout(n27105));
  jand g26937(.dina(n27063), .dinb(n27050), .dout(n27106));
  jnot g26938(.din(n27106), .dout(n27107));
  jand g26939(.dina(n27107), .dinb(n27105), .dout(n27108));
  jnot g26940(.din(n27108), .dout(n27109));
  jor  g26941(.dina(n27048), .dinb(n27040), .dout(n27110));
  jand g26942(.dina(n27049), .dinb(n26993), .dout(n27111));
  jnot g26943(.din(n27111), .dout(n27112));
  jand g26944(.dina(n27112), .dinb(n27110), .dout(n27113));
  jnot g26945(.din(n27113), .dout(n27114));
  jor  g26946(.dina(n27037), .dinb(n27029), .dout(n27115));
  jand g26947(.dina(n27038), .dinb(n26998), .dout(n27116));
  jnot g26948(.din(n27116), .dout(n27117));
  jand g26949(.dina(n27117), .dinb(n27115), .dout(n27118));
  jnot g26950(.din(n27118), .dout(n27119));
  jand g26951(.dina(n27019), .dinb(n27003), .dout(n27120));
  jand g26952(.dina(n27027), .dinb(n27020), .dout(n27121));
  jor  g26953(.dina(n27121), .dinb(n27120), .dout(n27122));
  jand g26954(.dina(n21355), .dinb(n5076), .dout(n27123));
  jand g26955(.dina(n21197), .dinb(n5084), .dout(n27124));
  jand g26956(.dina(n21198), .dinb(n5082), .dout(n27125));
  jand g26957(.dina(n20947), .dinb(n6050), .dout(n27126));
  jor  g26958(.dina(n27126), .dinb(n27125), .dout(n27127));
  jor  g26959(.dina(n27127), .dinb(n27124), .dout(n27128));
  jor  g26960(.dina(n27128), .dinb(n27123), .dout(n27129));
  jor  g26961(.dina(n27015), .dinb(n26777), .dout(n27130));
  jand g26962(.dina(n27018), .dinb(n27016), .dout(n27131));
  jnot g26963(.din(n27131), .dout(n27132));
  jand g26964(.dina(n27132), .dinb(n27130), .dout(n27133));
  jand g26965(.dina(n5248), .dinb(n622), .dout(n27134));
  jand g26966(.dina(n27134), .dinb(n6307), .dout(n27135));
  jand g26967(.dina(n27135), .dinb(n554), .dout(n27136));
  jand g26968(.dina(n27136), .dinb(n10381), .dout(n27137));
  jand g26969(.dina(n18359), .dinb(n9335), .dout(n27138));
  jand g26970(.dina(n3777), .dinb(n2042), .dout(n27139));
  jand g26971(.dina(n1360), .dinb(n351), .dout(n27140));
  jand g26972(.dina(n27140), .dinb(n1325), .dout(n27141));
  jand g26973(.dina(n27141), .dinb(n27139), .dout(n27142));
  jand g26974(.dina(n21772), .dinb(n514), .dout(n27143));
  jand g26975(.dina(n27143), .dinb(n1043), .dout(n27144));
  jand g26976(.dina(n27144), .dinb(n27142), .dout(n27145));
  jand g26977(.dina(n27145), .dinb(n27138), .dout(n27146));
  jand g26978(.dina(n27146), .dinb(n724), .dout(n27147));
  jand g26979(.dina(n27147), .dinb(n27137), .dout(n27148));
  jnot g26980(.din(n27148), .dout(n27149));
  jxor g26981(.dina(n27149), .dinb(n27133), .dout(n27150));
  jxor g26982(.dina(n27150), .dinb(n27129), .dout(n27151));
  jxor g26983(.dina(n27151), .dinb(n27122), .dout(n27152));
  jnot g26984(.din(n27152), .dout(n27153));
  jand g26985(.dina(n22291), .dinb(n2936), .dout(n27154));
  jand g26986(.dina(n21974), .dinb(n2940), .dout(n27155));
  jand g26987(.dina(n22164), .dinb(n2943), .dout(n27156));
  jor  g26988(.dina(n27156), .dinb(n27155), .dout(n27157));
  jand g26989(.dina(n21340), .dinb(n3684), .dout(n27158));
  jor  g26990(.dina(n27158), .dinb(n27157), .dout(n27159));
  jor  g26991(.dina(n27159), .dinb(n27154), .dout(n27160));
  jxor g26992(.dina(n27160), .dinb(n93), .dout(n27161));
  jxor g26993(.dina(n27161), .dinb(n27153), .dout(n27162));
  jxor g26994(.dina(n27162), .dinb(n27119), .dout(n27163));
  jnot g26995(.din(n27163), .dout(n27164));
  jand g26996(.dina(n22939), .dinb(n71), .dout(n27165));
  jand g26997(.dina(n22937), .dinb(n796), .dout(n27166));
  jand g26998(.dina(n22265), .dinb(n731), .dout(n27167));
  jand g26999(.dina(n22163), .dinb(n1806), .dout(n27168));
  jor  g27000(.dina(n27168), .dinb(n27167), .dout(n27169));
  jor  g27001(.dina(n27169), .dinb(n27166), .dout(n27170));
  jor  g27002(.dina(n27170), .dinb(n27165), .dout(n27171));
  jxor g27003(.dina(n27171), .dinb(n77), .dout(n27172));
  jxor g27004(.dina(n27172), .dinb(n27164), .dout(n27173));
  jxor g27005(.dina(n27173), .dinb(n27114), .dout(n27174));
  jnot g27006(.din(n27174), .dout(n27175));
  jand g27007(.dina(n23146), .dinb(n806), .dout(n27176));
  jand g27008(.dina(n23144), .dinb(n1620), .dout(n27177));
  jand g27009(.dina(n23079), .dinb(n1612), .dout(n27178));
  jand g27010(.dina(n23080), .dinb(n1644), .dout(n27179));
  jor  g27011(.dina(n27179), .dinb(n27178), .dout(n27180));
  jor  g27012(.dina(n27180), .dinb(n27177), .dout(n27181));
  jor  g27013(.dina(n27181), .dinb(n27176), .dout(n27182));
  jxor g27014(.dina(n27182), .dinb(n65), .dout(n27183));
  jxor g27015(.dina(n27183), .dinb(n27175), .dout(n27184));
  jxor g27016(.dina(n27184), .dinb(n27109), .dout(n27185));
  jnot g27017(.din(n27185), .dout(n27186));
  jor  g27018(.dina(n24302), .dinb(n1820), .dout(n27187));
  jor  g27019(.dina(n24266), .dinb(n2181), .dout(n27188));
  jor  g27020(.dina(n24304), .dinb(n2189), .dout(n27189));
  jand g27021(.dina(n27189), .dinb(n27188), .dout(n27190));
  jor  g27022(.dina(n24265), .dinb(n2186), .dout(n27191));
  jand g27023(.dina(n27191), .dinb(n27190), .dout(n27192));
  jand g27024(.dina(n27192), .dinb(n27187), .dout(n27193));
  jxor g27025(.dina(n27193), .dinb(\a[20] ), .dout(n27194));
  jxor g27026(.dina(n27194), .dinb(n27186), .dout(n27195));
  jxor g27027(.dina(n27195), .dinb(n27104), .dout(n27196));
  jor  g27028(.dina(n24932), .dinb(n2744), .dout(n27197));
  jor  g27029(.dina(n24738), .dinb(n2749), .dout(n27198));
  jor  g27030(.dina(n24930), .dinb(n2753), .dout(n27199));
  jand g27031(.dina(n27199), .dinb(n27198), .dout(n27200));
  jor  g27032(.dina(n24518), .dinb(n2758), .dout(n27201));
  jand g27033(.dina(n27201), .dinb(n27200), .dout(n27202));
  jand g27034(.dina(n27202), .dinb(n27197), .dout(n27203));
  jxor g27035(.dina(n27203), .dinb(\a[17] ), .dout(n27204));
  jxor g27036(.dina(n27204), .dinb(n27196), .dout(n27205));
  jxor g27037(.dina(n27205), .dinb(n27100), .dout(n27206));
  jxor g27038(.dina(n27206), .dinb(n27096), .dout(n27207));
  jxor g27039(.dina(n27207), .dinb(n27093), .dout(\result[20] ));
  jand g27040(.dina(n27207), .dinb(n27093), .dout(n27209));
  jnot g27041(.din(n27104), .dout(n27210));
  jand g27042(.dina(n27195), .dinb(n27210), .dout(n27211));
  jor  g27043(.dina(n27204), .dinb(n27196), .dout(n27212));
  jnot g27044(.din(n27212), .dout(n27213));
  jor  g27045(.dina(n27213), .dinb(n27211), .dout(n27214));
  jand g27046(.dina(n27184), .dinb(n27109), .dout(n27215));
  jnot g27047(.din(n27215), .dout(n27216));
  jor  g27048(.dina(n27194), .dinb(n27186), .dout(n27217));
  jand g27049(.dina(n27217), .dinb(n27216), .dout(n27218));
  jor  g27050(.dina(n25116), .dinb(n2744), .dout(n27219));
  jor  g27051(.dina(n24930), .dinb(n20969), .dout(n27220));
  jor  g27052(.dina(n24738), .dinb(n2758), .dout(n27221));
  jand g27053(.dina(n27221), .dinb(n27220), .dout(n27222));
  jand g27054(.dina(n27222), .dinb(n27219), .dout(n27223));
  jxor g27055(.dina(n27223), .dinb(\a[17] ), .dout(n27224));
  jxor g27056(.dina(n27224), .dinb(n27218), .dout(n27225));
  jand g27057(.dina(n27173), .dinb(n27114), .dout(n27226));
  jnot g27058(.din(n27226), .dout(n27227));
  jor  g27059(.dina(n27183), .dinb(n27175), .dout(n27228));
  jand g27060(.dina(n27228), .dinb(n27227), .dout(n27229));
  jnot g27061(.din(n27229), .dout(n27230));
  jand g27062(.dina(n27162), .dinb(n27119), .dout(n27231));
  jnot g27063(.din(n27231), .dout(n27232));
  jor  g27064(.dina(n27172), .dinb(n27164), .dout(n27233));
  jand g27065(.dina(n27233), .dinb(n27232), .dout(n27234));
  jnot g27066(.din(n27234), .dout(n27235));
  jand g27067(.dina(n27151), .dinb(n27122), .dout(n27236));
  jnot g27068(.din(n27236), .dout(n27237));
  jor  g27069(.dina(n27161), .dinb(n27153), .dout(n27238));
  jand g27070(.dina(n27238), .dinb(n27237), .dout(n27239));
  jnot g27071(.din(n27239), .dout(n27240));
  jand g27072(.dina(n21342), .dinb(n5076), .dout(n27241));
  jand g27073(.dina(n21340), .dinb(n5084), .dout(n27242));
  jand g27074(.dina(n21197), .dinb(n5082), .dout(n27243));
  jand g27075(.dina(n21198), .dinb(n6050), .dout(n27244));
  jor  g27076(.dina(n27244), .dinb(n27243), .dout(n27245));
  jor  g27077(.dina(n27245), .dinb(n27242), .dout(n27246));
  jor  g27078(.dina(n27246), .dinb(n27241), .dout(n27247));
  jnot g27079(.din(n27133), .dout(n27248));
  jand g27080(.dina(n27148), .dinb(n27248), .dout(n27249));
  jand g27081(.dina(n27150), .dinb(n27129), .dout(n27250));
  jor  g27082(.dina(n27250), .dinb(n27249), .dout(n27251));
  jand g27083(.dina(n15132), .dinb(n3066), .dout(n27252));
  jand g27084(.dina(n27252), .dinb(n1707), .dout(n27253));
  jand g27085(.dina(n270), .dinb(n901), .dout(n27254));
  jand g27086(.dina(n27254), .dinb(n179), .dout(n27255));
  jand g27087(.dina(n895), .dinb(n824), .dout(n27256));
  jand g27088(.dina(n645), .dinb(n555), .dout(n27257));
  jand g27089(.dina(n27257), .dinb(n27256), .dout(n27258));
  jand g27090(.dina(n27258), .dinb(n27255), .dout(n27259));
  jand g27091(.dina(n27259), .dinb(n1550), .dout(n27260));
  jand g27092(.dina(n27260), .dinb(n27253), .dout(n27261));
  jand g27093(.dina(n6224), .dinb(n1744), .dout(n27262));
  jand g27094(.dina(n27262), .dinb(n1229), .dout(n27263));
  jand g27095(.dina(n27263), .dinb(n27261), .dout(n27264));
  jand g27096(.dina(n27264), .dinb(n9553), .dout(n27265));
  jand g27097(.dina(n21133), .dinb(n14409), .dout(n27266));
  jand g27098(.dina(n27266), .dinb(n4004), .dout(n27267));
  jand g27099(.dina(n27267), .dinb(n27265), .dout(n27268));
  jxor g27100(.dina(n27268), .dinb(n27149), .dout(n27269));
  jxor g27101(.dina(n27269), .dinb(n27251), .dout(n27270));
  jxor g27102(.dina(n27270), .dinb(n27247), .dout(n27271));
  jnot g27103(.din(n27271), .dout(n27272));
  jand g27104(.dina(n22279), .dinb(n2936), .dout(n27273));
  jand g27105(.dina(n22163), .dinb(n2943), .dout(n27274));
  jand g27106(.dina(n22164), .dinb(n2940), .dout(n27275));
  jand g27107(.dina(n21974), .dinb(n3684), .dout(n27276));
  jor  g27108(.dina(n27276), .dinb(n27275), .dout(n27277));
  jor  g27109(.dina(n27277), .dinb(n27274), .dout(n27278));
  jor  g27110(.dina(n27278), .dinb(n27273), .dout(n27279));
  jxor g27111(.dina(n27279), .dinb(n93), .dout(n27280));
  jxor g27112(.dina(n27280), .dinb(n27272), .dout(n27281));
  jxor g27113(.dina(n27281), .dinb(n27240), .dout(n27282));
  jnot g27114(.din(n27282), .dout(n27283));
  jand g27115(.dina(n23172), .dinb(n71), .dout(n27284));
  jand g27116(.dina(n22937), .dinb(n731), .dout(n27285));
  jand g27117(.dina(n23080), .dinb(n796), .dout(n27286));
  jor  g27118(.dina(n27286), .dinb(n27285), .dout(n27287));
  jand g27119(.dina(n22265), .dinb(n1806), .dout(n27288));
  jor  g27120(.dina(n27288), .dinb(n27287), .dout(n27289));
  jor  g27121(.dina(n27289), .dinb(n27284), .dout(n27290));
  jxor g27122(.dina(n27290), .dinb(n77), .dout(n27291));
  jxor g27123(.dina(n27291), .dinb(n27283), .dout(n27292));
  jxor g27124(.dina(n27292), .dinb(n27235), .dout(n27293));
  jnot g27125(.din(n27293), .dout(n27294));
  jand g27126(.dina(n23847), .dinb(n806), .dout(n27295));
  jand g27127(.dina(n23144), .dinb(n1612), .dout(n27296));
  jand g27128(.dina(n23845), .dinb(n1620), .dout(n27297));
  jor  g27129(.dina(n27297), .dinb(n27296), .dout(n27298));
  jand g27130(.dina(n23079), .dinb(n1644), .dout(n27299));
  jor  g27131(.dina(n27299), .dinb(n27298), .dout(n27300));
  jor  g27132(.dina(n27300), .dinb(n27295), .dout(n27301));
  jxor g27133(.dina(n27301), .dinb(n65), .dout(n27302));
  jxor g27134(.dina(n27302), .dinb(n27294), .dout(n27303));
  jxor g27135(.dina(n27303), .dinb(n27230), .dout(n27304));
  jnot g27136(.din(n27304), .dout(n27305));
  jor  g27137(.dina(n24516), .dinb(n1820), .dout(n27306));
  jor  g27138(.dina(n24518), .dinb(n2189), .dout(n27307));
  jor  g27139(.dina(n24304), .dinb(n2181), .dout(n27308));
  jor  g27140(.dina(n24266), .dinb(n2186), .dout(n27309));
  jand g27141(.dina(n27309), .dinb(n27308), .dout(n27310));
  jand g27142(.dina(n27310), .dinb(n27307), .dout(n27311));
  jand g27143(.dina(n27311), .dinb(n27306), .dout(n27312));
  jxor g27144(.dina(n27312), .dinb(\a[20] ), .dout(n27313));
  jxor g27145(.dina(n27313), .dinb(n27305), .dout(n27314));
  jxor g27146(.dina(n27314), .dinb(n27225), .dout(n27315));
  jxor g27147(.dina(n27315), .dinb(n27214), .dout(n27316));
  jand g27148(.dina(n27205), .dinb(n27100), .dout(n27317));
  jand g27149(.dina(n27206), .dinb(n27096), .dout(n27318));
  jor  g27150(.dina(n27318), .dinb(n27317), .dout(n27319));
  jxor g27151(.dina(n27319), .dinb(n27316), .dout(n27320));
  jxor g27152(.dina(n27320), .dinb(n27209), .dout(\result[21] ));
  jand g27153(.dina(n27320), .dinb(n27209), .dout(n27322));
  jand g27154(.dina(n27315), .dinb(n27214), .dout(n27323));
  jand g27155(.dina(n27319), .dinb(n27316), .dout(n27324));
  jor  g27156(.dina(n27324), .dinb(n27323), .dout(n27325));
  jor  g27157(.dina(n27224), .dinb(n27218), .dout(n27326));
  jand g27158(.dina(n27314), .dinb(n27225), .dout(n27327));
  jnot g27159(.din(n27327), .dout(n27328));
  jand g27160(.dina(n27328), .dinb(n27326), .dout(n27329));
  jnot g27161(.din(n27329), .dout(n27330));
  jand g27162(.dina(n27292), .dinb(n27235), .dout(n27331));
  jnot g27163(.din(n27331), .dout(n27332));
  jor  g27164(.dina(n27302), .dinb(n27294), .dout(n27333));
  jand g27165(.dina(n27333), .dinb(n27332), .dout(n27334));
  jnot g27166(.din(n27334), .dout(n27335));
  jand g27167(.dina(n27281), .dinb(n27240), .dout(n27336));
  jnot g27168(.din(n27336), .dout(n27337));
  jor  g27169(.dina(n27291), .dinb(n27283), .dout(n27338));
  jand g27170(.dina(n27338), .dinb(n27337), .dout(n27339));
  jand g27171(.dina(n23159), .dinb(n71), .dout(n27340));
  jand g27172(.dina(n23079), .dinb(n796), .dout(n27341));
  jand g27173(.dina(n23080), .dinb(n731), .dout(n27342));
  jand g27174(.dina(n22937), .dinb(n1806), .dout(n27343));
  jor  g27175(.dina(n27343), .dinb(n27342), .dout(n27344));
  jor  g27176(.dina(n27344), .dinb(n27341), .dout(n27345));
  jor  g27177(.dina(n27345), .dinb(n27340), .dout(n27346));
  jxor g27178(.dina(n27346), .dinb(n77), .dout(n27347));
  jxor g27179(.dina(n27347), .dinb(n27339), .dout(n27348));
  jand g27180(.dina(n27270), .dinb(n27247), .dout(n27349));
  jnot g27181(.din(n27349), .dout(n27350));
  jor  g27182(.dina(n27280), .dinb(n27272), .dout(n27351));
  jand g27183(.dina(n27351), .dinb(n27350), .dout(n27352));
  jnot g27184(.din(n27352), .dout(n27353));
  jand g27185(.dina(n27268), .dinb(n27149), .dout(n27354));
  jand g27186(.dina(n27269), .dinb(n27251), .dout(n27355));
  jor  g27187(.dina(n27355), .dinb(n27354), .dout(n27356));
  jand g27188(.dina(n3879), .dinb(n628), .dout(n27357));
  jand g27189(.dina(n27357), .dinb(n21767), .dout(n27358));
  jand g27190(.dina(n27358), .dinb(n5205), .dout(n27359));
  jand g27191(.dina(n175), .dinb(n1226), .dout(n27360));
  jand g27192(.dina(n27360), .dinb(n5395), .dout(n27361));
  jand g27193(.dina(n1524), .dinb(n555), .dout(n27362));
  jand g27194(.dina(n27362), .dinb(n1575), .dout(n27363));
  jand g27195(.dina(n27363), .dinb(n27361), .dout(n27364));
  jand g27196(.dina(n27364), .dinb(n27359), .dout(n27365));
  jand g27197(.dina(n21252), .dinb(n4587), .dout(n27366));
  jand g27198(.dina(n27366), .dinb(n11406), .dout(n27367));
  jand g27199(.dina(n27367), .dinb(n12616), .dout(n27368));
  jand g27200(.dina(n27368), .dinb(n27365), .dout(n27369));
  jxor g27201(.dina(n27369), .dinb(n27268), .dout(n27370));
  jor  g27202(.dina(n24930), .dinb(n21142), .dout(n27371));
  jxor g27203(.dina(n27371), .dinb(\a[17] ), .dout(n27372));
  jxor g27204(.dina(n27372), .dinb(n27370), .dout(n27373));
  jand g27205(.dina(n21976), .dinb(n5076), .dout(n27374));
  jand g27206(.dina(n21974), .dinb(n5084), .dout(n27375));
  jand g27207(.dina(n21340), .dinb(n5082), .dout(n27376));
  jand g27208(.dina(n21197), .dinb(n6050), .dout(n27377));
  jor  g27209(.dina(n27377), .dinb(n27376), .dout(n27378));
  jor  g27210(.dina(n27378), .dinb(n27375), .dout(n27379));
  jor  g27211(.dina(n27379), .dinb(n27374), .dout(n27380));
  jxor g27212(.dina(n27380), .dinb(n27373), .dout(n27381));
  jxor g27213(.dina(n27381), .dinb(n27356), .dout(n27382));
  jxor g27214(.dina(n27382), .dinb(n27353), .dout(n27383));
  jnot g27215(.din(n27383), .dout(n27384));
  jand g27216(.dina(n22267), .dinb(n2936), .dout(n27385));
  jand g27217(.dina(n22163), .dinb(n2940), .dout(n27386));
  jand g27218(.dina(n22265), .dinb(n2943), .dout(n27387));
  jor  g27219(.dina(n27387), .dinb(n27386), .dout(n27388));
  jand g27220(.dina(n22164), .dinb(n3684), .dout(n27389));
  jor  g27221(.dina(n27389), .dinb(n27388), .dout(n27390));
  jor  g27222(.dina(n27390), .dinb(n27385), .dout(n27391));
  jxor g27223(.dina(n27391), .dinb(n93), .dout(n27392));
  jxor g27224(.dina(n27392), .dinb(n27384), .dout(n27393));
  jxor g27225(.dina(n27393), .dinb(n27348), .dout(n27394));
  jnot g27226(.din(n27394), .dout(n27395));
  jand g27227(.dina(n24077), .dinb(n806), .dout(n27396));
  jand g27228(.dina(n23845), .dinb(n1612), .dout(n27397));
  jand g27229(.dina(n24075), .dinb(n1620), .dout(n27398));
  jor  g27230(.dina(n27398), .dinb(n27397), .dout(n27399));
  jand g27231(.dina(n23144), .dinb(n1644), .dout(n27400));
  jor  g27232(.dina(n27400), .dinb(n27399), .dout(n27401));
  jor  g27233(.dina(n27401), .dinb(n27396), .dout(n27402));
  jxor g27234(.dina(n27402), .dinb(n65), .dout(n27403));
  jxor g27235(.dina(n27403), .dinb(n27395), .dout(n27404));
  jxor g27236(.dina(n27404), .dinb(n27335), .dout(n27405));
  jand g27237(.dina(n27303), .dinb(n27230), .dout(n27406));
  jnot g27238(.din(n27406), .dout(n27407));
  jor  g27239(.dina(n27313), .dinb(n27305), .dout(n27408));
  jand g27240(.dina(n27408), .dinb(n27407), .dout(n27409));
  jor  g27241(.dina(n24736), .dinb(n1820), .dout(n27410));
  jor  g27242(.dina(n24738), .dinb(n2189), .dout(n27411));
  jor  g27243(.dina(n24518), .dinb(n2181), .dout(n27412));
  jor  g27244(.dina(n24304), .dinb(n2186), .dout(n27413));
  jand g27245(.dina(n27413), .dinb(n27412), .dout(n27414));
  jand g27246(.dina(n27414), .dinb(n27411), .dout(n27415));
  jand g27247(.dina(n27415), .dinb(n27410), .dout(n27416));
  jxor g27248(.dina(n27416), .dinb(\a[20] ), .dout(n27417));
  jxor g27249(.dina(n27417), .dinb(n27409), .dout(n27418));
  jxor g27250(.dina(n27418), .dinb(n27405), .dout(n27419));
  jxor g27251(.dina(n27419), .dinb(n27330), .dout(n27420));
  jxor g27252(.dina(n27420), .dinb(n27325), .dout(n27421));
  jxor g27253(.dina(n27421), .dinb(n27322), .dout(\result[22] ));
  jand g27254(.dina(n27421), .dinb(n27322), .dout(n27423));
  jand g27255(.dina(n27419), .dinb(n27330), .dout(n27424));
  jand g27256(.dina(n27420), .dinb(n27325), .dout(n27425));
  jor  g27257(.dina(n27425), .dinb(n27424), .dout(n27426));
  jor  g27258(.dina(n27417), .dinb(n27409), .dout(n27427));
  jand g27259(.dina(n27418), .dinb(n27405), .dout(n27428));
  jnot g27260(.din(n27428), .dout(n27429));
  jand g27261(.dina(n27429), .dinb(n27427), .dout(n27430));
  jnot g27262(.din(n27430), .dout(n27431));
  jor  g27263(.dina(n27403), .dinb(n27395), .dout(n27432));
  jand g27264(.dina(n27404), .dinb(n27335), .dout(n27433));
  jnot g27265(.din(n27433), .dout(n27434));
  jand g27266(.dina(n27434), .dinb(n27432), .dout(n27435));
  jnot g27267(.din(n27435), .dout(n27436));
  jor  g27268(.dina(n27347), .dinb(n27339), .dout(n27437));
  jand g27269(.dina(n27393), .dinb(n27348), .dout(n27438));
  jnot g27270(.din(n27438), .dout(n27439));
  jand g27271(.dina(n27439), .dinb(n27437), .dout(n27440));
  jnot g27272(.din(n27440), .dout(n27441));
  jand g27273(.dina(n27382), .dinb(n27353), .dout(n27442));
  jnot g27274(.din(n27442), .dout(n27443));
  jor  g27275(.dina(n27392), .dinb(n27384), .dout(n27444));
  jand g27276(.dina(n27444), .dinb(n27443), .dout(n27445));
  jnot g27277(.din(n27445), .dout(n27446));
  jand g27278(.dina(n27380), .dinb(n27373), .dout(n27447));
  jand g27279(.dina(n27381), .dinb(n27356), .dout(n27448));
  jor  g27280(.dina(n27448), .dinb(n27447), .dout(n27449));
  jand g27281(.dina(n22291), .dinb(n5076), .dout(n27450));
  jand g27282(.dina(n22164), .dinb(n5084), .dout(n27451));
  jand g27283(.dina(n21974), .dinb(n5082), .dout(n27452));
  jand g27284(.dina(n21340), .dinb(n6050), .dout(n27453));
  jor  g27285(.dina(n27453), .dinb(n27452), .dout(n27454));
  jor  g27286(.dina(n27454), .dinb(n27451), .dout(n27455));
  jor  g27287(.dina(n27455), .dinb(n27450), .dout(n27456));
  jor  g27288(.dina(n27369), .dinb(n27268), .dout(n27457));
  jand g27289(.dina(n27372), .dinb(n27370), .dout(n27458));
  jnot g27290(.din(n27458), .dout(n27459));
  jand g27291(.dina(n27459), .dinb(n27457), .dout(n27460));
  jand g27292(.dina(n11394), .dinb(n2152), .dout(n27461));
  jand g27293(.dina(n27461), .dinb(n16554), .dout(n27462));
  jand g27294(.dina(n1409), .dinb(n1308), .dout(n27463));
  jand g27295(.dina(n27463), .dinb(n27462), .dout(n27464));
  jand g27296(.dina(n27464), .dinb(n26057), .dout(n27465));
  jand g27297(.dina(n630), .dinb(n271), .dout(n27466));
  jand g27298(.dina(n27466), .dinb(n1216), .dout(n27467));
  jand g27299(.dina(n1036), .dinb(n328), .dout(n27468));
  jand g27300(.dina(n27468), .dinb(n1531), .dout(n27469));
  jand g27301(.dina(n27469), .dinb(n641), .dout(n27470));
  jand g27302(.dina(n27470), .dinb(n5453), .dout(n27471));
  jand g27303(.dina(n27471), .dinb(n27467), .dout(n27472));
  jand g27304(.dina(n27472), .dinb(n8377), .dout(n27473));
  jand g27305(.dina(n27473), .dinb(n27465), .dout(n27474));
  jnot g27306(.din(n27474), .dout(n27475));
  jxor g27307(.dina(n27475), .dinb(n27460), .dout(n27476));
  jxor g27308(.dina(n27476), .dinb(n27456), .dout(n27477));
  jxor g27309(.dina(n27477), .dinb(n27449), .dout(n27478));
  jnot g27310(.din(n27478), .dout(n27479));
  jand g27311(.dina(n22939), .dinb(n2936), .dout(n27480));
  jand g27312(.dina(n22265), .dinb(n2940), .dout(n27481));
  jand g27313(.dina(n22937), .dinb(n2943), .dout(n27482));
  jor  g27314(.dina(n27482), .dinb(n27481), .dout(n27483));
  jand g27315(.dina(n22163), .dinb(n3684), .dout(n27484));
  jor  g27316(.dina(n27484), .dinb(n27483), .dout(n27485));
  jor  g27317(.dina(n27485), .dinb(n27480), .dout(n27486));
  jxor g27318(.dina(n27486), .dinb(n93), .dout(n27487));
  jxor g27319(.dina(n27487), .dinb(n27479), .dout(n27488));
  jxor g27320(.dina(n27488), .dinb(n27446), .dout(n27489));
  jnot g27321(.din(n27489), .dout(n27490));
  jand g27322(.dina(n23146), .dinb(n71), .dout(n27491));
  jand g27323(.dina(n23144), .dinb(n796), .dout(n27492));
  jand g27324(.dina(n23079), .dinb(n731), .dout(n27493));
  jand g27325(.dina(n23080), .dinb(n1806), .dout(n27494));
  jor  g27326(.dina(n27494), .dinb(n27493), .dout(n27495));
  jor  g27327(.dina(n27495), .dinb(n27492), .dout(n27496));
  jor  g27328(.dina(n27496), .dinb(n27491), .dout(n27497));
  jxor g27329(.dina(n27497), .dinb(n77), .dout(n27498));
  jxor g27330(.dina(n27498), .dinb(n27490), .dout(n27499));
  jxor g27331(.dina(n27499), .dinb(n27441), .dout(n27500));
  jnot g27332(.din(n27500), .dout(n27501));
  jor  g27333(.dina(n24302), .dinb(n807), .dout(n27502));
  jor  g27334(.dina(n24304), .dinb(n1621), .dout(n27503));
  jor  g27335(.dina(n24266), .dinb(n1613), .dout(n27504));
  jor  g27336(.dina(n24265), .dinb(n1617), .dout(n27505));
  jand g27337(.dina(n27505), .dinb(n27504), .dout(n27506));
  jand g27338(.dina(n27506), .dinb(n27503), .dout(n27507));
  jand g27339(.dina(n27507), .dinb(n27502), .dout(n27508));
  jxor g27340(.dina(n27508), .dinb(\a[23] ), .dout(n27509));
  jxor g27341(.dina(n27509), .dinb(n27501), .dout(n27510));
  jxor g27342(.dina(n27510), .dinb(n27436), .dout(n27511));
  jnot g27343(.din(n27511), .dout(n27512));
  jor  g27344(.dina(n24932), .dinb(n1820), .dout(n27513));
  jor  g27345(.dina(n24930), .dinb(n2189), .dout(n27514));
  jor  g27346(.dina(n24738), .dinb(n2181), .dout(n27515));
  jor  g27347(.dina(n24518), .dinb(n2186), .dout(n27516));
  jand g27348(.dina(n27516), .dinb(n27515), .dout(n27517));
  jand g27349(.dina(n27517), .dinb(n27514), .dout(n27518));
  jand g27350(.dina(n27518), .dinb(n27513), .dout(n27519));
  jxor g27351(.dina(n27519), .dinb(\a[20] ), .dout(n27520));
  jxor g27352(.dina(n27520), .dinb(n27512), .dout(n27521));
  jxor g27353(.dina(n27521), .dinb(n27431), .dout(n27522));
  jxor g27354(.dina(n27522), .dinb(n27426), .dout(n27523));
  jxor g27355(.dina(n27523), .dinb(n27423), .dout(\result[23] ));
  jand g27356(.dina(n27523), .dinb(n27423), .dout(n27525));
  jand g27357(.dina(n27510), .dinb(n27436), .dout(n27526));
  jnot g27358(.din(n27526), .dout(n27527));
  jor  g27359(.dina(n27520), .dinb(n27512), .dout(n27528));
  jand g27360(.dina(n27528), .dinb(n27527), .dout(n27529));
  jnot g27361(.din(n27529), .dout(n27530));
  jand g27362(.dina(n27499), .dinb(n27441), .dout(n27531));
  jnot g27363(.din(n27531), .dout(n27532));
  jor  g27364(.dina(n27509), .dinb(n27501), .dout(n27533));
  jand g27365(.dina(n27533), .dinb(n27532), .dout(n27534));
  jor  g27366(.dina(n25116), .dinb(n1820), .dout(n27535));
  jor  g27367(.dina(n24930), .dinb(n21882), .dout(n27536));
  jor  g27368(.dina(n24738), .dinb(n2186), .dout(n27537));
  jand g27369(.dina(n27537), .dinb(n27536), .dout(n27538));
  jand g27370(.dina(n27538), .dinb(n27535), .dout(n27539));
  jxor g27371(.dina(n27539), .dinb(\a[20] ), .dout(n27540));
  jxor g27372(.dina(n27540), .dinb(n27534), .dout(n27541));
  jand g27373(.dina(n27488), .dinb(n27446), .dout(n27542));
  jnot g27374(.din(n27542), .dout(n27543));
  jor  g27375(.dina(n27498), .dinb(n27490), .dout(n27544));
  jand g27376(.dina(n27544), .dinb(n27543), .dout(n27545));
  jnot g27377(.din(n27545), .dout(n27546));
  jnot g27378(.din(n27460), .dout(n27547));
  jand g27379(.dina(n27474), .dinb(n27547), .dout(n27548));
  jand g27380(.dina(n27476), .dinb(n27456), .dout(n27549));
  jor  g27381(.dina(n27549), .dinb(n27548), .dout(n27550));
  jand g27382(.dina(n22279), .dinb(n5076), .dout(n27551));
  jand g27383(.dina(n22163), .dinb(n5084), .dout(n27552));
  jand g27384(.dina(n22164), .dinb(n5082), .dout(n27553));
  jand g27385(.dina(n21974), .dinb(n6050), .dout(n27554));
  jor  g27386(.dina(n27554), .dinb(n27553), .dout(n27555));
  jor  g27387(.dina(n27555), .dinb(n27552), .dout(n27556));
  jor  g27388(.dina(n27556), .dinb(n27551), .dout(n27557));
  jand g27389(.dina(n673), .dinb(n1160), .dout(n27558));
  jand g27390(.dina(n27558), .dinb(n5228), .dout(n27559));
  jand g27391(.dina(n8141), .dinb(n1212), .dout(n27560));
  jand g27392(.dina(n21238), .dinb(n510), .dout(n27561));
  jand g27393(.dina(n27561), .dinb(n1189), .dout(n27562));
  jand g27394(.dina(n27562), .dinb(n25372), .dout(n27563));
  jand g27395(.dina(n27563), .dinb(n713), .dout(n27564));
  jand g27396(.dina(n27564), .dinb(n27560), .dout(n27565));
  jand g27397(.dina(n27255), .dinb(n12613), .dout(n27566));
  jand g27398(.dina(n27566), .dinb(n11543), .dout(n27567));
  jand g27399(.dina(n27567), .dinb(n5379), .dout(n27568));
  jand g27400(.dina(n27568), .dinb(n27565), .dout(n27569));
  jand g27401(.dina(n27569), .dinb(n27559), .dout(n27570));
  jxor g27402(.dina(n27570), .dinb(n27475), .dout(n27571));
  jxor g27403(.dina(n27571), .dinb(n27557), .dout(n27572));
  jxor g27404(.dina(n27572), .dinb(n27550), .dout(n27573));
  jnot g27405(.din(n27573), .dout(n27574));
  jand g27406(.dina(n27477), .dinb(n27449), .dout(n27575));
  jnot g27407(.din(n27575), .dout(n27576));
  jor  g27408(.dina(n27487), .dinb(n27479), .dout(n27577));
  jand g27409(.dina(n27577), .dinb(n27576), .dout(n27578));
  jxor g27410(.dina(n27578), .dinb(n27574), .dout(n27579));
  jnot g27411(.din(n27579), .dout(n27580));
  jand g27412(.dina(n23172), .dinb(n2936), .dout(n27581));
  jand g27413(.dina(n22937), .dinb(n2940), .dout(n27582));
  jand g27414(.dina(n23080), .dinb(n2943), .dout(n27583));
  jor  g27415(.dina(n27583), .dinb(n27582), .dout(n27584));
  jand g27416(.dina(n22265), .dinb(n3684), .dout(n27585));
  jor  g27417(.dina(n27585), .dinb(n27584), .dout(n27586));
  jor  g27418(.dina(n27586), .dinb(n27581), .dout(n27587));
  jxor g27419(.dina(n27587), .dinb(n93), .dout(n27588));
  jxor g27420(.dina(n27588), .dinb(n27580), .dout(n27589));
  jnot g27421(.din(n27589), .dout(n27590));
  jand g27422(.dina(n23847), .dinb(n71), .dout(n27591));
  jand g27423(.dina(n23144), .dinb(n731), .dout(n27592));
  jand g27424(.dina(n23845), .dinb(n796), .dout(n27593));
  jor  g27425(.dina(n27593), .dinb(n27592), .dout(n27594));
  jand g27426(.dina(n23079), .dinb(n1806), .dout(n27595));
  jor  g27427(.dina(n27595), .dinb(n27594), .dout(n27596));
  jor  g27428(.dina(n27596), .dinb(n27591), .dout(n27597));
  jxor g27429(.dina(n27597), .dinb(n77), .dout(n27598));
  jxor g27430(.dina(n27598), .dinb(n27590), .dout(n27599));
  jxor g27431(.dina(n27599), .dinb(n27546), .dout(n27600));
  jnot g27432(.din(n27600), .dout(n27601));
  jor  g27433(.dina(n24516), .dinb(n807), .dout(n27602));
  jor  g27434(.dina(n24304), .dinb(n1613), .dout(n27603));
  jor  g27435(.dina(n24518), .dinb(n1621), .dout(n27604));
  jand g27436(.dina(n27604), .dinb(n27603), .dout(n27605));
  jor  g27437(.dina(n24266), .dinb(n1617), .dout(n27606));
  jand g27438(.dina(n27606), .dinb(n27605), .dout(n27607));
  jand g27439(.dina(n27607), .dinb(n27602), .dout(n27608));
  jxor g27440(.dina(n27608), .dinb(\a[23] ), .dout(n27609));
  jxor g27441(.dina(n27609), .dinb(n27601), .dout(n27610));
  jxor g27442(.dina(n27610), .dinb(n27541), .dout(n27611));
  jxor g27443(.dina(n27611), .dinb(n27530), .dout(n27612));
  jand g27444(.dina(n27521), .dinb(n27431), .dout(n27613));
  jand g27445(.dina(n27522), .dinb(n27426), .dout(n27614));
  jor  g27446(.dina(n27614), .dinb(n27613), .dout(n27615));
  jxor g27447(.dina(n27615), .dinb(n27612), .dout(n27616));
  jxor g27448(.dina(n27616), .dinb(n27525), .dout(\result[24] ));
  jand g27449(.dina(n27616), .dinb(n27525), .dout(n27618));
  jand g27450(.dina(n27611), .dinb(n27530), .dout(n27619));
  jand g27451(.dina(n27615), .dinb(n27612), .dout(n27620));
  jor  g27452(.dina(n27620), .dinb(n27619), .dout(n27621));
  jor  g27453(.dina(n27540), .dinb(n27534), .dout(n27622));
  jand g27454(.dina(n27610), .dinb(n27541), .dout(n27623));
  jnot g27455(.din(n27623), .dout(n27624));
  jand g27456(.dina(n27624), .dinb(n27622), .dout(n27625));
  jnot g27457(.din(n27625), .dout(n27626));
  jor  g27458(.dina(n27588), .dinb(n27580), .dout(n27627));
  jor  g27459(.dina(n27598), .dinb(n27590), .dout(n27628));
  jand g27460(.dina(n27628), .dinb(n27627), .dout(n27629));
  jnot g27461(.din(n27629), .dout(n27630));
  jand g27462(.dina(n27572), .dinb(n27550), .dout(n27631));
  jnot g27463(.din(n27631), .dout(n27632));
  jor  g27464(.dina(n27578), .dinb(n27574), .dout(n27633));
  jand g27465(.dina(n27633), .dinb(n27632), .dout(n27634));
  jnot g27466(.din(n27634), .dout(n27635));
  jor  g27467(.dina(n27570), .dinb(n27475), .dout(n27636));
  jand g27468(.dina(n27571), .dinb(n27557), .dout(n27637));
  jnot g27469(.din(n27637), .dout(n27638));
  jand g27470(.dina(n27638), .dinb(n27636), .dout(n27639));
  jnot g27471(.din(n27639), .dout(n27640));
  jand g27472(.dina(n15654), .dinb(n6379), .dout(n27641));
  jand g27473(.dina(n1237), .dinb(n964), .dout(n27642));
  jand g27474(.dina(n27642), .dinb(n978), .dout(n27643));
  jand g27475(.dina(n7503), .dinb(n621), .dout(n27644));
  jand g27476(.dina(n27644), .dinb(n27643), .dout(n27645));
  jand g27477(.dina(n27645), .dinb(n1550), .dout(n27646));
  jand g27478(.dina(n27646), .dinb(n2522), .dout(n27647));
  jand g27479(.dina(n27647), .dinb(n27641), .dout(n27648));
  jand g27480(.dina(n27648), .dinb(n4447), .dout(n27649));
  jand g27481(.dina(n4528), .dinb(n137), .dout(n27650));
  jand g27482(.dina(n4668), .dinb(n325), .dout(n27651));
  jand g27483(.dina(n27651), .dinb(n17805), .dout(n27652));
  jand g27484(.dina(n5171), .dinb(n884), .dout(n27653));
  jand g27485(.dina(n27653), .dinb(n27652), .dout(n27654));
  jand g27486(.dina(n27654), .dinb(n27650), .dout(n27655));
  jand g27487(.dina(n27655), .dinb(n11215), .dout(n27656));
  jand g27488(.dina(n27656), .dinb(n27649), .dout(n27657));
  jxor g27489(.dina(n27657), .dinb(n27474), .dout(n27658));
  jor  g27490(.dina(n24930), .dinb(n22044), .dout(n27659));
  jxor g27491(.dina(n27659), .dinb(\a[20] ), .dout(n27660));
  jxor g27492(.dina(n27660), .dinb(n27658), .dout(n27661));
  jxor g27493(.dina(n27661), .dinb(n27640), .dout(n27662));
  jand g27494(.dina(n22267), .dinb(n5076), .dout(n27663));
  jand g27495(.dina(n22265), .dinb(n5084), .dout(n27664));
  jand g27496(.dina(n22163), .dinb(n5082), .dout(n27665));
  jand g27497(.dina(n22164), .dinb(n6050), .dout(n27666));
  jor  g27498(.dina(n27666), .dinb(n27665), .dout(n27667));
  jor  g27499(.dina(n27667), .dinb(n27664), .dout(n27668));
  jor  g27500(.dina(n27668), .dinb(n27663), .dout(n27669));
  jxor g27501(.dina(n27669), .dinb(n27662), .dout(n27670));
  jxor g27502(.dina(n27670), .dinb(n27635), .dout(n27671));
  jnot g27503(.din(n27671), .dout(n27672));
  jand g27504(.dina(n23159), .dinb(n2936), .dout(n27673));
  jand g27505(.dina(n23080), .dinb(n2940), .dout(n27674));
  jand g27506(.dina(n23079), .dinb(n2943), .dout(n27675));
  jor  g27507(.dina(n27675), .dinb(n27674), .dout(n27676));
  jand g27508(.dina(n22937), .dinb(n3684), .dout(n27677));
  jor  g27509(.dina(n27677), .dinb(n27676), .dout(n27678));
  jor  g27510(.dina(n27678), .dinb(n27673), .dout(n27679));
  jxor g27511(.dina(n27679), .dinb(n93), .dout(n27680));
  jxor g27512(.dina(n27680), .dinb(n27672), .dout(n27681));
  jnot g27513(.din(n27681), .dout(n27682));
  jand g27514(.dina(n24077), .dinb(n71), .dout(n27683));
  jand g27515(.dina(n24075), .dinb(n796), .dout(n27684));
  jand g27516(.dina(n23845), .dinb(n731), .dout(n27685));
  jand g27517(.dina(n23144), .dinb(n1806), .dout(n27686));
  jor  g27518(.dina(n27686), .dinb(n27685), .dout(n27687));
  jor  g27519(.dina(n27687), .dinb(n27684), .dout(n27688));
  jor  g27520(.dina(n27688), .dinb(n27683), .dout(n27689));
  jxor g27521(.dina(n27689), .dinb(n77), .dout(n27690));
  jxor g27522(.dina(n27690), .dinb(n27682), .dout(n27691));
  jxor g27523(.dina(n27691), .dinb(n27630), .dout(n27692));
  jand g27524(.dina(n27599), .dinb(n27546), .dout(n27693));
  jnot g27525(.din(n27693), .dout(n27694));
  jor  g27526(.dina(n27609), .dinb(n27601), .dout(n27695));
  jand g27527(.dina(n27695), .dinb(n27694), .dout(n27696));
  jor  g27528(.dina(n24736), .dinb(n807), .dout(n27697));
  jor  g27529(.dina(n24738), .dinb(n1621), .dout(n27698));
  jor  g27530(.dina(n24304), .dinb(n1617), .dout(n27699));
  jor  g27531(.dina(n24518), .dinb(n1613), .dout(n27700));
  jand g27532(.dina(n27700), .dinb(n27699), .dout(n27701));
  jand g27533(.dina(n27701), .dinb(n27698), .dout(n27702));
  jand g27534(.dina(n27702), .dinb(n27697), .dout(n27703));
  jxor g27535(.dina(n27703), .dinb(\a[23] ), .dout(n27704));
  jxor g27536(.dina(n27704), .dinb(n27696), .dout(n27705));
  jxor g27537(.dina(n27705), .dinb(n27692), .dout(n27706));
  jxor g27538(.dina(n27706), .dinb(n27626), .dout(n27707));
  jxor g27539(.dina(n27707), .dinb(n27621), .dout(n27708));
  jxor g27540(.dina(n27708), .dinb(n27618), .dout(\result[25] ));
  jand g27541(.dina(n27708), .dinb(n27618), .dout(n27710));
  jand g27542(.dina(n27706), .dinb(n27626), .dout(n27711));
  jand g27543(.dina(n27707), .dinb(n27621), .dout(n27712));
  jor  g27544(.dina(n27712), .dinb(n27711), .dout(n27713));
  jor  g27545(.dina(n27704), .dinb(n27696), .dout(n27714));
  jand g27546(.dina(n27705), .dinb(n27692), .dout(n27715));
  jnot g27547(.din(n27715), .dout(n27716));
  jand g27548(.dina(n27716), .dinb(n27714), .dout(n27717));
  jnot g27549(.din(n27717), .dout(n27718));
  jor  g27550(.dina(n27690), .dinb(n27682), .dout(n27719));
  jand g27551(.dina(n27691), .dinb(n27630), .dout(n27720));
  jnot g27552(.din(n27720), .dout(n27721));
  jand g27553(.dina(n27721), .dinb(n27719), .dout(n27722));
  jnot g27554(.din(n27722), .dout(n27723));
  jand g27555(.dina(n27670), .dinb(n27635), .dout(n27724));
  jnot g27556(.din(n27724), .dout(n27725));
  jor  g27557(.dina(n27680), .dinb(n27672), .dout(n27726));
  jand g27558(.dina(n27726), .dinb(n27725), .dout(n27727));
  jnot g27559(.din(n27727), .dout(n27728));
  jand g27560(.dina(n27661), .dinb(n27640), .dout(n27729));
  jand g27561(.dina(n27669), .dinb(n27662), .dout(n27730));
  jor  g27562(.dina(n27730), .dinb(n27729), .dout(n27731));
  jand g27563(.dina(n22939), .dinb(n5076), .dout(n27732));
  jand g27564(.dina(n22937), .dinb(n5084), .dout(n27733));
  jand g27565(.dina(n22265), .dinb(n5082), .dout(n27734));
  jand g27566(.dina(n22163), .dinb(n6050), .dout(n27735));
  jor  g27567(.dina(n27735), .dinb(n27734), .dout(n27736));
  jor  g27568(.dina(n27736), .dinb(n27733), .dout(n27737));
  jor  g27569(.dina(n27737), .dinb(n27732), .dout(n27738));
  jor  g27570(.dina(n27657), .dinb(n27474), .dout(n27739));
  jand g27571(.dina(n27660), .dinb(n27658), .dout(n27740));
  jnot g27572(.din(n27740), .dout(n27741));
  jand g27573(.dina(n27741), .dinb(n27739), .dout(n27742));
  jand g27574(.dina(n2701), .dinb(n2052), .dout(n27743));
  jand g27575(.dina(n1577), .dinb(n469), .dout(n27744));
  jand g27576(.dina(n27744), .dinb(n8362), .dout(n27745));
  jand g27577(.dina(n27745), .dinb(n1212), .dout(n27746));
  jand g27578(.dina(n27746), .dinb(n27743), .dout(n27747));
  jand g27579(.dina(n3214), .dinb(n1260), .dout(n27748));
  jand g27580(.dina(n27748), .dinb(n3179), .dout(n27749));
  jand g27581(.dina(n27749), .dinb(n670), .dout(n27750));
  jand g27582(.dina(n27750), .dinb(n27747), .dout(n27751));
  jand g27583(.dina(n27751), .dinb(n3106), .dout(n27752));
  jand g27584(.dina(n18385), .dinb(n14056), .dout(n27753));
  jand g27585(.dina(n13312), .dinb(n3274), .dout(n27754));
  jand g27586(.dina(n27754), .dinb(n27753), .dout(n27755));
  jand g27587(.dina(n27755), .dinb(n12616), .dout(n27756));
  jand g27588(.dina(n27756), .dinb(n27752), .dout(n27757));
  jnot g27589(.din(n27757), .dout(n27758));
  jxor g27590(.dina(n27758), .dinb(n27742), .dout(n27759));
  jxor g27591(.dina(n27759), .dinb(n27738), .dout(n27760));
  jxor g27592(.dina(n27760), .dinb(n27731), .dout(n27761));
  jnot g27593(.din(n27761), .dout(n27762));
  jand g27594(.dina(n23146), .dinb(n2936), .dout(n27763));
  jand g27595(.dina(n23079), .dinb(n2940), .dout(n27764));
  jand g27596(.dina(n23144), .dinb(n2943), .dout(n27765));
  jor  g27597(.dina(n27765), .dinb(n27764), .dout(n27766));
  jand g27598(.dina(n23080), .dinb(n3684), .dout(n27767));
  jor  g27599(.dina(n27767), .dinb(n27766), .dout(n27768));
  jor  g27600(.dina(n27768), .dinb(n27763), .dout(n27769));
  jxor g27601(.dina(n27769), .dinb(n93), .dout(n27770));
  jxor g27602(.dina(n27770), .dinb(n27762), .dout(n27771));
  jxor g27603(.dina(n27771), .dinb(n27728), .dout(n27772));
  jnot g27604(.din(n27772), .dout(n27773));
  jor  g27605(.dina(n24302), .dinb(n2303), .dout(n27774));
  jor  g27606(.dina(n24266), .dinb(n2306), .dout(n27775));
  jor  g27607(.dina(n24304), .dinb(n2309), .dout(n27776));
  jand g27608(.dina(n27776), .dinb(n27775), .dout(n27777));
  jor  g27609(.dina(n24265), .dinb(n1805), .dout(n27778));
  jand g27610(.dina(n27778), .dinb(n27777), .dout(n27779));
  jand g27611(.dina(n27779), .dinb(n27774), .dout(n27780));
  jxor g27612(.dina(n27780), .dinb(\a[26] ), .dout(n27781));
  jxor g27613(.dina(n27781), .dinb(n27773), .dout(n27782));
  jxor g27614(.dina(n27782), .dinb(n27723), .dout(n27783));
  jnot g27615(.din(n27783), .dout(n27784));
  jor  g27616(.dina(n24932), .dinb(n807), .dout(n27785));
  jor  g27617(.dina(n24930), .dinb(n1621), .dout(n27786));
  jor  g27618(.dina(n24738), .dinb(n1613), .dout(n27787));
  jor  g27619(.dina(n24518), .dinb(n1617), .dout(n27788));
  jand g27620(.dina(n27788), .dinb(n27787), .dout(n27789));
  jand g27621(.dina(n27789), .dinb(n27786), .dout(n27790));
  jand g27622(.dina(n27790), .dinb(n27785), .dout(n27791));
  jxor g27623(.dina(n27791), .dinb(\a[23] ), .dout(n27792));
  jxor g27624(.dina(n27792), .dinb(n27784), .dout(n27793));
  jxor g27625(.dina(n27793), .dinb(n27718), .dout(n27794));
  jxor g27626(.dina(n27794), .dinb(n27713), .dout(n27795));
  jxor g27627(.dina(n27795), .dinb(n27710), .dout(\result[26] ));
  jand g27628(.dina(n27795), .dinb(n27710), .dout(n27797));
  jnot g27629(.din(n27797), .dout(n27798));
  jand g27630(.dina(n27782), .dinb(n27723), .dout(n27799));
  jnot g27631(.din(n27799), .dout(n27800));
  jor  g27632(.dina(n27792), .dinb(n27784), .dout(n27801));
  jand g27633(.dina(n27801), .dinb(n27800), .dout(n27802));
  jnot g27634(.din(n27802), .dout(n27803));
  jand g27635(.dina(n27771), .dinb(n27728), .dout(n27804));
  jnot g27636(.din(n27804), .dout(n27805));
  jor  g27637(.dina(n27781), .dinb(n27773), .dout(n27806));
  jand g27638(.dina(n27806), .dinb(n27805), .dout(n27807));
  jor  g27639(.dina(n25116), .dinb(n807), .dout(n27808));
  jor  g27640(.dina(n24738), .dinb(n1617), .dout(n27809));
  jor  g27641(.dina(n24930), .dinb(n22185), .dout(n27810));
  jand g27642(.dina(n27810), .dinb(n27809), .dout(n27811));
  jand g27643(.dina(n27811), .dinb(n27808), .dout(n27812));
  jxor g27644(.dina(n27812), .dinb(\a[23] ), .dout(n27813));
  jxor g27645(.dina(n27813), .dinb(n27807), .dout(n27814));
  jand g27646(.dina(n27760), .dinb(n27731), .dout(n27815));
  jnot g27647(.din(n27815), .dout(n27816));
  jor  g27648(.dina(n27770), .dinb(n27762), .dout(n27817));
  jand g27649(.dina(n27817), .dinb(n27816), .dout(n27818));
  jnot g27650(.din(n27818), .dout(n27819));
  jand g27651(.dina(n23172), .dinb(n5076), .dout(n27820));
  jand g27652(.dina(n23080), .dinb(n5084), .dout(n27821));
  jand g27653(.dina(n22937), .dinb(n5082), .dout(n27822));
  jand g27654(.dina(n22265), .dinb(n6050), .dout(n27823));
  jor  g27655(.dina(n27823), .dinb(n27822), .dout(n27824));
  jor  g27656(.dina(n27824), .dinb(n27821), .dout(n27825));
  jor  g27657(.dina(n27825), .dinb(n27820), .dout(n27826));
  jnot g27658(.din(n27742), .dout(n27827));
  jand g27659(.dina(n27757), .dinb(n27827), .dout(n27828));
  jand g27660(.dina(n27759), .dinb(n27738), .dout(n27829));
  jor  g27661(.dina(n27829), .dinb(n27828), .dout(n27830));
  jand g27662(.dina(n808), .dinb(n907), .dout(n27831));
  jand g27663(.dina(n27831), .dinb(n5501), .dout(n27832));
  jand g27664(.dina(n27832), .dinb(n3827), .dout(n27833));
  jand g27665(.dina(n2052), .dinb(n1160), .dout(n27834));
  jand g27666(.dina(n27834), .dinb(n16565), .dout(n27835));
  jand g27667(.dina(n27835), .dinb(n27833), .dout(n27836));
  jand g27668(.dina(n16182), .dinb(n1247), .dout(n27837));
  jand g27669(.dina(n3989), .dinb(n1238), .dout(n27838));
  jand g27670(.dina(n27838), .dinb(n950), .dout(n27839));
  jand g27671(.dina(n27839), .dinb(n27837), .dout(n27840));
  jand g27672(.dina(n27840), .dinb(n27836), .dout(n27841));
  jand g27673(.dina(n27841), .dinb(n22972), .dout(n27842));
  jand g27674(.dina(n27842), .dinb(n11705), .dout(n27843));
  jand g27675(.dina(n26072), .dinb(n19697), .dout(n27844));
  jand g27676(.dina(n27844), .dinb(n27843), .dout(n27845));
  jxor g27677(.dina(n27845), .dinb(n27758), .dout(n27846));
  jxor g27678(.dina(n27846), .dinb(n27830), .dout(n27847));
  jxor g27679(.dina(n27847), .dinb(n27826), .dout(n27848));
  jxor g27680(.dina(n27848), .dinb(n27819), .dout(n27849));
  jnot g27681(.din(n27849), .dout(n27850));
  jand g27682(.dina(n23847), .dinb(n2936), .dout(n27851));
  jand g27683(.dina(n23845), .dinb(n2943), .dout(n27852));
  jand g27684(.dina(n23144), .dinb(n2940), .dout(n27853));
  jand g27685(.dina(n23079), .dinb(n3684), .dout(n27854));
  jor  g27686(.dina(n27854), .dinb(n27853), .dout(n27855));
  jor  g27687(.dina(n27855), .dinb(n27852), .dout(n27856));
  jor  g27688(.dina(n27856), .dinb(n27851), .dout(n27857));
  jxor g27689(.dina(n27857), .dinb(n93), .dout(n27858));
  jxor g27690(.dina(n27858), .dinb(n27850), .dout(n27859));
  jnot g27691(.din(n27859), .dout(n27860));
  jor  g27692(.dina(n24516), .dinb(n2303), .dout(n27861));
  jor  g27693(.dina(n24304), .dinb(n2306), .dout(n27862));
  jor  g27694(.dina(n24518), .dinb(n2309), .dout(n27863));
  jand g27695(.dina(n27863), .dinb(n27862), .dout(n27864));
  jor  g27696(.dina(n24266), .dinb(n1805), .dout(n27865));
  jand g27697(.dina(n27865), .dinb(n27864), .dout(n27866));
  jand g27698(.dina(n27866), .dinb(n27861), .dout(n27867));
  jxor g27699(.dina(n27867), .dinb(\a[26] ), .dout(n27868));
  jxor g27700(.dina(n27868), .dinb(n27860), .dout(n27869));
  jxor g27701(.dina(n27869), .dinb(n27814), .dout(n27870));
  jxor g27702(.dina(n27870), .dinb(n27803), .dout(n27871));
  jnot g27703(.din(n27871), .dout(n27872));
  jand g27704(.dina(n27793), .dinb(n27718), .dout(n27873));
  jand g27705(.dina(n27794), .dinb(n27713), .dout(n27874));
  jor  g27706(.dina(n27874), .dinb(n27873), .dout(n27875));
  jxor g27707(.dina(n27875), .dinb(n27872), .dout(n27876));
  jxor g27708(.dina(n27876), .dinb(n27798), .dout(\result[27] ));
  jor  g27709(.dina(n27876), .dinb(n27798), .dout(n27878));
  jnot g27710(.din(n27878), .dout(n27879));
  jand g27711(.dina(n27870), .dinb(n27803), .dout(n27880));
  jand g27712(.dina(n27875), .dinb(n27871), .dout(n27881));
  jor  g27713(.dina(n27881), .dinb(n27880), .dout(n27882));
  jor  g27714(.dina(n27813), .dinb(n27807), .dout(n27883));
  jand g27715(.dina(n27869), .dinb(n27814), .dout(n27884));
  jnot g27716(.din(n27884), .dout(n27885));
  jand g27717(.dina(n27885), .dinb(n27883), .dout(n27886));
  jnot g27718(.din(n27886), .dout(n27887));
  jor  g27719(.dina(n27858), .dinb(n27850), .dout(n27888));
  jor  g27720(.dina(n27868), .dinb(n27860), .dout(n27889));
  jand g27721(.dina(n27889), .dinb(n27888), .dout(n27890));
  jor  g27722(.dina(n24736), .dinb(n2303), .dout(n27891));
  jor  g27723(.dina(n24738), .dinb(n2309), .dout(n27892));
  jor  g27724(.dina(n24518), .dinb(n2306), .dout(n27893));
  jor  g27725(.dina(n24304), .dinb(n1805), .dout(n27894));
  jand g27726(.dina(n27894), .dinb(n27893), .dout(n27895));
  jand g27727(.dina(n27895), .dinb(n27892), .dout(n27896));
  jand g27728(.dina(n27896), .dinb(n27891), .dout(n27897));
  jxor g27729(.dina(n27897), .dinb(\a[26] ), .dout(n27898));
  jxor g27730(.dina(n27898), .dinb(n27890), .dout(n27899));
  jand g27731(.dina(n27847), .dinb(n27826), .dout(n27900));
  jand g27732(.dina(n27848), .dinb(n27819), .dout(n27901));
  jor  g27733(.dina(n27901), .dinb(n27900), .dout(n27902));
  jand g27734(.dina(n27845), .dinb(n27758), .dout(n27903));
  jand g27735(.dina(n27846), .dinb(n27830), .dout(n27904));
  jor  g27736(.dina(n27904), .dinb(n27903), .dout(n27905));
  jand g27737(.dina(n7231), .dinb(n1732), .dout(n27906));
  jand g27738(.dina(n27906), .dinb(n3392), .dout(n27907));
  jand g27739(.dina(n27907), .dinb(n8127), .dout(n27908));
  jand g27740(.dina(n27908), .dinb(n7656), .dout(n27909));
  jand g27741(.dina(n27909), .dinb(n7251), .dout(n27910));
  jand g27742(.dina(n925), .dinb(n871), .dout(n27911));
  jand g27743(.dina(n1473), .dinb(n870), .dout(n27912));
  jand g27744(.dina(n27912), .dinb(n27911), .dout(n27913));
  jand g27745(.dina(n27913), .dinb(n11367), .dout(n27914));
  jand g27746(.dina(n27914), .dinb(n563), .dout(n27915));
  jand g27747(.dina(n27915), .dinb(n27910), .dout(n27916));
  jand g27748(.dina(n27916), .dinb(n15532), .dout(n27917));
  jxor g27749(.dina(n27917), .dinb(n27845), .dout(n27918));
  jand g27750(.dina(n25199), .dinb(n22910), .dout(n27919));
  jxor g27751(.dina(n27919), .dinb(n65), .dout(n27920));
  jxor g27752(.dina(n27920), .dinb(n27918), .dout(n27921));
  jxor g27753(.dina(n27921), .dinb(n27905), .dout(n27922));
  jand g27754(.dina(n23159), .dinb(n5076), .dout(n27923));
  jand g27755(.dina(n23079), .dinb(n5084), .dout(n27924));
  jand g27756(.dina(n23080), .dinb(n5082), .dout(n27925));
  jand g27757(.dina(n22937), .dinb(n6050), .dout(n27926));
  jor  g27758(.dina(n27926), .dinb(n27925), .dout(n27927));
  jor  g27759(.dina(n27927), .dinb(n27924), .dout(n27928));
  jor  g27760(.dina(n27928), .dinb(n27923), .dout(n27929));
  jxor g27761(.dina(n27929), .dinb(n27922), .dout(n27930));
  jxor g27762(.dina(n27930), .dinb(n27902), .dout(n27931));
  jand g27763(.dina(n24077), .dinb(n2936), .dout(n27932));
  jand g27764(.dina(n24075), .dinb(n2943), .dout(n27933));
  jand g27765(.dina(n23845), .dinb(n2940), .dout(n27934));
  jand g27766(.dina(n23144), .dinb(n3684), .dout(n27935));
  jor  g27767(.dina(n27935), .dinb(n27934), .dout(n27936));
  jor  g27768(.dina(n27936), .dinb(n27933), .dout(n27937));
  jor  g27769(.dina(n27937), .dinb(n27932), .dout(n27938));
  jxor g27770(.dina(n27938), .dinb(n93), .dout(n27939));
  jnot g27771(.din(n27939), .dout(n27940));
  jxor g27772(.dina(n27940), .dinb(n27931), .dout(n27941));
  jxor g27773(.dina(n27941), .dinb(n27899), .dout(n27942));
  jxor g27774(.dina(n27942), .dinb(n27887), .dout(n27943));
  jxor g27775(.dina(n27943), .dinb(n27882), .dout(n27944));
  jxor g27776(.dina(n27944), .dinb(n27879), .dout(\result[28] ));
  jand g27777(.dina(n27944), .dinb(n27879), .dout(n27946));
  jand g27778(.dina(n27942), .dinb(n27887), .dout(n27947));
  jand g27779(.dina(n27943), .dinb(n27882), .dout(n27948));
  jor  g27780(.dina(n27948), .dinb(n27947), .dout(n27949));
  jor  g27781(.dina(n27898), .dinb(n27890), .dout(n27950));
  jand g27782(.dina(n27941), .dinb(n27899), .dout(n27951));
  jnot g27783(.din(n27951), .dout(n27952));
  jand g27784(.dina(n27952), .dinb(n27950), .dout(n27953));
  jnot g27785(.din(n27953), .dout(n27954));
  jand g27786(.dina(n27930), .dinb(n27902), .dout(n27955));
  jand g27787(.dina(n27940), .dinb(n27931), .dout(n27956));
  jor  g27788(.dina(n27956), .dinb(n27955), .dout(n27957));
  jand g27789(.dina(n27921), .dinb(n27905), .dout(n27958));
  jand g27790(.dina(n27929), .dinb(n27922), .dout(n27959));
  jor  g27791(.dina(n27959), .dinb(n27958), .dout(n27960));
  jand g27792(.dina(n23146), .dinb(n5076), .dout(n27961));
  jand g27793(.dina(n23144), .dinb(n5084), .dout(n27962));
  jand g27794(.dina(n23079), .dinb(n5082), .dout(n27963));
  jand g27795(.dina(n23080), .dinb(n6050), .dout(n27964));
  jor  g27796(.dina(n27964), .dinb(n27963), .dout(n27965));
  jor  g27797(.dina(n27965), .dinb(n27962), .dout(n27966));
  jor  g27798(.dina(n27966), .dinb(n27961), .dout(n27967));
  jor  g27799(.dina(n27917), .dinb(n27845), .dout(n27968));
  jand g27800(.dina(n27920), .dinb(n27918), .dout(n27969));
  jnot g27801(.din(n27969), .dout(n27970));
  jand g27802(.dina(n27970), .dinb(n27968), .dout(n27971));
  jand g27803(.dina(n1246), .dinb(n948), .dout(n27972));
  jand g27804(.dina(n27972), .dinb(n964), .dout(n27973));
  jand g27805(.dina(n1577), .dinb(n3185), .dout(n27974));
  jand g27806(.dina(n5415), .dinb(n1852), .dout(n27975));
  jand g27807(.dina(n27975), .dinb(n27974), .dout(n27976));
  jand g27808(.dina(n27976), .dinb(n27973), .dout(n27977));
  jand g27809(.dina(n27977), .dinb(n2331), .dout(n27978));
  jand g27810(.dina(n3758), .dinb(n554), .dout(n27979));
  jand g27811(.dina(n27979), .dinb(n6368), .dout(n27980));
  jand g27812(.dina(n27980), .dinb(n18825), .dout(n27981));
  jand g27813(.dina(n27981), .dinb(n7241), .dout(n27982));
  jand g27814(.dina(n27982), .dinb(n27978), .dout(n27983));
  jand g27815(.dina(n7813), .dinb(n6471), .dout(n27984));
  jand g27816(.dina(n27984), .dinb(n16198), .dout(n27985));
  jand g27817(.dina(n27985), .dinb(n27983), .dout(n27986));
  jand g27818(.dina(n27986), .dinb(n23106), .dout(n27987));
  jnot g27819(.din(n27987), .dout(n27988));
  jxor g27820(.dina(n27988), .dinb(n27971), .dout(n27989));
  jxor g27821(.dina(n27989), .dinb(n27967), .dout(n27990));
  jxor g27822(.dina(n27990), .dinb(n27960), .dout(n27991));
  jnot g27823(.din(n27991), .dout(n27992));
  jor  g27824(.dina(n24302), .dinb(n4343), .dout(n27993));
  jor  g27825(.dina(n24266), .dinb(n4346), .dout(n27994));
  jor  g27826(.dina(n24304), .dinb(n4348), .dout(n27995));
  jand g27827(.dina(n27995), .dinb(n27994), .dout(n27996));
  jor  g27828(.dina(n24265), .dinb(n3683), .dout(n27997));
  jand g27829(.dina(n27997), .dinb(n27996), .dout(n27998));
  jand g27830(.dina(n27998), .dinb(n27993), .dout(n27999));
  jxor g27831(.dina(n27999), .dinb(\a[29] ), .dout(n28000));
  jxor g27832(.dina(n28000), .dinb(n27992), .dout(n28001));
  jxor g27833(.dina(n28001), .dinb(n27957), .dout(n28002));
  jor  g27834(.dina(n24932), .dinb(n2303), .dout(n28003));
  jor  g27835(.dina(n24738), .dinb(n2306), .dout(n28004));
  jor  g27836(.dina(n24930), .dinb(n2309), .dout(n28005));
  jand g27837(.dina(n28005), .dinb(n28004), .dout(n28006));
  jor  g27838(.dina(n24518), .dinb(n1805), .dout(n28007));
  jand g27839(.dina(n28007), .dinb(n28006), .dout(n28008));
  jand g27840(.dina(n28008), .dinb(n28003), .dout(n28009));
  jxor g27841(.dina(n28009), .dinb(\a[26] ), .dout(n28010));
  jnot g27842(.din(n28010), .dout(n28011));
  jxor g27843(.dina(n28011), .dinb(n28002), .dout(n28012));
  jxor g27844(.dina(n28012), .dinb(n27954), .dout(n28013));
  jxor g27845(.dina(n28013), .dinb(n27949), .dout(n28014));
  jxor g27846(.dina(n28014), .dinb(n27946), .dout(\result[29] ));
  jnot g27847(.din(n27946), .dout(n28016));
  jnot g27848(.din(n28014), .dout(n28017));
  jor  g27849(.dina(n28017), .dinb(n28016), .dout(n28018));
  jand g27850(.dina(n28012), .dinb(n27954), .dout(n28019));
  jand g27851(.dina(n28013), .dinb(n27949), .dout(n28020));
  jor  g27852(.dina(n28020), .dinb(n28019), .dout(n28021));
  jand g27853(.dina(n28001), .dinb(n27957), .dout(n28022));
  jand g27854(.dina(n28011), .dinb(n28002), .dout(n28023));
  jor  g27855(.dina(n28023), .dinb(n28022), .dout(n28024));
  jand g27856(.dina(n27990), .dinb(n27960), .dout(n28025));
  jnot g27857(.din(n28025), .dout(n28026));
  jor  g27858(.dina(n28000), .dinb(n27992), .dout(n28027));
  jand g27859(.dina(n28027), .dinb(n28026), .dout(n28028));
  jnot g27860(.din(n28028), .dout(n28029));
  jand g27861(.dina(n23847), .dinb(n5076), .dout(n28030));
  jand g27862(.dina(n23845), .dinb(n5084), .dout(n28031));
  jand g27863(.dina(n23144), .dinb(n5082), .dout(n28032));
  jand g27864(.dina(n23079), .dinb(n6050), .dout(n28033));
  jor  g27865(.dina(n28033), .dinb(n28032), .dout(n28034));
  jor  g27866(.dina(n28034), .dinb(n28031), .dout(n28035));
  jor  g27867(.dina(n28035), .dinb(n28030), .dout(n28036));
  jnot g27868(.din(n27971), .dout(n28037));
  jand g27869(.dina(n27987), .dinb(n28037), .dout(n28038));
  jand g27870(.dina(n27989), .dinb(n27967), .dout(n28039));
  jor  g27871(.dina(n28039), .dinb(n28038), .dout(n28040));
  jnot g27872(.din(n27986), .dout(n28041));
  jand g27873(.dina(n7643), .dinb(n7272), .dout(n28042));
  jand g27874(.dina(n28042), .dinb(n1895), .dout(n28043));
  jand g27875(.dina(n28043), .dinb(n7677), .dout(n28044));
  jand g27876(.dina(n7261), .dinb(n1316), .dout(n28045));
  jand g27877(.dina(n28045), .dinb(n16329), .dout(n28046));
  jand g27878(.dina(n28046), .dinb(n28044), .dout(n28047));
  jand g27879(.dina(n28047), .dinb(n23106), .dout(n28048));
  jand g27880(.dina(n28048), .dinb(n28041), .dout(n28049));
  jnot g27881(.din(n28049), .dout(n28050));
  jor  g27882(.dina(n28047), .dinb(n27988), .dout(n28051));
  jand g27883(.dina(n28051), .dinb(n28050), .dout(n28052));
  jxor g27884(.dina(n28052), .dinb(n28040), .dout(n28053));
  jxor g27885(.dina(n28053), .dinb(n28036), .dout(n28054));
  jxor g27886(.dina(n28054), .dinb(n28029), .dout(n28055));
  jor  g27887(.dina(n25116), .dinb(n2303), .dout(n28056));
  jor  g27888(.dina(n24930), .dinb(n23060), .dout(n28057));
  jor  g27889(.dina(n24738), .dinb(n1805), .dout(n28058));
  jand g27890(.dina(n28058), .dinb(n28057), .dout(n28059));
  jand g27891(.dina(n28059), .dinb(n28056), .dout(n28060));
  jxor g27892(.dina(n28060), .dinb(\a[26] ), .dout(n28061));
  jor  g27893(.dina(n24516), .dinb(n4343), .dout(n28062));
  jor  g27894(.dina(n24304), .dinb(n4346), .dout(n28063));
  jor  g27895(.dina(n24518), .dinb(n4348), .dout(n28064));
  jand g27896(.dina(n28064), .dinb(n28063), .dout(n28065));
  jor  g27897(.dina(n24266), .dinb(n3683), .dout(n28066));
  jand g27898(.dina(n28066), .dinb(n28065), .dout(n28067));
  jand g27899(.dina(n28067), .dinb(n28062), .dout(n28068));
  jxor g27900(.dina(n28068), .dinb(\a[29] ), .dout(n28069));
  jxor g27901(.dina(n28069), .dinb(n28061), .dout(n28070));
  jxor g27902(.dina(n28070), .dinb(n28055), .dout(n28071));
  jxor g27903(.dina(n28071), .dinb(n28024), .dout(n28072));
  jnot g27904(.din(n28072), .dout(n28073));
  jxor g27905(.dina(n28073), .dinb(n28021), .dout(n28074));
  jxor g27906(.dina(n28074), .dinb(n28018), .dout(\result[30] ));
  jor  g27907(.dina(n28074), .dinb(n28018), .dout(n28076));
  jand g27908(.dina(n28071), .dinb(n28024), .dout(n28077));
  jand g27909(.dina(n28072), .dinb(n28021), .dout(n28078));
  jor  g27910(.dina(n28078), .dinb(n28077), .dout(n28079));
  jand g27911(.dina(n7997), .dinb(n7665), .dout(n28080));
  jxor g27912(.dina(n28080), .dinb(n27987), .dout(n28081));
  jxor g27913(.dina(n28081), .dinb(n77), .dout(n28082));
  jand g27914(.dina(n28053), .dinb(n28036), .dout(n28083));
  jand g27915(.dina(n28054), .dinb(n28029), .dout(n28084));
  jor  g27916(.dina(n28084), .dinb(n28083), .dout(n28085));
  jnot g27917(.din(n28051), .dout(n28086));
  jand g27918(.dina(n28052), .dinb(n28040), .dout(n28087));
  jor  g27919(.dina(n28087), .dinb(n28086), .dout(n28088));
  jand g27920(.dina(n24077), .dinb(n5076), .dout(n28089));
  jand g27921(.dina(n24075), .dinb(n5084), .dout(n28090));
  jand g27922(.dina(n23845), .dinb(n5082), .dout(n28091));
  jand g27923(.dina(n23144), .dinb(n6050), .dout(n28092));
  jor  g27924(.dina(n28092), .dinb(n28091), .dout(n28093));
  jor  g27925(.dina(n28093), .dinb(n28090), .dout(n28094));
  jor  g27926(.dina(n28094), .dinb(n28089), .dout(n28095));
  jor  g27927(.dina(n24736), .dinb(n4343), .dout(n28096));
  jor  g27928(.dina(n24738), .dinb(n4348), .dout(n28097));
  jor  g27929(.dina(n24518), .dinb(n4346), .dout(n28098));
  jor  g27930(.dina(n24304), .dinb(n3683), .dout(n28099));
  jand g27931(.dina(n28099), .dinb(n28098), .dout(n28100));
  jand g27932(.dina(n28100), .dinb(n28097), .dout(n28101));
  jand g27933(.dina(n28101), .dinb(n28096), .dout(n28102));
  jxor g27934(.dina(n28102), .dinb(n93), .dout(n28103));
  jxor g27935(.dina(n28103), .dinb(n28095), .dout(n28104));
  jxor g27936(.dina(n28104), .dinb(n28088), .dout(n28105));
  jxor g27937(.dina(n28105), .dinb(n28085), .dout(n28106));
  jxor g27938(.dina(n28106), .dinb(n28082), .dout(n28107));
  jor  g27939(.dina(n28069), .dinb(n28061), .dout(n28108));
  jnot g27940(.din(n28055), .dout(n28109));
  jnot g27941(.din(n28070), .dout(n28110));
  jor  g27942(.dina(n28110), .dinb(n28109), .dout(n28111));
  jand g27943(.dina(n28111), .dinb(n28108), .dout(n28112));
  jand g27944(.dina(n25199), .dinb(n23113), .dout(n28113));
  jxor g27945(.dina(n28113), .dinb(n28112), .dout(n28114));
  jxor g27946(.dina(n28114), .dinb(n28107), .dout(n28115));
  jxor g27947(.dina(n28115), .dinb(n28079), .dout(n28116));
  jxor g27948(.dina(n28116), .dinb(n28076), .dout(\result[31] ));
endmodule


