// Benchmark "c880" written by ABC on Sun May 24 21:28:53 2020

module c880 ( 
    G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat,
    G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat,
    G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat,
    G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat,
    G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat,
    G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat,
    G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat,
    G267gat, G268gat,
    G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat,
    G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat,
    G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat,
    G879gat, G880gat  );
  input  G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat,
    G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat,
    G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat,
    G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat,
    G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat,
    G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat,
    G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat,
    G261gat, G267gat, G268gat;
  output G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat,
    G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat,
    G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat,
    G878gat, G879gat, G880gat;
  wire n86, n88, n92, n93, n95, n96, n97, n98, n99, n100, n101, n103, n104,
    n105, n107, n108, n109, n111, n113, n115, n117, n119, n120, n122, n123,
    n126, n127, n128, n129, n130, n131, n132, n133, n135, n136, n137, n138,
    n139, n140, n141, n142, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431;
  jand g000(.dina(G75gat), .dinb(G29gat), .dout(n86));
  jand g001(.dina(n86), .dinb(G42gat), .dout(G388gat));
  jand g002(.dina(G36gat), .dinb(G29gat), .dout(n88));
  jand g003(.dina(n88), .dinb(G80gat), .dout(G389gat));
  jand g004(.dina(n88), .dinb(G42gat), .dout(G390gat));
  jand g005(.dina(G86gat), .dinb(G85gat), .dout(G391gat));
  jand g006(.dina(G8gat), .dinb(G1gat), .dout(n92));
  jand g007(.dina(n92), .dinb(G13gat), .dout(n93));
  jand g008(.dina(n93), .dinb(G17gat), .dout(G418gat));
  jnot g009(.din(G17gat), .dout(n95));
  jnot g010(.din(G13gat), .dout(n96));
  jnot g011(.din(G1gat), .dout(n97));
  jnot g012(.din(G26gat), .dout(n98));
  jor  g013(.dina(n98), .dinb(n97), .dout(n99));
  jor  g014(.dina(n99), .dinb(n96), .dout(n100));
  jor  g015(.dina(n100), .dinb(n95), .dout(n101));
  jor  g016(.dina(n101), .dinb(G390gat), .dout(G419gat));
  jnot g017(.din(G80gat), .dout(n103));
  jand g018(.dina(G75gat), .dinb(G59gat), .dout(n104));
  jnot g019(.din(n104), .dout(n105));
  jor  g020(.dina(n105), .dinb(n103), .dout(G420gat));
  jnot g021(.din(G36gat), .dout(n107));
  jnot g022(.din(G59gat), .dout(n108));
  jor  g023(.dina(n108), .dinb(n107), .dout(n109));
  jor  g024(.dina(n109), .dinb(n103), .dout(G421gat));
  jnot g025(.din(G42gat), .dout(n111));
  jor  g026(.dina(n109), .dinb(n111), .dout(G422gat));
  jor  g027(.dina(G88gat), .dinb(G87gat), .dout(n113));
  jand g028(.dina(n113), .dinb(G90gat), .dout(G423gat));
  jnot g029(.din(G390gat), .dout(n115));
  jor  g030(.dina(n101), .dinb(n115), .dout(G446gat));
  jand g031(.dina(G26gat), .dinb(G1gat), .dout(n117));
  jand g032(.dina(n117), .dinb(G51gat), .dout(G447gat));
  jand g033(.dina(n93), .dinb(G55gat), .dout(n119));
  jand g034(.dina(n119), .dinb(G29gat), .dout(n120));
  jand g035(.dina(n120), .dinb(G68gat), .dout(G448gat));
  jand g036(.dina(G68gat), .dinb(G59gat), .dout(n122));
  jand g037(.dina(n119), .dinb(G74gat), .dout(n123));
  jand g038(.dina(n123), .dinb(n122), .dout(G449gat));
  jand g039(.dina(n113), .dinb(G89gat), .dout(G450gat));
  jxor g040(.dina(G116gat), .dinb(G111gat), .dout(n126));
  jxor g041(.dina(n126), .dinb(G135gat), .dout(n127));
  jxor g042(.dina(G96gat), .dinb(G91gat), .dout(n128));
  jxor g043(.dina(n128), .dinb(G130gat), .dout(n129));
  jxor g044(.dina(G106gat), .dinb(G101gat), .dout(n130));
  jxor g045(.dina(G126gat), .dinb(G121gat), .dout(n131));
  jxor g046(.dina(n131), .dinb(n130), .dout(n132));
  jxor g047(.dina(n132), .dinb(n129), .dout(n133));
  jxor g048(.dina(n133), .dinb(n127), .dout(G767gat));
  jxor g049(.dina(G189gat), .dinb(G183gat), .dout(n135));
  jxor g050(.dina(n135), .dinb(G207gat), .dout(n136));
  jxor g051(.dina(G159gat), .dinb(G130gat), .dout(n137));
  jxor g052(.dina(n137), .dinb(G165gat), .dout(n138));
  jxor g053(.dina(G177gat), .dinb(G171gat), .dout(n139));
  jxor g054(.dina(G201gat), .dinb(G195gat), .dout(n140));
  jxor g055(.dina(n140), .dinb(n139), .dout(n141));
  jxor g056(.dina(n141), .dinb(n138), .dout(n142));
  jxor g057(.dina(n142), .dinb(n136), .dout(G768gat));
  jnot g058(.din(G268gat), .dout(n144));
  jand g059(.dina(G447gat), .dinb(G80gat), .dout(n145));
  jand g060(.dina(n145), .dinb(n86), .dout(n146));
  jand g061(.dina(n146), .dinb(G55gat), .dout(n147));
  jand g062(.dina(n147), .dinb(n144), .dout(n148));
  jand g063(.dina(n111), .dinb(n95), .dout(n149));
  jnot g064(.din(n149), .dout(n150));
  jand g065(.dina(G156gat), .dinb(G59gat), .dout(n151));
  jand g066(.dina(G42gat), .dinb(G17gat), .dout(n152));
  jnot g067(.din(n152), .dout(n153));
  jand g068(.dina(n153), .dinb(n151), .dout(n154));
  jand g069(.dina(n154), .dinb(G447gat), .dout(n155));
  jand g070(.dina(n155), .dinb(n150), .dout(n156));
  jnot g071(.din(n92), .dout(n157));
  jand g072(.dina(n104), .dinb(G42gat), .dout(n158));
  jand g073(.dina(G51gat), .dinb(G17gat), .dout(n159));
  jnot g074(.din(n159), .dout(n160));
  jor  g075(.dina(n160), .dinb(n158), .dout(n161));
  jor  g076(.dina(n161), .dinb(n157), .dout(n162));
  jnot g077(.din(n162), .dout(n163));
  jor  g078(.dina(n163), .dinb(n156), .dout(n164));
  jand g079(.dina(n164), .dinb(G126gat), .dout(n165));
  jnot g080(.din(G156gat), .dout(n166));
  jor  g081(.dina(n166), .dinb(n108), .dout(n167));
  jand g082(.dina(n167), .dinb(G447gat), .dout(n168));
  jand g083(.dina(n168), .dinb(G17gat), .dout(n169));
  jor  g084(.dina(n169), .dinb(n97), .dout(n170));
  jand g085(.dina(n170), .dinb(G153gat), .dout(n171));
  jor  g086(.dina(n171), .dinb(n165), .dout(n172));
  jor  g087(.dina(n172), .dinb(n148), .dout(n173));
  jand g088(.dina(n173), .dinb(G246gat), .dout(n174));
  jand g089(.dina(n122), .dinb(G42gat), .dout(n175));
  jand g090(.dina(G73gat), .dinb(G72gat), .dout(n176));
  jand g091(.dina(n176), .dinb(n175), .dout(n177));
  jand g092(.dina(n177), .dinb(n119), .dout(n178));
  jand g093(.dina(n178), .dinb(G201gat), .dout(n179));
  jor  g094(.dina(n179), .dinb(n174), .dout(n180));
  jnot g095(.din(G201gat), .dout(n181));
  jnot g096(.din(n148), .dout(n182));
  jnot g097(.din(G126gat), .dout(n183));
  jnot g098(.din(G51gat), .dout(n184));
  jor  g099(.dina(n99), .dinb(n184), .dout(n185));
  jor  g100(.dina(n152), .dinb(n167), .dout(n186));
  jor  g101(.dina(n186), .dinb(n185), .dout(n187));
  jor  g102(.dina(n187), .dinb(n149), .dout(n188));
  jand g103(.dina(n162), .dinb(n188), .dout(n189));
  jor  g104(.dina(n189), .dinb(n183), .dout(n190));
  jnot g105(.din(G153gat), .dout(n191));
  jor  g106(.dina(n151), .dinb(n185), .dout(n192));
  jor  g107(.dina(n192), .dinb(n95), .dout(n193));
  jand g108(.dina(n193), .dinb(G1gat), .dout(n194));
  jor  g109(.dina(n194), .dinb(n191), .dout(n195));
  jand g110(.dina(n195), .dinb(n190), .dout(n196));
  jand g111(.dina(n196), .dinb(n182), .dout(n197));
  jxor g112(.dina(n197), .dinb(n181), .dout(n198));
  jand g113(.dina(n198), .dinb(G228gat), .dout(n199));
  jand g114(.dina(n173), .dinb(G201gat), .dout(n200));
  jand g115(.dina(n200), .dinb(G237gat), .dout(n201));
  jand g116(.dina(G210gat), .dinb(G121gat), .dout(n202));
  jand g117(.dina(G267gat), .dinb(G255gat), .dout(n203));
  jor  g118(.dina(n203), .dinb(n202), .dout(n204));
  jor  g119(.dina(n204), .dinb(n201), .dout(n205));
  jor  g120(.dina(n205), .dinb(n199), .dout(n206));
  jor  g121(.dina(n206), .dinb(n180), .dout(n207));
  jor  g122(.dina(n198), .dinb(G261gat), .dout(n208));
  jnot g123(.din(G261gat), .dout(n209));
  jnot g124(.din(n198), .dout(n210));
  jor  g125(.dina(n210), .dinb(n209), .dout(n211));
  jand g126(.dina(n211), .dinb(G219gat), .dout(n212));
  jand g127(.dina(n212), .dinb(n208), .dout(n213));
  jor  g128(.dina(n213), .dinb(n207), .dout(G850gat));
  jand g129(.dina(n164), .dinb(G111gat), .dout(n215));
  jand g130(.dina(n170), .dinb(G143gat), .dout(n216));
  jor  g131(.dina(n216), .dinb(n148), .dout(n217));
  jor  g132(.dina(n217), .dinb(n215), .dout(n218));
  jxor g133(.dina(n218), .dinb(G183gat), .dout(n219));
  jand g134(.dina(n219), .dinb(G228gat), .dout(n220));
  jand g135(.dina(n178), .dinb(G183gat), .dout(n221));
  jand g136(.dina(n218), .dinb(G183gat), .dout(n222));
  jand g137(.dina(n222), .dinb(G237gat), .dout(n223));
  jand g138(.dina(n218), .dinb(G246gat), .dout(n224));
  jand g139(.dina(G210gat), .dinb(G106gat), .dout(n225));
  jor  g140(.dina(n225), .dinb(n224), .dout(n226));
  jor  g141(.dina(n226), .dinb(n223), .dout(n227));
  jor  g142(.dina(n227), .dinb(n221), .dout(n228));
  jor  g143(.dina(n228), .dinb(n220), .dout(n229));
  jand g144(.dina(n164), .dinb(G116gat), .dout(n230));
  jand g145(.dina(n170), .dinb(G146gat), .dout(n231));
  jor  g146(.dina(n231), .dinb(n148), .dout(n232));
  jor  g147(.dina(n232), .dinb(n230), .dout(n233));
  jand g148(.dina(n233), .dinb(G189gat), .dout(n234));
  jor  g149(.dina(n233), .dinb(G189gat), .dout(n235));
  jand g150(.dina(n164), .dinb(G121gat), .dout(n236));
  jand g151(.dina(n170), .dinb(G149gat), .dout(n237));
  jor  g152(.dina(n237), .dinb(n148), .dout(n238));
  jor  g153(.dina(n238), .dinb(n236), .dout(n239));
  jand g154(.dina(n239), .dinb(G195gat), .dout(n240));
  jor  g155(.dina(n239), .dinb(G195gat), .dout(n241));
  jand g156(.dina(n197), .dinb(n181), .dout(n242));
  jnot g157(.din(n242), .dout(n243));
  jor  g158(.dina(n200), .dinb(G261gat), .dout(n244));
  jand g159(.dina(n244), .dinb(n243), .dout(n245));
  jand g160(.dina(n245), .dinb(n241), .dout(n246));
  jor  g161(.dina(n246), .dinb(n240), .dout(n247));
  jand g162(.dina(n247), .dinb(n235), .dout(n248));
  jor  g163(.dina(n248), .dinb(n234), .dout(n249));
  jor  g164(.dina(n249), .dinb(n219), .dout(n250));
  jnot g165(.din(n219), .dout(n251));
  jnot g166(.din(n234), .dout(n252));
  jnot g167(.din(n235), .dout(n253));
  jnot g168(.din(n240), .dout(n254));
  jnot g169(.din(n241), .dout(n255));
  jor  g170(.dina(n197), .dinb(n181), .dout(n256));
  jand g171(.dina(n256), .dinb(n209), .dout(n257));
  jor  g172(.dina(n257), .dinb(n242), .dout(n258));
  jor  g173(.dina(n258), .dinb(n255), .dout(n259));
  jand g174(.dina(n259), .dinb(n254), .dout(n260));
  jor  g175(.dina(n260), .dinb(n253), .dout(n261));
  jand g176(.dina(n261), .dinb(n252), .dout(n262));
  jor  g177(.dina(n262), .dinb(n251), .dout(n263));
  jand g178(.dina(n263), .dinb(G219gat), .dout(n264));
  jand g179(.dina(n264), .dinb(n250), .dout(n265));
  jor  g180(.dina(n265), .dinb(n229), .dout(G863gat));
  jxor g181(.dina(n233), .dinb(G189gat), .dout(n267));
  jand g182(.dina(n267), .dinb(G228gat), .dout(n268));
  jand g183(.dina(G210gat), .dinb(G111gat), .dout(n269));
  jand g184(.dina(G237gat), .dinb(G189gat), .dout(n270));
  jor  g185(.dina(n270), .dinb(G246gat), .dout(n271));
  jand g186(.dina(n271), .dinb(n233), .dout(n272));
  jor  g187(.dina(n272), .dinb(n269), .dout(n273));
  jand g188(.dina(G259gat), .dinb(G255gat), .dout(n274));
  jand g189(.dina(n178), .dinb(G189gat), .dout(n275));
  jor  g190(.dina(n275), .dinb(n274), .dout(n276));
  jor  g191(.dina(n276), .dinb(n273), .dout(n277));
  jor  g192(.dina(n277), .dinb(n268), .dout(n278));
  jor  g193(.dina(n267), .dinb(n247), .dout(n279));
  jnot g194(.din(n267), .dout(n280));
  jor  g195(.dina(n280), .dinb(n260), .dout(n281));
  jand g196(.dina(n281), .dinb(G219gat), .dout(n282));
  jand g197(.dina(n282), .dinb(n279), .dout(n283));
  jor  g198(.dina(n283), .dinb(n278), .dout(G864gat));
  jxor g199(.dina(n239), .dinb(G195gat), .dout(n285));
  jand g200(.dina(n285), .dinb(G228gat), .dout(n286));
  jand g201(.dina(G210gat), .dinb(G116gat), .dout(n287));
  jand g202(.dina(G237gat), .dinb(G195gat), .dout(n288));
  jor  g203(.dina(n288), .dinb(G246gat), .dout(n289));
  jand g204(.dina(n289), .dinb(n239), .dout(n290));
  jor  g205(.dina(n290), .dinb(n287), .dout(n291));
  jand g206(.dina(n178), .dinb(G195gat), .dout(n292));
  jand g207(.dina(G260gat), .dinb(G255gat), .dout(n293));
  jor  g208(.dina(n293), .dinb(n292), .dout(n294));
  jor  g209(.dina(n294), .dinb(n291), .dout(n295));
  jor  g210(.dina(n295), .dinb(n286), .dout(n296));
  jor  g211(.dina(n285), .dinb(n245), .dout(n297));
  jnot g212(.din(n285), .dout(n298));
  jor  g213(.dina(n298), .dinb(n258), .dout(n299));
  jand g214(.dina(n299), .dinb(G219gat), .dout(n300));
  jand g215(.dina(n300), .dinb(n297), .dout(n301));
  jor  g216(.dina(n301), .dinb(n296), .dout(G865gat));
  jand g217(.dina(n168), .dinb(G55gat), .dout(n303));
  jand g218(.dina(n303), .dinb(G143gat), .dout(n304));
  jand g219(.dina(n146), .dinb(G17gat), .dout(n305));
  jand g220(.dina(n305), .dinb(n144), .dout(n306));
  jor  g221(.dina(n306), .dinb(n304), .dout(n307));
  jand g222(.dina(n164), .dinb(G91gat), .dout(n308));
  jand g223(.dina(G138gat), .dinb(G8gat), .dout(n309));
  jor  g224(.dina(n309), .dinb(n308), .dout(n310));
  jor  g225(.dina(n310), .dinb(n307), .dout(n311));
  jand g226(.dina(n311), .dinb(G159gat), .dout(n312));
  jor  g227(.dina(n311), .dinb(G159gat), .dout(n313));
  jand g228(.dina(n164), .dinb(G96gat), .dout(n314));
  jand g229(.dina(n303), .dinb(G146gat), .dout(n315));
  jand g230(.dina(G138gat), .dinb(G51gat), .dout(n316));
  jor  g231(.dina(n316), .dinb(n315), .dout(n317));
  jor  g232(.dina(n317), .dinb(n314), .dout(n318));
  jor  g233(.dina(n318), .dinb(n306), .dout(n319));
  jand g234(.dina(n319), .dinb(G165gat), .dout(n320));
  jor  g235(.dina(n319), .dinb(G165gat), .dout(n321));
  jand g236(.dina(n164), .dinb(G101gat), .dout(n322));
  jand g237(.dina(n303), .dinb(G149gat), .dout(n323));
  jand g238(.dina(G138gat), .dinb(G17gat), .dout(n324));
  jor  g239(.dina(n324), .dinb(n323), .dout(n325));
  jor  g240(.dina(n325), .dinb(n322), .dout(n326));
  jor  g241(.dina(n326), .dinb(n306), .dout(n327));
  jand g242(.dina(n327), .dinb(G171gat), .dout(n328));
  jor  g243(.dina(n327), .dinb(G171gat), .dout(n329));
  jand g244(.dina(n164), .dinb(G106gat), .dout(n330));
  jand g245(.dina(n303), .dinb(G153gat), .dout(n331));
  jand g246(.dina(G152gat), .dinb(G138gat), .dout(n332));
  jor  g247(.dina(n332), .dinb(n331), .dout(n333));
  jor  g248(.dina(n333), .dinb(n330), .dout(n334));
  jor  g249(.dina(n334), .dinb(n306), .dout(n335));
  jand g250(.dina(n335), .dinb(G177gat), .dout(n336));
  jnot g251(.din(G177gat), .dout(n337));
  jnot g252(.din(n335), .dout(n338));
  jand g253(.dina(n338), .dinb(n337), .dout(n339));
  jnot g254(.din(n339), .dout(n340));
  jnot g255(.din(G183gat), .dout(n341));
  jnot g256(.din(n218), .dout(n342));
  jand g257(.dina(n342), .dinb(n341), .dout(n343));
  jnot g258(.din(n343), .dout(n344));
  jand g259(.dina(n249), .dinb(n344), .dout(n345));
  jor  g260(.dina(n345), .dinb(n222), .dout(n346));
  jand g261(.dina(n346), .dinb(n340), .dout(n347));
  jor  g262(.dina(n347), .dinb(n336), .dout(n348));
  jand g263(.dina(n348), .dinb(n329), .dout(n349));
  jor  g264(.dina(n349), .dinb(n328), .dout(n350));
  jand g265(.dina(n350), .dinb(n321), .dout(n351));
  jor  g266(.dina(n351), .dinb(n320), .dout(n352));
  jand g267(.dina(n352), .dinb(n313), .dout(n353));
  jor  g268(.dina(n353), .dinb(n312), .dout(G866gat));
  jxor g269(.dina(n335), .dinb(G177gat), .dout(n355));
  jnot g270(.din(n355), .dout(n356));
  jand g271(.dina(n346), .dinb(G219gat), .dout(n357));
  jand g272(.dina(n357), .dinb(n356), .dout(n358));
  jnot g273(.din(n222), .dout(n359));
  jor  g274(.dina(n262), .dinb(n343), .dout(n360));
  jand g275(.dina(n360), .dinb(n359), .dout(n361));
  jand g276(.dina(n361), .dinb(G219gat), .dout(n362));
  jor  g277(.dina(n362), .dinb(G228gat), .dout(n363));
  jand g278(.dina(n363), .dinb(n355), .dout(n364));
  jand g279(.dina(n336), .dinb(G237gat), .dout(n365));
  jand g280(.dina(n335), .dinb(G246gat), .dout(n366));
  jand g281(.dina(G210gat), .dinb(G101gat), .dout(n367));
  jand g282(.dina(n178), .dinb(G177gat), .dout(n368));
  jor  g283(.dina(n368), .dinb(n367), .dout(n369));
  jor  g284(.dina(n369), .dinb(n366), .dout(n370));
  jor  g285(.dina(n370), .dinb(n365), .dout(n371));
  jor  g286(.dina(n371), .dinb(n364), .dout(n372));
  jor  g287(.dina(n372), .dinb(n358), .dout(G874gat));
  jand g288(.dina(n311), .dinb(G237gat), .dout(n374));
  jor  g289(.dina(n374), .dinb(n178), .dout(n375));
  jand g290(.dina(n375), .dinb(G159gat), .dout(n376));
  jxor g291(.dina(n311), .dinb(G159gat), .dout(n377));
  jand g292(.dina(n377), .dinb(G228gat), .dout(n378));
  jand g293(.dina(G268gat), .dinb(G210gat), .dout(n379));
  jor  g294(.dina(n379), .dinb(n378), .dout(n380));
  jand g295(.dina(n311), .dinb(G246gat), .dout(n381));
  jor  g296(.dina(n381), .dinb(n380), .dout(n382));
  jor  g297(.dina(n382), .dinb(n376), .dout(n383));
  jor  g298(.dina(n377), .dinb(n352), .dout(n384));
  jnot g299(.din(n320), .dout(n385));
  jnot g300(.din(n321), .dout(n386));
  jnot g301(.din(n328), .dout(n387));
  jnot g302(.din(n329), .dout(n388));
  jnot g303(.din(n336), .dout(n389));
  jor  g304(.dina(n361), .dinb(n339), .dout(n390));
  jand g305(.dina(n390), .dinb(n389), .dout(n391));
  jor  g306(.dina(n391), .dinb(n388), .dout(n392));
  jand g307(.dina(n392), .dinb(n387), .dout(n393));
  jor  g308(.dina(n393), .dinb(n386), .dout(n394));
  jand g309(.dina(n394), .dinb(n385), .dout(n395));
  jnot g310(.din(n377), .dout(n396));
  jor  g311(.dina(n396), .dinb(n395), .dout(n397));
  jand g312(.dina(n397), .dinb(G219gat), .dout(n398));
  jand g313(.dina(n398), .dinb(n384), .dout(n399));
  jor  g314(.dina(n399), .dinb(n383), .dout(G878gat));
  jand g315(.dina(n319), .dinb(G237gat), .dout(n401));
  jor  g316(.dina(n401), .dinb(n178), .dout(n402));
  jand g317(.dina(n402), .dinb(G165gat), .dout(n403));
  jxor g318(.dina(n319), .dinb(G165gat), .dout(n404));
  jand g319(.dina(n404), .dinb(G228gat), .dout(n405));
  jand g320(.dina(G210gat), .dinb(G91gat), .dout(n406));
  jor  g321(.dina(n406), .dinb(n405), .dout(n407));
  jand g322(.dina(n319), .dinb(G246gat), .dout(n408));
  jor  g323(.dina(n408), .dinb(n407), .dout(n409));
  jor  g324(.dina(n409), .dinb(n403), .dout(n410));
  jor  g325(.dina(n404), .dinb(n350), .dout(n411));
  jnot g326(.din(n404), .dout(n412));
  jor  g327(.dina(n412), .dinb(n393), .dout(n413));
  jand g328(.dina(n413), .dinb(G219gat), .dout(n414));
  jand g329(.dina(n414), .dinb(n411), .dout(n415));
  jor  g330(.dina(n415), .dinb(n410), .dout(G879gat));
  jand g331(.dina(n327), .dinb(G237gat), .dout(n417));
  jor  g332(.dina(n417), .dinb(n178), .dout(n418));
  jand g333(.dina(n418), .dinb(G171gat), .dout(n419));
  jxor g334(.dina(n327), .dinb(G171gat), .dout(n420));
  jand g335(.dina(n420), .dinb(G228gat), .dout(n421));
  jand g336(.dina(G210gat), .dinb(G96gat), .dout(n422));
  jor  g337(.dina(n422), .dinb(n421), .dout(n423));
  jand g338(.dina(n327), .dinb(G246gat), .dout(n424));
  jor  g339(.dina(n424), .dinb(n423), .dout(n425));
  jor  g340(.dina(n425), .dinb(n419), .dout(n426));
  jnot g341(.din(n420), .dout(n427));
  jor  g342(.dina(n427), .dinb(n391), .dout(n428));
  jor  g343(.dina(n420), .dinb(n348), .dout(n429));
  jand g344(.dina(n429), .dinb(G219gat), .dout(n430));
  jand g345(.dina(n430), .dinb(n428), .dout(n431));
  jor  g346(.dina(n431), .dinb(n426), .dout(G880gat));
endmodule


