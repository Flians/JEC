/*

c7552:
	jxor: 242
	jspl: 295
	jspl3: 359
	jnot: 215
	jdff: 3112
	jor: 391
	jand: 479

Summary:
	jxor: 242
	jspl: 295
	jspl3: 359
	jnot: 215
	jdff: 3112
	jor: 391
	jand: 479

The maximum logic level gap of any gate:
	c7552: 35
*/

module gf_c7552(gclk, G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399);
	input gclk;
	input G1;
	input G5;
	input G9;
	input G12;
	input G15;
	input G18;
	input G23;
	input G26;
	input G29;
	input G32;
	input G35;
	input G38;
	input G41;
	input G44;
	input G47;
	input G50;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G69;
	input G70;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G118;
	input G121;
	input G124;
	input G127;
	input G130;
	input G133;
	input G134;
	input G135;
	input G138;
	input G141;
	input G144;
	input G147;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G158;
	input G159;
	input G160;
	input G161;
	input G162;
	input G163;
	input G164;
	input G165;
	input G166;
	input G167;
	input G168;
	input G169;
	input G170;
	input G171;
	input G172;
	input G173;
	input G174;
	input G175;
	input G176;
	input G177;
	input G178;
	input G179;
	input G180;
	input G181;
	input G182;
	input G183;
	input G184;
	input G185;
	input G186;
	input G187;
	input G188;
	input G189;
	input G190;
	input G191;
	input G192;
	input G193;
	input G194;
	input G195;
	input G196;
	input G197;
	input G198;
	input G199;
	input G200;
	input G201;
	input G202;
	input G203;
	input G204;
	input G205;
	input G206;
	input G207;
	input G208;
	input G209;
	input G210;
	input G211;
	input G212;
	input G213;
	input G214;
	input G215;
	input G216;
	input G217;
	input G218;
	input G219;
	input G220;
	input G221;
	input G222;
	input G223;
	input G224;
	input G225;
	input G226;
	input G227;
	input G228;
	input G229;
	input G230;
	input G231;
	input G232;
	input G233;
	input G234;
	input G235;
	input G236;
	input G237;
	input G238;
	input G239;
	input G240;
	input G339;
	input G1197;
	input G1455;
	input G1459;
	input G1462;
	input G1469;
	input G1480;
	input G1486;
	input G1492;
	input G1496;
	input G2204;
	input G2208;
	input G2211;
	input G2218;
	input G2224;
	input G2230;
	input G2236;
	input G2239;
	input G2247;
	input G2253;
	input G2256;
	input G3698;
	input G3701;
	input G3705;
	input G3711;
	input G3717;
	input G3723;
	input G3729;
	input G3737;
	input G3743;
	input G3749;
	input G4393;
	input G4394;
	input G4400;
	input G4405;
	input G4410;
	input G4415;
	input G4420;
	input G4427;
	input G4432;
	input G4437;
	input G4526;
	input G4528;
	output G2;
	output G3;
	output G450;
	output G448;
	output G444;
	output G442;
	output G440;
	output G438;
	output G496;
	output G494;
	output G492;
	output G490;
	output G488;
	output G486;
	output G484;
	output G482;
	output G480;
	output G560;
	output G542;
	output G558;
	output G556;
	output G554;
	output G552;
	output G550;
	output G548;
	output G546;
	output G544;
	output G540;
	output G538;
	output G536;
	output G534;
	output G532;
	output G530;
	output G528;
	output G526;
	output G524;
	output G279;
	output G436;
	output G478;
	output G522;
	output G402;
	output G404;
	output G406;
	output G408;
	output G410;
	output G432;
	output G446;
	output G284;
	output G286;
	output G289;
	output G292;
	output G341;
	output G281;
	output G453;
	output G278;
	output G373;
	output G246;
	output G258;
	output G264;
	output G270;
	output G388;
	output G391;
	output G394;
	output G397;
	output G376;
	output G379;
	output G382;
	output G385;
	output G412;
	output G414;
	output G416;
	output G249;
	output G295;
	output G324;
	output G252;
	output G276;
	output G310;
	output G313;
	output G316;
	output G319;
	output G327;
	output G330;
	output G333;
	output G336;
	output G418;
	output G273;
	output G298;
	output G301;
	output G304;
	output G307;
	output G344;
	output G422;
	output G469;
	output G419;
	output G471;
	output G359;
	output G362;
	output G365;
	output G368;
	output G347;
	output G350;
	output G353;
	output G356;
	output G321;
	output G338;
	output G370;
	output G399;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n347;
	wire n348;
	wire n349;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1102;
	wire n1103;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1356;
	wire n1357;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1384;
	wire n1385;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1399;
	wire n1400;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1413;
	wire n1414;
	wire n1416;
	wire n1417;
	wire n1419;
	wire n1421;
	wire n1423;
	wire n1424;
	wire n1426;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[2:0] w_G5_0;
	wire[1:0] w_G5_1;
	wire[2:0] w_G15_0;
	wire[2:0] w_G18_0;
	wire[2:0] w_G18_1;
	wire[2:0] w_G18_2;
	wire[2:0] w_G18_3;
	wire[2:0] w_G18_4;
	wire[2:0] w_G18_5;
	wire[2:0] w_G18_6;
	wire[2:0] w_G18_7;
	wire[2:0] w_G18_8;
	wire[2:0] w_G18_9;
	wire[2:0] w_G18_10;
	wire[2:0] w_G18_11;
	wire[2:0] w_G18_12;
	wire[2:0] w_G18_13;
	wire[2:0] w_G18_14;
	wire[2:0] w_G18_15;
	wire[2:0] w_G18_16;
	wire[2:0] w_G18_17;
	wire[2:0] w_G18_18;
	wire[2:0] w_G18_19;
	wire[2:0] w_G18_20;
	wire[2:0] w_G18_21;
	wire[2:0] w_G18_22;
	wire[2:0] w_G18_23;
	wire[2:0] w_G18_24;
	wire[2:0] w_G18_25;
	wire[2:0] w_G18_26;
	wire[2:0] w_G18_27;
	wire[2:0] w_G18_28;
	wire[2:0] w_G18_29;
	wire[2:0] w_G18_30;
	wire[2:0] w_G18_31;
	wire[2:0] w_G18_32;
	wire[2:0] w_G18_33;
	wire[2:0] w_G18_34;
	wire[2:0] w_G18_35;
	wire[2:0] w_G18_36;
	wire[2:0] w_G18_37;
	wire[2:0] w_G18_38;
	wire[2:0] w_G18_39;
	wire[2:0] w_G18_40;
	wire[2:0] w_G18_41;
	wire[2:0] w_G18_42;
	wire[2:0] w_G18_43;
	wire[2:0] w_G18_44;
	wire[2:0] w_G18_45;
	wire[2:0] w_G18_46;
	wire[2:0] w_G18_47;
	wire[2:0] w_G18_48;
	wire[2:0] w_G18_49;
	wire[1:0] w_G29_0;
	wire[2:0] w_G38_0;
	wire[2:0] w_G38_1;
	wire[2:0] w_G38_2;
	wire[1:0] w_G41_0;
	wire[1:0] w_G70_0;
	wire[1:0] w_G89_0;
	wire[2:0] w_G106_0;
	wire[1:0] w_G106_1;
	wire[1:0] w_G209_0;
	wire[1:0] w_G238_0;
	wire[2:0] w_G1455_0;
	wire[1:0] w_G1459_0;
	wire[1:0] w_G1462_0;
	wire[1:0] w_G1469_0;
	wire[2:0] w_G1480_0;
	wire[1:0] w_G1486_0;
	wire[2:0] w_G1492_0;
	wire[1:0] w_G1492_1;
	wire[2:0] w_G1496_0;
	wire[1:0] w_G1496_1;
	wire[2:0] w_G2204_0;
	wire[1:0] w_G2208_0;
	wire[2:0] w_G2211_0;
	wire[2:0] w_G2218_0;
	wire[2:0] w_G2224_0;
	wire[1:0] w_G2224_1;
	wire[2:0] w_G2230_0;
	wire[2:0] w_G2236_0;
	wire[2:0] w_G2239_0;
	wire[1:0] w_G2239_1;
	wire[2:0] w_G2247_0;
	wire[2:0] w_G2253_0;
	wire[1:0] w_G2256_0;
	wire[1:0] w_G3698_0;
	wire[2:0] w_G3701_0;
	wire[1:0] w_G3701_1;
	wire[2:0] w_G3705_0;
	wire[2:0] w_G3705_1;
	wire[1:0] w_G3711_0;
	wire[2:0] w_G3717_0;
	wire[2:0] w_G3723_0;
	wire[2:0] w_G3729_0;
	wire[1:0] w_G3729_1;
	wire[2:0] w_G3737_0;
	wire[2:0] w_G3743_0;
	wire[2:0] w_G3749_0;
	wire[1:0] w_G4393_0;
	wire[2:0] w_G4394_0;
	wire[1:0] w_G4394_1;
	wire[2:0] w_G4400_0;
	wire[1:0] w_G4400_1;
	wire[2:0] w_G4405_0;
	wire[1:0] w_G4405_1;
	wire[2:0] w_G4410_0;
	wire[2:0] w_G4415_0;
	wire[1:0] w_G4415_1;
	wire[2:0] w_G4420_0;
	wire[1:0] w_G4420_1;
	wire[2:0] w_G4427_0;
	wire[2:0] w_G4432_0;
	wire[2:0] w_G4437_0;
	wire[2:0] w_G4526_0;
	wire[2:0] w_G4526_1;
	wire[2:0] w_G4526_2;
	wire[2:0] w_G4528_0;
	wire w_G404_0;
	wire G404_fa_;
	wire w_G406_0;
	wire G406_fa_;
	wire w_G408_0;
	wire G408_fa_;
	wire w_G410_0;
	wire G410_fa_;
	wire w_G412_0;
	wire G412_fa_;
	wire w_G414_0;
	wire G414_fa_;
	wire w_G416_0;
	wire G416_fa_;
	wire w_G252_0;
	wire G252_fa_;
	wire[1:0] w_n345_0;
	wire[1:0] w_n347_0;
	wire[1:0] w_n349_0;
	wire[1:0] w_n353_0;
	wire[2:0] w_n354_0;
	wire[2:0] w_n355_0;
	wire[2:0] w_n355_1;
	wire[2:0] w_n355_2;
	wire[2:0] w_n355_3;
	wire[2:0] w_n355_4;
	wire[2:0] w_n355_5;
	wire[2:0] w_n355_6;
	wire[2:0] w_n355_7;
	wire[2:0] w_n355_8;
	wire[2:0] w_n355_9;
	wire[2:0] w_n355_10;
	wire[2:0] w_n355_11;
	wire[2:0] w_n355_12;
	wire[2:0] w_n355_13;
	wire[2:0] w_n355_14;
	wire[2:0] w_n355_15;
	wire[2:0] w_n355_16;
	wire[2:0] w_n355_17;
	wire[2:0] w_n355_18;
	wire[2:0] w_n355_19;
	wire[2:0] w_n355_20;
	wire[2:0] w_n355_21;
	wire[2:0] w_n355_22;
	wire[2:0] w_n355_23;
	wire[2:0] w_n355_24;
	wire[2:0] w_n355_25;
	wire[2:0] w_n355_26;
	wire[2:0] w_n355_27;
	wire[2:0] w_n355_28;
	wire[2:0] w_n355_29;
	wire[2:0] w_n355_30;
	wire[2:0] w_n355_31;
	wire[2:0] w_n355_32;
	wire[2:0] w_n355_33;
	wire[2:0] w_n355_34;
	wire[2:0] w_n355_35;
	wire[1:0] w_n357_0;
	wire[1:0] w_n358_0;
	wire[2:0] w_n359_0;
	wire[1:0] w_n359_1;
	wire[2:0] w_n361_0;
	wire[2:0] w_n362_0;
	wire[2:0] w_n363_0;
	wire[2:0] w_n364_0;
	wire[2:0] w_n366_0;
	wire[1:0] w_n367_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n369_0;
	wire[2:0] w_n370_0;
	wire[2:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[2:0] w_n373_0;
	wire[2:0] w_n373_1;
	wire[2:0] w_n373_2;
	wire[2:0] w_n373_3;
	wire[2:0] w_n373_4;
	wire[2:0] w_n373_5;
	wire[2:0] w_n373_6;
	wire[2:0] w_n373_7;
	wire[2:0] w_n373_8;
	wire[2:0] w_n373_9;
	wire[1:0] w_n374_0;
	wire[2:0] w_n375_0;
	wire[2:0] w_n377_0;
	wire[2:0] w_n377_1;
	wire[1:0] w_n378_0;
	wire[2:0] w_n379_0;
	wire[1:0] w_n380_0;
	wire[2:0] w_n383_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[1:0] w_n387_1;
	wire[2:0] w_n388_0;
	wire[2:0] w_n388_1;
	wire[2:0] w_n389_0;
	wire[1:0] w_n389_1;
	wire[2:0] w_n391_0;
	wire[2:0] w_n392_0;
	wire[2:0] w_n393_0;
	wire[1:0] w_n393_1;
	wire[1:0] w_n394_0;
	wire[2:0] w_n395_0;
	wire[1:0] w_n395_1;
	wire[2:0] w_n396_0;
	wire[2:0] w_n396_1;
	wire[1:0] w_n397_0;
	wire[2:0] w_n405_0;
	wire[1:0] w_n407_0;
	wire[2:0] w_n409_0;
	wire[1:0] w_n409_1;
	wire[2:0] w_n411_0;
	wire[1:0] w_n411_1;
	wire[2:0] w_n413_0;
	wire[1:0] w_n413_1;
	wire[2:0] w_n414_0;
	wire[1:0] w_n414_1;
	wire[1:0] w_n415_0;
	wire[2:0] w_n416_0;
	wire[1:0] w_n418_0;
	wire[1:0] w_n419_0;
	wire[1:0] w_n420_0;
	wire[2:0] w_n421_0;
	wire[1:0] w_n422_0;
	wire[2:0] w_n423_0;
	wire[1:0] w_n424_0;
	wire[2:0] w_n425_0;
	wire[1:0] w_n425_1;
	wire[2:0] w_n426_0;
	wire[1:0] w_n427_0;
	wire[2:0] w_n428_0;
	wire[2:0] w_n429_0;
	wire[1:0] w_n430_0;
	wire[1:0] w_n431_0;
	wire[2:0] w_n432_0;
	wire[2:0] w_n433_0;
	wire[2:0] w_n433_1;
	wire[1:0] w_n434_0;
	wire[1:0] w_n435_0;
	wire[2:0] w_n436_0;
	wire[2:0] w_n437_0;
	wire[1:0] w_n438_0;
	wire[1:0] w_n440_0;
	wire[2:0] w_n444_0;
	wire[2:0] w_n445_0;
	wire[2:0] w_n447_0;
	wire[2:0] w_n449_0;
	wire[1:0] w_n449_1;
	wire[2:0] w_n450_0;
	wire[2:0] w_n451_0;
	wire[2:0] w_n453_0;
	wire[1:0] w_n453_1;
	wire[2:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[2:0] w_n459_0;
	wire[2:0] w_n460_0;
	wire[2:0] w_n460_1;
	wire[2:0] w_n462_0;
	wire[2:0] w_n463_0;
	wire[1:0] w_n463_1;
	wire[2:0] w_n464_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n466_0;
	wire[1:0] w_n467_0;
	wire[2:0] w_n469_0;
	wire[1:0] w_n469_1;
	wire[2:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[1:0] w_n472_0;
	wire[2:0] w_n474_0;
	wire[2:0] w_n475_0;
	wire[2:0] w_n476_0;
	wire[1:0] w_n477_0;
	wire[2:0] w_n479_0;
	wire[1:0] w_n479_1;
	wire[2:0] w_n480_0;
	wire[1:0] w_n480_1;
	wire[1:0] w_n481_0;
	wire[1:0] w_n485_0;
	wire[1:0] w_n486_0;
	wire[2:0] w_n487_0;
	wire[2:0] w_n489_0;
	wire[2:0] w_n491_0;
	wire[1:0] w_n491_1;
	wire[2:0] w_n495_0;
	wire[1:0] w_n495_1;
	wire[2:0] w_n496_0;
	wire[2:0] w_n497_0;
	wire[1:0] w_n497_1;
	wire[1:0] w_n499_0;
	wire[1:0] w_n500_0;
	wire[2:0] w_n501_0;
	wire[1:0] w_n503_0;
	wire[2:0] w_n504_0;
	wire[1:0] w_n504_1;
	wire[1:0] w_n505_0;
	wire[1:0] w_n507_0;
	wire[2:0] w_n509_0;
	wire[1:0] w_n511_0;
	wire[2:0] w_n512_0;
	wire[2:0] w_n513_0;
	wire[1:0] w_n513_1;
	wire[1:0] w_n514_0;
	wire[1:0] w_n516_0;
	wire[2:0] w_n517_0;
	wire[1:0] w_n517_1;
	wire[2:0] w_n518_0;
	wire[2:0] w_n518_1;
	wire[1:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[2:0] w_n524_0;
	wire[2:0] w_n524_1;
	wire[2:0] w_n526_0;
	wire[1:0] w_n528_0;
	wire[1:0] w_n530_0;
	wire[2:0] w_n531_0;
	wire[1:0] w_n531_1;
	wire[2:0] w_n536_0;
	wire[1:0] w_n538_0;
	wire[2:0] w_n539_0;
	wire[1:0] w_n539_1;
	wire[1:0] w_n544_0;
	wire[1:0] w_n546_0;
	wire[2:0] w_n547_0;
	wire[1:0] w_n547_1;
	wire[1:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n552_0;
	wire[1:0] w_n554_0;
	wire[2:0] w_n555_0;
	wire[1:0] w_n555_1;
	wire[2:0] w_n556_0;
	wire[1:0] w_n558_0;
	wire[1:0] w_n560_0;
	wire[1:0] w_n562_0;
	wire[2:0] w_n563_0;
	wire[1:0] w_n563_1;
	wire[2:0] w_n564_0;
	wire[1:0] w_n565_0;
	wire[2:0] w_n566_0;
	wire[2:0] w_n568_0;
	wire[2:0] w_n570_0;
	wire[2:0] w_n570_1;
	wire[2:0] w_n572_0;
	wire[1:0] w_n572_1;
	wire[2:0] w_n573_0;
	wire[1:0] w_n573_1;
	wire[2:0] w_n574_0;
	wire[2:0] w_n575_0;
	wire[1:0] w_n575_1;
	wire[2:0] w_n576_0;
	wire[1:0] w_n577_0;
	wire[2:0] w_n578_0;
	wire[2:0] w_n580_0;
	wire[2:0] w_n581_0;
	wire[2:0] w_n582_0;
	wire[1:0] w_n584_0;
	wire[2:0] w_n585_0;
	wire[1:0] w_n585_1;
	wire[2:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[2:0] w_n590_0;
	wire[1:0] w_n592_0;
	wire[2:0] w_n593_0;
	wire[1:0] w_n593_1;
	wire[2:0] w_n594_0;
	wire[2:0] w_n595_0;
	wire[1:0] w_n597_0;
	wire[2:0] w_n598_0;
	wire[1:0] w_n598_1;
	wire[2:0] w_n599_0;
	wire[1:0] w_n600_0;
	wire[1:0] w_n602_0;
	wire[2:0] w_n603_0;
	wire[1:0] w_n603_1;
	wire[1:0] w_n604_0;
	wire[2:0] w_n605_0;
	wire[1:0] w_n609_0;
	wire[1:0] w_n610_0;
	wire[1:0] w_n612_0;
	wire[2:0] w_n613_0;
	wire[2:0] w_n615_0;
	wire[1:0] w_n616_0;
	wire[2:0] w_n618_0;
	wire[2:0] w_n619_0;
	wire[2:0] w_n622_0;
	wire[1:0] w_n624_0;
	wire[2:0] w_n625_0;
	wire[1:0] w_n625_1;
	wire[2:0] w_n626_0;
	wire[1:0] w_n626_1;
	wire[2:0] w_n627_0;
	wire[1:0] w_n629_0;
	wire[2:0] w_n630_0;
	wire[2:0] w_n631_0;
	wire[2:0] w_n632_0;
	wire[1:0] w_n632_1;
	wire[1:0] w_n634_0;
	wire[2:0] w_n635_0;
	wire[1:0] w_n635_1;
	wire[2:0] w_n636_0;
	wire[2:0] w_n641_0;
	wire[2:0] w_n642_0;
	wire[1:0] w_n644_0;
	wire[1:0] w_n645_0;
	wire[1:0] w_n646_0;
	wire[1:0] w_n647_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n651_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n653_0;
	wire[2:0] w_n654_0;
	wire[1:0] w_n655_0;
	wire[1:0] w_n656_0;
	wire[2:0] w_n657_0;
	wire[1:0] w_n659_0;
	wire[2:0] w_n660_0;
	wire[2:0] w_n661_0;
	wire[1:0] w_n662_0;
	wire[2:0] w_n663_0;
	wire[1:0] w_n663_1;
	wire[1:0] w_n664_0;
	wire[1:0] w_n666_0;
	wire[1:0] w_n669_0;
	wire[1:0] w_n671_0;
	wire[2:0] w_n673_0;
	wire[1:0] w_n674_0;
	wire[2:0] w_n676_0;
	wire[1:0] w_n678_0;
	wire[2:0] w_n680_0;
	wire[2:0] w_n680_1;
	wire[2:0] w_n680_2;
	wire[1:0] w_n682_0;
	wire[1:0] w_n683_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[1:0] w_n695_0;
	wire[1:0] w_n696_0;
	wire[1:0] w_n698_0;
	wire[2:0] w_n700_0;
	wire[1:0] w_n700_1;
	wire[2:0] w_n703_0;
	wire[2:0] w_n703_1;
	wire[1:0] w_n705_0;
	wire[2:0] w_n707_0;
	wire[2:0] w_n707_1;
	wire[2:0] w_n709_0;
	wire[1:0] w_n709_1;
	wire[2:0] w_n711_0;
	wire[1:0] w_n711_1;
	wire[2:0] w_n712_0;
	wire[1:0] w_n713_0;
	wire[2:0] w_n715_0;
	wire[1:0] w_n715_1;
	wire[2:0] w_n718_0;
	wire[1:0] w_n719_0;
	wire[2:0] w_n720_0;
	wire[2:0] w_n723_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n725_0;
	wire[2:0] w_n726_0;
	wire[1:0] w_n726_1;
	wire[2:0] w_n729_0;
	wire[1:0] w_n729_1;
	wire[2:0] w_n734_0;
	wire[1:0] w_n736_0;
	wire[2:0] w_n737_0;
	wire[1:0] w_n737_1;
	wire[2:0] w_n741_0;
	wire[1:0] w_n741_1;
	wire[1:0] w_n743_0;
	wire[2:0] w_n744_0;
	wire[2:0] w_n747_0;
	wire[1:0] w_n749_0;
	wire[1:0] w_n754_0;
	wire[2:0] w_n755_0;
	wire[1:0] w_n755_1;
	wire[2:0] w_n758_0;
	wire[1:0] w_n758_1;
	wire[1:0] w_n760_0;
	wire[2:0] w_n761_0;
	wire[2:0] w_n764_0;
	wire[1:0] w_n766_0;
	wire[1:0] w_n767_0;
	wire[2:0] w_n768_0;
	wire[2:0] w_n772_0;
	wire[1:0] w_n773_0;
	wire[1:0] w_n774_0;
	wire[1:0] w_n775_0;
	wire[2:0] w_n776_0;
	wire[2:0] w_n780_0;
	wire[1:0] w_n781_0;
	wire[2:0] w_n796_0;
	wire[1:0] w_n796_1;
	wire[2:0] w_n800_0;
	wire[1:0] w_n800_1;
	wire[2:0] w_n803_0;
	wire[2:0] w_n806_0;
	wire[1:0] w_n808_0;
	wire[2:0] w_n810_0;
	wire[1:0] w_n810_1;
	wire[2:0] w_n814_0;
	wire[1:0] w_n814_1;
	wire[2:0] w_n817_0;
	wire[2:0] w_n820_0;
	wire[1:0] w_n822_0;
	wire[2:0] w_n824_0;
	wire[2:0] w_n827_0;
	wire[2:0] w_n845_0;
	wire[1:0] w_n845_1;
	wire[2:0] w_n848_0;
	wire[1:0] w_n848_1;
	wire[2:0] w_n851_0;
	wire[2:0] w_n854_0;
	wire[1:0] w_n856_0;
	wire[2:0] w_n858_0;
	wire[2:0] w_n862_0;
	wire[1:0] w_n863_0;
	wire[1:0] w_n864_0;
	wire[2:0] w_n866_0;
	wire[2:0] w_n870_0;
	wire[1:0] w_n871_0;
	wire[2:0] w_n885_0;
	wire[2:0] w_n888_0;
	wire[2:0] w_n891_0;
	wire[2:0] w_n894_0;
	wire[1:0] w_n895_0;
	wire[2:0] w_n900_0;
	wire[2:0] w_n903_0;
	wire[1:0] w_n905_0;
	wire[2:0] w_n916_0;
	wire[2:0] w_n919_0;
	wire[2:0] w_n926_0;
	wire[2:0] w_n930_0;
	wire[2:0] w_n935_0;
	wire[2:0] w_n938_0;
	wire[2:0] w_n944_0;
	wire[2:0] w_n947_0;
	wire[2:0] w_n950_0;
	wire[1:0] w_n950_1;
	wire[2:0] w_n953_0;
	wire[1:0] w_n953_1;
	wire[2:0] w_n966_0;
	wire[2:0] w_n970_0;
	wire[2:0] w_n973_0;
	wire[1:0] w_n973_1;
	wire[2:0] w_n977_0;
	wire[1:0] w_n977_1;
	wire[2:0] w_n980_0;
	wire[2:0] w_n983_0;
	wire[1:0] w_n985_0;
	wire[2:0] w_n987_0;
	wire[2:0] w_n991_0;
	wire[1:0] w_n992_0;
	wire[2:0] w_n995_0;
	wire[2:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1042_0;
	wire[2:0] w_n1059_0;
	wire[2:0] w_n1067_0;
	wire[2:0] w_n1069_0;
	wire[1:0] w_n1070_0;
	wire[1:0] w_n1073_0;
	wire[1:0] w_n1078_0;
	wire[2:0] w_n1084_0;
	wire[1:0] w_n1086_0;
	wire[1:0] w_n1090_0;
	wire[2:0] w_n1092_0;
	wire[2:0] w_n1094_0;
	wire[1:0] w_n1096_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1105_0;
	wire[1:0] w_n1106_0;
	wire[1:0] w_n1108_0;
	wire[1:0] w_n1113_0;
	wire[1:0] w_n1118_0;
	wire[1:0] w_n1127_0;
	wire[1:0] w_n1137_0;
	wire[1:0] w_n1150_0;
	wire[1:0] w_n1172_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1308_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1310_0;
	wire[2:0] w_n1312_0;
	wire[1:0] w_n1312_1;
	wire[1:0] w_n1316_0;
	wire[1:0] w_n1317_0;
	wire[2:0] w_n1321_0;
	wire[1:0] w_n1321_1;
	wire[1:0] w_n1323_0;
	wire[1:0] w_n1333_0;
	wire[2:0] w_n1337_0;
	wire[1:0] w_n1337_1;
	wire[2:0] w_n1340_0;
	wire[1:0] w_n1343_0;
	wire[1:0] w_n1344_0;
	wire[1:0] w_n1359_0;
	wire[1:0] w_n1364_0;
	wire[1:0] w_n1369_0;
	wire[1:0] w_n1370_0;
	wire[1:0] w_n1372_0;
	wire[1:0] w_n1387_0;
	wire[1:0] w_n1388_0;
	wire[1:0] w_n1396_0;
	wire[1:0] w_n1402_0;
	wire[1:0] w_n1408_0;
	wire[1:0] w_n1419_0;
	wire[1:0] w_n1426_0;
	wire[1:0] w_n1431_0;
	wire[1:0] w_n1433_0;
	wire[1:0] w_n1440_0;
	wire[2:0] w_n1452_0;
	wire[1:0] w_n1458_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1492_0;
	wire[1:0] w_n1506_0;
	wire[1:0] w_n1511_0;
	wire[1:0] w_n1518_0;
	wire[1:0] w_n1529_0;
	wire[1:0] w_n1531_0;
	wire[1:0] w_n1534_0;
	wire[1:0] w_n1536_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1554_0;
	wire[2:0] w_n1562_0;
	wire[1:0] w_n1587_0;
	wire[1:0] w_n1597_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1620_0;
	wire[1:0] w_n1624_0;
	wire w_dff_A_neoobXwD1_0;
	wire w_dff_B_dY68LMNi2_2;
	wire w_dff_B_c1VlsQ6b8_1;
	wire w_dff_B_LG1bYm0e9_1;
	wire w_dff_B_RPUVOxCn0_1;
	wire w_dff_B_TKq0mV5z9_1;
	wire w_dff_B_GqewLBi55_1;
	wire w_dff_B_GMI6467M9_1;
	wire w_dff_B_aAztm4hS6_1;
	wire w_dff_B_aQ5P1FDE8_1;
	wire w_dff_B_7qGpVZ1P4_1;
	wire w_dff_B_DEDLvIgL1_1;
	wire w_dff_B_I3uFP1fQ7_1;
	wire w_dff_B_NLE5NhC27_1;
	wire w_dff_B_vjfIi28Z3_1;
	wire w_dff_B_ZngyyZX71_1;
	wire w_dff_B_yodZqdA21_1;
	wire w_dff_B_rOvy3G2j8_1;
	wire w_dff_B_NI6Dgyqd3_1;
	wire w_dff_B_B6UBMEla4_1;
	wire w_dff_B_OsxWh6Gu4_0;
	wire w_dff_B_uAtrPtaT2_0;
	wire w_dff_B_CwMfwXe77_0;
	wire w_dff_B_vazfz53v6_0;
	wire w_dff_B_ZAryOtFP5_0;
	wire w_dff_B_0AWBxpFH7_0;
	wire w_dff_B_yoCuqTVD0_0;
	wire w_dff_B_8cVb4XS05_0;
	wire w_dff_B_qEBw09743_0;
	wire w_dff_B_UeaNXdH80_0;
	wire w_dff_B_2yWoyz8V1_0;
	wire w_dff_B_S7gC4XIz8_0;
	wire w_dff_B_iJsdmYZJ1_0;
	wire w_dff_B_yUS5D9F94_0;
	wire w_dff_B_HJqdpYuJ8_0;
	wire w_dff_B_POG4d9VZ1_0;
	wire w_dff_B_FddPjT129_0;
	wire w_dff_B_uJkImova9_0;
	wire w_dff_B_3Y8BuPAf9_0;
	wire w_dff_B_23I2t5e54_0;
	wire w_dff_B_u6M0AzWb0_0;
	wire w_dff_B_OhpzQVtd6_0;
	wire w_dff_B_ghqpiIah2_0;
	wire w_dff_B_5MmDMCKW7_0;
	wire w_dff_B_tVWczIsZ9_0;
	wire w_dff_B_BjwpQMHQ1_0;
	wire w_dff_B_ULDO8dqB2_0;
	wire w_dff_B_QlrdZJQH0_0;
	wire w_dff_B_IsgJckqP0_0;
	wire w_dff_B_eT6QaDVn0_0;
	wire w_dff_B_t0U6Pf0O4_0;
	wire w_dff_B_Dj7mkZ3I9_0;
	wire w_dff_B_T1d6BPOm2_0;
	wire w_dff_B_7M1lrMPW2_1;
	wire w_dff_B_XoG7i2o52_1;
	wire w_dff_B_3CM2afkW3_1;
	wire w_dff_B_5k0i0PCj5_1;
	wire w_dff_B_1RSpuAkh5_1;
	wire w_dff_B_vAg6SD5U8_1;
	wire w_dff_B_uD668HLK9_1;
	wire w_dff_B_GZuxk9lo6_1;
	wire w_dff_B_maC7SitY5_1;
	wire w_dff_B_SvJAykEn0_1;
	wire w_dff_B_WbhBj9pS6_1;
	wire w_dff_B_wEDlNkBH6_1;
	wire w_dff_B_RNc4U37m0_1;
	wire w_dff_B_brHvYuwj6_1;
	wire w_dff_B_u3oP7Dlo2_1;
	wire w_dff_B_6Us1o1PU5_1;
	wire w_dff_B_UA13COXH6_1;
	wire w_dff_B_BvbgFEcY5_1;
	wire w_dff_B_AlcbGVrj8_1;
	wire w_dff_B_vlmifdGp3_1;
	wire w_dff_B_91Pq6RVV2_1;
	wire w_dff_B_ifa296Kc3_1;
	wire w_dff_B_V1hcwmJH1_1;
	wire w_dff_B_Uqfl6Yaz1_1;
	wire w_dff_B_04WncmoK4_1;
	wire w_dff_B_qe1whFNV3_1;
	wire w_dff_B_hRWrvexO9_1;
	wire w_dff_B_gKcrzpjS8_1;
	wire w_dff_B_bWMxfGkw0_1;
	wire w_dff_B_NMFhvr9m9_1;
	wire w_dff_B_B2hLuiYn0_0;
	wire w_dff_B_38oiTr2l5_0;
	wire w_dff_B_uYbsBXlK2_0;
	wire w_dff_B_Zjqf0u0m4_0;
	wire w_dff_B_dyinEq376_0;
	wire w_dff_B_Wc4Ludv69_0;
	wire w_dff_B_zWrP37Rb6_0;
	wire w_dff_B_JH8UfnCm6_0;
	wire w_dff_B_l9PVMqNj6_0;
	wire w_dff_B_v02053He5_0;
	wire w_dff_B_paAqqfnL4_0;
	wire w_dff_B_QbAVlX530_0;
	wire w_dff_B_9VwHz3EU6_0;
	wire w_dff_B_y53gdfjG8_0;
	wire w_dff_B_7q9fuPJQ6_0;
	wire w_dff_B_9GcvIL8U1_0;
	wire w_dff_B_Gw1dYDfT7_1;
	wire w_dff_B_WKEClvuR0_1;
	wire w_dff_B_4Yixfr1f1_1;
	wire w_dff_B_Tax8CM1w1_1;
	wire w_dff_B_phUmAw6k9_1;
	wire w_dff_B_I5HoOQ6y8_1;
	wire w_dff_B_wcs81AfL4_1;
	wire w_dff_B_62W8pPqa8_1;
	wire w_dff_B_ZosEPnXn3_1;
	wire w_dff_B_FiXAGPcI3_1;
	wire w_dff_B_ZTSxbjnP1_1;
	wire w_dff_B_Bin7Hwuy9_1;
	wire w_dff_B_PYjbCfre1_1;
	wire w_dff_B_UPvoHW9n9_1;
	wire w_dff_B_UNZmtkoq5_1;
	wire w_dff_B_FF0x16jo9_1;
	wire w_dff_B_UDiyE8Cg4_1;
	wire w_dff_B_wQJCt7bC5_1;
	wire w_dff_B_EqioovOn5_1;
	wire w_dff_B_6PwXRHKg5_1;
	wire w_dff_B_tDZlnk9p1_1;
	wire w_dff_B_GV18tMPh4_1;
	wire w_dff_B_h38f78Fw0_1;
	wire w_dff_B_VeT2Yyaa5_1;
	wire w_dff_B_A5DwHN7y8_0;
	wire w_dff_B_gO0NL7DJ3_0;
	wire w_dff_B_Gf7KTZyb2_0;
	wire w_dff_B_IJO2BKKF0_0;
	wire w_dff_B_yFUpbVr59_0;
	wire w_dff_B_UqU1vpSG3_0;
	wire w_dff_B_3bY84fzm8_0;
	wire w_dff_B_BNtIyLIC8_0;
	wire w_dff_B_a6HOVMNp5_0;
	wire w_dff_B_VgNxVw340_0;
	wire w_dff_B_9dMiWYt69_0;
	wire w_dff_B_QbEwMlUz9_0;
	wire w_dff_B_CRsm53By6_0;
	wire w_dff_B_8loWY7PT9_0;
	wire w_dff_B_JuK41xEe3_3;
	wire w_dff_B_93SjQFsm5_3;
	wire w_dff_B_ie39DiEx3_3;
	wire w_dff_B_hpYgyyl18_3;
	wire w_dff_B_jMxuNleY0_3;
	wire w_dff_B_oXzYyErQ1_3;
	wire w_dff_B_xX8YJHkx6_3;
	wire w_dff_B_utu1s2SQ7_3;
	wire w_dff_B_7JPvDrLT9_3;
	wire w_dff_B_CV1ibV4a3_3;
	wire w_dff_B_7UuL3FUV5_3;
	wire w_dff_B_FZ91vWJ72_3;
	wire w_dff_B_hh9fC2uG3_3;
	wire w_dff_B_60DsptNY9_3;
	wire w_dff_B_BRdw5yBj8_3;
	wire w_dff_B_zeJQSlSZ3_3;
	wire w_dff_B_IdW8oNTG6_3;
	wire w_dff_B_QyolK1dE4_3;
	wire w_dff_B_Efdvrtbe2_3;
	wire w_dff_B_MSPwtXEF2_3;
	wire w_dff_B_u7PRntmF6_3;
	wire w_dff_B_bMaMMfOB6_3;
	wire w_dff_B_NcsPgPvU4_3;
	wire w_dff_B_4D5BXUHe7_3;
	wire w_dff_B_HzBoAF1D8_1;
	wire w_dff_B_tVLtNIMF4_1;
	wire w_dff_B_GuxoXpB74_1;
	wire w_dff_B_DTjEKTEt3_1;
	wire w_dff_B_rbx1awGU1_1;
	wire w_dff_B_OY0MOmnh6_1;
	wire w_dff_B_irR47WqU3_1;
	wire w_dff_B_SG1bO3fH1_1;
	wire w_dff_B_pJBwPVHu5_1;
	wire w_dff_B_DBJ1bMFB5_1;
	wire w_dff_B_evg1RF3N0_1;
	wire w_dff_B_7RYcBoPU1_1;
	wire w_dff_B_zXpsqUdH6_1;
	wire w_dff_B_Zob7ArHT6_1;
	wire w_dff_B_wc2eYW0k9_1;
	wire w_dff_B_hXe5Qo5m7_1;
	wire w_dff_B_3xjDdytG7_1;
	wire w_dff_B_eNvZU7tn2_1;
	wire w_dff_B_fHdbwiZG9_1;
	wire w_dff_B_UnqY7FVK3_1;
	wire w_dff_B_UZf5VXFx7_1;
	wire w_dff_B_MmUI7ZMm7_1;
	wire w_dff_B_uZ192TCG0_1;
	wire w_dff_B_WDf4wCSn8_1;
	wire w_dff_B_RznskHIj2_1;
	wire w_dff_B_Q5HzTztO4_1;
	wire w_dff_B_goT78SRU6_1;
	wire w_dff_B_WC0X31Ys1_1;
	wire w_dff_B_rM25Xr037_1;
	wire w_dff_B_nd1DUFUd8_1;
	wire w_dff_B_cU5aMtv53_1;
	wire w_dff_B_rDIOLzwH7_1;
	wire w_dff_B_ynMNMAMO9_1;
	wire w_dff_B_uozBSSLV5_1;
	wire w_dff_B_uaVUETXI5_1;
	wire w_dff_B_qaGvqW4J3_1;
	wire w_dff_B_sCoF3rCx2_1;
	wire w_dff_B_sqslCrcV6_1;
	wire w_dff_B_A7GEn0iK2_1;
	wire w_dff_B_i4FjaiwR6_1;
	wire w_dff_B_uWiypTGG0_1;
	wire w_dff_B_4tcwl7ig6_1;
	wire w_dff_B_opKgIT7H5_1;
	wire w_dff_B_TKf0P0eY2_1;
	wire w_dff_B_NiEoq66h7_1;
	wire w_dff_B_JyJ9ZyIc9_1;
	wire w_dff_B_le3aFNwW9_1;
	wire w_dff_B_yUTq1RZm8_1;
	wire w_dff_B_iV9Ty4gF7_1;
	wire w_dff_B_bhGoLnJM2_1;
	wire w_dff_B_XB3WTDsk3_1;
	wire w_dff_B_SFv6DJjw4_1;
	wire w_dff_B_e6bgyifi9_1;
	wire w_dff_B_fkChAObi7_1;
	wire w_dff_B_3eFE7fLM2_1;
	wire w_dff_B_LLmxIlqS9_1;
	wire w_dff_B_IOPm2ZGa5_1;
	wire w_dff_B_zz5BSZhW8_1;
	wire w_dff_B_39kMFezJ5_1;
	wire w_dff_B_q6WIcda37_1;
	wire w_dff_B_lNrZNO0Q0_1;
	wire w_dff_B_Z0sU4nZ85_1;
	wire w_dff_B_SBI04YPO6_1;
	wire w_dff_B_rUoPHGzb6_1;
	wire w_dff_B_qKGOuUOs9_1;
	wire w_dff_B_x4CrNFNp6_1;
	wire w_dff_B_avQhiC6t0_1;
	wire w_dff_B_7GMzqdeq9_0;
	wire w_dff_B_uRYSEkUI5_0;
	wire w_dff_B_bDaFGUFH9_0;
	wire w_dff_B_juw7xejP3_0;
	wire w_dff_B_BRxNbwkm8_0;
	wire w_dff_B_agVygko66_0;
	wire w_dff_B_RIw1Ilxk0_0;
	wire w_dff_A_76k9SREw6_0;
	wire w_dff_B_pbqrQltl6_3;
	wire w_dff_B_PUqrvXMC6_3;
	wire w_dff_B_K7hFgk7U8_3;
	wire w_dff_B_svD7A4pO2_3;
	wire w_dff_B_8xOSwhQ07_3;
	wire w_dff_B_nCKFztNW0_3;
	wire w_dff_B_biXxT3gb4_3;
	wire w_dff_B_dbVi2Z9V8_3;
	wire w_dff_B_1zBBAgAi3_3;
	wire w_dff_B_39clW5ga6_3;
	wire w_dff_B_ZkwrlPoR3_3;
	wire w_dff_B_NkFpvgDM0_3;
	wire w_dff_B_jpeCzUAy0_3;
	wire w_dff_B_MnmvRxqQ5_3;
	wire w_dff_B_DgBTPy9R6_3;
	wire w_dff_B_mRi94PP12_3;
	wire w_dff_B_QGxmCFnk2_3;
	wire w_dff_B_PDPdz2Yp4_3;
	wire w_dff_B_aLRc7sFK3_3;
	wire w_dff_B_hOhvEjaL4_3;
	wire w_dff_B_9w6MseZu9_3;
	wire w_dff_B_2xFQEemQ3_3;
	wire w_dff_B_YRuhaPUY8_3;
	wire w_dff_B_tXSifjvS6_3;
	wire w_dff_B_T6SfYfZx3_3;
	wire w_dff_B_S6FG1Isd3_3;
	wire w_dff_B_fv6XoOr35_3;
	wire w_dff_B_Ary4ZO6f5_3;
	wire w_dff_B_4LS7fqyE8_3;
	wire w_dff_B_dC65g0Go1_3;
	wire w_dff_B_VVFFn8WV7_3;
	wire w_dff_B_loIHxii74_3;
	wire w_dff_B_p6HvR6vZ2_3;
	wire w_dff_B_p1zgFYqg9_3;
	wire w_dff_B_7xfDQCrw4_0;
	wire w_dff_B_wJPTGXyJ2_0;
	wire w_dff_B_Ecfi3mhT0_0;
	wire w_dff_B_ilTnKteO2_1;
	wire w_dff_A_Dmc7a2bN2_1;
	wire w_dff_A_LLNBvJTM8_0;
	wire w_dff_A_GEvlkdsB5_0;
	wire w_dff_A_YaYzmZlX2_0;
	wire w_dff_A_FX0Iisaz5_0;
	wire w_dff_A_MIhcir4I6_0;
	wire w_dff_A_erFnwnth9_0;
	wire w_dff_A_bQzyhJSN6_0;
	wire w_dff_A_wLqUgbMr3_0;
	wire w_dff_A_uWI17KVJ3_0;
	wire w_dff_A_VB5iWxWM3_0;
	wire w_dff_A_zhbhsqta1_0;
	wire w_dff_A_gMEzPjoT8_0;
	wire w_dff_A_oAJOi9300_0;
	wire w_dff_A_FsicpojQ8_0;
	wire w_dff_A_mshP6Gmr6_0;
	wire w_dff_A_9ZwfPTf05_0;
	wire w_dff_A_N33t5uUQ4_0;
	wire w_dff_A_EbUD35wF7_0;
	wire w_dff_A_E3m7ZjeC2_0;
	wire w_dff_A_zVnf6q9a8_0;
	wire w_dff_A_Nq5hrONx9_0;
	wire w_dff_A_YqpFphdb8_0;
	wire w_dff_A_S5BJmosr8_0;
	wire w_dff_A_71RZnxKQ3_0;
	wire w_dff_A_6yMSafOb1_0;
	wire w_dff_A_jj6JeSgk7_0;
	wire w_dff_A_rGkCTCdA5_0;
	wire w_dff_A_hvCgOQpC5_0;
	wire w_dff_A_w7hDUjCD5_0;
	wire w_dff_A_TFlXIh2G6_0;
	wire w_dff_A_1n6ENcOU8_0;
	wire w_dff_A_6vJCtxEh0_0;
	wire w_dff_A_AUQvMz4w4_0;
	wire w_dff_A_ulmky10N1_0;
	wire w_dff_A_swuztbhy0_0;
	wire w_dff_A_v8D77aif1_0;
	wire w_dff_A_MzjyoJYC7_0;
	wire w_dff_A_LWM8mLPO1_0;
	wire w_dff_A_6v1KheBj0_1;
	wire w_dff_A_YY0xL0rk4_0;
	wire w_dff_A_3bF7dwZG0_0;
	wire w_dff_A_35PC5vQ83_0;
	wire w_dff_A_AJHmpnhH7_0;
	wire w_dff_A_CMwCjjRI2_0;
	wire w_dff_A_hqt01n107_0;
	wire w_dff_A_CnzwQmx13_0;
	wire w_dff_A_GN2WozW12_0;
	wire w_dff_A_sV4syeeH4_0;
	wire w_dff_A_jVx5KnoL8_0;
	wire w_dff_A_hCZEAIKm2_0;
	wire w_dff_A_ozKRS0Sp4_0;
	wire w_dff_A_QMaNV75Q3_0;
	wire w_dff_A_CqEIMk7e3_0;
	wire w_dff_A_9L2Rqvdx2_0;
	wire w_dff_A_XDt8ZnXd2_0;
	wire w_dff_A_MsXBp7Fd5_0;
	wire w_dff_A_Y12zr4vQ4_0;
	wire w_dff_A_YuVSPCiI7_0;
	wire w_dff_A_QTDWwmDk3_0;
	wire w_dff_A_6IZ5LgYS4_0;
	wire w_dff_A_8oR3DoJm0_0;
	wire w_dff_A_Nbl5VoIt6_0;
	wire w_dff_A_UY9cMqF68_0;
	wire w_dff_A_ybP7apAr7_0;
	wire w_dff_A_ovUm93dE4_0;
	wire w_dff_A_aayRUxMn9_0;
	wire w_dff_A_TzFmMYuV7_0;
	wire w_dff_A_yMHO25it0_0;
	wire w_dff_A_ED4QewEl8_0;
	wire w_dff_A_yCudmDL28_0;
	wire w_dff_A_MOmaS9wo9_0;
	wire w_dff_A_ZrhELOdn8_0;
	wire w_dff_A_JEg0rFPI8_0;
	wire w_dff_A_nsnh1dY66_0;
	wire w_dff_A_FMHQIao37_0;
	wire w_dff_A_5c5TmNXW1_0;
	wire w_dff_A_MkWXwYFV8_0;
	wire w_dff_A_P8WDRkB32_1;
	wire w_dff_A_KEHXtWQB4_0;
	wire w_dff_A_UJBNpKNU2_0;
	wire w_dff_A_CnjPptcQ8_0;
	wire w_dff_A_DJbw1rEN1_0;
	wire w_dff_A_vw3tfYfV2_0;
	wire w_dff_A_q63BVYZV5_0;
	wire w_dff_A_aTPQEO3a4_0;
	wire w_dff_A_6ZHdjy9k2_0;
	wire w_dff_A_s0xYhP2F4_0;
	wire w_dff_A_QZKpCIPp1_0;
	wire w_dff_A_jUL6YSMs4_0;
	wire w_dff_A_sFgDPNML0_0;
	wire w_dff_A_8kX9Yz7G6_0;
	wire w_dff_A_mcy3O4Vt9_0;
	wire w_dff_A_FoGZ3b4J6_0;
	wire w_dff_A_cqTPpmCQ6_0;
	wire w_dff_A_ys8UfOQC0_0;
	wire w_dff_A_k9OYpDMQ2_0;
	wire w_dff_A_7uDRE68t8_0;
	wire w_dff_A_qXWQFPdP2_0;
	wire w_dff_A_pwGBwSRd0_0;
	wire w_dff_A_oQ0QB7Ng0_0;
	wire w_dff_A_VU4g507v9_0;
	wire w_dff_A_Sn8GvQn42_0;
	wire w_dff_A_uKOB4OED5_0;
	wire w_dff_A_aYR3FIJa8_0;
	wire w_dff_A_6wknBOYK4_0;
	wire w_dff_A_8xsSwGYc3_0;
	wire w_dff_A_KTg2UkOS6_0;
	wire w_dff_A_1mGoiPaC2_0;
	wire w_dff_A_YNf3TYu26_0;
	wire w_dff_A_rR7wkgtB4_0;
	wire w_dff_A_R6k27Hmj9_0;
	wire w_dff_A_gANCoK860_0;
	wire w_dff_A_lLSRErtM9_0;
	wire w_dff_A_mSM3Ycj02_0;
	wire w_dff_A_0M3qaGI70_0;
	wire w_dff_A_dNfSPOfu6_0;
	wire w_dff_A_IflYUUBn6_1;
	wire w_dff_A_sRfM7A0E4_0;
	wire w_dff_A_MNfhiR7A3_0;
	wire w_dff_A_QkfOOnRg4_0;
	wire w_dff_A_g3qdOyMo7_0;
	wire w_dff_A_GAsH9soI5_0;
	wire w_dff_A_gJZmpSG89_0;
	wire w_dff_A_SfiU2wq33_0;
	wire w_dff_A_jMQZZB073_0;
	wire w_dff_A_rUdNl4IU4_0;
	wire w_dff_A_q7QZp0hU4_0;
	wire w_dff_A_k3Pyj5zi3_0;
	wire w_dff_A_GZjy3eqv4_0;
	wire w_dff_A_4ybbnZ511_0;
	wire w_dff_A_Lk4OfqAX8_0;
	wire w_dff_A_ceuXNrKz2_0;
	wire w_dff_A_Qla1hDku4_0;
	wire w_dff_A_qnhBl79k4_0;
	wire w_dff_A_H8FAlFuI8_0;
	wire w_dff_A_TMJ7B2sj0_0;
	wire w_dff_A_1E2AD5X72_0;
	wire w_dff_A_Yum01tnZ1_0;
	wire w_dff_A_riiZSMiM5_0;
	wire w_dff_A_Mo2MkYzG5_0;
	wire w_dff_A_uKon5cKx9_0;
	wire w_dff_A_2iCK4iSu6_0;
	wire w_dff_A_R7t4Bh989_0;
	wire w_dff_A_Me7Q28lX7_0;
	wire w_dff_A_g3Mop0g48_0;
	wire w_dff_A_sUHsZpr36_0;
	wire w_dff_A_loEuQvIp0_0;
	wire w_dff_A_2Di6GwsR7_0;
	wire w_dff_A_PZVXZ8I75_0;
	wire w_dff_A_SZ2yEkf29_0;
	wire w_dff_A_17KJYLmk1_0;
	wire w_dff_A_v9mhp5IQ1_0;
	wire w_dff_A_e2B9nFVc9_0;
	wire w_dff_A_eUhlLYI76_0;
	wire w_dff_A_F88TuU6w1_0;
	wire w_dff_A_U5TrYOk95_1;
	wire w_dff_A_Ha7yNAiw9_0;
	wire w_dff_A_slcV6hqE4_0;
	wire w_dff_A_7L2sUl0W4_0;
	wire w_dff_A_ZSx6VU495_0;
	wire w_dff_A_CX9L5Eh40_0;
	wire w_dff_A_W2hgN4rB7_0;
	wire w_dff_A_wBwQtfQe4_0;
	wire w_dff_A_OHemJ8Og7_0;
	wire w_dff_A_DOG31mfW3_0;
	wire w_dff_A_VFKnqIhs2_0;
	wire w_dff_A_x4nytnbj4_0;
	wire w_dff_A_uvOLy8EJ5_0;
	wire w_dff_A_mKXF3PJ13_0;
	wire w_dff_A_4xpbHIkx7_0;
	wire w_dff_A_fAI54q1Z8_0;
	wire w_dff_A_hHMApKnQ7_0;
	wire w_dff_A_Sc8i3oMz1_0;
	wire w_dff_A_EHHXM7mv5_0;
	wire w_dff_A_HgFIT1074_0;
	wire w_dff_A_tWKdS0U72_0;
	wire w_dff_A_JNmXtZol5_0;
	wire w_dff_A_A1wy8V5y0_0;
	wire w_dff_A_gRruVxYW7_0;
	wire w_dff_A_vAbBGfvT7_0;
	wire w_dff_A_cKuSHqRn2_0;
	wire w_dff_A_EphTaOWz2_0;
	wire w_dff_A_hA8FtDgM4_0;
	wire w_dff_A_BQAqS9To6_0;
	wire w_dff_A_GZ8iJtLX9_0;
	wire w_dff_A_yO26HhJC5_0;
	wire w_dff_A_9tAFCkcm5_0;
	wire w_dff_A_LM3GAe8w9_0;
	wire w_dff_A_Dl0QZvSs6_0;
	wire w_dff_A_8cOZigAO0_0;
	wire w_dff_A_I419XbQu8_0;
	wire w_dff_A_CZA5ch9p3_0;
	wire w_dff_A_5palj88r8_0;
	wire w_dff_A_WS0xxbFA7_0;
	wire w_dff_A_YONsQmPY7_1;
	wire w_dff_A_ANmmdNnK4_0;
	wire w_dff_A_ocVinIXo1_0;
	wire w_dff_A_r2jLnFdC5_0;
	wire w_dff_A_RxI2ZLu16_0;
	wire w_dff_A_IReLaPoU4_0;
	wire w_dff_A_plkQnMZJ0_0;
	wire w_dff_A_9AF9riub7_0;
	wire w_dff_A_aFM7aReY6_0;
	wire w_dff_A_fW4BfWbg9_0;
	wire w_dff_A_S7jIUXO43_0;
	wire w_dff_A_Bjv6ZlqM1_0;
	wire w_dff_A_pZYdD4oV8_0;
	wire w_dff_A_1EjCeFcd6_0;
	wire w_dff_A_tgDDu5xY7_0;
	wire w_dff_A_fn7e7yzk7_0;
	wire w_dff_A_Z28NkXa77_0;
	wire w_dff_A_dRqEIt030_0;
	wire w_dff_A_yyTncQKg7_0;
	wire w_dff_A_uBVxEl2A2_0;
	wire w_dff_A_HhUoXcMG6_0;
	wire w_dff_A_IX4uyESn0_0;
	wire w_dff_A_MpTDP1oo8_0;
	wire w_dff_A_ahQ8esOF0_0;
	wire w_dff_A_lAzi9spV8_0;
	wire w_dff_A_7CfKEnZE7_0;
	wire w_dff_A_B3sh92i29_0;
	wire w_dff_A_vHapubzK1_0;
	wire w_dff_A_RvlRpLbA4_0;
	wire w_dff_A_yUTz5umu0_0;
	wire w_dff_A_CVSsUflQ9_0;
	wire w_dff_A_IexcqqmL7_0;
	wire w_dff_A_A64mRuOH6_0;
	wire w_dff_A_NZNjYFxx6_0;
	wire w_dff_A_MZo8jf6F9_0;
	wire w_dff_A_A4fl1uXn7_0;
	wire w_dff_A_mT9j2k6k2_0;
	wire w_dff_A_esLmSjHq2_0;
	wire w_dff_A_ZdOEwVqN9_0;
	wire w_dff_A_7MrFhR7S7_1;
	wire w_dff_A_TAl1qSZX8_0;
	wire w_dff_A_EYxxYUb76_0;
	wire w_dff_A_jZhC1kvW8_0;
	wire w_dff_A_T53HvLAY2_0;
	wire w_dff_A_nORdTeXw7_0;
	wire w_dff_A_N8JPfGWk1_0;
	wire w_dff_A_isovUuZR6_0;
	wire w_dff_A_3QlqfaK12_0;
	wire w_dff_A_4ive3bFb7_0;
	wire w_dff_A_9n3qgERt5_0;
	wire w_dff_A_mRbFvcOQ5_0;
	wire w_dff_A_aDmuAb4J1_0;
	wire w_dff_A_CowIdsDB3_0;
	wire w_dff_A_DOjiXBQO1_0;
	wire w_dff_A_kL1awfcf6_0;
	wire w_dff_A_dUbhyRtm2_0;
	wire w_dff_A_foOBI6LB9_0;
	wire w_dff_A_OJkDzmtM1_0;
	wire w_dff_A_kwQgiElp5_0;
	wire w_dff_A_tzvoNRdm7_0;
	wire w_dff_A_0uDydB9g0_0;
	wire w_dff_A_9cVVqneJ3_0;
	wire w_dff_A_4EesM9SE6_0;
	wire w_dff_A_fmrxib7m7_0;
	wire w_dff_A_nmoeL7v56_0;
	wire w_dff_A_cKOyWVtE7_0;
	wire w_dff_A_ODhR2nVm7_0;
	wire w_dff_A_4mMJ0EFX4_0;
	wire w_dff_A_psWdfyE05_0;
	wire w_dff_A_SdQ5bftN2_0;
	wire w_dff_A_82CSJO2B4_0;
	wire w_dff_A_3RbBVgOa7_0;
	wire w_dff_A_2K8lkq8h9_0;
	wire w_dff_A_TZcd6i835_0;
	wire w_dff_A_gBHDVGLn4_0;
	wire w_dff_A_TgrAWO958_0;
	wire w_dff_A_39xY3sph6_0;
	wire w_dff_A_BvoqxjG86_0;
	wire w_dff_A_pV3lp2Th7_1;
	wire w_dff_A_KM9CCsM21_0;
	wire w_dff_A_Cz2Bgu0c8_0;
	wire w_dff_A_N2B4mVHN3_0;
	wire w_dff_A_IZCYFMx61_0;
	wire w_dff_A_JXMqe9UU5_0;
	wire w_dff_A_J6Y33yuM1_0;
	wire w_dff_A_dldMPbnL7_0;
	wire w_dff_A_B0MieEWu6_0;
	wire w_dff_A_fJhsAtbk0_0;
	wire w_dff_A_aYLOhwJI1_0;
	wire w_dff_A_tXbivGwa3_0;
	wire w_dff_A_rhnjMU0J6_0;
	wire w_dff_A_V7gHNQQU7_0;
	wire w_dff_A_3EpC6Hfn8_0;
	wire w_dff_A_uTMGRQJi3_0;
	wire w_dff_A_cx9rXWYN8_0;
	wire w_dff_A_hE08VOWD2_0;
	wire w_dff_A_uhHmn1Ot2_0;
	wire w_dff_A_etEJ1VS64_0;
	wire w_dff_A_kDuKOeZi7_0;
	wire w_dff_A_vzR2OpQl1_0;
	wire w_dff_A_f7dHFFwu5_0;
	wire w_dff_A_7SECabTb2_0;
	wire w_dff_A_TQVYDFq34_0;
	wire w_dff_A_ZiNYr72P0_0;
	wire w_dff_A_mwHNqASV5_0;
	wire w_dff_A_5VBQfUnU4_0;
	wire w_dff_A_WDBLBGzs7_0;
	wire w_dff_A_E6KjC8616_0;
	wire w_dff_A_cCK7Y65C8_0;
	wire w_dff_A_HYbqHw3Z4_0;
	wire w_dff_A_9i4A78N81_0;
	wire w_dff_A_gAQA6WhP8_0;
	wire w_dff_A_mBpUqUIy3_0;
	wire w_dff_A_E90cnU9I8_0;
	wire w_dff_A_uzXj0SC12_0;
	wire w_dff_A_PRY3VpPV8_0;
	wire w_dff_A_LzDIyGAn7_0;
	wire w_dff_A_GSYFA4ww3_1;
	wire w_dff_A_UCDwvfB98_0;
	wire w_dff_A_Xwd1dn5f9_0;
	wire w_dff_A_EYxB8Lc47_0;
	wire w_dff_A_xvxn9SEF2_0;
	wire w_dff_A_ivdgl1Ra8_0;
	wire w_dff_A_gjSGCExO3_0;
	wire w_dff_A_7O4fyjTs4_0;
	wire w_dff_A_RPIxa1pk0_0;
	wire w_dff_A_1WqGe35Z3_0;
	wire w_dff_A_UMCk5GSg1_0;
	wire w_dff_A_TJZAYtit9_0;
	wire w_dff_A_nYJVWxya9_0;
	wire w_dff_A_mlj9TEEr2_0;
	wire w_dff_A_q4Q1ISsF1_0;
	wire w_dff_A_qNyI5hBV7_0;
	wire w_dff_A_n0YcfmhI5_0;
	wire w_dff_A_yWCyAVIW2_0;
	wire w_dff_A_MAPhUM7N6_0;
	wire w_dff_A_8kmOKFZ74_0;
	wire w_dff_A_KRYGJYe34_0;
	wire w_dff_A_UkVafpsX8_0;
	wire w_dff_A_pYGMXtPG0_0;
	wire w_dff_A_qgOecMjz3_0;
	wire w_dff_A_AbMDtzDF4_0;
	wire w_dff_A_dOymBiyS4_0;
	wire w_dff_A_5Bc3xjBw8_0;
	wire w_dff_A_7gN0jQnA7_0;
	wire w_dff_A_8nqhAhPU0_0;
	wire w_dff_A_ukHPcTK93_0;
	wire w_dff_A_yMfo0Kd35_0;
	wire w_dff_A_620NMmt57_0;
	wire w_dff_A_PsVygU4V6_0;
	wire w_dff_A_is0H3t9B5_0;
	wire w_dff_A_nB6wTG6c9_0;
	wire w_dff_A_QLHHnaNR3_0;
	wire w_dff_A_rE57DQMO2_0;
	wire w_dff_A_3wSZ1bML4_0;
	wire w_dff_A_dljBLxcc5_0;
	wire w_dff_A_FBQkF7m74_1;
	wire w_dff_A_4fl1TdOT5_0;
	wire w_dff_A_7cGDXaDb1_0;
	wire w_dff_A_IuCW8esC3_0;
	wire w_dff_A_qb2SftNO3_0;
	wire w_dff_A_jf16ptjl6_0;
	wire w_dff_A_kXQcMjmI5_0;
	wire w_dff_A_MC9AYpHi9_0;
	wire w_dff_A_FU5lvZYK5_0;
	wire w_dff_A_G2AYCFir6_0;
	wire w_dff_A_Rj8jANqp8_0;
	wire w_dff_A_ZwqwohQk9_0;
	wire w_dff_A_JU4alewb1_0;
	wire w_dff_A_G1mKw5Sf3_0;
	wire w_dff_A_7F9hztQZ9_0;
	wire w_dff_A_Cm4q8UEB4_0;
	wire w_dff_A_XTssvDHE6_0;
	wire w_dff_A_OA9L6giI5_0;
	wire w_dff_A_sgdFz96H0_0;
	wire w_dff_A_eoSjGsmr2_0;
	wire w_dff_A_0of6W2W81_0;
	wire w_dff_A_pPwfNzyI9_0;
	wire w_dff_A_g3FQySvx7_0;
	wire w_dff_A_da3Hoaiz7_0;
	wire w_dff_A_DLICkPhl6_0;
	wire w_dff_A_q5vmGSpN0_0;
	wire w_dff_A_QgCp5rPq4_0;
	wire w_dff_A_0q3xGcbg7_0;
	wire w_dff_A_7mGhgGiY8_0;
	wire w_dff_A_wGuxlG9W7_0;
	wire w_dff_A_iXikGm2I1_0;
	wire w_dff_A_CrMsD6NM6_0;
	wire w_dff_A_fYF7LZEe3_0;
	wire w_dff_A_FXQNcGJm1_0;
	wire w_dff_A_OAluJ2xm7_0;
	wire w_dff_A_jZ7X0diM9_0;
	wire w_dff_A_Rnd37Xd55_0;
	wire w_dff_A_cFBAvjoj2_0;
	wire w_dff_A_pDcmaUo15_0;
	wire w_dff_A_YfYhlcZP8_1;
	wire w_dff_A_y2t7sUPu6_0;
	wire w_dff_A_42e3Nu0u0_0;
	wire w_dff_A_cMCizrwn5_0;
	wire w_dff_A_czJjS1ol4_0;
	wire w_dff_A_D8RA6Ehk1_0;
	wire w_dff_A_CGgXfMgQ3_0;
	wire w_dff_A_1z2gackJ6_0;
	wire w_dff_A_FzQssm2F1_0;
	wire w_dff_A_jOeeUuAC8_0;
	wire w_dff_A_Nzm3wD5c9_0;
	wire w_dff_A_aspOhlAV4_0;
	wire w_dff_A_gRwurW9b1_0;
	wire w_dff_A_C1R14Pgn4_0;
	wire w_dff_A_zOkywjSZ1_0;
	wire w_dff_A_6ITAj4yy4_0;
	wire w_dff_A_Ny8w7pGi1_0;
	wire w_dff_A_tgvazPQr9_0;
	wire w_dff_A_XssZaBn06_0;
	wire w_dff_A_HqNCbgsy7_0;
	wire w_dff_A_gmSWy4kD0_0;
	wire w_dff_A_NVJbwkiI8_0;
	wire w_dff_A_30yshV7O7_0;
	wire w_dff_A_ijbGCjpS9_0;
	wire w_dff_A_PyzddnWi8_0;
	wire w_dff_A_SQa6CXCT7_0;
	wire w_dff_A_BeRNFGHW5_0;
	wire w_dff_A_MAmaBNb15_0;
	wire w_dff_A_s6PzIUkA3_0;
	wire w_dff_A_peaBLIjd9_0;
	wire w_dff_A_ZpCw35dE1_0;
	wire w_dff_A_FZr2HDck5_0;
	wire w_dff_A_g3Sec77k9_0;
	wire w_dff_A_bjRPVOzQ3_0;
	wire w_dff_A_cEZkXk7w0_0;
	wire w_dff_A_cs3xDGtC2_0;
	wire w_dff_A_gUFwK4nh4_0;
	wire w_dff_A_ir4bMUJO9_0;
	wire w_dff_A_17fmTVMQ1_0;
	wire w_dff_A_tzhGpJqn6_1;
	wire w_dff_A_mfbW9HGd7_0;
	wire w_dff_A_1aixFJQK1_0;
	wire w_dff_A_qngvwCEc1_0;
	wire w_dff_A_sN0Z2cua7_0;
	wire w_dff_A_dYAtbBlm4_0;
	wire w_dff_A_fbKhrtWB5_0;
	wire w_dff_A_mHaWUr5G7_0;
	wire w_dff_A_RTmYkP9I4_0;
	wire w_dff_A_wmlkjIvu1_0;
	wire w_dff_A_NNIsZJ2s8_0;
	wire w_dff_A_PHJ6s1f81_0;
	wire w_dff_A_ymaG0ljj7_0;
	wire w_dff_A_ffOwCtHh2_0;
	wire w_dff_A_U9vRYRLH2_0;
	wire w_dff_A_eeKvm5xK3_0;
	wire w_dff_A_gBq5XAWp6_0;
	wire w_dff_A_6W7CEBAW1_0;
	wire w_dff_A_Xqke8QnJ7_0;
	wire w_dff_A_wzcgwqhc2_0;
	wire w_dff_A_jfkQr8Wy8_0;
	wire w_dff_A_jHi9cTO57_0;
	wire w_dff_A_hgLnWIsW6_0;
	wire w_dff_A_6POL6XvD0_0;
	wire w_dff_A_zIosLDnn4_0;
	wire w_dff_A_grINay6F3_0;
	wire w_dff_A_elW4YhXo0_0;
	wire w_dff_A_M9crSgu92_0;
	wire w_dff_A_PnGGQqeE7_0;
	wire w_dff_A_0EzfcwUL8_0;
	wire w_dff_A_uW7Lqxgf2_0;
	wire w_dff_A_eNYN0uf75_0;
	wire w_dff_A_TrpB85Je6_0;
	wire w_dff_A_EdtrBZVM6_0;
	wire w_dff_A_9DTXmvba8_0;
	wire w_dff_A_Q8ifz1Tj2_0;
	wire w_dff_A_kftT5qGG1_0;
	wire w_dff_A_M7JwIvUK5_0;
	wire w_dff_A_YJ2LTApK3_0;
	wire w_dff_A_Wdw6GYOZ5_1;
	wire w_dff_A_c6AG1F5e9_0;
	wire w_dff_A_FPU5Fyob7_0;
	wire w_dff_A_pZ0c0waE9_0;
	wire w_dff_A_BpMi0wnW0_0;
	wire w_dff_A_tzZuctiQ8_0;
	wire w_dff_A_j3PzZWYR8_0;
	wire w_dff_A_cYq2OVgH2_0;
	wire w_dff_A_h4eQE88U5_0;
	wire w_dff_A_bLkwVTOO0_0;
	wire w_dff_A_Wo661W4s3_0;
	wire w_dff_A_maEm4jcD8_0;
	wire w_dff_A_5zrgfV6c4_0;
	wire w_dff_A_IU2ndIBE5_0;
	wire w_dff_A_UjrdH04g4_0;
	wire w_dff_A_7Zzqu8E70_0;
	wire w_dff_A_9B2wsbLX2_0;
	wire w_dff_A_TunQH81q8_0;
	wire w_dff_A_vGfmp3lQ8_0;
	wire w_dff_A_UM1XqdFl8_0;
	wire w_dff_A_1TsuALWQ3_0;
	wire w_dff_A_wqoUCg256_0;
	wire w_dff_A_9Gj66eJi7_0;
	wire w_dff_A_r7DmmLKM8_0;
	wire w_dff_A_gJFqMbm18_0;
	wire w_dff_A_gBj7IIKO4_0;
	wire w_dff_A_GiRPAt5R9_0;
	wire w_dff_A_UJLviwNg7_0;
	wire w_dff_A_mYuPKgWy0_0;
	wire w_dff_A_i60DtdbK3_0;
	wire w_dff_A_JzBR7V1g5_0;
	wire w_dff_A_wC6rJ1v25_0;
	wire w_dff_A_tG6wXf507_0;
	wire w_dff_A_9F7I295l7_0;
	wire w_dff_A_oqspcb7P1_0;
	wire w_dff_A_L9RCra828_0;
	wire w_dff_A_Eu6vmsRB4_0;
	wire w_dff_A_NRpPcXoQ0_0;
	wire w_dff_A_QJOnwk5p7_0;
	wire w_dff_A_u6wSNtT59_1;
	wire w_dff_A_ogARaZaQ0_0;
	wire w_dff_A_rSFo8fLN2_0;
	wire w_dff_A_4QneGP4k5_0;
	wire w_dff_A_PPMO63dC6_0;
	wire w_dff_A_ZXuj7kq30_0;
	wire w_dff_A_G8RgCPor4_0;
	wire w_dff_A_u6fNNzz82_0;
	wire w_dff_A_kwW7jrr82_0;
	wire w_dff_A_kWwQTSAX4_0;
	wire w_dff_A_XwJzvhkQ0_0;
	wire w_dff_A_gIFPiC2d0_0;
	wire w_dff_A_vHNiVTO56_0;
	wire w_dff_A_9Jol0tfA5_0;
	wire w_dff_A_OKwI49SD0_0;
	wire w_dff_A_sxeuXXAK1_0;
	wire w_dff_A_R2KZCmJI7_0;
	wire w_dff_A_SY1HHCyC5_0;
	wire w_dff_A_JMwCNNkM2_0;
	wire w_dff_A_72IGDjn84_0;
	wire w_dff_A_LE4dsog42_0;
	wire w_dff_A_69ClauPI3_0;
	wire w_dff_A_gfnNGYZI6_0;
	wire w_dff_A_BWridLWQ5_0;
	wire w_dff_A_s3H1Qh1D8_0;
	wire w_dff_A_Gfz1pEMI3_0;
	wire w_dff_A_RdMaJqxI6_0;
	wire w_dff_A_MyygLSgm8_0;
	wire w_dff_A_X1f1yfy10_0;
	wire w_dff_A_Z68Fy68m6_0;
	wire w_dff_A_B9lpOEDx3_0;
	wire w_dff_A_EwgDJfKq0_0;
	wire w_dff_A_v9Ttm6UF0_0;
	wire w_dff_A_PiUU62Jp7_0;
	wire w_dff_A_caZpPZUH7_0;
	wire w_dff_A_SSOOoQON7_0;
	wire w_dff_A_2AzrEH9r2_0;
	wire w_dff_A_tEgdZ2YH3_0;
	wire w_dff_A_FEckNR5b8_0;
	wire w_dff_A_PWRWabNi9_1;
	wire w_dff_A_lgt7miUz1_0;
	wire w_dff_A_EoRT4ScD9_0;
	wire w_dff_A_ztQ7zwNs6_0;
	wire w_dff_A_yf8i2mg22_0;
	wire w_dff_A_k5GE9RK50_0;
	wire w_dff_A_jIOXscPi0_0;
	wire w_dff_A_jypcoECY8_0;
	wire w_dff_A_DZ1OtZQ91_0;
	wire w_dff_A_Gtz2kCmo4_0;
	wire w_dff_A_FLBYrJ0w6_0;
	wire w_dff_A_I2Tvambw9_0;
	wire w_dff_A_8zX5rKx91_0;
	wire w_dff_A_xROupiks4_0;
	wire w_dff_A_lZXXkAYH2_0;
	wire w_dff_A_skHUHohJ2_0;
	wire w_dff_A_SPGAQ09S7_0;
	wire w_dff_A_RyJSeOuc3_0;
	wire w_dff_A_9oAWMnwV5_0;
	wire w_dff_A_itbOQPyI8_0;
	wire w_dff_A_5sJ6YlhE0_0;
	wire w_dff_A_zQTQgKmI8_0;
	wire w_dff_A_YvDT5LJy2_0;
	wire w_dff_A_m5WIJLH01_0;
	wire w_dff_A_w9bbeijX5_0;
	wire w_dff_A_RCp7v3LI6_0;
	wire w_dff_A_hZ2y1I6z7_0;
	wire w_dff_A_O4NcS5zP9_0;
	wire w_dff_A_Ui8WGGKu5_0;
	wire w_dff_A_1mrLadKT3_0;
	wire w_dff_A_1me7KQPp4_0;
	wire w_dff_A_BusWKVox3_0;
	wire w_dff_A_qWhdg15Q7_0;
	wire w_dff_A_ZUpbi2yz0_0;
	wire w_dff_A_pcGYwQm57_0;
	wire w_dff_A_c8K4Cbv56_0;
	wire w_dff_A_9GYIiBBj0_0;
	wire w_dff_A_K0BXssRL8_0;
	wire w_dff_A_lQ0zgZkC0_0;
	wire w_dff_A_EMBTB4wN2_1;
	wire w_dff_A_IoHE6y2G1_0;
	wire w_dff_A_CRCKyV2J4_0;
	wire w_dff_A_It3jCPbb7_0;
	wire w_dff_A_EvQ6WAxz3_0;
	wire w_dff_A_tyTOJb811_0;
	wire w_dff_A_9jO1Pc4Z1_0;
	wire w_dff_A_i0eG4moB5_0;
	wire w_dff_A_PSmzHllw7_0;
	wire w_dff_A_Rj64f1GF7_0;
	wire w_dff_A_duSYX4qP7_0;
	wire w_dff_A_Y0bI5ljX6_0;
	wire w_dff_A_Sk5yPAOL4_0;
	wire w_dff_A_JOo7Meza7_0;
	wire w_dff_A_5MgsQhsR3_0;
	wire w_dff_A_32jWazju9_0;
	wire w_dff_A_OM6qYM0T6_0;
	wire w_dff_A_vhii8myx2_0;
	wire w_dff_A_kpomkAPO6_0;
	wire w_dff_A_qjRaUpfn9_0;
	wire w_dff_A_gSvF2GPJ4_0;
	wire w_dff_A_rccswgV80_0;
	wire w_dff_A_qcqOanec3_0;
	wire w_dff_A_tXEIIjLp2_0;
	wire w_dff_A_AtDqQuHg8_0;
	wire w_dff_A_Q2j1m7Ss5_0;
	wire w_dff_A_aaGHbAOQ6_0;
	wire w_dff_A_Cz7yroOU7_0;
	wire w_dff_A_HLh0ajyc6_0;
	wire w_dff_A_tJ1lhrs51_0;
	wire w_dff_A_nv8A5vB52_0;
	wire w_dff_A_lK8WX9Ux3_0;
	wire w_dff_A_Yc2GXOPw8_0;
	wire w_dff_A_lF1pILYu0_0;
	wire w_dff_A_BwcXCgqW6_0;
	wire w_dff_A_1qNGERZW3_0;
	wire w_dff_A_evvhmfus2_0;
	wire w_dff_A_tE92VkYX4_0;
	wire w_dff_A_1PhMdYyO0_0;
	wire w_dff_A_VAefslF47_1;
	wire w_dff_A_JBKSPWoC8_0;
	wire w_dff_A_OPPhVcSZ0_0;
	wire w_dff_A_a6NZlSbf6_0;
	wire w_dff_A_BXlAGvn60_0;
	wire w_dff_A_X1n7Qtwh0_0;
	wire w_dff_A_yucbsa8e4_0;
	wire w_dff_A_a2QxJeVJ6_0;
	wire w_dff_A_f85D9rMQ2_0;
	wire w_dff_A_64FeIGDE9_0;
	wire w_dff_A_MTcnVtGT9_0;
	wire w_dff_A_8VMW9GZG7_0;
	wire w_dff_A_6aRbW8xq3_0;
	wire w_dff_A_ERLEFsQR9_0;
	wire w_dff_A_FESRtSQO2_0;
	wire w_dff_A_WWBzT8wE6_0;
	wire w_dff_A_Xvy2JFTU7_0;
	wire w_dff_A_o13GDJGJ3_0;
	wire w_dff_A_bQmPcBNf4_0;
	wire w_dff_A_S86RJ6dr8_0;
	wire w_dff_A_5FIWgv9i7_0;
	wire w_dff_A_9qExALMw3_0;
	wire w_dff_A_cVaoeYiy3_0;
	wire w_dff_A_aDuNBe4C2_0;
	wire w_dff_A_9ezcKQ2K6_0;
	wire w_dff_A_sLJL2ump7_0;
	wire w_dff_A_GTgNNpKc9_0;
	wire w_dff_A_4qD0BJyu8_0;
	wire w_dff_A_aDrnXGyr2_0;
	wire w_dff_A_fnaRMI3b3_0;
	wire w_dff_A_ZWBFPxkZ0_0;
	wire w_dff_A_5IOP0DJc7_0;
	wire w_dff_A_OCtiaLFi3_0;
	wire w_dff_A_cUHbVPUs4_0;
	wire w_dff_A_asxETMYj4_0;
	wire w_dff_A_4FAYoMdA1_0;
	wire w_dff_A_dPzmdegS9_0;
	wire w_dff_A_XC1xLJcF0_0;
	wire w_dff_A_STVrNXob7_0;
	wire w_dff_A_upXkuxo17_1;
	wire w_dff_A_Wn9Unnih0_0;
	wire w_dff_A_aJvUgXFv1_0;
	wire w_dff_A_zNFZLKtX5_0;
	wire w_dff_A_rNj0B5FC6_0;
	wire w_dff_A_lb38hRM56_0;
	wire w_dff_A_dDTOJb5V5_0;
	wire w_dff_A_LBsMNjSL7_0;
	wire w_dff_A_NvktGuoa2_0;
	wire w_dff_A_APzxr2dN8_0;
	wire w_dff_A_SbKVvb031_0;
	wire w_dff_A_XRg64ZFO1_0;
	wire w_dff_A_1kMLIqZZ1_0;
	wire w_dff_A_5T4sD9UH3_0;
	wire w_dff_A_z66Swu4g2_0;
	wire w_dff_A_hv17DihY8_0;
	wire w_dff_A_S7WeAWGe3_0;
	wire w_dff_A_d5lJUpOD1_0;
	wire w_dff_A_WWdVHldh0_0;
	wire w_dff_A_ZqE2E6vf6_0;
	wire w_dff_A_pss353h47_0;
	wire w_dff_A_KU1ZnUpb4_0;
	wire w_dff_A_OfuAARV19_0;
	wire w_dff_A_ABqyipJf1_0;
	wire w_dff_A_ZKbfW3Cy0_0;
	wire w_dff_A_IbNmOxoV4_0;
	wire w_dff_A_FZcQF5jg5_0;
	wire w_dff_A_8BLrQC5q1_0;
	wire w_dff_A_wdIYs3126_0;
	wire w_dff_A_rVxrWfsv1_0;
	wire w_dff_A_cyJkNSPU9_0;
	wire w_dff_A_iwU0qOZu8_0;
	wire w_dff_A_D1RKJ3lC8_0;
	wire w_dff_A_NWpkGv7f6_0;
	wire w_dff_A_ixeIN3Wb2_0;
	wire w_dff_A_uumBwDeW0_0;
	wire w_dff_A_mWPf6GnF4_0;
	wire w_dff_A_5Q5DPuZB4_0;
	wire w_dff_A_9HkFBm2c0_0;
	wire w_dff_A_lj9ELOAr8_1;
	wire w_dff_A_6zCZWMoL3_0;
	wire w_dff_A_YSPSA9jN6_0;
	wire w_dff_A_yNx3sJVN3_0;
	wire w_dff_A_JeyC7pDw4_0;
	wire w_dff_A_fZblbgIO6_0;
	wire w_dff_A_6jMTSsvL1_0;
	wire w_dff_A_MqPguq3f9_0;
	wire w_dff_A_kg5IneT15_0;
	wire w_dff_A_olezRIXR0_0;
	wire w_dff_A_v8GcbxwV1_0;
	wire w_dff_A_PTbN5GtS4_0;
	wire w_dff_A_wSNhGyHy5_0;
	wire w_dff_A_ZjRMimW17_0;
	wire w_dff_A_5Tolaqjh3_0;
	wire w_dff_A_YAhmTbcy2_0;
	wire w_dff_A_Z6mvE0qT1_0;
	wire w_dff_A_MEeOtyWo3_0;
	wire w_dff_A_pvT1zztD0_0;
	wire w_dff_A_bGlGukqE6_0;
	wire w_dff_A_7BsqMZ3u1_0;
	wire w_dff_A_v2LvFqxO8_0;
	wire w_dff_A_tpJHmUX28_0;
	wire w_dff_A_S3wmCYtg5_0;
	wire w_dff_A_tE0tCvh50_0;
	wire w_dff_A_cHob9g9y3_0;
	wire w_dff_A_KLvQQeKS0_0;
	wire w_dff_A_kTq0Bqeq0_0;
	wire w_dff_A_rgFVGm4K0_0;
	wire w_dff_A_BqhQa66W8_0;
	wire w_dff_A_dedRN3x89_0;
	wire w_dff_A_G95fJe0B4_0;
	wire w_dff_A_5quZoQEu3_0;
	wire w_dff_A_RjUlvdqL7_0;
	wire w_dff_A_M4eR8Hkc6_0;
	wire w_dff_A_9srIdFhF1_0;
	wire w_dff_A_hTjntdic8_0;
	wire w_dff_A_AoQ929dH0_0;
	wire w_dff_A_PPqc7LGB7_0;
	wire w_dff_A_sDPgk8v97_1;
	wire w_dff_A_cFtTmN0o2_0;
	wire w_dff_A_kiiRQhBW5_0;
	wire w_dff_A_aCe00na87_0;
	wire w_dff_A_o7q1aemK9_0;
	wire w_dff_A_LkEF3ArN2_0;
	wire w_dff_A_qIhctuWI9_0;
	wire w_dff_A_9UhuZQLk7_0;
	wire w_dff_A_jh42ni1M2_0;
	wire w_dff_A_ZdjbCOHO3_0;
	wire w_dff_A_nI3iIqcp4_0;
	wire w_dff_A_mO0rfzEW8_0;
	wire w_dff_A_R41Q2i7T6_0;
	wire w_dff_A_wNCqBHlr2_0;
	wire w_dff_A_4tyyoAOk5_0;
	wire w_dff_A_KjDSevLa3_0;
	wire w_dff_A_A8oEypnS0_0;
	wire w_dff_A_jCSJLyrE3_0;
	wire w_dff_A_XtPCZB0c9_0;
	wire w_dff_A_uivzbkmY3_0;
	wire w_dff_A_UnZckhH29_0;
	wire w_dff_A_cfdmVm6c6_0;
	wire w_dff_A_g3R2Ld1J1_0;
	wire w_dff_A_sLMpOUEi6_0;
	wire w_dff_A_x4it03PW9_0;
	wire w_dff_A_6RVZL74B2_0;
	wire w_dff_A_xzRG97JL2_0;
	wire w_dff_A_UnLuVhtN9_0;
	wire w_dff_A_DGmXZjIi2_0;
	wire w_dff_A_CKi4v38a2_0;
	wire w_dff_A_abXsWAze8_0;
	wire w_dff_A_KoiKCyJb4_0;
	wire w_dff_A_MqFItUqQ6_0;
	wire w_dff_A_v0gvGUCS7_0;
	wire w_dff_A_wGcUSNGe5_0;
	wire w_dff_A_jafLSeyt9_0;
	wire w_dff_A_IytHxavg9_0;
	wire w_dff_A_dtEdkBdj1_0;
	wire w_dff_A_urSSzUsM1_0;
	wire w_dff_A_onEfvwvV6_1;
	wire w_dff_A_C0HUjNaI0_0;
	wire w_dff_A_mgP1VW8e0_0;
	wire w_dff_A_SxvRvK4p9_0;
	wire w_dff_A_tx07HFfa9_0;
	wire w_dff_A_JxFFZbCP5_0;
	wire w_dff_A_21UPNdX36_0;
	wire w_dff_A_b0JFeInU2_0;
	wire w_dff_A_lCUkQlQe8_0;
	wire w_dff_A_VhomK8Ca7_0;
	wire w_dff_A_5uZiJa7h7_0;
	wire w_dff_A_8tQoMJoe3_0;
	wire w_dff_A_Nfx7iYoX8_0;
	wire w_dff_A_Rprol9ET7_0;
	wire w_dff_A_2QPmdr2n1_0;
	wire w_dff_A_O9ojFsQs8_0;
	wire w_dff_A_4C5FZ3pB9_0;
	wire w_dff_A_nzP6p3E90_0;
	wire w_dff_A_R1PTbvuf4_0;
	wire w_dff_A_ogzJ2vlA4_0;
	wire w_dff_A_Ib00GUvM9_0;
	wire w_dff_A_tyVrybjw2_0;
	wire w_dff_A_okzfNU0q0_0;
	wire w_dff_A_dmrZLSd61_0;
	wire w_dff_A_sx9RMHmI6_0;
	wire w_dff_A_xRM73C7k6_0;
	wire w_dff_A_bnrbDias4_0;
	wire w_dff_A_9Qz45vB73_0;
	wire w_dff_A_s4JSap4n0_0;
	wire w_dff_A_CSwzjaeg9_0;
	wire w_dff_A_MeX7d2zu9_0;
	wire w_dff_A_iVJy5de78_0;
	wire w_dff_A_kpk24sAm7_0;
	wire w_dff_A_laKRt4fM5_0;
	wire w_dff_A_cIddYTD10_0;
	wire w_dff_A_HPZGDjGW3_0;
	wire w_dff_A_NaAAazET6_0;
	wire w_dff_A_MjseTzEz5_0;
	wire w_dff_A_OCoChaKG9_0;
	wire w_dff_A_XmweTCKr8_1;
	wire w_dff_A_EOGxKO371_0;
	wire w_dff_A_lUU18J799_0;
	wire w_dff_A_afXMxmPS7_0;
	wire w_dff_A_PBRVivZf7_0;
	wire w_dff_A_cLRFLt8e4_0;
	wire w_dff_A_4MjlSl9h2_0;
	wire w_dff_A_7D4SMPgx0_0;
	wire w_dff_A_L6EcYAQY8_0;
	wire w_dff_A_xWN4Yt747_0;
	wire w_dff_A_jha5NDAS0_0;
	wire w_dff_A_V6VZFrcV5_0;
	wire w_dff_A_GxTS27pS3_0;
	wire w_dff_A_6hAUldyh3_0;
	wire w_dff_A_ddzQnE3b7_0;
	wire w_dff_A_r17Fx0cV3_0;
	wire w_dff_A_zJstR2UV3_0;
	wire w_dff_A_ZZo8oM4s1_0;
	wire w_dff_A_uiHvil4E4_0;
	wire w_dff_A_OgxjZZWi3_0;
	wire w_dff_A_0DEc0Ifc7_0;
	wire w_dff_A_Hqlz0k4G8_0;
	wire w_dff_A_JFUymT810_0;
	wire w_dff_A_j4gFUobs9_0;
	wire w_dff_A_zCm0H4ih5_0;
	wire w_dff_A_l1HCIKy98_0;
	wire w_dff_A_ivmLM9J73_0;
	wire w_dff_A_e1PfDYZZ5_0;
	wire w_dff_A_EJOAexXK6_0;
	wire w_dff_A_5tUFrWPk6_0;
	wire w_dff_A_4WgN97nv7_0;
	wire w_dff_A_71mgfxK79_0;
	wire w_dff_A_2RKqtE8q8_0;
	wire w_dff_A_OQarV7mi0_0;
	wire w_dff_A_CXHTQpki3_0;
	wire w_dff_A_lOjk2tqx1_0;
	wire w_dff_A_UbleewQs0_0;
	wire w_dff_A_6RZk2ynx8_0;
	wire w_dff_A_r0VOjmTD7_0;
	wire w_dff_A_FwloGYnx1_1;
	wire w_dff_A_MpMoED0o2_0;
	wire w_dff_A_ch9L710B3_0;
	wire w_dff_A_ZdqSW84s7_0;
	wire w_dff_A_tpuMJF1Z5_0;
	wire w_dff_A_L19tyCWl8_0;
	wire w_dff_A_FfUc06ZZ5_0;
	wire w_dff_A_vJEhMdfj2_0;
	wire w_dff_A_xUBEpP752_0;
	wire w_dff_A_OU8g8YTV9_0;
	wire w_dff_A_jI4NSncm5_0;
	wire w_dff_A_ExDix2BP4_0;
	wire w_dff_A_d1PfQ0OE5_0;
	wire w_dff_A_kFxObhhO4_0;
	wire w_dff_A_ncMbpdAA2_0;
	wire w_dff_A_xgZvbUCQ1_0;
	wire w_dff_A_NcEbcPEE4_0;
	wire w_dff_A_cQBgkh7U3_0;
	wire w_dff_A_FmFIRANR1_0;
	wire w_dff_A_ihbKzhFi8_0;
	wire w_dff_A_mwdLyVdM1_0;
	wire w_dff_A_waHtKHPG7_0;
	wire w_dff_A_VK5CuF4n3_0;
	wire w_dff_A_BqFHOsmc8_0;
	wire w_dff_A_rcbVpIZv6_0;
	wire w_dff_A_9I9mWfGf7_0;
	wire w_dff_A_WKRtswHN5_0;
	wire w_dff_A_JSQxALEH2_0;
	wire w_dff_A_gpUwEeBL5_0;
	wire w_dff_A_ukvlCemw2_0;
	wire w_dff_A_KzXZROGU7_0;
	wire w_dff_A_TA578Zcc5_0;
	wire w_dff_A_4vJ2qQSY1_0;
	wire w_dff_A_IvvnpkiF6_0;
	wire w_dff_A_AyYapmSO7_0;
	wire w_dff_A_HsREqVyM5_0;
	wire w_dff_A_WOX5bTVf0_0;
	wire w_dff_A_Z0lg9tPg8_0;
	wire w_dff_A_QTMORFDm9_0;
	wire w_dff_A_gHt6hTma0_1;
	wire w_dff_A_nGPHs6QH5_0;
	wire w_dff_A_uOJwQ9EU1_0;
	wire w_dff_A_gfcJcOOx0_0;
	wire w_dff_A_F7mCBWlE7_0;
	wire w_dff_A_EBEOMbHW7_0;
	wire w_dff_A_9JseOFDB8_0;
	wire w_dff_A_o5nw1aGP8_0;
	wire w_dff_A_VnYT1duh6_0;
	wire w_dff_A_oWnjtQHt0_0;
	wire w_dff_A_Xs0om2bb3_0;
	wire w_dff_A_XxqiivVE8_0;
	wire w_dff_A_Wu7bGLzd4_0;
	wire w_dff_A_OSeIN3mp3_0;
	wire w_dff_A_drHUhbxT6_0;
	wire w_dff_A_YCZBGw692_0;
	wire w_dff_A_WAA0KjYz8_0;
	wire w_dff_A_ab9WmRfo5_0;
	wire w_dff_A_bHf2jcQN0_0;
	wire w_dff_A_JwPBoHa24_0;
	wire w_dff_A_mgby5pHw4_0;
	wire w_dff_A_LrOop5077_0;
	wire w_dff_A_lyPcdTvj1_0;
	wire w_dff_A_ZbaFq0o53_0;
	wire w_dff_A_c8rCM2qO0_0;
	wire w_dff_A_ZsWwFhcn1_0;
	wire w_dff_A_qJWzWsOf1_0;
	wire w_dff_A_0cU1KyT65_0;
	wire w_dff_A_tVbzCKHm5_0;
	wire w_dff_A_Izf5pvUg1_0;
	wire w_dff_A_42cxK4HZ5_0;
	wire w_dff_A_s2bNsu3r9_0;
	wire w_dff_A_mKO50t8y6_0;
	wire w_dff_A_NzuRFX0n9_0;
	wire w_dff_A_GeqN5l1K8_0;
	wire w_dff_A_5dImG5CV1_0;
	wire w_dff_A_GzHL9uzS9_0;
	wire w_dff_A_YCfI5aSf9_0;
	wire w_dff_A_sj9zNDpl1_0;
	wire w_dff_A_ljXzS98X0_1;
	wire w_dff_A_nOUr4nCw7_0;
	wire w_dff_A_BJFfyCt24_0;
	wire w_dff_A_NssCCimR2_0;
	wire w_dff_A_vPecCN0Y5_0;
	wire w_dff_A_f71xhcAR6_0;
	wire w_dff_A_PMB24OEl9_0;
	wire w_dff_A_gBHfUDLO7_0;
	wire w_dff_A_kwDnf1YH3_0;
	wire w_dff_A_q01KOlLi4_0;
	wire w_dff_A_t9nSfTNf9_0;
	wire w_dff_A_XqfoWssA8_0;
	wire w_dff_A_BTadeR402_0;
	wire w_dff_A_gX4cizWR7_0;
	wire w_dff_A_GnAbyRYC6_0;
	wire w_dff_A_MhZzZ5S27_0;
	wire w_dff_A_tdjnYDGm7_0;
	wire w_dff_A_cRn642oY2_0;
	wire w_dff_A_zQQKaLSp1_0;
	wire w_dff_A_fQvN1Xop9_0;
	wire w_dff_A_SIpWHAIr0_0;
	wire w_dff_A_vCCayale7_0;
	wire w_dff_A_fCk9bUh52_0;
	wire w_dff_A_tTQS9OPy8_0;
	wire w_dff_A_ut354afT3_0;
	wire w_dff_A_PTWxS2P06_0;
	wire w_dff_A_O9fVmEKK9_0;
	wire w_dff_A_QwLftZj48_0;
	wire w_dff_A_vsW6Xe1B0_0;
	wire w_dff_A_fn55Qm2Y0_0;
	wire w_dff_A_9eAIXyDp9_0;
	wire w_dff_A_VI4x1DKG9_0;
	wire w_dff_A_smGqW4zp3_0;
	wire w_dff_A_bb7P065s6_0;
	wire w_dff_A_bzO6WC0P9_0;
	wire w_dff_A_m2lgcgiZ9_0;
	wire w_dff_A_B6JKsWB17_0;
	wire w_dff_A_EulQXWeM5_0;
	wire w_dff_A_YPZ0QiCN5_0;
	wire w_dff_A_xShgKWs03_1;
	wire w_dff_A_kjO7M7KU8_0;
	wire w_dff_A_pGW84IGQ2_0;
	wire w_dff_A_1fWjeC0q6_0;
	wire w_dff_A_5MVLNlnI4_0;
	wire w_dff_A_wj4bYWy55_0;
	wire w_dff_A_fsKaOxVv5_0;
	wire w_dff_A_Yd3fyowR6_0;
	wire w_dff_A_4i3Q8WXZ6_0;
	wire w_dff_A_mxIET3BN6_0;
	wire w_dff_A_dGalxtaK2_0;
	wire w_dff_A_YkbXa5gH2_0;
	wire w_dff_A_lAMTkiGl1_0;
	wire w_dff_A_P2ywUzQV6_0;
	wire w_dff_A_WVY41mYz5_0;
	wire w_dff_A_GRi7oGyP1_0;
	wire w_dff_A_C0XZ1sFN3_0;
	wire w_dff_A_hi5RjgWL4_0;
	wire w_dff_A_A54dNGGp2_0;
	wire w_dff_A_xkBHSLTv2_0;
	wire w_dff_A_9NHPVGUc4_0;
	wire w_dff_A_gZE3wzeU3_0;
	wire w_dff_A_8ebbw5fz1_0;
	wire w_dff_A_rbnwV7Kj3_0;
	wire w_dff_A_Eh7rDtQW0_0;
	wire w_dff_A_9SWQ4wJ61_0;
	wire w_dff_A_qf0SmeG78_0;
	wire w_dff_A_Kkua1hZT1_0;
	wire w_dff_A_1tDb3pRP3_0;
	wire w_dff_A_surpiXqi2_0;
	wire w_dff_A_YXqfAoT57_0;
	wire w_dff_A_OO1CgwT00_0;
	wire w_dff_A_5TJHJzXw2_0;
	wire w_dff_A_LN9KTim27_0;
	wire w_dff_A_IzRFCL2H7_0;
	wire w_dff_A_GQC5mO9W5_0;
	wire w_dff_A_DaZSYZLk9_0;
	wire w_dff_A_Pqw0gOc15_0;
	wire w_dff_A_3IgEP2Jy8_0;
	wire w_dff_A_38sqavEp5_1;
	wire w_dff_A_Zs3qjdnn7_0;
	wire w_dff_A_1JT9aWSp4_0;
	wire w_dff_A_siffhDvj1_0;
	wire w_dff_A_4rQIcuBA1_0;
	wire w_dff_A_cSmseDur7_0;
	wire w_dff_A_H1OnigFP3_0;
	wire w_dff_A_czdYhQzf2_0;
	wire w_dff_A_ryuN8gsJ3_0;
	wire w_dff_A_pfTH7akb9_0;
	wire w_dff_A_QVSJHuk56_0;
	wire w_dff_A_MJXx3tXE2_0;
	wire w_dff_A_2VMtCcSr6_0;
	wire w_dff_A_Be2b51nP8_0;
	wire w_dff_A_Phgue6VH0_0;
	wire w_dff_A_zNKwNga97_0;
	wire w_dff_A_l3gqVx2B1_0;
	wire w_dff_A_w47ceNUJ4_0;
	wire w_dff_A_5uyAgXWX0_0;
	wire w_dff_A_TtWs1HRA1_0;
	wire w_dff_A_qsKlg1Qx5_0;
	wire w_dff_A_vu3d9g8D5_0;
	wire w_dff_A_xs121gWN4_0;
	wire w_dff_A_XvqHuXFx8_0;
	wire w_dff_A_WMIFTPsb4_0;
	wire w_dff_A_mKcd5Wzp7_0;
	wire w_dff_A_Znl8z9bx8_0;
	wire w_dff_A_ure21g7j4_0;
	wire w_dff_A_eaLZXhEP2_0;
	wire w_dff_A_wyt5FgrK6_0;
	wire w_dff_A_dFcjsN7R2_0;
	wire w_dff_A_WjliDwrF1_0;
	wire w_dff_A_Yz1i94GP0_0;
	wire w_dff_A_KCOoc4MH6_0;
	wire w_dff_A_a42OPxXh5_0;
	wire w_dff_A_S39VlzLt6_0;
	wire w_dff_A_uWsDV42Q3_0;
	wire w_dff_A_5csQeihD0_0;
	wire w_dff_A_qxYRl1AQ1_0;
	wire w_dff_A_DLdvL5Ht9_1;
	wire w_dff_A_HOcIIMqs8_0;
	wire w_dff_A_hoznheuJ8_0;
	wire w_dff_A_rAYN32AO2_0;
	wire w_dff_A_rLEFmK6y2_0;
	wire w_dff_A_L6XdCxsM8_0;
	wire w_dff_A_bWjUG67T1_0;
	wire w_dff_A_O5nDktmS3_0;
	wire w_dff_A_FLNitFLc8_0;
	wire w_dff_A_tMsHjJkH2_0;
	wire w_dff_A_UUhXu5p53_0;
	wire w_dff_A_2XVEdEIp7_0;
	wire w_dff_A_EpM0sfpu3_0;
	wire w_dff_A_z2ub1JVL2_0;
	wire w_dff_A_xjb6HRGR7_0;
	wire w_dff_A_jngDomR09_0;
	wire w_dff_A_K9nYleKo0_0;
	wire w_dff_A_YgD4JF749_0;
	wire w_dff_A_PatGGNCK5_0;
	wire w_dff_A_dsW7JR7S4_0;
	wire w_dff_A_jAR6E5a07_0;
	wire w_dff_A_bVnPyNSV0_0;
	wire w_dff_A_hwVmDXjr0_0;
	wire w_dff_A_Kzan7UU56_0;
	wire w_dff_A_yF40Rt5Y4_0;
	wire w_dff_A_DDAFCUvJ3_0;
	wire w_dff_A_xB6wulfQ6_0;
	wire w_dff_A_cNjKZeet2_0;
	wire w_dff_A_28m52jwX9_0;
	wire w_dff_A_9CZbkAR68_0;
	wire w_dff_A_qDRc3Jw05_0;
	wire w_dff_A_hxum9Leg2_0;
	wire w_dff_A_CF9t3HuT2_0;
	wire w_dff_A_ceVtjhnF2_0;
	wire w_dff_A_K4LptOkN3_0;
	wire w_dff_A_U4hyG6aO5_0;
	wire w_dff_A_ImkWfIsC8_0;
	wire w_dff_A_n0NYp1dL5_0;
	wire w_dff_A_b9rPRZxf7_0;
	wire w_dff_A_EW0imUD51_1;
	wire w_dff_A_26C0lEin4_0;
	wire w_dff_A_wINPRdya4_0;
	wire w_dff_A_pXTcFp8K9_0;
	wire w_dff_A_t3T7prDM5_0;
	wire w_dff_A_eBpafFru6_0;
	wire w_dff_A_oryNXrsh3_0;
	wire w_dff_A_pSLTGfiz8_0;
	wire w_dff_A_tPV5bS8u1_0;
	wire w_dff_A_GeGU1QUC8_0;
	wire w_dff_A_XiUMFY6i1_0;
	wire w_dff_A_w99GgYdx4_0;
	wire w_dff_A_s7QlhHlg1_0;
	wire w_dff_A_Etx7XtMV4_0;
	wire w_dff_A_lbbHW5266_0;
	wire w_dff_A_sKzts2hu5_0;
	wire w_dff_A_wqyYimta8_0;
	wire w_dff_A_uU8jEQhe4_0;
	wire w_dff_A_YYva5GVY8_0;
	wire w_dff_A_94xw8laE5_0;
	wire w_dff_A_dILC9Khq9_0;
	wire w_dff_A_2qdXm90B8_0;
	wire w_dff_A_q5P21ugw6_0;
	wire w_dff_A_3TlxiIuo9_0;
	wire w_dff_A_01JH3J1W4_0;
	wire w_dff_A_Ril6aFfp9_0;
	wire w_dff_A_FrqJ7RtD0_0;
	wire w_dff_A_b8kAt2EB8_0;
	wire w_dff_A_eatSQTXx9_0;
	wire w_dff_A_lZiGRDVi9_0;
	wire w_dff_A_PKa4odit5_0;
	wire w_dff_A_hzjcbEMe3_0;
	wire w_dff_A_JUIwAcP90_0;
	wire w_dff_A_7Zx8ASuy4_0;
	wire w_dff_A_vAl48w8K5_0;
	wire w_dff_A_KV5L78DF2_0;
	wire w_dff_A_NbQIdvFX0_0;
	wire w_dff_A_jANELNGQ5_0;
	wire w_dff_A_Wg2Zu0QT2_0;
	wire w_dff_A_pZScGDyA2_1;
	wire w_dff_A_Dz0znsbc8_0;
	wire w_dff_A_LJveWNLP7_0;
	wire w_dff_A_hYlLDHVy5_0;
	wire w_dff_A_oWA8x1w36_0;
	wire w_dff_A_4hhUBxVE4_0;
	wire w_dff_A_Sfop3p7p8_0;
	wire w_dff_A_PUMgXenJ7_0;
	wire w_dff_A_uc13hQny4_0;
	wire w_dff_A_toIw3Va90_0;
	wire w_dff_A_OK1tV9WE5_0;
	wire w_dff_A_e6k42ZkM0_0;
	wire w_dff_A_1uZx7O7X2_0;
	wire w_dff_A_SWTDTC4A3_0;
	wire w_dff_A_ATjbpP5w8_0;
	wire w_dff_A_F7bHCY530_0;
	wire w_dff_A_Bw9tKLlx7_0;
	wire w_dff_A_5aPjWhOc5_0;
	wire w_dff_A_OgSL8DjQ5_0;
	wire w_dff_A_7phPNwun4_0;
	wire w_dff_A_Gboaby8G3_0;
	wire w_dff_A_RTNloDsB1_0;
	wire w_dff_A_mZPJaOnL3_0;
	wire w_dff_A_cb0gjv0B3_0;
	wire w_dff_A_srQ33LFz4_0;
	wire w_dff_A_UAaU5ua07_0;
	wire w_dff_A_SESMrgmB8_0;
	wire w_dff_A_ttbdKH5X0_0;
	wire w_dff_A_w0xWYzyw2_0;
	wire w_dff_A_OuQnam1G8_0;
	wire w_dff_A_rzB2tTdl4_0;
	wire w_dff_A_74XDc4Gf3_0;
	wire w_dff_A_Hysq3mT26_0;
	wire w_dff_A_x2js2btP5_0;
	wire w_dff_A_8qxLEd5G3_0;
	wire w_dff_A_GoKdhjaH3_0;
	wire w_dff_A_xid1jguN1_0;
	wire w_dff_A_nvwqbOaQ0_0;
	wire w_dff_A_uAzFVU012_0;
	wire w_dff_A_s9CBI2X99_1;
	wire w_dff_A_5j4X6org3_0;
	wire w_dff_A_o8iTZWdY2_0;
	wire w_dff_A_P4vQ4pzD5_0;
	wire w_dff_A_unbKZawH9_0;
	wire w_dff_A_35C307ns7_0;
	wire w_dff_A_tV1Kezob9_0;
	wire w_dff_A_REkXp1r70_0;
	wire w_dff_A_WUrqD82e6_0;
	wire w_dff_A_5x2nP9jM6_0;
	wire w_dff_A_GzdYYtnu4_0;
	wire w_dff_A_M8ltJ3DN2_0;
	wire w_dff_A_YAhXaJ6b0_0;
	wire w_dff_A_586ElPPZ2_0;
	wire w_dff_A_rS5yQATm5_0;
	wire w_dff_A_yI3DnthI3_0;
	wire w_dff_A_0OP8pJvZ1_0;
	wire w_dff_A_m5xsyH0s3_0;
	wire w_dff_A_B2gofKCl5_0;
	wire w_dff_A_H6WoT1RM1_0;
	wire w_dff_A_LvF4yQfq3_0;
	wire w_dff_A_nE6UP5G59_0;
	wire w_dff_A_APzV3JU79_0;
	wire w_dff_A_FdlJiHep2_0;
	wire w_dff_A_sumutRLf2_0;
	wire w_dff_A_Fmc8i1Op4_0;
	wire w_dff_A_saZHOdSU0_0;
	wire w_dff_A_3GP0EtA17_0;
	wire w_dff_A_4GEYyXez1_0;
	wire w_dff_A_VxlFqlQU1_0;
	wire w_dff_A_AUPmesxs4_0;
	wire w_dff_A_8xehiPFf6_0;
	wire w_dff_A_zWkRpF5C4_0;
	wire w_dff_A_LM15TwUm5_0;
	wire w_dff_A_YVNYLe6J0_0;
	wire w_dff_A_ijOsg7Oa3_0;
	wire w_dff_A_EXZmuuH19_0;
	wire w_dff_A_3zZ4H4rX1_0;
	wire w_dff_A_FmHOqaXh5_0;
	wire w_dff_A_ltJWpPGm4_1;
	wire w_dff_A_bTj4dEHH2_0;
	wire w_dff_A_n8ApaKVc7_0;
	wire w_dff_A_KcfK5MyF3_0;
	wire w_dff_A_pE7lSduZ5_0;
	wire w_dff_A_YiQbfKdg3_0;
	wire w_dff_A_D69IDZIi1_0;
	wire w_dff_A_yRF65uNC9_0;
	wire w_dff_A_YjkzyKuc2_0;
	wire w_dff_A_TWTwWK5n6_0;
	wire w_dff_A_yPgFgPSA9_0;
	wire w_dff_A_sGQUdmmi7_0;
	wire w_dff_A_i6TZp9aW1_0;
	wire w_dff_A_N7DxbTFP1_0;
	wire w_dff_A_PP9eikLr5_0;
	wire w_dff_A_VLGLq12v6_0;
	wire w_dff_A_Wu7GTIuA1_0;
	wire w_dff_A_EY5H5PSt2_0;
	wire w_dff_A_VTdLg4rc3_0;
	wire w_dff_A_ZSDcuK9b9_0;
	wire w_dff_A_hMNeXxaf3_0;
	wire w_dff_A_Yvj76dXK0_0;
	wire w_dff_A_Oxxn2wMM0_0;
	wire w_dff_A_73939TPZ4_0;
	wire w_dff_A_cCQA6j7L3_0;
	wire w_dff_A_PF9gHu5I0_0;
	wire w_dff_A_PjWrK1Ch8_0;
	wire w_dff_A_bz0hL5Dy8_0;
	wire w_dff_A_PF4f4Foc7_0;
	wire w_dff_A_TmwLJyQp7_0;
	wire w_dff_A_nJBGiABp0_0;
	wire w_dff_A_orQpsPhc2_0;
	wire w_dff_A_7A4MWDON8_0;
	wire w_dff_A_vbzK9DWS0_0;
	wire w_dff_A_SrlVGlhG1_0;
	wire w_dff_A_6cxfcSvs8_0;
	wire w_dff_A_hGP8F4OX5_0;
	wire w_dff_A_i6mFKTzI7_0;
	wire w_dff_A_KDNPJ6ir4_0;
	wire w_dff_A_YJS1iCK09_1;
	wire w_dff_A_TbVdD3vB2_0;
	wire w_dff_A_NnG0DdCZ7_0;
	wire w_dff_A_0Mw1IltL6_0;
	wire w_dff_A_KMqhhc703_0;
	wire w_dff_A_UgpTv6zH6_0;
	wire w_dff_A_gagAgT4D0_0;
	wire w_dff_A_X9OInrxT8_0;
	wire w_dff_A_edachBqU8_0;
	wire w_dff_A_o8L9tTTP2_0;
	wire w_dff_A_t5yS1FMO9_0;
	wire w_dff_A_2QeghzNY7_0;
	wire w_dff_A_uiJ2ECX90_0;
	wire w_dff_A_ZESKld5F3_0;
	wire w_dff_A_qddnKWYm6_0;
	wire w_dff_A_QmZJafKr2_0;
	wire w_dff_A_Ia459EA71_0;
	wire w_dff_A_P4GwI2Vz9_0;
	wire w_dff_A_8dHBC7Oa4_0;
	wire w_dff_A_1CPyePqK3_0;
	wire w_dff_A_XVkRIzdC1_0;
	wire w_dff_A_17zQs4O20_0;
	wire w_dff_A_2ih7ywQW7_0;
	wire w_dff_A_3VKPvNBR8_0;
	wire w_dff_A_wJWYmI1s0_0;
	wire w_dff_A_46ZLSEbS5_0;
	wire w_dff_A_ejOkQggK5_0;
	wire w_dff_A_S9o3y3cQ1_0;
	wire w_dff_A_jO09T9Oj6_0;
	wire w_dff_A_s1PEjzWx4_0;
	wire w_dff_A_J4QPgZ4j4_0;
	wire w_dff_A_UyQeu1gk3_0;
	wire w_dff_A_jf9T34HT1_0;
	wire w_dff_A_0lHXl7NV9_0;
	wire w_dff_A_EV38FxhT5_0;
	wire w_dff_A_PKVQcffY0_0;
	wire w_dff_A_8hyZE7070_0;
	wire w_dff_A_0FAgAEJO9_0;
	wire w_dff_A_SnNak6mp8_0;
	wire w_dff_A_ThUKi2cH2_1;
	wire w_dff_A_xn8OdA137_0;
	wire w_dff_A_VX6DQ02v2_0;
	wire w_dff_A_qQFbfMUI1_0;
	wire w_dff_A_SZZlzdoY1_0;
	wire w_dff_A_9x1ZqXLj1_0;
	wire w_dff_A_lZ8gwEzV6_0;
	wire w_dff_A_TTy78zse9_0;
	wire w_dff_A_dkYbxvAD5_0;
	wire w_dff_A_rVubgCGZ7_0;
	wire w_dff_A_u0KJr7cm1_0;
	wire w_dff_A_iHkEg4030_0;
	wire w_dff_A_67zJikhZ5_0;
	wire w_dff_A_ARQmbsby9_0;
	wire w_dff_A_SvRG6qyz2_0;
	wire w_dff_A_hS4mnYRb5_0;
	wire w_dff_A_UmqymFCp1_0;
	wire w_dff_A_uCk6lHbm7_0;
	wire w_dff_A_OR48rN5f0_0;
	wire w_dff_A_9RxGd0mk4_0;
	wire w_dff_A_0t1bdfl26_0;
	wire w_dff_A_VhCp261p1_0;
	wire w_dff_A_ILBL7SRY2_0;
	wire w_dff_A_j3mpOVkK7_0;
	wire w_dff_A_2AhICZnV6_0;
	wire w_dff_A_Xqm8grg42_0;
	wire w_dff_A_byw5h8b02_0;
	wire w_dff_A_ftFp8D6W9_0;
	wire w_dff_A_j2sNVIHr0_0;
	wire w_dff_A_8nDB3CRG2_0;
	wire w_dff_A_B5AJLaOR1_0;
	wire w_dff_A_nZcpkXBO8_0;
	wire w_dff_A_5U2Bz5y88_0;
	wire w_dff_A_uEbCVBHr1_0;
	wire w_dff_A_oQb8kAjb1_0;
	wire w_dff_A_IywEnK069_0;
	wire w_dff_A_vEQNVOj77_0;
	wire w_dff_A_pRi1a1yi5_0;
	wire w_dff_A_27Rgy5BW4_0;
	wire w_dff_A_7DWNk9T28_1;
	wire w_dff_A_GPbwSp8Y7_0;
	wire w_dff_A_MS3QaBnO0_0;
	wire w_dff_A_RCPFmIum0_0;
	wire w_dff_A_neqVBslu4_0;
	wire w_dff_A_KmsC0oP25_0;
	wire w_dff_A_MILeSvMh8_0;
	wire w_dff_A_KOgqUn8M5_0;
	wire w_dff_A_h9b3Mp9F5_0;
	wire w_dff_A_eDz3EFhw6_0;
	wire w_dff_A_quOz00uA6_0;
	wire w_dff_A_nBPxCYg98_0;
	wire w_dff_A_3t2382n48_0;
	wire w_dff_A_QvNZENNn7_0;
	wire w_dff_A_2AnsEprB6_0;
	wire w_dff_A_ZHgUQeHx9_0;
	wire w_dff_A_nRGZjNJJ2_0;
	wire w_dff_A_oOCp26wR0_0;
	wire w_dff_A_jAfaHDjI4_0;
	wire w_dff_A_92NsBwqc2_0;
	wire w_dff_A_D6IxUAoF9_0;
	wire w_dff_A_VBz9XKmS4_0;
	wire w_dff_A_1YgUQNqL8_0;
	wire w_dff_A_S6Jrppwh8_0;
	wire w_dff_A_qHubb2Kl7_0;
	wire w_dff_A_5yPzmDu28_0;
	wire w_dff_A_po4c7hv07_0;
	wire w_dff_A_zpz9j1RA2_0;
	wire w_dff_A_jumjBDQd2_0;
	wire w_dff_A_L8x3EYEC8_0;
	wire w_dff_A_XFamfHR42_0;
	wire w_dff_A_gLD2oU346_0;
	wire w_dff_A_R8nDrZIW9_0;
	wire w_dff_A_020cK1fd5_0;
	wire w_dff_A_qRr5YlwW2_0;
	wire w_dff_A_yHEuMzV22_0;
	wire w_dff_A_miszG4F57_0;
	wire w_dff_A_iZWM93os3_0;
	wire w_dff_A_lXXplaG52_0;
	wire w_dff_A_KWb9btUV8_1;
	wire w_dff_A_7wQgQEAD2_0;
	wire w_dff_A_1QoJXjGR3_0;
	wire w_dff_A_QFdvQS6w0_0;
	wire w_dff_A_A9KPtago5_0;
	wire w_dff_A_WdZgDvQ91_0;
	wire w_dff_A_Ok5dBrgs0_0;
	wire w_dff_A_f2s49wTY3_0;
	wire w_dff_A_pOfHl5DV2_0;
	wire w_dff_A_T4dIaOIi1_0;
	wire w_dff_A_FTgag51p5_0;
	wire w_dff_A_czAU8MEn8_0;
	wire w_dff_A_I7yfueF96_0;
	wire w_dff_A_fdwEG1Nz3_0;
	wire w_dff_A_ZniZFP1Y8_0;
	wire w_dff_A_23MY2xiG1_0;
	wire w_dff_A_UpeCYdxG6_0;
	wire w_dff_A_WyfAiTCP8_0;
	wire w_dff_A_ElcTUQB91_0;
	wire w_dff_A_EDpJjPvG1_0;
	wire w_dff_A_AkCpCpk23_0;
	wire w_dff_A_sImYZN0Z7_0;
	wire w_dff_A_Dcmsywqt3_0;
	wire w_dff_A_G17aN4Ui6_0;
	wire w_dff_A_ihS8N92j6_0;
	wire w_dff_A_chl4Yehu0_0;
	wire w_dff_A_g5guW00w0_0;
	wire w_dff_A_PCZMgcec4_0;
	wire w_dff_A_CyN3oALh9_0;
	wire w_dff_A_NuqozF7E7_0;
	wire w_dff_A_1IEEYlq61_0;
	wire w_dff_A_jGiIuj499_0;
	wire w_dff_A_bGbD4Y8e4_0;
	wire w_dff_A_pREiaToH1_0;
	wire w_dff_A_9fqtvgvi1_0;
	wire w_dff_A_k6cdTKzc3_0;
	wire w_dff_A_4MMsdCtT3_0;
	wire w_dff_A_kDXVf9032_0;
	wire w_dff_A_oCouwUys8_0;
	wire w_dff_A_Ecw3XE0C8_1;
	wire w_dff_A_JxtG2gM51_0;
	wire w_dff_A_w9givJGQ5_0;
	wire w_dff_A_BX5t45CH8_0;
	wire w_dff_A_eAeQP5g77_0;
	wire w_dff_A_dkTfI9qz8_0;
	wire w_dff_A_y4j5juJP0_0;
	wire w_dff_A_6D3O5RuW5_0;
	wire w_dff_A_8zl4laL25_0;
	wire w_dff_A_F9zbjyzh8_0;
	wire w_dff_A_fRURxQSj2_0;
	wire w_dff_A_ZcNOHpNk4_0;
	wire w_dff_A_Pyr9ZYRo9_0;
	wire w_dff_A_hvojzIHa4_0;
	wire w_dff_A_E8yhJQnZ7_0;
	wire w_dff_A_8GVBXo291_0;
	wire w_dff_A_9lKYjnjk7_0;
	wire w_dff_A_cmNluERk6_0;
	wire w_dff_A_CZQDbA8H0_0;
	wire w_dff_A_wQK9nt550_0;
	wire w_dff_A_G9kc5lVR6_0;
	wire w_dff_A_Augx0A7H8_0;
	wire w_dff_A_MsGYMzO90_0;
	wire w_dff_A_rzFpPzJV4_0;
	wire w_dff_A_E9msK8wW2_0;
	wire w_dff_A_r2Lmlu2r1_0;
	wire w_dff_A_V6c6oLjl9_0;
	wire w_dff_A_pCm67LpO3_0;
	wire w_dff_A_wznbd0EH2_0;
	wire w_dff_A_9z0AByg69_0;
	wire w_dff_A_gEiuKOGj2_0;
	wire w_dff_A_xArsL7LR1_0;
	wire w_dff_A_p6iOJAju7_0;
	wire w_dff_A_tadBGjSV2_0;
	wire w_dff_A_A14g1eR75_0;
	wire w_dff_A_3BrMdQ0f5_0;
	wire w_dff_A_XzfZhxu66_0;
	wire w_dff_A_uxlMMV2T6_0;
	wire w_dff_A_mkapjFNr2_1;
	wire w_dff_A_gseXjABl7_0;
	wire w_dff_A_VSopTJoF1_0;
	wire w_dff_A_M1BkhQtZ6_0;
	wire w_dff_A_5PH3PAnc6_0;
	wire w_dff_A_5St6i9pA1_0;
	wire w_dff_A_DaujxEGc1_0;
	wire w_dff_A_OeMst2Un4_0;
	wire w_dff_A_HAbOU5VZ0_0;
	wire w_dff_A_zZBKXntg1_0;
	wire w_dff_A_u9PKfo3T1_0;
	wire w_dff_A_p9LCjROE3_0;
	wire w_dff_A_9c6bRCCB5_0;
	wire w_dff_A_62APR6QZ6_0;
	wire w_dff_A_MGYQNllt8_0;
	wire w_dff_A_QL6RY0b14_0;
	wire w_dff_A_mMvxT7Yz4_0;
	wire w_dff_A_CwAxFP3j3_0;
	wire w_dff_A_jmiroCuE7_0;
	wire w_dff_A_eEITPnr53_0;
	wire w_dff_A_DVJWp4ud6_0;
	wire w_dff_A_XpqYFIWo5_0;
	wire w_dff_A_g3P4FDHU6_0;
	wire w_dff_A_Zl2UCqnZ8_0;
	wire w_dff_A_ExnCMEin5_0;
	wire w_dff_A_MbZyLN2u2_0;
	wire w_dff_A_OZJ01zsz1_0;
	wire w_dff_A_MQ7WdUvN5_0;
	wire w_dff_A_yAiHocCZ2_0;
	wire w_dff_A_JCq70if10_0;
	wire w_dff_A_wLat4gce2_0;
	wire w_dff_A_Dsfqz4gA9_0;
	wire w_dff_A_0JEkb5Ut9_0;
	wire w_dff_A_COggvmzL5_0;
	wire w_dff_A_Ap4Dv5kD4_0;
	wire w_dff_A_RBEDV1Rf6_0;
	wire w_dff_A_KQ4WqkKx5_0;
	wire w_dff_A_F62O6jpF7_0;
	wire w_dff_A_SAgjieT26_0;
	wire w_dff_A_JNSQA5WW0_1;
	wire w_dff_A_sZ2Ye7S04_0;
	wire w_dff_A_p9J2VSBu8_0;
	wire w_dff_A_fCUDzCgx7_0;
	wire w_dff_A_UxmXelcD8_0;
	wire w_dff_A_dd5dwjNi9_0;
	wire w_dff_A_IJyDPoxj6_0;
	wire w_dff_A_Ukr7kAib5_0;
	wire w_dff_A_t0MR3e8e7_0;
	wire w_dff_A_mZb1Kx5i2_0;
	wire w_dff_A_sbK9BLBZ5_0;
	wire w_dff_A_I68zm5vB6_0;
	wire w_dff_A_Zso0yqaY5_0;
	wire w_dff_A_CSt4kDh24_0;
	wire w_dff_A_uC9RWX2K2_0;
	wire w_dff_A_Pc6eUPN04_0;
	wire w_dff_A_tUeVAjnK3_0;
	wire w_dff_A_1MuqX2YZ2_0;
	wire w_dff_A_twvCwRQT9_0;
	wire w_dff_A_7x8xuhKI4_0;
	wire w_dff_A_ewI8G7jQ8_0;
	wire w_dff_A_ktRMidhS3_0;
	wire w_dff_A_rERIW63D6_0;
	wire w_dff_A_Y6T4ICtY3_0;
	wire w_dff_A_1TIdyplS2_0;
	wire w_dff_A_4rFqcHvh3_0;
	wire w_dff_A_0f0qnMpj7_0;
	wire w_dff_A_79ZePbnR8_0;
	wire w_dff_A_g5sNgMBQ3_0;
	wire w_dff_A_6jAGtIOk9_0;
	wire w_dff_A_vSpJVBrE1_0;
	wire w_dff_A_mYbgiXqX8_0;
	wire w_dff_A_bEvidwvA1_0;
	wire w_dff_A_46ntLdMS0_0;
	wire w_dff_A_V98IpRcV3_0;
	wire w_dff_A_a57WLguh3_0;
	wire w_dff_A_qWkNnZEb1_0;
	wire w_dff_A_zzpcdWs51_0;
	wire w_dff_A_bK1yUz2T7_0;
	wire w_dff_A_UcGMKMoa0_1;
	wire w_dff_A_Jx3pVlHg4_0;
	wire w_dff_A_EoD5PMn01_0;
	wire w_dff_A_zJgKbrJK3_0;
	wire w_dff_A_SXVwpqOM7_0;
	wire w_dff_A_0AU0VOUP1_0;
	wire w_dff_A_5jMvbd6v9_0;
	wire w_dff_A_oJQSa3TH1_0;
	wire w_dff_A_JEC6AGJ29_0;
	wire w_dff_A_4risWdAi4_0;
	wire w_dff_A_p7yvjMcI6_0;
	wire w_dff_A_QxRaRArh5_0;
	wire w_dff_A_1MaeLNCf7_0;
	wire w_dff_A_hJV1y4ok9_0;
	wire w_dff_A_Bpyenhtu7_0;
	wire w_dff_A_bMwFIHxA3_0;
	wire w_dff_A_7L91PiaT8_0;
	wire w_dff_A_ZHMStFjQ9_0;
	wire w_dff_A_HiyQfKje3_0;
	wire w_dff_A_t08A0Wh90_0;
	wire w_dff_A_yYxBmyyI7_0;
	wire w_dff_A_uHsWKiTq6_0;
	wire w_dff_A_COmVAiYt6_0;
	wire w_dff_A_OB4xrie35_0;
	wire w_dff_A_4cazQZu34_0;
	wire w_dff_A_Azxin5gJ9_0;
	wire w_dff_A_uNKUOqjj9_0;
	wire w_dff_A_nUDK1cDz3_0;
	wire w_dff_A_YKtJb5iH1_0;
	wire w_dff_A_AB1fkHal0_0;
	wire w_dff_A_YJKu4n7R1_0;
	wire w_dff_A_JQOtpg7T5_0;
	wire w_dff_A_2l7LCQqd5_0;
	wire w_dff_A_xLawbqg44_0;
	wire w_dff_A_TI0CfsI76_0;
	wire w_dff_A_TyRnyetE3_0;
	wire w_dff_A_EjvaFcqK0_0;
	wire w_dff_A_RImng3S02_0;
	wire w_dff_A_0zcSSwgI6_0;
	wire w_dff_A_l29pao1a2_2;
	wire w_dff_A_vpHsIN2M8_0;
	wire w_dff_A_twkstNKm7_0;
	wire w_dff_A_o8UYQHkv5_0;
	wire w_dff_A_Z72aivL71_0;
	wire w_dff_A_VR5xCiLY6_0;
	wire w_dff_A_puoj0En35_0;
	wire w_dff_A_ftHEnxS79_0;
	wire w_dff_A_CW0krvaF6_0;
	wire w_dff_A_trhOOQNj2_0;
	wire w_dff_A_onFXXuws4_0;
	wire w_dff_A_cvvdYd0z6_0;
	wire w_dff_A_qDjEyS7M6_0;
	wire w_dff_A_qHCHfUXE1_0;
	wire w_dff_A_RhaAMeBP5_0;
	wire w_dff_A_MbwJ5eIo9_0;
	wire w_dff_A_r595fPhb1_0;
	wire w_dff_A_aODRENxC7_0;
	wire w_dff_A_Y3mPe2o84_0;
	wire w_dff_A_LKkzhW2h4_0;
	wire w_dff_A_O1Uh8qCm5_0;
	wire w_dff_A_IMhJg36c7_0;
	wire w_dff_A_NS5V6sgc8_0;
	wire w_dff_A_ip84immA1_0;
	wire w_dff_A_1ua8GXzo3_0;
	wire w_dff_A_mVzlf2gk4_0;
	wire w_dff_A_eI88lScm7_0;
	wire w_dff_A_w4tfmbqf3_0;
	wire w_dff_A_TtIABepv9_0;
	wire w_dff_A_EJj0UGy71_0;
	wire w_dff_A_ZCSFIX2b7_0;
	wire w_dff_A_xPWT8kjR8_0;
	wire w_dff_A_IlJbGYVQ9_0;
	wire w_dff_A_7mNEW4CC9_0;
	wire w_dff_A_II3vq1OJ0_0;
	wire w_dff_A_KOVwRCJu8_0;
	wire w_dff_A_SeCEcx126_0;
	wire w_dff_A_fskGHtJ71_0;
	wire w_dff_A_f9BvEB0p2_1;
	wire w_dff_A_QmFN9ecY0_0;
	wire w_dff_A_ABvL59jj2_0;
	wire w_dff_A_2Q5aWDyp0_0;
	wire w_dff_A_G2h1cVhs3_0;
	wire w_dff_A_9x4m3eGD3_0;
	wire w_dff_A_QTuckQAp2_0;
	wire w_dff_A_ChHE3GpA4_0;
	wire w_dff_A_uL8ms4jz8_0;
	wire w_dff_A_rz2Tsc6i4_0;
	wire w_dff_A_4s3dByA95_0;
	wire w_dff_A_04nuj0MO6_0;
	wire w_dff_A_lq2F7Xmy0_0;
	wire w_dff_A_hayGb6pg4_0;
	wire w_dff_A_sGDSKULh9_0;
	wire w_dff_A_N6ev3BFD3_0;
	wire w_dff_A_8Oaw93Af3_0;
	wire w_dff_A_S4oO2WE52_0;
	wire w_dff_A_vdtiLAcA9_0;
	wire w_dff_A_OLhZKdKE8_0;
	wire w_dff_A_jnYdKqCs7_0;
	wire w_dff_A_skrNjDKt5_0;
	wire w_dff_A_PcC3T0l90_0;
	wire w_dff_A_eHZ51nIy2_0;
	wire w_dff_A_e7UtXRq43_0;
	wire w_dff_A_B5iqlsxA6_0;
	wire w_dff_A_UCla0D5N8_0;
	wire w_dff_A_AVUd1WYq7_0;
	wire w_dff_A_sWaSxgmF6_0;
	wire w_dff_A_JshhyMeG4_0;
	wire w_dff_A_WPCzSxIp7_0;
	wire w_dff_A_fRz2Ewyi3_0;
	wire w_dff_A_nNAPGyfd0_0;
	wire w_dff_A_n9nueMw50_0;
	wire w_dff_A_q3x932343_0;
	wire w_dff_A_mGOYjGEC3_0;
	wire w_dff_A_cVJigQ0M0_1;
	wire w_dff_A_UUcobrs82_0;
	wire w_dff_A_DK6Wrpyk9_0;
	wire w_dff_A_7G9uf8QO5_0;
	wire w_dff_A_nkDNo1se6_0;
	wire w_dff_A_h81KICLp8_0;
	wire w_dff_A_nioisLAD5_0;
	wire w_dff_A_LJlZtDij9_0;
	wire w_dff_A_813iFHv09_0;
	wire w_dff_A_axJ7XbcL9_0;
	wire w_dff_A_0oRzjyim8_0;
	wire w_dff_A_Vdx44zb02_0;
	wire w_dff_A_nMldML9W4_0;
	wire w_dff_A_kc4iEzfq2_0;
	wire w_dff_A_HeU802GO1_0;
	wire w_dff_A_xoKHy0wl1_0;
	wire w_dff_A_jneBexU33_0;
	wire w_dff_A_DZpTgcTD7_0;
	wire w_dff_A_kaSynU7e8_0;
	wire w_dff_A_AzYZCCN58_0;
	wire w_dff_A_GlViQ2a47_0;
	wire w_dff_A_DDb3mBxp7_0;
	wire w_dff_A_IWg0Q6zc7_0;
	wire w_dff_A_NafJUaX61_0;
	wire w_dff_A_MuXb125O4_0;
	wire w_dff_A_w8SPfYI32_0;
	wire w_dff_A_ctGLWZTc9_0;
	wire w_dff_A_RMUWSGP52_0;
	wire w_dff_A_9tM1MDuc0_0;
	wire w_dff_A_A7nEpr661_0;
	wire w_dff_A_VHpXnndZ9_0;
	wire w_dff_A_ooj0XJgm7_0;
	wire w_dff_A_vCu00N991_0;
	wire w_dff_A_HlqCQLAY6_0;
	wire w_dff_A_rg1a1AVl8_0;
	wire w_dff_A_7zVj4Qf74_0;
	wire w_dff_A_uXZKF6Yh3_1;
	wire w_dff_A_QAPZCd5D5_0;
	wire w_dff_A_wGjYtbn99_0;
	wire w_dff_A_p4seJZne1_0;
	wire w_dff_A_dzeNiATj5_0;
	wire w_dff_A_NzNxO6yS0_0;
	wire w_dff_A_ABdOXtSb4_0;
	wire w_dff_A_BE4Jz0VU6_0;
	wire w_dff_A_hpHsj7jz7_0;
	wire w_dff_A_6NEzPVXR5_0;
	wire w_dff_A_UFzQSGYo5_0;
	wire w_dff_A_CzELws3Q1_0;
	wire w_dff_A_lu92C5VG8_0;
	wire w_dff_A_fVmzrn5z1_0;
	wire w_dff_A_FjVfwBkm4_0;
	wire w_dff_A_2CaVv1wK5_0;
	wire w_dff_A_jTZG1E9T2_0;
	wire w_dff_A_LgsP8qEz8_0;
	wire w_dff_A_cPj50RB71_0;
	wire w_dff_A_9BFB27r18_0;
	wire w_dff_A_pMPG5zP03_0;
	wire w_dff_A_XaLre3FV2_0;
	wire w_dff_A_6Ei26ZAL3_0;
	wire w_dff_A_cKqrvQBg8_0;
	wire w_dff_A_HJRmcQFq0_0;
	wire w_dff_A_FQcqCSdl9_0;
	wire w_dff_A_OvIeQQXb0_0;
	wire w_dff_A_qXxicUeF3_0;
	wire w_dff_A_ms99laM27_0;
	wire w_dff_A_OjMdN8nn0_0;
	wire w_dff_A_SSDbt0Ut6_0;
	wire w_dff_A_gZ5rN5JU7_0;
	wire w_dff_A_1KAVeFYD7_0;
	wire w_dff_A_oG7cPQNU3_0;
	wire w_dff_A_A0RuoFMe1_0;
	wire w_dff_A_SzsJbbxU2_0;
	wire w_dff_A_vLRVPHpJ9_1;
	wire w_dff_A_pETu6NWu8_0;
	wire w_dff_A_0q4VzV568_0;
	wire w_dff_A_LCWWeUNO3_0;
	wire w_dff_A_x6jMIy466_0;
	wire w_dff_A_fKMs039R1_0;
	wire w_dff_A_ZtjpM78x7_0;
	wire w_dff_A_l4xmYpXr7_0;
	wire w_dff_A_90B53fqI6_0;
	wire w_dff_A_VorGZjvp6_0;
	wire w_dff_A_MF5KCvsH8_0;
	wire w_dff_A_3KFt32vo5_0;
	wire w_dff_A_Bygal0ww1_0;
	wire w_dff_A_OLmDZgpm8_0;
	wire w_dff_A_WFWLv4Ef7_0;
	wire w_dff_A_yCfeM25i3_0;
	wire w_dff_A_RafLgjDR8_0;
	wire w_dff_A_VngPkwI53_0;
	wire w_dff_A_vsN2pBpa8_0;
	wire w_dff_A_8nALCqNr5_0;
	wire w_dff_A_bUTpaOBi0_0;
	wire w_dff_A_jBOyfPDn4_0;
	wire w_dff_A_LvD3dYgc2_0;
	wire w_dff_A_ze9uco4J0_0;
	wire w_dff_A_1mImsz3t5_0;
	wire w_dff_A_zdcSQLJZ4_0;
	wire w_dff_A_CSmIodxh4_0;
	wire w_dff_A_QauGlLGA8_0;
	wire w_dff_A_ajnPqiCO0_0;
	wire w_dff_A_VGbi1yME3_0;
	wire w_dff_A_JNv0kTSU6_0;
	wire w_dff_A_larRg07u8_0;
	wire w_dff_A_CBsy12Sx9_0;
	wire w_dff_A_Txxc89Ca1_0;
	wire w_dff_A_ZeCSr41v6_0;
	wire w_dff_A_BviXlD0x7_0;
	wire w_dff_A_UmRpndW02_1;
	wire w_dff_A_g6aYWzKz7_0;
	wire w_dff_A_iNeR9I6u7_0;
	wire w_dff_A_SgN08v1v3_0;
	wire w_dff_A_rINHG92u2_0;
	wire w_dff_A_lNY9aq9L3_0;
	wire w_dff_A_PU6oLifR3_0;
	wire w_dff_A_PplyFSli5_0;
	wire w_dff_A_7Ie371jD9_0;
	wire w_dff_A_tQiVhEhr4_0;
	wire w_dff_A_ECIM6ThG5_0;
	wire w_dff_A_lxKSkcwZ0_0;
	wire w_dff_A_7idhb0VO5_0;
	wire w_dff_A_CYtfvawb0_0;
	wire w_dff_A_dC8Rr2P03_0;
	wire w_dff_A_7QABMPlQ5_0;
	wire w_dff_A_36BMpCoG5_0;
	wire w_dff_A_s1jtSIvt7_0;
	wire w_dff_A_gnEyxGXA9_0;
	wire w_dff_A_4mUNCGDX5_0;
	wire w_dff_A_EerkGR6q7_0;
	wire w_dff_A_jKNmD0wk7_0;
	wire w_dff_A_cFHSo8kd3_0;
	wire w_dff_A_5hlrKPv12_0;
	wire w_dff_A_HzBBmX0l4_0;
	wire w_dff_A_P24sqcHi5_0;
	wire w_dff_A_GtbN2OiQ3_0;
	wire w_dff_A_AVkXWHZx7_0;
	wire w_dff_A_156IjwjA0_0;
	wire w_dff_A_13QnXjkB8_0;
	wire w_dff_A_0D7KPyRq7_0;
	wire w_dff_A_8JSeBPHl2_0;
	wire w_dff_A_Jkjwe1l57_0;
	wire w_dff_A_yOBfpf2J7_0;
	wire w_dff_A_8zlEVCJZ9_0;
	wire w_dff_A_XZm1WecU4_0;
	wire w_dff_A_wXxqaB6A9_0;
	wire w_dff_A_AtyoT8ZO0_0;
	wire w_dff_A_olSL7hVn3_0;
	wire w_dff_A_GvhcWMRm2_1;
	wire w_dff_A_8Nfw95BS7_0;
	wire w_dff_A_sYlMZort9_0;
	wire w_dff_A_LPUJtTLt0_0;
	wire w_dff_A_Mu5BzN2u8_0;
	wire w_dff_A_8znLl8dS8_0;
	wire w_dff_A_HZ15V9MR7_0;
	wire w_dff_A_HXvb78Tb1_0;
	wire w_dff_A_NhK5mDNZ6_0;
	wire w_dff_A_7LhMwXib8_0;
	wire w_dff_A_69w0CmSt1_0;
	wire w_dff_A_0qmWonwJ3_0;
	wire w_dff_A_asimPkSb1_0;
	wire w_dff_A_4eGrZ8K15_0;
	wire w_dff_A_8QLY8DaK4_0;
	wire w_dff_A_EF3nEqlO5_0;
	wire w_dff_A_IqDXQpKH1_0;
	wire w_dff_A_GIZWvFyN2_0;
	wire w_dff_A_HV7wdW6r1_0;
	wire w_dff_A_X6gXpop32_0;
	wire w_dff_A_d0h6NpRa9_0;
	wire w_dff_A_RDD70BOP3_0;
	wire w_dff_A_bHDwJCfG7_0;
	wire w_dff_A_YN49zphR2_0;
	wire w_dff_A_ch18PvVw0_0;
	wire w_dff_A_YowinJjM0_0;
	wire w_dff_A_nifW53gz9_0;
	wire w_dff_A_pzh1n70A3_0;
	wire w_dff_A_MfXwBtvq8_0;
	wire w_dff_A_teoyOoBm3_0;
	wire w_dff_A_RF3bfCx54_0;
	wire w_dff_A_N9sllnDa5_0;
	wire w_dff_A_z4GtcDGJ2_0;
	wire w_dff_A_3iHvKG7B1_0;
	wire w_dff_A_4k6m9DqR5_0;
	wire w_dff_A_B1CqK4mr5_0;
	wire w_dff_A_ebVxtHs96_0;
	wire w_dff_A_StI7oTcp7_0;
	wire w_dff_A_u4outPN43_0;
	wire w_dff_A_shAXd2VJ7_2;
	wire w_dff_A_sBOX5pMf4_0;
	wire w_dff_A_d8gA6SAU7_0;
	wire w_dff_A_POQLqnuM1_0;
	wire w_dff_A_eSQrbb492_0;
	wire w_dff_A_8Ea9HJjE5_0;
	wire w_dff_A_Yixjxbt06_0;
	wire w_dff_A_vXgtixgr3_0;
	wire w_dff_A_psz6UQtf2_0;
	wire w_dff_A_4tNNQwRC4_0;
	wire w_dff_A_qhHSbbHM5_0;
	wire w_dff_A_wFFAiIgn5_0;
	wire w_dff_A_axaXoooe0_0;
	wire w_dff_A_AmH0nBOK3_0;
	wire w_dff_A_mj3N1yxe0_0;
	wire w_dff_A_cyfgnMUv7_0;
	wire w_dff_A_ZptR4TQq8_0;
	wire w_dff_A_ZK6uJmzb0_0;
	wire w_dff_A_VZSmSLFH6_0;
	wire w_dff_A_GmlhfgGs2_0;
	wire w_dff_A_87i4wdCQ9_0;
	wire w_dff_A_5jRbM2bp8_0;
	wire w_dff_A_kv8hPPfP8_0;
	wire w_dff_A_CHkdAiIW0_0;
	wire w_dff_A_BzQBSkrh8_0;
	wire w_dff_A_lKYiOSZv8_0;
	wire w_dff_A_rB1y8qcf4_0;
	wire w_dff_A_5jWupdvD4_0;
	wire w_dff_A_557gGvBh8_0;
	wire w_dff_A_GhHtLrJ53_0;
	wire w_dff_A_F8mbicrI9_0;
	wire w_dff_A_6USjyokI4_0;
	wire w_dff_A_jLUQKHfc6_0;
	wire w_dff_A_L5JoTiLQ0_0;
	wire w_dff_A_uFMOIDk74_0;
	wire w_dff_A_TD9z5fXV5_0;
	wire w_dff_A_gOSHElLu0_0;
	wire w_dff_A_80dpXEcR8_1;
	wire w_dff_A_QtRn1iNZ1_0;
	wire w_dff_A_6f9MzD7l5_0;
	wire w_dff_A_pyRvFWsR5_0;
	wire w_dff_A_iVauyqfL4_0;
	wire w_dff_A_ivkVRNC56_0;
	wire w_dff_A_UlF54cb87_0;
	wire w_dff_A_tkhvg9TS1_0;
	wire w_dff_A_10xolld75_0;
	wire w_dff_A_EVz7tDW14_0;
	wire w_dff_A_iax3o9Jk5_0;
	wire w_dff_A_ULKJWwH77_0;
	wire w_dff_A_nrke1Mab4_0;
	wire w_dff_A_9oXUnIOz7_0;
	wire w_dff_A_8LNW5BtM0_0;
	wire w_dff_A_TK7FDZtd3_0;
	wire w_dff_A_nNm2M1T17_0;
	wire w_dff_A_ikf2zKF11_0;
	wire w_dff_A_VFjj4J008_0;
	wire w_dff_A_Uhod3cOY3_0;
	wire w_dff_A_zpKaUDB92_0;
	wire w_dff_A_LGuYaKgw8_0;
	wire w_dff_A_UlWOZn0M5_0;
	wire w_dff_A_hIFWfd6U2_0;
	wire w_dff_A_WBICRSrf0_0;
	wire w_dff_A_MlfVKyUe7_0;
	wire w_dff_A_O1RgAoCZ5_0;
	wire w_dff_A_9t05lWiJ1_0;
	wire w_dff_A_8e3Ab73a8_0;
	wire w_dff_A_IOr5R2l06_0;
	wire w_dff_A_OhjlDZ687_0;
	wire w_dff_A_PVC1HXKf8_0;
	wire w_dff_A_BhGFb2IV8_0;
	wire w_dff_A_BeLrqKEh3_0;
	wire w_dff_A_3DQjD6g93_0;
	wire w_dff_A_9Uq65EFi0_0;
	wire w_dff_A_AniK33Dp4_0;
	wire w_dff_A_gJN29yv56_0;
	wire w_dff_A_2ffOjGSw0_2;
	wire w_dff_A_lZwHf6R40_0;
	wire w_dff_A_y4g9cm1v4_0;
	wire w_dff_A_pvsCAZDH1_0;
	wire w_dff_A_SBvcXEsb3_0;
	wire w_dff_A_KeUUZKkh9_0;
	wire w_dff_A_D0XsJf9x0_0;
	wire w_dff_A_LO9zKj3B5_0;
	wire w_dff_A_RsJhGyoV5_0;
	wire w_dff_A_9DeQYJjo2_0;
	wire w_dff_A_B2c7gVPS9_0;
	wire w_dff_A_UrI4DLaB7_0;
	wire w_dff_A_Z5WxMyim5_0;
	wire w_dff_A_zQC6m5t67_0;
	wire w_dff_A_fgLj68N53_0;
	wire w_dff_A_qbGJPf7C7_0;
	wire w_dff_A_SpMBQ90i0_0;
	wire w_dff_A_w6PG7JqV9_0;
	wire w_dff_A_rUAgz0BP6_0;
	wire w_dff_A_lTS3vKVH0_0;
	wire w_dff_A_A5gke3At5_0;
	wire w_dff_A_ZtR7t5VX8_0;
	wire w_dff_A_ZDWOUPiC8_0;
	wire w_dff_A_hoafLdX80_0;
	wire w_dff_A_5racRmi43_0;
	wire w_dff_A_ijAeR4rh3_0;
	wire w_dff_A_ImcgR7xm9_0;
	wire w_dff_A_Sd58F3UK2_0;
	wire w_dff_A_cQ8qT2dE3_0;
	wire w_dff_A_G3kR2pin3_0;
	wire w_dff_A_E4NHioB47_0;
	wire w_dff_A_CptaiCnM7_0;
	wire w_dff_A_9TQb8tTY9_0;
	wire w_dff_A_tyy4Ebdq7_0;
	wire w_dff_A_xxyNTzB67_0;
	wire w_dff_A_BJDi9gcw9_0;
	wire w_dff_A_I9mtoSGP1_0;
	wire w_dff_A_5CWJDb799_2;
	wire w_dff_A_gBIXloda6_0;
	wire w_dff_A_lmqIViUF0_0;
	wire w_dff_A_JSXejjHQ0_0;
	wire w_dff_A_d7GRBcPd6_0;
	wire w_dff_A_lHw19Lfd9_0;
	wire w_dff_A_1enBGeNJ6_0;
	wire w_dff_A_T9eJqdRv8_0;
	wire w_dff_A_RvoX3PVw5_0;
	wire w_dff_A_sAWPyZ7B9_0;
	wire w_dff_A_6bQx5k2h2_0;
	wire w_dff_A_MIMuAJRc2_0;
	wire w_dff_A_G7bHtZWK7_0;
	wire w_dff_A_VI3Fp35F9_0;
	wire w_dff_A_bk9s3Rj58_0;
	wire w_dff_A_JWuAjjag5_0;
	wire w_dff_A_TXvXQldr2_0;
	wire w_dff_A_fwdvcNeG0_0;
	wire w_dff_A_yAH4vpjM2_0;
	wire w_dff_A_wMQptCx18_0;
	wire w_dff_A_amkVk9Oq1_0;
	wire w_dff_A_j40ug4rP7_0;
	wire w_dff_A_MBybOkkQ0_0;
	wire w_dff_A_v7DppBZp6_0;
	wire w_dff_A_Zb9ekEIH1_0;
	wire w_dff_A_v48GulAq7_0;
	wire w_dff_A_vteSKWGg3_0;
	wire w_dff_A_TTWLxi272_0;
	wire w_dff_A_wRXPZGqq9_0;
	wire w_dff_A_hYG6VFTD3_0;
	wire w_dff_A_6UpMiI3Z2_0;
	wire w_dff_A_pCuZM0lV5_0;
	wire w_dff_A_rKqX1lhP6_0;
	wire w_dff_A_4scZZCVe2_0;
	wire w_dff_A_KuyJyPJT5_0;
	wire w_dff_A_NYKCgtdD7_0;
	wire w_dff_A_5UJxVmwi0_1;
	wire w_dff_A_b2XBNgqA6_0;
	wire w_dff_A_eEgdHU7Q1_0;
	wire w_dff_A_OPwWvTME9_0;
	wire w_dff_A_XxpWVlXX4_0;
	wire w_dff_A_M4ISSJIz9_0;
	wire w_dff_A_sR6jGFbd4_0;
	wire w_dff_A_F7t6vG9k5_0;
	wire w_dff_A_YTEGXAvm4_0;
	wire w_dff_A_qluAPOsF2_0;
	wire w_dff_A_HA1Jo9N09_0;
	wire w_dff_A_R1xys3UN0_0;
	wire w_dff_A_YuGT2vLL5_0;
	wire w_dff_A_yhE1oluh6_0;
	wire w_dff_A_57palikL4_0;
	wire w_dff_A_nRMANwxx1_0;
	wire w_dff_A_Ci6ruBFk3_0;
	wire w_dff_A_wI9VE5U23_0;
	wire w_dff_A_UOulhVea0_0;
	wire w_dff_A_KfzX7r6E1_0;
	wire w_dff_A_zitRS7j84_0;
	wire w_dff_A_m58o1jfZ3_0;
	wire w_dff_A_oTpXEnrE9_0;
	wire w_dff_A_ve2dmMk57_0;
	wire w_dff_A_CFovSXlD4_0;
	wire w_dff_A_63Jd9I6I5_0;
	wire w_dff_A_72UBYXcW8_0;
	wire w_dff_A_VMcvQswL1_0;
	wire w_dff_A_gIB7J3tz4_0;
	wire w_dff_A_pUXQxgje3_0;
	wire w_dff_A_aVMdw0M67_0;
	wire w_dff_A_rYW2m9Lx6_0;
	wire w_dff_A_5SGfGcPQ0_0;
	wire w_dff_A_Brk5I6Kr5_0;
	wire w_dff_A_cChG1fMn0_0;
	wire w_dff_A_z1L8L5Ah3_0;
	wire w_dff_A_THGPqgYF5_0;
	wire w_dff_A_UkS5GTox6_0;
	wire w_dff_A_LYTWwnQT3_2;
	wire w_dff_A_rOhaXiQu9_0;
	wire w_dff_A_qSnjebqh5_0;
	wire w_dff_A_axO0PiAe0_0;
	wire w_dff_A_qag10fA49_0;
	wire w_dff_A_Jfcy6ivk8_0;
	wire w_dff_A_e9npHuAR1_0;
	wire w_dff_A_M4OBSOlH5_0;
	wire w_dff_A_sp0YFyoC1_0;
	wire w_dff_A_npVOn1jy5_0;
	wire w_dff_A_RzB7xMFP5_0;
	wire w_dff_A_kS9mjGrh5_0;
	wire w_dff_A_UWfax2q97_0;
	wire w_dff_A_PZlZX5CP8_0;
	wire w_dff_A_6k2aV4Wv5_0;
	wire w_dff_A_x7H4R5ju3_0;
	wire w_dff_A_JWp8zvp55_0;
	wire w_dff_A_U4U6aH6s4_0;
	wire w_dff_A_4ZuLP4ev6_0;
	wire w_dff_A_1OYAlXSC9_0;
	wire w_dff_A_7RyYZd4j5_0;
	wire w_dff_A_7CBFCoj75_0;
	wire w_dff_A_xtSKDinO3_0;
	wire w_dff_A_YBmOpkG23_0;
	wire w_dff_A_njEXYHq94_0;
	wire w_dff_A_l9zCHjn00_0;
	wire w_dff_A_y6mXuzjy1_0;
	wire w_dff_A_SqhIIYuN3_0;
	wire w_dff_A_Fy68E4ri0_0;
	wire w_dff_A_MMhPxFZC5_0;
	wire w_dff_A_5ICq8oAh5_0;
	wire w_dff_A_cSWnvPqz8_0;
	wire w_dff_A_tTnXYDlF1_0;
	wire w_dff_A_AxbIMWhd7_0;
	wire w_dff_A_JtGuUzYo4_0;
	wire w_dff_A_XXnkcJya1_0;
	wire w_dff_A_v6D1FION8_1;
	wire w_dff_A_WXnqrcDo0_0;
	wire w_dff_A_h4wWoAuY3_0;
	wire w_dff_A_J2Y6GuVK3_0;
	wire w_dff_A_GrZzI1TX9_0;
	wire w_dff_A_oAmrXrWR6_0;
	wire w_dff_A_vz6SqLEs1_0;
	wire w_dff_A_riF2gTTT2_0;
	wire w_dff_A_txUkHtJJ7_0;
	wire w_dff_A_tfPqtxZD4_0;
	wire w_dff_A_GqLnxeAP1_0;
	wire w_dff_A_a3qliUqZ3_0;
	wire w_dff_A_YsXibD2e5_0;
	wire w_dff_A_jxRaui4Z3_0;
	wire w_dff_A_UXIeOfXk5_0;
	wire w_dff_A_QXgHYmff0_0;
	wire w_dff_A_HchAHDuA6_0;
	wire w_dff_A_FiyQ8NZB0_0;
	wire w_dff_A_85hrb3iP2_0;
	wire w_dff_A_9tsud5Bl6_0;
	wire w_dff_A_wZehHiKb2_0;
	wire w_dff_A_1Oqsl1bb5_0;
	wire w_dff_A_oflB3tYa7_0;
	wire w_dff_A_asaIc2GR5_0;
	wire w_dff_A_6tFU48pa8_0;
	wire w_dff_A_A77uKbXu1_0;
	wire w_dff_A_uplEs2uz3_0;
	wire w_dff_A_l7IEkgS81_0;
	wire w_dff_A_HHM2aAnN1_0;
	wire w_dff_A_K3LEQtDj6_0;
	wire w_dff_A_bk1vyzJA0_0;
	wire w_dff_A_ZthzvxHl9_0;
	wire w_dff_A_pIUJ1OB06_0;
	wire w_dff_A_5zKAxaVt0_0;
	wire w_dff_A_1OuSgU3z5_0;
	wire w_dff_A_FD6u7nH66_0;
	wire w_dff_A_VmfczGuC8_0;
	wire w_dff_A_6j1uDAKw2_0;
	wire w_dff_A_yULD7g5r5_0;
	wire w_dff_A_6JNnbqa23_2;
	wire w_dff_A_TgSBmCTr9_0;
	wire w_dff_A_nsEkwB1u2_0;
	wire w_dff_A_xENo23u41_0;
	wire w_dff_A_J1Wq44AT9_0;
	wire w_dff_A_WwNDomRU8_0;
	wire w_dff_A_MZuE6uKN3_0;
	wire w_dff_A_uDcMwWqz3_0;
	wire w_dff_A_jnpnw1D61_0;
	wire w_dff_A_tJ1NdhgQ2_0;
	wire w_dff_A_iyNZ2jFh6_0;
	wire w_dff_A_lbjLwgey2_0;
	wire w_dff_A_UMBV82v74_0;
	wire w_dff_A_mboFH9Xs4_0;
	wire w_dff_A_NU65Fn1J5_0;
	wire w_dff_A_evzEM4tN1_0;
	wire w_dff_A_UbO1NeX40_0;
	wire w_dff_A_UmRaH5YV2_0;
	wire w_dff_A_njncPKZm2_0;
	wire w_dff_A_RcIDBfhq2_0;
	wire w_dff_A_64X2WlhV8_0;
	wire w_dff_A_j9qVIGQX3_0;
	wire w_dff_A_y4Cspc1X9_0;
	wire w_dff_A_bi8BWD2L9_0;
	wire w_dff_A_tpnaq9my9_0;
	wire w_dff_A_uXa5h7pz6_0;
	wire w_dff_A_byOiI9Mn9_0;
	wire w_dff_A_rCz93Nd91_0;
	wire w_dff_A_JJJQY4Cb6_0;
	wire w_dff_A_0LPf6fYh5_0;
	wire w_dff_A_hrYBhWcf5_0;
	wire w_dff_A_qrCIzEHB0_0;
	wire w_dff_A_uIzUog2C5_0;
	wire w_dff_A_Da6qkFV23_0;
	wire w_dff_A_2BUrEj0k5_0;
	wire w_dff_A_75b2Pduh5_0;
	wire w_dff_A_YFaS9lDM2_0;
	wire w_dff_A_nnznEvcV8_0;
	wire w_dff_A_JUhLnoel6_2;
	wire w_dff_A_YIPQoqhU6_0;
	wire w_dff_A_xU9CMkso1_0;
	wire w_dff_A_fWTD6whD3_0;
	wire w_dff_A_WwJWWjDG7_0;
	wire w_dff_A_WUQ9TBw92_0;
	wire w_dff_A_Rmjp52Px5_0;
	wire w_dff_A_7HILhU292_0;
	wire w_dff_A_pB5TzMQF2_0;
	wire w_dff_A_5WNYiVIZ8_0;
	wire w_dff_A_r269STCO2_0;
	wire w_dff_A_t7zpBKCr2_0;
	wire w_dff_A_c8nFuvde7_0;
	wire w_dff_A_steTrupJ0_0;
	wire w_dff_A_sHvWjVfY7_0;
	wire w_dff_A_3qGhr6OA7_0;
	wire w_dff_A_L2wcn2YN5_0;
	wire w_dff_A_S7Ay9VY61_0;
	wire w_dff_A_HFCc6Y289_0;
	wire w_dff_A_vz9gJvBL0_0;
	wire w_dff_A_OgeEnrSc8_0;
	wire w_dff_A_DhQvmmJb6_0;
	wire w_dff_A_yWxvpk0L9_0;
	wire w_dff_A_LeDvghwO5_0;
	wire w_dff_A_uAscGIOG7_0;
	wire w_dff_A_2fGdQq3H6_0;
	wire w_dff_A_OOpz2K8o9_0;
	wire w_dff_A_IsIB4EQA3_0;
	wire w_dff_A_8Ch04RuM5_0;
	wire w_dff_A_HffPPdwN1_0;
	wire w_dff_A_U6TSY54Z8_0;
	wire w_dff_A_wp0QpJAL5_0;
	wire w_dff_A_UzUYjMgM6_0;
	wire w_dff_A_WgdesOxS6_2;
	wire w_dff_A_0MAjtAZX9_0;
	wire w_dff_A_XnWGpai63_0;
	wire w_dff_A_uPiXm35k8_0;
	wire w_dff_A_Jpk3n4926_0;
	wire w_dff_A_MiuRKQMd9_0;
	wire w_dff_A_h8e3CzGx6_0;
	wire w_dff_A_JjFLABj79_0;
	wire w_dff_A_iGD8WHOb0_0;
	wire w_dff_A_4rCrF3xX4_0;
	wire w_dff_A_6dZOUxLq7_0;
	wire w_dff_A_gVGYXbAZ9_2;
	wire w_dff_A_NqrjpIF95_0;
	wire w_dff_A_HNivIQsl8_0;
	wire w_dff_A_QY9Wrn8O2_0;
	wire w_dff_A_TuTty8EX9_0;
	wire w_dff_A_LX2u7u419_0;
	wire w_dff_A_yAKUWmNi4_0;
	wire w_dff_A_7HlLi65N3_0;
	wire w_dff_A_qsajmEeY3_0;
	wire w_dff_A_J8pd6cwc7_0;
	wire w_dff_A_52ewoE7D6_0;
	wire w_dff_A_hPnAfq4F4_2;
	wire w_dff_A_iNwMUUHK5_0;
	wire w_dff_A_PFOM2LhJ2_0;
	wire w_dff_A_nWiicRqs2_0;
	wire w_dff_A_rnXX74dU7_0;
	wire w_dff_A_a49ATBdq9_0;
	wire w_dff_A_xbkIkvNl6_0;
	wire w_dff_A_APefuJA21_0;
	wire w_dff_A_r4f54s5A3_0;
	wire w_dff_A_heXjPChd8_0;
	wire w_dff_A_Vz7q3ErZ5_0;
	wire w_dff_A_1OtQR8rD3_0;
	wire w_dff_A_MIaF2AKB6_0;
	wire w_dff_A_nGmhZ0yO2_0;
	wire w_dff_A_EdCsBd2c5_0;
	wire w_dff_A_T4b63vDR7_0;
	wire w_dff_A_A1kwbq6i9_0;
	wire w_dff_A_QY6wIL7V5_0;
	wire w_dff_A_oyuiGHus1_0;
	wire w_dff_A_FoXPssr27_0;
	wire w_dff_A_L2IfLhs72_0;
	wire w_dff_A_chT3XV4f0_0;
	wire w_dff_A_fumqalSS2_0;
	wire w_dff_A_2nnZdTm25_0;
	wire w_dff_A_2wIBugvy5_0;
	wire w_dff_A_gTjHNFqz8_2;
	wire w_dff_A_WKNUtcIs5_0;
	wire w_dff_A_rbcDPmp47_0;
	wire w_dff_A_Wn738bAv0_0;
	wire w_dff_A_tevt4oG43_0;
	wire w_dff_A_gMkcfKNc5_0;
	wire w_dff_A_hA6kEm0g5_0;
	wire w_dff_A_n20VkMtD0_0;
	wire w_dff_A_HeVyyHWm8_0;
	wire w_dff_A_OEhLT8dJ8_0;
	wire w_dff_A_QxwFQzQX8_0;
	wire w_dff_A_u5vFU4tv9_0;
	wire w_dff_A_LiReZLmP4_0;
	wire w_dff_A_Vlzubrbv1_0;
	wire w_dff_A_h0zZEJrs3_0;
	wire w_dff_A_7VuxU29p2_0;
	wire w_dff_A_lKhtrzhY2_0;
	wire w_dff_A_TmBXw6hR3_0;
	wire w_dff_A_peZAriNm4_0;
	wire w_dff_A_xZMnHIwy8_0;
	wire w_dff_A_4uGXzQWa7_0;
	wire w_dff_A_Wyp9HWKV7_0;
	wire w_dff_A_MAcM2TRw3_0;
	wire w_dff_A_lwhkvxhm6_0;
	wire w_dff_A_5wo7rnwH5_0;
	wire w_dff_A_CYQWdov97_0;
	wire w_dff_A_z7yc9I0i3_0;
	wire w_dff_A_5B1bkyF47_2;
	wire w_dff_A_Ttn95e517_0;
	wire w_dff_A_8t703pIG5_0;
	wire w_dff_A_qUGBXbCV2_0;
	wire w_dff_A_L8C51wfk8_0;
	wire w_dff_A_sJCoUQNH1_0;
	wire w_dff_A_GmKIpH9Y4_0;
	wire w_dff_A_rNfIFAE02_0;
	wire w_dff_A_4f4qySzM1_0;
	wire w_dff_A_3ncSnTUK7_0;
	wire w_dff_A_2eEKXkb91_0;
	wire w_dff_A_MyHPrs2b8_0;
	wire w_dff_A_5VaeJNyz4_0;
	wire w_dff_A_h2PRlNUO8_0;
	wire w_dff_A_LUECO1XC8_0;
	wire w_dff_A_vnvenVbj8_0;
	wire w_dff_A_qhYYZH6r5_0;
	wire w_dff_A_nT7D9dZC8_0;
	wire w_dff_A_EX1eb4ry4_0;
	wire w_dff_A_lk9Gz33w6_0;
	wire w_dff_A_RcZ9vyPH6_0;
	wire w_dff_A_5XM4gxYI7_0;
	wire w_dff_A_nj0FVd7u8_0;
	wire w_dff_A_UFeAFPWr9_0;
	wire w_dff_A_B9QL6Qe05_0;
	wire w_dff_A_ped9jlaL8_0;
	wire w_dff_A_IokUSfhx5_0;
	wire w_dff_A_b6l6bhqQ5_0;
	wire w_dff_A_gIFno2YV5_0;
	wire w_dff_A_zTDeMC165_0;
	wire w_dff_A_fpenTOu76_2;
	wire w_dff_A_cwWDxqXY1_0;
	wire w_dff_A_CAivFeWN1_0;
	wire w_dff_A_5BBLyt4O1_0;
	wire w_dff_A_PuUG3zsC7_0;
	wire w_dff_A_LscEx0BE1_0;
	wire w_dff_A_7GqgwZiS1_0;
	wire w_dff_A_v8dGGnxG1_0;
	wire w_dff_A_6jUbPnNn8_0;
	wire w_dff_A_jWCE1zxJ0_0;
	wire w_dff_A_djldMywr3_0;
	wire w_dff_A_H2nKMvgE4_0;
	wire w_dff_A_5eLdNyu16_0;
	wire w_dff_A_DLAr7g077_0;
	wire w_dff_A_HlNsc1Mn2_0;
	wire w_dff_A_CA924rQb5_0;
	wire w_dff_A_IhlIqXHJ2_0;
	wire w_dff_A_GtW6pevU5_0;
	wire w_dff_A_AT9S9VJt0_0;
	wire w_dff_A_wKFIr6Cp0_0;
	wire w_dff_A_dDURwMH97_0;
	wire w_dff_A_2RcdRk0R1_0;
	wire w_dff_A_uR8sQkJh2_0;
	wire w_dff_A_aVhbpkvT9_0;
	wire w_dff_A_tGUeM6AL7_0;
	wire w_dff_A_JGTVUj4L7_0;
	wire w_dff_A_5YcxzyGN2_0;
	wire w_dff_A_MNdxUWzQ8_0;
	wire w_dff_A_yF8MwC7r1_0;
	wire w_dff_A_AMEMdVHP1_0;
	wire w_dff_A_ttfj0vH04_0;
	wire w_dff_A_TNQcEwwd4_2;
	wire w_dff_A_RRZKL7iL4_0;
	wire w_dff_A_3P5NaF2r5_0;
	wire w_dff_A_YonoLV990_0;
	wire w_dff_A_oHh0BOtM0_0;
	wire w_dff_A_3nrLiEVZ3_0;
	wire w_dff_A_RIjcep6Q8_0;
	wire w_dff_A_g23pRVwW7_0;
	wire w_dff_A_neoHDwvD0_0;
	wire w_dff_A_ZISIHtAJ1_0;
	wire w_dff_A_qlxHZB3k5_0;
	wire w_dff_A_nLYwuqj32_0;
	wire w_dff_A_qSlaXN8l8_0;
	wire w_dff_A_itfXPfYC3_0;
	wire w_dff_A_vwKU9xyl8_0;
	wire w_dff_A_1DnrtLmJ0_0;
	wire w_dff_A_HZeatMJE7_0;
	wire w_dff_A_4xjDzBpk8_0;
	wire w_dff_A_Wfi1tSMF9_0;
	wire w_dff_A_4arLJuD57_0;
	wire w_dff_A_RCtQWRw62_2;
	wire w_dff_A_wcCPGPVJ7_0;
	wire w_dff_A_YvBnnsTX1_0;
	wire w_dff_A_2S5E8xlm4_0;
	wire w_dff_A_F3SD8t3w8_0;
	wire w_dff_A_CozWiyfC4_0;
	wire w_dff_A_pkWkkBzf1_0;
	wire w_dff_A_ROpv3ED38_0;
	wire w_dff_A_9gQuaPxf8_0;
	wire w_dff_A_LH8pqbTX2_0;
	wire w_dff_A_x10gWTsH5_0;
	wire w_dff_A_TxYwJokZ6_0;
	wire w_dff_A_cN0aZ28w5_0;
	wire w_dff_A_s8ahpQih9_0;
	wire w_dff_A_qs21yKio3_0;
	wire w_dff_A_6o22pCvI9_0;
	wire w_dff_A_pEagct3R1_0;
	wire w_dff_A_ItHBpcHd1_0;
	wire w_dff_A_hR0gFTZn6_0;
	wire w_dff_A_VP3xdPTV0_0;
	wire w_dff_A_pqvkgzNJ8_0;
	wire w_dff_A_WPg6b8Tt1_0;
	wire w_dff_A_OwLg3vyW3_2;
	wire w_dff_A_fvxalksz5_0;
	wire w_dff_A_rC8rH8iX2_0;
	wire w_dff_A_srhtw1sZ8_0;
	wire w_dff_A_D8D7JTuH6_0;
	wire w_dff_A_BeNOCHJK7_0;
	wire w_dff_A_y8Nwq1Ec0_0;
	wire w_dff_A_vu1tZF2J9_0;
	wire w_dff_A_1hAiqw6U1_0;
	wire w_dff_A_wTmaZm8A1_0;
	wire w_dff_A_qoAP9IPY5_0;
	wire w_dff_A_Vn4DOyHy3_0;
	wire w_dff_A_BkJWTfI02_0;
	wire w_dff_A_JoP7uMAJ8_0;
	wire w_dff_A_Eo61JeLz8_0;
	wire w_dff_A_h2gs3CPy0_0;
	wire w_dff_A_3hektXhU1_0;
	wire w_dff_A_8z8TXkf17_0;
	wire w_dff_A_b83fJIyn8_0;
	wire w_dff_A_SeBPHW0r9_0;
	wire w_dff_A_ksVtyhS00_0;
	wire w_dff_A_4eq7X4Hm1_0;
	wire w_dff_A_BjAxq4mU0_2;
	wire w_dff_A_AlaYxrBK0_0;
	wire w_dff_A_8Np7gqqZ4_0;
	wire w_dff_A_FjVQ1N0P3_0;
	wire w_dff_A_YizKHwPR9_0;
	wire w_dff_A_wMP8YfKD9_0;
	wire w_dff_A_ktN8mmT99_0;
	wire w_dff_A_JtAFwv1D8_0;
	wire w_dff_A_GBlqMzBr5_0;
	wire w_dff_A_IV9sS5hg3_0;
	wire w_dff_A_tkCW5NPm9_0;
	wire w_dff_A_yYfyuP0p9_0;
	wire w_dff_A_JcOduGcL3_0;
	wire w_dff_A_GqbmMOa65_0;
	wire w_dff_A_UW2H3DRS7_0;
	wire w_dff_A_30Z7lW6x8_0;
	wire w_dff_A_e1uFaW1d9_0;
	wire w_dff_A_Yz3OiWn37_0;
	wire w_dff_A_AlUDMGWd7_0;
	wire w_dff_A_Ml85E7gs4_0;
	wire w_dff_A_rT4QnQEg1_0;
	wire w_dff_A_aUq1rw834_0;
	wire w_dff_A_08KUKXUt9_0;
	wire w_dff_A_7nAMY1rS0_0;
	wire w_dff_A_2m0EwwEg5_1;
	wire w_dff_A_I79e2AdF7_0;
	wire w_dff_A_6GkCo1DY6_0;
	wire w_dff_A_Lzey1E5Q1_0;
	wire w_dff_A_vCziq13r3_0;
	wire w_dff_A_GyxDS2LV9_0;
	wire w_dff_A_zjVysDTQ8_0;
	wire w_dff_A_kvqK0fIk0_0;
	wire w_dff_A_cugCo0mY1_0;
	wire w_dff_A_yswv97vH4_0;
	wire w_dff_A_OTfUuAtz5_0;
	wire w_dff_A_znDqZmWn2_0;
	wire w_dff_A_AnYQczUh4_0;
	wire w_dff_A_21UXCDvQ8_0;
	wire w_dff_A_2JPM1RxN1_0;
	wire w_dff_A_EPkzaIMr8_0;
	wire w_dff_A_3Zt31WK36_0;
	wire w_dff_A_PY7L3h4w1_0;
	wire w_dff_A_JT2Qq6Wb8_0;
	wire w_dff_A_UeYTx0wR9_0;
	wire w_dff_A_619BqzGV5_0;
	wire w_dff_A_jSmQNULw3_0;
	wire w_dff_A_B36V9xMd3_0;
	wire w_dff_A_hSejvORY1_0;
	wire w_dff_A_mRNqj3FC6_0;
	wire w_dff_A_WTjy3ssg7_0;
	wire w_dff_A_3zbxlb3T1_0;
	wire w_dff_A_ktr9uM4W4_0;
	wire w_dff_A_67FtK3pA2_1;
	wire w_dff_A_9dgE1jca0_0;
	wire w_dff_A_EP3B2JAi3_0;
	wire w_dff_A_73V960tj1_0;
	wire w_dff_A_9E9W0fdr0_0;
	wire w_dff_A_D1dyQpxn2_0;
	wire w_dff_A_GXm1967f7_0;
	wire w_dff_A_XfvMSRI60_0;
	wire w_dff_A_LEh3Tolj0_0;
	wire w_dff_A_8dce071Y0_0;
	wire w_dff_A_bh23YbnF9_0;
	wire w_dff_A_Sx3YBwK79_0;
	wire w_dff_A_TMjMIq1m6_0;
	wire w_dff_A_fDoeD3mO3_0;
	wire w_dff_A_BrM7y7Wq4_0;
	wire w_dff_A_MyPP7GLA4_0;
	wire w_dff_A_5QZCV04S1_0;
	wire w_dff_A_szl0iRQX2_0;
	wire w_dff_A_PpeJRPJC2_0;
	wire w_dff_A_alQXCNca7_0;
	wire w_dff_A_qpNJ4XxK8_0;
	wire w_dff_A_iltF4K2b2_0;
	wire w_dff_A_PGClOh0e2_0;
	wire w_dff_A_QXLh2RUm6_0;
	wire w_dff_A_Y1iaUumO9_0;
	wire w_dff_A_JNrj9jQy8_0;
	wire w_dff_A_tvKswgPv6_0;
	wire w_dff_A_wyNujQAN6_0;
	wire w_dff_A_gUc6hg5Q3_0;
	wire w_dff_A_Prsmcg8I7_0;
	wire w_dff_A_uaKJXgnV6_1;
	wire w_dff_A_h5JBuQF76_0;
	wire w_dff_A_2ZJ62Hke8_0;
	wire w_dff_A_ZNUX4UNg4_0;
	wire w_dff_A_WIkNu8zs2_0;
	wire w_dff_A_rS9ARH322_0;
	wire w_dff_A_i0Hh5bi44_0;
	wire w_dff_A_3I0MAEwU7_0;
	wire w_dff_A_LwMR0Vku3_0;
	wire w_dff_A_P2s9Y6sz8_0;
	wire w_dff_A_iWZ45yAQ5_0;
	wire w_dff_A_uTKPxXnP2_0;
	wire w_dff_A_EkrwcEyk3_0;
	wire w_dff_A_K5yjHLD10_0;
	wire w_dff_A_WJi3thGz1_0;
	wire w_dff_A_uxlGiOiS8_0;
	wire w_dff_A_hUpOauQa6_0;
	wire w_dff_A_PiMq0HRz4_0;
	wire w_dff_A_ignETw157_0;
	wire w_dff_A_sJCbjRRJ7_0;
	wire w_dff_A_hsKkG99B8_0;
	wire w_dff_A_iDVVtPbT9_0;
	wire w_dff_A_LHAjMOk64_0;
	wire w_dff_A_VIofv5Dt7_0;
	wire w_dff_A_ZaDQpY7l0_0;
	wire w_dff_A_6bOOtbGN8_0;
	wire w_dff_A_pMyue93u8_0;
	wire w_dff_A_AerFbYG80_0;
	wire w_dff_A_4Eh9CV0b4_0;
	wire w_dff_A_82ekGnhb0_2;
	wire w_dff_A_mKWthDho3_0;
	wire w_dff_A_FsWRfJGQ1_0;
	wire w_dff_A_GLDRUKkP5_0;
	wire w_dff_A_mMq5Lym85_0;
	wire w_dff_A_jigFhaxh6_0;
	wire w_dff_A_f8nkZmKJ0_0;
	wire w_dff_A_UsT9TBU19_0;
	wire w_dff_A_3HsUEeS55_0;
	wire w_dff_A_UMuR8MuL9_0;
	wire w_dff_A_pO8AZ6KA9_0;
	wire w_dff_A_ZJcOyy2e3_2;
	wire w_dff_A_COdxG20V3_0;
	wire w_dff_A_143LnfCB1_0;
	wire w_dff_A_GkHFLnsU3_0;
	wire w_dff_A_5KTqZrHY2_0;
	wire w_dff_A_jc0uY5c56_0;
	wire w_dff_A_dCB0pl8P9_0;
	wire w_dff_A_Xza456590_0;
	wire w_dff_A_QxziYi5t2_0;
	wire w_dff_A_yn8UVNzb7_0;
	wire w_dff_A_2F7OlOpe4_0;
	wire w_dff_A_fhIVqjCk4_2;
	wire w_dff_A_NchF0ExF4_0;
	wire w_dff_A_MF4fZL7G0_0;
	wire w_dff_A_WEzBVKBl6_0;
	wire w_dff_A_V1fSan9U2_1;
	wire w_dff_A_Ns3mTjbj3_0;
	wire w_dff_A_bvZgs5WK5_0;
	wire w_dff_A_wIVhEDTH4_0;
	wire w_dff_A_WyUpv4VO2_0;
	wire w_dff_A_8yYfWPyb3_0;
	wire w_dff_A_8LWQXudB1_0;
	wire w_dff_A_L4X1tgIA8_0;
	wire w_dff_A_1LZTMBJY8_0;
	wire w_dff_A_TxdXcCOk2_0;
	wire w_dff_A_on29UYq85_0;
	wire w_dff_A_2IKsu5tu1_0;
	wire w_dff_A_JCARljA63_0;
	wire w_dff_A_W2uEw8W79_0;
	wire w_dff_A_5ijsCaKo7_0;
	wire w_dff_A_yVOnFs1x9_0;
	wire w_dff_A_eoMt9YBF5_0;
	wire w_dff_A_62aXicn74_0;
	wire w_dff_A_3y16qGmv6_0;
	wire w_dff_A_lBVvOCYB5_0;
	wire w_dff_A_MXthOtod9_0;
	wire w_dff_A_GCOhVMYb7_2;
	wire w_dff_A_N3V3GSHY4_0;
	wire w_dff_A_WheD8US29_0;
	wire w_dff_A_mzqW7H6v3_0;
	wire w_dff_A_fn9tgkcG9_0;
	wire w_dff_A_OoLH6zQG7_0;
	wire w_dff_A_bWmbwUsV7_2;
	wire w_dff_A_fEr1VKOp6_0;
	wire w_dff_A_XgVXNhuH4_0;
	wire w_dff_A_QMRmzlLC3_0;
	wire w_dff_A_LTETGmhr2_0;
	wire w_dff_A_Zs4DPBih4_2;
	wire w_dff_A_7yna31FM6_0;
	wire w_dff_A_Epkq8GxI7_0;
	wire w_dff_A_j3fxXw7N2_0;
	wire w_dff_A_mNPRPVNR2_0;
	wire w_dff_A_d3U8Z1yA2_0;
	wire w_dff_A_8O4ZoJvT0_0;
	wire w_dff_A_b15N8rKA5_0;
	wire w_dff_A_uF1Aix0e0_0;
	wire w_dff_A_A2Ayl1W59_2;
	wire w_dff_A_6QfHv3ah8_0;
	wire w_dff_A_t4yerWQ56_0;
	wire w_dff_A_k8SIRAVT3_0;
	wire w_dff_A_mWHsMMDK2_0;
	wire w_dff_A_B914WQtK6_0;
	wire w_dff_A_Thea6Efg8_0;
	wire w_dff_A_9GdNTB9o9_0;
	wire w_dff_A_JEMRoawf2_0;
	wire w_dff_A_Di2h08h34_2;
	wire w_dff_A_cGtTuxfP2_0;
	wire w_dff_A_mrhQvpES1_2;
	wire w_dff_A_zDkIfLAq2_0;
	wire w_dff_A_iQ4quPVT4_2;
	wire w_dff_A_awmdFMC91_0;
	wire w_dff_A_bYZjOR4l8_2;
	wire w_dff_A_Sg8h2GHg4_0;
	wire w_dff_A_xodhc1gd3_0;
	wire w_dff_A_zhCzkvGB9_0;
	wire w_dff_A_4Rt6owKt7_0;
	wire w_dff_A_v9kVG2yQ4_0;
	wire w_dff_A_XgARWpSg8_0;
	wire w_dff_A_YMDJDxIo4_0;
	wire w_dff_A_0mQReEc72_0;
	wire w_dff_A_9SM2rFlR4_0;
	wire w_dff_A_QWXKn5Ug5_0;
	wire w_dff_A_s8pf0N6O3_0;
	wire w_dff_A_DRWXHmrG5_0;
	wire w_dff_A_2lVtROAw7_0;
	wire w_dff_A_ut142qF65_0;
	wire w_dff_A_Kf58cNfz8_0;
	wire w_dff_A_aPeUoKoA8_0;
	wire w_dff_A_SEuCHR110_0;
	wire w_dff_A_0APREGL63_0;
	wire w_dff_A_4unxHd6X7_0;
	wire w_dff_A_fpSu00BN5_0;
	wire w_dff_A_VsyDl8U20_0;
	wire w_dff_A_aMAuTsPq4_0;
	wire w_dff_A_pU2kcv4h2_0;
	wire w_dff_A_HbeBnZqG9_0;
	wire w_dff_A_xYcOwCKE4_2;
	wire w_dff_A_lp4BZ3Ra3_0;
	wire w_dff_A_MNWCFF3m6_0;
	wire w_dff_A_S8kL1AYv6_0;
	wire w_dff_A_9QEweryx9_0;
	wire w_dff_A_cWJs2vos8_0;
	wire w_dff_A_DKHFtTxw2_2;
	wire w_dff_A_GYaUbAuZ3_0;
	wire w_dff_A_5z2Rx1GY8_0;
	wire w_dff_A_v62LrHl38_0;
	wire w_dff_A_o6GMIi889_0;
	wire w_dff_A_FFhDPAqN4_0;
	wire w_dff_A_xHBLP3f76_2;
	wire w_dff_A_AcBhlfou6_0;
	wire w_dff_A_ftPGgdGO7_0;
	wire w_dff_A_Vd1u5Ds90_0;
	wire w_dff_A_WUj3Bhz24_0;
	wire w_dff_A_5FgrVi0f7_0;
	wire w_dff_A_kmbXyAx51_2;
	wire w_dff_A_6Xe8z1hJ0_0;
	wire w_dff_A_k7mUY3ae4_0;
	wire w_dff_A_gyjqWEac6_0;
	wire w_dff_A_n2xGXPLM7_0;
	wire w_dff_A_RAwpjRFA3_0;
	wire w_dff_A_KCAQtB6M2_0;
	wire w_dff_A_CNeCHZog3_0;
	wire w_dff_A_g9igXi8t2_2;
	wire w_dff_A_QWF5MNSI7_0;
	wire w_dff_A_JiJS0Jb39_0;
	wire w_dff_A_QvmVZT986_0;
	wire w_dff_A_YT14wwP74_0;
	wire w_dff_A_reEqvgj73_0;
	wire w_dff_A_4lwNbUNa5_0;
	wire w_dff_A_7YGOf3Tg3_0;
	wire w_dff_A_Q3YppFAk3_0;
	wire w_dff_A_guZB8wGF9_0;
	wire w_dff_A_22TNwHTZ8_0;
	wire w_dff_A_dz8hkwqB1_0;
	wire w_dff_A_mDA0UIXU1_0;
	wire w_dff_A_OrLuNpyR6_0;
	wire w_dff_A_7PDWFlxK6_0;
	wire w_dff_A_sizJU5Kv2_0;
	wire w_dff_A_w8OodaHw7_0;
	wire w_dff_A_bNDGyu6c7_0;
	wire w_dff_A_TGOisIUX3_0;
	wire w_dff_A_CsRxIJfP3_0;
	wire w_dff_A_DGJTufCb5_2;
	wire w_dff_A_4jJHDijp6_0;
	wire w_dff_A_RDG8Zhod6_2;
	wire w_dff_A_7lbDtceC0_0;
	wire w_dff_A_Snttc1Yu1_2;
	wire w_dff_A_j4qyzTbw6_0;
	wire w_dff_A_zInl2alh1_0;
	wire w_dff_A_t3ajAGXb6_0;
	wire w_dff_A_2MmhuD854_0;
	wire w_dff_A_WSPM8UuE1_0;
	wire w_dff_A_ffCIwah64_0;
	wire w_dff_A_M1ogNM1q4_0;
	wire w_dff_A_wvPK4jcW6_0;
	wire w_dff_A_Ay7YtLpr7_0;
	wire w_dff_A_n09qDzQp9_0;
	wire w_dff_A_cFBNnqgR7_0;
	wire w_dff_A_BqNKQ9v92_0;
	wire w_dff_A_NTodMKiG3_0;
	wire w_dff_A_PP7ucWkp5_0;
	wire w_dff_A_1ZcJDa6n1_0;
	wire w_dff_A_8bC3HfEN8_0;
	wire w_dff_A_iJoqc8sB5_0;
	wire w_dff_A_T4PMdRc97_2;
	wire w_dff_A_TKO326SN7_0;
	wire w_dff_A_PKXtIPsC3_0;
	wire w_dff_A_UMRMhsY89_0;
	wire w_dff_A_Yh1FBwUM8_0;
	wire w_dff_A_Z3HXBjD97_0;
	wire w_dff_A_vDcxGj9e0_0;
	wire w_dff_A_KTcEJu3D9_0;
	wire w_dff_A_iDMvqfhM1_0;
	wire w_dff_A_k7cGj2179_0;
	wire w_dff_A_dRvmNNQ72_0;
	wire w_dff_A_YJfnu9sG4_0;
	wire w_dff_A_R1B35dN19_0;
	wire w_dff_A_Abow7xoR7_0;
	wire w_dff_A_qP62sMNU0_0;
	wire w_dff_A_iy0AUKON6_0;
	wire w_dff_A_LXYKvGO26_0;
	wire w_dff_A_zt3cnxgn0_0;
	wire w_dff_A_B7P868BX1_2;
	wire w_dff_A_twqNrC4O3_0;
	wire w_dff_A_r2E4A33R4_0;
	wire w_dff_A_eimFmXYt7_0;
	wire w_dff_A_VKBRRyAn1_0;
	wire w_dff_A_puVLSrGL2_0;
	wire w_dff_A_z9J559Ir9_0;
	wire w_dff_A_2Rw37lrH3_0;
	wire w_dff_A_ATgClKxn7_0;
	wire w_dff_A_yzPcVvkx7_0;
	wire w_dff_A_RvmMBtZn8_0;
	wire w_dff_A_YXZXptmH8_0;
	wire w_dff_A_qXK4AFGg4_0;
	wire w_dff_A_UJlvFUtW7_0;
	wire w_dff_A_MSYfMvN65_0;
	wire w_dff_A_d14eUvhp3_0;
	wire w_dff_A_2PjQjbGr0_0;
	wire w_dff_A_JRksjT0Y4_0;
	wire w_dff_A_eHl8FGiB3_2;
	wire w_dff_A_ymbhNT8k6_0;
	wire w_dff_A_mGxwTEWz5_0;
	wire w_dff_A_9CU3jchR9_0;
	wire w_dff_A_pClrmOfj1_0;
	wire w_dff_A_KUfJE5t25_0;
	wire w_dff_A_sfMyqbEA3_0;
	wire w_dff_A_hr863h1V0_0;
	wire w_dff_A_6owKjLva0_0;
	wire w_dff_A_86LP1u9I2_0;
	wire w_dff_A_qmNOK5M19_0;
	wire w_dff_A_kYOh8TQN1_0;
	wire w_dff_A_3V49KIAp6_0;
	wire w_dff_A_OFiyNJQp4_0;
	wire w_dff_A_x1IFlwdf7_0;
	wire w_dff_A_9Qe4mkAm0_0;
	wire w_dff_A_SAGprpq54_0;
	wire w_dff_A_CTqnyzxH1_0;
	wire w_dff_A_5mhHFufl9_2;
	wire w_dff_A_19WJnn0R1_0;
	wire w_dff_A_duRybRl99_0;
	wire w_dff_A_SLFzaVaZ8_0;
	wire w_dff_A_aZmbzrCo5_0;
	wire w_dff_A_LJOtiIoB9_0;
	wire w_dff_A_GgEsdxbu5_0;
	wire w_dff_A_BiWMoxcW3_0;
	wire w_dff_A_l5BLak9X0_0;
	wire w_dff_A_XIjrMCKd7_0;
	wire w_dff_A_4OEcOAsP4_0;
	wire w_dff_A_tSCJWxxE3_0;
	wire w_dff_A_Yj5j4oGV8_0;
	wire w_dff_A_xY7oVWid9_2;
	wire w_dff_A_H7Bpe8DN4_0;
	wire w_dff_A_0aNFDEvN2_0;
	wire w_dff_A_KFanRTyL6_0;
	wire w_dff_A_yNWv5jkV2_0;
	wire w_dff_A_hieiPy7B8_0;
	wire w_dff_A_D2G9Ea7L4_0;
	wire w_dff_A_oykV85p26_0;
	wire w_dff_A_Lm3IZnW65_0;
	wire w_dff_A_g0i1D3m36_0;
	wire w_dff_A_eUYqKwrW7_0;
	wire w_dff_A_6YL5nnzd4_0;
	wire w_dff_A_pimnF4Yg8_0;
	wire w_dff_A_WzTSYKqK5_0;
	wire w_dff_A_fHXgdtt22_2;
	wire w_dff_A_gTNWBnM93_0;
	wire w_dff_A_TdsFmoIP6_0;
	wire w_dff_A_gAUiuOrl9_0;
	wire w_dff_A_Muibnq176_0;
	wire w_dff_A_oVp5WkuG8_0;
	wire w_dff_A_xtkFZcCD1_0;
	wire w_dff_A_qQDQ2b2E7_0;
	wire w_dff_A_qJXakTve7_0;
	wire w_dff_A_WlpHqxfu4_0;
	wire w_dff_A_ybmJz2dY0_0;
	wire w_dff_A_4uaK6ABo8_0;
	wire w_dff_A_Q2BsnpJv6_0;
	wire w_dff_A_YEAUu2gz1_0;
	wire w_dff_A_xXTSCJ4S6_0;
	wire w_dff_A_VECBTTSw6_0;
	wire w_dff_A_DuDkDjYi5_2;
	wire w_dff_A_dDB7qp5P3_0;
	wire w_dff_A_ujPwQOr92_0;
	wire w_dff_A_uv51KXtt9_0;
	wire w_dff_A_8SNbUtTT7_0;
	wire w_dff_A_VDkiLel90_0;
	wire w_dff_A_Xq16iuJx4_0;
	wire w_dff_A_EmpRYlBd5_0;
	wire w_dff_A_zQ4WrqJF6_0;
	wire w_dff_A_TaBkhPJf7_0;
	wire w_dff_A_Xnsx3GZd2_0;
	wire w_dff_A_qPoyoRLT4_0;
	wire w_dff_A_7PqEaO3n3_0;
	wire w_dff_A_WYwLRXyU9_0;
	wire w_dff_A_LxYwAEA64_0;
	wire w_dff_A_TAKFhnAa9_0;
	wire w_dff_A_NVjqnmDu3_0;
	wire w_dff_A_xgoaf3wx5_0;
	wire w_dff_A_jSAFT7W59_2;
	wire w_dff_A_ithHaM9Q9_0;
	wire w_dff_A_v6w6Ftd80_0;
	wire w_dff_A_Vl2GIAja8_0;
	wire w_dff_A_Cmblx7ZX3_0;
	wire w_dff_A_t9rU1ift3_0;
	wire w_dff_A_ViLkVnO16_2;
	wire w_dff_A_zgLAj29Z1_2;
	wire w_dff_A_8Py4PAuS1_0;
	wire w_dff_A_i0vAyBVg6_0;
	wire w_dff_A_LbjnRCS27_0;
	wire w_dff_A_n8oqx6re5_0;
	wire w_dff_A_00ppykpA8_0;
	wire w_dff_A_kaB0RiT85_0;
	wire w_dff_A_rcSvvZI04_0;
	wire w_dff_A_GfgDLexN6_0;
	wire w_dff_A_OWNeayUu7_0;
	wire w_dff_A_bquQDG432_0;
	wire w_dff_A_kOGCfB0W4_0;
	wire w_dff_A_xkYPtzHz6_0;
	wire w_dff_A_I849F7qj0_0;
	wire w_dff_A_jfGPZSUK9_0;
	wire w_dff_A_EJgYPLe23_0;
	wire w_dff_A_tx596gK83_0;
	wire w_dff_A_h2dOt8HR5_2;
	wire w_dff_A_hqGjitwK4_0;
	wire w_dff_A_jjcjwSm05_0;
	wire w_dff_A_F75Ogi0B6_0;
	wire w_dff_A_FU5Di0Jo4_0;
	wire w_dff_A_sOfyeLFc0_0;
	wire w_dff_A_4JhhMymf1_0;
	wire w_dff_A_Y3P78nY31_0;
	wire w_dff_A_aNI955nh5_0;
	wire w_dff_A_aU3f0mlL2_0;
	wire w_dff_A_n6MTmMDB2_0;
	wire w_dff_A_YGVnJeVP7_0;
	wire w_dff_A_MYi7ROnW9_0;
	wire w_dff_A_EIJTCDdr0_0;
	wire w_dff_A_n1wO9CLk5_0;
	wire w_dff_A_hRfp8CU42_0;
	wire w_dff_A_YlkdBaCC6_0;
	wire w_dff_A_uxLl9poC2_0;
	wire w_dff_A_MmJRikpF7_0;
	wire w_dff_A_X5aQ5GJ57_0;
	wire w_dff_A_vRhT0YsU5_0;
	jnot g0000(.din(w_G15_0[2]),.dout(w_dff_A_Ecw3XE0C8_1),.clk(gclk));
	jor g0001(.dina(G57),.dinb(w_G5_1[1]),.dout(w_dff_A_l29pao1a2_2),.clk(gclk));
	jnot g0002(.din(G184),.dout(n317),.clk(gclk));
	jnot g0003(.din(G228),.dout(n318),.clk(gclk));
	jor g0004(.dina(n318),.dinb(n317),.dout(n319),.clk(gclk));
	jnot g0005(.din(G150),.dout(n320),.clk(gclk));
	jnot g0006(.din(G240),.dout(n321),.clk(gclk));
	jor g0007(.dina(n321),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0008(.dina(n322),.dinb(n319),.dout(G404_fa_),.clk(gclk));
	jnot g0009(.din(G210),.dout(n324),.clk(gclk));
	jnot g0010(.din(G218),.dout(n325),.clk(gclk));
	jor g0011(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jnot g0012(.din(G152),.dout(n327),.clk(gclk));
	jnot g0013(.din(G230),.dout(n328),.clk(gclk));
	jor g0014(.dina(n328),.dinb(n327),.dout(n329),.clk(gclk));
	jor g0015(.dina(n329),.dinb(n326),.dout(G406_fa_),.clk(gclk));
	jnot g0016(.din(G183),.dout(n331),.clk(gclk));
	jnot g0017(.din(G185),.dout(n332),.clk(gclk));
	jor g0018(.dina(n332),.dinb(n331),.dout(n333),.clk(gclk));
	jnot g0019(.din(G182),.dout(n334),.clk(gclk));
	jnot g0020(.din(G186),.dout(n335),.clk(gclk));
	jor g0021(.dina(n335),.dinb(n334),.dout(n336),.clk(gclk));
	jor g0022(.dina(n336),.dinb(n333),.dout(G408_fa_),.clk(gclk));
	jnot g0023(.din(G172),.dout(n338),.clk(gclk));
	jnot g0024(.din(G188),.dout(n339),.clk(gclk));
	jor g0025(.dina(n339),.dinb(n338),.dout(n340),.clk(gclk));
	jnot g0026(.din(G162),.dout(n341),.clk(gclk));
	jnot g0027(.din(G199),.dout(n342),.clk(gclk));
	jor g0028(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jor g0029(.dina(n343),.dinb(n340),.dout(G410_fa_),.clk(gclk));
	jnot g0030(.din(G1197),.dout(n345),.clk(gclk));
	jor g0031(.dina(w_n345_0[1]),.dinb(w_G5_1[0]),.dout(w_dff_A_shAXd2VJ7_2),.clk(gclk));
	jnot g0032(.din(G134),.dout(n347),.clk(gclk));
	jnot g0033(.din(G133),.dout(n348),.clk(gclk));
	jor g0034(.dina(n348),.dinb(w_G5_0[2]),.dout(n349),.clk(gclk));
	jor g0035(.dina(w_n349_0[1]),.dinb(w_n347_0[1]),.dout(w_dff_A_5CWJDb799_2),.clk(gclk));
	jand g0036(.dina(G163),.dinb(w_G1_1[2]),.dout(w_dff_A_6JNnbqa23_2),.clk(gclk));
	jnot g0037(.din(w_G41_0[1]),.dout(n352),.clk(gclk));
	jor g0038(.dina(n352),.dinb(w_G18_49[2]),.dout(n353),.clk(gclk));
	jor g0039(.dina(w_n353_0[1]),.dinb(w_G3701_1[1]),.dout(n354),.clk(gclk));
	jnot g0040(.din(w_G18_49[1]),.dout(n355),.clk(gclk));
	jand g0041(.dina(w_G3701_1[0]),.dinb(w_n355_35[2]),.dout(n356),.clk(gclk));
	jand g0042(.dina(n356),.dinb(w_n353_0[0]),.dout(n357),.clk(gclk));
	jnot g0043(.din(w_n357_0[1]),.dout(n358),.clk(gclk));
	jand g0044(.dina(w_n358_0[1]),.dinb(w_n354_0[2]),.dout(n359),.clk(gclk));
	jxor g0045(.dina(w_n359_1[1]),.dinb(w_G4526_2[2]),.dout(w_dff_A_JUhLnoel6_2),.clk(gclk));
	jnot g0046(.din(w_G38_2[2]),.dout(n361),.clk(gclk));
	jand g0047(.dina(w_G4528_0[2]),.dinb(w_G1492_1[1]),.dout(n362),.clk(gclk));
	jxor g0048(.dina(w_n362_0[2]),.dinb(w_n361_0[2]),.dout(n363),.clk(gclk));
	jand g0049(.dina(w_G4528_0[1]),.dinb(w_G1496_1[1]),.dout(n364),.clk(gclk));
	jor g0050(.dina(w_n364_0[2]),.dinb(w_n361_0[1]),.dout(n365),.clk(gclk));
	jnot g0051(.din(w_G1496_1[0]),.dout(n366),.clk(gclk));
	jnot g0052(.din(w_G4528_0[0]),.dout(n367),.clk(gclk));
	jor g0053(.dina(w_n367_0[1]),.dinb(w_G38_2[1]),.dout(n368),.clk(gclk));
	jor g0054(.dina(w_n368_0[1]),.dinb(w_n366_0[2]),.dout(n369),.clk(gclk));
	jand g0055(.dina(w_n369_0[1]),.dinb(n365),.dout(n370),.clk(gclk));
	jnot g0056(.din(w_G1486_0[1]),.dout(n371),.clk(gclk));
	jand g0057(.dina(G12),.dinb(G9),.dout(n372),.clk(gclk));
	jnot g0058(.din(w_n372_0[1]),.dout(n373),.clk(gclk));
	jor g0059(.dina(G213),.dinb(w_n355_35[1]),.dout(n374),.clk(gclk));
	jand g0060(.dina(w_n374_0[1]),.dinb(w_n373_9[2]),.dout(n375),.clk(gclk));
	jand g0061(.dina(w_n375_0[2]),.dinb(w_n371_0[2]),.dout(n376),.clk(gclk));
	jxor g0062(.dina(w_n375_0[1]),.dinb(w_n371_0[1]),.dout(n377),.clk(gclk));
	jor g0063(.dina(G214),.dinb(w_n355_35[0]),.dout(n378),.clk(gclk));
	jand g0064(.dina(w_n378_0[1]),.dinb(w_n373_9[1]),.dout(n379),.clk(gclk));
	jnot g0065(.din(w_n379_0[2]),.dout(n380),.clk(gclk));
	jand g0066(.dina(w_n380_0[1]),.dinb(w_G1480_0[2]),.dout(n381),.clk(gclk));
	jnot g0067(.din(n381),.dout(n382),.clk(gclk));
	jnot g0068(.din(w_G1480_0[1]),.dout(n383),.clk(gclk));
	jand g0069(.dina(w_n379_0[1]),.dinb(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g0070(.din(w_G106_1[1]),.dout(n385),.clk(gclk));
	jor g0071(.dina(G215),.dinb(w_n355_34[2]),.dout(n386),.clk(gclk));
	jand g0072(.dina(w_n386_0[1]),.dinb(w_n373_9[0]),.dout(n387),.clk(gclk));
	jxor g0073(.dina(w_n387_1[1]),.dinb(w_n385_0[1]),.dout(n388),.clk(gclk));
	jnot g0074(.din(w_G1462_0[1]),.dout(n389),.clk(gclk));
	jor g0075(.dina(w_G209_0[1]),.dinb(w_n355_34[1]),.dout(n390),.clk(gclk));
	jand g0076(.dina(n390),.dinb(w_n373_8[2]),.dout(n391),.clk(gclk));
	jand g0077(.dina(w_n391_0[2]),.dinb(w_n389_1[1]),.dout(n392),.clk(gclk));
	jnot g0078(.din(w_G1469_0[1]),.dout(n393),.clk(gclk));
	jor g0079(.dina(G216),.dinb(w_n355_34[0]),.dout(n394),.clk(gclk));
	jand g0080(.dina(w_n394_0[1]),.dinb(w_n373_8[1]),.dout(n395),.clk(gclk));
	jxor g0081(.dina(w_n395_1[1]),.dinb(w_n393_1[1]),.dout(n396),.clk(gclk));
	jand g0082(.dina(w_n396_1[2]),.dinb(w_n392_0[2]),.dout(n397),.clk(gclk));
	jand g0083(.dina(w_n397_0[1]),.dinb(w_n388_1[2]),.dout(n398),.clk(gclk));
	jnot g0084(.din(n398),.dout(n399),.clk(gclk));
	jand g0085(.dina(w_n387_1[0]),.dinb(w_n385_0[0]),.dout(n400),.clk(gclk));
	jnot g0086(.din(n400),.dout(n401),.clk(gclk));
	jnot g0087(.din(w_n387_0[2]),.dout(n402),.clk(gclk));
	jand g0088(.dina(n402),.dinb(w_G106_1[0]),.dout(n403),.clk(gclk));
	jand g0089(.dina(w_n395_1[0]),.dinb(w_n393_1[0]),.dout(n404),.clk(gclk));
	jnot g0090(.din(n404),.dout(n405),.clk(gclk));
	jor g0091(.dina(w_n405_0[2]),.dinb(n403),.dout(n406),.clk(gclk));
	jand g0092(.dina(n406),.dinb(n401),.dout(n407),.clk(gclk));
	jand g0093(.dina(w_n407_0[1]),.dinb(n399),.dout(n408),.clk(gclk));
	jnot g0094(.din(n408),.dout(n409),.clk(gclk));
	jor g0095(.dina(w_n409_1[1]),.dinb(n384),.dout(n410),.clk(gclk));
	jand g0096(.dina(n410),.dinb(n382),.dout(n411),.clk(gclk));
	jand g0097(.dina(w_n411_1[1]),.dinb(w_n377_1[2]),.dout(n412),.clk(gclk));
	jor g0098(.dina(n412),.dinb(n376),.dout(n413),.clk(gclk));
	jxor g0099(.dina(w_n391_0[1]),.dinb(w_n389_1[0]),.dout(n414),.clk(gclk));
	jand g0100(.dina(w_n414_1[1]),.dinb(w_n396_1[1]),.dout(n415),.clk(gclk));
	jxor g0101(.dina(w_n379_0[0]),.dinb(w_n383_0[1]),.dout(n416),.clk(gclk));
	jand g0102(.dina(w_n416_0[2]),.dinb(w_n388_1[1]),.dout(n417),.clk(gclk));
	jand g0103(.dina(n417),.dinb(w_n415_0[1]),.dout(n418),.clk(gclk));
	jand g0104(.dina(w_n418_0[1]),.dinb(w_n377_1[1]),.dout(n419),.clk(gclk));
	jor g0105(.dina(w_n419_0[1]),.dinb(w_n413_1[1]),.dout(n420),.clk(gclk));
	jnot g0106(.din(w_G2256_0[1]),.dout(n421),.clk(gclk));
	jor g0107(.dina(G153),.dinb(w_n355_33[2]),.dout(n422),.clk(gclk));
	jand g0108(.dina(w_n422_0[1]),.dinb(w_n373_8[0]),.dout(n423),.clk(gclk));
	jand g0109(.dina(w_n423_0[2]),.dinb(w_n421_0[2]),.dout(n424),.clk(gclk));
	jxor g0110(.dina(w_n423_0[1]),.dinb(w_n421_0[1]),.dout(n425),.clk(gclk));
	jnot g0111(.din(w_G2253_0[2]),.dout(n426),.clk(gclk));
	jor g0112(.dina(G154),.dinb(w_n355_33[1]),.dout(n427),.clk(gclk));
	jand g0113(.dina(w_n427_0[1]),.dinb(w_n373_7[2]),.dout(n428),.clk(gclk));
	jxor g0114(.dina(w_n428_0[2]),.dinb(w_n426_0[2]),.dout(n429),.clk(gclk));
	jnot g0115(.din(w_G2247_0[2]),.dout(n430),.clk(gclk));
	jor g0116(.dina(G155),.dinb(w_n355_33[0]),.dout(n431),.clk(gclk));
	jand g0117(.dina(w_n431_0[1]),.dinb(w_n373_7[1]),.dout(n432),.clk(gclk));
	jxor g0118(.dina(w_n432_0[2]),.dinb(w_n430_0[1]),.dout(n433),.clk(gclk));
	jnot g0119(.din(w_G2239_1[1]),.dout(n434),.clk(gclk));
	jor g0120(.dina(G156),.dinb(w_n355_32[2]),.dout(n435),.clk(gclk));
	jand g0121(.dina(w_n435_0[1]),.dinb(w_n373_7[0]),.dout(n436),.clk(gclk));
	jxor g0122(.dina(w_n436_0[2]),.dinb(w_n434_0[1]),.dout(n437),.clk(gclk));
	jand g0123(.dina(w_n437_0[2]),.dinb(w_n433_1[2]),.dout(n438),.clk(gclk));
	jand g0124(.dina(w_n438_0[1]),.dinb(w_n429_0[2]),.dout(n439),.clk(gclk));
	jnot g0125(.din(w_n428_0[1]),.dout(n440),.clk(gclk));
	jand g0126(.dina(w_n440_0[1]),.dinb(w_G2253_0[1]),.dout(n441),.clk(gclk));
	jnot g0127(.din(n441),.dout(n442),.clk(gclk));
	jand g0128(.dina(w_n428_0[0]),.dinb(w_n426_0[1]),.dout(n443),.clk(gclk));
	jand g0129(.dina(w_n432_0[1]),.dinb(w_n430_0[0]),.dout(n444),.clk(gclk));
	jand g0130(.dina(w_n436_0[1]),.dinb(w_n434_0[0]),.dout(n445),.clk(gclk));
	jand g0131(.dina(w_n445_0[2]),.dinb(w_n433_1[1]),.dout(n446),.clk(gclk));
	jor g0132(.dina(n446),.dinb(w_n444_0[2]),.dout(n447),.clk(gclk));
	jor g0133(.dina(w_n447_0[2]),.dinb(n443),.dout(n448),.clk(gclk));
	jand g0134(.dina(n448),.dinb(n442),.dout(n449),.clk(gclk));
	jor g0135(.dina(w_n449_1[1]),.dinb(n439),.dout(n450),.clk(gclk));
	jnot g0136(.din(w_G2236_0[2]),.dout(n451),.clk(gclk));
	jor g0137(.dina(G157),.dinb(w_n355_32[1]),.dout(n452),.clk(gclk));
	jand g0138(.dina(n452),.dinb(w_n373_6[2]),.dout(n453),.clk(gclk));
	jand g0139(.dina(w_n453_1[1]),.dinb(w_n451_0[2]),.dout(n454),.clk(gclk));
	jor g0140(.dina(w_n453_1[0]),.dinb(w_n451_0[1]),.dout(n455),.clk(gclk));
	jnot g0141(.din(w_G2230_0[2]),.dout(n456),.clk(gclk));
	jand g0142(.dina(G135),.dinb(w_n355_32[0]),.dout(n457),.clk(gclk));
	jand g0143(.dina(G158),.dinb(w_G18_49[0]),.dout(n458),.clk(gclk));
	jor g0144(.dina(n458),.dinb(w_n457_0[1]),.dout(n459),.clk(gclk));
	jand g0145(.dina(w_n459_0[2]),.dinb(w_n456_0[2]),.dout(n460),.clk(gclk));
	jand g0146(.dina(w_n460_1[2]),.dinb(n455),.dout(n461),.clk(gclk));
	jor g0147(.dina(n461),.dinb(n454),.dout(n462),.clk(gclk));
	jxor g0148(.dina(w_n453_0[2]),.dinb(w_n451_0[0]),.dout(n463),.clk(gclk));
	jxor g0149(.dina(w_n459_0[1]),.dinb(w_n456_0[1]),.dout(n464),.clk(gclk));
	jand g0150(.dina(w_n464_0[2]),.dinb(w_n463_1[1]),.dout(n465),.clk(gclk));
	jnot g0151(.din(w_G2224_1[1]),.dout(n466),.clk(gclk));
	jand g0152(.dina(G144),.dinb(w_n355_31[2]),.dout(n467),.clk(gclk));
	jand g0153(.dina(G159),.dinb(w_G18_48[2]),.dout(n468),.clk(gclk));
	jor g0154(.dina(n468),.dinb(w_n467_0[1]),.dout(n469),.clk(gclk));
	jxor g0155(.dina(w_n469_1[1]),.dinb(w_n466_0[1]),.dout(n470),.clk(gclk));
	jnot g0156(.din(w_G2218_0[2]),.dout(n471),.clk(gclk));
	jand g0157(.dina(G138),.dinb(w_n355_31[1]),.dout(n472),.clk(gclk));
	jand g0158(.dina(G160),.dinb(w_G18_48[1]),.dout(n473),.clk(gclk));
	jor g0159(.dina(n473),.dinb(w_n472_0[1]),.dout(n474),.clk(gclk));
	jxor g0160(.dina(w_n474_0[2]),.dinb(w_n471_0[2]),.dout(n475),.clk(gclk));
	jnot g0161(.din(w_G2211_0[2]),.dout(n476),.clk(gclk));
	jand g0162(.dina(G147),.dinb(w_n355_31[0]),.dout(n477),.clk(gclk));
	jand g0163(.dina(G151),.dinb(w_G18_48[0]),.dout(n478),.clk(gclk));
	jor g0164(.dina(n478),.dinb(w_n477_0[1]),.dout(n479),.clk(gclk));
	jxor g0165(.dina(w_n479_1[1]),.dinb(w_n476_0[2]),.dout(n480),.clk(gclk));
	jand g0166(.dina(w_n480_1[1]),.dinb(w_n475_0[2]),.dout(n481),.clk(gclk));
	jand g0167(.dina(w_n481_0[1]),.dinb(w_n470_0[2]),.dout(n482),.clk(gclk));
	jnot g0168(.din(w_n469_1[0]),.dout(n483),.clk(gclk));
	jand g0169(.dina(n483),.dinb(w_G2224_1[0]),.dout(n484),.clk(gclk));
	jnot g0170(.din(w_n474_0[1]),.dout(n485),.clk(gclk));
	jand g0171(.dina(w_n485_0[1]),.dinb(w_G2218_0[1]),.dout(n486),.clk(gclk));
	jand g0172(.dina(w_n479_1[0]),.dinb(w_n476_0[1]),.dout(n487),.clk(gclk));
	jnot g0173(.din(w_n487_0[2]),.dout(n488),.clk(gclk));
	jor g0174(.dina(n488),.dinb(w_n486_0[1]),.dout(n489),.clk(gclk));
	jand g0175(.dina(w_n469_0[2]),.dinb(w_n466_0[0]),.dout(n490),.clk(gclk));
	jand g0176(.dina(w_n474_0[0]),.dinb(w_n471_0[1]),.dout(n491),.clk(gclk));
	jor g0177(.dina(w_n491_1[1]),.dinb(n490),.dout(n492),.clk(gclk));
	jnot g0178(.din(n492),.dout(n493),.clk(gclk));
	jand g0179(.dina(n493),.dinb(w_n489_0[2]),.dout(n494),.clk(gclk));
	jor g0180(.dina(n494),.dinb(n484),.dout(n495),.clk(gclk));
	jnot g0181(.din(w_n495_1[1]),.dout(n496),.clk(gclk));
	jor g0182(.dina(w_n496_0[2]),.dinb(n482),.dout(n497),.clk(gclk));
	jand g0183(.dina(w_n497_1[1]),.dinb(w_n465_0[1]),.dout(n498),.clk(gclk));
	jor g0184(.dina(n498),.dinb(w_n462_0[2]),.dout(n499),.clk(gclk));
	jand g0185(.dina(w_n496_0[1]),.dinb(w_n465_0[0]),.dout(n500),.clk(gclk));
	jnot g0186(.din(w_G4437_0[2]),.dout(n501),.clk(gclk));
	jand g0187(.dina(G219),.dinb(w_G18_47[2]),.dout(n502),.clk(gclk));
	jand g0188(.dina(G66),.dinb(w_n355_30[2]),.dout(n503),.clk(gclk));
	jor g0189(.dina(w_n503_0[1]),.dinb(n502),.dout(n504),.clk(gclk));
	jand g0190(.dina(w_n504_1[1]),.dinb(w_n501_0[2]),.dout(n505),.clk(gclk));
	jnot g0191(.din(w_n504_1[0]),.dout(n506),.clk(gclk));
	jand g0192(.dina(n506),.dinb(w_G4437_0[1]),.dout(n507),.clk(gclk));
	jnot g0193(.din(w_n507_0[1]),.dout(n508),.clk(gclk));
	jnot g0194(.din(w_G4432_0[2]),.dout(n509),.clk(gclk));
	jand g0195(.dina(G220),.dinb(w_G18_47[1]),.dout(n510),.clk(gclk));
	jand g0196(.dina(G50),.dinb(w_n355_30[1]),.dout(n511),.clk(gclk));
	jor g0197(.dina(w_n511_0[1]),.dinb(n510),.dout(n512),.clk(gclk));
	jxor g0198(.dina(w_n512_0[2]),.dinb(w_n509_0[2]),.dout(n513),.clk(gclk));
	jnot g0199(.din(w_G4420_1[1]),.dout(n514),.clk(gclk));
	jand g0200(.dina(G222),.dinb(w_G18_47[0]),.dout(n515),.clk(gclk));
	jand g0201(.dina(G35),.dinb(w_n355_30[0]),.dout(n516),.clk(gclk));
	jor g0202(.dina(w_n516_0[1]),.dinb(n515),.dout(n517),.clk(gclk));
	jand g0203(.dina(w_n517_1[1]),.dinb(w_n514_0[1]),.dout(n518),.clk(gclk));
	jnot g0204(.din(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0205(.din(w_G4427_0[2]),.dout(n520),.clk(gclk));
	jand g0206(.dina(G221),.dinb(w_G18_46[2]),.dout(n521),.clk(gclk));
	jand g0207(.dina(G32),.dinb(w_n355_29[2]),.dout(n522),.clk(gclk));
	jor g0208(.dina(w_n522_0[1]),.dinb(n521),.dout(n523),.clk(gclk));
	jxor g0209(.dina(w_n523_0[2]),.dinb(w_n520_0[1]),.dout(n524),.clk(gclk));
	jnot g0210(.din(w_n517_1[0]),.dout(n525),.clk(gclk));
	jand g0211(.dina(n525),.dinb(w_G4420_1[0]),.dout(n526),.clk(gclk));
	jnot g0212(.din(w_n526_0[2]),.dout(n527),.clk(gclk));
	jnot g0213(.din(w_G4415_1[1]),.dout(n528),.clk(gclk));
	jand g0214(.dina(G223),.dinb(w_G18_46[1]),.dout(n529),.clk(gclk));
	jand g0215(.dina(G47),.dinb(w_n355_29[1]),.dout(n530),.clk(gclk));
	jor g0216(.dina(w_n530_0[1]),.dinb(n529),.dout(n531),.clk(gclk));
	jand g0217(.dina(w_n531_1[1]),.dinb(w_n528_0[1]),.dout(n532),.clk(gclk));
	jnot g0218(.din(w_n531_1[0]),.dout(n533),.clk(gclk));
	jand g0219(.dina(n533),.dinb(w_G4415_1[0]),.dout(n534),.clk(gclk));
	jnot g0220(.din(n534),.dout(n535),.clk(gclk));
	jnot g0221(.din(w_G4410_0[2]),.dout(n536),.clk(gclk));
	jand g0222(.dina(G224),.dinb(w_G18_46[0]),.dout(n537),.clk(gclk));
	jand g0223(.dina(G121),.dinb(w_n355_29[0]),.dout(n538),.clk(gclk));
	jor g0224(.dina(w_n538_0[1]),.dinb(n537),.dout(n539),.clk(gclk));
	jand g0225(.dina(w_n539_1[1]),.dinb(w_n536_0[2]),.dout(n540),.clk(gclk));
	jnot g0226(.din(w_n539_1[0]),.dout(n541),.clk(gclk));
	jand g0227(.dina(n541),.dinb(w_G4410_0[1]),.dout(n542),.clk(gclk));
	jnot g0228(.din(n542),.dout(n543),.clk(gclk));
	jnot g0229(.din(w_G4405_1[1]),.dout(n544),.clk(gclk));
	jand g0230(.dina(G225),.dinb(w_G18_45[2]),.dout(n545),.clk(gclk));
	jand g0231(.dina(G94),.dinb(w_n355_28[2]),.dout(n546),.clk(gclk));
	jor g0232(.dina(w_n546_0[1]),.dinb(n545),.dout(n547),.clk(gclk));
	jand g0233(.dina(w_n547_1[1]),.dinb(w_n544_0[1]),.dout(n548),.clk(gclk));
	jnot g0234(.din(w_n547_1[0]),.dout(n549),.clk(gclk));
	jand g0235(.dina(n549),.dinb(w_G4405_1[0]),.dout(n550),.clk(gclk));
	jnot g0236(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0237(.din(w_G4400_1[1]),.dout(n552),.clk(gclk));
	jand g0238(.dina(G226),.dinb(w_G18_45[1]),.dout(n553),.clk(gclk));
	jand g0239(.dina(G97),.dinb(w_n355_28[1]),.dout(n554),.clk(gclk));
	jor g0240(.dina(w_n554_0[1]),.dinb(n553),.dout(n555),.clk(gclk));
	jand g0241(.dina(w_n555_1[1]),.dinb(w_n552_0[1]),.dout(n556),.clk(gclk));
	jnot g0242(.din(w_n555_1[0]),.dout(n557),.clk(gclk));
	jand g0243(.dina(n557),.dinb(w_G4400_1[0]),.dout(n558),.clk(gclk));
	jnot g0244(.din(w_n558_0[1]),.dout(n559),.clk(gclk));
	jnot g0245(.din(w_G4394_1[1]),.dout(n560),.clk(gclk));
	jand g0246(.dina(G217),.dinb(w_G18_45[0]),.dout(n561),.clk(gclk));
	jand g0247(.dina(G118),.dinb(w_n355_28[0]),.dout(n562),.clk(gclk));
	jor g0248(.dina(w_n562_0[1]),.dinb(n561),.dout(n563),.clk(gclk));
	jand g0249(.dina(w_n563_1[1]),.dinb(w_n560_0[1]),.dout(n564),.clk(gclk));
	jand g0250(.dina(w_n564_0[2]),.dinb(n559),.dout(n565),.clk(gclk));
	jor g0251(.dina(w_n565_0[1]),.dinb(w_n556_0[2]),.dout(n566),.clk(gclk));
	jand g0252(.dina(w_n566_0[2]),.dinb(n551),.dout(n567),.clk(gclk));
	jor g0253(.dina(n567),.dinb(w_n548_0[1]),.dout(n568),.clk(gclk));
	jand g0254(.dina(w_n568_0[2]),.dinb(n543),.dout(n569),.clk(gclk));
	jor g0255(.dina(n569),.dinb(n540),.dout(n570),.clk(gclk));
	jand g0256(.dina(w_n570_1[2]),.dinb(n535),.dout(n571),.clk(gclk));
	jor g0257(.dina(n571),.dinb(n532),.dout(n572),.clk(gclk));
	jxor g0258(.dina(w_n531_0[2]),.dinb(w_n528_0[0]),.dout(n573),.clk(gclk));
	jxor g0259(.dina(w_n555_0[2]),.dinb(w_n552_0[0]),.dout(n574),.clk(gclk));
	jxor g0260(.dina(w_n563_1[0]),.dinb(w_n560_0[0]),.dout(n575),.clk(gclk));
	jand g0261(.dina(w_n575_1[1]),.dinb(w_n574_0[2]),.dout(n576),.clk(gclk));
	jxor g0262(.dina(w_n539_0[2]),.dinb(w_n536_0[1]),.dout(n577),.clk(gclk));
	jxor g0263(.dina(w_n547_0[2]),.dinb(w_n544_0[0]),.dout(n578),.clk(gclk));
	jand g0264(.dina(w_n578_0[2]),.dinb(w_n577_0[1]),.dout(n579),.clk(gclk));
	jand g0265(.dina(n579),.dinb(w_n576_0[2]),.dout(n580),.clk(gclk));
	jand g0266(.dina(w_n580_0[2]),.dinb(w_n573_1[1]),.dout(n581),.clk(gclk));
	jnot g0267(.din(w_G3749_0[2]),.dout(n582),.clk(gclk));
	jand g0268(.dina(G231),.dinb(w_G18_44[2]),.dout(n583),.clk(gclk));
	jand g0269(.dina(G100),.dinb(w_n355_27[2]),.dout(n584),.clk(gclk));
	jor g0270(.dina(w_n584_0[1]),.dinb(n583),.dout(n585),.clk(gclk));
	jand g0271(.dina(w_n585_1[1]),.dinb(w_n582_0[2]),.dout(n586),.clk(gclk));
	jnot g0272(.din(w_n585_1[0]),.dout(n587),.clk(gclk));
	jand g0273(.dina(n587),.dinb(w_G3749_0[1]),.dout(n588),.clk(gclk));
	jnot g0274(.din(w_n588_0[1]),.dout(n589),.clk(gclk));
	jnot g0275(.din(w_G3743_0[2]),.dout(n590),.clk(gclk));
	jand g0276(.dina(G232),.dinb(w_G18_44[1]),.dout(n591),.clk(gclk));
	jand g0277(.dina(G124),.dinb(w_n355_27[1]),.dout(n592),.clk(gclk));
	jor g0278(.dina(w_n592_0[1]),.dinb(n591),.dout(n593),.clk(gclk));
	jxor g0279(.dina(w_n593_1[1]),.dinb(w_n590_0[2]),.dout(n594),.clk(gclk));
	jnot g0280(.din(w_G3737_0[2]),.dout(n595),.clk(gclk));
	jand g0281(.dina(G233),.dinb(w_G18_44[0]),.dout(n596),.clk(gclk));
	jand g0282(.dina(G127),.dinb(w_n355_27[0]),.dout(n597),.clk(gclk));
	jor g0283(.dina(w_n597_0[1]),.dinb(n596),.dout(n598),.clk(gclk));
	jxor g0284(.dina(w_n598_1[1]),.dinb(w_n595_0[2]),.dout(n599),.clk(gclk));
	jnot g0285(.din(w_G3729_1[1]),.dout(n600),.clk(gclk));
	jand g0286(.dina(G234),.dinb(w_G18_43[2]),.dout(n601),.clk(gclk));
	jand g0287(.dina(G130),.dinb(w_n355_26[2]),.dout(n602),.clk(gclk));
	jor g0288(.dina(w_n602_0[1]),.dinb(n601),.dout(n603),.clk(gclk));
	jxor g0289(.dina(w_n603_1[1]),.dinb(w_n600_0[1]),.dout(n604),.clk(gclk));
	jand g0290(.dina(w_n604_0[1]),.dinb(w_n599_0[2]),.dout(n605),.clk(gclk));
	jand g0291(.dina(w_n605_0[2]),.dinb(w_n594_0[2]),.dout(n606),.clk(gclk));
	jnot g0292(.din(n606),.dout(n607),.clk(gclk));
	jnot g0293(.din(w_n593_1[0]),.dout(n608),.clk(gclk));
	jand g0294(.dina(n608),.dinb(w_G3743_0[1]),.dout(n609),.clk(gclk));
	jand g0295(.dina(w_n593_0[2]),.dinb(w_n590_0[1]),.dout(n610),.clk(gclk));
	jnot g0296(.din(w_n610_0[1]),.dout(n611),.clk(gclk));
	jand g0297(.dina(w_n598_1[0]),.dinb(w_n595_0[1]),.dout(n612),.clk(gclk));
	jand g0298(.dina(w_n603_1[0]),.dinb(w_n600_0[0]),.dout(n613),.clk(gclk));
	jand g0299(.dina(w_n613_0[2]),.dinb(w_n599_0[1]),.dout(n614),.clk(gclk));
	jor g0300(.dina(n614),.dinb(w_n612_0[1]),.dout(n615),.clk(gclk));
	jnot g0301(.din(w_n615_0[2]),.dout(n616),.clk(gclk));
	jand g0302(.dina(w_n616_0[1]),.dinb(n611),.dout(n617),.clk(gclk));
	jor g0303(.dina(n617),.dinb(w_n609_0[1]),.dout(n618),.clk(gclk));
	jand g0304(.dina(w_n618_0[2]),.dinb(n607),.dout(n619),.clk(gclk));
	jnot g0305(.din(w_n619_0[2]),.dout(n620),.clk(gclk));
	jnot g0306(.din(w_n618_0[1]),.dout(n621),.clk(gclk));
	jnot g0307(.din(w_G3723_0[2]),.dout(n622),.clk(gclk));
	jand g0308(.dina(G235),.dinb(w_G18_43[1]),.dout(n623),.clk(gclk));
	jand g0309(.dina(G103),.dinb(w_n355_26[1]),.dout(n624),.clk(gclk));
	jor g0310(.dina(w_n624_0[1]),.dinb(n623),.dout(n625),.clk(gclk));
	jxor g0311(.dina(w_n625_1[1]),.dinb(w_n622_0[2]),.dout(n626),.clk(gclk));
	jnot g0312(.din(w_G3717_0[2]),.dout(n627),.clk(gclk));
	jand g0313(.dina(G236),.dinb(w_G18_43[0]),.dout(n628),.clk(gclk));
	jand g0314(.dina(G23),.dinb(w_n355_26[0]),.dout(n629),.clk(gclk));
	jor g0315(.dina(w_n629_0[1]),.dinb(n628),.dout(n630),.clk(gclk));
	jxor g0316(.dina(w_n630_0[2]),.dinb(w_n627_0[2]),.dout(n631),.clk(gclk));
	jnot g0317(.din(w_G3711_0[1]),.dout(n632),.clk(gclk));
	jand g0318(.dina(G237),.dinb(w_G18_42[2]),.dout(n633),.clk(gclk));
	jand g0319(.dina(G26),.dinb(w_n355_25[2]),.dout(n634),.clk(gclk));
	jor g0320(.dina(w_n634_0[1]),.dinb(n633),.dout(n635),.clk(gclk));
	jxor g0321(.dina(w_n635_1[1]),.dinb(w_n632_1[1]),.dout(n636),.clk(gclk));
	jnot g0322(.din(w_G238_0[1]),.dout(n637),.clk(gclk));
	jor g0323(.dina(n637),.dinb(w_n355_25[1]),.dout(n638),.clk(gclk));
	jnot g0324(.din(w_G29_0[1]),.dout(n639),.clk(gclk));
	jor g0325(.dina(n639),.dinb(w_G18_42[1]),.dout(n640),.clk(gclk));
	jand g0326(.dina(n640),.dinb(n638),.dout(n641),.clk(gclk));
	jxor g0327(.dina(w_n641_0[2]),.dinb(w_G3705_1[2]),.dout(n642),.clk(gclk));
	jand g0328(.dina(w_n642_0[2]),.dinb(w_n359_1[0]),.dout(n643),.clk(gclk));
	jand g0329(.dina(n643),.dinb(w_n636_0[2]),.dout(n644),.clk(gclk));
	jand g0330(.dina(w_n644_0[1]),.dinb(w_n631_0[2]),.dout(n645),.clk(gclk));
	jand g0331(.dina(w_n645_0[1]),.dinb(w_n626_1[1]),.dout(n646),.clk(gclk));
	jand g0332(.dina(w_n625_1[0]),.dinb(w_n622_0[1]),.dout(n647),.clk(gclk));
	jnot g0333(.din(w_n625_0[2]),.dout(n648),.clk(gclk));
	jand g0334(.dina(n648),.dinb(w_G3723_0[1]),.dout(n649),.clk(gclk));
	jnot g0335(.din(w_n649_0[1]),.dout(n650),.clk(gclk));
	jnot g0336(.din(w_n630_0[1]),.dout(n651),.clk(gclk));
	jand g0337(.dina(w_n651_0[1]),.dinb(w_G3717_0[1]),.dout(n652),.clk(gclk));
	jnot g0338(.din(w_n652_0[1]),.dout(n653),.clk(gclk));
	jand g0339(.dina(w_n630_0[0]),.dinb(w_n627_0[1]),.dout(n654),.clk(gclk));
	jand g0340(.dina(w_n635_1[0]),.dinb(w_n632_1[0]),.dout(n655),.clk(gclk));
	jor g0341(.dina(w_n635_0[2]),.dinb(w_n632_0[2]),.dout(n656),.clk(gclk));
	jnot g0342(.din(w_G3705_1[1]),.dout(n657),.clk(gclk));
	jand g0343(.dina(w_G238_0[0]),.dinb(w_G18_42[0]),.dout(n658),.clk(gclk));
	jand g0344(.dina(w_G29_0[0]),.dinb(w_n355_25[0]),.dout(n659),.clk(gclk));
	jor g0345(.dina(w_n659_0[1]),.dinb(n658),.dout(n660),.clk(gclk));
	jor g0346(.dina(w_n660_0[2]),.dinb(w_n657_0[2]),.dout(n661),.clk(gclk));
	jnot g0347(.din(w_G3701_0[2]),.dout(n662),.clk(gclk));
	jand g0348(.dina(w_G41_0[0]),.dinb(w_n355_24[2]),.dout(n663),.clk(gclk));
	jand g0349(.dina(w_n663_1[1]),.dinb(w_n662_0[1]),.dout(n664),.clk(gclk));
	jand g0350(.dina(w_n660_0[1]),.dinb(w_n657_0[1]),.dout(n665),.clk(gclk));
	jor g0351(.dina(n665),.dinb(w_n664_0[1]),.dout(n666),.clk(gclk));
	jand g0352(.dina(w_n666_0[1]),.dinb(w_n661_0[2]),.dout(n667),.clk(gclk));
	jand g0353(.dina(n667),.dinb(w_n656_0[1]),.dout(n668),.clk(gclk));
	jor g0354(.dina(n668),.dinb(w_n655_0[1]),.dout(n669),.clk(gclk));
	jor g0355(.dina(w_n669_0[1]),.dinb(w_n654_0[2]),.dout(n670),.clk(gclk));
	jand g0356(.dina(n670),.dinb(w_n653_0[1]),.dout(n671),.clk(gclk));
	jand g0357(.dina(w_n671_0[1]),.dinb(n650),.dout(n672),.clk(gclk));
	jor g0358(.dina(n672),.dinb(w_n647_0[1]),.dout(n673),.clk(gclk));
	jor g0359(.dina(w_n673_0[2]),.dinb(w_n646_0[1]),.dout(n674),.clk(gclk));
	jor g0360(.dina(w_n673_0[1]),.dinb(w_G4526_2[1]),.dout(n675),.clk(gclk));
	jand g0361(.dina(n675),.dinb(w_n674_0[1]),.dout(n676),.clk(gclk));
	jor g0362(.dina(w_n676_0[2]),.dinb(n621),.dout(n677),.clk(gclk));
	jand g0363(.dina(n677),.dinb(n620),.dout(n678),.clk(gclk));
	jand g0364(.dina(w_n678_0[1]),.dinb(n589),.dout(n679),.clk(gclk));
	jor g0365(.dina(n679),.dinb(w_n586_0[2]),.dout(n680),.clk(gclk));
	jand g0366(.dina(w_n680_2[2]),.dinb(w_n581_0[2]),.dout(n681),.clk(gclk));
	jor g0367(.dina(n681),.dinb(w_n572_1[1]),.dout(n682),.clk(gclk));
	jand g0368(.dina(w_n682_0[1]),.dinb(n527),.dout(n683),.clk(gclk));
	jand g0369(.dina(w_n683_0[1]),.dinb(w_n524_1[2]),.dout(n684),.clk(gclk));
	jand g0370(.dina(n684),.dinb(n519),.dout(n685),.clk(gclk));
	jand g0371(.dina(n685),.dinb(w_n513_1[1]),.dout(n686),.clk(gclk));
	jand g0372(.dina(w_n512_0[1]),.dinb(w_n509_0[1]),.dout(n687),.clk(gclk));
	jnot g0373(.din(w_n687_0[1]),.dout(n688),.clk(gclk));
	jnot g0374(.din(w_n512_0[0]),.dout(n689),.clk(gclk));
	jand g0375(.dina(w_n689_0[1]),.dinb(w_G4432_0[1]),.dout(n690),.clk(gclk));
	jand g0376(.dina(w_n523_0[1]),.dinb(w_n520_0[0]),.dout(n691),.clk(gclk));
	jand g0377(.dina(w_n524_1[1]),.dinb(w_n518_1[1]),.dout(n692),.clk(gclk));
	jor g0378(.dina(n692),.dinb(n691),.dout(n693),.clk(gclk));
	jnot g0379(.din(w_n693_0[1]),.dout(n694),.clk(gclk));
	jor g0380(.dina(w_n694_0[1]),.dinb(w_n690_0[1]),.dout(n695),.clk(gclk));
	jand g0381(.dina(w_n695_0[1]),.dinb(n688),.dout(n696),.clk(gclk));
	jnot g0382(.din(w_n696_0[1]),.dout(n697),.clk(gclk));
	jor g0383(.dina(n697),.dinb(n686),.dout(n698),.clk(gclk));
	jand g0384(.dina(w_n698_0[1]),.dinb(n508),.dout(n699),.clk(gclk));
	jor g0385(.dina(n699),.dinb(w_n505_0[1]),.dout(n700),.clk(gclk));
	jor g0386(.dina(w_n700_1[1]),.dinb(w_n462_0[1]),.dout(n701),.clk(gclk));
	jor g0387(.dina(n701),.dinb(w_n500_0[1]),.dout(n702),.clk(gclk));
	jand g0388(.dina(n702),.dinb(w_n499_0[1]),.dout(n703),.clk(gclk));
	jor g0389(.dina(w_n703_1[2]),.dinb(w_n449_1[0]),.dout(n704),.clk(gclk));
	jand g0390(.dina(n704),.dinb(w_n450_0[2]),.dout(n705),.clk(gclk));
	jand g0391(.dina(w_n705_0[1]),.dinb(w_n425_1[1]),.dout(n706),.clk(gclk));
	jor g0392(.dina(n706),.dinb(w_n424_0[1]),.dout(n707),.clk(gclk));
	jor g0393(.dina(w_n707_1[2]),.dinb(w_n413_1[0]),.dout(n708),.clk(gclk));
	jand g0394(.dina(n708),.dinb(w_n420_0[1]),.dout(n709),.clk(gclk));
	jand g0395(.dina(w_n709_1[1]),.dinb(w_n370_0[2]),.dout(n710),.clk(gclk));
	jand g0396(.dina(n710),.dinb(w_n363_0[2]),.dout(n711),.clk(gclk));
	jnot g0397(.din(w_n362_0[1]),.dout(n712),.clk(gclk));
	jand g0398(.dina(w_n712_0[2]),.dinb(w_G38_2[0]),.dout(n713),.clk(gclk));
	jand g0399(.dina(w_n366_0[1]),.dinb(w_G38_1[2]),.dout(n714),.clk(gclk));
	jor g0400(.dina(n714),.dinb(w_n713_0[1]),.dout(n715),.clk(gclk));
	jor g0401(.dina(w_n715_1[1]),.dinb(w_n711_1[1]),.dout(G246),.clk(gclk));
	jand g0402(.dina(w_G2204_0[2]),.dinb(w_G1455_0[2]),.dout(n717),.clk(gclk));
	jor g0403(.dina(n717),.dinb(w_n368_0[0]),.dout(n718),.clk(gclk));
	jor g0404(.dina(G166),.dinb(w_n355_24[1]),.dout(n719),.clk(gclk));
	jand g0405(.dina(w_n719_0[1]),.dinb(w_n373_6[1]),.dout(n720),.clk(gclk));
	jor g0406(.dina(w_n371_0[0]),.dinb(w_n355_24[0]),.dout(n721),.clk(gclk));
	jor g0407(.dina(G88),.dinb(w_G18_41[2]),.dout(n722),.clk(gclk));
	jand g0408(.dina(n722),.dinb(n721),.dout(n723),.clk(gclk));
	jxor g0409(.dina(w_n723_0[2]),.dinb(w_n720_0[2]),.dout(n724),.clk(gclk));
	jor g0410(.dina(G167),.dinb(w_n355_23[2]),.dout(n725),.clk(gclk));
	jand g0411(.dina(w_n725_0[1]),.dinb(w_n373_6[0]),.dout(n726),.clk(gclk));
	jor g0412(.dina(w_n383_0[0]),.dinb(w_n355_23[1]),.dout(n727),.clk(gclk));
	jor g0413(.dina(G112),.dinb(w_G18_41[1]),.dout(n728),.clk(gclk));
	jand g0414(.dina(n728),.dinb(n727),.dout(n729),.clk(gclk));
	jor g0415(.dina(w_n729_1[1]),.dinb(w_n726_1[1]),.dout(n730),.clk(gclk));
	jand g0416(.dina(w_n729_1[0]),.dinb(w_n726_1[0]),.dout(n731),.clk(gclk));
	jor g0417(.dina(w_n389_0[2]),.dinb(w_n355_23[0]),.dout(n732),.clk(gclk));
	jor g0418(.dina(G113),.dinb(w_G18_41[0]),.dout(n733),.clk(gclk));
	jand g0419(.dina(n733),.dinb(n732),.dout(n734),.clk(gclk));
	jand g0420(.dina(w_n734_0[2]),.dinb(w_n373_5[2]),.dout(n735),.clk(gclk));
	jor g0421(.dina(G168),.dinb(w_n355_22[2]),.dout(n736),.clk(gclk));
	jand g0422(.dina(w_n736_0[1]),.dinb(w_n373_5[1]),.dout(n737),.clk(gclk));
	jand g0423(.dina(w_G106_0[2]),.dinb(w_G18_40[2]),.dout(n738),.clk(gclk));
	jnot g0424(.din(n738),.dout(n739),.clk(gclk));
	jor g0425(.dina(G87),.dinb(w_G18_40[1]),.dout(n740),.clk(gclk));
	jand g0426(.dina(n740),.dinb(n739),.dout(n741),.clk(gclk));
	jxor g0427(.dina(w_n741_1[1]),.dinb(w_n737_1[1]),.dout(n742),.clk(gclk));
	jor g0428(.dina(G169),.dinb(w_n355_22[1]),.dout(n743),.clk(gclk));
	jand g0429(.dina(w_n743_0[1]),.dinb(w_n373_5[0]),.dout(n744),.clk(gclk));
	jor g0430(.dina(w_n393_0[2]),.dinb(w_n355_22[0]),.dout(n745),.clk(gclk));
	jor g0431(.dina(G111),.dinb(w_G18_40[0]),.dout(n746),.clk(gclk));
	jand g0432(.dina(n746),.dinb(n745),.dout(n747),.clk(gclk));
	jxor g0433(.dina(w_n747_0[2]),.dinb(w_n744_0[2]),.dout(n748),.clk(gclk));
	jand g0434(.dina(n748),.dinb(n742),.dout(n749),.clk(gclk));
	jand g0435(.dina(w_n749_0[1]),.dinb(n735),.dout(n750),.clk(gclk));
	jor g0436(.dina(n750),.dinb(n731),.dout(n751),.clk(gclk));
	jand g0437(.dina(n751),.dinb(n730),.dout(n752),.clk(gclk));
	jand g0438(.dina(n752),.dinb(w_n724_0[1]),.dout(n753),.clk(gclk));
	jor g0439(.dina(G173),.dinb(w_n355_21[2]),.dout(n754),.clk(gclk));
	jand g0440(.dina(w_n754_0[1]),.dinb(w_n373_4[2]),.dout(n755),.clk(gclk));
	jor g0441(.dina(w_n421_0[0]),.dinb(w_n355_21[1]),.dout(n756),.clk(gclk));
	jor g0442(.dina(G110),.dinb(w_G18_39[2]),.dout(n757),.clk(gclk));
	jand g0443(.dina(n757),.dinb(n756),.dout(n758),.clk(gclk));
	jxor g0444(.dina(w_n758_1[1]),.dinb(w_n755_1[1]),.dout(n759),.clk(gclk));
	jor g0445(.dina(G174),.dinb(w_n355_21[0]),.dout(n760),.clk(gclk));
	jand g0446(.dina(w_n760_0[1]),.dinb(w_n373_4[1]),.dout(n761),.clk(gclk));
	jor g0447(.dina(w_n426_0[0]),.dinb(w_n355_20[2]),.dout(n762),.clk(gclk));
	jor g0448(.dina(G109),.dinb(w_G18_39[1]),.dout(n763),.clk(gclk));
	jand g0449(.dina(n763),.dinb(n762),.dout(n764),.clk(gclk));
	jxor g0450(.dina(w_n764_0[2]),.dinb(w_n761_0[2]),.dout(n765),.clk(gclk));
	jand g0451(.dina(n765),.dinb(n759),.dout(n766),.clk(gclk));
	jor g0452(.dina(G175),.dinb(w_n355_20[1]),.dout(n767),.clk(gclk));
	jand g0453(.dina(w_n767_0[1]),.dinb(w_n373_4[0]),.dout(n768),.clk(gclk));
	jand g0454(.dina(w_G2247_0[1]),.dinb(w_G18_39[0]),.dout(n769),.clk(gclk));
	jnot g0455(.din(n769),.dout(n770),.clk(gclk));
	jor g0456(.dina(G86),.dinb(w_G18_38[2]),.dout(n771),.clk(gclk));
	jand g0457(.dina(n771),.dinb(n770),.dout(n772),.clk(gclk));
	jand g0458(.dina(w_n772_0[2]),.dinb(w_n768_0[2]),.dout(n773),.clk(gclk));
	jor g0459(.dina(w_n772_0[1]),.dinb(w_n768_0[1]),.dout(n774),.clk(gclk));
	jor g0460(.dina(G176),.dinb(w_n355_20[0]),.dout(n775),.clk(gclk));
	jand g0461(.dina(w_n775_0[1]),.dinb(w_n373_3[2]),.dout(n776),.clk(gclk));
	jand g0462(.dina(w_G2239_1[0]),.dinb(w_G18_38[1]),.dout(n777),.clk(gclk));
	jnot g0463(.din(n777),.dout(n778),.clk(gclk));
	jor g0464(.dina(G63),.dinb(w_G18_38[0]),.dout(n779),.clk(gclk));
	jand g0465(.dina(n779),.dinb(n778),.dout(n780),.clk(gclk));
	jand g0466(.dina(w_n780_0[2]),.dinb(w_n776_0[2]),.dout(n781),.clk(gclk));
	jand g0467(.dina(w_n781_0[1]),.dinb(w_n774_0[1]),.dout(n782),.clk(gclk));
	jor g0468(.dina(n782),.dinb(w_n773_0[1]),.dout(n783),.clk(gclk));
	jand g0469(.dina(n783),.dinb(w_n766_0[1]),.dout(n784),.clk(gclk));
	jand g0470(.dina(w_n758_1[0]),.dinb(w_n755_1[0]),.dout(n785),.clk(gclk));
	jor g0471(.dina(w_n758_0[2]),.dinb(w_n755_0[2]),.dout(n786),.clk(gclk));
	jand g0472(.dina(w_n764_0[1]),.dinb(w_n761_0[1]),.dout(n787),.clk(gclk));
	jand g0473(.dina(n787),.dinb(n786),.dout(n788),.clk(gclk));
	jor g0474(.dina(n788),.dinb(n785),.dout(n789),.clk(gclk));
	jor g0475(.dina(n789),.dinb(n784),.dout(n790),.clk(gclk));
	jnot g0476(.din(w_n773_0[0]),.dout(n791),.clk(gclk));
	jnot g0477(.din(w_n781_0[0]),.dout(n792),.clk(gclk));
	jand g0478(.dina(n792),.dinb(n791),.dout(n793),.clk(gclk));
	jand g0479(.dina(n793),.dinb(w_n766_0[0]),.dout(n794),.clk(gclk));
	jor g0480(.dina(G177),.dinb(w_n355_19[2]),.dout(n795),.clk(gclk));
	jand g0481(.dina(n795),.dinb(w_n373_3[1]),.dout(n796),.clk(gclk));
	jand g0482(.dina(w_G2236_0[1]),.dinb(w_G18_37[2]),.dout(n797),.clk(gclk));
	jnot g0483(.din(n797),.dout(n798),.clk(gclk));
	jor g0484(.dina(G64),.dinb(w_G18_37[1]),.dout(n799),.clk(gclk));
	jand g0485(.dina(n799),.dinb(n798),.dout(n800),.clk(gclk));
	jxor g0486(.dina(w_n800_1[1]),.dinb(w_n796_1[1]),.dout(n801),.clk(gclk));
	jand g0487(.dina(G178),.dinb(w_G18_37[0]),.dout(n802),.clk(gclk));
	jor g0488(.dina(n802),.dinb(w_n457_0[0]),.dout(n803),.clk(gclk));
	jor g0489(.dina(w_n456_0[0]),.dinb(w_n355_19[1]),.dout(n804),.clk(gclk));
	jor g0490(.dina(G85),.dinb(w_G18_36[2]),.dout(n805),.clk(gclk));
	jand g0491(.dina(n805),.dinb(n804),.dout(n806),.clk(gclk));
	jxor g0492(.dina(w_n806_0[2]),.dinb(w_n803_0[2]),.dout(n807),.clk(gclk));
	jand g0493(.dina(n807),.dinb(n801),.dout(n808),.clk(gclk));
	jand g0494(.dina(G179),.dinb(w_G18_36[1]),.dout(n809),.clk(gclk));
	jor g0495(.dina(n809),.dinb(w_n467_0[0]),.dout(n810),.clk(gclk));
	jand g0496(.dina(w_G2224_0[2]),.dinb(w_G18_36[0]),.dout(n811),.clk(gclk));
	jnot g0497(.din(n811),.dout(n812),.clk(gclk));
	jor g0498(.dina(G84),.dinb(w_G18_35[2]),.dout(n813),.clk(gclk));
	jand g0499(.dina(n813),.dinb(n812),.dout(n814),.clk(gclk));
	jxor g0500(.dina(w_n814_1[1]),.dinb(w_n810_1[1]),.dout(n815),.clk(gclk));
	jand g0501(.dina(G180),.dinb(w_G18_35[1]),.dout(n816),.clk(gclk));
	jor g0502(.dina(n816),.dinb(w_n472_0[0]),.dout(n817),.clk(gclk));
	jor g0503(.dina(w_n471_0[0]),.dinb(w_n355_19[0]),.dout(n818),.clk(gclk));
	jor g0504(.dina(G83),.dinb(w_G18_35[0]),.dout(n819),.clk(gclk));
	jand g0505(.dina(n819),.dinb(n818),.dout(n820),.clk(gclk));
	jxor g0506(.dina(w_n820_0[2]),.dinb(w_n817_0[2]),.dout(n821),.clk(gclk));
	jand g0507(.dina(n821),.dinb(n815),.dout(n822),.clk(gclk));
	jand g0508(.dina(G171),.dinb(w_G18_34[2]),.dout(n823),.clk(gclk));
	jor g0509(.dina(n823),.dinb(w_n477_0[0]),.dout(n824),.clk(gclk));
	jor g0510(.dina(w_n476_0[0]),.dinb(w_n355_18[2]),.dout(n825),.clk(gclk));
	jor g0511(.dina(G65),.dinb(w_G18_34[1]),.dout(n826),.clk(gclk));
	jand g0512(.dina(n826),.dinb(n825),.dout(n827),.clk(gclk));
	jand g0513(.dina(w_n827_0[2]),.dinb(w_n824_0[2]),.dout(n828),.clk(gclk));
	jand g0514(.dina(n828),.dinb(w_n822_0[1]),.dout(n829),.clk(gclk));
	jand g0515(.dina(w_n814_1[0]),.dinb(w_n810_1[0]),.dout(n830),.clk(gclk));
	jor g0516(.dina(w_n814_0[2]),.dinb(w_n810_0[2]),.dout(n831),.clk(gclk));
	jand g0517(.dina(w_n820_0[1]),.dinb(w_n817_0[1]),.dout(n832),.clk(gclk));
	jand g0518(.dina(n832),.dinb(n831),.dout(n833),.clk(gclk));
	jor g0519(.dina(n833),.dinb(n830),.dout(n834),.clk(gclk));
	jor g0520(.dina(n834),.dinb(n829),.dout(n835),.clk(gclk));
	jand g0521(.dina(n835),.dinb(w_n808_0[1]),.dout(n836),.clk(gclk));
	jand g0522(.dina(w_n800_1[0]),.dinb(w_n796_1[0]),.dout(n837),.clk(gclk));
	jor g0523(.dina(w_n800_0[2]),.dinb(w_n796_0[2]),.dout(n838),.clk(gclk));
	jand g0524(.dina(w_n806_0[1]),.dinb(w_n803_0[1]),.dout(n839),.clk(gclk));
	jand g0525(.dina(n839),.dinb(n838),.dout(n840),.clk(gclk));
	jor g0526(.dina(n840),.dinb(n837),.dout(n841),.clk(gclk));
	jor g0527(.dina(n841),.dinb(n836),.dout(n842),.clk(gclk));
	jand g0528(.dina(w_n822_0[0]),.dinb(w_n808_0[0]),.dout(n843),.clk(gclk));
	jand g0529(.dina(G189),.dinb(w_G18_34[0]),.dout(n844),.clk(gclk));
	jor g0530(.dina(n844),.dinb(w_n503_0[0]),.dout(n845),.clk(gclk));
	jor g0531(.dina(w_n501_0[1]),.dinb(w_n355_18[1]),.dout(n846),.clk(gclk));
	jor g0532(.dina(G62),.dinb(w_G18_33[2]),.dout(n847),.clk(gclk));
	jand g0533(.dina(n847),.dinb(n846),.dout(n848),.clk(gclk));
	jxor g0534(.dina(w_n848_1[1]),.dinb(w_n845_1[1]),.dout(n849),.clk(gclk));
	jand g0535(.dina(G190),.dinb(w_G18_33[1]),.dout(n850),.clk(gclk));
	jor g0536(.dina(n850),.dinb(w_n511_0[0]),.dout(n851),.clk(gclk));
	jor g0537(.dina(w_n509_0[0]),.dinb(w_n355_18[0]),.dout(n852),.clk(gclk));
	jor g0538(.dina(G61),.dinb(w_G18_33[0]),.dout(n853),.clk(gclk));
	jand g0539(.dina(n853),.dinb(n852),.dout(n854),.clk(gclk));
	jxor g0540(.dina(w_n854_0[2]),.dinb(w_n851_0[2]),.dout(n855),.clk(gclk));
	jand g0541(.dina(n855),.dinb(n849),.dout(n856),.clk(gclk));
	jand g0542(.dina(G191),.dinb(w_G18_32[2]),.dout(n857),.clk(gclk));
	jor g0543(.dina(n857),.dinb(w_n522_0[0]),.dout(n858),.clk(gclk));
	jand g0544(.dina(w_G4427_0[1]),.dinb(w_G18_32[1]),.dout(n859),.clk(gclk));
	jnot g0545(.din(n859),.dout(n860),.clk(gclk));
	jor g0546(.dina(G60),.dinb(w_G18_32[0]),.dout(n861),.clk(gclk));
	jand g0547(.dina(n861),.dinb(n860),.dout(n862),.clk(gclk));
	jand g0548(.dina(w_n862_0[2]),.dinb(w_n858_0[2]),.dout(n863),.clk(gclk));
	jor g0549(.dina(w_n862_0[1]),.dinb(w_n858_0[1]),.dout(n864),.clk(gclk));
	jand g0550(.dina(G192),.dinb(w_G18_31[2]),.dout(n865),.clk(gclk));
	jor g0551(.dina(n865),.dinb(w_n516_0[0]),.dout(n866),.clk(gclk));
	jand g0552(.dina(w_G4420_0[2]),.dinb(w_G18_31[1]),.dout(n867),.clk(gclk));
	jnot g0553(.din(n867),.dout(n868),.clk(gclk));
	jor g0554(.dina(G79),.dinb(w_G18_31[0]),.dout(n869),.clk(gclk));
	jand g0555(.dina(n869),.dinb(n868),.dout(n870),.clk(gclk));
	jand g0556(.dina(w_n870_0[2]),.dinb(w_n866_0[2]),.dout(n871),.clk(gclk));
	jand g0557(.dina(w_n871_0[1]),.dinb(w_n864_0[1]),.dout(n872),.clk(gclk));
	jor g0558(.dina(n872),.dinb(w_n863_0[1]),.dout(n873),.clk(gclk));
	jand g0559(.dina(n873),.dinb(w_n856_0[1]),.dout(n874),.clk(gclk));
	jand g0560(.dina(w_n848_1[0]),.dinb(w_n845_1[0]),.dout(n875),.clk(gclk));
	jor g0561(.dina(w_n848_0[2]),.dinb(w_n845_0[2]),.dout(n876),.clk(gclk));
	jand g0562(.dina(w_n854_0[1]),.dinb(w_n851_0[1]),.dout(n877),.clk(gclk));
	jand g0563(.dina(n877),.dinb(n876),.dout(n878),.clk(gclk));
	jor g0564(.dina(n878),.dinb(n875),.dout(n879),.clk(gclk));
	jor g0565(.dina(n879),.dinb(n874),.dout(n880),.clk(gclk));
	jor g0566(.dina(w_n870_0[1]),.dinb(w_n866_0[1]),.dout(n881),.clk(gclk));
	jand g0567(.dina(n881),.dinb(w_n864_0[0]),.dout(n882),.clk(gclk));
	jand g0568(.dina(n882),.dinb(w_n856_0[0]),.dout(n883),.clk(gclk));
	jand g0569(.dina(G205),.dinb(w_G18_30[2]),.dout(n884),.clk(gclk));
	jor g0570(.dina(n884),.dinb(w_n629_0[0]),.dout(n885),.clk(gclk));
	jor g0571(.dina(w_n627_0[0]),.dinb(w_n355_17[2]),.dout(n886),.clk(gclk));
	jor g0572(.dina(G75),.dinb(w_G18_30[1]),.dout(n887),.clk(gclk));
	jand g0573(.dina(n887),.dinb(n886),.dout(n888),.clk(gclk));
	jor g0574(.dina(w_n888_0[2]),.dinb(w_n885_0[2]),.dout(n889),.clk(gclk));
	jand g0575(.dina(G206),.dinb(w_G18_30[0]),.dout(n890),.clk(gclk));
	jor g0576(.dina(n890),.dinb(w_n634_0[0]),.dout(n891),.clk(gclk));
	jor g0577(.dina(w_n632_0[1]),.dinb(w_n355_17[1]),.dout(n892),.clk(gclk));
	jor g0578(.dina(G76),.dinb(w_G18_29[2]),.dout(n893),.clk(gclk));
	jand g0579(.dina(n893),.dinb(n892),.dout(n894),.clk(gclk));
	jand g0580(.dina(w_n894_0[2]),.dinb(w_n891_0[2]),.dout(n895),.clk(gclk));
	jor g0581(.dina(w_G89_0[1]),.dinb(w_G70_0[1]),.dout(n896),.clk(gclk));
	jand g0582(.dina(n896),.dinb(w_n663_1[0]),.dout(n897),.clk(gclk));
	jor g0583(.dina(n897),.dinb(w_n895_0[1]),.dout(n898),.clk(gclk));
	jand g0584(.dina(G207),.dinb(w_G18_29[1]),.dout(n899),.clk(gclk));
	jor g0585(.dina(n899),.dinb(w_n659_0[0]),.dout(n900),.clk(gclk));
	jor g0586(.dina(w_n657_0[0]),.dinb(w_n355_17[0]),.dout(n901),.clk(gclk));
	jor g0587(.dina(G74),.dinb(w_G18_29[0]),.dout(n902),.clk(gclk));
	jand g0588(.dina(n902),.dinb(n901),.dout(n903),.clk(gclk));
	jand g0589(.dina(w_n903_0[2]),.dinb(w_n900_0[2]),.dout(n904),.clk(gclk));
	jor g0590(.dina(w_G70_0[0]),.dinb(w_G18_28[2]),.dout(n905),.clk(gclk));
	jand g0591(.dina(w_n905_0[1]),.dinb(w_G89_0[0]),.dout(n906),.clk(gclk));
	jor g0592(.dina(n906),.dinb(n904),.dout(n907),.clk(gclk));
	jor g0593(.dina(n907),.dinb(n898),.dout(n908),.clk(gclk));
	jor g0594(.dina(w_n903_0[1]),.dinb(w_n900_0[1]),.dout(n909),.clk(gclk));
	jor g0595(.dina(w_n894_0[1]),.dinb(w_n891_0[1]),.dout(n910),.clk(gclk));
	jand g0596(.dina(n910),.dinb(n909),.dout(n911),.clk(gclk));
	jor g0597(.dina(n911),.dinb(w_n895_0[0]),.dout(n912),.clk(gclk));
	jand g0598(.dina(n912),.dinb(n908),.dout(n913),.clk(gclk));
	jand g0599(.dina(n913),.dinb(n889),.dout(n914),.clk(gclk));
	jand g0600(.dina(G204),.dinb(w_G18_28[1]),.dout(n915),.clk(gclk));
	jor g0601(.dina(n915),.dinb(w_n624_0[0]),.dout(n916),.clk(gclk));
	jor g0602(.dina(w_n622_0[0]),.dinb(w_n355_16[2]),.dout(n917),.clk(gclk));
	jor g0603(.dina(G73),.dinb(w_G18_28[0]),.dout(n918),.clk(gclk));
	jand g0604(.dina(n918),.dinb(n917),.dout(n919),.clk(gclk));
	jand g0605(.dina(w_n919_0[2]),.dinb(w_n916_0[2]),.dout(n920),.clk(gclk));
	jand g0606(.dina(w_n888_0[1]),.dinb(w_n885_0[1]),.dout(n921),.clk(gclk));
	jor g0607(.dina(n921),.dinb(n920),.dout(n922),.clk(gclk));
	jor g0608(.dina(n922),.dinb(n914),.dout(n923),.clk(gclk));
	jor g0609(.dina(w_n919_0[1]),.dinb(w_n916_0[1]),.dout(n924),.clk(gclk));
	jand g0610(.dina(G203),.dinb(w_G18_27[2]),.dout(n925),.clk(gclk));
	jor g0611(.dina(n925),.dinb(w_n602_0[0]),.dout(n926),.clk(gclk));
	jand g0612(.dina(w_G3729_1[0]),.dinb(w_G18_27[1]),.dout(n927),.clk(gclk));
	jnot g0613(.din(n927),.dout(n928),.clk(gclk));
	jor g0614(.dina(G53),.dinb(w_G18_27[0]),.dout(n929),.clk(gclk));
	jand g0615(.dina(n929),.dinb(n928),.dout(n930),.clk(gclk));
	jor g0616(.dina(w_n930_0[2]),.dinb(w_n926_0[2]),.dout(n931),.clk(gclk));
	jand g0617(.dina(n931),.dinb(n924),.dout(n932),.clk(gclk));
	jand g0618(.dina(n932),.dinb(n923),.dout(n933),.clk(gclk));
	jand g0619(.dina(G202),.dinb(w_G18_26[2]),.dout(n934),.clk(gclk));
	jor g0620(.dina(n934),.dinb(w_n597_0[0]),.dout(n935),.clk(gclk));
	jor g0621(.dina(w_n595_0[0]),.dinb(w_n355_16[1]),.dout(n936),.clk(gclk));
	jor g0622(.dina(G54),.dinb(w_G18_26[1]),.dout(n937),.clk(gclk));
	jand g0623(.dina(n937),.dinb(n936),.dout(n938),.clk(gclk));
	jand g0624(.dina(w_n938_0[2]),.dinb(w_n935_0[2]),.dout(n939),.clk(gclk));
	jand g0625(.dina(w_n930_0[1]),.dinb(w_n926_0[1]),.dout(n940),.clk(gclk));
	jor g0626(.dina(n940),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0627(.dina(n941),.dinb(n933),.dout(n942),.clk(gclk));
	jand g0628(.dina(G201),.dinb(w_G18_26[0]),.dout(n943),.clk(gclk));
	jor g0629(.dina(n943),.dinb(w_n592_0[0]),.dout(n944),.clk(gclk));
	jor g0630(.dina(w_n590_0[0]),.dinb(w_n355_16[0]),.dout(n945),.clk(gclk));
	jor g0631(.dina(G55),.dinb(w_G18_25[2]),.dout(n946),.clk(gclk));
	jand g0632(.dina(n946),.dinb(n945),.dout(n947),.clk(gclk));
	jxor g0633(.dina(w_n947_0[2]),.dinb(w_n944_0[2]),.dout(n948),.clk(gclk));
	jand g0634(.dina(G200),.dinb(w_G18_25[1]),.dout(n949),.clk(gclk));
	jor g0635(.dina(n949),.dinb(w_n584_0[0]),.dout(n950),.clk(gclk));
	jor g0636(.dina(w_n582_0[1]),.dinb(w_n355_15[2]),.dout(n951),.clk(gclk));
	jor g0637(.dina(G56),.dinb(w_G18_25[0]),.dout(n952),.clk(gclk));
	jand g0638(.dina(n952),.dinb(n951),.dout(n953),.clk(gclk));
	jxor g0639(.dina(w_n953_1[1]),.dinb(w_n950_1[1]),.dout(n954),.clk(gclk));
	jand g0640(.dina(n954),.dinb(n948),.dout(n955),.clk(gclk));
	jor g0641(.dina(w_n938_0[1]),.dinb(w_n935_0[1]),.dout(n956),.clk(gclk));
	jand g0642(.dina(n956),.dinb(n955),.dout(n957),.clk(gclk));
	jand g0643(.dina(n957),.dinb(n942),.dout(n958),.clk(gclk));
	jand g0644(.dina(w_n953_1[0]),.dinb(w_n950_1[0]),.dout(n959),.clk(gclk));
	jand g0645(.dina(w_n947_0[1]),.dinb(w_n944_0[1]),.dout(n960),.clk(gclk));
	jor g0646(.dina(w_n953_0[2]),.dinb(w_n950_0[2]),.dout(n961),.clk(gclk));
	jand g0647(.dina(n961),.dinb(n960),.dout(n962),.clk(gclk));
	jor g0648(.dina(n962),.dinb(n959),.dout(n963),.clk(gclk));
	jor g0649(.dina(n963),.dinb(n958),.dout(n964),.clk(gclk));
	jand g0650(.dina(G187),.dinb(w_G18_24[2]),.dout(n965),.clk(gclk));
	jor g0651(.dina(n965),.dinb(w_n562_0[0]),.dout(n966),.clk(gclk));
	jand g0652(.dina(w_G4394_1[0]),.dinb(w_G18_24[1]),.dout(n967),.clk(gclk));
	jnot g0653(.din(n967),.dout(n968),.clk(gclk));
	jor g0654(.dina(G77),.dinb(w_G18_24[0]),.dout(n969),.clk(gclk));
	jand g0655(.dina(n969),.dinb(n968),.dout(n970),.clk(gclk));
	jor g0656(.dina(w_n970_0[2]),.dinb(w_n966_0[2]),.dout(n971),.clk(gclk));
	jand g0657(.dina(G193),.dinb(w_G18_23[2]),.dout(n972),.clk(gclk));
	jor g0658(.dina(n972),.dinb(w_n530_0[0]),.dout(n973),.clk(gclk));
	jand g0659(.dina(w_G4415_0[2]),.dinb(w_G18_23[1]),.dout(n974),.clk(gclk));
	jnot g0660(.din(n974),.dout(n975),.clk(gclk));
	jor g0661(.dina(G80),.dinb(w_G18_23[0]),.dout(n976),.clk(gclk));
	jand g0662(.dina(n976),.dinb(n975),.dout(n977),.clk(gclk));
	jxor g0663(.dina(w_n977_1[1]),.dinb(w_n973_1[1]),.dout(n978),.clk(gclk));
	jand g0664(.dina(G194),.dinb(w_G18_22[2]),.dout(n979),.clk(gclk));
	jor g0665(.dina(n979),.dinb(w_n538_0[0]),.dout(n980),.clk(gclk));
	jor g0666(.dina(w_n536_0[0]),.dinb(w_n355_15[1]),.dout(n981),.clk(gclk));
	jor g0667(.dina(G81),.dinb(w_G18_22[1]),.dout(n982),.clk(gclk));
	jand g0668(.dina(n982),.dinb(n981),.dout(n983),.clk(gclk));
	jxor g0669(.dina(w_n983_0[2]),.dinb(w_n980_0[2]),.dout(n984),.clk(gclk));
	jand g0670(.dina(n984),.dinb(n978),.dout(n985),.clk(gclk));
	jand g0671(.dina(G196),.dinb(w_G18_22[0]),.dout(n986),.clk(gclk));
	jor g0672(.dina(n986),.dinb(w_n554_0[0]),.dout(n987),.clk(gclk));
	jand g0673(.dina(w_G4400_0[2]),.dinb(w_G18_21[2]),.dout(n988),.clk(gclk));
	jnot g0674(.din(n988),.dout(n989),.clk(gclk));
	jor g0675(.dina(G78),.dinb(w_G18_21[1]),.dout(n990),.clk(gclk));
	jand g0676(.dina(n990),.dinb(n989),.dout(n991),.clk(gclk));
	jand g0677(.dina(w_n991_0[2]),.dinb(w_n987_0[2]),.dout(n992),.clk(gclk));
	jnot g0678(.din(w_n992_0[1]),.dout(n993),.clk(gclk));
	jand g0679(.dina(G195),.dinb(w_G18_21[0]),.dout(n994),.clk(gclk));
	jor g0680(.dina(n994),.dinb(w_n546_0[0]),.dout(n995),.clk(gclk));
	jand g0681(.dina(w_G4405_0[2]),.dinb(w_G18_20[2]),.dout(n996),.clk(gclk));
	jnot g0682(.din(n996),.dout(n997),.clk(gclk));
	jor g0683(.dina(G59),.dinb(w_G18_20[1]),.dout(n998),.clk(gclk));
	jand g0684(.dina(n998),.dinb(n997),.dout(n999),.clk(gclk));
	jor g0685(.dina(w_n999_0[2]),.dinb(w_n995_0[2]),.dout(n1000),.clk(gclk));
	jand g0686(.dina(w_n1000_0[1]),.dinb(n993),.dout(n1001),.clk(gclk));
	jor g0687(.dina(w_n991_0[1]),.dinb(w_n987_0[1]),.dout(n1002),.clk(gclk));
	jand g0688(.dina(w_n999_0[1]),.dinb(w_n995_0[1]),.dout(n1003),.clk(gclk));
	jnot g0689(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0690(.dina(n1004),.dinb(n1002),.dout(n1005),.clk(gclk));
	jand g0691(.dina(n1005),.dinb(n1001),.dout(n1006),.clk(gclk));
	jand g0692(.dina(n1006),.dinb(w_n985_0[1]),.dout(n1007),.clk(gclk));
	jand g0693(.dina(w_n970_0[1]),.dinb(w_n966_0[1]),.dout(n1008),.clk(gclk));
	jnot g0694(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jand g0695(.dina(n1009),.dinb(w_n1007_0[1]),.dout(n1010),.clk(gclk));
	jand g0696(.dina(n1010),.dinb(n971),.dout(n1011),.clk(gclk));
	jand g0697(.dina(n1011),.dinb(n964),.dout(n1012),.clk(gclk));
	jand g0698(.dina(w_n977_1[0]),.dinb(w_n973_1[0]),.dout(n1013),.clk(gclk));
	jor g0699(.dina(w_n977_0[2]),.dinb(w_n973_0[2]),.dout(n1014),.clk(gclk));
	jand g0700(.dina(w_n983_0[1]),.dinb(w_n980_0[1]),.dout(n1015),.clk(gclk));
	jand g0701(.dina(n1015),.dinb(n1014),.dout(n1016),.clk(gclk));
	jor g0702(.dina(n1016),.dinb(n1013),.dout(n1017),.clk(gclk));
	jand g0703(.dina(w_n1008_0[0]),.dinb(w_n1007_0[0]),.dout(n1018),.clk(gclk));
	jand g0704(.dina(w_n1000_0[0]),.dinb(w_n992_0[0]),.dout(n1019),.clk(gclk));
	jor g0705(.dina(n1019),.dinb(w_n1003_0[0]),.dout(n1020),.clk(gclk));
	jand g0706(.dina(n1020),.dinb(w_n985_0[0]),.dout(n1021),.clk(gclk));
	jor g0707(.dina(n1021),.dinb(n1018),.dout(n1022),.clk(gclk));
	jor g0708(.dina(n1022),.dinb(n1017),.dout(n1023),.clk(gclk));
	jor g0709(.dina(n1023),.dinb(n1012),.dout(n1024),.clk(gclk));
	jnot g0710(.din(w_n863_0[0]),.dout(n1025),.clk(gclk));
	jnot g0711(.din(w_n871_0[0]),.dout(n1026),.clk(gclk));
	jand g0712(.dina(n1026),.dinb(n1025),.dout(n1027),.clk(gclk));
	jand g0713(.dina(n1027),.dinb(n1024),.dout(n1028),.clk(gclk));
	jand g0714(.dina(n1028),.dinb(n883),.dout(n1029),.clk(gclk));
	jor g0715(.dina(n1029),.dinb(n880),.dout(G252_fa_),.clk(gclk));
	jxor g0716(.dina(w_n827_0[1]),.dinb(w_n824_0[1]),.dout(n1031),.clk(gclk));
	jand g0717(.dina(w_dff_B_8loWY7PT9_0),.dinb(w_G252_0),.dout(n1032),.clk(gclk));
	jand g0718(.dina(n1032),.dinb(w_dff_B_VeT2Yyaa5_1),.dout(n1033),.clk(gclk));
	jor g0719(.dina(n1033),.dinb(w_dff_B_ZTSxbjnP1_1),.dout(n1034),.clk(gclk));
	jor g0720(.dina(w_n780_0[1]),.dinb(w_n776_0[1]),.dout(n1035),.clk(gclk));
	jand g0721(.dina(n1035),.dinb(w_n774_0[0]),.dout(n1036),.clk(gclk));
	jand g0722(.dina(w_dff_B_9GcvIL8U1_0),.dinb(n1034),.dout(n1037),.clk(gclk));
	jand g0723(.dina(n1037),.dinb(w_dff_B_NMFhvr9m9_1),.dout(n1038),.clk(gclk));
	jor g0724(.dina(n1038),.dinb(w_dff_B_u3oP7Dlo2_1),.dout(n1039),.clk(gclk));
	jxor g0725(.dina(w_n734_0[1]),.dinb(w_n373_3[0]),.dout(n1040),.clk(gclk));
	jxor g0726(.dina(w_n729_0[2]),.dinb(w_n726_0[2]),.dout(n1041),.clk(gclk));
	jand g0727(.dina(n1041),.dinb(w_n724_0[0]),.dout(n1042),.clk(gclk));
	jand g0728(.dina(w_n1042_0[1]),.dinb(w_n749_0[0]),.dout(n1043),.clk(gclk));
	jand g0729(.dina(n1043),.dinb(n1040),.dout(n1044),.clk(gclk));
	jand g0730(.dina(w_dff_B_T1d6BPOm2_0),.dinb(n1039),.dout(n1045),.clk(gclk));
	jor g0731(.dina(w_G2204_0[1]),.dinb(w_G1455_0[1]),.dout(n1046),.clk(gclk));
	jor g0732(.dina(n1046),.dinb(w_n367_0[0]),.dout(n1047),.clk(gclk));
	jand g0733(.dina(n1047),.dinb(w_G38_1[1]),.dout(n1048),.clk(gclk));
	jand g0734(.dina(w_n723_0[1]),.dinb(w_n720_0[1]),.dout(n1049),.clk(gclk));
	jand g0735(.dina(w_n741_1[0]),.dinb(w_n737_1[0]),.dout(n1050),.clk(gclk));
	jor g0736(.dina(w_n741_0[2]),.dinb(w_n737_0[2]),.dout(n1051),.clk(gclk));
	jand g0737(.dina(w_n747_0[1]),.dinb(w_n744_0[1]),.dout(n1052),.clk(gclk));
	jand g0738(.dina(n1052),.dinb(n1051),.dout(n1053),.clk(gclk));
	jor g0739(.dina(n1053),.dinb(n1050),.dout(n1054),.clk(gclk));
	jand g0740(.dina(n1054),.dinb(w_n1042_0[0]),.dout(n1055),.clk(gclk));
	jor g0741(.dina(n1055),.dinb(n1049),.dout(n1056),.clk(gclk));
	jor g0742(.dina(n1056),.dinb(n1048),.dout(n1057),.clk(gclk));
	jor g0743(.dina(w_dff_B_POG4d9VZ1_0),.dinb(n1045),.dout(n1058),.clk(gclk));
	jor g0744(.dina(n1058),.dinb(w_dff_B_B6UBMEla4_1),.dout(n1059),.clk(gclk));
	jand g0745(.dina(w_n1059_0[2]),.dinb(w_n718_0[2]),.dout(w_dff_A_WgdesOxS6_2),.clk(gclk));
	jnot g0746(.din(w_n644_0[0]),.dout(n1061),.clk(gclk));
	jnot g0747(.din(w_n655_0[0]),.dout(n1062),.clk(gclk));
	jnot g0748(.din(w_n656_0[0]),.dout(n1063),.clk(gclk));
	jand g0749(.dina(w_n641_0[1]),.dinb(w_G3705_1[0]),.dout(n1064),.clk(gclk));
	jor g0750(.dina(w_n641_0[0]),.dinb(w_G3705_0[2]),.dout(n1065),.clk(gclk));
	jand g0751(.dina(n1065),.dinb(w_n354_0[1]),.dout(n1066),.clk(gclk));
	jor g0752(.dina(n1066),.dinb(n1064),.dout(n1067),.clk(gclk));
	jor g0753(.dina(w_n1067_0[2]),.dinb(n1063),.dout(n1068),.clk(gclk));
	jand g0754(.dina(n1068),.dinb(n1062),.dout(n1069),.clk(gclk));
	jand g0755(.dina(w_n1069_0[2]),.dinb(n1061),.dout(n1070),.clk(gclk));
	jnot g0756(.din(w_n1070_0[1]),.dout(n1071),.clk(gclk));
	jor g0757(.dina(w_n669_0[0]),.dinb(w_G4526_2[0]),.dout(n1072),.clk(gclk));
	jand g0758(.dina(n1072),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0759(.dina(w_n1073_0[1]),.dinb(w_n654_0[1]),.dout(n1074),.clk(gclk));
	jand g0760(.dina(n1074),.dinb(w_n653_0[0]),.dout(n1075),.clk(gclk));
	jxor g0761(.dina(n1075),.dinb(w_n626_1[0]),.dout(w_dff_A_hPnAfq4F4_2),.clk(gclk));
	jxor g0762(.dina(w_n1073_0[0]),.dinb(w_n631_0[1]),.dout(w_dff_A_gTjHNFqz8_2),.clk(gclk));
	jand g0763(.dina(w_n359_0[2]),.dinb(w_G4526_1[2]),.dout(n1078),.clk(gclk));
	jor g0764(.dina(w_n666_0[0]),.dinb(w_n1078_0[1]),.dout(n1079),.clk(gclk));
	jand g0765(.dina(n1079),.dinb(w_n661_0[1]),.dout(n1080),.clk(gclk));
	jxor g0766(.dina(n1080),.dinb(w_n636_0[1]),.dout(w_dff_A_5B1bkyF47_2),.clk(gclk));
	jor g0767(.dina(w_n1078_0[0]),.dinb(w_n664_0[0]),.dout(n1082),.clk(gclk));
	jxor g0768(.dina(n1082),.dinb(w_n642_0[1]),.dout(w_dff_A_fpenTOu76_2),.clk(gclk));
	jxor g0769(.dina(w_n585_0[2]),.dinb(w_n582_0[0]),.dout(n1084),.clk(gclk));
	jor g0770(.dina(w_n1084_0[2]),.dinb(w_n678_0[0]),.dout(n1085),.clk(gclk));
	jnot g0771(.din(w_n646_0[0]),.dout(n1086),.clk(gclk));
	jnot g0772(.din(w_n647_0[0]),.dout(n1087),.clk(gclk));
	jnot g0773(.din(w_n654_0[0]),.dout(n1088),.clk(gclk));
	jand g0774(.dina(w_n1069_0[1]),.dinb(n1088),.dout(n1089),.clk(gclk));
	jor g0775(.dina(n1089),.dinb(w_n652_0[0]),.dout(n1090),.clk(gclk));
	jor g0776(.dina(w_n1090_0[1]),.dinb(w_n649_0[0]),.dout(n1091),.clk(gclk));
	jand g0777(.dina(n1091),.dinb(n1087),.dout(n1092),.clk(gclk));
	jand g0778(.dina(w_n1092_0[2]),.dinb(w_n1086_0[1]),.dout(n1093),.clk(gclk));
	jnot g0779(.din(w_G4526_1[1]),.dout(n1094),.clk(gclk));
	jand g0780(.dina(w_n1092_0[1]),.dinb(w_n1094_0[2]),.dout(n1095),.clk(gclk));
	jor g0781(.dina(n1095),.dinb(n1093),.dout(n1096),.clk(gclk));
	jand g0782(.dina(w_n1096_0[1]),.dinb(w_n618_0[0]),.dout(n1097),.clk(gclk));
	jor g0783(.dina(n1097),.dinb(w_n619_0[1]),.dout(n1098),.clk(gclk));
	jor g0784(.dina(n1098),.dinb(w_n588_0[0]),.dout(n1099),.clk(gclk));
	jor g0785(.dina(w_n1099_0[1]),.dinb(w_n586_0[1]),.dout(n1100),.clk(gclk));
	jand g0786(.dina(n1100),.dinb(w_dff_B_c1VlsQ6b8_1),.dout(w_dff_A_TNQcEwwd4_2),.clk(gclk));
	jand g0787(.dina(w_n676_0[1]),.dinb(w_n605_0[1]),.dout(n1102),.clk(gclk));
	jor g0788(.dina(n1102),.dinb(w_n615_0[1]),.dout(n1103),.clk(gclk));
	jxor g0789(.dina(n1103),.dinb(w_n594_0[1]),.dout(w_dff_A_RCtQWRw62_2),.clk(gclk));
	jnot g0790(.din(w_n599_0[0]),.dout(n1105),.clk(gclk));
	jnot g0791(.din(w_n613_0[1]),.dout(n1106),.clk(gclk));
	jnot g0792(.din(w_n603_0[2]),.dout(n1107),.clk(gclk));
	jand g0793(.dina(n1107),.dinb(w_G3729_0[2]),.dout(n1108),.clk(gclk));
	jor g0794(.dina(w_n1096_0[0]),.dinb(w_n1108_0[1]),.dout(n1109),.clk(gclk));
	jand g0795(.dina(n1109),.dinb(w_n1106_0[1]),.dout(n1110),.clk(gclk));
	jxor g0796(.dina(n1110),.dinb(w_n1105_0[1]),.dout(w_dff_A_OwLg3vyW3_2),.clk(gclk));
	jxor g0797(.dina(w_n676_0[0]),.dinb(w_n604_0[0]),.dout(w_dff_A_BjAxq4mU0_2),.clk(gclk));
	jnot g0798(.din(w_n436_0[0]),.dout(n1113),.clk(gclk));
	jor g0799(.dina(w_n1113_0[1]),.dinb(w_n431_0[0]),.dout(n1114),.clk(gclk));
	jnot g0800(.din(w_n432_0[0]),.dout(n1115),.clk(gclk));
	jor g0801(.dina(w_n435_0[0]),.dinb(n1115),.dout(n1116),.clk(gclk));
	jand g0802(.dina(n1116),.dinb(n1114),.dout(n1117),.clk(gclk));
	jnot g0803(.din(w_n459_0[0]),.dout(n1118),.clk(gclk));
	jxor g0804(.dina(w_n1118_0[1]),.dinb(w_n453_0[1]),.dout(n1119),.clk(gclk));
	jxor g0805(.dina(n1119),.dinb(n1117),.dout(n1120),.clk(gclk));
	jxor g0806(.dina(w_n485_0[0]),.dinb(w_n469_0[1]),.dout(n1121),.clk(gclk));
	jor g0807(.dina(w_n440_0[0]),.dinb(w_n422_0[0]),.dout(n1122),.clk(gclk));
	jnot g0808(.din(w_n423_0[0]),.dout(n1123),.clk(gclk));
	jor g0809(.dina(w_n427_0[0]),.dinb(n1123),.dout(n1124),.clk(gclk));
	jand g0810(.dina(n1124),.dinb(n1122),.dout(n1125),.clk(gclk));
	jnot g0811(.din(G141),.dout(n1126),.clk(gclk));
	jor g0812(.dina(n1126),.dinb(w_G18_20[0]),.dout(n1127),.clk(gclk));
	jnot g0813(.din(G161),.dout(n1128),.clk(gclk));
	jor g0814(.dina(n1128),.dinb(w_n355_15[0]),.dout(n1129),.clk(gclk));
	jand g0815(.dina(n1129),.dinb(w_n1127_0[1]),.dout(n1130),.clk(gclk));
	jxor g0816(.dina(n1130),.dinb(w_n479_0[2]),.dout(n1131),.clk(gclk));
	jxor g0817(.dina(n1131),.dinb(n1125),.dout(n1132),.clk(gclk));
	jxor g0818(.dina(n1132),.dinb(n1121),.dout(n1133),.clk(gclk));
	jxor g0819(.dina(n1133),.dinb(n1120),.dout(n1134),.clk(gclk));
	jxor g0820(.dina(w_n603_0[1]),.dinb(w_n598_0[2]),.dout(n1135),.clk(gclk));
	jand g0821(.dina(G239),.dinb(w_G18_19[2]),.dout(n1136),.clk(gclk));
	jand g0822(.dina(G44),.dinb(w_n355_14[2]),.dout(n1137),.clk(gclk));
	jor g0823(.dina(w_n1137_0[1]),.dinb(n1136),.dout(n1138),.clk(gclk));
	jxor g0824(.dina(n1138),.dinb(w_n651_0[0]),.dout(n1139),.clk(gclk));
	jxor g0825(.dina(n1139),.dinb(n1135),.dout(n1140),.clk(gclk));
	jand g0826(.dina(G229),.dinb(w_G18_19[1]),.dout(n1141),.clk(gclk));
	jor g0827(.dina(n1141),.dinb(w_n663_0[2]),.dout(n1142),.clk(gclk));
	jxor g0828(.dina(n1142),.dinb(w_n660_0[0]),.dout(n1143),.clk(gclk));
	jxor g0829(.dina(w_n635_0[1]),.dinb(w_n625_0[1]),.dout(n1144),.clk(gclk));
	jxor g0830(.dina(n1144),.dinb(n1143),.dout(n1145),.clk(gclk));
	jxor g0831(.dina(w_n593_0[1]),.dinb(w_n585_0[1]),.dout(n1146),.clk(gclk));
	jxor g0832(.dina(n1146),.dinb(n1145),.dout(n1147),.clk(gclk));
	jxor g0833(.dina(n1147),.dinb(n1140),.dout(n1148),.clk(gclk));
	jor g0834(.dina(n1148),.dinb(n1134),.dout(n1149),.clk(gclk));
	jor g0835(.dina(w_n372_0[0]),.dinb(w_n355_14[1]),.dout(n1150),.clk(gclk));
	jxor g0836(.dina(G212),.dinb(G211),.dout(n1151),.clk(gclk));
	jxor g0837(.dina(n1151),.dinb(w_G209_0[0]),.dout(n1152),.clk(gclk));
	jor g0838(.dina(n1152),.dinb(w_n1150_0[1]),.dout(n1153),.clk(gclk));
	jnot g0839(.din(w_n386_0[0]),.dout(n1154),.clk(gclk));
	jand g0840(.dina(w_n395_0[2]),.dinb(n1154),.dout(n1155),.clk(gclk));
	jnot g0841(.din(w_n394_0[0]),.dout(n1156),.clk(gclk));
	jand g0842(.dina(n1156),.dinb(w_n387_0[1]),.dout(n1157),.clk(gclk));
	jor g0843(.dina(n1157),.dinb(n1155),.dout(n1158),.clk(gclk));
	jor g0844(.dina(w_n380_0[0]),.dinb(w_n374_0[0]),.dout(n1159),.clk(gclk));
	jnot g0845(.din(w_n375_0[0]),.dout(n1160),.clk(gclk));
	jor g0846(.dina(w_n378_0[0]),.dinb(n1160),.dout(n1161),.clk(gclk));
	jand g0847(.dina(n1161),.dinb(n1159),.dout(n1162),.clk(gclk));
	jxor g0848(.dina(n1162),.dinb(n1158),.dout(n1163),.clk(gclk));
	jxor g0849(.dina(n1163),.dinb(n1153),.dout(n1164),.clk(gclk));
	jxor g0850(.dina(w_n689_0[0]),.dinb(w_n504_0[2]),.dout(n1165),.clk(gclk));
	jxor g0851(.dina(w_n523_0[0]),.dinb(w_n517_0[2]),.dout(n1166),.clk(gclk));
	jxor g0852(.dina(n1166),.dinb(n1165),.dout(n1167),.clk(gclk));
	jxor g0853(.dina(w_n555_0[1]),.dinb(w_n539_0[1]),.dout(n1168),.clk(gclk));
	jxor g0854(.dina(w_n547_0[1]),.dinb(w_n531_0[1]),.dout(n1169),.clk(gclk));
	jxor g0855(.dina(n1169),.dinb(n1168),.dout(n1170),.clk(gclk));
	jand g0856(.dina(G227),.dinb(w_G18_19[0]),.dout(n1171),.clk(gclk));
	jand g0857(.dina(G115),.dinb(w_n355_14[0]),.dout(n1172),.clk(gclk));
	jor g0858(.dina(w_n1172_0[1]),.dinb(n1171),.dout(n1173),.clk(gclk));
	jxor g0859(.dina(n1173),.dinb(w_n563_0[2]),.dout(n1174),.clk(gclk));
	jxor g0860(.dina(n1174),.dinb(n1170),.dout(n1175),.clk(gclk));
	jxor g0861(.dina(n1175),.dinb(n1167),.dout(n1176),.clk(gclk));
	jor g0862(.dina(n1176),.dinb(n1164),.dout(n1177),.clk(gclk));
	jor g0863(.dina(n1177),.dinb(n1149),.dout(G412_fa_),.clk(gclk));
	jnot g0864(.din(w_n772_0[0]),.dout(n1179),.clk(gclk));
	jxor g0865(.dina(w_n780_0[0]),.dinb(n1179),.dout(n1180),.clk(gclk));
	jnot g0866(.din(w_G2208_0[1]),.dout(n1181),.clk(gclk));
	jor g0867(.dina(n1181),.dinb(w_n355_13[2]),.dout(n1182),.clk(gclk));
	jor g0868(.dina(G82),.dinb(w_G18_18[2]),.dout(n1183),.clk(gclk));
	jand g0869(.dina(n1183),.dinb(n1182),.dout(n1184),.clk(gclk));
	jxor g0870(.dina(n1184),.dinb(w_n827_0[0]),.dout(n1185),.clk(gclk));
	jxor g0871(.dina(n1185),.dinb(n1180),.dout(n1186),.clk(gclk));
	jxor g0872(.dina(w_n806_0[0]),.dinb(w_n800_0[1]),.dout(n1187),.clk(gclk));
	jxor g0873(.dina(w_n820_0[0]),.dinb(w_n814_0[1]),.dout(n1188),.clk(gclk));
	jxor g0874(.dina(n1188),.dinb(n1187),.dout(n1189),.clk(gclk));
	jxor g0875(.dina(w_n764_0[0]),.dinb(w_n758_0[1]),.dout(n1190),.clk(gclk));
	jxor g0876(.dina(n1190),.dinb(n1189),.dout(n1191),.clk(gclk));
	jxor g0877(.dina(n1191),.dinb(n1186),.dout(n1192),.clk(gclk));
	jxor g0878(.dina(w_n953_0[1]),.dinb(w_n947_0[0]),.dout(n1193),.clk(gclk));
	jxor g0879(.dina(w_n903_0[0]),.dinb(w_n894_0[0]),.dout(n1194),.clk(gclk));
	jxor g0880(.dina(n1194),.dinb(n1193),.dout(n1195),.clk(gclk));
	jnot g0881(.din(w_G3698_0[1]),.dout(n1196),.clk(gclk));
	jor g0882(.dina(n1196),.dinb(w_n355_13[1]),.dout(n1197),.clk(gclk));
	jor g0883(.dina(G69),.dinb(w_G18_18[1]),.dout(n1198),.clk(gclk));
	jand g0884(.dina(n1198),.dinb(n1197),.dout(n1199),.clk(gclk));
	jxor g0885(.dina(n1199),.dinb(w_n888_0[0]),.dout(n1200),.clk(gclk));
	jor g0886(.dina(w_n662_0[0]),.dinb(w_n355_13[0]),.dout(n1201),.clk(gclk));
	jand g0887(.dina(n1201),.dinb(w_n905_0[0]),.dout(n1202),.clk(gclk));
	jxor g0888(.dina(n1202),.dinb(w_n919_0[0]),.dout(n1203),.clk(gclk));
	jxor g0889(.dina(n1203),.dinb(n1200),.dout(n1204),.clk(gclk));
	jnot g0890(.din(w_n930_0[0]),.dout(n1205),.clk(gclk));
	jxor g0891(.dina(w_n938_0[0]),.dinb(n1205),.dout(n1206),.clk(gclk));
	jxor g0892(.dina(n1206),.dinb(n1204),.dout(n1207),.clk(gclk));
	jxor g0893(.dina(n1207),.dinb(n1195),.dout(n1208),.clk(gclk));
	jor g0894(.dina(n1208),.dinb(n1192),.dout(n1209),.clk(gclk));
	jxor g0895(.dina(w_n854_0[0]),.dinb(w_n848_0[1]),.dout(n1210),.clk(gclk));
	jxor g0896(.dina(w_n870_0[0]),.dinb(w_n862_0[0]),.dout(n1211),.clk(gclk));
	jxor g0897(.dina(n1211),.dinb(n1210),.dout(n1212),.clk(gclk));
	jxor g0898(.dina(w_n983_0[0]),.dinb(w_n977_0[1]),.dout(n1213),.clk(gclk));
	jand g0899(.dina(w_G4393_0[1]),.dinb(w_G18_18[0]),.dout(n1214),.clk(gclk));
	jnot g0900(.din(G58),.dout(n1215),.clk(gclk));
	jand g0901(.dina(n1215),.dinb(w_n355_12[2]),.dout(n1216),.clk(gclk));
	jor g0902(.dina(n1216),.dinb(n1214),.dout(n1217),.clk(gclk));
	jxor g0903(.dina(n1217),.dinb(w_n970_0[0]),.dout(n1218),.clk(gclk));
	jxor g0904(.dina(w_n999_0[0]),.dinb(w_n991_0[0]),.dout(n1219),.clk(gclk));
	jxor g0905(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jxor g0906(.dina(n1220),.dinb(n1213),.dout(n1221),.clk(gclk));
	jxor g0907(.dina(n1221),.dinb(n1212),.dout(n1222),.clk(gclk));
	jxor g0908(.dina(w_n366_0[0]),.dinb(w_G1492_1[0]),.dout(n1223),.clk(gclk));
	jor g0909(.dina(n1223),.dinb(w_n355_12[1]),.dout(n1224),.clk(gclk));
	jnot g0910(.din(w_G1455_0[0]),.dout(n1225),.clk(gclk));
	jxor g0911(.dina(w_G2204_0[0]),.dinb(n1225),.dout(n1226),.clk(gclk));
	jor g0912(.dina(n1226),.dinb(w_G18_17[2]),.dout(n1227),.clk(gclk));
	jand g0913(.dina(n1227),.dinb(n1224),.dout(n1228),.clk(gclk));
	jxor g0914(.dina(w_n729_0[1]),.dinb(w_n723_0[0]),.dout(n1229),.clk(gclk));
	jxor g0915(.dina(w_n747_0[0]),.dinb(w_n741_0[1]),.dout(n1230),.clk(gclk));
	jxor g0916(.dina(n1230),.dinb(n1229),.dout(n1231),.clk(gclk));
	jnot g0917(.din(w_G1459_0[1]),.dout(n1232),.clk(gclk));
	jor g0918(.dina(n1232),.dinb(w_n355_12[0]),.dout(n1233),.clk(gclk));
	jor g0919(.dina(G114),.dinb(w_G18_17[1]),.dout(n1234),.clk(gclk));
	jand g0920(.dina(n1234),.dinb(n1233),.dout(n1235),.clk(gclk));
	jxor g0921(.dina(n1235),.dinb(w_n734_0[0]),.dout(n1236),.clk(gclk));
	jxor g0922(.dina(n1236),.dinb(n1231),.dout(n1237),.clk(gclk));
	jxor g0923(.dina(n1237),.dinb(n1228),.dout(n1238),.clk(gclk));
	jor g0924(.dina(n1238),.dinb(n1222),.dout(n1239),.clk(gclk));
	jor g0925(.dina(n1239),.dinb(n1209),.dout(G414_fa_),.clk(gclk));
	jnot g0926(.din(w_n935_0[0]),.dout(n1241),.clk(gclk));
	jxor g0927(.dina(n1241),.dinb(w_n926_0[0]),.dout(n1242),.clk(gclk));
	jxor g0928(.dina(w_n950_0[1]),.dinb(w_n944_0[0]),.dout(n1243),.clk(gclk));
	jxor g0929(.dina(n1243),.dinb(n1242),.dout(n1244),.clk(gclk));
	jand g0930(.dina(G208),.dinb(w_G18_17[0]),.dout(n1245),.clk(gclk));
	jor g0931(.dina(n1245),.dinb(w_n1137_0[0]),.dout(n1246),.clk(gclk));
	jand g0932(.dina(G198),.dinb(w_G18_16[2]),.dout(n1247),.clk(gclk));
	jor g0933(.dina(n1247),.dinb(w_n663_0[1]),.dout(n1248),.clk(gclk));
	jxor g0934(.dina(n1248),.dinb(n1246),.dout(n1249),.clk(gclk));
	jxor g0935(.dina(w_n916_0[0]),.dinb(w_n885_0[0]),.dout(n1250),.clk(gclk));
	jxor g0936(.dina(n1250),.dinb(n1249),.dout(n1251),.clk(gclk));
	jxor g0937(.dina(w_n900_0[0]),.dinb(w_n891_0[0]),.dout(n1252),.clk(gclk));
	jxor g0938(.dina(n1252),.dinb(n1251),.dout(n1253),.clk(gclk));
	jxor g0939(.dina(n1253),.dinb(n1244),.dout(n1254),.clk(gclk));
	jxor g0940(.dina(w_n866_0[0]),.dinb(w_n858_0[0]),.dout(n1255),.clk(gclk));
	jxor g0941(.dina(w_n995_0[0]),.dinb(w_n987_0[0]),.dout(n1256),.clk(gclk));
	jxor g0942(.dina(n1256),.dinb(n1255),.dout(n1257),.clk(gclk));
	jxor g0943(.dina(w_n980_0[0]),.dinb(w_n973_0[1]),.dout(n1258),.clk(gclk));
	jand g0944(.dina(G197),.dinb(w_G18_16[1]),.dout(n1259),.clk(gclk));
	jor g0945(.dina(n1259),.dinb(w_n1172_0[0]),.dout(n1260),.clk(gclk));
	jxor g0946(.dina(n1260),.dinb(w_n966_0[0]),.dout(n1261),.clk(gclk));
	jxor g0947(.dina(n1261),.dinb(n1258),.dout(n1262),.clk(gclk));
	jnot g0948(.din(w_n851_0[0]),.dout(n1263),.clk(gclk));
	jxor g0949(.dina(n1263),.dinb(w_n845_0[1]),.dout(n1264),.clk(gclk));
	jxor g0950(.dina(n1264),.dinb(n1262),.dout(n1265),.clk(gclk));
	jxor g0951(.dina(n1265),.dinb(n1257),.dout(n1266),.clk(gclk));
	jor g0952(.dina(n1266),.dinb(n1254),.dout(n1267),.clk(gclk));
	jxor g0953(.dina(G165),.dinb(G164),.dout(n1268),.clk(gclk));
	jxor g0954(.dina(n1268),.dinb(G170),.dout(n1269),.clk(gclk));
	jor g0955(.dina(n1269),.dinb(w_n1150_0[0]),.dout(n1270),.clk(gclk));
	jnot g0956(.din(w_n736_0[0]),.dout(n1271),.clk(gclk));
	jand g0957(.dina(w_n744_0[0]),.dinb(n1271),.dout(n1272),.clk(gclk));
	jnot g0958(.din(w_n743_0[0]),.dout(n1273),.clk(gclk));
	jand g0959(.dina(n1273),.dinb(w_n737_0[1]),.dout(n1274),.clk(gclk));
	jor g0960(.dina(n1274),.dinb(n1272),.dout(n1275),.clk(gclk));
	jnot g0961(.din(w_n726_0[1]),.dout(n1276),.clk(gclk));
	jor g0962(.dina(n1276),.dinb(w_n719_0[0]),.dout(n1277),.clk(gclk));
	jnot g0963(.din(w_n720_0[0]),.dout(n1278),.clk(gclk));
	jor g0964(.dina(w_n725_0[0]),.dinb(n1278),.dout(n1279),.clk(gclk));
	jand g0965(.dina(n1279),.dinb(n1277),.dout(n1280),.clk(gclk));
	jxor g0966(.dina(n1280),.dinb(n1275),.dout(n1281),.clk(gclk));
	jxor g0967(.dina(n1281),.dinb(n1270),.dout(n1282),.clk(gclk));
	jor g0968(.dina(n1282),.dinb(n1267),.dout(n1283),.clk(gclk));
	jnot g0969(.din(G181),.dout(n1284),.clk(gclk));
	jor g0970(.dina(n1284),.dinb(w_n355_11[2]),.dout(n1285),.clk(gclk));
	jand g0971(.dina(n1285),.dinb(w_n1127_0[0]),.dout(n1286),.clk(gclk));
	jxor g0972(.dina(n1286),.dinb(w_n824_0[0]),.dout(n1287),.clk(gclk));
	jxor g0973(.dina(w_n803_0[0]),.dinb(w_n796_0[1]),.dout(n1288),.clk(gclk));
	jxor g0974(.dina(n1288),.dinb(n1287),.dout(n1289),.clk(gclk));
	jnot g0975(.din(w_n767_0[0]),.dout(n1290),.clk(gclk));
	jand g0976(.dina(w_n776_0[0]),.dinb(n1290),.dout(n1291),.clk(gclk));
	jnot g0977(.din(w_n775_0[0]),.dout(n1292),.clk(gclk));
	jand g0978(.dina(n1292),.dinb(w_n768_0[0]),.dout(n1293),.clk(gclk));
	jor g0979(.dina(n1293),.dinb(n1291),.dout(n1294),.clk(gclk));
	jnot g0980(.din(w_n754_0[0]),.dout(n1295),.clk(gclk));
	jand g0981(.dina(w_n761_0[0]),.dinb(n1295),.dout(n1296),.clk(gclk));
	jnot g0982(.din(w_n760_0[0]),.dout(n1297),.clk(gclk));
	jand g0983(.dina(n1297),.dinb(w_n755_0[1]),.dout(n1298),.clk(gclk));
	jor g0984(.dina(n1298),.dinb(n1296),.dout(n1299),.clk(gclk));
	jxor g0985(.dina(n1299),.dinb(n1294),.dout(n1300),.clk(gclk));
	jxor g0986(.dina(w_n817_0[0]),.dinb(w_n810_0[1]),.dout(n1301),.clk(gclk));
	jxor g0987(.dina(n1301),.dinb(n1300),.dout(n1302),.clk(gclk));
	jxor g0988(.dina(n1302),.dinb(n1289),.dout(n1303),.clk(gclk));
	jor g0989(.dina(n1303),.dinb(n1283),.dout(G416_fa_),.clk(gclk));
	jnot g0990(.din(w_n480_1[0]),.dout(n1305),.clk(gclk));
	jnot g0991(.din(w_n505_0[0]),.dout(n1306),.clk(gclk));
	jnot g0992(.din(w_n513_1[0]),.dout(n1307),.clk(gclk));
	jnot g0993(.din(w_n524_1[0]),.dout(n1308),.clk(gclk));
	jnot g0994(.din(w_n572_1[0]),.dout(n1309),.clk(gclk));
	jnot g0995(.din(w_n581_0[1]),.dout(n1310),.clk(gclk));
	jnot g0996(.din(w_n586_0[0]),.dout(n1311),.clk(gclk));
	jand g0997(.dina(w_n1099_0[0]),.dinb(n1311),.dout(n1312),.clk(gclk));
	jor g0998(.dina(w_n1312_1[1]),.dinb(w_n1310_0[1]),.dout(n1313),.clk(gclk));
	jand g0999(.dina(n1313),.dinb(w_n1309_0[1]),.dout(n1314),.clk(gclk));
	jor g1000(.dina(n1314),.dinb(w_n526_0[1]),.dout(n1315),.clk(gclk));
	jor g1001(.dina(n1315),.dinb(w_n1308_0[1]),.dout(n1316),.clk(gclk));
	jor g1002(.dina(w_n1316_0[1]),.dinb(w_n518_1[0]),.dout(n1317),.clk(gclk));
	jor g1003(.dina(w_n1317_0[1]),.dinb(w_n1307_0[1]),.dout(n1318),.clk(gclk));
	jand g1004(.dina(w_n696_0[0]),.dinb(n1318),.dout(n1319),.clk(gclk));
	jor g1005(.dina(n1319),.dinb(w_n507_0[0]),.dout(n1320),.clk(gclk));
	jand g1006(.dina(n1320),.dinb(n1306),.dout(n1321),.clk(gclk));
	jxor g1007(.dina(w_n1321_1[1]),.dinb(w_dff_B_MmUI7ZMm7_1),.dout(w_dff_A_ZJcOyy2e3_2),.clk(gclk));
	jnot g1008(.din(w_n414_1[0]),.dout(n1323),.clk(gclk));
	jnot g1009(.din(w_n424_0[0]),.dout(n1324),.clk(gclk));
	jnot g1010(.din(w_n425_1[0]),.dout(n1325),.clk(gclk));
	jnot g1011(.din(w_n450_0[1]),.dout(n1326),.clk(gclk));
	jnot g1012(.din(w_n449_0[2]),.dout(n1327),.clk(gclk));
	jnot g1013(.din(w_n499_0[0]),.dout(n1328),.clk(gclk));
	jnot g1014(.din(w_n500_0[0]),.dout(n1329),.clk(gclk));
	jnot g1015(.din(w_n462_0[0]),.dout(n1330),.clk(gclk));
	jand g1016(.dina(w_n1321_1[0]),.dinb(n1330),.dout(n1331),.clk(gclk));
	jand g1017(.dina(n1331),.dinb(n1329),.dout(n1332),.clk(gclk));
	jor g1018(.dina(n1332),.dinb(n1328),.dout(n1333),.clk(gclk));
	jand g1019(.dina(w_n1333_0[1]),.dinb(n1327),.dout(n1334),.clk(gclk));
	jor g1020(.dina(n1334),.dinb(n1326),.dout(n1335),.clk(gclk));
	jor g1021(.dina(n1335),.dinb(n1325),.dout(n1336),.clk(gclk));
	jand g1022(.dina(n1336),.dinb(n1324),.dout(n1337),.clk(gclk));
	jxor g1023(.dina(w_n1337_1[1]),.dinb(w_n1323_0[1]),.dout(w_dff_A_fhIVqjCk4_2),.clk(gclk));
	jand g1024(.dina(w_n1118_0[0]),.dinb(w_G2230_0[1]),.dout(n1339),.clk(gclk));
	jnot g1025(.din(n1339),.dout(n1340),.clk(gclk));
	jand g1026(.dina(w_n1321_0[2]),.dinb(w_n495_1[0]),.dout(n1341),.clk(gclk));
	jnot g1027(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1028(.dina(n1342),.dinb(w_n497_1[0]),.dout(n1343),.clk(gclk));
	jand g1029(.dina(w_n1343_0[1]),.dinb(w_n1340_0[2]),.dout(n1344),.clk(gclk));
	jor g1030(.dina(w_n1344_0[1]),.dinb(w_n460_1[1]),.dout(n1345),.clk(gclk));
	jxor g1031(.dina(n1345),.dinb(w_n463_1[0]),.dout(w_dff_A_GCOhVMYb7_2),.clk(gclk));
	jor g1032(.dina(w_n1343_0[0]),.dinb(w_n464_0[1]),.dout(n1347),.clk(gclk));
	jnot g1033(.din(w_n1344_0[0]),.dout(n1348),.clk(gclk));
	jor g1034(.dina(n1348),.dinb(w_n460_1[0]),.dout(n1349),.clk(gclk));
	jand g1035(.dina(n1349),.dinb(w_dff_B_WDf4wCSn8_1),.dout(w_dff_A_bWmbwUsV7_2),.clk(gclk));
	jnot g1036(.din(w_n489_0[1]),.dout(n1351),.clk(gclk));
	jor g1037(.dina(n1351),.dinb(w_n491_1[0]),.dout(n1352),.clk(gclk));
	jand g1038(.dina(w_n700_1[0]),.dinb(w_n481_0[0]),.dout(n1353),.clk(gclk));
	jor g1039(.dina(n1353),.dinb(n1352),.dout(n1354),.clk(gclk));
	jxor g1040(.dina(n1354),.dinb(w_n470_0[1]),.dout(w_dff_A_Zs4DPBih4_2),.clk(gclk));
	jand g1041(.dina(w_n700_0[2]),.dinb(w_n480_0[2]),.dout(n1356),.clk(gclk));
	jor g1042(.dina(n1356),.dinb(w_n487_0[1]),.dout(n1357),.clk(gclk));
	jxor g1043(.dina(n1357),.dinb(w_n475_0[1]),.dout(w_dff_A_A2Ayl1W59_2),.clk(gclk));
	jor g1044(.dina(w_n418_0[0]),.dinb(w_n411_1[0]),.dout(n1359),.clk(gclk));
	jor g1045(.dina(w_n707_1[1]),.dinb(w_n411_0[2]),.dout(n1360),.clk(gclk));
	jand g1046(.dina(n1360),.dinb(w_n1359_0[1]),.dout(n1361),.clk(gclk));
	jxor g1047(.dina(n1361),.dinb(w_n377_1[0]),.dout(w_dff_A_Di2h08h34_2),.clk(gclk));
	jand g1048(.dina(w_n415_0[0]),.dinb(w_n388_1[0]),.dout(n1363),.clk(gclk));
	jor g1049(.dina(n1363),.dinb(w_n409_1[0]),.dout(n1364),.clk(gclk));
	jor g1050(.dina(w_n707_1[0]),.dinb(w_n409_0[2]),.dout(n1365),.clk(gclk));
	jand g1051(.dina(n1365),.dinb(w_n1364_0[1]),.dout(n1366),.clk(gclk));
	jxor g1052(.dina(n1366),.dinb(w_n416_0[1]),.dout(w_dff_A_mrhQvpES1_2),.clk(gclk));
	jnot g1053(.din(w_n388_0[2]),.dout(n1368),.clk(gclk));
	jnot g1054(.din(w_n396_1[0]),.dout(n1369),.clk(gclk));
	jnot g1055(.din(w_n392_0[1]),.dout(n1370),.clk(gclk));
	jor g1056(.dina(w_n1337_1[0]),.dinb(w_n1323_0[0]),.dout(n1371),.clk(gclk));
	jand g1057(.dina(n1371),.dinb(w_n1370_0[1]),.dout(n1372),.clk(gclk));
	jor g1058(.dina(w_n1372_0[1]),.dinb(w_n1369_0[1]),.dout(n1373),.clk(gclk));
	jand g1059(.dina(n1373),.dinb(w_n405_0[1]),.dout(n1374),.clk(gclk));
	jxor g1060(.dina(n1374),.dinb(w_dff_B_IOPm2ZGa5_1),.dout(G333),.clk(gclk));
	jxor g1061(.dina(w_n1372_0[0]),.dinb(w_n1369_0[0]),.dout(w_dff_A_iQ4quPVT4_2),.clk(gclk));
	jor g1062(.dina(w_G416_0),.dinb(w_G414_0),.dout(n1377),.clk(gclk));
	jor g1063(.dina(w_G408_0),.dinb(w_G404_0),.dout(n1378),.clk(gclk));
	jor g1064(.dina(w_G410_0),.dinb(w_G406_0),.dout(n1379),.clk(gclk));
	jor g1065(.dina(w_dff_B_RIw1Ilxk0_0),.dinb(w_G412_0),.dout(n1380),.clk(gclk));
	jor g1066(.dina(n1380),.dinb(w_dff_B_avQhiC6t0_1),.dout(n1381),.clk(gclk));
	jor g1067(.dina(n1381),.dinb(w_dff_B_39kMFezJ5_1),.dout(w_dff_A_bYZjOR4l8_2),.clk(gclk));
	jxor g1068(.dina(w_n705_0[0]),.dinb(w_n425_0[2]),.dout(w_dff_A_xYcOwCKE4_2),.clk(gclk));
	jand g1069(.dina(w_n703_1[1]),.dinb(w_n438_0[0]),.dout(n1384),.clk(gclk));
	jor g1070(.dina(n1384),.dinb(w_n447_0[1]),.dout(n1385),.clk(gclk));
	jxor g1071(.dina(n1385),.dinb(w_n429_0[1]),.dout(w_dff_A_DKHFtTxw2_2),.clk(gclk));
	jand g1072(.dina(w_n1113_0[0]),.dinb(w_G2239_0[2]),.dout(n1387),.clk(gclk));
	jnot g1073(.din(w_n1387_0[1]),.dout(n1388),.clk(gclk));
	jor g1074(.dina(w_n703_1[0]),.dinb(w_n445_0[1]),.dout(n1389),.clk(gclk));
	jand g1075(.dina(n1389),.dinb(w_n1388_0[1]),.dout(n1390),.clk(gclk));
	jxor g1076(.dina(n1390),.dinb(w_n433_1[0]),.dout(w_dff_A_xHBLP3f76_2),.clk(gclk));
	jxor g1077(.dina(w_n703_0[2]),.dinb(w_n437_0[1]),.dout(w_dff_A_kmbXyAx51_2),.clk(gclk));
	jxor g1078(.dina(w_n680_2[1]),.dinb(w_n575_1[0]),.dout(w_dff_A_g9igXi8t2_2),.clk(gclk));
	jor g1079(.dina(w_n712_0[1]),.dinb(w_G38_1[0]),.dout(n1394),.clk(gclk));
	jor g1080(.dina(w_n713_0[0]),.dinb(w_n709_1[0]),.dout(n1395),.clk(gclk));
	jand g1081(.dina(n1395),.dinb(n1394),.dout(n1396),.clk(gclk));
	jxor g1082(.dina(w_n1396_0[1]),.dinb(w_n370_0[1]),.dout(G422),.clk(gclk));
	jxor g1083(.dina(w_n709_0[2]),.dinb(w_n363_0[1]),.dout(w_dff_A_DGJTufCb5_2),.clk(gclk));
	jand g1084(.dina(w_n680_2[0]),.dinb(w_n580_0[1]),.dout(n1399),.clk(gclk));
	jor g1085(.dina(n1399),.dinb(w_n570_1[1]),.dout(n1400),.clk(gclk));
	jxor g1086(.dina(n1400),.dinb(w_n573_1[0]),.dout(w_dff_A_Snttc1Yu1_2),.clk(gclk));
	jnot g1087(.din(w_n577_0[0]),.dout(n1402),.clk(gclk));
	jnot g1088(.din(w_n548_0[0]),.dout(n1403),.clk(gclk));
	jnot g1089(.din(w_n566_0[1]),.dout(n1404),.clk(gclk));
	jnot g1090(.din(w_n576_0[1]),.dout(n1405),.clk(gclk));
	jand g1091(.dina(n1405),.dinb(n1404),.dout(n1406),.clk(gclk));
	jor g1092(.dina(n1406),.dinb(w_n550_0[0]),.dout(n1407),.clk(gclk));
	jand g1093(.dina(n1407),.dinb(n1403),.dout(n1408),.clk(gclk));
	jnot g1094(.din(w_n568_0[1]),.dout(n1409),.clk(gclk));
	jand g1095(.dina(w_n1312_1[0]),.dinb(n1409),.dout(n1410),.clk(gclk));
	jor g1096(.dina(n1410),.dinb(w_n1408_0[1]),.dout(n1411),.clk(gclk));
	jxor g1097(.dina(n1411),.dinb(w_n1402_0[1]),.dout(w_dff_A_T4PMdRc97_2),.clk(gclk));
	jand g1098(.dina(w_n680_1[2]),.dinb(w_n576_0[0]),.dout(n1413),.clk(gclk));
	jor g1099(.dina(n1413),.dinb(w_n566_0[0]),.dout(n1414),.clk(gclk));
	jxor g1100(.dina(n1414),.dinb(w_n578_0[1]),.dout(w_dff_A_B7P868BX1_2),.clk(gclk));
	jand g1101(.dina(w_n680_1[1]),.dinb(w_n575_0[2]),.dout(n1416),.clk(gclk));
	jor g1102(.dina(n1416),.dinb(w_n564_0[1]),.dout(n1417),.clk(gclk));
	jxor g1103(.dina(n1417),.dinb(w_n574_0[1]),.dout(w_dff_A_eHl8FGiB3_2),.clk(gclk));
	jxor g1104(.dina(w_n504_0[1]),.dinb(w_n501_0[0]),.dout(n1419),.clk(gclk));
	jxor g1105(.dina(w_n1419_0[1]),.dinb(w_n698_0[0]),.dout(w_dff_A_5mhHFufl9_2),.clk(gclk));
	jand g1106(.dina(w_n694_0[0]),.dinb(w_n1317_0[0]),.dout(n1421),.clk(gclk));
	jxor g1107(.dina(n1421),.dinb(w_n1307_0[0]),.dout(w_dff_A_xY7oVWid9_2),.clk(gclk));
	jxor g1108(.dina(w_n524_0[2]),.dinb(w_n518_0[2]),.dout(n1423),.clk(gclk));
	jor g1109(.dina(n1423),.dinb(w_n683_0[0]),.dout(n1424),.clk(gclk));
	jand g1110(.dina(n1424),.dinb(w_n1316_0[0]),.dout(w_dff_A_fHXgdtt22_2),.clk(gclk));
	jxor g1111(.dina(w_n517_0[1]),.dinb(w_n514_0[0]),.dout(n1426),.clk(gclk));
	jxor g1112(.dina(w_n1426_0[1]),.dinb(w_n682_0[0]),.dout(w_dff_A_DuDkDjYi5_2),.clk(gclk));
	jxor g1113(.dina(w_n429_0[0]),.dinb(w_n425_0[1]),.dout(n1431),.clk(gclk));
	jor g1114(.dina(w_n1388_0[0]),.dinb(w_n444_0[1]),.dout(n1432),.clk(gclk));
	jnot g1115(.din(w_n447_0[0]),.dout(n1433),.clk(gclk));
	jor g1116(.dina(w_n1433_0[1]),.dinb(w_n1387_0[0]),.dout(n1434),.clk(gclk));
	jand g1117(.dina(n1434),.dinb(n1432),.dout(n1435),.clk(gclk));
	jxor g1118(.dina(n1435),.dinb(w_n1431_0[1]),.dout(n1436),.clk(gclk));
	jxor g1119(.dina(w_n449_0[1]),.dinb(w_n433_0[2]),.dout(n1437),.clk(gclk));
	jxor g1120(.dina(n1437),.dinb(n1436),.dout(n1438),.clk(gclk));
	jand g1121(.dina(n1438),.dinb(w_n1333_0[0]),.dout(n1439),.clk(gclk));
	jxor g1122(.dina(w_n445_0[0]),.dinb(w_n433_0[1]),.dout(n1440),.clk(gclk));
	jnot g1123(.din(w_n1440_0[1]),.dout(n1441),.clk(gclk));
	jand g1124(.dina(n1441),.dinb(w_n1433_0[0]),.dout(n1442),.clk(gclk));
	jor g1125(.dina(w_n437_0[0]),.dinb(w_n444_0[0]),.dout(n1443),.clk(gclk));
	jand g1126(.dina(n1443),.dinb(w_n1440_0[0]),.dout(n1444),.clk(gclk));
	jor g1127(.dina(n1444),.dinb(n1442),.dout(n1445),.clk(gclk));
	jxor g1128(.dina(w_n1431_0[0]),.dinb(w_n450_0[0]),.dout(n1446),.clk(gclk));
	jxor g1129(.dina(n1446),.dinb(n1445),.dout(n1447),.clk(gclk));
	jand g1130(.dina(n1447),.dinb(w_n703_0[1]),.dout(n1448),.clk(gclk));
	jor g1131(.dina(n1448),.dinb(n1439),.dout(n1449),.clk(gclk));
	jand g1132(.dina(w_n497_0[2]),.dinb(w_n1340_0[1]),.dout(n1450),.clk(gclk));
	jor g1133(.dina(n1450),.dinb(w_n460_0[2]),.dout(n1451),.clk(gclk));
	jxor g1134(.dina(w_n480_0[1]),.dinb(w_n475_0[0]),.dout(n1452),.clk(gclk));
	jand g1135(.dina(w_n1452_0[2]),.dinb(w_n495_0[2]),.dout(n1453),.clk(gclk));
	jnot g1136(.din(w_n1452_0[1]),.dout(n1454),.clk(gclk));
	jand g1137(.dina(n1454),.dinb(w_n497_0[1]),.dout(n1455),.clk(gclk));
	jor g1138(.dina(n1455),.dinb(n1453),.dout(n1456),.clk(gclk));
	jnot g1139(.din(w_n479_0[1]),.dout(n1457),.clk(gclk));
	jand g1140(.dina(n1457),.dinb(w_G2211_0[1]),.dout(n1458),.clk(gclk));
	jnot g1141(.din(w_n1458_0[1]),.dout(n1459),.clk(gclk));
	jor g1142(.dina(n1459),.dinb(w_n491_0[2]),.dout(n1460),.clk(gclk));
	jor g1143(.dina(w_n1458_0[0]),.dinb(w_n486_0[0]),.dout(n1461),.clk(gclk));
	jand g1144(.dina(n1461),.dinb(n1460),.dout(n1462),.clk(gclk));
	jxor g1145(.dina(n1462),.dinb(w_n463_0[2]),.dout(n1463),.clk(gclk));
	jxor g1146(.dina(n1463),.dinb(n1456),.dout(n1464),.clk(gclk));
	jxor g1147(.dina(n1464),.dinb(n1451),.dout(n1465),.clk(gclk));
	jand g1148(.dina(n1465),.dinb(w_n700_0[1]),.dout(n1466),.clk(gclk));
	jand g1149(.dina(w_n496_0[0]),.dinb(w_n1340_0[0]),.dout(n1467),.clk(gclk));
	jor g1150(.dina(n1467),.dinb(w_n460_0[1]),.dout(n1468),.clk(gclk));
	jor g1151(.dina(w_n487_0[0]),.dinb(w_n491_0[1]),.dout(n1469),.clk(gclk));
	jand g1152(.dina(n1469),.dinb(w_n489_0[0]),.dout(n1470),.clk(gclk));
	jxor g1153(.dina(n1470),.dinb(w_n463_0[1]),.dout(n1471),.clk(gclk));
	jxor g1154(.dina(n1471),.dinb(w_n495_0[1]),.dout(n1472),.clk(gclk));
	jxor g1155(.dina(n1472),.dinb(w_n1452_0[0]),.dout(n1473),.clk(gclk));
	jxor g1156(.dina(n1473),.dinb(n1468),.dout(n1474),.clk(gclk));
	jand g1157(.dina(n1474),.dinb(w_n1321_0[1]),.dout(n1475),.clk(gclk));
	jor g1158(.dina(n1475),.dinb(n1466),.dout(n1476),.clk(gclk));
	jxor g1159(.dina(w_n470_0[0]),.dinb(w_n464_0[0]),.dout(n1477),.clk(gclk));
	jxor g1160(.dina(n1477),.dinb(n1476),.dout(n1478),.clk(gclk));
	jxor g1161(.dina(w_dff_B_wJPTGXyJ2_0),.dinb(n1449),.dout(w_dff_A_jSAFT7W59_2),.clk(gclk));
	jxor g1162(.dina(w_n416_0[0]),.dinb(w_n388_0[1]),.dout(n1480),.clk(gclk));
	jxor g1163(.dina(w_n411_0[1]),.dinb(w_n377_0[2]),.dout(n1481),.clk(gclk));
	jand g1164(.dina(w_n407_0[0]),.dinb(w_n1370_0[0]),.dout(n1482),.clk(gclk));
	jand g1165(.dina(w_n409_0[1]),.dinb(w_n392_0[0]),.dout(n1483),.clk(gclk));
	jor g1166(.dina(n1483),.dinb(n1482),.dout(n1484),.clk(gclk));
	jnot g1167(.din(w_n397_0[0]),.dout(n1485),.clk(gclk));
	jand g1168(.dina(n1485),.dinb(w_n405_0[0]),.dout(n1486),.clk(gclk));
	jxor g1169(.dina(w_n414_0[2]),.dinb(w_n396_0[2]),.dout(n1487),.clk(gclk));
	jxor g1170(.dina(n1487),.dinb(w_n1486_0[1]),.dout(n1488),.clk(gclk));
	jxor g1171(.dina(n1488),.dinb(n1484),.dout(n1489),.clk(gclk));
	jxor g1172(.dina(n1489),.dinb(n1481),.dout(n1490),.clk(gclk));
	jor g1173(.dina(n1490),.dinb(w_n707_0[2]),.dout(n1491),.clk(gclk));
	jor g1174(.dina(w_n391_0[0]),.dinb(w_n389_0[1]),.dout(n1492),.clk(gclk));
	jor g1175(.dina(w_n395_0[1]),.dinb(w_n393_0[1]),.dout(n1493),.clk(gclk));
	jand g1176(.dina(n1493),.dinb(w_n1492_0[1]),.dout(n1494),.clk(gclk));
	jnot g1177(.din(w_n1492_0[0]),.dout(n1495),.clk(gclk));
	jand g1178(.dina(w_n1486_0[0]),.dinb(n1495),.dout(n1496),.clk(gclk));
	jor g1179(.dina(n1496),.dinb(n1494),.dout(n1497),.clk(gclk));
	jxor g1180(.dina(w_n396_0[1]),.dinb(w_n377_0[1]),.dout(n1498),.clk(gclk));
	jxor g1181(.dina(n1498),.dinb(w_n1364_0[0]),.dout(n1499),.clk(gclk));
	jxor g1182(.dina(n1499),.dinb(n1497),.dout(n1500),.clk(gclk));
	jxor g1183(.dina(n1500),.dinb(w_n414_0[1]),.dout(n1501),.clk(gclk));
	jxor g1184(.dina(n1501),.dinb(w_n1359_0[0]),.dout(n1502),.clk(gclk));
	jor g1185(.dina(n1502),.dinb(w_n1337_0[2]),.dout(n1503),.clk(gclk));
	jand g1186(.dina(n1503),.dinb(n1491),.dout(n1504),.clk(gclk));
	jxor g1187(.dina(n1504),.dinb(n1480),.dout(n1505),.clk(gclk));
	jand g1188(.dina(w_n362_0[0]),.dinb(w_G38_0[2]),.dout(n1506),.clk(gclk));
	jnot g1189(.din(w_n364_0[1]),.dout(n1507),.clk(gclk));
	jor g1190(.dina(n1507),.dinb(w_n1506_0[1]),.dout(n1508),.clk(gclk));
	jnot g1191(.din(w_n1506_0[0]),.dout(n1509),.clk(gclk));
	jor g1192(.dina(n1509),.dinb(w_G1496_0[2]),.dout(n1510),.clk(gclk));
	jand g1193(.dina(n1510),.dinb(n1508),.dout(n1511),.clk(gclk));
	jand g1194(.dina(w_n1511_0[1]),.dinb(w_n413_0[2]),.dout(n1512),.clk(gclk));
	jnot g1195(.din(w_n413_0[1]),.dout(n1513),.clk(gclk));
	jand g1196(.dina(w_n712_0[0]),.dinb(w_n361_0[0]),.dout(n1514),.clk(gclk));
	jor g1197(.dina(w_n364_0[0]),.dinb(n1514),.dout(n1515),.clk(gclk));
	jor g1198(.dina(w_n369_0[0]),.dinb(w_G1492_0[2]),.dout(n1516),.clk(gclk));
	jand g1199(.dina(n1516),.dinb(n1515),.dout(n1517),.clk(gclk));
	jand g1200(.dina(n1517),.dinb(n1513),.dout(n1518),.clk(gclk));
	jor g1201(.dina(w_n1518_0[1]),.dinb(n1512),.dout(n1519),.clk(gclk));
	jor g1202(.dina(n1519),.dinb(w_n707_0[1]),.dout(n1520),.clk(gclk));
	jnot g1203(.din(w_n419_0[0]),.dout(n1521),.clk(gclk));
	jand g1204(.dina(w_n1518_0[0]),.dinb(n1521),.dout(n1522),.clk(gclk));
	jand g1205(.dina(w_n1511_0[0]),.dinb(w_n420_0[0]),.dout(n1523),.clk(gclk));
	jor g1206(.dina(n1523),.dinb(n1522),.dout(n1524),.clk(gclk));
	jor g1207(.dina(n1524),.dinb(w_n1337_0[1]),.dout(n1525),.clk(gclk));
	jand g1208(.dina(n1525),.dinb(n1520),.dout(n1526),.clk(gclk));
	jxor g1209(.dina(w_dff_B_Ecfi3mhT0_0),.dinb(n1505),.dout(w_dff_A_ViLkVnO16_2),.clk(gclk));
	jor g1210(.dina(w_n693_0[0]),.dinb(w_n687_0[0]),.dout(n1528),.clk(gclk));
	jand g1211(.dina(n1528),.dinb(w_n695_0[0]),.dout(n1529),.clk(gclk));
	jor g1212(.dina(w_n1529_0[1]),.dinb(w_n513_0[2]),.dout(n1530),.clk(gclk));
	jxor g1213(.dina(w_n1419_0[0]),.dinb(w_n1308_0[0]),.dout(n1531),.clk(gclk));
	jxor g1214(.dina(w_n1531_0[1]),.dinb(w_n526_0[0]),.dout(n1532),.clk(gclk));
	jxor g1215(.dina(n1532),.dinb(n1530),.dout(n1533),.clk(gclk));
	jand g1216(.dina(n1533),.dinb(w_n1309_0[0]),.dout(n1534),.clk(gclk));
	jand g1217(.dina(w_n1534_0[1]),.dinb(w_n1310_0[0]),.dout(n1535),.clk(gclk));
	jand g1218(.dina(w_n1426_0[0]),.dinb(w_n524_0[1]),.dout(n1536),.clk(gclk));
	jnot g1219(.din(w_n1536_0[1]),.dout(n1537),.clk(gclk));
	jor g1220(.dina(n1537),.dinb(w_n690_0[0]),.dout(n1538),.clk(gclk));
	jor g1221(.dina(w_n1536_0[0]),.dinb(w_n1529_0[0]),.dout(n1539),.clk(gclk));
	jand g1222(.dina(n1539),.dinb(n1538),.dout(n1540),.clk(gclk));
	jxor g1223(.dina(w_n518_0[1]),.dinb(w_n513_0[1]),.dout(n1541),.clk(gclk));
	jxor g1224(.dina(n1541),.dinb(w_n1531_0[0]),.dout(n1542),.clk(gclk));
	jxor g1225(.dina(n1542),.dinb(n1540),.dout(n1543),.clk(gclk));
	jor g1226(.dina(w_n581_0[0]),.dinb(w_n572_0[2]),.dout(n1544),.clk(gclk));
	jand g1227(.dina(n1544),.dinb(w_n1543_0[1]),.dout(n1545),.clk(gclk));
	jor g1228(.dina(n1545),.dinb(n1535),.dout(n1546),.clk(gclk));
	jand g1229(.dina(n1546),.dinb(w_n680_1[0]),.dout(n1547),.clk(gclk));
	jand g1230(.dina(w_n1543_0[0]),.dinb(w_n572_0[1]),.dout(n1548),.clk(gclk));
	jor g1231(.dina(n1548),.dinb(w_n1534_0[0]),.dout(n1549),.clk(gclk));
	jand g1232(.dina(n1549),.dinb(w_n1312_0[2]),.dout(n1550),.clk(gclk));
	jor g1233(.dina(n1550),.dinb(n1547),.dout(n1551),.clk(gclk));
	jxor g1234(.dina(w_n578_0[0]),.dinb(w_n1402_0[0]),.dout(n1552),.clk(gclk));
	jnot g1235(.din(w_n563_0[1]),.dout(n1553),.clk(gclk));
	jand g1236(.dina(n1553),.dinb(w_G4394_0[2]),.dout(n1554),.clk(gclk));
	jnot g1237(.din(w_n1554_0[1]),.dout(n1555),.clk(gclk));
	jand g1238(.dina(n1555),.dinb(w_n558_0[0]),.dout(n1556),.clk(gclk));
	jand g1239(.dina(w_n1554_0[0]),.dinb(w_n556_0[1]),.dout(n1557),.clk(gclk));
	jor g1240(.dina(n1557),.dinb(n1556),.dout(n1558),.clk(gclk));
	jxor g1241(.dina(n1558),.dinb(w_n573_0[2]),.dout(n1559),.clk(gclk));
	jxor g1242(.dina(n1559),.dinb(w_n1408_0[0]),.dout(n1560),.clk(gclk));
	jnot g1243(.din(w_n570_1[0]),.dout(n1561),.clk(gclk));
	jxor g1244(.dina(w_n575_0[1]),.dinb(w_n574_0[0]),.dout(n1562),.clk(gclk));
	jnot g1245(.din(w_n1562_0[2]),.dout(n1563),.clk(gclk));
	jor g1246(.dina(n1563),.dinb(n1561),.dout(n1564),.clk(gclk));
	jor g1247(.dina(w_n1562_0[1]),.dinb(w_n570_0[2]),.dout(n1565),.clk(gclk));
	jor g1248(.dina(n1565),.dinb(w_n580_0[0]),.dout(n1566),.clk(gclk));
	jand g1249(.dina(n1566),.dinb(n1564),.dout(n1567),.clk(gclk));
	jxor g1250(.dina(n1567),.dinb(n1560),.dout(n1568),.clk(gclk));
	jor g1251(.dina(n1568),.dinb(w_n1312_0[1]),.dout(n1569),.clk(gclk));
	jxor g1252(.dina(w_n1562_0[0]),.dinb(w_n570_0[1]),.dout(n1570),.clk(gclk));
	jnot g1253(.din(w_n565_0[0]),.dout(n1571),.clk(gclk));
	jor g1254(.dina(w_n564_0[0]),.dinb(w_n556_0[0]),.dout(n1572),.clk(gclk));
	jand g1255(.dina(n1572),.dinb(n1571),.dout(n1573),.clk(gclk));
	jxor g1256(.dina(n1573),.dinb(w_n573_0[1]),.dout(n1574),.clk(gclk));
	jxor g1257(.dina(n1574),.dinb(w_n568_0[0]),.dout(n1575),.clk(gclk));
	jxor g1258(.dina(n1575),.dinb(n1570),.dout(n1576),.clk(gclk));
	jor g1259(.dina(n1576),.dinb(w_n680_0[2]),.dout(n1577),.clk(gclk));
	jand g1260(.dina(n1577),.dinb(n1569),.dout(n1578),.clk(gclk));
	jxor g1261(.dina(n1578),.dinb(n1552),.dout(n1579),.clk(gclk));
	jxor g1262(.dina(n1579),.dinb(w_dff_B_ilTnKteO2_1),.dout(w_dff_A_zgLAj29Z1_2),.clk(gclk));
	jxor g1263(.dina(w_n1084_0[1]),.dinb(w_n1108_0[0]),.dout(n1581),.clk(gclk));
	jxor g1264(.dina(n1581),.dinb(w_n1105_0[0]),.dout(n1582),.clk(gclk));
	jand g1265(.dina(w_n616_0[0]),.dinb(w_n609_0[0]),.dout(n1583),.clk(gclk));
	jand g1266(.dina(w_n615_0[0]),.dinb(w_n610_0[0]),.dout(n1584),.clk(gclk));
	jor g1267(.dina(n1584),.dinb(n1583),.dout(n1585),.clk(gclk));
	jxor g1268(.dina(n1585),.dinb(n1582),.dout(n1586),.clk(gclk));
	jand g1269(.dina(n1586),.dinb(w_n1092_0[0]),.dout(n1587),.clk(gclk));
	jand g1270(.dina(w_n1587_0[1]),.dinb(w_n1086_0[0]),.dout(n1588),.clk(gclk));
	jnot g1271(.din(w_n598_0[1]),.dout(n1589),.clk(gclk));
	jand g1272(.dina(n1589),.dinb(w_G3737_0[1]),.dout(n1590),.clk(gclk));
	jand g1273(.dina(w_n1106_0[0]),.dinb(n1590),.dout(n1591),.clk(gclk));
	jand g1274(.dina(w_n613_0[0]),.dinb(w_n612_0[0]),.dout(n1592),.clk(gclk));
	jor g1275(.dina(n1592),.dinb(n1591),.dout(n1593),.clk(gclk));
	jor g1276(.dina(n1593),.dinb(w_n605_0[0]),.dout(n1594),.clk(gclk));
	jxor g1277(.dina(w_n1084_0[0]),.dinb(w_n594_0[0]),.dout(n1595),.clk(gclk));
	jxor g1278(.dina(n1595),.dinb(n1594),.dout(n1596),.clk(gclk));
	jxor g1279(.dina(n1596),.dinb(w_n619_0[0]),.dout(n1597),.clk(gclk));
	jand g1280(.dina(w_n1597_0[1]),.dinb(w_n674_0[0]),.dout(n1598),.clk(gclk));
	jor g1281(.dina(n1598),.dinb(w_n1094_0[1]),.dout(n1599),.clk(gclk));
	jor g1282(.dina(n1599),.dinb(n1588),.dout(n1600),.clk(gclk));
	jand g1283(.dina(w_n1597_0[0]),.dinb(w_n673_0[0]),.dout(n1601),.clk(gclk));
	jor g1284(.dina(n1601),.dinb(w_n1587_0[0]),.dout(n1602),.clk(gclk));
	jor g1285(.dina(n1602),.dinb(w_G4526_1[0]),.dout(n1603),.clk(gclk));
	jand g1286(.dina(n1603),.dinb(n1600),.dout(n1604),.clk(gclk));
	jxor g1287(.dina(w_n642_0[0]),.dinb(w_n359_0[1]),.dout(n1605),.clk(gclk));
	jxor g1288(.dina(w_n1605_0[1]),.dinb(w_n1067_0[1]),.dout(n1606),.clk(gclk));
	jxor g1289(.dina(n1606),.dinb(w_n1069_0[0]),.dout(n1607),.clk(gclk));
	jnot g1290(.din(w_n1607_0[1]),.dout(n1608),.clk(gclk));
	jxor g1291(.dina(w_n626_0[2]),.dinb(w_n354_0[0]),.dout(n1609),.clk(gclk));
	jxor g1292(.dina(n1609),.dinb(w_n671_0[0]),.dout(n1610),.clk(gclk));
	jor g1293(.dina(w_n1610_0[1]),.dinb(n1608),.dout(n1611),.clk(gclk));
	jnot g1294(.din(w_n1610_0[0]),.dout(n1612),.clk(gclk));
	jor g1295(.dina(n1612),.dinb(w_n1607_0[0]),.dout(n1613),.clk(gclk));
	jand g1296(.dina(n1613),.dinb(w_n1094_0[0]),.dout(n1614),.clk(gclk));
	jand g1297(.dina(n1614),.dinb(n1611),.dout(n1615),.clk(gclk));
	jand g1298(.dina(w_n1067_0[0]),.dinb(w_n357_0[0]),.dout(n1616),.clk(gclk));
	jand g1299(.dina(w_n661_0[0]),.dinb(w_n358_0[0]),.dout(n1617),.clk(gclk));
	jor g1300(.dina(n1617),.dinb(n1616),.dout(n1618),.clk(gclk));
	jxor g1301(.dina(n1618),.dinb(w_n626_0[1]),.dout(n1619),.clk(gclk));
	jxor g1302(.dina(n1619),.dinb(w_n1070_0[0]),.dout(n1620),.clk(gclk));
	jnot g1303(.din(w_n1620_0[1]),.dout(n1621),.clk(gclk));
	jnot g1304(.din(w_n645_0[0]),.dout(n1622),.clk(gclk));
	jand g1305(.dina(w_n1090_0[0]),.dinb(n1622),.dout(n1623),.clk(gclk));
	jxor g1306(.dina(n1623),.dinb(w_n1605_0[0]),.dout(n1624),.clk(gclk));
	jnot g1307(.din(w_n1624_0[1]),.dout(n1625),.clk(gclk));
	jor g1308(.dina(n1625),.dinb(n1621),.dout(n1626),.clk(gclk));
	jor g1309(.dina(w_n1624_0[0]),.dinb(w_n1620_0[0]),.dout(n1627),.clk(gclk));
	jand g1310(.dina(n1627),.dinb(w_G4526_0[2]),.dout(n1628),.clk(gclk));
	jand g1311(.dina(n1628),.dinb(n1626),.dout(n1629),.clk(gclk));
	jor g1312(.dina(n1629),.dinb(n1615),.dout(n1630),.clk(gclk));
	jxor g1313(.dina(w_n636_0[0]),.dinb(w_n631_0[0]),.dout(n1631),.clk(gclk));
	jxor g1314(.dina(n1631),.dinb(n1630),.dout(n1632),.clk(gclk));
	jxor g1315(.dina(n1632),.dinb(n1604),.dout(w_dff_A_h2dOt8HR5_2),.clk(gclk));
	jdff g1316(.din(w_G1_1[1]),.dout(w_dff_A_Dmc7a2bN2_1));
	jdff g1317(.din(w_G1_1[0]),.dout(w_dff_A_6v1KheBj0_1));
	jdff g1318(.din(w_G1459_0[0]),.dout(w_dff_A_P8WDRkB32_1));
	jdff g1319(.din(w_G1469_0[0]),.dout(w_dff_A_IflYUUBn6_1));
	jdff g1320(.din(w_G1480_0[0]),.dout(w_dff_A_U5TrYOk95_1));
	jdff g1321(.din(w_G1486_0[0]),.dout(w_dff_A_YONsQmPY7_1));
	jdff g1322(.din(w_G1492_0[1]),.dout(w_dff_A_7MrFhR7S7_1));
	jdff g1323(.din(w_G1496_0[1]),.dout(w_dff_A_pV3lp2Th7_1));
	jdff g1324(.din(w_G2208_0[0]),.dout(w_dff_A_GSYFA4ww3_1));
	jdff g1325(.din(w_G2218_0[0]),.dout(w_dff_A_FBQkF7m74_1));
	jdff g1326(.din(w_G2224_0[1]),.dout(w_dff_A_YfYhlcZP8_1));
	jdff g1327(.din(w_G2230_0[0]),.dout(w_dff_A_tzhGpJqn6_1));
	jdff g1328(.din(w_G2236_0[0]),.dout(w_dff_A_Wdw6GYOZ5_1));
	jdff g1329(.din(w_G2239_0[1]),.dout(w_dff_A_u6wSNtT59_1));
	jdff g1330(.din(w_G2247_0[0]),.dout(w_dff_A_PWRWabNi9_1));
	jdff g1331(.din(w_G2253_0[0]),.dout(w_dff_A_EMBTB4wN2_1));
	jdff g1332(.din(w_G2256_0[0]),.dout(w_dff_A_VAefslF47_1));
	jdff g1333(.din(w_G3698_0[0]),.dout(w_dff_A_upXkuxo17_1));
	jdff g1334(.din(w_G3701_0[1]),.dout(w_dff_A_lj9ELOAr8_1));
	jdff g1335(.din(w_G3705_0[1]),.dout(w_dff_A_sDPgk8v97_1));
	jdff g1336(.din(w_G3711_0[0]),.dout(w_dff_A_onEfvwvV6_1));
	jdff g1337(.din(w_G3717_0[0]),.dout(w_dff_A_XmweTCKr8_1));
	jdff g1338(.din(w_G3723_0[0]),.dout(w_dff_A_FwloGYnx1_1));
	jdff g1339(.din(w_G3729_0[1]),.dout(w_dff_A_gHt6hTma0_1));
	jdff g1340(.din(w_G3737_0[0]),.dout(w_dff_A_ljXzS98X0_1));
	jdff g1341(.din(w_G3743_0[0]),.dout(w_dff_A_xShgKWs03_1));
	jdff g1342(.din(w_G3749_0[0]),.dout(w_dff_A_38sqavEp5_1));
	jdff g1343(.din(w_G4393_0[0]),.dout(w_dff_A_DLdvL5Ht9_1));
	jdff g1344(.din(w_G4400_0[1]),.dout(w_dff_A_EW0imUD51_1));
	jdff g1345(.din(w_G4405_0[1]),.dout(w_dff_A_pZScGDyA2_1));
	jdff g1346(.din(w_G4410_0[0]),.dout(w_dff_A_s9CBI2X99_1));
	jdff g1347(.din(w_G4415_0[1]),.dout(w_dff_A_ltJWpPGm4_1));
	jdff g1348(.din(w_G4420_0[1]),.dout(w_dff_A_YJS1iCK09_1));
	jdff g1349(.din(w_G4427_0[0]),.dout(w_dff_A_ThUKi2cH2_1));
	jdff g1350(.din(w_G4432_0[0]),.dout(w_dff_A_7DWNk9T28_1));
	jdff g1351(.din(w_G4437_0[0]),.dout(w_dff_A_KWb9btUV8_1));
	jdff g1352(.din(w_G1462_0[0]),.dout(w_dff_A_mkapjFNr2_1));
	jdff g1353(.din(w_G2211_0[0]),.dout(w_dff_A_JNSQA5WW0_1));
	jdff g1354(.din(w_G4394_0[1]),.dout(w_dff_A_UcGMKMoa0_1));
	jdff g1355(.din(w_G1_0[2]),.dout(w_dff_A_UmRpndW02_1));
	jdff g1356(.din(w_G106_0[1]),.dout(w_dff_A_GvhcWMRm2_1));
	jnot g1357(.din(w_G15_0[1]),.dout(w_dff_A_80dpXEcR8_1),.clk(gclk));
	jor g1358(.dina(w_n345_0[0]),.dinb(w_G5_0[1]),.dout(w_dff_A_2ffOjGSw0_2),.clk(gclk));
	jnot g1359(.din(w_G15_0[0]),.dout(w_dff_A_5UJxVmwi0_1),.clk(gclk));
	jor g1360(.dina(w_n349_0[0]),.dinb(w_n347_0[0]),.dout(w_dff_A_LYTWwnQT3_2),.clk(gclk));
	jdff g1361(.din(w_G1_0[1]),.dout(w_dff_A_v6D1FION8_1));
	jand g1362(.dina(w_n1059_0[1]),.dinb(w_n718_0[1]),.dout(w_dff_A_gVGYXbAZ9_2),.clk(gclk));
	jor g1363(.dina(w_n715_1[0]),.dinb(w_n711_1[0]),.dout(G270),.clk(gclk));
	jand g1364(.dina(w_n1059_0[0]),.dinb(w_n718_0[0]),.dout(w_dff_A_82ekGnhb0_2),.clk(gclk));
	jor g1365(.dina(w_n715_0[2]),.dinb(w_n711_0[2]),.dout(G276),.clk(gclk));
	jor g1366(.dina(w_n715_0[1]),.dinb(w_n711_0[1]),.dout(G273),.clk(gclk));
	jxor g1367(.dina(w_n1396_0[0]),.dinb(w_n370_0[0]),.dout(G469),.clk(gclk));
	jxor g1368(.dina(w_n709_0[1]),.dinb(w_n363_0[0]),.dout(w_dff_A_RDG8Zhod6_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G5_0(.douta(w_G5_0[0]),.doutb(w_G5_0[1]),.doutc(w_G5_0[2]),.din(G5));
	jspl jspl_w_G5_1(.douta(w_dff_A_neoobXwD1_0),.doutb(w_G5_1[1]),.din(w_G5_0[0]));
	jspl3 jspl3_w_G15_0(.douta(w_G15_0[0]),.doutb(w_G15_0[1]),.doutc(w_G15_0[2]),.din(G15));
	jspl3 jspl3_w_G18_0(.douta(w_G18_0[0]),.doutb(w_G18_0[1]),.doutc(w_G18_0[2]),.din(G18));
	jspl3 jspl3_w_G18_1(.douta(w_G18_1[0]),.doutb(w_G18_1[1]),.doutc(w_G18_1[2]),.din(w_G18_0[0]));
	jspl3 jspl3_w_G18_2(.douta(w_G18_2[0]),.doutb(w_G18_2[1]),.doutc(w_G18_2[2]),.din(w_G18_0[1]));
	jspl3 jspl3_w_G18_3(.douta(w_G18_3[0]),.doutb(w_G18_3[1]),.doutc(w_G18_3[2]),.din(w_G18_0[2]));
	jspl3 jspl3_w_G18_4(.douta(w_G18_4[0]),.doutb(w_G18_4[1]),.doutc(w_G18_4[2]),.din(w_G18_1[0]));
	jspl3 jspl3_w_G18_5(.douta(w_G18_5[0]),.doutb(w_G18_5[1]),.doutc(w_G18_5[2]),.din(w_G18_1[1]));
	jspl3 jspl3_w_G18_6(.douta(w_G18_6[0]),.doutb(w_G18_6[1]),.doutc(w_G18_6[2]),.din(w_G18_1[2]));
	jspl3 jspl3_w_G18_7(.douta(w_G18_7[0]),.doutb(w_G18_7[1]),.doutc(w_G18_7[2]),.din(w_G18_2[0]));
	jspl3 jspl3_w_G18_8(.douta(w_G18_8[0]),.doutb(w_G18_8[1]),.doutc(w_G18_8[2]),.din(w_G18_2[1]));
	jspl3 jspl3_w_G18_9(.douta(w_G18_9[0]),.doutb(w_G18_9[1]),.doutc(w_G18_9[2]),.din(w_G18_2[2]));
	jspl3 jspl3_w_G18_10(.douta(w_G18_10[0]),.doutb(w_G18_10[1]),.doutc(w_G18_10[2]),.din(w_G18_3[0]));
	jspl3 jspl3_w_G18_11(.douta(w_G18_11[0]),.doutb(w_G18_11[1]),.doutc(w_G18_11[2]),.din(w_G18_3[1]));
	jspl3 jspl3_w_G18_12(.douta(w_G18_12[0]),.doutb(w_G18_12[1]),.doutc(w_G18_12[2]),.din(w_G18_3[2]));
	jspl3 jspl3_w_G18_13(.douta(w_G18_13[0]),.doutb(w_G18_13[1]),.doutc(w_G18_13[2]),.din(w_G18_4[0]));
	jspl3 jspl3_w_G18_14(.douta(w_G18_14[0]),.doutb(w_G18_14[1]),.doutc(w_G18_14[2]),.din(w_G18_4[1]));
	jspl3 jspl3_w_G18_15(.douta(w_G18_15[0]),.doutb(w_G18_15[1]),.doutc(w_G18_15[2]),.din(w_G18_4[2]));
	jspl3 jspl3_w_G18_16(.douta(w_G18_16[0]),.doutb(w_G18_16[1]),.doutc(w_G18_16[2]),.din(w_G18_5[0]));
	jspl3 jspl3_w_G18_17(.douta(w_G18_17[0]),.doutb(w_G18_17[1]),.doutc(w_G18_17[2]),.din(w_G18_5[1]));
	jspl3 jspl3_w_G18_18(.douta(w_G18_18[0]),.doutb(w_G18_18[1]),.doutc(w_G18_18[2]),.din(w_G18_5[2]));
	jspl3 jspl3_w_G18_19(.douta(w_G18_19[0]),.doutb(w_G18_19[1]),.doutc(w_G18_19[2]),.din(w_G18_6[0]));
	jspl3 jspl3_w_G18_20(.douta(w_G18_20[0]),.doutb(w_G18_20[1]),.doutc(w_G18_20[2]),.din(w_G18_6[1]));
	jspl3 jspl3_w_G18_21(.douta(w_G18_21[0]),.doutb(w_G18_21[1]),.doutc(w_G18_21[2]),.din(w_G18_6[2]));
	jspl3 jspl3_w_G18_22(.douta(w_G18_22[0]),.doutb(w_G18_22[1]),.doutc(w_G18_22[2]),.din(w_G18_7[0]));
	jspl3 jspl3_w_G18_23(.douta(w_G18_23[0]),.doutb(w_G18_23[1]),.doutc(w_G18_23[2]),.din(w_G18_7[1]));
	jspl3 jspl3_w_G18_24(.douta(w_G18_24[0]),.doutb(w_G18_24[1]),.doutc(w_G18_24[2]),.din(w_G18_7[2]));
	jspl3 jspl3_w_G18_25(.douta(w_G18_25[0]),.doutb(w_G18_25[1]),.doutc(w_G18_25[2]),.din(w_G18_8[0]));
	jspl3 jspl3_w_G18_26(.douta(w_G18_26[0]),.doutb(w_G18_26[1]),.doutc(w_G18_26[2]),.din(w_G18_8[1]));
	jspl3 jspl3_w_G18_27(.douta(w_G18_27[0]),.doutb(w_G18_27[1]),.doutc(w_G18_27[2]),.din(w_G18_8[2]));
	jspl3 jspl3_w_G18_28(.douta(w_G18_28[0]),.doutb(w_G18_28[1]),.doutc(w_G18_28[2]),.din(w_G18_9[0]));
	jspl3 jspl3_w_G18_29(.douta(w_G18_29[0]),.doutb(w_G18_29[1]),.doutc(w_G18_29[2]),.din(w_G18_9[1]));
	jspl3 jspl3_w_G18_30(.douta(w_G18_30[0]),.doutb(w_G18_30[1]),.doutc(w_G18_30[2]),.din(w_G18_9[2]));
	jspl3 jspl3_w_G18_31(.douta(w_G18_31[0]),.doutb(w_G18_31[1]),.doutc(w_G18_31[2]),.din(w_G18_10[0]));
	jspl3 jspl3_w_G18_32(.douta(w_G18_32[0]),.doutb(w_G18_32[1]),.doutc(w_G18_32[2]),.din(w_G18_10[1]));
	jspl3 jspl3_w_G18_33(.douta(w_G18_33[0]),.doutb(w_G18_33[1]),.doutc(w_G18_33[2]),.din(w_G18_10[2]));
	jspl3 jspl3_w_G18_34(.douta(w_G18_34[0]),.doutb(w_G18_34[1]),.doutc(w_G18_34[2]),.din(w_G18_11[0]));
	jspl3 jspl3_w_G18_35(.douta(w_G18_35[0]),.doutb(w_G18_35[1]),.doutc(w_G18_35[2]),.din(w_G18_11[1]));
	jspl3 jspl3_w_G18_36(.douta(w_G18_36[0]),.doutb(w_G18_36[1]),.doutc(w_G18_36[2]),.din(w_G18_11[2]));
	jspl3 jspl3_w_G18_37(.douta(w_G18_37[0]),.doutb(w_G18_37[1]),.doutc(w_G18_37[2]),.din(w_G18_12[0]));
	jspl3 jspl3_w_G18_38(.douta(w_G18_38[0]),.doutb(w_G18_38[1]),.doutc(w_G18_38[2]),.din(w_G18_12[1]));
	jspl3 jspl3_w_G18_39(.douta(w_G18_39[0]),.doutb(w_G18_39[1]),.doutc(w_G18_39[2]),.din(w_G18_12[2]));
	jspl3 jspl3_w_G18_40(.douta(w_G18_40[0]),.doutb(w_G18_40[1]),.doutc(w_G18_40[2]),.din(w_G18_13[0]));
	jspl3 jspl3_w_G18_41(.douta(w_G18_41[0]),.doutb(w_G18_41[1]),.doutc(w_G18_41[2]),.din(w_G18_13[1]));
	jspl3 jspl3_w_G18_42(.douta(w_G18_42[0]),.doutb(w_G18_42[1]),.doutc(w_G18_42[2]),.din(w_G18_13[2]));
	jspl3 jspl3_w_G18_43(.douta(w_G18_43[0]),.doutb(w_G18_43[1]),.doutc(w_G18_43[2]),.din(w_G18_14[0]));
	jspl3 jspl3_w_G18_44(.douta(w_G18_44[0]),.doutb(w_G18_44[1]),.doutc(w_G18_44[2]),.din(w_G18_14[1]));
	jspl3 jspl3_w_G18_45(.douta(w_G18_45[0]),.doutb(w_G18_45[1]),.doutc(w_G18_45[2]),.din(w_G18_14[2]));
	jspl3 jspl3_w_G18_46(.douta(w_G18_46[0]),.doutb(w_G18_46[1]),.doutc(w_G18_46[2]),.din(w_G18_15[0]));
	jspl3 jspl3_w_G18_47(.douta(w_G18_47[0]),.doutb(w_G18_47[1]),.doutc(w_G18_47[2]),.din(w_G18_15[1]));
	jspl3 jspl3_w_G18_48(.douta(w_G18_48[0]),.doutb(w_G18_48[1]),.doutc(w_G18_48[2]),.din(w_G18_15[2]));
	jspl3 jspl3_w_G18_49(.douta(w_G18_49[0]),.doutb(w_G18_49[1]),.doutc(w_G18_49[2]),.din(w_G18_16[0]));
	jspl jspl_w_G29_0(.douta(w_G29_0[0]),.doutb(w_G29_0[1]),.din(G29));
	jspl3 jspl3_w_G38_0(.douta(w_G38_0[0]),.doutb(w_G38_0[1]),.doutc(w_G38_0[2]),.din(G38));
	jspl3 jspl3_w_G38_1(.douta(w_G38_1[0]),.doutb(w_G38_1[1]),.doutc(w_G38_1[2]),.din(w_G38_0[0]));
	jspl3 jspl3_w_G38_2(.douta(w_G38_2[0]),.doutb(w_G38_2[1]),.doutc(w_G38_2[2]),.din(w_G38_0[1]));
	jspl jspl_w_G41_0(.douta(w_G41_0[0]),.doutb(w_G41_0[1]),.din(G41));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl jspl_w_G89_0(.douta(w_G89_0[0]),.doutb(w_G89_0[1]),.din(G89));
	jspl3 jspl3_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.doutc(w_G106_0[2]),.din(G106));
	jspl jspl_w_G106_1(.douta(w_G106_1[0]),.doutb(w_G106_1[1]),.din(w_G106_0[0]));
	jspl jspl_w_G209_0(.douta(w_G209_0[0]),.doutb(w_G209_0[1]),.din(G209));
	jspl jspl_w_G238_0(.douta(w_G238_0[0]),.doutb(w_G238_0[1]),.din(G238));
	jspl3 jspl3_w_G1455_0(.douta(w_G1455_0[0]),.doutb(w_G1455_0[1]),.doutc(w_G1455_0[2]),.din(G1455));
	jspl jspl_w_G1459_0(.douta(w_G1459_0[0]),.doutb(w_G1459_0[1]),.din(G1459));
	jspl jspl_w_G1462_0(.douta(w_G1462_0[0]),.doutb(w_G1462_0[1]),.din(G1462));
	jspl jspl_w_G1469_0(.douta(w_G1469_0[0]),.doutb(w_G1469_0[1]),.din(G1469));
	jspl3 jspl3_w_G1480_0(.douta(w_G1480_0[0]),.doutb(w_G1480_0[1]),.doutc(w_G1480_0[2]),.din(G1480));
	jspl jspl_w_G1486_0(.douta(w_G1486_0[0]),.doutb(w_G1486_0[1]),.din(G1486));
	jspl3 jspl3_w_G1492_0(.douta(w_G1492_0[0]),.doutb(w_G1492_0[1]),.doutc(w_G1492_0[2]),.din(G1492));
	jspl jspl_w_G1492_1(.douta(w_G1492_1[0]),.doutb(w_G1492_1[1]),.din(w_G1492_0[0]));
	jspl3 jspl3_w_G1496_0(.douta(w_G1496_0[0]),.doutb(w_G1496_0[1]),.doutc(w_G1496_0[2]),.din(G1496));
	jspl jspl_w_G1496_1(.douta(w_G1496_1[0]),.doutb(w_G1496_1[1]),.din(w_G1496_0[0]));
	jspl3 jspl3_w_G2204_0(.douta(w_G2204_0[0]),.doutb(w_G2204_0[1]),.doutc(w_G2204_0[2]),.din(G2204));
	jspl jspl_w_G2208_0(.douta(w_G2208_0[0]),.doutb(w_G2208_0[1]),.din(G2208));
	jspl3 jspl3_w_G2211_0(.douta(w_G2211_0[0]),.doutb(w_G2211_0[1]),.doutc(w_G2211_0[2]),.din(G2211));
	jspl3 jspl3_w_G2218_0(.douta(w_G2218_0[0]),.doutb(w_G2218_0[1]),.doutc(w_G2218_0[2]),.din(G2218));
	jspl3 jspl3_w_G2224_0(.douta(w_G2224_0[0]),.doutb(w_G2224_0[1]),.doutc(w_G2224_0[2]),.din(G2224));
	jspl jspl_w_G2224_1(.douta(w_G2224_1[0]),.doutb(w_G2224_1[1]),.din(w_G2224_0[0]));
	jspl3 jspl3_w_G2230_0(.douta(w_G2230_0[0]),.doutb(w_G2230_0[1]),.doutc(w_G2230_0[2]),.din(G2230));
	jspl3 jspl3_w_G2236_0(.douta(w_G2236_0[0]),.doutb(w_G2236_0[1]),.doutc(w_G2236_0[2]),.din(G2236));
	jspl3 jspl3_w_G2239_0(.douta(w_G2239_0[0]),.doutb(w_G2239_0[1]),.doutc(w_G2239_0[2]),.din(G2239));
	jspl jspl_w_G2239_1(.douta(w_G2239_1[0]),.doutb(w_G2239_1[1]),.din(w_G2239_0[0]));
	jspl3 jspl3_w_G2247_0(.douta(w_G2247_0[0]),.doutb(w_G2247_0[1]),.doutc(w_G2247_0[2]),.din(G2247));
	jspl3 jspl3_w_G2253_0(.douta(w_G2253_0[0]),.doutb(w_G2253_0[1]),.doutc(w_G2253_0[2]),.din(G2253));
	jspl jspl_w_G2256_0(.douta(w_G2256_0[0]),.doutb(w_G2256_0[1]),.din(G2256));
	jspl jspl_w_G3698_0(.douta(w_G3698_0[0]),.doutb(w_G3698_0[1]),.din(G3698));
	jspl3 jspl3_w_G3701_0(.douta(w_G3701_0[0]),.doutb(w_G3701_0[1]),.doutc(w_G3701_0[2]),.din(G3701));
	jspl jspl_w_G3701_1(.douta(w_G3701_1[0]),.doutb(w_G3701_1[1]),.din(w_G3701_0[0]));
	jspl3 jspl3_w_G3705_0(.douta(w_G3705_0[0]),.doutb(w_G3705_0[1]),.doutc(w_G3705_0[2]),.din(G3705));
	jspl3 jspl3_w_G3705_1(.douta(w_G3705_1[0]),.doutb(w_G3705_1[1]),.doutc(w_G3705_1[2]),.din(w_G3705_0[0]));
	jspl jspl_w_G3711_0(.douta(w_G3711_0[0]),.doutb(w_G3711_0[1]),.din(G3711));
	jspl3 jspl3_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_G3717_0[1]),.doutc(w_G3717_0[2]),.din(G3717));
	jspl3 jspl3_w_G3723_0(.douta(w_G3723_0[0]),.doutb(w_G3723_0[1]),.doutc(w_G3723_0[2]),.din(G3723));
	jspl3 jspl3_w_G3729_0(.douta(w_G3729_0[0]),.doutb(w_G3729_0[1]),.doutc(w_G3729_0[2]),.din(G3729));
	jspl jspl_w_G3729_1(.douta(w_G3729_1[0]),.doutb(w_G3729_1[1]),.din(w_G3729_0[0]));
	jspl3 jspl3_w_G3737_0(.douta(w_G3737_0[0]),.doutb(w_G3737_0[1]),.doutc(w_G3737_0[2]),.din(G3737));
	jspl3 jspl3_w_G3743_0(.douta(w_G3743_0[0]),.doutb(w_G3743_0[1]),.doutc(w_G3743_0[2]),.din(G3743));
	jspl3 jspl3_w_G3749_0(.douta(w_G3749_0[0]),.doutb(w_G3749_0[1]),.doutc(w_G3749_0[2]),.din(G3749));
	jspl jspl_w_G4393_0(.douta(w_G4393_0[0]),.doutb(w_G4393_0[1]),.din(G4393));
	jspl3 jspl3_w_G4394_0(.douta(w_G4394_0[0]),.doutb(w_G4394_0[1]),.doutc(w_G4394_0[2]),.din(G4394));
	jspl jspl_w_G4394_1(.douta(w_G4394_1[0]),.doutb(w_G4394_1[1]),.din(w_G4394_0[0]));
	jspl3 jspl3_w_G4400_0(.douta(w_G4400_0[0]),.doutb(w_G4400_0[1]),.doutc(w_G4400_0[2]),.din(G4400));
	jspl jspl_w_G4400_1(.douta(w_G4400_1[0]),.doutb(w_G4400_1[1]),.din(w_G4400_0[0]));
	jspl3 jspl3_w_G4405_0(.douta(w_G4405_0[0]),.doutb(w_G4405_0[1]),.doutc(w_G4405_0[2]),.din(G4405));
	jspl jspl_w_G4405_1(.douta(w_G4405_1[0]),.doutb(w_G4405_1[1]),.din(w_G4405_0[0]));
	jspl3 jspl3_w_G4410_0(.douta(w_G4410_0[0]),.doutb(w_G4410_0[1]),.doutc(w_G4410_0[2]),.din(G4410));
	jspl3 jspl3_w_G4415_0(.douta(w_G4415_0[0]),.doutb(w_G4415_0[1]),.doutc(w_G4415_0[2]),.din(G4415));
	jspl jspl_w_G4415_1(.douta(w_G4415_1[0]),.doutb(w_G4415_1[1]),.din(w_G4415_0[0]));
	jspl3 jspl3_w_G4420_0(.douta(w_G4420_0[0]),.doutb(w_G4420_0[1]),.doutc(w_G4420_0[2]),.din(G4420));
	jspl jspl_w_G4420_1(.douta(w_G4420_1[0]),.doutb(w_G4420_1[1]),.din(w_G4420_0[0]));
	jspl3 jspl3_w_G4427_0(.douta(w_G4427_0[0]),.doutb(w_G4427_0[1]),.doutc(w_G4427_0[2]),.din(G4427));
	jspl3 jspl3_w_G4432_0(.douta(w_G4432_0[0]),.doutb(w_G4432_0[1]),.doutc(w_G4432_0[2]),.din(G4432));
	jspl3 jspl3_w_G4437_0(.douta(w_G4437_0[0]),.doutb(w_G4437_0[1]),.doutc(w_G4437_0[2]),.din(G4437));
	jspl3 jspl3_w_G4526_0(.douta(w_G4526_0[0]),.doutb(w_G4526_0[1]),.doutc(w_G4526_0[2]),.din(G4526));
	jspl3 jspl3_w_G4526_1(.douta(w_G4526_1[0]),.doutb(w_G4526_1[1]),.doutc(w_G4526_1[2]),.din(w_G4526_0[0]));
	jspl3 jspl3_w_G4526_2(.douta(w_G4526_2[0]),.doutb(w_G4526_2[1]),.doutc(w_G4526_2[2]),.din(w_G4526_0[1]));
	jspl3 jspl3_w_G4528_0(.douta(w_G4528_0[0]),.doutb(w_G4528_0[1]),.doutc(w_G4528_0[2]),.din(G4528));
	jspl jspl_w_G404_0(.douta(w_G404_0),.doutb(w_dff_A_f9BvEB0p2_1),.din(G404_fa_));
	jspl jspl_w_G406_0(.douta(w_G406_0),.doutb(w_dff_A_cVJigQ0M0_1),.din(G406_fa_));
	jspl jspl_w_G408_0(.douta(w_G408_0),.doutb(w_dff_A_uXZKF6Yh3_1),.din(G408_fa_));
	jspl jspl_w_G410_0(.douta(w_G410_0),.doutb(w_dff_A_vLRVPHpJ9_1),.din(G410_fa_));
	jspl jspl_w_G412_0(.douta(w_G412_0),.doutb(w_dff_A_2m0EwwEg5_1),.din(G412_fa_));
	jspl jspl_w_G414_0(.douta(w_dff_A_76k9SREw6_0),.doutb(w_dff_A_67FtK3pA2_1),.din(G414_fa_));
	jspl jspl_w_G416_0(.douta(w_G416_0),.doutb(w_dff_A_uaKJXgnV6_1),.din(G416_fa_));
	jspl jspl_w_G252_0(.douta(w_G252_0),.doutb(w_dff_A_V1fSan9U2_1),.din(G252_fa_));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n347_0(.douta(w_n347_0[0]),.doutb(w_n347_0[1]),.din(w_dff_B_dY68LMNi2_2));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(n353));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(n354));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl3 jspl3_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.doutc(w_n355_1[2]),.din(w_n355_0[0]));
	jspl3 jspl3_w_n355_2(.douta(w_n355_2[0]),.doutb(w_n355_2[1]),.doutc(w_n355_2[2]),.din(w_n355_0[1]));
	jspl3 jspl3_w_n355_3(.douta(w_n355_3[0]),.doutb(w_n355_3[1]),.doutc(w_n355_3[2]),.din(w_n355_0[2]));
	jspl3 jspl3_w_n355_4(.douta(w_n355_4[0]),.doutb(w_n355_4[1]),.doutc(w_n355_4[2]),.din(w_n355_1[0]));
	jspl3 jspl3_w_n355_5(.douta(w_n355_5[0]),.doutb(w_n355_5[1]),.doutc(w_n355_5[2]),.din(w_n355_1[1]));
	jspl3 jspl3_w_n355_6(.douta(w_n355_6[0]),.doutb(w_n355_6[1]),.doutc(w_n355_6[2]),.din(w_n355_1[2]));
	jspl3 jspl3_w_n355_7(.douta(w_n355_7[0]),.doutb(w_n355_7[1]),.doutc(w_n355_7[2]),.din(w_n355_2[0]));
	jspl3 jspl3_w_n355_8(.douta(w_n355_8[0]),.doutb(w_n355_8[1]),.doutc(w_n355_8[2]),.din(w_n355_2[1]));
	jspl3 jspl3_w_n355_9(.douta(w_n355_9[0]),.doutb(w_n355_9[1]),.doutc(w_n355_9[2]),.din(w_n355_2[2]));
	jspl3 jspl3_w_n355_10(.douta(w_n355_10[0]),.doutb(w_n355_10[1]),.doutc(w_n355_10[2]),.din(w_n355_3[0]));
	jspl3 jspl3_w_n355_11(.douta(w_n355_11[0]),.doutb(w_n355_11[1]),.doutc(w_n355_11[2]),.din(w_n355_3[1]));
	jspl3 jspl3_w_n355_12(.douta(w_n355_12[0]),.doutb(w_n355_12[1]),.doutc(w_n355_12[2]),.din(w_n355_3[2]));
	jspl3 jspl3_w_n355_13(.douta(w_n355_13[0]),.doutb(w_n355_13[1]),.doutc(w_n355_13[2]),.din(w_n355_4[0]));
	jspl3 jspl3_w_n355_14(.douta(w_n355_14[0]),.doutb(w_n355_14[1]),.doutc(w_n355_14[2]),.din(w_n355_4[1]));
	jspl3 jspl3_w_n355_15(.douta(w_n355_15[0]),.doutb(w_n355_15[1]),.doutc(w_n355_15[2]),.din(w_n355_4[2]));
	jspl3 jspl3_w_n355_16(.douta(w_n355_16[0]),.doutb(w_n355_16[1]),.doutc(w_n355_16[2]),.din(w_n355_5[0]));
	jspl3 jspl3_w_n355_17(.douta(w_n355_17[0]),.doutb(w_n355_17[1]),.doutc(w_n355_17[2]),.din(w_n355_5[1]));
	jspl3 jspl3_w_n355_18(.douta(w_n355_18[0]),.doutb(w_n355_18[1]),.doutc(w_n355_18[2]),.din(w_n355_5[2]));
	jspl3 jspl3_w_n355_19(.douta(w_n355_19[0]),.doutb(w_n355_19[1]),.doutc(w_n355_19[2]),.din(w_n355_6[0]));
	jspl3 jspl3_w_n355_20(.douta(w_n355_20[0]),.doutb(w_n355_20[1]),.doutc(w_n355_20[2]),.din(w_n355_6[1]));
	jspl3 jspl3_w_n355_21(.douta(w_n355_21[0]),.doutb(w_n355_21[1]),.doutc(w_n355_21[2]),.din(w_n355_6[2]));
	jspl3 jspl3_w_n355_22(.douta(w_n355_22[0]),.doutb(w_n355_22[1]),.doutc(w_n355_22[2]),.din(w_n355_7[0]));
	jspl3 jspl3_w_n355_23(.douta(w_n355_23[0]),.doutb(w_n355_23[1]),.doutc(w_n355_23[2]),.din(w_n355_7[1]));
	jspl3 jspl3_w_n355_24(.douta(w_n355_24[0]),.doutb(w_n355_24[1]),.doutc(w_n355_24[2]),.din(w_n355_7[2]));
	jspl3 jspl3_w_n355_25(.douta(w_n355_25[0]),.doutb(w_n355_25[1]),.doutc(w_n355_25[2]),.din(w_n355_8[0]));
	jspl3 jspl3_w_n355_26(.douta(w_n355_26[0]),.doutb(w_n355_26[1]),.doutc(w_n355_26[2]),.din(w_n355_8[1]));
	jspl3 jspl3_w_n355_27(.douta(w_n355_27[0]),.doutb(w_n355_27[1]),.doutc(w_n355_27[2]),.din(w_n355_8[2]));
	jspl3 jspl3_w_n355_28(.douta(w_n355_28[0]),.doutb(w_n355_28[1]),.doutc(w_n355_28[2]),.din(w_n355_9[0]));
	jspl3 jspl3_w_n355_29(.douta(w_n355_29[0]),.doutb(w_n355_29[1]),.doutc(w_n355_29[2]),.din(w_n355_9[1]));
	jspl3 jspl3_w_n355_30(.douta(w_n355_30[0]),.doutb(w_n355_30[1]),.doutc(w_n355_30[2]),.din(w_n355_9[2]));
	jspl3 jspl3_w_n355_31(.douta(w_n355_31[0]),.doutb(w_n355_31[1]),.doutc(w_n355_31[2]),.din(w_n355_10[0]));
	jspl3 jspl3_w_n355_32(.douta(w_n355_32[0]),.doutb(w_n355_32[1]),.doutc(w_n355_32[2]),.din(w_n355_10[1]));
	jspl3 jspl3_w_n355_33(.douta(w_n355_33[0]),.doutb(w_n355_33[1]),.doutc(w_n355_33[2]),.din(w_n355_10[2]));
	jspl3 jspl3_w_n355_34(.douta(w_n355_34[0]),.doutb(w_n355_34[1]),.doutc(w_n355_34[2]),.din(w_n355_11[0]));
	jspl3 jspl3_w_n355_35(.douta(w_n355_35[0]),.doutb(w_n355_35[1]),.doutc(w_n355_35[2]),.din(w_n355_11[1]));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl3 jspl3_w_n359_0(.douta(w_n359_0[0]),.doutb(w_n359_0[1]),.doutc(w_n359_0[2]),.din(n359));
	jspl jspl_w_n359_1(.douta(w_n359_1[0]),.doutb(w_n359_1[1]),.din(w_n359_0[0]));
	jspl3 jspl3_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.doutc(w_n361_0[2]),.din(n361));
	jspl3 jspl3_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.doutc(w_n362_0[2]),.din(n362));
	jspl3 jspl3_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.doutc(w_n363_0[2]),.din(n363));
	jspl3 jspl3_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.doutc(w_n364_0[2]),.din(n364));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl3 jspl3_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.doutc(w_n370_0[2]),.din(n370));
	jspl3 jspl3_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.doutc(w_n371_0[2]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.doutc(w_n373_0[2]),.din(n373));
	jspl3 jspl3_w_n373_1(.douta(w_n373_1[0]),.doutb(w_n373_1[1]),.doutc(w_n373_1[2]),.din(w_n373_0[0]));
	jspl3 jspl3_w_n373_2(.douta(w_n373_2[0]),.doutb(w_n373_2[1]),.doutc(w_n373_2[2]),.din(w_n373_0[1]));
	jspl3 jspl3_w_n373_3(.douta(w_n373_3[0]),.doutb(w_n373_3[1]),.doutc(w_n373_3[2]),.din(w_n373_0[2]));
	jspl3 jspl3_w_n373_4(.douta(w_n373_4[0]),.doutb(w_n373_4[1]),.doutc(w_n373_4[2]),.din(w_n373_1[0]));
	jspl3 jspl3_w_n373_5(.douta(w_n373_5[0]),.doutb(w_n373_5[1]),.doutc(w_n373_5[2]),.din(w_n373_1[1]));
	jspl3 jspl3_w_n373_6(.douta(w_n373_6[0]),.doutb(w_n373_6[1]),.doutc(w_n373_6[2]),.din(w_n373_1[2]));
	jspl3 jspl3_w_n373_7(.douta(w_n373_7[0]),.doutb(w_n373_7[1]),.doutc(w_n373_7[2]),.din(w_n373_2[0]));
	jspl3 jspl3_w_n373_8(.douta(w_n373_8[0]),.doutb(w_n373_8[1]),.doutc(w_n373_8[2]),.din(w_n373_2[1]));
	jspl3 jspl3_w_n373_9(.douta(w_n373_9[0]),.doutb(w_n373_9[1]),.doutc(w_n373_9[2]),.din(w_n373_2[2]));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.din(n374));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_n377_0[2]),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.doutc(w_n377_1[2]),.din(w_n377_0[0]));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl3 jspl3_w_n379_0(.douta(w_n379_0[0]),.doutb(w_n379_0[1]),.doutc(w_n379_0[2]),.din(n379));
	jspl jspl_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.din(n380));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_n388_0[2]),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_n388_1[0]),.doutb(w_n388_1[1]),.doutc(w_n388_1[2]),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl jspl_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl3 jspl3_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.doutc(w_n392_0[2]),.din(n392));
	jspl3 jspl3_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.doutc(w_n393_0[2]),.din(n393));
	jspl jspl_w_n393_1(.douta(w_n393_1[0]),.doutb(w_n393_1[1]),.din(w_n393_0[0]));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl3 jspl3_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl jspl_w_n395_1(.douta(w_n395_1[0]),.doutb(w_n395_1[1]),.din(w_n395_0[0]));
	jspl3 jspl3_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.doutc(w_n396_0[2]),.din(n396));
	jspl3 jspl3_w_n396_1(.douta(w_n396_1[0]),.doutb(w_n396_1[1]),.doutc(w_n396_1[2]),.din(w_n396_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl3 jspl3_w_n409_0(.douta(w_n409_0[0]),.doutb(w_n409_0[1]),.doutc(w_n409_0[2]),.din(n409));
	jspl jspl_w_n409_1(.douta(w_n409_1[0]),.doutb(w_n409_1[1]),.din(w_n409_0[0]));
	jspl3 jspl3_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.doutc(w_n411_0[2]),.din(n411));
	jspl jspl_w_n411_1(.douta(w_n411_1[0]),.doutb(w_n411_1[1]),.din(w_n411_0[0]));
	jspl3 jspl3_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.doutc(w_n413_0[2]),.din(n413));
	jspl jspl_w_n413_1(.douta(w_n413_1[0]),.doutb(w_n413_1[1]),.din(w_n413_0[0]));
	jspl3 jspl3_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.doutc(w_n414_0[2]),.din(n414));
	jspl jspl_w_n414_1(.douta(w_n414_1[0]),.doutb(w_n414_1[1]),.din(w_n414_0[0]));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.doutc(w_n416_0[2]),.din(n416));
	jspl jspl_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.din(n418));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.din(n419));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl3 jspl3_w_n421_0(.douta(w_n421_0[0]),.doutb(w_n421_0[1]),.doutc(w_n421_0[2]),.din(n421));
	jspl jspl_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.din(n422));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl jspl_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.din(n424));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl jspl_w_n425_1(.douta(w_n425_1[0]),.doutb(w_n425_1[1]),.din(w_n425_0[0]));
	jspl3 jspl3_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.doutc(w_n426_0[2]),.din(n426));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(n427));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.doutc(w_n429_0[2]),.din(n429));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n431_0(.douta(w_n431_0[0]),.doutb(w_n431_0[1]),.din(n431));
	jspl3 jspl3_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.doutc(w_n432_0[2]),.din(n432));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_n433_0[2]),.din(n433));
	jspl3 jspl3_w_n433_1(.douta(w_n433_1[0]),.doutb(w_n433_1[1]),.doutc(w_n433_1[2]),.din(w_n433_0[0]));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.doutc(w_n437_0[2]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl3 jspl3_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.doutc(w_n444_0[2]),.din(n444));
	jspl3 jspl3_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.doutc(w_n445_0[2]),.din(n445));
	jspl3 jspl3_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.doutc(w_n447_0[2]),.din(n447));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl jspl_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.doutc(w_n450_0[2]),.din(n450));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.doutc(w_n451_0[2]),.din(n451));
	jspl3 jspl3_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.doutc(w_n453_0[2]),.din(n453));
	jspl jspl_w_n453_1(.douta(w_n453_1[0]),.doutb(w_n453_1[1]),.din(w_n453_0[0]));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.doutc(w_n456_0[2]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.doutc(w_n459_0[2]),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl3 jspl3_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.doutc(w_n463_0[2]),.din(n463));
	jspl jspl_w_n463_1(.douta(w_n463_1[0]),.doutb(w_n463_1[1]),.din(w_n463_0[0]));
	jspl3 jspl3_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.doutc(w_n464_0[2]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl3 jspl3_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.doutc(w_n469_0[2]),.din(n469));
	jspl jspl_w_n469_1(.douta(w_n469_1[0]),.doutb(w_n469_1[1]),.din(w_n469_0[0]));
	jspl3 jspl3_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.doutc(w_n470_0[2]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl3 jspl3_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.doutc(w_n474_0[2]),.din(n474));
	jspl3 jspl3_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.doutc(w_n475_0[2]),.din(n475));
	jspl3 jspl3_w_n476_0(.douta(w_n476_0[0]),.doutb(w_n476_0[1]),.doutc(w_n476_0[2]),.din(n476));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.doutc(w_n479_0[2]),.din(n479));
	jspl jspl_w_n479_1(.douta(w_n479_1[0]),.doutb(w_n479_1[1]),.din(w_n479_0[0]));
	jspl3 jspl3_w_n480_0(.douta(w_n480_0[0]),.doutb(w_n480_0[1]),.doutc(w_n480_0[2]),.din(n480));
	jspl jspl_w_n480_1(.douta(w_n480_1[0]),.doutb(w_n480_1[1]),.din(w_n480_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl jspl_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.din(n485));
	jspl jspl_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.din(n486));
	jspl3 jspl3_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.doutc(w_n487_0[2]),.din(n487));
	jspl3 jspl3_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.doutc(w_n489_0[2]),.din(n489));
	jspl3 jspl3_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.doutc(w_n491_0[2]),.din(n491));
	jspl jspl_w_n491_1(.douta(w_n491_1[0]),.doutb(w_n491_1[1]),.din(w_n491_0[0]));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl jspl_w_n495_1(.douta(w_n495_1[0]),.doutb(w_n495_1[1]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_n496_0[2]),.din(n496));
	jspl3 jspl3_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.doutc(w_n497_0[2]),.din(n497));
	jspl jspl_w_n497_1(.douta(w_n497_1[0]),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.din(n500));
	jspl3 jspl3_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.doutc(w_n501_0[2]),.din(n501));
	jspl jspl_w_n503_0(.douta(w_n503_0[0]),.doutb(w_n503_0[1]),.din(n503));
	jspl3 jspl3_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.doutc(w_n504_0[2]),.din(n504));
	jspl jspl_w_n504_1(.douta(w_n504_1[0]),.doutb(w_n504_1[1]),.din(w_n504_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl3 jspl3_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.doutc(w_n509_0[2]),.din(n509));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl3 jspl3_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.doutc(w_n512_0[2]),.din(n512));
	jspl3 jspl3_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.doutc(w_n513_0[2]),.din(n513));
	jspl jspl_w_n513_1(.douta(w_n513_1[0]),.doutb(w_n513_1[1]),.din(w_n513_0[0]));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl3 jspl3_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.doutc(w_n517_0[2]),.din(n517));
	jspl jspl_w_n517_1(.douta(w_n517_1[0]),.doutb(w_n517_1[1]),.din(w_n517_0[0]));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl3 jspl3_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.doutc(w_n524_0[2]),.din(n524));
	jspl3 jspl3_w_n524_1(.douta(w_n524_1[0]),.doutb(w_n524_1[1]),.doutc(w_n524_1[2]),.din(w_n524_0[0]));
	jspl3 jspl3_w_n526_0(.douta(w_n526_0[0]),.doutb(w_n526_0[1]),.doutc(w_n526_0[2]),.din(n526));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(n530));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.doutc(w_n531_0[2]),.din(n531));
	jspl jspl_w_n531_1(.douta(w_n531_1[0]),.doutb(w_n531_1[1]),.din(w_n531_0[0]));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.doutc(w_n536_0[2]),.din(n536));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl jspl_w_n539_1(.douta(w_n539_1[0]),.doutb(w_n539_1[1]),.din(w_n539_0[0]));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n546_0(.douta(w_n546_0[0]),.doutb(w_n546_0[1]),.din(n546));
	jspl3 jspl3_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.doutc(w_n547_0[2]),.din(n547));
	jspl jspl_w_n547_1(.douta(w_n547_1[0]),.doutb(w_n547_1[1]),.din(w_n547_0[0]));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(n552));
	jspl jspl_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.din(n554));
	jspl3 jspl3_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.doutc(w_n555_0[2]),.din(n555));
	jspl jspl_w_n555_1(.douta(w_n555_1[0]),.doutb(w_n555_1[1]),.din(w_n555_0[0]));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl jspl_w_n558_0(.douta(w_n558_0[0]),.doutb(w_n558_0[1]),.din(n558));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.doutc(w_n563_0[2]),.din(n563));
	jspl jspl_w_n563_1(.douta(w_n563_1[0]),.doutb(w_n563_1[1]),.din(w_n563_0[0]));
	jspl3 jspl3_w_n564_0(.douta(w_n564_0[0]),.doutb(w_n564_0[1]),.doutc(w_n564_0[2]),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.doutc(w_n568_0[2]),.din(n568));
	jspl3 jspl3_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.doutc(w_n570_0[2]),.din(n570));
	jspl3 jspl3_w_n570_1(.douta(w_n570_1[0]),.doutb(w_n570_1[1]),.doutc(w_n570_1[2]),.din(w_n570_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl jspl_w_n572_1(.douta(w_n572_1[0]),.doutb(w_n572_1[1]),.din(w_n572_0[0]));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl jspl_w_n573_1(.douta(w_n573_1[0]),.doutb(w_n573_1[1]),.din(w_n573_0[0]));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.doutc(w_n575_0[2]),.din(n575));
	jspl jspl_w_n575_1(.douta(w_n575_1[0]),.doutb(w_n575_1[1]),.din(w_n575_0[0]));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.doutc(w_n580_0[2]),.din(n580));
	jspl3 jspl3_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.doutc(w_n581_0[2]),.din(n581));
	jspl3 jspl3_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.doutc(w_n582_0[2]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl3 jspl3_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.doutc(w_n585_0[2]),.din(n585));
	jspl jspl_w_n585_1(.douta(w_n585_1[0]),.doutb(w_n585_1[1]),.din(w_n585_0[0]));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(n588));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.doutc(w_n590_0[2]),.din(n590));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(n592));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n593_1(.douta(w_n593_1[0]),.doutb(w_n593_1[1]),.din(w_n593_0[0]));
	jspl3 jspl3_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.doutc(w_n594_0[2]),.din(n594));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl3 jspl3_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.doutc(w_n598_0[2]),.din(n598));
	jspl jspl_w_n598_1(.douta(w_n598_1[0]),.doutb(w_n598_1[1]),.din(w_n598_0[0]));
	jspl3 jspl3_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.doutc(w_n599_0[2]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.doutc(w_n603_0[2]),.din(n603));
	jspl jspl_w_n603_1(.douta(w_n603_1[0]),.doutb(w_n603_1[1]),.din(w_n603_0[0]));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n610_0(.douta(w_n610_0[0]),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.doutc(w_n615_0[2]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n625_1(.douta(w_n625_1[0]),.doutb(w_n625_1[1]),.din(w_n625_0[0]));
	jspl3 jspl3_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.doutc(w_n626_0[2]),.din(n626));
	jspl jspl_w_n626_1(.douta(w_n626_1[0]),.doutb(w_n626_1[1]),.din(w_n626_0[0]));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.doutc(w_n631_0[2]),.din(n631));
	jspl3 jspl3_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.doutc(w_n632_0[2]),.din(n632));
	jspl jspl_w_n632_1(.douta(w_n632_1[0]),.doutb(w_n632_1[1]),.din(w_n632_0[0]));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_n635_1[0]),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_n641_0[2]),.din(n641));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.doutc(w_n642_0[2]),.din(n642));
	jspl jspl_w_n644_0(.douta(w_n644_0[0]),.doutb(w_n644_0[1]),.din(n644));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.din(n646));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.din(n653));
	jspl3 jspl3_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.doutc(w_n654_0[2]),.din(n654));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n656_0(.douta(w_n656_0[0]),.doutb(w_n656_0[1]),.din(n656));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.doutc(w_n657_0[2]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_n660_0[2]),.din(n660));
	jspl3 jspl3_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.doutc(w_n661_0[2]),.din(n661));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl3 jspl3_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.doutc(w_n663_0[2]),.din(n663));
	jspl jspl_w_n663_1(.douta(w_n663_1[0]),.doutb(w_n663_1[1]),.din(w_n663_0[0]));
	jspl jspl_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.din(n664));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(n669));
	jspl jspl_w_n671_0(.douta(w_n671_0[0]),.doutb(w_n671_0[1]),.din(n671));
	jspl3 jspl3_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.doutc(w_n673_0[2]),.din(n673));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(n674));
	jspl3 jspl3_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.doutc(w_n680_0[2]),.din(n680));
	jspl3 jspl3_w_n680_1(.douta(w_n680_1[0]),.doutb(w_n680_1[1]),.doutc(w_n680_1[2]),.din(w_n680_0[0]));
	jspl3 jspl3_w_n680_2(.douta(w_n680_2[0]),.doutb(w_n680_2[1]),.doutc(w_n680_2[2]),.din(w_n680_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.din(n694));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(n696));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl3 jspl3_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.doutc(w_n700_0[2]),.din(n700));
	jspl jspl_w_n700_1(.douta(w_n700_1[0]),.doutb(w_n700_1[1]),.din(w_n700_0[0]));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl3 jspl3_w_n703_1(.douta(w_n703_1[0]),.doutb(w_n703_1[1]),.doutc(w_n703_1[2]),.din(w_n703_0[0]));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl3 jspl3_w_n707_1(.douta(w_n707_1[0]),.doutb(w_n707_1[1]),.doutc(w_n707_1[2]),.din(w_n707_0[0]));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl3 jspl3_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.doutc(w_n711_0[2]),.din(n711));
	jspl jspl_w_n711_1(.douta(w_n711_1[0]),.doutb(w_n711_1[1]),.din(w_n711_0[0]));
	jspl3 jspl3_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.doutc(w_n712_0[2]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(w_dff_B_p1zgFYqg9_3));
	jspl jspl_w_n715_1(.douta(w_n715_1[0]),.doutb(w_n715_1[1]),.din(w_n715_0[0]));
	jspl3 jspl3_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.doutc(w_n718_0[2]),.din(w_dff_B_4D5BXUHe7_3));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(n719));
	jspl3 jspl3_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.doutc(w_n720_0[2]),.din(n720));
	jspl3 jspl3_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.doutc(w_n723_0[2]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.din(n725));
	jspl3 jspl3_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.doutc(w_n726_0[2]),.din(n726));
	jspl jspl_w_n726_1(.douta(w_n726_1[0]),.doutb(w_n726_1[1]),.din(w_n726_0[0]));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.doutc(w_n734_0[2]),.din(n734));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl jspl_w_n737_1(.douta(w_n737_1[0]),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n741_1(.douta(w_n741_1[0]),.doutb(w_n741_1[1]),.din(w_n741_0[0]));
	jspl jspl_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.din(n743));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_n744_0[2]),.din(n744));
	jspl3 jspl3_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.doutc(w_n747_0[2]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(n749));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.doutc(w_n755_0[2]),.din(n755));
	jspl jspl_w_n755_1(.douta(w_n755_1[0]),.doutb(w_n755_1[1]),.din(w_n755_0[0]));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_n758_1[1]),.din(w_n758_0[0]));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.doutc(w_n761_0[2]),.din(n761));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_n764_0[2]),.din(n764));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(n766));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl3 jspl3_w_n768_0(.douta(w_n768_0[0]),.doutb(w_n768_0[1]),.doutc(w_n768_0[2]),.din(n768));
	jspl3 jspl3_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.doutc(w_n772_0[2]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl3 jspl3_w_n776_0(.douta(w_n776_0[0]),.doutb(w_n776_0[1]),.doutc(w_n776_0[2]),.din(n776));
	jspl3 jspl3_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.doutc(w_n780_0[2]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(n781));
	jspl3 jspl3_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.doutc(w_n796_0[2]),.din(n796));
	jspl jspl_w_n796_1(.douta(w_n796_1[0]),.doutb(w_n796_1[1]),.din(w_n796_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.doutc(w_n800_0[2]),.din(n800));
	jspl jspl_w_n800_1(.douta(w_n800_1[0]),.doutb(w_n800_1[1]),.din(w_n800_0[0]));
	jspl3 jspl3_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.doutc(w_n803_0[2]),.din(n803));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl3 jspl3_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.doutc(w_n810_0[2]),.din(n810));
	jspl jspl_w_n810_1(.douta(w_n810_1[0]),.doutb(w_n810_1[1]),.din(w_n810_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.doutc(w_n814_0[2]),.din(n814));
	jspl jspl_w_n814_1(.douta(w_n814_1[0]),.doutb(w_n814_1[1]),.din(w_n814_0[0]));
	jspl3 jspl3_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.doutc(w_n817_0[2]),.din(n817));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl3 jspl3_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.doutc(w_n824_0[2]),.din(n824));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.doutc(w_n845_0[2]),.din(n845));
	jspl jspl_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n848_0(.douta(w_n848_0[0]),.doutb(w_n848_0[1]),.doutc(w_n848_0[2]),.din(n848));
	jspl jspl_w_n848_1(.douta(w_n848_1[0]),.doutb(w_n848_1[1]),.din(w_n848_0[0]));
	jspl3 jspl3_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.doutc(w_n851_0[2]),.din(n851));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.doutc(w_n854_0[2]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl3 jspl3_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.doutc(w_n858_0[2]),.din(n858));
	jspl3 jspl3_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.doutc(w_n862_0[2]),.din(n862));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl3 jspl3_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.doutc(w_n866_0[2]),.din(n866));
	jspl3 jspl3_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.doutc(w_n870_0[2]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl3 jspl3_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.doutc(w_n885_0[2]),.din(n885));
	jspl3 jspl3_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.doutc(w_n888_0[2]),.din(n888));
	jspl3 jspl3_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.doutc(w_n891_0[2]),.din(n891));
	jspl3 jspl3_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.doutc(w_n894_0[2]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.doutc(w_n900_0[2]),.din(n900));
	jspl3 jspl3_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.doutc(w_n903_0[2]),.din(n903));
	jspl jspl_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.din(n905));
	jspl3 jspl3_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.doutc(w_n916_0[2]),.din(n916));
	jspl3 jspl3_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.doutc(w_n919_0[2]),.din(n919));
	jspl3 jspl3_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.doutc(w_n926_0[2]),.din(n926));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_n930_0[2]),.din(n930));
	jspl3 jspl3_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.doutc(w_n935_0[2]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.doutc(w_n938_0[2]),.din(n938));
	jspl3 jspl3_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.doutc(w_n944_0[2]),.din(n944));
	jspl3 jspl3_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.doutc(w_n947_0[2]),.din(n947));
	jspl3 jspl3_w_n950_0(.douta(w_n950_0[0]),.doutb(w_n950_0[1]),.doutc(w_n950_0[2]),.din(n950));
	jspl jspl_w_n950_1(.douta(w_n950_1[0]),.doutb(w_n950_1[1]),.din(w_n950_0[0]));
	jspl3 jspl3_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.doutc(w_n953_0[2]),.din(n953));
	jspl jspl_w_n953_1(.douta(w_n953_1[0]),.doutb(w_n953_1[1]),.din(w_n953_0[0]));
	jspl3 jspl3_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.doutc(w_n966_0[2]),.din(n966));
	jspl3 jspl3_w_n970_0(.douta(w_n970_0[0]),.doutb(w_n970_0[1]),.doutc(w_n970_0[2]),.din(n970));
	jspl3 jspl3_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.doutc(w_n973_0[2]),.din(n973));
	jspl jspl_w_n973_1(.douta(w_n973_1[0]),.doutb(w_n973_1[1]),.din(w_n973_0[0]));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n977_1(.douta(w_n977_1[0]),.doutb(w_n977_1[1]),.din(w_n977_0[0]));
	jspl3 jspl3_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.doutc(w_n980_0[2]),.din(n980));
	jspl3 jspl3_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.doutc(w_n983_0[2]),.din(n983));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.doutc(w_n995_0[2]),.din(n995));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1042_0(.douta(w_n1042_0[0]),.doutb(w_n1042_0[1]),.din(n1042));
	jspl3 jspl3_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.doutc(w_n1059_0[2]),.din(n1059));
	jspl3 jspl3_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.doutc(w_n1067_0[2]),.din(n1067));
	jspl3 jspl3_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.doutc(w_n1069_0[2]),.din(n1069));
	jspl jspl_w_n1070_0(.douta(w_n1070_0[0]),.doutb(w_n1070_0[1]),.din(n1070));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(n1073));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl3 jspl3_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.doutc(w_n1084_0[2]),.din(n1084));
	jspl jspl_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.din(n1086));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl3 jspl3_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.doutc(w_n1092_0[2]),.din(n1092));
	jspl3 jspl3_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.doutc(w_n1094_0[2]),.din(n1094));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_n1106_0[1]),.din(n1106));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_n1108_0[1]),.din(n1108));
	jspl jspl_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_n1113_0[1]),.din(n1113));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(n1127));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1150_0(.douta(w_n1150_0[0]),.doutb(w_n1150_0[1]),.din(n1150));
	jspl jspl_w_n1172_0(.douta(w_n1172_0[0]),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_n1308_0[1]),.din(n1308));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl3 jspl3_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.doutc(w_n1312_0[2]),.din(n1312));
	jspl jspl_w_n1312_1(.douta(w_n1312_1[0]),.doutb(w_n1312_1[1]),.din(w_n1312_0[0]));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(n1316));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl3 jspl3_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.doutc(w_n1321_0[2]),.din(n1321));
	jspl jspl_w_n1321_1(.douta(w_n1321_1[0]),.doutb(w_n1321_1[1]),.din(w_n1321_0[0]));
	jspl jspl_w_n1323_0(.douta(w_n1323_0[0]),.doutb(w_n1323_0[1]),.din(n1323));
	jspl jspl_w_n1333_0(.douta(w_n1333_0[0]),.doutb(w_n1333_0[1]),.din(n1333));
	jspl3 jspl3_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.doutc(w_n1337_0[2]),.din(n1337));
	jspl jspl_w_n1337_1(.douta(w_n1337_1[0]),.doutb(w_n1337_1[1]),.din(w_n1337_0[0]));
	jspl3 jspl3_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.doutc(w_n1340_0[2]),.din(n1340));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(n1343));
	jspl jspl_w_n1344_0(.douta(w_n1344_0[0]),.doutb(w_n1344_0[1]),.din(n1344));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(n1364));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_n1370_0[1]),.din(n1370));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1387_0(.douta(w_n1387_0[0]),.doutb(w_n1387_0[1]),.din(n1387));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.din(n1388));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.din(n1402));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_n1408_0[1]),.din(n1408));
	jspl jspl_w_n1419_0(.douta(w_n1419_0[0]),.doutb(w_n1419_0[1]),.din(n1419));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(n1426));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(n1431));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(n1440));
	jspl3 jspl3_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.doutc(w_n1452_0[2]),.din(n1452));
	jspl jspl_w_n1458_0(.douta(w_n1458_0[0]),.doutb(w_n1458_0[1]),.din(n1458));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl jspl_w_n1492_0(.douta(w_n1492_0[0]),.doutb(w_n1492_0[1]),.din(n1492));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1511_0(.douta(w_n1511_0[0]),.doutb(w_n1511_0[1]),.din(n1511));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(n1531));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1536_0(.douta(w_n1536_0[0]),.doutb(w_n1536_0[1]),.din(n1536));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl3 jspl3_w_n1562_0(.douta(w_n1562_0[0]),.doutb(w_n1562_0[1]),.doutc(w_n1562_0[2]),.din(n1562));
	jspl jspl_w_n1587_0(.douta(w_n1587_0[0]),.doutb(w_n1587_0[1]),.din(n1587));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1620_0(.douta(w_n1620_0[0]),.doutb(w_n1620_0[1]),.din(n1620));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(n1624));
	jdff dff_A_neoobXwD1_0(.dout(w_G5_1[0]),.din(w_dff_A_neoobXwD1_0),.clk(gclk));
	jdff dff_B_dY68LMNi2_2(.din(n347),.dout(w_dff_B_dY68LMNi2_2),.clk(gclk));
	jdff dff_B_c1VlsQ6b8_1(.din(n1085),.dout(w_dff_B_c1VlsQ6b8_1),.clk(gclk));
	jdff dff_B_LG1bYm0e9_1(.din(n753),.dout(w_dff_B_LG1bYm0e9_1),.clk(gclk));
	jdff dff_B_RPUVOxCn0_1(.din(w_dff_B_LG1bYm0e9_1),.dout(w_dff_B_RPUVOxCn0_1),.clk(gclk));
	jdff dff_B_TKq0mV5z9_1(.din(w_dff_B_RPUVOxCn0_1),.dout(w_dff_B_TKq0mV5z9_1),.clk(gclk));
	jdff dff_B_GqewLBi55_1(.din(w_dff_B_TKq0mV5z9_1),.dout(w_dff_B_GqewLBi55_1),.clk(gclk));
	jdff dff_B_GMI6467M9_1(.din(w_dff_B_GqewLBi55_1),.dout(w_dff_B_GMI6467M9_1),.clk(gclk));
	jdff dff_B_aAztm4hS6_1(.din(w_dff_B_GMI6467M9_1),.dout(w_dff_B_aAztm4hS6_1),.clk(gclk));
	jdff dff_B_aQ5P1FDE8_1(.din(w_dff_B_aAztm4hS6_1),.dout(w_dff_B_aQ5P1FDE8_1),.clk(gclk));
	jdff dff_B_7qGpVZ1P4_1(.din(w_dff_B_aQ5P1FDE8_1),.dout(w_dff_B_7qGpVZ1P4_1),.clk(gclk));
	jdff dff_B_DEDLvIgL1_1(.din(w_dff_B_7qGpVZ1P4_1),.dout(w_dff_B_DEDLvIgL1_1),.clk(gclk));
	jdff dff_B_I3uFP1fQ7_1(.din(w_dff_B_DEDLvIgL1_1),.dout(w_dff_B_I3uFP1fQ7_1),.clk(gclk));
	jdff dff_B_NLE5NhC27_1(.din(w_dff_B_I3uFP1fQ7_1),.dout(w_dff_B_NLE5NhC27_1),.clk(gclk));
	jdff dff_B_vjfIi28Z3_1(.din(w_dff_B_NLE5NhC27_1),.dout(w_dff_B_vjfIi28Z3_1),.clk(gclk));
	jdff dff_B_ZngyyZX71_1(.din(w_dff_B_vjfIi28Z3_1),.dout(w_dff_B_ZngyyZX71_1),.clk(gclk));
	jdff dff_B_yodZqdA21_1(.din(w_dff_B_ZngyyZX71_1),.dout(w_dff_B_yodZqdA21_1),.clk(gclk));
	jdff dff_B_rOvy3G2j8_1(.din(w_dff_B_yodZqdA21_1),.dout(w_dff_B_rOvy3G2j8_1),.clk(gclk));
	jdff dff_B_NI6Dgyqd3_1(.din(w_dff_B_rOvy3G2j8_1),.dout(w_dff_B_NI6Dgyqd3_1),.clk(gclk));
	jdff dff_B_B6UBMEla4_1(.din(w_dff_B_NI6Dgyqd3_1),.dout(w_dff_B_B6UBMEla4_1),.clk(gclk));
	jdff dff_B_OsxWh6Gu4_0(.din(n1057),.dout(w_dff_B_OsxWh6Gu4_0),.clk(gclk));
	jdff dff_B_uAtrPtaT2_0(.din(w_dff_B_OsxWh6Gu4_0),.dout(w_dff_B_uAtrPtaT2_0),.clk(gclk));
	jdff dff_B_CwMfwXe77_0(.din(w_dff_B_uAtrPtaT2_0),.dout(w_dff_B_CwMfwXe77_0),.clk(gclk));
	jdff dff_B_vazfz53v6_0(.din(w_dff_B_CwMfwXe77_0),.dout(w_dff_B_vazfz53v6_0),.clk(gclk));
	jdff dff_B_ZAryOtFP5_0(.din(w_dff_B_vazfz53v6_0),.dout(w_dff_B_ZAryOtFP5_0),.clk(gclk));
	jdff dff_B_0AWBxpFH7_0(.din(w_dff_B_ZAryOtFP5_0),.dout(w_dff_B_0AWBxpFH7_0),.clk(gclk));
	jdff dff_B_yoCuqTVD0_0(.din(w_dff_B_0AWBxpFH7_0),.dout(w_dff_B_yoCuqTVD0_0),.clk(gclk));
	jdff dff_B_8cVb4XS05_0(.din(w_dff_B_yoCuqTVD0_0),.dout(w_dff_B_8cVb4XS05_0),.clk(gclk));
	jdff dff_B_qEBw09743_0(.din(w_dff_B_8cVb4XS05_0),.dout(w_dff_B_qEBw09743_0),.clk(gclk));
	jdff dff_B_UeaNXdH80_0(.din(w_dff_B_qEBw09743_0),.dout(w_dff_B_UeaNXdH80_0),.clk(gclk));
	jdff dff_B_2yWoyz8V1_0(.din(w_dff_B_UeaNXdH80_0),.dout(w_dff_B_2yWoyz8V1_0),.clk(gclk));
	jdff dff_B_S7gC4XIz8_0(.din(w_dff_B_2yWoyz8V1_0),.dout(w_dff_B_S7gC4XIz8_0),.clk(gclk));
	jdff dff_B_iJsdmYZJ1_0(.din(w_dff_B_S7gC4XIz8_0),.dout(w_dff_B_iJsdmYZJ1_0),.clk(gclk));
	jdff dff_B_yUS5D9F94_0(.din(w_dff_B_iJsdmYZJ1_0),.dout(w_dff_B_yUS5D9F94_0),.clk(gclk));
	jdff dff_B_HJqdpYuJ8_0(.din(w_dff_B_yUS5D9F94_0),.dout(w_dff_B_HJqdpYuJ8_0),.clk(gclk));
	jdff dff_B_POG4d9VZ1_0(.din(w_dff_B_HJqdpYuJ8_0),.dout(w_dff_B_POG4d9VZ1_0),.clk(gclk));
	jdff dff_B_FddPjT129_0(.din(n1044),.dout(w_dff_B_FddPjT129_0),.clk(gclk));
	jdff dff_B_uJkImova9_0(.din(w_dff_B_FddPjT129_0),.dout(w_dff_B_uJkImova9_0),.clk(gclk));
	jdff dff_B_3Y8BuPAf9_0(.din(w_dff_B_uJkImova9_0),.dout(w_dff_B_3Y8BuPAf9_0),.clk(gclk));
	jdff dff_B_23I2t5e54_0(.din(w_dff_B_3Y8BuPAf9_0),.dout(w_dff_B_23I2t5e54_0),.clk(gclk));
	jdff dff_B_u6M0AzWb0_0(.din(w_dff_B_23I2t5e54_0),.dout(w_dff_B_u6M0AzWb0_0),.clk(gclk));
	jdff dff_B_OhpzQVtd6_0(.din(w_dff_B_u6M0AzWb0_0),.dout(w_dff_B_OhpzQVtd6_0),.clk(gclk));
	jdff dff_B_ghqpiIah2_0(.din(w_dff_B_OhpzQVtd6_0),.dout(w_dff_B_ghqpiIah2_0),.clk(gclk));
	jdff dff_B_5MmDMCKW7_0(.din(w_dff_B_ghqpiIah2_0),.dout(w_dff_B_5MmDMCKW7_0),.clk(gclk));
	jdff dff_B_tVWczIsZ9_0(.din(w_dff_B_5MmDMCKW7_0),.dout(w_dff_B_tVWczIsZ9_0),.clk(gclk));
	jdff dff_B_BjwpQMHQ1_0(.din(w_dff_B_tVWczIsZ9_0),.dout(w_dff_B_BjwpQMHQ1_0),.clk(gclk));
	jdff dff_B_ULDO8dqB2_0(.din(w_dff_B_BjwpQMHQ1_0),.dout(w_dff_B_ULDO8dqB2_0),.clk(gclk));
	jdff dff_B_QlrdZJQH0_0(.din(w_dff_B_ULDO8dqB2_0),.dout(w_dff_B_QlrdZJQH0_0),.clk(gclk));
	jdff dff_B_IsgJckqP0_0(.din(w_dff_B_QlrdZJQH0_0),.dout(w_dff_B_IsgJckqP0_0),.clk(gclk));
	jdff dff_B_eT6QaDVn0_0(.din(w_dff_B_IsgJckqP0_0),.dout(w_dff_B_eT6QaDVn0_0),.clk(gclk));
	jdff dff_B_t0U6Pf0O4_0(.din(w_dff_B_eT6QaDVn0_0),.dout(w_dff_B_t0U6Pf0O4_0),.clk(gclk));
	jdff dff_B_Dj7mkZ3I9_0(.din(w_dff_B_t0U6Pf0O4_0),.dout(w_dff_B_Dj7mkZ3I9_0),.clk(gclk));
	jdff dff_B_T1d6BPOm2_0(.din(w_dff_B_Dj7mkZ3I9_0),.dout(w_dff_B_T1d6BPOm2_0),.clk(gclk));
	jdff dff_B_7M1lrMPW2_1(.din(n790),.dout(w_dff_B_7M1lrMPW2_1),.clk(gclk));
	jdff dff_B_XoG7i2o52_1(.din(w_dff_B_7M1lrMPW2_1),.dout(w_dff_B_XoG7i2o52_1),.clk(gclk));
	jdff dff_B_3CM2afkW3_1(.din(w_dff_B_XoG7i2o52_1),.dout(w_dff_B_3CM2afkW3_1),.clk(gclk));
	jdff dff_B_5k0i0PCj5_1(.din(w_dff_B_3CM2afkW3_1),.dout(w_dff_B_5k0i0PCj5_1),.clk(gclk));
	jdff dff_B_1RSpuAkh5_1(.din(w_dff_B_5k0i0PCj5_1),.dout(w_dff_B_1RSpuAkh5_1),.clk(gclk));
	jdff dff_B_vAg6SD5U8_1(.din(w_dff_B_1RSpuAkh5_1),.dout(w_dff_B_vAg6SD5U8_1),.clk(gclk));
	jdff dff_B_uD668HLK9_1(.din(w_dff_B_vAg6SD5U8_1),.dout(w_dff_B_uD668HLK9_1),.clk(gclk));
	jdff dff_B_GZuxk9lo6_1(.din(w_dff_B_uD668HLK9_1),.dout(w_dff_B_GZuxk9lo6_1),.clk(gclk));
	jdff dff_B_maC7SitY5_1(.din(w_dff_B_GZuxk9lo6_1),.dout(w_dff_B_maC7SitY5_1),.clk(gclk));
	jdff dff_B_SvJAykEn0_1(.din(w_dff_B_maC7SitY5_1),.dout(w_dff_B_SvJAykEn0_1),.clk(gclk));
	jdff dff_B_WbhBj9pS6_1(.din(w_dff_B_SvJAykEn0_1),.dout(w_dff_B_WbhBj9pS6_1),.clk(gclk));
	jdff dff_B_wEDlNkBH6_1(.din(w_dff_B_WbhBj9pS6_1),.dout(w_dff_B_wEDlNkBH6_1),.clk(gclk));
	jdff dff_B_RNc4U37m0_1(.din(w_dff_B_wEDlNkBH6_1),.dout(w_dff_B_RNc4U37m0_1),.clk(gclk));
	jdff dff_B_brHvYuwj6_1(.din(w_dff_B_RNc4U37m0_1),.dout(w_dff_B_brHvYuwj6_1),.clk(gclk));
	jdff dff_B_u3oP7Dlo2_1(.din(w_dff_B_brHvYuwj6_1),.dout(w_dff_B_u3oP7Dlo2_1),.clk(gclk));
	jdff dff_B_6Us1o1PU5_1(.din(n794),.dout(w_dff_B_6Us1o1PU5_1),.clk(gclk));
	jdff dff_B_UA13COXH6_1(.din(w_dff_B_6Us1o1PU5_1),.dout(w_dff_B_UA13COXH6_1),.clk(gclk));
	jdff dff_B_BvbgFEcY5_1(.din(w_dff_B_UA13COXH6_1),.dout(w_dff_B_BvbgFEcY5_1),.clk(gclk));
	jdff dff_B_AlcbGVrj8_1(.din(w_dff_B_BvbgFEcY5_1),.dout(w_dff_B_AlcbGVrj8_1),.clk(gclk));
	jdff dff_B_vlmifdGp3_1(.din(w_dff_B_AlcbGVrj8_1),.dout(w_dff_B_vlmifdGp3_1),.clk(gclk));
	jdff dff_B_91Pq6RVV2_1(.din(w_dff_B_vlmifdGp3_1),.dout(w_dff_B_91Pq6RVV2_1),.clk(gclk));
	jdff dff_B_ifa296Kc3_1(.din(w_dff_B_91Pq6RVV2_1),.dout(w_dff_B_ifa296Kc3_1),.clk(gclk));
	jdff dff_B_V1hcwmJH1_1(.din(w_dff_B_ifa296Kc3_1),.dout(w_dff_B_V1hcwmJH1_1),.clk(gclk));
	jdff dff_B_Uqfl6Yaz1_1(.din(w_dff_B_V1hcwmJH1_1),.dout(w_dff_B_Uqfl6Yaz1_1),.clk(gclk));
	jdff dff_B_04WncmoK4_1(.din(w_dff_B_Uqfl6Yaz1_1),.dout(w_dff_B_04WncmoK4_1),.clk(gclk));
	jdff dff_B_qe1whFNV3_1(.din(w_dff_B_04WncmoK4_1),.dout(w_dff_B_qe1whFNV3_1),.clk(gclk));
	jdff dff_B_hRWrvexO9_1(.din(w_dff_B_qe1whFNV3_1),.dout(w_dff_B_hRWrvexO9_1),.clk(gclk));
	jdff dff_B_gKcrzpjS8_1(.din(w_dff_B_hRWrvexO9_1),.dout(w_dff_B_gKcrzpjS8_1),.clk(gclk));
	jdff dff_B_bWMxfGkw0_1(.din(w_dff_B_gKcrzpjS8_1),.dout(w_dff_B_bWMxfGkw0_1),.clk(gclk));
	jdff dff_B_NMFhvr9m9_1(.din(w_dff_B_bWMxfGkw0_1),.dout(w_dff_B_NMFhvr9m9_1),.clk(gclk));
	jdff dff_B_B2hLuiYn0_0(.din(n1036),.dout(w_dff_B_B2hLuiYn0_0),.clk(gclk));
	jdff dff_B_38oiTr2l5_0(.din(w_dff_B_B2hLuiYn0_0),.dout(w_dff_B_38oiTr2l5_0),.clk(gclk));
	jdff dff_B_uYbsBXlK2_0(.din(w_dff_B_38oiTr2l5_0),.dout(w_dff_B_uYbsBXlK2_0),.clk(gclk));
	jdff dff_B_Zjqf0u0m4_0(.din(w_dff_B_uYbsBXlK2_0),.dout(w_dff_B_Zjqf0u0m4_0),.clk(gclk));
	jdff dff_B_dyinEq376_0(.din(w_dff_B_Zjqf0u0m4_0),.dout(w_dff_B_dyinEq376_0),.clk(gclk));
	jdff dff_B_Wc4Ludv69_0(.din(w_dff_B_dyinEq376_0),.dout(w_dff_B_Wc4Ludv69_0),.clk(gclk));
	jdff dff_B_zWrP37Rb6_0(.din(w_dff_B_Wc4Ludv69_0),.dout(w_dff_B_zWrP37Rb6_0),.clk(gclk));
	jdff dff_B_JH8UfnCm6_0(.din(w_dff_B_zWrP37Rb6_0),.dout(w_dff_B_JH8UfnCm6_0),.clk(gclk));
	jdff dff_B_l9PVMqNj6_0(.din(w_dff_B_JH8UfnCm6_0),.dout(w_dff_B_l9PVMqNj6_0),.clk(gclk));
	jdff dff_B_v02053He5_0(.din(w_dff_B_l9PVMqNj6_0),.dout(w_dff_B_v02053He5_0),.clk(gclk));
	jdff dff_B_paAqqfnL4_0(.din(w_dff_B_v02053He5_0),.dout(w_dff_B_paAqqfnL4_0),.clk(gclk));
	jdff dff_B_QbAVlX530_0(.din(w_dff_B_paAqqfnL4_0),.dout(w_dff_B_QbAVlX530_0),.clk(gclk));
	jdff dff_B_9VwHz3EU6_0(.din(w_dff_B_QbAVlX530_0),.dout(w_dff_B_9VwHz3EU6_0),.clk(gclk));
	jdff dff_B_y53gdfjG8_0(.din(w_dff_B_9VwHz3EU6_0),.dout(w_dff_B_y53gdfjG8_0),.clk(gclk));
	jdff dff_B_7q9fuPJQ6_0(.din(w_dff_B_y53gdfjG8_0),.dout(w_dff_B_7q9fuPJQ6_0),.clk(gclk));
	jdff dff_B_9GcvIL8U1_0(.din(w_dff_B_7q9fuPJQ6_0),.dout(w_dff_B_9GcvIL8U1_0),.clk(gclk));
	jdff dff_B_Gw1dYDfT7_1(.din(n842),.dout(w_dff_B_Gw1dYDfT7_1),.clk(gclk));
	jdff dff_B_WKEClvuR0_1(.din(w_dff_B_Gw1dYDfT7_1),.dout(w_dff_B_WKEClvuR0_1),.clk(gclk));
	jdff dff_B_4Yixfr1f1_1(.din(w_dff_B_WKEClvuR0_1),.dout(w_dff_B_4Yixfr1f1_1),.clk(gclk));
	jdff dff_B_Tax8CM1w1_1(.din(w_dff_B_4Yixfr1f1_1),.dout(w_dff_B_Tax8CM1w1_1),.clk(gclk));
	jdff dff_B_phUmAw6k9_1(.din(w_dff_B_Tax8CM1w1_1),.dout(w_dff_B_phUmAw6k9_1),.clk(gclk));
	jdff dff_B_I5HoOQ6y8_1(.din(w_dff_B_phUmAw6k9_1),.dout(w_dff_B_I5HoOQ6y8_1),.clk(gclk));
	jdff dff_B_wcs81AfL4_1(.din(w_dff_B_I5HoOQ6y8_1),.dout(w_dff_B_wcs81AfL4_1),.clk(gclk));
	jdff dff_B_62W8pPqa8_1(.din(w_dff_B_wcs81AfL4_1),.dout(w_dff_B_62W8pPqa8_1),.clk(gclk));
	jdff dff_B_ZosEPnXn3_1(.din(w_dff_B_62W8pPqa8_1),.dout(w_dff_B_ZosEPnXn3_1),.clk(gclk));
	jdff dff_B_FiXAGPcI3_1(.din(w_dff_B_ZosEPnXn3_1),.dout(w_dff_B_FiXAGPcI3_1),.clk(gclk));
	jdff dff_B_ZTSxbjnP1_1(.din(w_dff_B_FiXAGPcI3_1),.dout(w_dff_B_ZTSxbjnP1_1),.clk(gclk));
	jdff dff_B_Bin7Hwuy9_1(.din(n843),.dout(w_dff_B_Bin7Hwuy9_1),.clk(gclk));
	jdff dff_B_PYjbCfre1_1(.din(w_dff_B_Bin7Hwuy9_1),.dout(w_dff_B_PYjbCfre1_1),.clk(gclk));
	jdff dff_B_UPvoHW9n9_1(.din(w_dff_B_PYjbCfre1_1),.dout(w_dff_B_UPvoHW9n9_1),.clk(gclk));
	jdff dff_B_UNZmtkoq5_1(.din(w_dff_B_UPvoHW9n9_1),.dout(w_dff_B_UNZmtkoq5_1),.clk(gclk));
	jdff dff_B_FF0x16jo9_1(.din(w_dff_B_UNZmtkoq5_1),.dout(w_dff_B_FF0x16jo9_1),.clk(gclk));
	jdff dff_B_UDiyE8Cg4_1(.din(w_dff_B_FF0x16jo9_1),.dout(w_dff_B_UDiyE8Cg4_1),.clk(gclk));
	jdff dff_B_wQJCt7bC5_1(.din(w_dff_B_UDiyE8Cg4_1),.dout(w_dff_B_wQJCt7bC5_1),.clk(gclk));
	jdff dff_B_EqioovOn5_1(.din(w_dff_B_wQJCt7bC5_1),.dout(w_dff_B_EqioovOn5_1),.clk(gclk));
	jdff dff_B_6PwXRHKg5_1(.din(w_dff_B_EqioovOn5_1),.dout(w_dff_B_6PwXRHKg5_1),.clk(gclk));
	jdff dff_B_tDZlnk9p1_1(.din(w_dff_B_6PwXRHKg5_1),.dout(w_dff_B_tDZlnk9p1_1),.clk(gclk));
	jdff dff_B_GV18tMPh4_1(.din(w_dff_B_tDZlnk9p1_1),.dout(w_dff_B_GV18tMPh4_1),.clk(gclk));
	jdff dff_B_h38f78Fw0_1(.din(w_dff_B_GV18tMPh4_1),.dout(w_dff_B_h38f78Fw0_1),.clk(gclk));
	jdff dff_B_VeT2Yyaa5_1(.din(w_dff_B_h38f78Fw0_1),.dout(w_dff_B_VeT2Yyaa5_1),.clk(gclk));
	jdff dff_B_A5DwHN7y8_0(.din(n1031),.dout(w_dff_B_A5DwHN7y8_0),.clk(gclk));
	jdff dff_B_gO0NL7DJ3_0(.din(w_dff_B_A5DwHN7y8_0),.dout(w_dff_B_gO0NL7DJ3_0),.clk(gclk));
	jdff dff_B_Gf7KTZyb2_0(.din(w_dff_B_gO0NL7DJ3_0),.dout(w_dff_B_Gf7KTZyb2_0),.clk(gclk));
	jdff dff_B_IJO2BKKF0_0(.din(w_dff_B_Gf7KTZyb2_0),.dout(w_dff_B_IJO2BKKF0_0),.clk(gclk));
	jdff dff_B_yFUpbVr59_0(.din(w_dff_B_IJO2BKKF0_0),.dout(w_dff_B_yFUpbVr59_0),.clk(gclk));
	jdff dff_B_UqU1vpSG3_0(.din(w_dff_B_yFUpbVr59_0),.dout(w_dff_B_UqU1vpSG3_0),.clk(gclk));
	jdff dff_B_3bY84fzm8_0(.din(w_dff_B_UqU1vpSG3_0),.dout(w_dff_B_3bY84fzm8_0),.clk(gclk));
	jdff dff_B_BNtIyLIC8_0(.din(w_dff_B_3bY84fzm8_0),.dout(w_dff_B_BNtIyLIC8_0),.clk(gclk));
	jdff dff_B_a6HOVMNp5_0(.din(w_dff_B_BNtIyLIC8_0),.dout(w_dff_B_a6HOVMNp5_0),.clk(gclk));
	jdff dff_B_VgNxVw340_0(.din(w_dff_B_a6HOVMNp5_0),.dout(w_dff_B_VgNxVw340_0),.clk(gclk));
	jdff dff_B_9dMiWYt69_0(.din(w_dff_B_VgNxVw340_0),.dout(w_dff_B_9dMiWYt69_0),.clk(gclk));
	jdff dff_B_QbEwMlUz9_0(.din(w_dff_B_9dMiWYt69_0),.dout(w_dff_B_QbEwMlUz9_0),.clk(gclk));
	jdff dff_B_CRsm53By6_0(.din(w_dff_B_QbEwMlUz9_0),.dout(w_dff_B_CRsm53By6_0),.clk(gclk));
	jdff dff_B_8loWY7PT9_0(.din(w_dff_B_CRsm53By6_0),.dout(w_dff_B_8loWY7PT9_0),.clk(gclk));
	jdff dff_B_JuK41xEe3_3(.din(n718),.dout(w_dff_B_JuK41xEe3_3),.clk(gclk));
	jdff dff_B_93SjQFsm5_3(.din(w_dff_B_JuK41xEe3_3),.dout(w_dff_B_93SjQFsm5_3),.clk(gclk));
	jdff dff_B_ie39DiEx3_3(.din(w_dff_B_93SjQFsm5_3),.dout(w_dff_B_ie39DiEx3_3),.clk(gclk));
	jdff dff_B_hpYgyyl18_3(.din(w_dff_B_ie39DiEx3_3),.dout(w_dff_B_hpYgyyl18_3),.clk(gclk));
	jdff dff_B_jMxuNleY0_3(.din(w_dff_B_hpYgyyl18_3),.dout(w_dff_B_jMxuNleY0_3),.clk(gclk));
	jdff dff_B_oXzYyErQ1_3(.din(w_dff_B_jMxuNleY0_3),.dout(w_dff_B_oXzYyErQ1_3),.clk(gclk));
	jdff dff_B_xX8YJHkx6_3(.din(w_dff_B_oXzYyErQ1_3),.dout(w_dff_B_xX8YJHkx6_3),.clk(gclk));
	jdff dff_B_utu1s2SQ7_3(.din(w_dff_B_xX8YJHkx6_3),.dout(w_dff_B_utu1s2SQ7_3),.clk(gclk));
	jdff dff_B_7JPvDrLT9_3(.din(w_dff_B_utu1s2SQ7_3),.dout(w_dff_B_7JPvDrLT9_3),.clk(gclk));
	jdff dff_B_CV1ibV4a3_3(.din(w_dff_B_7JPvDrLT9_3),.dout(w_dff_B_CV1ibV4a3_3),.clk(gclk));
	jdff dff_B_7UuL3FUV5_3(.din(w_dff_B_CV1ibV4a3_3),.dout(w_dff_B_7UuL3FUV5_3),.clk(gclk));
	jdff dff_B_FZ91vWJ72_3(.din(w_dff_B_7UuL3FUV5_3),.dout(w_dff_B_FZ91vWJ72_3),.clk(gclk));
	jdff dff_B_hh9fC2uG3_3(.din(w_dff_B_FZ91vWJ72_3),.dout(w_dff_B_hh9fC2uG3_3),.clk(gclk));
	jdff dff_B_60DsptNY9_3(.din(w_dff_B_hh9fC2uG3_3),.dout(w_dff_B_60DsptNY9_3),.clk(gclk));
	jdff dff_B_BRdw5yBj8_3(.din(w_dff_B_60DsptNY9_3),.dout(w_dff_B_BRdw5yBj8_3),.clk(gclk));
	jdff dff_B_zeJQSlSZ3_3(.din(w_dff_B_BRdw5yBj8_3),.dout(w_dff_B_zeJQSlSZ3_3),.clk(gclk));
	jdff dff_B_IdW8oNTG6_3(.din(w_dff_B_zeJQSlSZ3_3),.dout(w_dff_B_IdW8oNTG6_3),.clk(gclk));
	jdff dff_B_QyolK1dE4_3(.din(w_dff_B_IdW8oNTG6_3),.dout(w_dff_B_QyolK1dE4_3),.clk(gclk));
	jdff dff_B_Efdvrtbe2_3(.din(w_dff_B_QyolK1dE4_3),.dout(w_dff_B_Efdvrtbe2_3),.clk(gclk));
	jdff dff_B_MSPwtXEF2_3(.din(w_dff_B_Efdvrtbe2_3),.dout(w_dff_B_MSPwtXEF2_3),.clk(gclk));
	jdff dff_B_u7PRntmF6_3(.din(w_dff_B_MSPwtXEF2_3),.dout(w_dff_B_u7PRntmF6_3),.clk(gclk));
	jdff dff_B_bMaMMfOB6_3(.din(w_dff_B_u7PRntmF6_3),.dout(w_dff_B_bMaMMfOB6_3),.clk(gclk));
	jdff dff_B_NcsPgPvU4_3(.din(w_dff_B_bMaMMfOB6_3),.dout(w_dff_B_NcsPgPvU4_3),.clk(gclk));
	jdff dff_B_4D5BXUHe7_3(.din(w_dff_B_NcsPgPvU4_3),.dout(w_dff_B_4D5BXUHe7_3),.clk(gclk));
	jdff dff_B_HzBoAF1D8_1(.din(n1305),.dout(w_dff_B_HzBoAF1D8_1),.clk(gclk));
	jdff dff_B_tVLtNIMF4_1(.din(w_dff_B_HzBoAF1D8_1),.dout(w_dff_B_tVLtNIMF4_1),.clk(gclk));
	jdff dff_B_GuxoXpB74_1(.din(w_dff_B_tVLtNIMF4_1),.dout(w_dff_B_GuxoXpB74_1),.clk(gclk));
	jdff dff_B_DTjEKTEt3_1(.din(w_dff_B_GuxoXpB74_1),.dout(w_dff_B_DTjEKTEt3_1),.clk(gclk));
	jdff dff_B_rbx1awGU1_1(.din(w_dff_B_DTjEKTEt3_1),.dout(w_dff_B_rbx1awGU1_1),.clk(gclk));
	jdff dff_B_OY0MOmnh6_1(.din(w_dff_B_rbx1awGU1_1),.dout(w_dff_B_OY0MOmnh6_1),.clk(gclk));
	jdff dff_B_irR47WqU3_1(.din(w_dff_B_OY0MOmnh6_1),.dout(w_dff_B_irR47WqU3_1),.clk(gclk));
	jdff dff_B_SG1bO3fH1_1(.din(w_dff_B_irR47WqU3_1),.dout(w_dff_B_SG1bO3fH1_1),.clk(gclk));
	jdff dff_B_pJBwPVHu5_1(.din(w_dff_B_SG1bO3fH1_1),.dout(w_dff_B_pJBwPVHu5_1),.clk(gclk));
	jdff dff_B_DBJ1bMFB5_1(.din(w_dff_B_pJBwPVHu5_1),.dout(w_dff_B_DBJ1bMFB5_1),.clk(gclk));
	jdff dff_B_evg1RF3N0_1(.din(w_dff_B_DBJ1bMFB5_1),.dout(w_dff_B_evg1RF3N0_1),.clk(gclk));
	jdff dff_B_7RYcBoPU1_1(.din(w_dff_B_evg1RF3N0_1),.dout(w_dff_B_7RYcBoPU1_1),.clk(gclk));
	jdff dff_B_zXpsqUdH6_1(.din(w_dff_B_7RYcBoPU1_1),.dout(w_dff_B_zXpsqUdH6_1),.clk(gclk));
	jdff dff_B_Zob7ArHT6_1(.din(w_dff_B_zXpsqUdH6_1),.dout(w_dff_B_Zob7ArHT6_1),.clk(gclk));
	jdff dff_B_wc2eYW0k9_1(.din(w_dff_B_Zob7ArHT6_1),.dout(w_dff_B_wc2eYW0k9_1),.clk(gclk));
	jdff dff_B_hXe5Qo5m7_1(.din(w_dff_B_wc2eYW0k9_1),.dout(w_dff_B_hXe5Qo5m7_1),.clk(gclk));
	jdff dff_B_3xjDdytG7_1(.din(w_dff_B_hXe5Qo5m7_1),.dout(w_dff_B_3xjDdytG7_1),.clk(gclk));
	jdff dff_B_eNvZU7tn2_1(.din(w_dff_B_3xjDdytG7_1),.dout(w_dff_B_eNvZU7tn2_1),.clk(gclk));
	jdff dff_B_fHdbwiZG9_1(.din(w_dff_B_eNvZU7tn2_1),.dout(w_dff_B_fHdbwiZG9_1),.clk(gclk));
	jdff dff_B_UnqY7FVK3_1(.din(w_dff_B_fHdbwiZG9_1),.dout(w_dff_B_UnqY7FVK3_1),.clk(gclk));
	jdff dff_B_UZf5VXFx7_1(.din(w_dff_B_UnqY7FVK3_1),.dout(w_dff_B_UZf5VXFx7_1),.clk(gclk));
	jdff dff_B_MmUI7ZMm7_1(.din(w_dff_B_UZf5VXFx7_1),.dout(w_dff_B_MmUI7ZMm7_1),.clk(gclk));
	jdff dff_B_uZ192TCG0_1(.din(n1347),.dout(w_dff_B_uZ192TCG0_1),.clk(gclk));
	jdff dff_B_WDf4wCSn8_1(.din(w_dff_B_uZ192TCG0_1),.dout(w_dff_B_WDf4wCSn8_1),.clk(gclk));
	jdff dff_B_RznskHIj2_1(.din(n1368),.dout(w_dff_B_RznskHIj2_1),.clk(gclk));
	jdff dff_B_Q5HzTztO4_1(.din(w_dff_B_RznskHIj2_1),.dout(w_dff_B_Q5HzTztO4_1),.clk(gclk));
	jdff dff_B_goT78SRU6_1(.din(w_dff_B_Q5HzTztO4_1),.dout(w_dff_B_goT78SRU6_1),.clk(gclk));
	jdff dff_B_WC0X31Ys1_1(.din(w_dff_B_goT78SRU6_1),.dout(w_dff_B_WC0X31Ys1_1),.clk(gclk));
	jdff dff_B_rM25Xr037_1(.din(w_dff_B_WC0X31Ys1_1),.dout(w_dff_B_rM25Xr037_1),.clk(gclk));
	jdff dff_B_nd1DUFUd8_1(.din(w_dff_B_rM25Xr037_1),.dout(w_dff_B_nd1DUFUd8_1),.clk(gclk));
	jdff dff_B_cU5aMtv53_1(.din(w_dff_B_nd1DUFUd8_1),.dout(w_dff_B_cU5aMtv53_1),.clk(gclk));
	jdff dff_B_rDIOLzwH7_1(.din(w_dff_B_cU5aMtv53_1),.dout(w_dff_B_rDIOLzwH7_1),.clk(gclk));
	jdff dff_B_ynMNMAMO9_1(.din(w_dff_B_rDIOLzwH7_1),.dout(w_dff_B_ynMNMAMO9_1),.clk(gclk));
	jdff dff_B_uozBSSLV5_1(.din(w_dff_B_ynMNMAMO9_1),.dout(w_dff_B_uozBSSLV5_1),.clk(gclk));
	jdff dff_B_uaVUETXI5_1(.din(w_dff_B_uozBSSLV5_1),.dout(w_dff_B_uaVUETXI5_1),.clk(gclk));
	jdff dff_B_qaGvqW4J3_1(.din(w_dff_B_uaVUETXI5_1),.dout(w_dff_B_qaGvqW4J3_1),.clk(gclk));
	jdff dff_B_sCoF3rCx2_1(.din(w_dff_B_qaGvqW4J3_1),.dout(w_dff_B_sCoF3rCx2_1),.clk(gclk));
	jdff dff_B_sqslCrcV6_1(.din(w_dff_B_sCoF3rCx2_1),.dout(w_dff_B_sqslCrcV6_1),.clk(gclk));
	jdff dff_B_A7GEn0iK2_1(.din(w_dff_B_sqslCrcV6_1),.dout(w_dff_B_A7GEn0iK2_1),.clk(gclk));
	jdff dff_B_i4FjaiwR6_1(.din(w_dff_B_A7GEn0iK2_1),.dout(w_dff_B_i4FjaiwR6_1),.clk(gclk));
	jdff dff_B_uWiypTGG0_1(.din(w_dff_B_i4FjaiwR6_1),.dout(w_dff_B_uWiypTGG0_1),.clk(gclk));
	jdff dff_B_4tcwl7ig6_1(.din(w_dff_B_uWiypTGG0_1),.dout(w_dff_B_4tcwl7ig6_1),.clk(gclk));
	jdff dff_B_opKgIT7H5_1(.din(w_dff_B_4tcwl7ig6_1),.dout(w_dff_B_opKgIT7H5_1),.clk(gclk));
	jdff dff_B_TKf0P0eY2_1(.din(w_dff_B_opKgIT7H5_1),.dout(w_dff_B_TKf0P0eY2_1),.clk(gclk));
	jdff dff_B_NiEoq66h7_1(.din(w_dff_B_TKf0P0eY2_1),.dout(w_dff_B_NiEoq66h7_1),.clk(gclk));
	jdff dff_B_JyJ9ZyIc9_1(.din(w_dff_B_NiEoq66h7_1),.dout(w_dff_B_JyJ9ZyIc9_1),.clk(gclk));
	jdff dff_B_le3aFNwW9_1(.din(w_dff_B_JyJ9ZyIc9_1),.dout(w_dff_B_le3aFNwW9_1),.clk(gclk));
	jdff dff_B_yUTq1RZm8_1(.din(w_dff_B_le3aFNwW9_1),.dout(w_dff_B_yUTq1RZm8_1),.clk(gclk));
	jdff dff_B_iV9Ty4gF7_1(.din(w_dff_B_yUTq1RZm8_1),.dout(w_dff_B_iV9Ty4gF7_1),.clk(gclk));
	jdff dff_B_bhGoLnJM2_1(.din(w_dff_B_iV9Ty4gF7_1),.dout(w_dff_B_bhGoLnJM2_1),.clk(gclk));
	jdff dff_B_XB3WTDsk3_1(.din(w_dff_B_bhGoLnJM2_1),.dout(w_dff_B_XB3WTDsk3_1),.clk(gclk));
	jdff dff_B_SFv6DJjw4_1(.din(w_dff_B_XB3WTDsk3_1),.dout(w_dff_B_SFv6DJjw4_1),.clk(gclk));
	jdff dff_B_e6bgyifi9_1(.din(w_dff_B_SFv6DJjw4_1),.dout(w_dff_B_e6bgyifi9_1),.clk(gclk));
	jdff dff_B_fkChAObi7_1(.din(w_dff_B_e6bgyifi9_1),.dout(w_dff_B_fkChAObi7_1),.clk(gclk));
	jdff dff_B_3eFE7fLM2_1(.din(w_dff_B_fkChAObi7_1),.dout(w_dff_B_3eFE7fLM2_1),.clk(gclk));
	jdff dff_B_LLmxIlqS9_1(.din(w_dff_B_3eFE7fLM2_1),.dout(w_dff_B_LLmxIlqS9_1),.clk(gclk));
	jdff dff_B_IOPm2ZGa5_1(.din(w_dff_B_LLmxIlqS9_1),.dout(w_dff_B_IOPm2ZGa5_1),.clk(gclk));
	jdff dff_B_zz5BSZhW8_1(.din(n1377),.dout(w_dff_B_zz5BSZhW8_1),.clk(gclk));
	jdff dff_B_39kMFezJ5_1(.din(w_dff_B_zz5BSZhW8_1),.dout(w_dff_B_39kMFezJ5_1),.clk(gclk));
	jdff dff_B_q6WIcda37_1(.din(n1378),.dout(w_dff_B_q6WIcda37_1),.clk(gclk));
	jdff dff_B_lNrZNO0Q0_1(.din(w_dff_B_q6WIcda37_1),.dout(w_dff_B_lNrZNO0Q0_1),.clk(gclk));
	jdff dff_B_Z0sU4nZ85_1(.din(w_dff_B_lNrZNO0Q0_1),.dout(w_dff_B_Z0sU4nZ85_1),.clk(gclk));
	jdff dff_B_SBI04YPO6_1(.din(w_dff_B_Z0sU4nZ85_1),.dout(w_dff_B_SBI04YPO6_1),.clk(gclk));
	jdff dff_B_rUoPHGzb6_1(.din(w_dff_B_SBI04YPO6_1),.dout(w_dff_B_rUoPHGzb6_1),.clk(gclk));
	jdff dff_B_qKGOuUOs9_1(.din(w_dff_B_rUoPHGzb6_1),.dout(w_dff_B_qKGOuUOs9_1),.clk(gclk));
	jdff dff_B_x4CrNFNp6_1(.din(w_dff_B_qKGOuUOs9_1),.dout(w_dff_B_x4CrNFNp6_1),.clk(gclk));
	jdff dff_B_avQhiC6t0_1(.din(w_dff_B_x4CrNFNp6_1),.dout(w_dff_B_avQhiC6t0_1),.clk(gclk));
	jdff dff_B_7GMzqdeq9_0(.din(n1379),.dout(w_dff_B_7GMzqdeq9_0),.clk(gclk));
	jdff dff_B_uRYSEkUI5_0(.din(w_dff_B_7GMzqdeq9_0),.dout(w_dff_B_uRYSEkUI5_0),.clk(gclk));
	jdff dff_B_bDaFGUFH9_0(.din(w_dff_B_uRYSEkUI5_0),.dout(w_dff_B_bDaFGUFH9_0),.clk(gclk));
	jdff dff_B_juw7xejP3_0(.din(w_dff_B_bDaFGUFH9_0),.dout(w_dff_B_juw7xejP3_0),.clk(gclk));
	jdff dff_B_BRxNbwkm8_0(.din(w_dff_B_juw7xejP3_0),.dout(w_dff_B_BRxNbwkm8_0),.clk(gclk));
	jdff dff_B_agVygko66_0(.din(w_dff_B_BRxNbwkm8_0),.dout(w_dff_B_agVygko66_0),.clk(gclk));
	jdff dff_B_RIw1Ilxk0_0(.din(w_dff_B_agVygko66_0),.dout(w_dff_B_RIw1Ilxk0_0),.clk(gclk));
	jdff dff_A_76k9SREw6_0(.dout(w_G414_0),.din(w_dff_A_76k9SREw6_0),.clk(gclk));
	jdff dff_B_pbqrQltl6_3(.din(n715),.dout(w_dff_B_pbqrQltl6_3),.clk(gclk));
	jdff dff_B_PUqrvXMC6_3(.din(w_dff_B_pbqrQltl6_3),.dout(w_dff_B_PUqrvXMC6_3),.clk(gclk));
	jdff dff_B_K7hFgk7U8_3(.din(w_dff_B_PUqrvXMC6_3),.dout(w_dff_B_K7hFgk7U8_3),.clk(gclk));
	jdff dff_B_svD7A4pO2_3(.din(w_dff_B_K7hFgk7U8_3),.dout(w_dff_B_svD7A4pO2_3),.clk(gclk));
	jdff dff_B_8xOSwhQ07_3(.din(w_dff_B_svD7A4pO2_3),.dout(w_dff_B_8xOSwhQ07_3),.clk(gclk));
	jdff dff_B_nCKFztNW0_3(.din(w_dff_B_8xOSwhQ07_3),.dout(w_dff_B_nCKFztNW0_3),.clk(gclk));
	jdff dff_B_biXxT3gb4_3(.din(w_dff_B_nCKFztNW0_3),.dout(w_dff_B_biXxT3gb4_3),.clk(gclk));
	jdff dff_B_dbVi2Z9V8_3(.din(w_dff_B_biXxT3gb4_3),.dout(w_dff_B_dbVi2Z9V8_3),.clk(gclk));
	jdff dff_B_1zBBAgAi3_3(.din(w_dff_B_dbVi2Z9V8_3),.dout(w_dff_B_1zBBAgAi3_3),.clk(gclk));
	jdff dff_B_39clW5ga6_3(.din(w_dff_B_1zBBAgAi3_3),.dout(w_dff_B_39clW5ga6_3),.clk(gclk));
	jdff dff_B_ZkwrlPoR3_3(.din(w_dff_B_39clW5ga6_3),.dout(w_dff_B_ZkwrlPoR3_3),.clk(gclk));
	jdff dff_B_NkFpvgDM0_3(.din(w_dff_B_ZkwrlPoR3_3),.dout(w_dff_B_NkFpvgDM0_3),.clk(gclk));
	jdff dff_B_jpeCzUAy0_3(.din(w_dff_B_NkFpvgDM0_3),.dout(w_dff_B_jpeCzUAy0_3),.clk(gclk));
	jdff dff_B_MnmvRxqQ5_3(.din(w_dff_B_jpeCzUAy0_3),.dout(w_dff_B_MnmvRxqQ5_3),.clk(gclk));
	jdff dff_B_DgBTPy9R6_3(.din(w_dff_B_MnmvRxqQ5_3),.dout(w_dff_B_DgBTPy9R6_3),.clk(gclk));
	jdff dff_B_mRi94PP12_3(.din(w_dff_B_DgBTPy9R6_3),.dout(w_dff_B_mRi94PP12_3),.clk(gclk));
	jdff dff_B_QGxmCFnk2_3(.din(w_dff_B_mRi94PP12_3),.dout(w_dff_B_QGxmCFnk2_3),.clk(gclk));
	jdff dff_B_PDPdz2Yp4_3(.din(w_dff_B_QGxmCFnk2_3),.dout(w_dff_B_PDPdz2Yp4_3),.clk(gclk));
	jdff dff_B_aLRc7sFK3_3(.din(w_dff_B_PDPdz2Yp4_3),.dout(w_dff_B_aLRc7sFK3_3),.clk(gclk));
	jdff dff_B_hOhvEjaL4_3(.din(w_dff_B_aLRc7sFK3_3),.dout(w_dff_B_hOhvEjaL4_3),.clk(gclk));
	jdff dff_B_9w6MseZu9_3(.din(w_dff_B_hOhvEjaL4_3),.dout(w_dff_B_9w6MseZu9_3),.clk(gclk));
	jdff dff_B_2xFQEemQ3_3(.din(w_dff_B_9w6MseZu9_3),.dout(w_dff_B_2xFQEemQ3_3),.clk(gclk));
	jdff dff_B_YRuhaPUY8_3(.din(w_dff_B_2xFQEemQ3_3),.dout(w_dff_B_YRuhaPUY8_3),.clk(gclk));
	jdff dff_B_tXSifjvS6_3(.din(w_dff_B_YRuhaPUY8_3),.dout(w_dff_B_tXSifjvS6_3),.clk(gclk));
	jdff dff_B_T6SfYfZx3_3(.din(w_dff_B_tXSifjvS6_3),.dout(w_dff_B_T6SfYfZx3_3),.clk(gclk));
	jdff dff_B_S6FG1Isd3_3(.din(w_dff_B_T6SfYfZx3_3),.dout(w_dff_B_S6FG1Isd3_3),.clk(gclk));
	jdff dff_B_fv6XoOr35_3(.din(w_dff_B_S6FG1Isd3_3),.dout(w_dff_B_fv6XoOr35_3),.clk(gclk));
	jdff dff_B_Ary4ZO6f5_3(.din(w_dff_B_fv6XoOr35_3),.dout(w_dff_B_Ary4ZO6f5_3),.clk(gclk));
	jdff dff_B_4LS7fqyE8_3(.din(w_dff_B_Ary4ZO6f5_3),.dout(w_dff_B_4LS7fqyE8_3),.clk(gclk));
	jdff dff_B_dC65g0Go1_3(.din(w_dff_B_4LS7fqyE8_3),.dout(w_dff_B_dC65g0Go1_3),.clk(gclk));
	jdff dff_B_VVFFn8WV7_3(.din(w_dff_B_dC65g0Go1_3),.dout(w_dff_B_VVFFn8WV7_3),.clk(gclk));
	jdff dff_B_loIHxii74_3(.din(w_dff_B_VVFFn8WV7_3),.dout(w_dff_B_loIHxii74_3),.clk(gclk));
	jdff dff_B_p6HvR6vZ2_3(.din(w_dff_B_loIHxii74_3),.dout(w_dff_B_p6HvR6vZ2_3),.clk(gclk));
	jdff dff_B_p1zgFYqg9_3(.din(w_dff_B_p6HvR6vZ2_3),.dout(w_dff_B_p1zgFYqg9_3),.clk(gclk));
	jdff dff_B_7xfDQCrw4_0(.din(n1478),.dout(w_dff_B_7xfDQCrw4_0),.clk(gclk));
	jdff dff_B_wJPTGXyJ2_0(.din(w_dff_B_7xfDQCrw4_0),.dout(w_dff_B_wJPTGXyJ2_0),.clk(gclk));
	jdff dff_B_Ecfi3mhT0_0(.din(n1526),.dout(w_dff_B_Ecfi3mhT0_0),.clk(gclk));
	jdff dff_B_ilTnKteO2_1(.din(n1551),.dout(w_dff_B_ilTnKteO2_1),.clk(gclk));
	jdff dff_A_Dmc7a2bN2_1(.dout(w_dff_A_LLNBvJTM8_0),.din(w_dff_A_Dmc7a2bN2_1),.clk(gclk));
	jdff dff_A_LLNBvJTM8_0(.dout(w_dff_A_GEvlkdsB5_0),.din(w_dff_A_LLNBvJTM8_0),.clk(gclk));
	jdff dff_A_GEvlkdsB5_0(.dout(w_dff_A_YaYzmZlX2_0),.din(w_dff_A_GEvlkdsB5_0),.clk(gclk));
	jdff dff_A_YaYzmZlX2_0(.dout(w_dff_A_FX0Iisaz5_0),.din(w_dff_A_YaYzmZlX2_0),.clk(gclk));
	jdff dff_A_FX0Iisaz5_0(.dout(w_dff_A_MIhcir4I6_0),.din(w_dff_A_FX0Iisaz5_0),.clk(gclk));
	jdff dff_A_MIhcir4I6_0(.dout(w_dff_A_erFnwnth9_0),.din(w_dff_A_MIhcir4I6_0),.clk(gclk));
	jdff dff_A_erFnwnth9_0(.dout(w_dff_A_bQzyhJSN6_0),.din(w_dff_A_erFnwnth9_0),.clk(gclk));
	jdff dff_A_bQzyhJSN6_0(.dout(w_dff_A_wLqUgbMr3_0),.din(w_dff_A_bQzyhJSN6_0),.clk(gclk));
	jdff dff_A_wLqUgbMr3_0(.dout(w_dff_A_uWI17KVJ3_0),.din(w_dff_A_wLqUgbMr3_0),.clk(gclk));
	jdff dff_A_uWI17KVJ3_0(.dout(w_dff_A_VB5iWxWM3_0),.din(w_dff_A_uWI17KVJ3_0),.clk(gclk));
	jdff dff_A_VB5iWxWM3_0(.dout(w_dff_A_zhbhsqta1_0),.din(w_dff_A_VB5iWxWM3_0),.clk(gclk));
	jdff dff_A_zhbhsqta1_0(.dout(w_dff_A_gMEzPjoT8_0),.din(w_dff_A_zhbhsqta1_0),.clk(gclk));
	jdff dff_A_gMEzPjoT8_0(.dout(w_dff_A_oAJOi9300_0),.din(w_dff_A_gMEzPjoT8_0),.clk(gclk));
	jdff dff_A_oAJOi9300_0(.dout(w_dff_A_FsicpojQ8_0),.din(w_dff_A_oAJOi9300_0),.clk(gclk));
	jdff dff_A_FsicpojQ8_0(.dout(w_dff_A_mshP6Gmr6_0),.din(w_dff_A_FsicpojQ8_0),.clk(gclk));
	jdff dff_A_mshP6Gmr6_0(.dout(w_dff_A_9ZwfPTf05_0),.din(w_dff_A_mshP6Gmr6_0),.clk(gclk));
	jdff dff_A_9ZwfPTf05_0(.dout(w_dff_A_N33t5uUQ4_0),.din(w_dff_A_9ZwfPTf05_0),.clk(gclk));
	jdff dff_A_N33t5uUQ4_0(.dout(w_dff_A_EbUD35wF7_0),.din(w_dff_A_N33t5uUQ4_0),.clk(gclk));
	jdff dff_A_EbUD35wF7_0(.dout(w_dff_A_E3m7ZjeC2_0),.din(w_dff_A_EbUD35wF7_0),.clk(gclk));
	jdff dff_A_E3m7ZjeC2_0(.dout(w_dff_A_zVnf6q9a8_0),.din(w_dff_A_E3m7ZjeC2_0),.clk(gclk));
	jdff dff_A_zVnf6q9a8_0(.dout(w_dff_A_Nq5hrONx9_0),.din(w_dff_A_zVnf6q9a8_0),.clk(gclk));
	jdff dff_A_Nq5hrONx9_0(.dout(w_dff_A_YqpFphdb8_0),.din(w_dff_A_Nq5hrONx9_0),.clk(gclk));
	jdff dff_A_YqpFphdb8_0(.dout(w_dff_A_S5BJmosr8_0),.din(w_dff_A_YqpFphdb8_0),.clk(gclk));
	jdff dff_A_S5BJmosr8_0(.dout(w_dff_A_71RZnxKQ3_0),.din(w_dff_A_S5BJmosr8_0),.clk(gclk));
	jdff dff_A_71RZnxKQ3_0(.dout(w_dff_A_6yMSafOb1_0),.din(w_dff_A_71RZnxKQ3_0),.clk(gclk));
	jdff dff_A_6yMSafOb1_0(.dout(w_dff_A_jj6JeSgk7_0),.din(w_dff_A_6yMSafOb1_0),.clk(gclk));
	jdff dff_A_jj6JeSgk7_0(.dout(w_dff_A_rGkCTCdA5_0),.din(w_dff_A_jj6JeSgk7_0),.clk(gclk));
	jdff dff_A_rGkCTCdA5_0(.dout(w_dff_A_hvCgOQpC5_0),.din(w_dff_A_rGkCTCdA5_0),.clk(gclk));
	jdff dff_A_hvCgOQpC5_0(.dout(w_dff_A_w7hDUjCD5_0),.din(w_dff_A_hvCgOQpC5_0),.clk(gclk));
	jdff dff_A_w7hDUjCD5_0(.dout(w_dff_A_TFlXIh2G6_0),.din(w_dff_A_w7hDUjCD5_0),.clk(gclk));
	jdff dff_A_TFlXIh2G6_0(.dout(w_dff_A_1n6ENcOU8_0),.din(w_dff_A_TFlXIh2G6_0),.clk(gclk));
	jdff dff_A_1n6ENcOU8_0(.dout(w_dff_A_6vJCtxEh0_0),.din(w_dff_A_1n6ENcOU8_0),.clk(gclk));
	jdff dff_A_6vJCtxEh0_0(.dout(w_dff_A_AUQvMz4w4_0),.din(w_dff_A_6vJCtxEh0_0),.clk(gclk));
	jdff dff_A_AUQvMz4w4_0(.dout(w_dff_A_ulmky10N1_0),.din(w_dff_A_AUQvMz4w4_0),.clk(gclk));
	jdff dff_A_ulmky10N1_0(.dout(w_dff_A_swuztbhy0_0),.din(w_dff_A_ulmky10N1_0),.clk(gclk));
	jdff dff_A_swuztbhy0_0(.dout(w_dff_A_v8D77aif1_0),.din(w_dff_A_swuztbhy0_0),.clk(gclk));
	jdff dff_A_v8D77aif1_0(.dout(w_dff_A_MzjyoJYC7_0),.din(w_dff_A_v8D77aif1_0),.clk(gclk));
	jdff dff_A_MzjyoJYC7_0(.dout(w_dff_A_LWM8mLPO1_0),.din(w_dff_A_MzjyoJYC7_0),.clk(gclk));
	jdff dff_A_LWM8mLPO1_0(.dout(G2),.din(w_dff_A_LWM8mLPO1_0),.clk(gclk));
	jdff dff_A_6v1KheBj0_1(.dout(w_dff_A_YY0xL0rk4_0),.din(w_dff_A_6v1KheBj0_1),.clk(gclk));
	jdff dff_A_YY0xL0rk4_0(.dout(w_dff_A_3bF7dwZG0_0),.din(w_dff_A_YY0xL0rk4_0),.clk(gclk));
	jdff dff_A_3bF7dwZG0_0(.dout(w_dff_A_35PC5vQ83_0),.din(w_dff_A_3bF7dwZG0_0),.clk(gclk));
	jdff dff_A_35PC5vQ83_0(.dout(w_dff_A_AJHmpnhH7_0),.din(w_dff_A_35PC5vQ83_0),.clk(gclk));
	jdff dff_A_AJHmpnhH7_0(.dout(w_dff_A_CMwCjjRI2_0),.din(w_dff_A_AJHmpnhH7_0),.clk(gclk));
	jdff dff_A_CMwCjjRI2_0(.dout(w_dff_A_hqt01n107_0),.din(w_dff_A_CMwCjjRI2_0),.clk(gclk));
	jdff dff_A_hqt01n107_0(.dout(w_dff_A_CnzwQmx13_0),.din(w_dff_A_hqt01n107_0),.clk(gclk));
	jdff dff_A_CnzwQmx13_0(.dout(w_dff_A_GN2WozW12_0),.din(w_dff_A_CnzwQmx13_0),.clk(gclk));
	jdff dff_A_GN2WozW12_0(.dout(w_dff_A_sV4syeeH4_0),.din(w_dff_A_GN2WozW12_0),.clk(gclk));
	jdff dff_A_sV4syeeH4_0(.dout(w_dff_A_jVx5KnoL8_0),.din(w_dff_A_sV4syeeH4_0),.clk(gclk));
	jdff dff_A_jVx5KnoL8_0(.dout(w_dff_A_hCZEAIKm2_0),.din(w_dff_A_jVx5KnoL8_0),.clk(gclk));
	jdff dff_A_hCZEAIKm2_0(.dout(w_dff_A_ozKRS0Sp4_0),.din(w_dff_A_hCZEAIKm2_0),.clk(gclk));
	jdff dff_A_ozKRS0Sp4_0(.dout(w_dff_A_QMaNV75Q3_0),.din(w_dff_A_ozKRS0Sp4_0),.clk(gclk));
	jdff dff_A_QMaNV75Q3_0(.dout(w_dff_A_CqEIMk7e3_0),.din(w_dff_A_QMaNV75Q3_0),.clk(gclk));
	jdff dff_A_CqEIMk7e3_0(.dout(w_dff_A_9L2Rqvdx2_0),.din(w_dff_A_CqEIMk7e3_0),.clk(gclk));
	jdff dff_A_9L2Rqvdx2_0(.dout(w_dff_A_XDt8ZnXd2_0),.din(w_dff_A_9L2Rqvdx2_0),.clk(gclk));
	jdff dff_A_XDt8ZnXd2_0(.dout(w_dff_A_MsXBp7Fd5_0),.din(w_dff_A_XDt8ZnXd2_0),.clk(gclk));
	jdff dff_A_MsXBp7Fd5_0(.dout(w_dff_A_Y12zr4vQ4_0),.din(w_dff_A_MsXBp7Fd5_0),.clk(gclk));
	jdff dff_A_Y12zr4vQ4_0(.dout(w_dff_A_YuVSPCiI7_0),.din(w_dff_A_Y12zr4vQ4_0),.clk(gclk));
	jdff dff_A_YuVSPCiI7_0(.dout(w_dff_A_QTDWwmDk3_0),.din(w_dff_A_YuVSPCiI7_0),.clk(gclk));
	jdff dff_A_QTDWwmDk3_0(.dout(w_dff_A_6IZ5LgYS4_0),.din(w_dff_A_QTDWwmDk3_0),.clk(gclk));
	jdff dff_A_6IZ5LgYS4_0(.dout(w_dff_A_8oR3DoJm0_0),.din(w_dff_A_6IZ5LgYS4_0),.clk(gclk));
	jdff dff_A_8oR3DoJm0_0(.dout(w_dff_A_Nbl5VoIt6_0),.din(w_dff_A_8oR3DoJm0_0),.clk(gclk));
	jdff dff_A_Nbl5VoIt6_0(.dout(w_dff_A_UY9cMqF68_0),.din(w_dff_A_Nbl5VoIt6_0),.clk(gclk));
	jdff dff_A_UY9cMqF68_0(.dout(w_dff_A_ybP7apAr7_0),.din(w_dff_A_UY9cMqF68_0),.clk(gclk));
	jdff dff_A_ybP7apAr7_0(.dout(w_dff_A_ovUm93dE4_0),.din(w_dff_A_ybP7apAr7_0),.clk(gclk));
	jdff dff_A_ovUm93dE4_0(.dout(w_dff_A_aayRUxMn9_0),.din(w_dff_A_ovUm93dE4_0),.clk(gclk));
	jdff dff_A_aayRUxMn9_0(.dout(w_dff_A_TzFmMYuV7_0),.din(w_dff_A_aayRUxMn9_0),.clk(gclk));
	jdff dff_A_TzFmMYuV7_0(.dout(w_dff_A_yMHO25it0_0),.din(w_dff_A_TzFmMYuV7_0),.clk(gclk));
	jdff dff_A_yMHO25it0_0(.dout(w_dff_A_ED4QewEl8_0),.din(w_dff_A_yMHO25it0_0),.clk(gclk));
	jdff dff_A_ED4QewEl8_0(.dout(w_dff_A_yCudmDL28_0),.din(w_dff_A_ED4QewEl8_0),.clk(gclk));
	jdff dff_A_yCudmDL28_0(.dout(w_dff_A_MOmaS9wo9_0),.din(w_dff_A_yCudmDL28_0),.clk(gclk));
	jdff dff_A_MOmaS9wo9_0(.dout(w_dff_A_ZrhELOdn8_0),.din(w_dff_A_MOmaS9wo9_0),.clk(gclk));
	jdff dff_A_ZrhELOdn8_0(.dout(w_dff_A_JEg0rFPI8_0),.din(w_dff_A_ZrhELOdn8_0),.clk(gclk));
	jdff dff_A_JEg0rFPI8_0(.dout(w_dff_A_nsnh1dY66_0),.din(w_dff_A_JEg0rFPI8_0),.clk(gclk));
	jdff dff_A_nsnh1dY66_0(.dout(w_dff_A_FMHQIao37_0),.din(w_dff_A_nsnh1dY66_0),.clk(gclk));
	jdff dff_A_FMHQIao37_0(.dout(w_dff_A_5c5TmNXW1_0),.din(w_dff_A_FMHQIao37_0),.clk(gclk));
	jdff dff_A_5c5TmNXW1_0(.dout(w_dff_A_MkWXwYFV8_0),.din(w_dff_A_5c5TmNXW1_0),.clk(gclk));
	jdff dff_A_MkWXwYFV8_0(.dout(G3),.din(w_dff_A_MkWXwYFV8_0),.clk(gclk));
	jdff dff_A_P8WDRkB32_1(.dout(w_dff_A_KEHXtWQB4_0),.din(w_dff_A_P8WDRkB32_1),.clk(gclk));
	jdff dff_A_KEHXtWQB4_0(.dout(w_dff_A_UJBNpKNU2_0),.din(w_dff_A_KEHXtWQB4_0),.clk(gclk));
	jdff dff_A_UJBNpKNU2_0(.dout(w_dff_A_CnjPptcQ8_0),.din(w_dff_A_UJBNpKNU2_0),.clk(gclk));
	jdff dff_A_CnjPptcQ8_0(.dout(w_dff_A_DJbw1rEN1_0),.din(w_dff_A_CnjPptcQ8_0),.clk(gclk));
	jdff dff_A_DJbw1rEN1_0(.dout(w_dff_A_vw3tfYfV2_0),.din(w_dff_A_DJbw1rEN1_0),.clk(gclk));
	jdff dff_A_vw3tfYfV2_0(.dout(w_dff_A_q63BVYZV5_0),.din(w_dff_A_vw3tfYfV2_0),.clk(gclk));
	jdff dff_A_q63BVYZV5_0(.dout(w_dff_A_aTPQEO3a4_0),.din(w_dff_A_q63BVYZV5_0),.clk(gclk));
	jdff dff_A_aTPQEO3a4_0(.dout(w_dff_A_6ZHdjy9k2_0),.din(w_dff_A_aTPQEO3a4_0),.clk(gclk));
	jdff dff_A_6ZHdjy9k2_0(.dout(w_dff_A_s0xYhP2F4_0),.din(w_dff_A_6ZHdjy9k2_0),.clk(gclk));
	jdff dff_A_s0xYhP2F4_0(.dout(w_dff_A_QZKpCIPp1_0),.din(w_dff_A_s0xYhP2F4_0),.clk(gclk));
	jdff dff_A_QZKpCIPp1_0(.dout(w_dff_A_jUL6YSMs4_0),.din(w_dff_A_QZKpCIPp1_0),.clk(gclk));
	jdff dff_A_jUL6YSMs4_0(.dout(w_dff_A_sFgDPNML0_0),.din(w_dff_A_jUL6YSMs4_0),.clk(gclk));
	jdff dff_A_sFgDPNML0_0(.dout(w_dff_A_8kX9Yz7G6_0),.din(w_dff_A_sFgDPNML0_0),.clk(gclk));
	jdff dff_A_8kX9Yz7G6_0(.dout(w_dff_A_mcy3O4Vt9_0),.din(w_dff_A_8kX9Yz7G6_0),.clk(gclk));
	jdff dff_A_mcy3O4Vt9_0(.dout(w_dff_A_FoGZ3b4J6_0),.din(w_dff_A_mcy3O4Vt9_0),.clk(gclk));
	jdff dff_A_FoGZ3b4J6_0(.dout(w_dff_A_cqTPpmCQ6_0),.din(w_dff_A_FoGZ3b4J6_0),.clk(gclk));
	jdff dff_A_cqTPpmCQ6_0(.dout(w_dff_A_ys8UfOQC0_0),.din(w_dff_A_cqTPpmCQ6_0),.clk(gclk));
	jdff dff_A_ys8UfOQC0_0(.dout(w_dff_A_k9OYpDMQ2_0),.din(w_dff_A_ys8UfOQC0_0),.clk(gclk));
	jdff dff_A_k9OYpDMQ2_0(.dout(w_dff_A_7uDRE68t8_0),.din(w_dff_A_k9OYpDMQ2_0),.clk(gclk));
	jdff dff_A_7uDRE68t8_0(.dout(w_dff_A_qXWQFPdP2_0),.din(w_dff_A_7uDRE68t8_0),.clk(gclk));
	jdff dff_A_qXWQFPdP2_0(.dout(w_dff_A_pwGBwSRd0_0),.din(w_dff_A_qXWQFPdP2_0),.clk(gclk));
	jdff dff_A_pwGBwSRd0_0(.dout(w_dff_A_oQ0QB7Ng0_0),.din(w_dff_A_pwGBwSRd0_0),.clk(gclk));
	jdff dff_A_oQ0QB7Ng0_0(.dout(w_dff_A_VU4g507v9_0),.din(w_dff_A_oQ0QB7Ng0_0),.clk(gclk));
	jdff dff_A_VU4g507v9_0(.dout(w_dff_A_Sn8GvQn42_0),.din(w_dff_A_VU4g507v9_0),.clk(gclk));
	jdff dff_A_Sn8GvQn42_0(.dout(w_dff_A_uKOB4OED5_0),.din(w_dff_A_Sn8GvQn42_0),.clk(gclk));
	jdff dff_A_uKOB4OED5_0(.dout(w_dff_A_aYR3FIJa8_0),.din(w_dff_A_uKOB4OED5_0),.clk(gclk));
	jdff dff_A_aYR3FIJa8_0(.dout(w_dff_A_6wknBOYK4_0),.din(w_dff_A_aYR3FIJa8_0),.clk(gclk));
	jdff dff_A_6wknBOYK4_0(.dout(w_dff_A_8xsSwGYc3_0),.din(w_dff_A_6wknBOYK4_0),.clk(gclk));
	jdff dff_A_8xsSwGYc3_0(.dout(w_dff_A_KTg2UkOS6_0),.din(w_dff_A_8xsSwGYc3_0),.clk(gclk));
	jdff dff_A_KTg2UkOS6_0(.dout(w_dff_A_1mGoiPaC2_0),.din(w_dff_A_KTg2UkOS6_0),.clk(gclk));
	jdff dff_A_1mGoiPaC2_0(.dout(w_dff_A_YNf3TYu26_0),.din(w_dff_A_1mGoiPaC2_0),.clk(gclk));
	jdff dff_A_YNf3TYu26_0(.dout(w_dff_A_rR7wkgtB4_0),.din(w_dff_A_YNf3TYu26_0),.clk(gclk));
	jdff dff_A_rR7wkgtB4_0(.dout(w_dff_A_R6k27Hmj9_0),.din(w_dff_A_rR7wkgtB4_0),.clk(gclk));
	jdff dff_A_R6k27Hmj9_0(.dout(w_dff_A_gANCoK860_0),.din(w_dff_A_R6k27Hmj9_0),.clk(gclk));
	jdff dff_A_gANCoK860_0(.dout(w_dff_A_lLSRErtM9_0),.din(w_dff_A_gANCoK860_0),.clk(gclk));
	jdff dff_A_lLSRErtM9_0(.dout(w_dff_A_mSM3Ycj02_0),.din(w_dff_A_lLSRErtM9_0),.clk(gclk));
	jdff dff_A_mSM3Ycj02_0(.dout(w_dff_A_0M3qaGI70_0),.din(w_dff_A_mSM3Ycj02_0),.clk(gclk));
	jdff dff_A_0M3qaGI70_0(.dout(w_dff_A_dNfSPOfu6_0),.din(w_dff_A_0M3qaGI70_0),.clk(gclk));
	jdff dff_A_dNfSPOfu6_0(.dout(G450),.din(w_dff_A_dNfSPOfu6_0),.clk(gclk));
	jdff dff_A_IflYUUBn6_1(.dout(w_dff_A_sRfM7A0E4_0),.din(w_dff_A_IflYUUBn6_1),.clk(gclk));
	jdff dff_A_sRfM7A0E4_0(.dout(w_dff_A_MNfhiR7A3_0),.din(w_dff_A_sRfM7A0E4_0),.clk(gclk));
	jdff dff_A_MNfhiR7A3_0(.dout(w_dff_A_QkfOOnRg4_0),.din(w_dff_A_MNfhiR7A3_0),.clk(gclk));
	jdff dff_A_QkfOOnRg4_0(.dout(w_dff_A_g3qdOyMo7_0),.din(w_dff_A_QkfOOnRg4_0),.clk(gclk));
	jdff dff_A_g3qdOyMo7_0(.dout(w_dff_A_GAsH9soI5_0),.din(w_dff_A_g3qdOyMo7_0),.clk(gclk));
	jdff dff_A_GAsH9soI5_0(.dout(w_dff_A_gJZmpSG89_0),.din(w_dff_A_GAsH9soI5_0),.clk(gclk));
	jdff dff_A_gJZmpSG89_0(.dout(w_dff_A_SfiU2wq33_0),.din(w_dff_A_gJZmpSG89_0),.clk(gclk));
	jdff dff_A_SfiU2wq33_0(.dout(w_dff_A_jMQZZB073_0),.din(w_dff_A_SfiU2wq33_0),.clk(gclk));
	jdff dff_A_jMQZZB073_0(.dout(w_dff_A_rUdNl4IU4_0),.din(w_dff_A_jMQZZB073_0),.clk(gclk));
	jdff dff_A_rUdNl4IU4_0(.dout(w_dff_A_q7QZp0hU4_0),.din(w_dff_A_rUdNl4IU4_0),.clk(gclk));
	jdff dff_A_q7QZp0hU4_0(.dout(w_dff_A_k3Pyj5zi3_0),.din(w_dff_A_q7QZp0hU4_0),.clk(gclk));
	jdff dff_A_k3Pyj5zi3_0(.dout(w_dff_A_GZjy3eqv4_0),.din(w_dff_A_k3Pyj5zi3_0),.clk(gclk));
	jdff dff_A_GZjy3eqv4_0(.dout(w_dff_A_4ybbnZ511_0),.din(w_dff_A_GZjy3eqv4_0),.clk(gclk));
	jdff dff_A_4ybbnZ511_0(.dout(w_dff_A_Lk4OfqAX8_0),.din(w_dff_A_4ybbnZ511_0),.clk(gclk));
	jdff dff_A_Lk4OfqAX8_0(.dout(w_dff_A_ceuXNrKz2_0),.din(w_dff_A_Lk4OfqAX8_0),.clk(gclk));
	jdff dff_A_ceuXNrKz2_0(.dout(w_dff_A_Qla1hDku4_0),.din(w_dff_A_ceuXNrKz2_0),.clk(gclk));
	jdff dff_A_Qla1hDku4_0(.dout(w_dff_A_qnhBl79k4_0),.din(w_dff_A_Qla1hDku4_0),.clk(gclk));
	jdff dff_A_qnhBl79k4_0(.dout(w_dff_A_H8FAlFuI8_0),.din(w_dff_A_qnhBl79k4_0),.clk(gclk));
	jdff dff_A_H8FAlFuI8_0(.dout(w_dff_A_TMJ7B2sj0_0),.din(w_dff_A_H8FAlFuI8_0),.clk(gclk));
	jdff dff_A_TMJ7B2sj0_0(.dout(w_dff_A_1E2AD5X72_0),.din(w_dff_A_TMJ7B2sj0_0),.clk(gclk));
	jdff dff_A_1E2AD5X72_0(.dout(w_dff_A_Yum01tnZ1_0),.din(w_dff_A_1E2AD5X72_0),.clk(gclk));
	jdff dff_A_Yum01tnZ1_0(.dout(w_dff_A_riiZSMiM5_0),.din(w_dff_A_Yum01tnZ1_0),.clk(gclk));
	jdff dff_A_riiZSMiM5_0(.dout(w_dff_A_Mo2MkYzG5_0),.din(w_dff_A_riiZSMiM5_0),.clk(gclk));
	jdff dff_A_Mo2MkYzG5_0(.dout(w_dff_A_uKon5cKx9_0),.din(w_dff_A_Mo2MkYzG5_0),.clk(gclk));
	jdff dff_A_uKon5cKx9_0(.dout(w_dff_A_2iCK4iSu6_0),.din(w_dff_A_uKon5cKx9_0),.clk(gclk));
	jdff dff_A_2iCK4iSu6_0(.dout(w_dff_A_R7t4Bh989_0),.din(w_dff_A_2iCK4iSu6_0),.clk(gclk));
	jdff dff_A_R7t4Bh989_0(.dout(w_dff_A_Me7Q28lX7_0),.din(w_dff_A_R7t4Bh989_0),.clk(gclk));
	jdff dff_A_Me7Q28lX7_0(.dout(w_dff_A_g3Mop0g48_0),.din(w_dff_A_Me7Q28lX7_0),.clk(gclk));
	jdff dff_A_g3Mop0g48_0(.dout(w_dff_A_sUHsZpr36_0),.din(w_dff_A_g3Mop0g48_0),.clk(gclk));
	jdff dff_A_sUHsZpr36_0(.dout(w_dff_A_loEuQvIp0_0),.din(w_dff_A_sUHsZpr36_0),.clk(gclk));
	jdff dff_A_loEuQvIp0_0(.dout(w_dff_A_2Di6GwsR7_0),.din(w_dff_A_loEuQvIp0_0),.clk(gclk));
	jdff dff_A_2Di6GwsR7_0(.dout(w_dff_A_PZVXZ8I75_0),.din(w_dff_A_2Di6GwsR7_0),.clk(gclk));
	jdff dff_A_PZVXZ8I75_0(.dout(w_dff_A_SZ2yEkf29_0),.din(w_dff_A_PZVXZ8I75_0),.clk(gclk));
	jdff dff_A_SZ2yEkf29_0(.dout(w_dff_A_17KJYLmk1_0),.din(w_dff_A_SZ2yEkf29_0),.clk(gclk));
	jdff dff_A_17KJYLmk1_0(.dout(w_dff_A_v9mhp5IQ1_0),.din(w_dff_A_17KJYLmk1_0),.clk(gclk));
	jdff dff_A_v9mhp5IQ1_0(.dout(w_dff_A_e2B9nFVc9_0),.din(w_dff_A_v9mhp5IQ1_0),.clk(gclk));
	jdff dff_A_e2B9nFVc9_0(.dout(w_dff_A_eUhlLYI76_0),.din(w_dff_A_e2B9nFVc9_0),.clk(gclk));
	jdff dff_A_eUhlLYI76_0(.dout(w_dff_A_F88TuU6w1_0),.din(w_dff_A_eUhlLYI76_0),.clk(gclk));
	jdff dff_A_F88TuU6w1_0(.dout(G448),.din(w_dff_A_F88TuU6w1_0),.clk(gclk));
	jdff dff_A_U5TrYOk95_1(.dout(w_dff_A_Ha7yNAiw9_0),.din(w_dff_A_U5TrYOk95_1),.clk(gclk));
	jdff dff_A_Ha7yNAiw9_0(.dout(w_dff_A_slcV6hqE4_0),.din(w_dff_A_Ha7yNAiw9_0),.clk(gclk));
	jdff dff_A_slcV6hqE4_0(.dout(w_dff_A_7L2sUl0W4_0),.din(w_dff_A_slcV6hqE4_0),.clk(gclk));
	jdff dff_A_7L2sUl0W4_0(.dout(w_dff_A_ZSx6VU495_0),.din(w_dff_A_7L2sUl0W4_0),.clk(gclk));
	jdff dff_A_ZSx6VU495_0(.dout(w_dff_A_CX9L5Eh40_0),.din(w_dff_A_ZSx6VU495_0),.clk(gclk));
	jdff dff_A_CX9L5Eh40_0(.dout(w_dff_A_W2hgN4rB7_0),.din(w_dff_A_CX9L5Eh40_0),.clk(gclk));
	jdff dff_A_W2hgN4rB7_0(.dout(w_dff_A_wBwQtfQe4_0),.din(w_dff_A_W2hgN4rB7_0),.clk(gclk));
	jdff dff_A_wBwQtfQe4_0(.dout(w_dff_A_OHemJ8Og7_0),.din(w_dff_A_wBwQtfQe4_0),.clk(gclk));
	jdff dff_A_OHemJ8Og7_0(.dout(w_dff_A_DOG31mfW3_0),.din(w_dff_A_OHemJ8Og7_0),.clk(gclk));
	jdff dff_A_DOG31mfW3_0(.dout(w_dff_A_VFKnqIhs2_0),.din(w_dff_A_DOG31mfW3_0),.clk(gclk));
	jdff dff_A_VFKnqIhs2_0(.dout(w_dff_A_x4nytnbj4_0),.din(w_dff_A_VFKnqIhs2_0),.clk(gclk));
	jdff dff_A_x4nytnbj4_0(.dout(w_dff_A_uvOLy8EJ5_0),.din(w_dff_A_x4nytnbj4_0),.clk(gclk));
	jdff dff_A_uvOLy8EJ5_0(.dout(w_dff_A_mKXF3PJ13_0),.din(w_dff_A_uvOLy8EJ5_0),.clk(gclk));
	jdff dff_A_mKXF3PJ13_0(.dout(w_dff_A_4xpbHIkx7_0),.din(w_dff_A_mKXF3PJ13_0),.clk(gclk));
	jdff dff_A_4xpbHIkx7_0(.dout(w_dff_A_fAI54q1Z8_0),.din(w_dff_A_4xpbHIkx7_0),.clk(gclk));
	jdff dff_A_fAI54q1Z8_0(.dout(w_dff_A_hHMApKnQ7_0),.din(w_dff_A_fAI54q1Z8_0),.clk(gclk));
	jdff dff_A_hHMApKnQ7_0(.dout(w_dff_A_Sc8i3oMz1_0),.din(w_dff_A_hHMApKnQ7_0),.clk(gclk));
	jdff dff_A_Sc8i3oMz1_0(.dout(w_dff_A_EHHXM7mv5_0),.din(w_dff_A_Sc8i3oMz1_0),.clk(gclk));
	jdff dff_A_EHHXM7mv5_0(.dout(w_dff_A_HgFIT1074_0),.din(w_dff_A_EHHXM7mv5_0),.clk(gclk));
	jdff dff_A_HgFIT1074_0(.dout(w_dff_A_tWKdS0U72_0),.din(w_dff_A_HgFIT1074_0),.clk(gclk));
	jdff dff_A_tWKdS0U72_0(.dout(w_dff_A_JNmXtZol5_0),.din(w_dff_A_tWKdS0U72_0),.clk(gclk));
	jdff dff_A_JNmXtZol5_0(.dout(w_dff_A_A1wy8V5y0_0),.din(w_dff_A_JNmXtZol5_0),.clk(gclk));
	jdff dff_A_A1wy8V5y0_0(.dout(w_dff_A_gRruVxYW7_0),.din(w_dff_A_A1wy8V5y0_0),.clk(gclk));
	jdff dff_A_gRruVxYW7_0(.dout(w_dff_A_vAbBGfvT7_0),.din(w_dff_A_gRruVxYW7_0),.clk(gclk));
	jdff dff_A_vAbBGfvT7_0(.dout(w_dff_A_cKuSHqRn2_0),.din(w_dff_A_vAbBGfvT7_0),.clk(gclk));
	jdff dff_A_cKuSHqRn2_0(.dout(w_dff_A_EphTaOWz2_0),.din(w_dff_A_cKuSHqRn2_0),.clk(gclk));
	jdff dff_A_EphTaOWz2_0(.dout(w_dff_A_hA8FtDgM4_0),.din(w_dff_A_EphTaOWz2_0),.clk(gclk));
	jdff dff_A_hA8FtDgM4_0(.dout(w_dff_A_BQAqS9To6_0),.din(w_dff_A_hA8FtDgM4_0),.clk(gclk));
	jdff dff_A_BQAqS9To6_0(.dout(w_dff_A_GZ8iJtLX9_0),.din(w_dff_A_BQAqS9To6_0),.clk(gclk));
	jdff dff_A_GZ8iJtLX9_0(.dout(w_dff_A_yO26HhJC5_0),.din(w_dff_A_GZ8iJtLX9_0),.clk(gclk));
	jdff dff_A_yO26HhJC5_0(.dout(w_dff_A_9tAFCkcm5_0),.din(w_dff_A_yO26HhJC5_0),.clk(gclk));
	jdff dff_A_9tAFCkcm5_0(.dout(w_dff_A_LM3GAe8w9_0),.din(w_dff_A_9tAFCkcm5_0),.clk(gclk));
	jdff dff_A_LM3GAe8w9_0(.dout(w_dff_A_Dl0QZvSs6_0),.din(w_dff_A_LM3GAe8w9_0),.clk(gclk));
	jdff dff_A_Dl0QZvSs6_0(.dout(w_dff_A_8cOZigAO0_0),.din(w_dff_A_Dl0QZvSs6_0),.clk(gclk));
	jdff dff_A_8cOZigAO0_0(.dout(w_dff_A_I419XbQu8_0),.din(w_dff_A_8cOZigAO0_0),.clk(gclk));
	jdff dff_A_I419XbQu8_0(.dout(w_dff_A_CZA5ch9p3_0),.din(w_dff_A_I419XbQu8_0),.clk(gclk));
	jdff dff_A_CZA5ch9p3_0(.dout(w_dff_A_5palj88r8_0),.din(w_dff_A_CZA5ch9p3_0),.clk(gclk));
	jdff dff_A_5palj88r8_0(.dout(w_dff_A_WS0xxbFA7_0),.din(w_dff_A_5palj88r8_0),.clk(gclk));
	jdff dff_A_WS0xxbFA7_0(.dout(G444),.din(w_dff_A_WS0xxbFA7_0),.clk(gclk));
	jdff dff_A_YONsQmPY7_1(.dout(w_dff_A_ANmmdNnK4_0),.din(w_dff_A_YONsQmPY7_1),.clk(gclk));
	jdff dff_A_ANmmdNnK4_0(.dout(w_dff_A_ocVinIXo1_0),.din(w_dff_A_ANmmdNnK4_0),.clk(gclk));
	jdff dff_A_ocVinIXo1_0(.dout(w_dff_A_r2jLnFdC5_0),.din(w_dff_A_ocVinIXo1_0),.clk(gclk));
	jdff dff_A_r2jLnFdC5_0(.dout(w_dff_A_RxI2ZLu16_0),.din(w_dff_A_r2jLnFdC5_0),.clk(gclk));
	jdff dff_A_RxI2ZLu16_0(.dout(w_dff_A_IReLaPoU4_0),.din(w_dff_A_RxI2ZLu16_0),.clk(gclk));
	jdff dff_A_IReLaPoU4_0(.dout(w_dff_A_plkQnMZJ0_0),.din(w_dff_A_IReLaPoU4_0),.clk(gclk));
	jdff dff_A_plkQnMZJ0_0(.dout(w_dff_A_9AF9riub7_0),.din(w_dff_A_plkQnMZJ0_0),.clk(gclk));
	jdff dff_A_9AF9riub7_0(.dout(w_dff_A_aFM7aReY6_0),.din(w_dff_A_9AF9riub7_0),.clk(gclk));
	jdff dff_A_aFM7aReY6_0(.dout(w_dff_A_fW4BfWbg9_0),.din(w_dff_A_aFM7aReY6_0),.clk(gclk));
	jdff dff_A_fW4BfWbg9_0(.dout(w_dff_A_S7jIUXO43_0),.din(w_dff_A_fW4BfWbg9_0),.clk(gclk));
	jdff dff_A_S7jIUXO43_0(.dout(w_dff_A_Bjv6ZlqM1_0),.din(w_dff_A_S7jIUXO43_0),.clk(gclk));
	jdff dff_A_Bjv6ZlqM1_0(.dout(w_dff_A_pZYdD4oV8_0),.din(w_dff_A_Bjv6ZlqM1_0),.clk(gclk));
	jdff dff_A_pZYdD4oV8_0(.dout(w_dff_A_1EjCeFcd6_0),.din(w_dff_A_pZYdD4oV8_0),.clk(gclk));
	jdff dff_A_1EjCeFcd6_0(.dout(w_dff_A_tgDDu5xY7_0),.din(w_dff_A_1EjCeFcd6_0),.clk(gclk));
	jdff dff_A_tgDDu5xY7_0(.dout(w_dff_A_fn7e7yzk7_0),.din(w_dff_A_tgDDu5xY7_0),.clk(gclk));
	jdff dff_A_fn7e7yzk7_0(.dout(w_dff_A_Z28NkXa77_0),.din(w_dff_A_fn7e7yzk7_0),.clk(gclk));
	jdff dff_A_Z28NkXa77_0(.dout(w_dff_A_dRqEIt030_0),.din(w_dff_A_Z28NkXa77_0),.clk(gclk));
	jdff dff_A_dRqEIt030_0(.dout(w_dff_A_yyTncQKg7_0),.din(w_dff_A_dRqEIt030_0),.clk(gclk));
	jdff dff_A_yyTncQKg7_0(.dout(w_dff_A_uBVxEl2A2_0),.din(w_dff_A_yyTncQKg7_0),.clk(gclk));
	jdff dff_A_uBVxEl2A2_0(.dout(w_dff_A_HhUoXcMG6_0),.din(w_dff_A_uBVxEl2A2_0),.clk(gclk));
	jdff dff_A_HhUoXcMG6_0(.dout(w_dff_A_IX4uyESn0_0),.din(w_dff_A_HhUoXcMG6_0),.clk(gclk));
	jdff dff_A_IX4uyESn0_0(.dout(w_dff_A_MpTDP1oo8_0),.din(w_dff_A_IX4uyESn0_0),.clk(gclk));
	jdff dff_A_MpTDP1oo8_0(.dout(w_dff_A_ahQ8esOF0_0),.din(w_dff_A_MpTDP1oo8_0),.clk(gclk));
	jdff dff_A_ahQ8esOF0_0(.dout(w_dff_A_lAzi9spV8_0),.din(w_dff_A_ahQ8esOF0_0),.clk(gclk));
	jdff dff_A_lAzi9spV8_0(.dout(w_dff_A_7CfKEnZE7_0),.din(w_dff_A_lAzi9spV8_0),.clk(gclk));
	jdff dff_A_7CfKEnZE7_0(.dout(w_dff_A_B3sh92i29_0),.din(w_dff_A_7CfKEnZE7_0),.clk(gclk));
	jdff dff_A_B3sh92i29_0(.dout(w_dff_A_vHapubzK1_0),.din(w_dff_A_B3sh92i29_0),.clk(gclk));
	jdff dff_A_vHapubzK1_0(.dout(w_dff_A_RvlRpLbA4_0),.din(w_dff_A_vHapubzK1_0),.clk(gclk));
	jdff dff_A_RvlRpLbA4_0(.dout(w_dff_A_yUTz5umu0_0),.din(w_dff_A_RvlRpLbA4_0),.clk(gclk));
	jdff dff_A_yUTz5umu0_0(.dout(w_dff_A_CVSsUflQ9_0),.din(w_dff_A_yUTz5umu0_0),.clk(gclk));
	jdff dff_A_CVSsUflQ9_0(.dout(w_dff_A_IexcqqmL7_0),.din(w_dff_A_CVSsUflQ9_0),.clk(gclk));
	jdff dff_A_IexcqqmL7_0(.dout(w_dff_A_A64mRuOH6_0),.din(w_dff_A_IexcqqmL7_0),.clk(gclk));
	jdff dff_A_A64mRuOH6_0(.dout(w_dff_A_NZNjYFxx6_0),.din(w_dff_A_A64mRuOH6_0),.clk(gclk));
	jdff dff_A_NZNjYFxx6_0(.dout(w_dff_A_MZo8jf6F9_0),.din(w_dff_A_NZNjYFxx6_0),.clk(gclk));
	jdff dff_A_MZo8jf6F9_0(.dout(w_dff_A_A4fl1uXn7_0),.din(w_dff_A_MZo8jf6F9_0),.clk(gclk));
	jdff dff_A_A4fl1uXn7_0(.dout(w_dff_A_mT9j2k6k2_0),.din(w_dff_A_A4fl1uXn7_0),.clk(gclk));
	jdff dff_A_mT9j2k6k2_0(.dout(w_dff_A_esLmSjHq2_0),.din(w_dff_A_mT9j2k6k2_0),.clk(gclk));
	jdff dff_A_esLmSjHq2_0(.dout(w_dff_A_ZdOEwVqN9_0),.din(w_dff_A_esLmSjHq2_0),.clk(gclk));
	jdff dff_A_ZdOEwVqN9_0(.dout(G442),.din(w_dff_A_ZdOEwVqN9_0),.clk(gclk));
	jdff dff_A_7MrFhR7S7_1(.dout(w_dff_A_TAl1qSZX8_0),.din(w_dff_A_7MrFhR7S7_1),.clk(gclk));
	jdff dff_A_TAl1qSZX8_0(.dout(w_dff_A_EYxxYUb76_0),.din(w_dff_A_TAl1qSZX8_0),.clk(gclk));
	jdff dff_A_EYxxYUb76_0(.dout(w_dff_A_jZhC1kvW8_0),.din(w_dff_A_EYxxYUb76_0),.clk(gclk));
	jdff dff_A_jZhC1kvW8_0(.dout(w_dff_A_T53HvLAY2_0),.din(w_dff_A_jZhC1kvW8_0),.clk(gclk));
	jdff dff_A_T53HvLAY2_0(.dout(w_dff_A_nORdTeXw7_0),.din(w_dff_A_T53HvLAY2_0),.clk(gclk));
	jdff dff_A_nORdTeXw7_0(.dout(w_dff_A_N8JPfGWk1_0),.din(w_dff_A_nORdTeXw7_0),.clk(gclk));
	jdff dff_A_N8JPfGWk1_0(.dout(w_dff_A_isovUuZR6_0),.din(w_dff_A_N8JPfGWk1_0),.clk(gclk));
	jdff dff_A_isovUuZR6_0(.dout(w_dff_A_3QlqfaK12_0),.din(w_dff_A_isovUuZR6_0),.clk(gclk));
	jdff dff_A_3QlqfaK12_0(.dout(w_dff_A_4ive3bFb7_0),.din(w_dff_A_3QlqfaK12_0),.clk(gclk));
	jdff dff_A_4ive3bFb7_0(.dout(w_dff_A_9n3qgERt5_0),.din(w_dff_A_4ive3bFb7_0),.clk(gclk));
	jdff dff_A_9n3qgERt5_0(.dout(w_dff_A_mRbFvcOQ5_0),.din(w_dff_A_9n3qgERt5_0),.clk(gclk));
	jdff dff_A_mRbFvcOQ5_0(.dout(w_dff_A_aDmuAb4J1_0),.din(w_dff_A_mRbFvcOQ5_0),.clk(gclk));
	jdff dff_A_aDmuAb4J1_0(.dout(w_dff_A_CowIdsDB3_0),.din(w_dff_A_aDmuAb4J1_0),.clk(gclk));
	jdff dff_A_CowIdsDB3_0(.dout(w_dff_A_DOjiXBQO1_0),.din(w_dff_A_CowIdsDB3_0),.clk(gclk));
	jdff dff_A_DOjiXBQO1_0(.dout(w_dff_A_kL1awfcf6_0),.din(w_dff_A_DOjiXBQO1_0),.clk(gclk));
	jdff dff_A_kL1awfcf6_0(.dout(w_dff_A_dUbhyRtm2_0),.din(w_dff_A_kL1awfcf6_0),.clk(gclk));
	jdff dff_A_dUbhyRtm2_0(.dout(w_dff_A_foOBI6LB9_0),.din(w_dff_A_dUbhyRtm2_0),.clk(gclk));
	jdff dff_A_foOBI6LB9_0(.dout(w_dff_A_OJkDzmtM1_0),.din(w_dff_A_foOBI6LB9_0),.clk(gclk));
	jdff dff_A_OJkDzmtM1_0(.dout(w_dff_A_kwQgiElp5_0),.din(w_dff_A_OJkDzmtM1_0),.clk(gclk));
	jdff dff_A_kwQgiElp5_0(.dout(w_dff_A_tzvoNRdm7_0),.din(w_dff_A_kwQgiElp5_0),.clk(gclk));
	jdff dff_A_tzvoNRdm7_0(.dout(w_dff_A_0uDydB9g0_0),.din(w_dff_A_tzvoNRdm7_0),.clk(gclk));
	jdff dff_A_0uDydB9g0_0(.dout(w_dff_A_9cVVqneJ3_0),.din(w_dff_A_0uDydB9g0_0),.clk(gclk));
	jdff dff_A_9cVVqneJ3_0(.dout(w_dff_A_4EesM9SE6_0),.din(w_dff_A_9cVVqneJ3_0),.clk(gclk));
	jdff dff_A_4EesM9SE6_0(.dout(w_dff_A_fmrxib7m7_0),.din(w_dff_A_4EesM9SE6_0),.clk(gclk));
	jdff dff_A_fmrxib7m7_0(.dout(w_dff_A_nmoeL7v56_0),.din(w_dff_A_fmrxib7m7_0),.clk(gclk));
	jdff dff_A_nmoeL7v56_0(.dout(w_dff_A_cKOyWVtE7_0),.din(w_dff_A_nmoeL7v56_0),.clk(gclk));
	jdff dff_A_cKOyWVtE7_0(.dout(w_dff_A_ODhR2nVm7_0),.din(w_dff_A_cKOyWVtE7_0),.clk(gclk));
	jdff dff_A_ODhR2nVm7_0(.dout(w_dff_A_4mMJ0EFX4_0),.din(w_dff_A_ODhR2nVm7_0),.clk(gclk));
	jdff dff_A_4mMJ0EFX4_0(.dout(w_dff_A_psWdfyE05_0),.din(w_dff_A_4mMJ0EFX4_0),.clk(gclk));
	jdff dff_A_psWdfyE05_0(.dout(w_dff_A_SdQ5bftN2_0),.din(w_dff_A_psWdfyE05_0),.clk(gclk));
	jdff dff_A_SdQ5bftN2_0(.dout(w_dff_A_82CSJO2B4_0),.din(w_dff_A_SdQ5bftN2_0),.clk(gclk));
	jdff dff_A_82CSJO2B4_0(.dout(w_dff_A_3RbBVgOa7_0),.din(w_dff_A_82CSJO2B4_0),.clk(gclk));
	jdff dff_A_3RbBVgOa7_0(.dout(w_dff_A_2K8lkq8h9_0),.din(w_dff_A_3RbBVgOa7_0),.clk(gclk));
	jdff dff_A_2K8lkq8h9_0(.dout(w_dff_A_TZcd6i835_0),.din(w_dff_A_2K8lkq8h9_0),.clk(gclk));
	jdff dff_A_TZcd6i835_0(.dout(w_dff_A_gBHDVGLn4_0),.din(w_dff_A_TZcd6i835_0),.clk(gclk));
	jdff dff_A_gBHDVGLn4_0(.dout(w_dff_A_TgrAWO958_0),.din(w_dff_A_gBHDVGLn4_0),.clk(gclk));
	jdff dff_A_TgrAWO958_0(.dout(w_dff_A_39xY3sph6_0),.din(w_dff_A_TgrAWO958_0),.clk(gclk));
	jdff dff_A_39xY3sph6_0(.dout(w_dff_A_BvoqxjG86_0),.din(w_dff_A_39xY3sph6_0),.clk(gclk));
	jdff dff_A_BvoqxjG86_0(.dout(G440),.din(w_dff_A_BvoqxjG86_0),.clk(gclk));
	jdff dff_A_pV3lp2Th7_1(.dout(w_dff_A_KM9CCsM21_0),.din(w_dff_A_pV3lp2Th7_1),.clk(gclk));
	jdff dff_A_KM9CCsM21_0(.dout(w_dff_A_Cz2Bgu0c8_0),.din(w_dff_A_KM9CCsM21_0),.clk(gclk));
	jdff dff_A_Cz2Bgu0c8_0(.dout(w_dff_A_N2B4mVHN3_0),.din(w_dff_A_Cz2Bgu0c8_0),.clk(gclk));
	jdff dff_A_N2B4mVHN3_0(.dout(w_dff_A_IZCYFMx61_0),.din(w_dff_A_N2B4mVHN3_0),.clk(gclk));
	jdff dff_A_IZCYFMx61_0(.dout(w_dff_A_JXMqe9UU5_0),.din(w_dff_A_IZCYFMx61_0),.clk(gclk));
	jdff dff_A_JXMqe9UU5_0(.dout(w_dff_A_J6Y33yuM1_0),.din(w_dff_A_JXMqe9UU5_0),.clk(gclk));
	jdff dff_A_J6Y33yuM1_0(.dout(w_dff_A_dldMPbnL7_0),.din(w_dff_A_J6Y33yuM1_0),.clk(gclk));
	jdff dff_A_dldMPbnL7_0(.dout(w_dff_A_B0MieEWu6_0),.din(w_dff_A_dldMPbnL7_0),.clk(gclk));
	jdff dff_A_B0MieEWu6_0(.dout(w_dff_A_fJhsAtbk0_0),.din(w_dff_A_B0MieEWu6_0),.clk(gclk));
	jdff dff_A_fJhsAtbk0_0(.dout(w_dff_A_aYLOhwJI1_0),.din(w_dff_A_fJhsAtbk0_0),.clk(gclk));
	jdff dff_A_aYLOhwJI1_0(.dout(w_dff_A_tXbivGwa3_0),.din(w_dff_A_aYLOhwJI1_0),.clk(gclk));
	jdff dff_A_tXbivGwa3_0(.dout(w_dff_A_rhnjMU0J6_0),.din(w_dff_A_tXbivGwa3_0),.clk(gclk));
	jdff dff_A_rhnjMU0J6_0(.dout(w_dff_A_V7gHNQQU7_0),.din(w_dff_A_rhnjMU0J6_0),.clk(gclk));
	jdff dff_A_V7gHNQQU7_0(.dout(w_dff_A_3EpC6Hfn8_0),.din(w_dff_A_V7gHNQQU7_0),.clk(gclk));
	jdff dff_A_3EpC6Hfn8_0(.dout(w_dff_A_uTMGRQJi3_0),.din(w_dff_A_3EpC6Hfn8_0),.clk(gclk));
	jdff dff_A_uTMGRQJi3_0(.dout(w_dff_A_cx9rXWYN8_0),.din(w_dff_A_uTMGRQJi3_0),.clk(gclk));
	jdff dff_A_cx9rXWYN8_0(.dout(w_dff_A_hE08VOWD2_0),.din(w_dff_A_cx9rXWYN8_0),.clk(gclk));
	jdff dff_A_hE08VOWD2_0(.dout(w_dff_A_uhHmn1Ot2_0),.din(w_dff_A_hE08VOWD2_0),.clk(gclk));
	jdff dff_A_uhHmn1Ot2_0(.dout(w_dff_A_etEJ1VS64_0),.din(w_dff_A_uhHmn1Ot2_0),.clk(gclk));
	jdff dff_A_etEJ1VS64_0(.dout(w_dff_A_kDuKOeZi7_0),.din(w_dff_A_etEJ1VS64_0),.clk(gclk));
	jdff dff_A_kDuKOeZi7_0(.dout(w_dff_A_vzR2OpQl1_0),.din(w_dff_A_kDuKOeZi7_0),.clk(gclk));
	jdff dff_A_vzR2OpQl1_0(.dout(w_dff_A_f7dHFFwu5_0),.din(w_dff_A_vzR2OpQl1_0),.clk(gclk));
	jdff dff_A_f7dHFFwu5_0(.dout(w_dff_A_7SECabTb2_0),.din(w_dff_A_f7dHFFwu5_0),.clk(gclk));
	jdff dff_A_7SECabTb2_0(.dout(w_dff_A_TQVYDFq34_0),.din(w_dff_A_7SECabTb2_0),.clk(gclk));
	jdff dff_A_TQVYDFq34_0(.dout(w_dff_A_ZiNYr72P0_0),.din(w_dff_A_TQVYDFq34_0),.clk(gclk));
	jdff dff_A_ZiNYr72P0_0(.dout(w_dff_A_mwHNqASV5_0),.din(w_dff_A_ZiNYr72P0_0),.clk(gclk));
	jdff dff_A_mwHNqASV5_0(.dout(w_dff_A_5VBQfUnU4_0),.din(w_dff_A_mwHNqASV5_0),.clk(gclk));
	jdff dff_A_5VBQfUnU4_0(.dout(w_dff_A_WDBLBGzs7_0),.din(w_dff_A_5VBQfUnU4_0),.clk(gclk));
	jdff dff_A_WDBLBGzs7_0(.dout(w_dff_A_E6KjC8616_0),.din(w_dff_A_WDBLBGzs7_0),.clk(gclk));
	jdff dff_A_E6KjC8616_0(.dout(w_dff_A_cCK7Y65C8_0),.din(w_dff_A_E6KjC8616_0),.clk(gclk));
	jdff dff_A_cCK7Y65C8_0(.dout(w_dff_A_HYbqHw3Z4_0),.din(w_dff_A_cCK7Y65C8_0),.clk(gclk));
	jdff dff_A_HYbqHw3Z4_0(.dout(w_dff_A_9i4A78N81_0),.din(w_dff_A_HYbqHw3Z4_0),.clk(gclk));
	jdff dff_A_9i4A78N81_0(.dout(w_dff_A_gAQA6WhP8_0),.din(w_dff_A_9i4A78N81_0),.clk(gclk));
	jdff dff_A_gAQA6WhP8_0(.dout(w_dff_A_mBpUqUIy3_0),.din(w_dff_A_gAQA6WhP8_0),.clk(gclk));
	jdff dff_A_mBpUqUIy3_0(.dout(w_dff_A_E90cnU9I8_0),.din(w_dff_A_mBpUqUIy3_0),.clk(gclk));
	jdff dff_A_E90cnU9I8_0(.dout(w_dff_A_uzXj0SC12_0),.din(w_dff_A_E90cnU9I8_0),.clk(gclk));
	jdff dff_A_uzXj0SC12_0(.dout(w_dff_A_PRY3VpPV8_0),.din(w_dff_A_uzXj0SC12_0),.clk(gclk));
	jdff dff_A_PRY3VpPV8_0(.dout(w_dff_A_LzDIyGAn7_0),.din(w_dff_A_PRY3VpPV8_0),.clk(gclk));
	jdff dff_A_LzDIyGAn7_0(.dout(G438),.din(w_dff_A_LzDIyGAn7_0),.clk(gclk));
	jdff dff_A_GSYFA4ww3_1(.dout(w_dff_A_UCDwvfB98_0),.din(w_dff_A_GSYFA4ww3_1),.clk(gclk));
	jdff dff_A_UCDwvfB98_0(.dout(w_dff_A_Xwd1dn5f9_0),.din(w_dff_A_UCDwvfB98_0),.clk(gclk));
	jdff dff_A_Xwd1dn5f9_0(.dout(w_dff_A_EYxB8Lc47_0),.din(w_dff_A_Xwd1dn5f9_0),.clk(gclk));
	jdff dff_A_EYxB8Lc47_0(.dout(w_dff_A_xvxn9SEF2_0),.din(w_dff_A_EYxB8Lc47_0),.clk(gclk));
	jdff dff_A_xvxn9SEF2_0(.dout(w_dff_A_ivdgl1Ra8_0),.din(w_dff_A_xvxn9SEF2_0),.clk(gclk));
	jdff dff_A_ivdgl1Ra8_0(.dout(w_dff_A_gjSGCExO3_0),.din(w_dff_A_ivdgl1Ra8_0),.clk(gclk));
	jdff dff_A_gjSGCExO3_0(.dout(w_dff_A_7O4fyjTs4_0),.din(w_dff_A_gjSGCExO3_0),.clk(gclk));
	jdff dff_A_7O4fyjTs4_0(.dout(w_dff_A_RPIxa1pk0_0),.din(w_dff_A_7O4fyjTs4_0),.clk(gclk));
	jdff dff_A_RPIxa1pk0_0(.dout(w_dff_A_1WqGe35Z3_0),.din(w_dff_A_RPIxa1pk0_0),.clk(gclk));
	jdff dff_A_1WqGe35Z3_0(.dout(w_dff_A_UMCk5GSg1_0),.din(w_dff_A_1WqGe35Z3_0),.clk(gclk));
	jdff dff_A_UMCk5GSg1_0(.dout(w_dff_A_TJZAYtit9_0),.din(w_dff_A_UMCk5GSg1_0),.clk(gclk));
	jdff dff_A_TJZAYtit9_0(.dout(w_dff_A_nYJVWxya9_0),.din(w_dff_A_TJZAYtit9_0),.clk(gclk));
	jdff dff_A_nYJVWxya9_0(.dout(w_dff_A_mlj9TEEr2_0),.din(w_dff_A_nYJVWxya9_0),.clk(gclk));
	jdff dff_A_mlj9TEEr2_0(.dout(w_dff_A_q4Q1ISsF1_0),.din(w_dff_A_mlj9TEEr2_0),.clk(gclk));
	jdff dff_A_q4Q1ISsF1_0(.dout(w_dff_A_qNyI5hBV7_0),.din(w_dff_A_q4Q1ISsF1_0),.clk(gclk));
	jdff dff_A_qNyI5hBV7_0(.dout(w_dff_A_n0YcfmhI5_0),.din(w_dff_A_qNyI5hBV7_0),.clk(gclk));
	jdff dff_A_n0YcfmhI5_0(.dout(w_dff_A_yWCyAVIW2_0),.din(w_dff_A_n0YcfmhI5_0),.clk(gclk));
	jdff dff_A_yWCyAVIW2_0(.dout(w_dff_A_MAPhUM7N6_0),.din(w_dff_A_yWCyAVIW2_0),.clk(gclk));
	jdff dff_A_MAPhUM7N6_0(.dout(w_dff_A_8kmOKFZ74_0),.din(w_dff_A_MAPhUM7N6_0),.clk(gclk));
	jdff dff_A_8kmOKFZ74_0(.dout(w_dff_A_KRYGJYe34_0),.din(w_dff_A_8kmOKFZ74_0),.clk(gclk));
	jdff dff_A_KRYGJYe34_0(.dout(w_dff_A_UkVafpsX8_0),.din(w_dff_A_KRYGJYe34_0),.clk(gclk));
	jdff dff_A_UkVafpsX8_0(.dout(w_dff_A_pYGMXtPG0_0),.din(w_dff_A_UkVafpsX8_0),.clk(gclk));
	jdff dff_A_pYGMXtPG0_0(.dout(w_dff_A_qgOecMjz3_0),.din(w_dff_A_pYGMXtPG0_0),.clk(gclk));
	jdff dff_A_qgOecMjz3_0(.dout(w_dff_A_AbMDtzDF4_0),.din(w_dff_A_qgOecMjz3_0),.clk(gclk));
	jdff dff_A_AbMDtzDF4_0(.dout(w_dff_A_dOymBiyS4_0),.din(w_dff_A_AbMDtzDF4_0),.clk(gclk));
	jdff dff_A_dOymBiyS4_0(.dout(w_dff_A_5Bc3xjBw8_0),.din(w_dff_A_dOymBiyS4_0),.clk(gclk));
	jdff dff_A_5Bc3xjBw8_0(.dout(w_dff_A_7gN0jQnA7_0),.din(w_dff_A_5Bc3xjBw8_0),.clk(gclk));
	jdff dff_A_7gN0jQnA7_0(.dout(w_dff_A_8nqhAhPU0_0),.din(w_dff_A_7gN0jQnA7_0),.clk(gclk));
	jdff dff_A_8nqhAhPU0_0(.dout(w_dff_A_ukHPcTK93_0),.din(w_dff_A_8nqhAhPU0_0),.clk(gclk));
	jdff dff_A_ukHPcTK93_0(.dout(w_dff_A_yMfo0Kd35_0),.din(w_dff_A_ukHPcTK93_0),.clk(gclk));
	jdff dff_A_yMfo0Kd35_0(.dout(w_dff_A_620NMmt57_0),.din(w_dff_A_yMfo0Kd35_0),.clk(gclk));
	jdff dff_A_620NMmt57_0(.dout(w_dff_A_PsVygU4V6_0),.din(w_dff_A_620NMmt57_0),.clk(gclk));
	jdff dff_A_PsVygU4V6_0(.dout(w_dff_A_is0H3t9B5_0),.din(w_dff_A_PsVygU4V6_0),.clk(gclk));
	jdff dff_A_is0H3t9B5_0(.dout(w_dff_A_nB6wTG6c9_0),.din(w_dff_A_is0H3t9B5_0),.clk(gclk));
	jdff dff_A_nB6wTG6c9_0(.dout(w_dff_A_QLHHnaNR3_0),.din(w_dff_A_nB6wTG6c9_0),.clk(gclk));
	jdff dff_A_QLHHnaNR3_0(.dout(w_dff_A_rE57DQMO2_0),.din(w_dff_A_QLHHnaNR3_0),.clk(gclk));
	jdff dff_A_rE57DQMO2_0(.dout(w_dff_A_3wSZ1bML4_0),.din(w_dff_A_rE57DQMO2_0),.clk(gclk));
	jdff dff_A_3wSZ1bML4_0(.dout(w_dff_A_dljBLxcc5_0),.din(w_dff_A_3wSZ1bML4_0),.clk(gclk));
	jdff dff_A_dljBLxcc5_0(.dout(G496),.din(w_dff_A_dljBLxcc5_0),.clk(gclk));
	jdff dff_A_FBQkF7m74_1(.dout(w_dff_A_4fl1TdOT5_0),.din(w_dff_A_FBQkF7m74_1),.clk(gclk));
	jdff dff_A_4fl1TdOT5_0(.dout(w_dff_A_7cGDXaDb1_0),.din(w_dff_A_4fl1TdOT5_0),.clk(gclk));
	jdff dff_A_7cGDXaDb1_0(.dout(w_dff_A_IuCW8esC3_0),.din(w_dff_A_7cGDXaDb1_0),.clk(gclk));
	jdff dff_A_IuCW8esC3_0(.dout(w_dff_A_qb2SftNO3_0),.din(w_dff_A_IuCW8esC3_0),.clk(gclk));
	jdff dff_A_qb2SftNO3_0(.dout(w_dff_A_jf16ptjl6_0),.din(w_dff_A_qb2SftNO3_0),.clk(gclk));
	jdff dff_A_jf16ptjl6_0(.dout(w_dff_A_kXQcMjmI5_0),.din(w_dff_A_jf16ptjl6_0),.clk(gclk));
	jdff dff_A_kXQcMjmI5_0(.dout(w_dff_A_MC9AYpHi9_0),.din(w_dff_A_kXQcMjmI5_0),.clk(gclk));
	jdff dff_A_MC9AYpHi9_0(.dout(w_dff_A_FU5lvZYK5_0),.din(w_dff_A_MC9AYpHi9_0),.clk(gclk));
	jdff dff_A_FU5lvZYK5_0(.dout(w_dff_A_G2AYCFir6_0),.din(w_dff_A_FU5lvZYK5_0),.clk(gclk));
	jdff dff_A_G2AYCFir6_0(.dout(w_dff_A_Rj8jANqp8_0),.din(w_dff_A_G2AYCFir6_0),.clk(gclk));
	jdff dff_A_Rj8jANqp8_0(.dout(w_dff_A_ZwqwohQk9_0),.din(w_dff_A_Rj8jANqp8_0),.clk(gclk));
	jdff dff_A_ZwqwohQk9_0(.dout(w_dff_A_JU4alewb1_0),.din(w_dff_A_ZwqwohQk9_0),.clk(gclk));
	jdff dff_A_JU4alewb1_0(.dout(w_dff_A_G1mKw5Sf3_0),.din(w_dff_A_JU4alewb1_0),.clk(gclk));
	jdff dff_A_G1mKw5Sf3_0(.dout(w_dff_A_7F9hztQZ9_0),.din(w_dff_A_G1mKw5Sf3_0),.clk(gclk));
	jdff dff_A_7F9hztQZ9_0(.dout(w_dff_A_Cm4q8UEB4_0),.din(w_dff_A_7F9hztQZ9_0),.clk(gclk));
	jdff dff_A_Cm4q8UEB4_0(.dout(w_dff_A_XTssvDHE6_0),.din(w_dff_A_Cm4q8UEB4_0),.clk(gclk));
	jdff dff_A_XTssvDHE6_0(.dout(w_dff_A_OA9L6giI5_0),.din(w_dff_A_XTssvDHE6_0),.clk(gclk));
	jdff dff_A_OA9L6giI5_0(.dout(w_dff_A_sgdFz96H0_0),.din(w_dff_A_OA9L6giI5_0),.clk(gclk));
	jdff dff_A_sgdFz96H0_0(.dout(w_dff_A_eoSjGsmr2_0),.din(w_dff_A_sgdFz96H0_0),.clk(gclk));
	jdff dff_A_eoSjGsmr2_0(.dout(w_dff_A_0of6W2W81_0),.din(w_dff_A_eoSjGsmr2_0),.clk(gclk));
	jdff dff_A_0of6W2W81_0(.dout(w_dff_A_pPwfNzyI9_0),.din(w_dff_A_0of6W2W81_0),.clk(gclk));
	jdff dff_A_pPwfNzyI9_0(.dout(w_dff_A_g3FQySvx7_0),.din(w_dff_A_pPwfNzyI9_0),.clk(gclk));
	jdff dff_A_g3FQySvx7_0(.dout(w_dff_A_da3Hoaiz7_0),.din(w_dff_A_g3FQySvx7_0),.clk(gclk));
	jdff dff_A_da3Hoaiz7_0(.dout(w_dff_A_DLICkPhl6_0),.din(w_dff_A_da3Hoaiz7_0),.clk(gclk));
	jdff dff_A_DLICkPhl6_0(.dout(w_dff_A_q5vmGSpN0_0),.din(w_dff_A_DLICkPhl6_0),.clk(gclk));
	jdff dff_A_q5vmGSpN0_0(.dout(w_dff_A_QgCp5rPq4_0),.din(w_dff_A_q5vmGSpN0_0),.clk(gclk));
	jdff dff_A_QgCp5rPq4_0(.dout(w_dff_A_0q3xGcbg7_0),.din(w_dff_A_QgCp5rPq4_0),.clk(gclk));
	jdff dff_A_0q3xGcbg7_0(.dout(w_dff_A_7mGhgGiY8_0),.din(w_dff_A_0q3xGcbg7_0),.clk(gclk));
	jdff dff_A_7mGhgGiY8_0(.dout(w_dff_A_wGuxlG9W7_0),.din(w_dff_A_7mGhgGiY8_0),.clk(gclk));
	jdff dff_A_wGuxlG9W7_0(.dout(w_dff_A_iXikGm2I1_0),.din(w_dff_A_wGuxlG9W7_0),.clk(gclk));
	jdff dff_A_iXikGm2I1_0(.dout(w_dff_A_CrMsD6NM6_0),.din(w_dff_A_iXikGm2I1_0),.clk(gclk));
	jdff dff_A_CrMsD6NM6_0(.dout(w_dff_A_fYF7LZEe3_0),.din(w_dff_A_CrMsD6NM6_0),.clk(gclk));
	jdff dff_A_fYF7LZEe3_0(.dout(w_dff_A_FXQNcGJm1_0),.din(w_dff_A_fYF7LZEe3_0),.clk(gclk));
	jdff dff_A_FXQNcGJm1_0(.dout(w_dff_A_OAluJ2xm7_0),.din(w_dff_A_FXQNcGJm1_0),.clk(gclk));
	jdff dff_A_OAluJ2xm7_0(.dout(w_dff_A_jZ7X0diM9_0),.din(w_dff_A_OAluJ2xm7_0),.clk(gclk));
	jdff dff_A_jZ7X0diM9_0(.dout(w_dff_A_Rnd37Xd55_0),.din(w_dff_A_jZ7X0diM9_0),.clk(gclk));
	jdff dff_A_Rnd37Xd55_0(.dout(w_dff_A_cFBAvjoj2_0),.din(w_dff_A_Rnd37Xd55_0),.clk(gclk));
	jdff dff_A_cFBAvjoj2_0(.dout(w_dff_A_pDcmaUo15_0),.din(w_dff_A_cFBAvjoj2_0),.clk(gclk));
	jdff dff_A_pDcmaUo15_0(.dout(G494),.din(w_dff_A_pDcmaUo15_0),.clk(gclk));
	jdff dff_A_YfYhlcZP8_1(.dout(w_dff_A_y2t7sUPu6_0),.din(w_dff_A_YfYhlcZP8_1),.clk(gclk));
	jdff dff_A_y2t7sUPu6_0(.dout(w_dff_A_42e3Nu0u0_0),.din(w_dff_A_y2t7sUPu6_0),.clk(gclk));
	jdff dff_A_42e3Nu0u0_0(.dout(w_dff_A_cMCizrwn5_0),.din(w_dff_A_42e3Nu0u0_0),.clk(gclk));
	jdff dff_A_cMCizrwn5_0(.dout(w_dff_A_czJjS1ol4_0),.din(w_dff_A_cMCizrwn5_0),.clk(gclk));
	jdff dff_A_czJjS1ol4_0(.dout(w_dff_A_D8RA6Ehk1_0),.din(w_dff_A_czJjS1ol4_0),.clk(gclk));
	jdff dff_A_D8RA6Ehk1_0(.dout(w_dff_A_CGgXfMgQ3_0),.din(w_dff_A_D8RA6Ehk1_0),.clk(gclk));
	jdff dff_A_CGgXfMgQ3_0(.dout(w_dff_A_1z2gackJ6_0),.din(w_dff_A_CGgXfMgQ3_0),.clk(gclk));
	jdff dff_A_1z2gackJ6_0(.dout(w_dff_A_FzQssm2F1_0),.din(w_dff_A_1z2gackJ6_0),.clk(gclk));
	jdff dff_A_FzQssm2F1_0(.dout(w_dff_A_jOeeUuAC8_0),.din(w_dff_A_FzQssm2F1_0),.clk(gclk));
	jdff dff_A_jOeeUuAC8_0(.dout(w_dff_A_Nzm3wD5c9_0),.din(w_dff_A_jOeeUuAC8_0),.clk(gclk));
	jdff dff_A_Nzm3wD5c9_0(.dout(w_dff_A_aspOhlAV4_0),.din(w_dff_A_Nzm3wD5c9_0),.clk(gclk));
	jdff dff_A_aspOhlAV4_0(.dout(w_dff_A_gRwurW9b1_0),.din(w_dff_A_aspOhlAV4_0),.clk(gclk));
	jdff dff_A_gRwurW9b1_0(.dout(w_dff_A_C1R14Pgn4_0),.din(w_dff_A_gRwurW9b1_0),.clk(gclk));
	jdff dff_A_C1R14Pgn4_0(.dout(w_dff_A_zOkywjSZ1_0),.din(w_dff_A_C1R14Pgn4_0),.clk(gclk));
	jdff dff_A_zOkywjSZ1_0(.dout(w_dff_A_6ITAj4yy4_0),.din(w_dff_A_zOkywjSZ1_0),.clk(gclk));
	jdff dff_A_6ITAj4yy4_0(.dout(w_dff_A_Ny8w7pGi1_0),.din(w_dff_A_6ITAj4yy4_0),.clk(gclk));
	jdff dff_A_Ny8w7pGi1_0(.dout(w_dff_A_tgvazPQr9_0),.din(w_dff_A_Ny8w7pGi1_0),.clk(gclk));
	jdff dff_A_tgvazPQr9_0(.dout(w_dff_A_XssZaBn06_0),.din(w_dff_A_tgvazPQr9_0),.clk(gclk));
	jdff dff_A_XssZaBn06_0(.dout(w_dff_A_HqNCbgsy7_0),.din(w_dff_A_XssZaBn06_0),.clk(gclk));
	jdff dff_A_HqNCbgsy7_0(.dout(w_dff_A_gmSWy4kD0_0),.din(w_dff_A_HqNCbgsy7_0),.clk(gclk));
	jdff dff_A_gmSWy4kD0_0(.dout(w_dff_A_NVJbwkiI8_0),.din(w_dff_A_gmSWy4kD0_0),.clk(gclk));
	jdff dff_A_NVJbwkiI8_0(.dout(w_dff_A_30yshV7O7_0),.din(w_dff_A_NVJbwkiI8_0),.clk(gclk));
	jdff dff_A_30yshV7O7_0(.dout(w_dff_A_ijbGCjpS9_0),.din(w_dff_A_30yshV7O7_0),.clk(gclk));
	jdff dff_A_ijbGCjpS9_0(.dout(w_dff_A_PyzddnWi8_0),.din(w_dff_A_ijbGCjpS9_0),.clk(gclk));
	jdff dff_A_PyzddnWi8_0(.dout(w_dff_A_SQa6CXCT7_0),.din(w_dff_A_PyzddnWi8_0),.clk(gclk));
	jdff dff_A_SQa6CXCT7_0(.dout(w_dff_A_BeRNFGHW5_0),.din(w_dff_A_SQa6CXCT7_0),.clk(gclk));
	jdff dff_A_BeRNFGHW5_0(.dout(w_dff_A_MAmaBNb15_0),.din(w_dff_A_BeRNFGHW5_0),.clk(gclk));
	jdff dff_A_MAmaBNb15_0(.dout(w_dff_A_s6PzIUkA3_0),.din(w_dff_A_MAmaBNb15_0),.clk(gclk));
	jdff dff_A_s6PzIUkA3_0(.dout(w_dff_A_peaBLIjd9_0),.din(w_dff_A_s6PzIUkA3_0),.clk(gclk));
	jdff dff_A_peaBLIjd9_0(.dout(w_dff_A_ZpCw35dE1_0),.din(w_dff_A_peaBLIjd9_0),.clk(gclk));
	jdff dff_A_ZpCw35dE1_0(.dout(w_dff_A_FZr2HDck5_0),.din(w_dff_A_ZpCw35dE1_0),.clk(gclk));
	jdff dff_A_FZr2HDck5_0(.dout(w_dff_A_g3Sec77k9_0),.din(w_dff_A_FZr2HDck5_0),.clk(gclk));
	jdff dff_A_g3Sec77k9_0(.dout(w_dff_A_bjRPVOzQ3_0),.din(w_dff_A_g3Sec77k9_0),.clk(gclk));
	jdff dff_A_bjRPVOzQ3_0(.dout(w_dff_A_cEZkXk7w0_0),.din(w_dff_A_bjRPVOzQ3_0),.clk(gclk));
	jdff dff_A_cEZkXk7w0_0(.dout(w_dff_A_cs3xDGtC2_0),.din(w_dff_A_cEZkXk7w0_0),.clk(gclk));
	jdff dff_A_cs3xDGtC2_0(.dout(w_dff_A_gUFwK4nh4_0),.din(w_dff_A_cs3xDGtC2_0),.clk(gclk));
	jdff dff_A_gUFwK4nh4_0(.dout(w_dff_A_ir4bMUJO9_0),.din(w_dff_A_gUFwK4nh4_0),.clk(gclk));
	jdff dff_A_ir4bMUJO9_0(.dout(w_dff_A_17fmTVMQ1_0),.din(w_dff_A_ir4bMUJO9_0),.clk(gclk));
	jdff dff_A_17fmTVMQ1_0(.dout(G492),.din(w_dff_A_17fmTVMQ1_0),.clk(gclk));
	jdff dff_A_tzhGpJqn6_1(.dout(w_dff_A_mfbW9HGd7_0),.din(w_dff_A_tzhGpJqn6_1),.clk(gclk));
	jdff dff_A_mfbW9HGd7_0(.dout(w_dff_A_1aixFJQK1_0),.din(w_dff_A_mfbW9HGd7_0),.clk(gclk));
	jdff dff_A_1aixFJQK1_0(.dout(w_dff_A_qngvwCEc1_0),.din(w_dff_A_1aixFJQK1_0),.clk(gclk));
	jdff dff_A_qngvwCEc1_0(.dout(w_dff_A_sN0Z2cua7_0),.din(w_dff_A_qngvwCEc1_0),.clk(gclk));
	jdff dff_A_sN0Z2cua7_0(.dout(w_dff_A_dYAtbBlm4_0),.din(w_dff_A_sN0Z2cua7_0),.clk(gclk));
	jdff dff_A_dYAtbBlm4_0(.dout(w_dff_A_fbKhrtWB5_0),.din(w_dff_A_dYAtbBlm4_0),.clk(gclk));
	jdff dff_A_fbKhrtWB5_0(.dout(w_dff_A_mHaWUr5G7_0),.din(w_dff_A_fbKhrtWB5_0),.clk(gclk));
	jdff dff_A_mHaWUr5G7_0(.dout(w_dff_A_RTmYkP9I4_0),.din(w_dff_A_mHaWUr5G7_0),.clk(gclk));
	jdff dff_A_RTmYkP9I4_0(.dout(w_dff_A_wmlkjIvu1_0),.din(w_dff_A_RTmYkP9I4_0),.clk(gclk));
	jdff dff_A_wmlkjIvu1_0(.dout(w_dff_A_NNIsZJ2s8_0),.din(w_dff_A_wmlkjIvu1_0),.clk(gclk));
	jdff dff_A_NNIsZJ2s8_0(.dout(w_dff_A_PHJ6s1f81_0),.din(w_dff_A_NNIsZJ2s8_0),.clk(gclk));
	jdff dff_A_PHJ6s1f81_0(.dout(w_dff_A_ymaG0ljj7_0),.din(w_dff_A_PHJ6s1f81_0),.clk(gclk));
	jdff dff_A_ymaG0ljj7_0(.dout(w_dff_A_ffOwCtHh2_0),.din(w_dff_A_ymaG0ljj7_0),.clk(gclk));
	jdff dff_A_ffOwCtHh2_0(.dout(w_dff_A_U9vRYRLH2_0),.din(w_dff_A_ffOwCtHh2_0),.clk(gclk));
	jdff dff_A_U9vRYRLH2_0(.dout(w_dff_A_eeKvm5xK3_0),.din(w_dff_A_U9vRYRLH2_0),.clk(gclk));
	jdff dff_A_eeKvm5xK3_0(.dout(w_dff_A_gBq5XAWp6_0),.din(w_dff_A_eeKvm5xK3_0),.clk(gclk));
	jdff dff_A_gBq5XAWp6_0(.dout(w_dff_A_6W7CEBAW1_0),.din(w_dff_A_gBq5XAWp6_0),.clk(gclk));
	jdff dff_A_6W7CEBAW1_0(.dout(w_dff_A_Xqke8QnJ7_0),.din(w_dff_A_6W7CEBAW1_0),.clk(gclk));
	jdff dff_A_Xqke8QnJ7_0(.dout(w_dff_A_wzcgwqhc2_0),.din(w_dff_A_Xqke8QnJ7_0),.clk(gclk));
	jdff dff_A_wzcgwqhc2_0(.dout(w_dff_A_jfkQr8Wy8_0),.din(w_dff_A_wzcgwqhc2_0),.clk(gclk));
	jdff dff_A_jfkQr8Wy8_0(.dout(w_dff_A_jHi9cTO57_0),.din(w_dff_A_jfkQr8Wy8_0),.clk(gclk));
	jdff dff_A_jHi9cTO57_0(.dout(w_dff_A_hgLnWIsW6_0),.din(w_dff_A_jHi9cTO57_0),.clk(gclk));
	jdff dff_A_hgLnWIsW6_0(.dout(w_dff_A_6POL6XvD0_0),.din(w_dff_A_hgLnWIsW6_0),.clk(gclk));
	jdff dff_A_6POL6XvD0_0(.dout(w_dff_A_zIosLDnn4_0),.din(w_dff_A_6POL6XvD0_0),.clk(gclk));
	jdff dff_A_zIosLDnn4_0(.dout(w_dff_A_grINay6F3_0),.din(w_dff_A_zIosLDnn4_0),.clk(gclk));
	jdff dff_A_grINay6F3_0(.dout(w_dff_A_elW4YhXo0_0),.din(w_dff_A_grINay6F3_0),.clk(gclk));
	jdff dff_A_elW4YhXo0_0(.dout(w_dff_A_M9crSgu92_0),.din(w_dff_A_elW4YhXo0_0),.clk(gclk));
	jdff dff_A_M9crSgu92_0(.dout(w_dff_A_PnGGQqeE7_0),.din(w_dff_A_M9crSgu92_0),.clk(gclk));
	jdff dff_A_PnGGQqeE7_0(.dout(w_dff_A_0EzfcwUL8_0),.din(w_dff_A_PnGGQqeE7_0),.clk(gclk));
	jdff dff_A_0EzfcwUL8_0(.dout(w_dff_A_uW7Lqxgf2_0),.din(w_dff_A_0EzfcwUL8_0),.clk(gclk));
	jdff dff_A_uW7Lqxgf2_0(.dout(w_dff_A_eNYN0uf75_0),.din(w_dff_A_uW7Lqxgf2_0),.clk(gclk));
	jdff dff_A_eNYN0uf75_0(.dout(w_dff_A_TrpB85Je6_0),.din(w_dff_A_eNYN0uf75_0),.clk(gclk));
	jdff dff_A_TrpB85Je6_0(.dout(w_dff_A_EdtrBZVM6_0),.din(w_dff_A_TrpB85Je6_0),.clk(gclk));
	jdff dff_A_EdtrBZVM6_0(.dout(w_dff_A_9DTXmvba8_0),.din(w_dff_A_EdtrBZVM6_0),.clk(gclk));
	jdff dff_A_9DTXmvba8_0(.dout(w_dff_A_Q8ifz1Tj2_0),.din(w_dff_A_9DTXmvba8_0),.clk(gclk));
	jdff dff_A_Q8ifz1Tj2_0(.dout(w_dff_A_kftT5qGG1_0),.din(w_dff_A_Q8ifz1Tj2_0),.clk(gclk));
	jdff dff_A_kftT5qGG1_0(.dout(w_dff_A_M7JwIvUK5_0),.din(w_dff_A_kftT5qGG1_0),.clk(gclk));
	jdff dff_A_M7JwIvUK5_0(.dout(w_dff_A_YJ2LTApK3_0),.din(w_dff_A_M7JwIvUK5_0),.clk(gclk));
	jdff dff_A_YJ2LTApK3_0(.dout(G490),.din(w_dff_A_YJ2LTApK3_0),.clk(gclk));
	jdff dff_A_Wdw6GYOZ5_1(.dout(w_dff_A_c6AG1F5e9_0),.din(w_dff_A_Wdw6GYOZ5_1),.clk(gclk));
	jdff dff_A_c6AG1F5e9_0(.dout(w_dff_A_FPU5Fyob7_0),.din(w_dff_A_c6AG1F5e9_0),.clk(gclk));
	jdff dff_A_FPU5Fyob7_0(.dout(w_dff_A_pZ0c0waE9_0),.din(w_dff_A_FPU5Fyob7_0),.clk(gclk));
	jdff dff_A_pZ0c0waE9_0(.dout(w_dff_A_BpMi0wnW0_0),.din(w_dff_A_pZ0c0waE9_0),.clk(gclk));
	jdff dff_A_BpMi0wnW0_0(.dout(w_dff_A_tzZuctiQ8_0),.din(w_dff_A_BpMi0wnW0_0),.clk(gclk));
	jdff dff_A_tzZuctiQ8_0(.dout(w_dff_A_j3PzZWYR8_0),.din(w_dff_A_tzZuctiQ8_0),.clk(gclk));
	jdff dff_A_j3PzZWYR8_0(.dout(w_dff_A_cYq2OVgH2_0),.din(w_dff_A_j3PzZWYR8_0),.clk(gclk));
	jdff dff_A_cYq2OVgH2_0(.dout(w_dff_A_h4eQE88U5_0),.din(w_dff_A_cYq2OVgH2_0),.clk(gclk));
	jdff dff_A_h4eQE88U5_0(.dout(w_dff_A_bLkwVTOO0_0),.din(w_dff_A_h4eQE88U5_0),.clk(gclk));
	jdff dff_A_bLkwVTOO0_0(.dout(w_dff_A_Wo661W4s3_0),.din(w_dff_A_bLkwVTOO0_0),.clk(gclk));
	jdff dff_A_Wo661W4s3_0(.dout(w_dff_A_maEm4jcD8_0),.din(w_dff_A_Wo661W4s3_0),.clk(gclk));
	jdff dff_A_maEm4jcD8_0(.dout(w_dff_A_5zrgfV6c4_0),.din(w_dff_A_maEm4jcD8_0),.clk(gclk));
	jdff dff_A_5zrgfV6c4_0(.dout(w_dff_A_IU2ndIBE5_0),.din(w_dff_A_5zrgfV6c4_0),.clk(gclk));
	jdff dff_A_IU2ndIBE5_0(.dout(w_dff_A_UjrdH04g4_0),.din(w_dff_A_IU2ndIBE5_0),.clk(gclk));
	jdff dff_A_UjrdH04g4_0(.dout(w_dff_A_7Zzqu8E70_0),.din(w_dff_A_UjrdH04g4_0),.clk(gclk));
	jdff dff_A_7Zzqu8E70_0(.dout(w_dff_A_9B2wsbLX2_0),.din(w_dff_A_7Zzqu8E70_0),.clk(gclk));
	jdff dff_A_9B2wsbLX2_0(.dout(w_dff_A_TunQH81q8_0),.din(w_dff_A_9B2wsbLX2_0),.clk(gclk));
	jdff dff_A_TunQH81q8_0(.dout(w_dff_A_vGfmp3lQ8_0),.din(w_dff_A_TunQH81q8_0),.clk(gclk));
	jdff dff_A_vGfmp3lQ8_0(.dout(w_dff_A_UM1XqdFl8_0),.din(w_dff_A_vGfmp3lQ8_0),.clk(gclk));
	jdff dff_A_UM1XqdFl8_0(.dout(w_dff_A_1TsuALWQ3_0),.din(w_dff_A_UM1XqdFl8_0),.clk(gclk));
	jdff dff_A_1TsuALWQ3_0(.dout(w_dff_A_wqoUCg256_0),.din(w_dff_A_1TsuALWQ3_0),.clk(gclk));
	jdff dff_A_wqoUCg256_0(.dout(w_dff_A_9Gj66eJi7_0),.din(w_dff_A_wqoUCg256_0),.clk(gclk));
	jdff dff_A_9Gj66eJi7_0(.dout(w_dff_A_r7DmmLKM8_0),.din(w_dff_A_9Gj66eJi7_0),.clk(gclk));
	jdff dff_A_r7DmmLKM8_0(.dout(w_dff_A_gJFqMbm18_0),.din(w_dff_A_r7DmmLKM8_0),.clk(gclk));
	jdff dff_A_gJFqMbm18_0(.dout(w_dff_A_gBj7IIKO4_0),.din(w_dff_A_gJFqMbm18_0),.clk(gclk));
	jdff dff_A_gBj7IIKO4_0(.dout(w_dff_A_GiRPAt5R9_0),.din(w_dff_A_gBj7IIKO4_0),.clk(gclk));
	jdff dff_A_GiRPAt5R9_0(.dout(w_dff_A_UJLviwNg7_0),.din(w_dff_A_GiRPAt5R9_0),.clk(gclk));
	jdff dff_A_UJLviwNg7_0(.dout(w_dff_A_mYuPKgWy0_0),.din(w_dff_A_UJLviwNg7_0),.clk(gclk));
	jdff dff_A_mYuPKgWy0_0(.dout(w_dff_A_i60DtdbK3_0),.din(w_dff_A_mYuPKgWy0_0),.clk(gclk));
	jdff dff_A_i60DtdbK3_0(.dout(w_dff_A_JzBR7V1g5_0),.din(w_dff_A_i60DtdbK3_0),.clk(gclk));
	jdff dff_A_JzBR7V1g5_0(.dout(w_dff_A_wC6rJ1v25_0),.din(w_dff_A_JzBR7V1g5_0),.clk(gclk));
	jdff dff_A_wC6rJ1v25_0(.dout(w_dff_A_tG6wXf507_0),.din(w_dff_A_wC6rJ1v25_0),.clk(gclk));
	jdff dff_A_tG6wXf507_0(.dout(w_dff_A_9F7I295l7_0),.din(w_dff_A_tG6wXf507_0),.clk(gclk));
	jdff dff_A_9F7I295l7_0(.dout(w_dff_A_oqspcb7P1_0),.din(w_dff_A_9F7I295l7_0),.clk(gclk));
	jdff dff_A_oqspcb7P1_0(.dout(w_dff_A_L9RCra828_0),.din(w_dff_A_oqspcb7P1_0),.clk(gclk));
	jdff dff_A_L9RCra828_0(.dout(w_dff_A_Eu6vmsRB4_0),.din(w_dff_A_L9RCra828_0),.clk(gclk));
	jdff dff_A_Eu6vmsRB4_0(.dout(w_dff_A_NRpPcXoQ0_0),.din(w_dff_A_Eu6vmsRB4_0),.clk(gclk));
	jdff dff_A_NRpPcXoQ0_0(.dout(w_dff_A_QJOnwk5p7_0),.din(w_dff_A_NRpPcXoQ0_0),.clk(gclk));
	jdff dff_A_QJOnwk5p7_0(.dout(G488),.din(w_dff_A_QJOnwk5p7_0),.clk(gclk));
	jdff dff_A_u6wSNtT59_1(.dout(w_dff_A_ogARaZaQ0_0),.din(w_dff_A_u6wSNtT59_1),.clk(gclk));
	jdff dff_A_ogARaZaQ0_0(.dout(w_dff_A_rSFo8fLN2_0),.din(w_dff_A_ogARaZaQ0_0),.clk(gclk));
	jdff dff_A_rSFo8fLN2_0(.dout(w_dff_A_4QneGP4k5_0),.din(w_dff_A_rSFo8fLN2_0),.clk(gclk));
	jdff dff_A_4QneGP4k5_0(.dout(w_dff_A_PPMO63dC6_0),.din(w_dff_A_4QneGP4k5_0),.clk(gclk));
	jdff dff_A_PPMO63dC6_0(.dout(w_dff_A_ZXuj7kq30_0),.din(w_dff_A_PPMO63dC6_0),.clk(gclk));
	jdff dff_A_ZXuj7kq30_0(.dout(w_dff_A_G8RgCPor4_0),.din(w_dff_A_ZXuj7kq30_0),.clk(gclk));
	jdff dff_A_G8RgCPor4_0(.dout(w_dff_A_u6fNNzz82_0),.din(w_dff_A_G8RgCPor4_0),.clk(gclk));
	jdff dff_A_u6fNNzz82_0(.dout(w_dff_A_kwW7jrr82_0),.din(w_dff_A_u6fNNzz82_0),.clk(gclk));
	jdff dff_A_kwW7jrr82_0(.dout(w_dff_A_kWwQTSAX4_0),.din(w_dff_A_kwW7jrr82_0),.clk(gclk));
	jdff dff_A_kWwQTSAX4_0(.dout(w_dff_A_XwJzvhkQ0_0),.din(w_dff_A_kWwQTSAX4_0),.clk(gclk));
	jdff dff_A_XwJzvhkQ0_0(.dout(w_dff_A_gIFPiC2d0_0),.din(w_dff_A_XwJzvhkQ0_0),.clk(gclk));
	jdff dff_A_gIFPiC2d0_0(.dout(w_dff_A_vHNiVTO56_0),.din(w_dff_A_gIFPiC2d0_0),.clk(gclk));
	jdff dff_A_vHNiVTO56_0(.dout(w_dff_A_9Jol0tfA5_0),.din(w_dff_A_vHNiVTO56_0),.clk(gclk));
	jdff dff_A_9Jol0tfA5_0(.dout(w_dff_A_OKwI49SD0_0),.din(w_dff_A_9Jol0tfA5_0),.clk(gclk));
	jdff dff_A_OKwI49SD0_0(.dout(w_dff_A_sxeuXXAK1_0),.din(w_dff_A_OKwI49SD0_0),.clk(gclk));
	jdff dff_A_sxeuXXAK1_0(.dout(w_dff_A_R2KZCmJI7_0),.din(w_dff_A_sxeuXXAK1_0),.clk(gclk));
	jdff dff_A_R2KZCmJI7_0(.dout(w_dff_A_SY1HHCyC5_0),.din(w_dff_A_R2KZCmJI7_0),.clk(gclk));
	jdff dff_A_SY1HHCyC5_0(.dout(w_dff_A_JMwCNNkM2_0),.din(w_dff_A_SY1HHCyC5_0),.clk(gclk));
	jdff dff_A_JMwCNNkM2_0(.dout(w_dff_A_72IGDjn84_0),.din(w_dff_A_JMwCNNkM2_0),.clk(gclk));
	jdff dff_A_72IGDjn84_0(.dout(w_dff_A_LE4dsog42_0),.din(w_dff_A_72IGDjn84_0),.clk(gclk));
	jdff dff_A_LE4dsog42_0(.dout(w_dff_A_69ClauPI3_0),.din(w_dff_A_LE4dsog42_0),.clk(gclk));
	jdff dff_A_69ClauPI3_0(.dout(w_dff_A_gfnNGYZI6_0),.din(w_dff_A_69ClauPI3_0),.clk(gclk));
	jdff dff_A_gfnNGYZI6_0(.dout(w_dff_A_BWridLWQ5_0),.din(w_dff_A_gfnNGYZI6_0),.clk(gclk));
	jdff dff_A_BWridLWQ5_0(.dout(w_dff_A_s3H1Qh1D8_0),.din(w_dff_A_BWridLWQ5_0),.clk(gclk));
	jdff dff_A_s3H1Qh1D8_0(.dout(w_dff_A_Gfz1pEMI3_0),.din(w_dff_A_s3H1Qh1D8_0),.clk(gclk));
	jdff dff_A_Gfz1pEMI3_0(.dout(w_dff_A_RdMaJqxI6_0),.din(w_dff_A_Gfz1pEMI3_0),.clk(gclk));
	jdff dff_A_RdMaJqxI6_0(.dout(w_dff_A_MyygLSgm8_0),.din(w_dff_A_RdMaJqxI6_0),.clk(gclk));
	jdff dff_A_MyygLSgm8_0(.dout(w_dff_A_X1f1yfy10_0),.din(w_dff_A_MyygLSgm8_0),.clk(gclk));
	jdff dff_A_X1f1yfy10_0(.dout(w_dff_A_Z68Fy68m6_0),.din(w_dff_A_X1f1yfy10_0),.clk(gclk));
	jdff dff_A_Z68Fy68m6_0(.dout(w_dff_A_B9lpOEDx3_0),.din(w_dff_A_Z68Fy68m6_0),.clk(gclk));
	jdff dff_A_B9lpOEDx3_0(.dout(w_dff_A_EwgDJfKq0_0),.din(w_dff_A_B9lpOEDx3_0),.clk(gclk));
	jdff dff_A_EwgDJfKq0_0(.dout(w_dff_A_v9Ttm6UF0_0),.din(w_dff_A_EwgDJfKq0_0),.clk(gclk));
	jdff dff_A_v9Ttm6UF0_0(.dout(w_dff_A_PiUU62Jp7_0),.din(w_dff_A_v9Ttm6UF0_0),.clk(gclk));
	jdff dff_A_PiUU62Jp7_0(.dout(w_dff_A_caZpPZUH7_0),.din(w_dff_A_PiUU62Jp7_0),.clk(gclk));
	jdff dff_A_caZpPZUH7_0(.dout(w_dff_A_SSOOoQON7_0),.din(w_dff_A_caZpPZUH7_0),.clk(gclk));
	jdff dff_A_SSOOoQON7_0(.dout(w_dff_A_2AzrEH9r2_0),.din(w_dff_A_SSOOoQON7_0),.clk(gclk));
	jdff dff_A_2AzrEH9r2_0(.dout(w_dff_A_tEgdZ2YH3_0),.din(w_dff_A_2AzrEH9r2_0),.clk(gclk));
	jdff dff_A_tEgdZ2YH3_0(.dout(w_dff_A_FEckNR5b8_0),.din(w_dff_A_tEgdZ2YH3_0),.clk(gclk));
	jdff dff_A_FEckNR5b8_0(.dout(G486),.din(w_dff_A_FEckNR5b8_0),.clk(gclk));
	jdff dff_A_PWRWabNi9_1(.dout(w_dff_A_lgt7miUz1_0),.din(w_dff_A_PWRWabNi9_1),.clk(gclk));
	jdff dff_A_lgt7miUz1_0(.dout(w_dff_A_EoRT4ScD9_0),.din(w_dff_A_lgt7miUz1_0),.clk(gclk));
	jdff dff_A_EoRT4ScD9_0(.dout(w_dff_A_ztQ7zwNs6_0),.din(w_dff_A_EoRT4ScD9_0),.clk(gclk));
	jdff dff_A_ztQ7zwNs6_0(.dout(w_dff_A_yf8i2mg22_0),.din(w_dff_A_ztQ7zwNs6_0),.clk(gclk));
	jdff dff_A_yf8i2mg22_0(.dout(w_dff_A_k5GE9RK50_0),.din(w_dff_A_yf8i2mg22_0),.clk(gclk));
	jdff dff_A_k5GE9RK50_0(.dout(w_dff_A_jIOXscPi0_0),.din(w_dff_A_k5GE9RK50_0),.clk(gclk));
	jdff dff_A_jIOXscPi0_0(.dout(w_dff_A_jypcoECY8_0),.din(w_dff_A_jIOXscPi0_0),.clk(gclk));
	jdff dff_A_jypcoECY8_0(.dout(w_dff_A_DZ1OtZQ91_0),.din(w_dff_A_jypcoECY8_0),.clk(gclk));
	jdff dff_A_DZ1OtZQ91_0(.dout(w_dff_A_Gtz2kCmo4_0),.din(w_dff_A_DZ1OtZQ91_0),.clk(gclk));
	jdff dff_A_Gtz2kCmo4_0(.dout(w_dff_A_FLBYrJ0w6_0),.din(w_dff_A_Gtz2kCmo4_0),.clk(gclk));
	jdff dff_A_FLBYrJ0w6_0(.dout(w_dff_A_I2Tvambw9_0),.din(w_dff_A_FLBYrJ0w6_0),.clk(gclk));
	jdff dff_A_I2Tvambw9_0(.dout(w_dff_A_8zX5rKx91_0),.din(w_dff_A_I2Tvambw9_0),.clk(gclk));
	jdff dff_A_8zX5rKx91_0(.dout(w_dff_A_xROupiks4_0),.din(w_dff_A_8zX5rKx91_0),.clk(gclk));
	jdff dff_A_xROupiks4_0(.dout(w_dff_A_lZXXkAYH2_0),.din(w_dff_A_xROupiks4_0),.clk(gclk));
	jdff dff_A_lZXXkAYH2_0(.dout(w_dff_A_skHUHohJ2_0),.din(w_dff_A_lZXXkAYH2_0),.clk(gclk));
	jdff dff_A_skHUHohJ2_0(.dout(w_dff_A_SPGAQ09S7_0),.din(w_dff_A_skHUHohJ2_0),.clk(gclk));
	jdff dff_A_SPGAQ09S7_0(.dout(w_dff_A_RyJSeOuc3_0),.din(w_dff_A_SPGAQ09S7_0),.clk(gclk));
	jdff dff_A_RyJSeOuc3_0(.dout(w_dff_A_9oAWMnwV5_0),.din(w_dff_A_RyJSeOuc3_0),.clk(gclk));
	jdff dff_A_9oAWMnwV5_0(.dout(w_dff_A_itbOQPyI8_0),.din(w_dff_A_9oAWMnwV5_0),.clk(gclk));
	jdff dff_A_itbOQPyI8_0(.dout(w_dff_A_5sJ6YlhE0_0),.din(w_dff_A_itbOQPyI8_0),.clk(gclk));
	jdff dff_A_5sJ6YlhE0_0(.dout(w_dff_A_zQTQgKmI8_0),.din(w_dff_A_5sJ6YlhE0_0),.clk(gclk));
	jdff dff_A_zQTQgKmI8_0(.dout(w_dff_A_YvDT5LJy2_0),.din(w_dff_A_zQTQgKmI8_0),.clk(gclk));
	jdff dff_A_YvDT5LJy2_0(.dout(w_dff_A_m5WIJLH01_0),.din(w_dff_A_YvDT5LJy2_0),.clk(gclk));
	jdff dff_A_m5WIJLH01_0(.dout(w_dff_A_w9bbeijX5_0),.din(w_dff_A_m5WIJLH01_0),.clk(gclk));
	jdff dff_A_w9bbeijX5_0(.dout(w_dff_A_RCp7v3LI6_0),.din(w_dff_A_w9bbeijX5_0),.clk(gclk));
	jdff dff_A_RCp7v3LI6_0(.dout(w_dff_A_hZ2y1I6z7_0),.din(w_dff_A_RCp7v3LI6_0),.clk(gclk));
	jdff dff_A_hZ2y1I6z7_0(.dout(w_dff_A_O4NcS5zP9_0),.din(w_dff_A_hZ2y1I6z7_0),.clk(gclk));
	jdff dff_A_O4NcS5zP9_0(.dout(w_dff_A_Ui8WGGKu5_0),.din(w_dff_A_O4NcS5zP9_0),.clk(gclk));
	jdff dff_A_Ui8WGGKu5_0(.dout(w_dff_A_1mrLadKT3_0),.din(w_dff_A_Ui8WGGKu5_0),.clk(gclk));
	jdff dff_A_1mrLadKT3_0(.dout(w_dff_A_1me7KQPp4_0),.din(w_dff_A_1mrLadKT3_0),.clk(gclk));
	jdff dff_A_1me7KQPp4_0(.dout(w_dff_A_BusWKVox3_0),.din(w_dff_A_1me7KQPp4_0),.clk(gclk));
	jdff dff_A_BusWKVox3_0(.dout(w_dff_A_qWhdg15Q7_0),.din(w_dff_A_BusWKVox3_0),.clk(gclk));
	jdff dff_A_qWhdg15Q7_0(.dout(w_dff_A_ZUpbi2yz0_0),.din(w_dff_A_qWhdg15Q7_0),.clk(gclk));
	jdff dff_A_ZUpbi2yz0_0(.dout(w_dff_A_pcGYwQm57_0),.din(w_dff_A_ZUpbi2yz0_0),.clk(gclk));
	jdff dff_A_pcGYwQm57_0(.dout(w_dff_A_c8K4Cbv56_0),.din(w_dff_A_pcGYwQm57_0),.clk(gclk));
	jdff dff_A_c8K4Cbv56_0(.dout(w_dff_A_9GYIiBBj0_0),.din(w_dff_A_c8K4Cbv56_0),.clk(gclk));
	jdff dff_A_9GYIiBBj0_0(.dout(w_dff_A_K0BXssRL8_0),.din(w_dff_A_9GYIiBBj0_0),.clk(gclk));
	jdff dff_A_K0BXssRL8_0(.dout(w_dff_A_lQ0zgZkC0_0),.din(w_dff_A_K0BXssRL8_0),.clk(gclk));
	jdff dff_A_lQ0zgZkC0_0(.dout(G484),.din(w_dff_A_lQ0zgZkC0_0),.clk(gclk));
	jdff dff_A_EMBTB4wN2_1(.dout(w_dff_A_IoHE6y2G1_0),.din(w_dff_A_EMBTB4wN2_1),.clk(gclk));
	jdff dff_A_IoHE6y2G1_0(.dout(w_dff_A_CRCKyV2J4_0),.din(w_dff_A_IoHE6y2G1_0),.clk(gclk));
	jdff dff_A_CRCKyV2J4_0(.dout(w_dff_A_It3jCPbb7_0),.din(w_dff_A_CRCKyV2J4_0),.clk(gclk));
	jdff dff_A_It3jCPbb7_0(.dout(w_dff_A_EvQ6WAxz3_0),.din(w_dff_A_It3jCPbb7_0),.clk(gclk));
	jdff dff_A_EvQ6WAxz3_0(.dout(w_dff_A_tyTOJb811_0),.din(w_dff_A_EvQ6WAxz3_0),.clk(gclk));
	jdff dff_A_tyTOJb811_0(.dout(w_dff_A_9jO1Pc4Z1_0),.din(w_dff_A_tyTOJb811_0),.clk(gclk));
	jdff dff_A_9jO1Pc4Z1_0(.dout(w_dff_A_i0eG4moB5_0),.din(w_dff_A_9jO1Pc4Z1_0),.clk(gclk));
	jdff dff_A_i0eG4moB5_0(.dout(w_dff_A_PSmzHllw7_0),.din(w_dff_A_i0eG4moB5_0),.clk(gclk));
	jdff dff_A_PSmzHllw7_0(.dout(w_dff_A_Rj64f1GF7_0),.din(w_dff_A_PSmzHllw7_0),.clk(gclk));
	jdff dff_A_Rj64f1GF7_0(.dout(w_dff_A_duSYX4qP7_0),.din(w_dff_A_Rj64f1GF7_0),.clk(gclk));
	jdff dff_A_duSYX4qP7_0(.dout(w_dff_A_Y0bI5ljX6_0),.din(w_dff_A_duSYX4qP7_0),.clk(gclk));
	jdff dff_A_Y0bI5ljX6_0(.dout(w_dff_A_Sk5yPAOL4_0),.din(w_dff_A_Y0bI5ljX6_0),.clk(gclk));
	jdff dff_A_Sk5yPAOL4_0(.dout(w_dff_A_JOo7Meza7_0),.din(w_dff_A_Sk5yPAOL4_0),.clk(gclk));
	jdff dff_A_JOo7Meza7_0(.dout(w_dff_A_5MgsQhsR3_0),.din(w_dff_A_JOo7Meza7_0),.clk(gclk));
	jdff dff_A_5MgsQhsR3_0(.dout(w_dff_A_32jWazju9_0),.din(w_dff_A_5MgsQhsR3_0),.clk(gclk));
	jdff dff_A_32jWazju9_0(.dout(w_dff_A_OM6qYM0T6_0),.din(w_dff_A_32jWazju9_0),.clk(gclk));
	jdff dff_A_OM6qYM0T6_0(.dout(w_dff_A_vhii8myx2_0),.din(w_dff_A_OM6qYM0T6_0),.clk(gclk));
	jdff dff_A_vhii8myx2_0(.dout(w_dff_A_kpomkAPO6_0),.din(w_dff_A_vhii8myx2_0),.clk(gclk));
	jdff dff_A_kpomkAPO6_0(.dout(w_dff_A_qjRaUpfn9_0),.din(w_dff_A_kpomkAPO6_0),.clk(gclk));
	jdff dff_A_qjRaUpfn9_0(.dout(w_dff_A_gSvF2GPJ4_0),.din(w_dff_A_qjRaUpfn9_0),.clk(gclk));
	jdff dff_A_gSvF2GPJ4_0(.dout(w_dff_A_rccswgV80_0),.din(w_dff_A_gSvF2GPJ4_0),.clk(gclk));
	jdff dff_A_rccswgV80_0(.dout(w_dff_A_qcqOanec3_0),.din(w_dff_A_rccswgV80_0),.clk(gclk));
	jdff dff_A_qcqOanec3_0(.dout(w_dff_A_tXEIIjLp2_0),.din(w_dff_A_qcqOanec3_0),.clk(gclk));
	jdff dff_A_tXEIIjLp2_0(.dout(w_dff_A_AtDqQuHg8_0),.din(w_dff_A_tXEIIjLp2_0),.clk(gclk));
	jdff dff_A_AtDqQuHg8_0(.dout(w_dff_A_Q2j1m7Ss5_0),.din(w_dff_A_AtDqQuHg8_0),.clk(gclk));
	jdff dff_A_Q2j1m7Ss5_0(.dout(w_dff_A_aaGHbAOQ6_0),.din(w_dff_A_Q2j1m7Ss5_0),.clk(gclk));
	jdff dff_A_aaGHbAOQ6_0(.dout(w_dff_A_Cz7yroOU7_0),.din(w_dff_A_aaGHbAOQ6_0),.clk(gclk));
	jdff dff_A_Cz7yroOU7_0(.dout(w_dff_A_HLh0ajyc6_0),.din(w_dff_A_Cz7yroOU7_0),.clk(gclk));
	jdff dff_A_HLh0ajyc6_0(.dout(w_dff_A_tJ1lhrs51_0),.din(w_dff_A_HLh0ajyc6_0),.clk(gclk));
	jdff dff_A_tJ1lhrs51_0(.dout(w_dff_A_nv8A5vB52_0),.din(w_dff_A_tJ1lhrs51_0),.clk(gclk));
	jdff dff_A_nv8A5vB52_0(.dout(w_dff_A_lK8WX9Ux3_0),.din(w_dff_A_nv8A5vB52_0),.clk(gclk));
	jdff dff_A_lK8WX9Ux3_0(.dout(w_dff_A_Yc2GXOPw8_0),.din(w_dff_A_lK8WX9Ux3_0),.clk(gclk));
	jdff dff_A_Yc2GXOPw8_0(.dout(w_dff_A_lF1pILYu0_0),.din(w_dff_A_Yc2GXOPw8_0),.clk(gclk));
	jdff dff_A_lF1pILYu0_0(.dout(w_dff_A_BwcXCgqW6_0),.din(w_dff_A_lF1pILYu0_0),.clk(gclk));
	jdff dff_A_BwcXCgqW6_0(.dout(w_dff_A_1qNGERZW3_0),.din(w_dff_A_BwcXCgqW6_0),.clk(gclk));
	jdff dff_A_1qNGERZW3_0(.dout(w_dff_A_evvhmfus2_0),.din(w_dff_A_1qNGERZW3_0),.clk(gclk));
	jdff dff_A_evvhmfus2_0(.dout(w_dff_A_tE92VkYX4_0),.din(w_dff_A_evvhmfus2_0),.clk(gclk));
	jdff dff_A_tE92VkYX4_0(.dout(w_dff_A_1PhMdYyO0_0),.din(w_dff_A_tE92VkYX4_0),.clk(gclk));
	jdff dff_A_1PhMdYyO0_0(.dout(G482),.din(w_dff_A_1PhMdYyO0_0),.clk(gclk));
	jdff dff_A_VAefslF47_1(.dout(w_dff_A_JBKSPWoC8_0),.din(w_dff_A_VAefslF47_1),.clk(gclk));
	jdff dff_A_JBKSPWoC8_0(.dout(w_dff_A_OPPhVcSZ0_0),.din(w_dff_A_JBKSPWoC8_0),.clk(gclk));
	jdff dff_A_OPPhVcSZ0_0(.dout(w_dff_A_a6NZlSbf6_0),.din(w_dff_A_OPPhVcSZ0_0),.clk(gclk));
	jdff dff_A_a6NZlSbf6_0(.dout(w_dff_A_BXlAGvn60_0),.din(w_dff_A_a6NZlSbf6_0),.clk(gclk));
	jdff dff_A_BXlAGvn60_0(.dout(w_dff_A_X1n7Qtwh0_0),.din(w_dff_A_BXlAGvn60_0),.clk(gclk));
	jdff dff_A_X1n7Qtwh0_0(.dout(w_dff_A_yucbsa8e4_0),.din(w_dff_A_X1n7Qtwh0_0),.clk(gclk));
	jdff dff_A_yucbsa8e4_0(.dout(w_dff_A_a2QxJeVJ6_0),.din(w_dff_A_yucbsa8e4_0),.clk(gclk));
	jdff dff_A_a2QxJeVJ6_0(.dout(w_dff_A_f85D9rMQ2_0),.din(w_dff_A_a2QxJeVJ6_0),.clk(gclk));
	jdff dff_A_f85D9rMQ2_0(.dout(w_dff_A_64FeIGDE9_0),.din(w_dff_A_f85D9rMQ2_0),.clk(gclk));
	jdff dff_A_64FeIGDE9_0(.dout(w_dff_A_MTcnVtGT9_0),.din(w_dff_A_64FeIGDE9_0),.clk(gclk));
	jdff dff_A_MTcnVtGT9_0(.dout(w_dff_A_8VMW9GZG7_0),.din(w_dff_A_MTcnVtGT9_0),.clk(gclk));
	jdff dff_A_8VMW9GZG7_0(.dout(w_dff_A_6aRbW8xq3_0),.din(w_dff_A_8VMW9GZG7_0),.clk(gclk));
	jdff dff_A_6aRbW8xq3_0(.dout(w_dff_A_ERLEFsQR9_0),.din(w_dff_A_6aRbW8xq3_0),.clk(gclk));
	jdff dff_A_ERLEFsQR9_0(.dout(w_dff_A_FESRtSQO2_0),.din(w_dff_A_ERLEFsQR9_0),.clk(gclk));
	jdff dff_A_FESRtSQO2_0(.dout(w_dff_A_WWBzT8wE6_0),.din(w_dff_A_FESRtSQO2_0),.clk(gclk));
	jdff dff_A_WWBzT8wE6_0(.dout(w_dff_A_Xvy2JFTU7_0),.din(w_dff_A_WWBzT8wE6_0),.clk(gclk));
	jdff dff_A_Xvy2JFTU7_0(.dout(w_dff_A_o13GDJGJ3_0),.din(w_dff_A_Xvy2JFTU7_0),.clk(gclk));
	jdff dff_A_o13GDJGJ3_0(.dout(w_dff_A_bQmPcBNf4_0),.din(w_dff_A_o13GDJGJ3_0),.clk(gclk));
	jdff dff_A_bQmPcBNf4_0(.dout(w_dff_A_S86RJ6dr8_0),.din(w_dff_A_bQmPcBNf4_0),.clk(gclk));
	jdff dff_A_S86RJ6dr8_0(.dout(w_dff_A_5FIWgv9i7_0),.din(w_dff_A_S86RJ6dr8_0),.clk(gclk));
	jdff dff_A_5FIWgv9i7_0(.dout(w_dff_A_9qExALMw3_0),.din(w_dff_A_5FIWgv9i7_0),.clk(gclk));
	jdff dff_A_9qExALMw3_0(.dout(w_dff_A_cVaoeYiy3_0),.din(w_dff_A_9qExALMw3_0),.clk(gclk));
	jdff dff_A_cVaoeYiy3_0(.dout(w_dff_A_aDuNBe4C2_0),.din(w_dff_A_cVaoeYiy3_0),.clk(gclk));
	jdff dff_A_aDuNBe4C2_0(.dout(w_dff_A_9ezcKQ2K6_0),.din(w_dff_A_aDuNBe4C2_0),.clk(gclk));
	jdff dff_A_9ezcKQ2K6_0(.dout(w_dff_A_sLJL2ump7_0),.din(w_dff_A_9ezcKQ2K6_0),.clk(gclk));
	jdff dff_A_sLJL2ump7_0(.dout(w_dff_A_GTgNNpKc9_0),.din(w_dff_A_sLJL2ump7_0),.clk(gclk));
	jdff dff_A_GTgNNpKc9_0(.dout(w_dff_A_4qD0BJyu8_0),.din(w_dff_A_GTgNNpKc9_0),.clk(gclk));
	jdff dff_A_4qD0BJyu8_0(.dout(w_dff_A_aDrnXGyr2_0),.din(w_dff_A_4qD0BJyu8_0),.clk(gclk));
	jdff dff_A_aDrnXGyr2_0(.dout(w_dff_A_fnaRMI3b3_0),.din(w_dff_A_aDrnXGyr2_0),.clk(gclk));
	jdff dff_A_fnaRMI3b3_0(.dout(w_dff_A_ZWBFPxkZ0_0),.din(w_dff_A_fnaRMI3b3_0),.clk(gclk));
	jdff dff_A_ZWBFPxkZ0_0(.dout(w_dff_A_5IOP0DJc7_0),.din(w_dff_A_ZWBFPxkZ0_0),.clk(gclk));
	jdff dff_A_5IOP0DJc7_0(.dout(w_dff_A_OCtiaLFi3_0),.din(w_dff_A_5IOP0DJc7_0),.clk(gclk));
	jdff dff_A_OCtiaLFi3_0(.dout(w_dff_A_cUHbVPUs4_0),.din(w_dff_A_OCtiaLFi3_0),.clk(gclk));
	jdff dff_A_cUHbVPUs4_0(.dout(w_dff_A_asxETMYj4_0),.din(w_dff_A_cUHbVPUs4_0),.clk(gclk));
	jdff dff_A_asxETMYj4_0(.dout(w_dff_A_4FAYoMdA1_0),.din(w_dff_A_asxETMYj4_0),.clk(gclk));
	jdff dff_A_4FAYoMdA1_0(.dout(w_dff_A_dPzmdegS9_0),.din(w_dff_A_4FAYoMdA1_0),.clk(gclk));
	jdff dff_A_dPzmdegS9_0(.dout(w_dff_A_XC1xLJcF0_0),.din(w_dff_A_dPzmdegS9_0),.clk(gclk));
	jdff dff_A_XC1xLJcF0_0(.dout(w_dff_A_STVrNXob7_0),.din(w_dff_A_XC1xLJcF0_0),.clk(gclk));
	jdff dff_A_STVrNXob7_0(.dout(G480),.din(w_dff_A_STVrNXob7_0),.clk(gclk));
	jdff dff_A_upXkuxo17_1(.dout(w_dff_A_Wn9Unnih0_0),.din(w_dff_A_upXkuxo17_1),.clk(gclk));
	jdff dff_A_Wn9Unnih0_0(.dout(w_dff_A_aJvUgXFv1_0),.din(w_dff_A_Wn9Unnih0_0),.clk(gclk));
	jdff dff_A_aJvUgXFv1_0(.dout(w_dff_A_zNFZLKtX5_0),.din(w_dff_A_aJvUgXFv1_0),.clk(gclk));
	jdff dff_A_zNFZLKtX5_0(.dout(w_dff_A_rNj0B5FC6_0),.din(w_dff_A_zNFZLKtX5_0),.clk(gclk));
	jdff dff_A_rNj0B5FC6_0(.dout(w_dff_A_lb38hRM56_0),.din(w_dff_A_rNj0B5FC6_0),.clk(gclk));
	jdff dff_A_lb38hRM56_0(.dout(w_dff_A_dDTOJb5V5_0),.din(w_dff_A_lb38hRM56_0),.clk(gclk));
	jdff dff_A_dDTOJb5V5_0(.dout(w_dff_A_LBsMNjSL7_0),.din(w_dff_A_dDTOJb5V5_0),.clk(gclk));
	jdff dff_A_LBsMNjSL7_0(.dout(w_dff_A_NvktGuoa2_0),.din(w_dff_A_LBsMNjSL7_0),.clk(gclk));
	jdff dff_A_NvktGuoa2_0(.dout(w_dff_A_APzxr2dN8_0),.din(w_dff_A_NvktGuoa2_0),.clk(gclk));
	jdff dff_A_APzxr2dN8_0(.dout(w_dff_A_SbKVvb031_0),.din(w_dff_A_APzxr2dN8_0),.clk(gclk));
	jdff dff_A_SbKVvb031_0(.dout(w_dff_A_XRg64ZFO1_0),.din(w_dff_A_SbKVvb031_0),.clk(gclk));
	jdff dff_A_XRg64ZFO1_0(.dout(w_dff_A_1kMLIqZZ1_0),.din(w_dff_A_XRg64ZFO1_0),.clk(gclk));
	jdff dff_A_1kMLIqZZ1_0(.dout(w_dff_A_5T4sD9UH3_0),.din(w_dff_A_1kMLIqZZ1_0),.clk(gclk));
	jdff dff_A_5T4sD9UH3_0(.dout(w_dff_A_z66Swu4g2_0),.din(w_dff_A_5T4sD9UH3_0),.clk(gclk));
	jdff dff_A_z66Swu4g2_0(.dout(w_dff_A_hv17DihY8_0),.din(w_dff_A_z66Swu4g2_0),.clk(gclk));
	jdff dff_A_hv17DihY8_0(.dout(w_dff_A_S7WeAWGe3_0),.din(w_dff_A_hv17DihY8_0),.clk(gclk));
	jdff dff_A_S7WeAWGe3_0(.dout(w_dff_A_d5lJUpOD1_0),.din(w_dff_A_S7WeAWGe3_0),.clk(gclk));
	jdff dff_A_d5lJUpOD1_0(.dout(w_dff_A_WWdVHldh0_0),.din(w_dff_A_d5lJUpOD1_0),.clk(gclk));
	jdff dff_A_WWdVHldh0_0(.dout(w_dff_A_ZqE2E6vf6_0),.din(w_dff_A_WWdVHldh0_0),.clk(gclk));
	jdff dff_A_ZqE2E6vf6_0(.dout(w_dff_A_pss353h47_0),.din(w_dff_A_ZqE2E6vf6_0),.clk(gclk));
	jdff dff_A_pss353h47_0(.dout(w_dff_A_KU1ZnUpb4_0),.din(w_dff_A_pss353h47_0),.clk(gclk));
	jdff dff_A_KU1ZnUpb4_0(.dout(w_dff_A_OfuAARV19_0),.din(w_dff_A_KU1ZnUpb4_0),.clk(gclk));
	jdff dff_A_OfuAARV19_0(.dout(w_dff_A_ABqyipJf1_0),.din(w_dff_A_OfuAARV19_0),.clk(gclk));
	jdff dff_A_ABqyipJf1_0(.dout(w_dff_A_ZKbfW3Cy0_0),.din(w_dff_A_ABqyipJf1_0),.clk(gclk));
	jdff dff_A_ZKbfW3Cy0_0(.dout(w_dff_A_IbNmOxoV4_0),.din(w_dff_A_ZKbfW3Cy0_0),.clk(gclk));
	jdff dff_A_IbNmOxoV4_0(.dout(w_dff_A_FZcQF5jg5_0),.din(w_dff_A_IbNmOxoV4_0),.clk(gclk));
	jdff dff_A_FZcQF5jg5_0(.dout(w_dff_A_8BLrQC5q1_0),.din(w_dff_A_FZcQF5jg5_0),.clk(gclk));
	jdff dff_A_8BLrQC5q1_0(.dout(w_dff_A_wdIYs3126_0),.din(w_dff_A_8BLrQC5q1_0),.clk(gclk));
	jdff dff_A_wdIYs3126_0(.dout(w_dff_A_rVxrWfsv1_0),.din(w_dff_A_wdIYs3126_0),.clk(gclk));
	jdff dff_A_rVxrWfsv1_0(.dout(w_dff_A_cyJkNSPU9_0),.din(w_dff_A_rVxrWfsv1_0),.clk(gclk));
	jdff dff_A_cyJkNSPU9_0(.dout(w_dff_A_iwU0qOZu8_0),.din(w_dff_A_cyJkNSPU9_0),.clk(gclk));
	jdff dff_A_iwU0qOZu8_0(.dout(w_dff_A_D1RKJ3lC8_0),.din(w_dff_A_iwU0qOZu8_0),.clk(gclk));
	jdff dff_A_D1RKJ3lC8_0(.dout(w_dff_A_NWpkGv7f6_0),.din(w_dff_A_D1RKJ3lC8_0),.clk(gclk));
	jdff dff_A_NWpkGv7f6_0(.dout(w_dff_A_ixeIN3Wb2_0),.din(w_dff_A_NWpkGv7f6_0),.clk(gclk));
	jdff dff_A_ixeIN3Wb2_0(.dout(w_dff_A_uumBwDeW0_0),.din(w_dff_A_ixeIN3Wb2_0),.clk(gclk));
	jdff dff_A_uumBwDeW0_0(.dout(w_dff_A_mWPf6GnF4_0),.din(w_dff_A_uumBwDeW0_0),.clk(gclk));
	jdff dff_A_mWPf6GnF4_0(.dout(w_dff_A_5Q5DPuZB4_0),.din(w_dff_A_mWPf6GnF4_0),.clk(gclk));
	jdff dff_A_5Q5DPuZB4_0(.dout(w_dff_A_9HkFBm2c0_0),.din(w_dff_A_5Q5DPuZB4_0),.clk(gclk));
	jdff dff_A_9HkFBm2c0_0(.dout(G560),.din(w_dff_A_9HkFBm2c0_0),.clk(gclk));
	jdff dff_A_lj9ELOAr8_1(.dout(w_dff_A_6zCZWMoL3_0),.din(w_dff_A_lj9ELOAr8_1),.clk(gclk));
	jdff dff_A_6zCZWMoL3_0(.dout(w_dff_A_YSPSA9jN6_0),.din(w_dff_A_6zCZWMoL3_0),.clk(gclk));
	jdff dff_A_YSPSA9jN6_0(.dout(w_dff_A_yNx3sJVN3_0),.din(w_dff_A_YSPSA9jN6_0),.clk(gclk));
	jdff dff_A_yNx3sJVN3_0(.dout(w_dff_A_JeyC7pDw4_0),.din(w_dff_A_yNx3sJVN3_0),.clk(gclk));
	jdff dff_A_JeyC7pDw4_0(.dout(w_dff_A_fZblbgIO6_0),.din(w_dff_A_JeyC7pDw4_0),.clk(gclk));
	jdff dff_A_fZblbgIO6_0(.dout(w_dff_A_6jMTSsvL1_0),.din(w_dff_A_fZblbgIO6_0),.clk(gclk));
	jdff dff_A_6jMTSsvL1_0(.dout(w_dff_A_MqPguq3f9_0),.din(w_dff_A_6jMTSsvL1_0),.clk(gclk));
	jdff dff_A_MqPguq3f9_0(.dout(w_dff_A_kg5IneT15_0),.din(w_dff_A_MqPguq3f9_0),.clk(gclk));
	jdff dff_A_kg5IneT15_0(.dout(w_dff_A_olezRIXR0_0),.din(w_dff_A_kg5IneT15_0),.clk(gclk));
	jdff dff_A_olezRIXR0_0(.dout(w_dff_A_v8GcbxwV1_0),.din(w_dff_A_olezRIXR0_0),.clk(gclk));
	jdff dff_A_v8GcbxwV1_0(.dout(w_dff_A_PTbN5GtS4_0),.din(w_dff_A_v8GcbxwV1_0),.clk(gclk));
	jdff dff_A_PTbN5GtS4_0(.dout(w_dff_A_wSNhGyHy5_0),.din(w_dff_A_PTbN5GtS4_0),.clk(gclk));
	jdff dff_A_wSNhGyHy5_0(.dout(w_dff_A_ZjRMimW17_0),.din(w_dff_A_wSNhGyHy5_0),.clk(gclk));
	jdff dff_A_ZjRMimW17_0(.dout(w_dff_A_5Tolaqjh3_0),.din(w_dff_A_ZjRMimW17_0),.clk(gclk));
	jdff dff_A_5Tolaqjh3_0(.dout(w_dff_A_YAhmTbcy2_0),.din(w_dff_A_5Tolaqjh3_0),.clk(gclk));
	jdff dff_A_YAhmTbcy2_0(.dout(w_dff_A_Z6mvE0qT1_0),.din(w_dff_A_YAhmTbcy2_0),.clk(gclk));
	jdff dff_A_Z6mvE0qT1_0(.dout(w_dff_A_MEeOtyWo3_0),.din(w_dff_A_Z6mvE0qT1_0),.clk(gclk));
	jdff dff_A_MEeOtyWo3_0(.dout(w_dff_A_pvT1zztD0_0),.din(w_dff_A_MEeOtyWo3_0),.clk(gclk));
	jdff dff_A_pvT1zztD0_0(.dout(w_dff_A_bGlGukqE6_0),.din(w_dff_A_pvT1zztD0_0),.clk(gclk));
	jdff dff_A_bGlGukqE6_0(.dout(w_dff_A_7BsqMZ3u1_0),.din(w_dff_A_bGlGukqE6_0),.clk(gclk));
	jdff dff_A_7BsqMZ3u1_0(.dout(w_dff_A_v2LvFqxO8_0),.din(w_dff_A_7BsqMZ3u1_0),.clk(gclk));
	jdff dff_A_v2LvFqxO8_0(.dout(w_dff_A_tpJHmUX28_0),.din(w_dff_A_v2LvFqxO8_0),.clk(gclk));
	jdff dff_A_tpJHmUX28_0(.dout(w_dff_A_S3wmCYtg5_0),.din(w_dff_A_tpJHmUX28_0),.clk(gclk));
	jdff dff_A_S3wmCYtg5_0(.dout(w_dff_A_tE0tCvh50_0),.din(w_dff_A_S3wmCYtg5_0),.clk(gclk));
	jdff dff_A_tE0tCvh50_0(.dout(w_dff_A_cHob9g9y3_0),.din(w_dff_A_tE0tCvh50_0),.clk(gclk));
	jdff dff_A_cHob9g9y3_0(.dout(w_dff_A_KLvQQeKS0_0),.din(w_dff_A_cHob9g9y3_0),.clk(gclk));
	jdff dff_A_KLvQQeKS0_0(.dout(w_dff_A_kTq0Bqeq0_0),.din(w_dff_A_KLvQQeKS0_0),.clk(gclk));
	jdff dff_A_kTq0Bqeq0_0(.dout(w_dff_A_rgFVGm4K0_0),.din(w_dff_A_kTq0Bqeq0_0),.clk(gclk));
	jdff dff_A_rgFVGm4K0_0(.dout(w_dff_A_BqhQa66W8_0),.din(w_dff_A_rgFVGm4K0_0),.clk(gclk));
	jdff dff_A_BqhQa66W8_0(.dout(w_dff_A_dedRN3x89_0),.din(w_dff_A_BqhQa66W8_0),.clk(gclk));
	jdff dff_A_dedRN3x89_0(.dout(w_dff_A_G95fJe0B4_0),.din(w_dff_A_dedRN3x89_0),.clk(gclk));
	jdff dff_A_G95fJe0B4_0(.dout(w_dff_A_5quZoQEu3_0),.din(w_dff_A_G95fJe0B4_0),.clk(gclk));
	jdff dff_A_5quZoQEu3_0(.dout(w_dff_A_RjUlvdqL7_0),.din(w_dff_A_5quZoQEu3_0),.clk(gclk));
	jdff dff_A_RjUlvdqL7_0(.dout(w_dff_A_M4eR8Hkc6_0),.din(w_dff_A_RjUlvdqL7_0),.clk(gclk));
	jdff dff_A_M4eR8Hkc6_0(.dout(w_dff_A_9srIdFhF1_0),.din(w_dff_A_M4eR8Hkc6_0),.clk(gclk));
	jdff dff_A_9srIdFhF1_0(.dout(w_dff_A_hTjntdic8_0),.din(w_dff_A_9srIdFhF1_0),.clk(gclk));
	jdff dff_A_hTjntdic8_0(.dout(w_dff_A_AoQ929dH0_0),.din(w_dff_A_hTjntdic8_0),.clk(gclk));
	jdff dff_A_AoQ929dH0_0(.dout(w_dff_A_PPqc7LGB7_0),.din(w_dff_A_AoQ929dH0_0),.clk(gclk));
	jdff dff_A_PPqc7LGB7_0(.dout(G542),.din(w_dff_A_PPqc7LGB7_0),.clk(gclk));
	jdff dff_A_sDPgk8v97_1(.dout(w_dff_A_cFtTmN0o2_0),.din(w_dff_A_sDPgk8v97_1),.clk(gclk));
	jdff dff_A_cFtTmN0o2_0(.dout(w_dff_A_kiiRQhBW5_0),.din(w_dff_A_cFtTmN0o2_0),.clk(gclk));
	jdff dff_A_kiiRQhBW5_0(.dout(w_dff_A_aCe00na87_0),.din(w_dff_A_kiiRQhBW5_0),.clk(gclk));
	jdff dff_A_aCe00na87_0(.dout(w_dff_A_o7q1aemK9_0),.din(w_dff_A_aCe00na87_0),.clk(gclk));
	jdff dff_A_o7q1aemK9_0(.dout(w_dff_A_LkEF3ArN2_0),.din(w_dff_A_o7q1aemK9_0),.clk(gclk));
	jdff dff_A_LkEF3ArN2_0(.dout(w_dff_A_qIhctuWI9_0),.din(w_dff_A_LkEF3ArN2_0),.clk(gclk));
	jdff dff_A_qIhctuWI9_0(.dout(w_dff_A_9UhuZQLk7_0),.din(w_dff_A_qIhctuWI9_0),.clk(gclk));
	jdff dff_A_9UhuZQLk7_0(.dout(w_dff_A_jh42ni1M2_0),.din(w_dff_A_9UhuZQLk7_0),.clk(gclk));
	jdff dff_A_jh42ni1M2_0(.dout(w_dff_A_ZdjbCOHO3_0),.din(w_dff_A_jh42ni1M2_0),.clk(gclk));
	jdff dff_A_ZdjbCOHO3_0(.dout(w_dff_A_nI3iIqcp4_0),.din(w_dff_A_ZdjbCOHO3_0),.clk(gclk));
	jdff dff_A_nI3iIqcp4_0(.dout(w_dff_A_mO0rfzEW8_0),.din(w_dff_A_nI3iIqcp4_0),.clk(gclk));
	jdff dff_A_mO0rfzEW8_0(.dout(w_dff_A_R41Q2i7T6_0),.din(w_dff_A_mO0rfzEW8_0),.clk(gclk));
	jdff dff_A_R41Q2i7T6_0(.dout(w_dff_A_wNCqBHlr2_0),.din(w_dff_A_R41Q2i7T6_0),.clk(gclk));
	jdff dff_A_wNCqBHlr2_0(.dout(w_dff_A_4tyyoAOk5_0),.din(w_dff_A_wNCqBHlr2_0),.clk(gclk));
	jdff dff_A_4tyyoAOk5_0(.dout(w_dff_A_KjDSevLa3_0),.din(w_dff_A_4tyyoAOk5_0),.clk(gclk));
	jdff dff_A_KjDSevLa3_0(.dout(w_dff_A_A8oEypnS0_0),.din(w_dff_A_KjDSevLa3_0),.clk(gclk));
	jdff dff_A_A8oEypnS0_0(.dout(w_dff_A_jCSJLyrE3_0),.din(w_dff_A_A8oEypnS0_0),.clk(gclk));
	jdff dff_A_jCSJLyrE3_0(.dout(w_dff_A_XtPCZB0c9_0),.din(w_dff_A_jCSJLyrE3_0),.clk(gclk));
	jdff dff_A_XtPCZB0c9_0(.dout(w_dff_A_uivzbkmY3_0),.din(w_dff_A_XtPCZB0c9_0),.clk(gclk));
	jdff dff_A_uivzbkmY3_0(.dout(w_dff_A_UnZckhH29_0),.din(w_dff_A_uivzbkmY3_0),.clk(gclk));
	jdff dff_A_UnZckhH29_0(.dout(w_dff_A_cfdmVm6c6_0),.din(w_dff_A_UnZckhH29_0),.clk(gclk));
	jdff dff_A_cfdmVm6c6_0(.dout(w_dff_A_g3R2Ld1J1_0),.din(w_dff_A_cfdmVm6c6_0),.clk(gclk));
	jdff dff_A_g3R2Ld1J1_0(.dout(w_dff_A_sLMpOUEi6_0),.din(w_dff_A_g3R2Ld1J1_0),.clk(gclk));
	jdff dff_A_sLMpOUEi6_0(.dout(w_dff_A_x4it03PW9_0),.din(w_dff_A_sLMpOUEi6_0),.clk(gclk));
	jdff dff_A_x4it03PW9_0(.dout(w_dff_A_6RVZL74B2_0),.din(w_dff_A_x4it03PW9_0),.clk(gclk));
	jdff dff_A_6RVZL74B2_0(.dout(w_dff_A_xzRG97JL2_0),.din(w_dff_A_6RVZL74B2_0),.clk(gclk));
	jdff dff_A_xzRG97JL2_0(.dout(w_dff_A_UnLuVhtN9_0),.din(w_dff_A_xzRG97JL2_0),.clk(gclk));
	jdff dff_A_UnLuVhtN9_0(.dout(w_dff_A_DGmXZjIi2_0),.din(w_dff_A_UnLuVhtN9_0),.clk(gclk));
	jdff dff_A_DGmXZjIi2_0(.dout(w_dff_A_CKi4v38a2_0),.din(w_dff_A_DGmXZjIi2_0),.clk(gclk));
	jdff dff_A_CKi4v38a2_0(.dout(w_dff_A_abXsWAze8_0),.din(w_dff_A_CKi4v38a2_0),.clk(gclk));
	jdff dff_A_abXsWAze8_0(.dout(w_dff_A_KoiKCyJb4_0),.din(w_dff_A_abXsWAze8_0),.clk(gclk));
	jdff dff_A_KoiKCyJb4_0(.dout(w_dff_A_MqFItUqQ6_0),.din(w_dff_A_KoiKCyJb4_0),.clk(gclk));
	jdff dff_A_MqFItUqQ6_0(.dout(w_dff_A_v0gvGUCS7_0),.din(w_dff_A_MqFItUqQ6_0),.clk(gclk));
	jdff dff_A_v0gvGUCS7_0(.dout(w_dff_A_wGcUSNGe5_0),.din(w_dff_A_v0gvGUCS7_0),.clk(gclk));
	jdff dff_A_wGcUSNGe5_0(.dout(w_dff_A_jafLSeyt9_0),.din(w_dff_A_wGcUSNGe5_0),.clk(gclk));
	jdff dff_A_jafLSeyt9_0(.dout(w_dff_A_IytHxavg9_0),.din(w_dff_A_jafLSeyt9_0),.clk(gclk));
	jdff dff_A_IytHxavg9_0(.dout(w_dff_A_dtEdkBdj1_0),.din(w_dff_A_IytHxavg9_0),.clk(gclk));
	jdff dff_A_dtEdkBdj1_0(.dout(w_dff_A_urSSzUsM1_0),.din(w_dff_A_dtEdkBdj1_0),.clk(gclk));
	jdff dff_A_urSSzUsM1_0(.dout(G558),.din(w_dff_A_urSSzUsM1_0),.clk(gclk));
	jdff dff_A_onEfvwvV6_1(.dout(w_dff_A_C0HUjNaI0_0),.din(w_dff_A_onEfvwvV6_1),.clk(gclk));
	jdff dff_A_C0HUjNaI0_0(.dout(w_dff_A_mgP1VW8e0_0),.din(w_dff_A_C0HUjNaI0_0),.clk(gclk));
	jdff dff_A_mgP1VW8e0_0(.dout(w_dff_A_SxvRvK4p9_0),.din(w_dff_A_mgP1VW8e0_0),.clk(gclk));
	jdff dff_A_SxvRvK4p9_0(.dout(w_dff_A_tx07HFfa9_0),.din(w_dff_A_SxvRvK4p9_0),.clk(gclk));
	jdff dff_A_tx07HFfa9_0(.dout(w_dff_A_JxFFZbCP5_0),.din(w_dff_A_tx07HFfa9_0),.clk(gclk));
	jdff dff_A_JxFFZbCP5_0(.dout(w_dff_A_21UPNdX36_0),.din(w_dff_A_JxFFZbCP5_0),.clk(gclk));
	jdff dff_A_21UPNdX36_0(.dout(w_dff_A_b0JFeInU2_0),.din(w_dff_A_21UPNdX36_0),.clk(gclk));
	jdff dff_A_b0JFeInU2_0(.dout(w_dff_A_lCUkQlQe8_0),.din(w_dff_A_b0JFeInU2_0),.clk(gclk));
	jdff dff_A_lCUkQlQe8_0(.dout(w_dff_A_VhomK8Ca7_0),.din(w_dff_A_lCUkQlQe8_0),.clk(gclk));
	jdff dff_A_VhomK8Ca7_0(.dout(w_dff_A_5uZiJa7h7_0),.din(w_dff_A_VhomK8Ca7_0),.clk(gclk));
	jdff dff_A_5uZiJa7h7_0(.dout(w_dff_A_8tQoMJoe3_0),.din(w_dff_A_5uZiJa7h7_0),.clk(gclk));
	jdff dff_A_8tQoMJoe3_0(.dout(w_dff_A_Nfx7iYoX8_0),.din(w_dff_A_8tQoMJoe3_0),.clk(gclk));
	jdff dff_A_Nfx7iYoX8_0(.dout(w_dff_A_Rprol9ET7_0),.din(w_dff_A_Nfx7iYoX8_0),.clk(gclk));
	jdff dff_A_Rprol9ET7_0(.dout(w_dff_A_2QPmdr2n1_0),.din(w_dff_A_Rprol9ET7_0),.clk(gclk));
	jdff dff_A_2QPmdr2n1_0(.dout(w_dff_A_O9ojFsQs8_0),.din(w_dff_A_2QPmdr2n1_0),.clk(gclk));
	jdff dff_A_O9ojFsQs8_0(.dout(w_dff_A_4C5FZ3pB9_0),.din(w_dff_A_O9ojFsQs8_0),.clk(gclk));
	jdff dff_A_4C5FZ3pB9_0(.dout(w_dff_A_nzP6p3E90_0),.din(w_dff_A_4C5FZ3pB9_0),.clk(gclk));
	jdff dff_A_nzP6p3E90_0(.dout(w_dff_A_R1PTbvuf4_0),.din(w_dff_A_nzP6p3E90_0),.clk(gclk));
	jdff dff_A_R1PTbvuf4_0(.dout(w_dff_A_ogzJ2vlA4_0),.din(w_dff_A_R1PTbvuf4_0),.clk(gclk));
	jdff dff_A_ogzJ2vlA4_0(.dout(w_dff_A_Ib00GUvM9_0),.din(w_dff_A_ogzJ2vlA4_0),.clk(gclk));
	jdff dff_A_Ib00GUvM9_0(.dout(w_dff_A_tyVrybjw2_0),.din(w_dff_A_Ib00GUvM9_0),.clk(gclk));
	jdff dff_A_tyVrybjw2_0(.dout(w_dff_A_okzfNU0q0_0),.din(w_dff_A_tyVrybjw2_0),.clk(gclk));
	jdff dff_A_okzfNU0q0_0(.dout(w_dff_A_dmrZLSd61_0),.din(w_dff_A_okzfNU0q0_0),.clk(gclk));
	jdff dff_A_dmrZLSd61_0(.dout(w_dff_A_sx9RMHmI6_0),.din(w_dff_A_dmrZLSd61_0),.clk(gclk));
	jdff dff_A_sx9RMHmI6_0(.dout(w_dff_A_xRM73C7k6_0),.din(w_dff_A_sx9RMHmI6_0),.clk(gclk));
	jdff dff_A_xRM73C7k6_0(.dout(w_dff_A_bnrbDias4_0),.din(w_dff_A_xRM73C7k6_0),.clk(gclk));
	jdff dff_A_bnrbDias4_0(.dout(w_dff_A_9Qz45vB73_0),.din(w_dff_A_bnrbDias4_0),.clk(gclk));
	jdff dff_A_9Qz45vB73_0(.dout(w_dff_A_s4JSap4n0_0),.din(w_dff_A_9Qz45vB73_0),.clk(gclk));
	jdff dff_A_s4JSap4n0_0(.dout(w_dff_A_CSwzjaeg9_0),.din(w_dff_A_s4JSap4n0_0),.clk(gclk));
	jdff dff_A_CSwzjaeg9_0(.dout(w_dff_A_MeX7d2zu9_0),.din(w_dff_A_CSwzjaeg9_0),.clk(gclk));
	jdff dff_A_MeX7d2zu9_0(.dout(w_dff_A_iVJy5de78_0),.din(w_dff_A_MeX7d2zu9_0),.clk(gclk));
	jdff dff_A_iVJy5de78_0(.dout(w_dff_A_kpk24sAm7_0),.din(w_dff_A_iVJy5de78_0),.clk(gclk));
	jdff dff_A_kpk24sAm7_0(.dout(w_dff_A_laKRt4fM5_0),.din(w_dff_A_kpk24sAm7_0),.clk(gclk));
	jdff dff_A_laKRt4fM5_0(.dout(w_dff_A_cIddYTD10_0),.din(w_dff_A_laKRt4fM5_0),.clk(gclk));
	jdff dff_A_cIddYTD10_0(.dout(w_dff_A_HPZGDjGW3_0),.din(w_dff_A_cIddYTD10_0),.clk(gclk));
	jdff dff_A_HPZGDjGW3_0(.dout(w_dff_A_NaAAazET6_0),.din(w_dff_A_HPZGDjGW3_0),.clk(gclk));
	jdff dff_A_NaAAazET6_0(.dout(w_dff_A_MjseTzEz5_0),.din(w_dff_A_NaAAazET6_0),.clk(gclk));
	jdff dff_A_MjseTzEz5_0(.dout(w_dff_A_OCoChaKG9_0),.din(w_dff_A_MjseTzEz5_0),.clk(gclk));
	jdff dff_A_OCoChaKG9_0(.dout(G556),.din(w_dff_A_OCoChaKG9_0),.clk(gclk));
	jdff dff_A_XmweTCKr8_1(.dout(w_dff_A_EOGxKO371_0),.din(w_dff_A_XmweTCKr8_1),.clk(gclk));
	jdff dff_A_EOGxKO371_0(.dout(w_dff_A_lUU18J799_0),.din(w_dff_A_EOGxKO371_0),.clk(gclk));
	jdff dff_A_lUU18J799_0(.dout(w_dff_A_afXMxmPS7_0),.din(w_dff_A_lUU18J799_0),.clk(gclk));
	jdff dff_A_afXMxmPS7_0(.dout(w_dff_A_PBRVivZf7_0),.din(w_dff_A_afXMxmPS7_0),.clk(gclk));
	jdff dff_A_PBRVivZf7_0(.dout(w_dff_A_cLRFLt8e4_0),.din(w_dff_A_PBRVivZf7_0),.clk(gclk));
	jdff dff_A_cLRFLt8e4_0(.dout(w_dff_A_4MjlSl9h2_0),.din(w_dff_A_cLRFLt8e4_0),.clk(gclk));
	jdff dff_A_4MjlSl9h2_0(.dout(w_dff_A_7D4SMPgx0_0),.din(w_dff_A_4MjlSl9h2_0),.clk(gclk));
	jdff dff_A_7D4SMPgx0_0(.dout(w_dff_A_L6EcYAQY8_0),.din(w_dff_A_7D4SMPgx0_0),.clk(gclk));
	jdff dff_A_L6EcYAQY8_0(.dout(w_dff_A_xWN4Yt747_0),.din(w_dff_A_L6EcYAQY8_0),.clk(gclk));
	jdff dff_A_xWN4Yt747_0(.dout(w_dff_A_jha5NDAS0_0),.din(w_dff_A_xWN4Yt747_0),.clk(gclk));
	jdff dff_A_jha5NDAS0_0(.dout(w_dff_A_V6VZFrcV5_0),.din(w_dff_A_jha5NDAS0_0),.clk(gclk));
	jdff dff_A_V6VZFrcV5_0(.dout(w_dff_A_GxTS27pS3_0),.din(w_dff_A_V6VZFrcV5_0),.clk(gclk));
	jdff dff_A_GxTS27pS3_0(.dout(w_dff_A_6hAUldyh3_0),.din(w_dff_A_GxTS27pS3_0),.clk(gclk));
	jdff dff_A_6hAUldyh3_0(.dout(w_dff_A_ddzQnE3b7_0),.din(w_dff_A_6hAUldyh3_0),.clk(gclk));
	jdff dff_A_ddzQnE3b7_0(.dout(w_dff_A_r17Fx0cV3_0),.din(w_dff_A_ddzQnE3b7_0),.clk(gclk));
	jdff dff_A_r17Fx0cV3_0(.dout(w_dff_A_zJstR2UV3_0),.din(w_dff_A_r17Fx0cV3_0),.clk(gclk));
	jdff dff_A_zJstR2UV3_0(.dout(w_dff_A_ZZo8oM4s1_0),.din(w_dff_A_zJstR2UV3_0),.clk(gclk));
	jdff dff_A_ZZo8oM4s1_0(.dout(w_dff_A_uiHvil4E4_0),.din(w_dff_A_ZZo8oM4s1_0),.clk(gclk));
	jdff dff_A_uiHvil4E4_0(.dout(w_dff_A_OgxjZZWi3_0),.din(w_dff_A_uiHvil4E4_0),.clk(gclk));
	jdff dff_A_OgxjZZWi3_0(.dout(w_dff_A_0DEc0Ifc7_0),.din(w_dff_A_OgxjZZWi3_0),.clk(gclk));
	jdff dff_A_0DEc0Ifc7_0(.dout(w_dff_A_Hqlz0k4G8_0),.din(w_dff_A_0DEc0Ifc7_0),.clk(gclk));
	jdff dff_A_Hqlz0k4G8_0(.dout(w_dff_A_JFUymT810_0),.din(w_dff_A_Hqlz0k4G8_0),.clk(gclk));
	jdff dff_A_JFUymT810_0(.dout(w_dff_A_j4gFUobs9_0),.din(w_dff_A_JFUymT810_0),.clk(gclk));
	jdff dff_A_j4gFUobs9_0(.dout(w_dff_A_zCm0H4ih5_0),.din(w_dff_A_j4gFUobs9_0),.clk(gclk));
	jdff dff_A_zCm0H4ih5_0(.dout(w_dff_A_l1HCIKy98_0),.din(w_dff_A_zCm0H4ih5_0),.clk(gclk));
	jdff dff_A_l1HCIKy98_0(.dout(w_dff_A_ivmLM9J73_0),.din(w_dff_A_l1HCIKy98_0),.clk(gclk));
	jdff dff_A_ivmLM9J73_0(.dout(w_dff_A_e1PfDYZZ5_0),.din(w_dff_A_ivmLM9J73_0),.clk(gclk));
	jdff dff_A_e1PfDYZZ5_0(.dout(w_dff_A_EJOAexXK6_0),.din(w_dff_A_e1PfDYZZ5_0),.clk(gclk));
	jdff dff_A_EJOAexXK6_0(.dout(w_dff_A_5tUFrWPk6_0),.din(w_dff_A_EJOAexXK6_0),.clk(gclk));
	jdff dff_A_5tUFrWPk6_0(.dout(w_dff_A_4WgN97nv7_0),.din(w_dff_A_5tUFrWPk6_0),.clk(gclk));
	jdff dff_A_4WgN97nv7_0(.dout(w_dff_A_71mgfxK79_0),.din(w_dff_A_4WgN97nv7_0),.clk(gclk));
	jdff dff_A_71mgfxK79_0(.dout(w_dff_A_2RKqtE8q8_0),.din(w_dff_A_71mgfxK79_0),.clk(gclk));
	jdff dff_A_2RKqtE8q8_0(.dout(w_dff_A_OQarV7mi0_0),.din(w_dff_A_2RKqtE8q8_0),.clk(gclk));
	jdff dff_A_OQarV7mi0_0(.dout(w_dff_A_CXHTQpki3_0),.din(w_dff_A_OQarV7mi0_0),.clk(gclk));
	jdff dff_A_CXHTQpki3_0(.dout(w_dff_A_lOjk2tqx1_0),.din(w_dff_A_CXHTQpki3_0),.clk(gclk));
	jdff dff_A_lOjk2tqx1_0(.dout(w_dff_A_UbleewQs0_0),.din(w_dff_A_lOjk2tqx1_0),.clk(gclk));
	jdff dff_A_UbleewQs0_0(.dout(w_dff_A_6RZk2ynx8_0),.din(w_dff_A_UbleewQs0_0),.clk(gclk));
	jdff dff_A_6RZk2ynx8_0(.dout(w_dff_A_r0VOjmTD7_0),.din(w_dff_A_6RZk2ynx8_0),.clk(gclk));
	jdff dff_A_r0VOjmTD7_0(.dout(G554),.din(w_dff_A_r0VOjmTD7_0),.clk(gclk));
	jdff dff_A_FwloGYnx1_1(.dout(w_dff_A_MpMoED0o2_0),.din(w_dff_A_FwloGYnx1_1),.clk(gclk));
	jdff dff_A_MpMoED0o2_0(.dout(w_dff_A_ch9L710B3_0),.din(w_dff_A_MpMoED0o2_0),.clk(gclk));
	jdff dff_A_ch9L710B3_0(.dout(w_dff_A_ZdqSW84s7_0),.din(w_dff_A_ch9L710B3_0),.clk(gclk));
	jdff dff_A_ZdqSW84s7_0(.dout(w_dff_A_tpuMJF1Z5_0),.din(w_dff_A_ZdqSW84s7_0),.clk(gclk));
	jdff dff_A_tpuMJF1Z5_0(.dout(w_dff_A_L19tyCWl8_0),.din(w_dff_A_tpuMJF1Z5_0),.clk(gclk));
	jdff dff_A_L19tyCWl8_0(.dout(w_dff_A_FfUc06ZZ5_0),.din(w_dff_A_L19tyCWl8_0),.clk(gclk));
	jdff dff_A_FfUc06ZZ5_0(.dout(w_dff_A_vJEhMdfj2_0),.din(w_dff_A_FfUc06ZZ5_0),.clk(gclk));
	jdff dff_A_vJEhMdfj2_0(.dout(w_dff_A_xUBEpP752_0),.din(w_dff_A_vJEhMdfj2_0),.clk(gclk));
	jdff dff_A_xUBEpP752_0(.dout(w_dff_A_OU8g8YTV9_0),.din(w_dff_A_xUBEpP752_0),.clk(gclk));
	jdff dff_A_OU8g8YTV9_0(.dout(w_dff_A_jI4NSncm5_0),.din(w_dff_A_OU8g8YTV9_0),.clk(gclk));
	jdff dff_A_jI4NSncm5_0(.dout(w_dff_A_ExDix2BP4_0),.din(w_dff_A_jI4NSncm5_0),.clk(gclk));
	jdff dff_A_ExDix2BP4_0(.dout(w_dff_A_d1PfQ0OE5_0),.din(w_dff_A_ExDix2BP4_0),.clk(gclk));
	jdff dff_A_d1PfQ0OE5_0(.dout(w_dff_A_kFxObhhO4_0),.din(w_dff_A_d1PfQ0OE5_0),.clk(gclk));
	jdff dff_A_kFxObhhO4_0(.dout(w_dff_A_ncMbpdAA2_0),.din(w_dff_A_kFxObhhO4_0),.clk(gclk));
	jdff dff_A_ncMbpdAA2_0(.dout(w_dff_A_xgZvbUCQ1_0),.din(w_dff_A_ncMbpdAA2_0),.clk(gclk));
	jdff dff_A_xgZvbUCQ1_0(.dout(w_dff_A_NcEbcPEE4_0),.din(w_dff_A_xgZvbUCQ1_0),.clk(gclk));
	jdff dff_A_NcEbcPEE4_0(.dout(w_dff_A_cQBgkh7U3_0),.din(w_dff_A_NcEbcPEE4_0),.clk(gclk));
	jdff dff_A_cQBgkh7U3_0(.dout(w_dff_A_FmFIRANR1_0),.din(w_dff_A_cQBgkh7U3_0),.clk(gclk));
	jdff dff_A_FmFIRANR1_0(.dout(w_dff_A_ihbKzhFi8_0),.din(w_dff_A_FmFIRANR1_0),.clk(gclk));
	jdff dff_A_ihbKzhFi8_0(.dout(w_dff_A_mwdLyVdM1_0),.din(w_dff_A_ihbKzhFi8_0),.clk(gclk));
	jdff dff_A_mwdLyVdM1_0(.dout(w_dff_A_waHtKHPG7_0),.din(w_dff_A_mwdLyVdM1_0),.clk(gclk));
	jdff dff_A_waHtKHPG7_0(.dout(w_dff_A_VK5CuF4n3_0),.din(w_dff_A_waHtKHPG7_0),.clk(gclk));
	jdff dff_A_VK5CuF4n3_0(.dout(w_dff_A_BqFHOsmc8_0),.din(w_dff_A_VK5CuF4n3_0),.clk(gclk));
	jdff dff_A_BqFHOsmc8_0(.dout(w_dff_A_rcbVpIZv6_0),.din(w_dff_A_BqFHOsmc8_0),.clk(gclk));
	jdff dff_A_rcbVpIZv6_0(.dout(w_dff_A_9I9mWfGf7_0),.din(w_dff_A_rcbVpIZv6_0),.clk(gclk));
	jdff dff_A_9I9mWfGf7_0(.dout(w_dff_A_WKRtswHN5_0),.din(w_dff_A_9I9mWfGf7_0),.clk(gclk));
	jdff dff_A_WKRtswHN5_0(.dout(w_dff_A_JSQxALEH2_0),.din(w_dff_A_WKRtswHN5_0),.clk(gclk));
	jdff dff_A_JSQxALEH2_0(.dout(w_dff_A_gpUwEeBL5_0),.din(w_dff_A_JSQxALEH2_0),.clk(gclk));
	jdff dff_A_gpUwEeBL5_0(.dout(w_dff_A_ukvlCemw2_0),.din(w_dff_A_gpUwEeBL5_0),.clk(gclk));
	jdff dff_A_ukvlCemw2_0(.dout(w_dff_A_KzXZROGU7_0),.din(w_dff_A_ukvlCemw2_0),.clk(gclk));
	jdff dff_A_KzXZROGU7_0(.dout(w_dff_A_TA578Zcc5_0),.din(w_dff_A_KzXZROGU7_0),.clk(gclk));
	jdff dff_A_TA578Zcc5_0(.dout(w_dff_A_4vJ2qQSY1_0),.din(w_dff_A_TA578Zcc5_0),.clk(gclk));
	jdff dff_A_4vJ2qQSY1_0(.dout(w_dff_A_IvvnpkiF6_0),.din(w_dff_A_4vJ2qQSY1_0),.clk(gclk));
	jdff dff_A_IvvnpkiF6_0(.dout(w_dff_A_AyYapmSO7_0),.din(w_dff_A_IvvnpkiF6_0),.clk(gclk));
	jdff dff_A_AyYapmSO7_0(.dout(w_dff_A_HsREqVyM5_0),.din(w_dff_A_AyYapmSO7_0),.clk(gclk));
	jdff dff_A_HsREqVyM5_0(.dout(w_dff_A_WOX5bTVf0_0),.din(w_dff_A_HsREqVyM5_0),.clk(gclk));
	jdff dff_A_WOX5bTVf0_0(.dout(w_dff_A_Z0lg9tPg8_0),.din(w_dff_A_WOX5bTVf0_0),.clk(gclk));
	jdff dff_A_Z0lg9tPg8_0(.dout(w_dff_A_QTMORFDm9_0),.din(w_dff_A_Z0lg9tPg8_0),.clk(gclk));
	jdff dff_A_QTMORFDm9_0(.dout(G552),.din(w_dff_A_QTMORFDm9_0),.clk(gclk));
	jdff dff_A_gHt6hTma0_1(.dout(w_dff_A_nGPHs6QH5_0),.din(w_dff_A_gHt6hTma0_1),.clk(gclk));
	jdff dff_A_nGPHs6QH5_0(.dout(w_dff_A_uOJwQ9EU1_0),.din(w_dff_A_nGPHs6QH5_0),.clk(gclk));
	jdff dff_A_uOJwQ9EU1_0(.dout(w_dff_A_gfcJcOOx0_0),.din(w_dff_A_uOJwQ9EU1_0),.clk(gclk));
	jdff dff_A_gfcJcOOx0_0(.dout(w_dff_A_F7mCBWlE7_0),.din(w_dff_A_gfcJcOOx0_0),.clk(gclk));
	jdff dff_A_F7mCBWlE7_0(.dout(w_dff_A_EBEOMbHW7_0),.din(w_dff_A_F7mCBWlE7_0),.clk(gclk));
	jdff dff_A_EBEOMbHW7_0(.dout(w_dff_A_9JseOFDB8_0),.din(w_dff_A_EBEOMbHW7_0),.clk(gclk));
	jdff dff_A_9JseOFDB8_0(.dout(w_dff_A_o5nw1aGP8_0),.din(w_dff_A_9JseOFDB8_0),.clk(gclk));
	jdff dff_A_o5nw1aGP8_0(.dout(w_dff_A_VnYT1duh6_0),.din(w_dff_A_o5nw1aGP8_0),.clk(gclk));
	jdff dff_A_VnYT1duh6_0(.dout(w_dff_A_oWnjtQHt0_0),.din(w_dff_A_VnYT1duh6_0),.clk(gclk));
	jdff dff_A_oWnjtQHt0_0(.dout(w_dff_A_Xs0om2bb3_0),.din(w_dff_A_oWnjtQHt0_0),.clk(gclk));
	jdff dff_A_Xs0om2bb3_0(.dout(w_dff_A_XxqiivVE8_0),.din(w_dff_A_Xs0om2bb3_0),.clk(gclk));
	jdff dff_A_XxqiivVE8_0(.dout(w_dff_A_Wu7bGLzd4_0),.din(w_dff_A_XxqiivVE8_0),.clk(gclk));
	jdff dff_A_Wu7bGLzd4_0(.dout(w_dff_A_OSeIN3mp3_0),.din(w_dff_A_Wu7bGLzd4_0),.clk(gclk));
	jdff dff_A_OSeIN3mp3_0(.dout(w_dff_A_drHUhbxT6_0),.din(w_dff_A_OSeIN3mp3_0),.clk(gclk));
	jdff dff_A_drHUhbxT6_0(.dout(w_dff_A_YCZBGw692_0),.din(w_dff_A_drHUhbxT6_0),.clk(gclk));
	jdff dff_A_YCZBGw692_0(.dout(w_dff_A_WAA0KjYz8_0),.din(w_dff_A_YCZBGw692_0),.clk(gclk));
	jdff dff_A_WAA0KjYz8_0(.dout(w_dff_A_ab9WmRfo5_0),.din(w_dff_A_WAA0KjYz8_0),.clk(gclk));
	jdff dff_A_ab9WmRfo5_0(.dout(w_dff_A_bHf2jcQN0_0),.din(w_dff_A_ab9WmRfo5_0),.clk(gclk));
	jdff dff_A_bHf2jcQN0_0(.dout(w_dff_A_JwPBoHa24_0),.din(w_dff_A_bHf2jcQN0_0),.clk(gclk));
	jdff dff_A_JwPBoHa24_0(.dout(w_dff_A_mgby5pHw4_0),.din(w_dff_A_JwPBoHa24_0),.clk(gclk));
	jdff dff_A_mgby5pHw4_0(.dout(w_dff_A_LrOop5077_0),.din(w_dff_A_mgby5pHw4_0),.clk(gclk));
	jdff dff_A_LrOop5077_0(.dout(w_dff_A_lyPcdTvj1_0),.din(w_dff_A_LrOop5077_0),.clk(gclk));
	jdff dff_A_lyPcdTvj1_0(.dout(w_dff_A_ZbaFq0o53_0),.din(w_dff_A_lyPcdTvj1_0),.clk(gclk));
	jdff dff_A_ZbaFq0o53_0(.dout(w_dff_A_c8rCM2qO0_0),.din(w_dff_A_ZbaFq0o53_0),.clk(gclk));
	jdff dff_A_c8rCM2qO0_0(.dout(w_dff_A_ZsWwFhcn1_0),.din(w_dff_A_c8rCM2qO0_0),.clk(gclk));
	jdff dff_A_ZsWwFhcn1_0(.dout(w_dff_A_qJWzWsOf1_0),.din(w_dff_A_ZsWwFhcn1_0),.clk(gclk));
	jdff dff_A_qJWzWsOf1_0(.dout(w_dff_A_0cU1KyT65_0),.din(w_dff_A_qJWzWsOf1_0),.clk(gclk));
	jdff dff_A_0cU1KyT65_0(.dout(w_dff_A_tVbzCKHm5_0),.din(w_dff_A_0cU1KyT65_0),.clk(gclk));
	jdff dff_A_tVbzCKHm5_0(.dout(w_dff_A_Izf5pvUg1_0),.din(w_dff_A_tVbzCKHm5_0),.clk(gclk));
	jdff dff_A_Izf5pvUg1_0(.dout(w_dff_A_42cxK4HZ5_0),.din(w_dff_A_Izf5pvUg1_0),.clk(gclk));
	jdff dff_A_42cxK4HZ5_0(.dout(w_dff_A_s2bNsu3r9_0),.din(w_dff_A_42cxK4HZ5_0),.clk(gclk));
	jdff dff_A_s2bNsu3r9_0(.dout(w_dff_A_mKO50t8y6_0),.din(w_dff_A_s2bNsu3r9_0),.clk(gclk));
	jdff dff_A_mKO50t8y6_0(.dout(w_dff_A_NzuRFX0n9_0),.din(w_dff_A_mKO50t8y6_0),.clk(gclk));
	jdff dff_A_NzuRFX0n9_0(.dout(w_dff_A_GeqN5l1K8_0),.din(w_dff_A_NzuRFX0n9_0),.clk(gclk));
	jdff dff_A_GeqN5l1K8_0(.dout(w_dff_A_5dImG5CV1_0),.din(w_dff_A_GeqN5l1K8_0),.clk(gclk));
	jdff dff_A_5dImG5CV1_0(.dout(w_dff_A_GzHL9uzS9_0),.din(w_dff_A_5dImG5CV1_0),.clk(gclk));
	jdff dff_A_GzHL9uzS9_0(.dout(w_dff_A_YCfI5aSf9_0),.din(w_dff_A_GzHL9uzS9_0),.clk(gclk));
	jdff dff_A_YCfI5aSf9_0(.dout(w_dff_A_sj9zNDpl1_0),.din(w_dff_A_YCfI5aSf9_0),.clk(gclk));
	jdff dff_A_sj9zNDpl1_0(.dout(G550),.din(w_dff_A_sj9zNDpl1_0),.clk(gclk));
	jdff dff_A_ljXzS98X0_1(.dout(w_dff_A_nOUr4nCw7_0),.din(w_dff_A_ljXzS98X0_1),.clk(gclk));
	jdff dff_A_nOUr4nCw7_0(.dout(w_dff_A_BJFfyCt24_0),.din(w_dff_A_nOUr4nCw7_0),.clk(gclk));
	jdff dff_A_BJFfyCt24_0(.dout(w_dff_A_NssCCimR2_0),.din(w_dff_A_BJFfyCt24_0),.clk(gclk));
	jdff dff_A_NssCCimR2_0(.dout(w_dff_A_vPecCN0Y5_0),.din(w_dff_A_NssCCimR2_0),.clk(gclk));
	jdff dff_A_vPecCN0Y5_0(.dout(w_dff_A_f71xhcAR6_0),.din(w_dff_A_vPecCN0Y5_0),.clk(gclk));
	jdff dff_A_f71xhcAR6_0(.dout(w_dff_A_PMB24OEl9_0),.din(w_dff_A_f71xhcAR6_0),.clk(gclk));
	jdff dff_A_PMB24OEl9_0(.dout(w_dff_A_gBHfUDLO7_0),.din(w_dff_A_PMB24OEl9_0),.clk(gclk));
	jdff dff_A_gBHfUDLO7_0(.dout(w_dff_A_kwDnf1YH3_0),.din(w_dff_A_gBHfUDLO7_0),.clk(gclk));
	jdff dff_A_kwDnf1YH3_0(.dout(w_dff_A_q01KOlLi4_0),.din(w_dff_A_kwDnf1YH3_0),.clk(gclk));
	jdff dff_A_q01KOlLi4_0(.dout(w_dff_A_t9nSfTNf9_0),.din(w_dff_A_q01KOlLi4_0),.clk(gclk));
	jdff dff_A_t9nSfTNf9_0(.dout(w_dff_A_XqfoWssA8_0),.din(w_dff_A_t9nSfTNf9_0),.clk(gclk));
	jdff dff_A_XqfoWssA8_0(.dout(w_dff_A_BTadeR402_0),.din(w_dff_A_XqfoWssA8_0),.clk(gclk));
	jdff dff_A_BTadeR402_0(.dout(w_dff_A_gX4cizWR7_0),.din(w_dff_A_BTadeR402_0),.clk(gclk));
	jdff dff_A_gX4cizWR7_0(.dout(w_dff_A_GnAbyRYC6_0),.din(w_dff_A_gX4cizWR7_0),.clk(gclk));
	jdff dff_A_GnAbyRYC6_0(.dout(w_dff_A_MhZzZ5S27_0),.din(w_dff_A_GnAbyRYC6_0),.clk(gclk));
	jdff dff_A_MhZzZ5S27_0(.dout(w_dff_A_tdjnYDGm7_0),.din(w_dff_A_MhZzZ5S27_0),.clk(gclk));
	jdff dff_A_tdjnYDGm7_0(.dout(w_dff_A_cRn642oY2_0),.din(w_dff_A_tdjnYDGm7_0),.clk(gclk));
	jdff dff_A_cRn642oY2_0(.dout(w_dff_A_zQQKaLSp1_0),.din(w_dff_A_cRn642oY2_0),.clk(gclk));
	jdff dff_A_zQQKaLSp1_0(.dout(w_dff_A_fQvN1Xop9_0),.din(w_dff_A_zQQKaLSp1_0),.clk(gclk));
	jdff dff_A_fQvN1Xop9_0(.dout(w_dff_A_SIpWHAIr0_0),.din(w_dff_A_fQvN1Xop9_0),.clk(gclk));
	jdff dff_A_SIpWHAIr0_0(.dout(w_dff_A_vCCayale7_0),.din(w_dff_A_SIpWHAIr0_0),.clk(gclk));
	jdff dff_A_vCCayale7_0(.dout(w_dff_A_fCk9bUh52_0),.din(w_dff_A_vCCayale7_0),.clk(gclk));
	jdff dff_A_fCk9bUh52_0(.dout(w_dff_A_tTQS9OPy8_0),.din(w_dff_A_fCk9bUh52_0),.clk(gclk));
	jdff dff_A_tTQS9OPy8_0(.dout(w_dff_A_ut354afT3_0),.din(w_dff_A_tTQS9OPy8_0),.clk(gclk));
	jdff dff_A_ut354afT3_0(.dout(w_dff_A_PTWxS2P06_0),.din(w_dff_A_ut354afT3_0),.clk(gclk));
	jdff dff_A_PTWxS2P06_0(.dout(w_dff_A_O9fVmEKK9_0),.din(w_dff_A_PTWxS2P06_0),.clk(gclk));
	jdff dff_A_O9fVmEKK9_0(.dout(w_dff_A_QwLftZj48_0),.din(w_dff_A_O9fVmEKK9_0),.clk(gclk));
	jdff dff_A_QwLftZj48_0(.dout(w_dff_A_vsW6Xe1B0_0),.din(w_dff_A_QwLftZj48_0),.clk(gclk));
	jdff dff_A_vsW6Xe1B0_0(.dout(w_dff_A_fn55Qm2Y0_0),.din(w_dff_A_vsW6Xe1B0_0),.clk(gclk));
	jdff dff_A_fn55Qm2Y0_0(.dout(w_dff_A_9eAIXyDp9_0),.din(w_dff_A_fn55Qm2Y0_0),.clk(gclk));
	jdff dff_A_9eAIXyDp9_0(.dout(w_dff_A_VI4x1DKG9_0),.din(w_dff_A_9eAIXyDp9_0),.clk(gclk));
	jdff dff_A_VI4x1DKG9_0(.dout(w_dff_A_smGqW4zp3_0),.din(w_dff_A_VI4x1DKG9_0),.clk(gclk));
	jdff dff_A_smGqW4zp3_0(.dout(w_dff_A_bb7P065s6_0),.din(w_dff_A_smGqW4zp3_0),.clk(gclk));
	jdff dff_A_bb7P065s6_0(.dout(w_dff_A_bzO6WC0P9_0),.din(w_dff_A_bb7P065s6_0),.clk(gclk));
	jdff dff_A_bzO6WC0P9_0(.dout(w_dff_A_m2lgcgiZ9_0),.din(w_dff_A_bzO6WC0P9_0),.clk(gclk));
	jdff dff_A_m2lgcgiZ9_0(.dout(w_dff_A_B6JKsWB17_0),.din(w_dff_A_m2lgcgiZ9_0),.clk(gclk));
	jdff dff_A_B6JKsWB17_0(.dout(w_dff_A_EulQXWeM5_0),.din(w_dff_A_B6JKsWB17_0),.clk(gclk));
	jdff dff_A_EulQXWeM5_0(.dout(w_dff_A_YPZ0QiCN5_0),.din(w_dff_A_EulQXWeM5_0),.clk(gclk));
	jdff dff_A_YPZ0QiCN5_0(.dout(G548),.din(w_dff_A_YPZ0QiCN5_0),.clk(gclk));
	jdff dff_A_xShgKWs03_1(.dout(w_dff_A_kjO7M7KU8_0),.din(w_dff_A_xShgKWs03_1),.clk(gclk));
	jdff dff_A_kjO7M7KU8_0(.dout(w_dff_A_pGW84IGQ2_0),.din(w_dff_A_kjO7M7KU8_0),.clk(gclk));
	jdff dff_A_pGW84IGQ2_0(.dout(w_dff_A_1fWjeC0q6_0),.din(w_dff_A_pGW84IGQ2_0),.clk(gclk));
	jdff dff_A_1fWjeC0q6_0(.dout(w_dff_A_5MVLNlnI4_0),.din(w_dff_A_1fWjeC0q6_0),.clk(gclk));
	jdff dff_A_5MVLNlnI4_0(.dout(w_dff_A_wj4bYWy55_0),.din(w_dff_A_5MVLNlnI4_0),.clk(gclk));
	jdff dff_A_wj4bYWy55_0(.dout(w_dff_A_fsKaOxVv5_0),.din(w_dff_A_wj4bYWy55_0),.clk(gclk));
	jdff dff_A_fsKaOxVv5_0(.dout(w_dff_A_Yd3fyowR6_0),.din(w_dff_A_fsKaOxVv5_0),.clk(gclk));
	jdff dff_A_Yd3fyowR6_0(.dout(w_dff_A_4i3Q8WXZ6_0),.din(w_dff_A_Yd3fyowR6_0),.clk(gclk));
	jdff dff_A_4i3Q8WXZ6_0(.dout(w_dff_A_mxIET3BN6_0),.din(w_dff_A_4i3Q8WXZ6_0),.clk(gclk));
	jdff dff_A_mxIET3BN6_0(.dout(w_dff_A_dGalxtaK2_0),.din(w_dff_A_mxIET3BN6_0),.clk(gclk));
	jdff dff_A_dGalxtaK2_0(.dout(w_dff_A_YkbXa5gH2_0),.din(w_dff_A_dGalxtaK2_0),.clk(gclk));
	jdff dff_A_YkbXa5gH2_0(.dout(w_dff_A_lAMTkiGl1_0),.din(w_dff_A_YkbXa5gH2_0),.clk(gclk));
	jdff dff_A_lAMTkiGl1_0(.dout(w_dff_A_P2ywUzQV6_0),.din(w_dff_A_lAMTkiGl1_0),.clk(gclk));
	jdff dff_A_P2ywUzQV6_0(.dout(w_dff_A_WVY41mYz5_0),.din(w_dff_A_P2ywUzQV6_0),.clk(gclk));
	jdff dff_A_WVY41mYz5_0(.dout(w_dff_A_GRi7oGyP1_0),.din(w_dff_A_WVY41mYz5_0),.clk(gclk));
	jdff dff_A_GRi7oGyP1_0(.dout(w_dff_A_C0XZ1sFN3_0),.din(w_dff_A_GRi7oGyP1_0),.clk(gclk));
	jdff dff_A_C0XZ1sFN3_0(.dout(w_dff_A_hi5RjgWL4_0),.din(w_dff_A_C0XZ1sFN3_0),.clk(gclk));
	jdff dff_A_hi5RjgWL4_0(.dout(w_dff_A_A54dNGGp2_0),.din(w_dff_A_hi5RjgWL4_0),.clk(gclk));
	jdff dff_A_A54dNGGp2_0(.dout(w_dff_A_xkBHSLTv2_0),.din(w_dff_A_A54dNGGp2_0),.clk(gclk));
	jdff dff_A_xkBHSLTv2_0(.dout(w_dff_A_9NHPVGUc4_0),.din(w_dff_A_xkBHSLTv2_0),.clk(gclk));
	jdff dff_A_9NHPVGUc4_0(.dout(w_dff_A_gZE3wzeU3_0),.din(w_dff_A_9NHPVGUc4_0),.clk(gclk));
	jdff dff_A_gZE3wzeU3_0(.dout(w_dff_A_8ebbw5fz1_0),.din(w_dff_A_gZE3wzeU3_0),.clk(gclk));
	jdff dff_A_8ebbw5fz1_0(.dout(w_dff_A_rbnwV7Kj3_0),.din(w_dff_A_8ebbw5fz1_0),.clk(gclk));
	jdff dff_A_rbnwV7Kj3_0(.dout(w_dff_A_Eh7rDtQW0_0),.din(w_dff_A_rbnwV7Kj3_0),.clk(gclk));
	jdff dff_A_Eh7rDtQW0_0(.dout(w_dff_A_9SWQ4wJ61_0),.din(w_dff_A_Eh7rDtQW0_0),.clk(gclk));
	jdff dff_A_9SWQ4wJ61_0(.dout(w_dff_A_qf0SmeG78_0),.din(w_dff_A_9SWQ4wJ61_0),.clk(gclk));
	jdff dff_A_qf0SmeG78_0(.dout(w_dff_A_Kkua1hZT1_0),.din(w_dff_A_qf0SmeG78_0),.clk(gclk));
	jdff dff_A_Kkua1hZT1_0(.dout(w_dff_A_1tDb3pRP3_0),.din(w_dff_A_Kkua1hZT1_0),.clk(gclk));
	jdff dff_A_1tDb3pRP3_0(.dout(w_dff_A_surpiXqi2_0),.din(w_dff_A_1tDb3pRP3_0),.clk(gclk));
	jdff dff_A_surpiXqi2_0(.dout(w_dff_A_YXqfAoT57_0),.din(w_dff_A_surpiXqi2_0),.clk(gclk));
	jdff dff_A_YXqfAoT57_0(.dout(w_dff_A_OO1CgwT00_0),.din(w_dff_A_YXqfAoT57_0),.clk(gclk));
	jdff dff_A_OO1CgwT00_0(.dout(w_dff_A_5TJHJzXw2_0),.din(w_dff_A_OO1CgwT00_0),.clk(gclk));
	jdff dff_A_5TJHJzXw2_0(.dout(w_dff_A_LN9KTim27_0),.din(w_dff_A_5TJHJzXw2_0),.clk(gclk));
	jdff dff_A_LN9KTim27_0(.dout(w_dff_A_IzRFCL2H7_0),.din(w_dff_A_LN9KTim27_0),.clk(gclk));
	jdff dff_A_IzRFCL2H7_0(.dout(w_dff_A_GQC5mO9W5_0),.din(w_dff_A_IzRFCL2H7_0),.clk(gclk));
	jdff dff_A_GQC5mO9W5_0(.dout(w_dff_A_DaZSYZLk9_0),.din(w_dff_A_GQC5mO9W5_0),.clk(gclk));
	jdff dff_A_DaZSYZLk9_0(.dout(w_dff_A_Pqw0gOc15_0),.din(w_dff_A_DaZSYZLk9_0),.clk(gclk));
	jdff dff_A_Pqw0gOc15_0(.dout(w_dff_A_3IgEP2Jy8_0),.din(w_dff_A_Pqw0gOc15_0),.clk(gclk));
	jdff dff_A_3IgEP2Jy8_0(.dout(G546),.din(w_dff_A_3IgEP2Jy8_0),.clk(gclk));
	jdff dff_A_38sqavEp5_1(.dout(w_dff_A_Zs3qjdnn7_0),.din(w_dff_A_38sqavEp5_1),.clk(gclk));
	jdff dff_A_Zs3qjdnn7_0(.dout(w_dff_A_1JT9aWSp4_0),.din(w_dff_A_Zs3qjdnn7_0),.clk(gclk));
	jdff dff_A_1JT9aWSp4_0(.dout(w_dff_A_siffhDvj1_0),.din(w_dff_A_1JT9aWSp4_0),.clk(gclk));
	jdff dff_A_siffhDvj1_0(.dout(w_dff_A_4rQIcuBA1_0),.din(w_dff_A_siffhDvj1_0),.clk(gclk));
	jdff dff_A_4rQIcuBA1_0(.dout(w_dff_A_cSmseDur7_0),.din(w_dff_A_4rQIcuBA1_0),.clk(gclk));
	jdff dff_A_cSmseDur7_0(.dout(w_dff_A_H1OnigFP3_0),.din(w_dff_A_cSmseDur7_0),.clk(gclk));
	jdff dff_A_H1OnigFP3_0(.dout(w_dff_A_czdYhQzf2_0),.din(w_dff_A_H1OnigFP3_0),.clk(gclk));
	jdff dff_A_czdYhQzf2_0(.dout(w_dff_A_ryuN8gsJ3_0),.din(w_dff_A_czdYhQzf2_0),.clk(gclk));
	jdff dff_A_ryuN8gsJ3_0(.dout(w_dff_A_pfTH7akb9_0),.din(w_dff_A_ryuN8gsJ3_0),.clk(gclk));
	jdff dff_A_pfTH7akb9_0(.dout(w_dff_A_QVSJHuk56_0),.din(w_dff_A_pfTH7akb9_0),.clk(gclk));
	jdff dff_A_QVSJHuk56_0(.dout(w_dff_A_MJXx3tXE2_0),.din(w_dff_A_QVSJHuk56_0),.clk(gclk));
	jdff dff_A_MJXx3tXE2_0(.dout(w_dff_A_2VMtCcSr6_0),.din(w_dff_A_MJXx3tXE2_0),.clk(gclk));
	jdff dff_A_2VMtCcSr6_0(.dout(w_dff_A_Be2b51nP8_0),.din(w_dff_A_2VMtCcSr6_0),.clk(gclk));
	jdff dff_A_Be2b51nP8_0(.dout(w_dff_A_Phgue6VH0_0),.din(w_dff_A_Be2b51nP8_0),.clk(gclk));
	jdff dff_A_Phgue6VH0_0(.dout(w_dff_A_zNKwNga97_0),.din(w_dff_A_Phgue6VH0_0),.clk(gclk));
	jdff dff_A_zNKwNga97_0(.dout(w_dff_A_l3gqVx2B1_0),.din(w_dff_A_zNKwNga97_0),.clk(gclk));
	jdff dff_A_l3gqVx2B1_0(.dout(w_dff_A_w47ceNUJ4_0),.din(w_dff_A_l3gqVx2B1_0),.clk(gclk));
	jdff dff_A_w47ceNUJ4_0(.dout(w_dff_A_5uyAgXWX0_0),.din(w_dff_A_w47ceNUJ4_0),.clk(gclk));
	jdff dff_A_5uyAgXWX0_0(.dout(w_dff_A_TtWs1HRA1_0),.din(w_dff_A_5uyAgXWX0_0),.clk(gclk));
	jdff dff_A_TtWs1HRA1_0(.dout(w_dff_A_qsKlg1Qx5_0),.din(w_dff_A_TtWs1HRA1_0),.clk(gclk));
	jdff dff_A_qsKlg1Qx5_0(.dout(w_dff_A_vu3d9g8D5_0),.din(w_dff_A_qsKlg1Qx5_0),.clk(gclk));
	jdff dff_A_vu3d9g8D5_0(.dout(w_dff_A_xs121gWN4_0),.din(w_dff_A_vu3d9g8D5_0),.clk(gclk));
	jdff dff_A_xs121gWN4_0(.dout(w_dff_A_XvqHuXFx8_0),.din(w_dff_A_xs121gWN4_0),.clk(gclk));
	jdff dff_A_XvqHuXFx8_0(.dout(w_dff_A_WMIFTPsb4_0),.din(w_dff_A_XvqHuXFx8_0),.clk(gclk));
	jdff dff_A_WMIFTPsb4_0(.dout(w_dff_A_mKcd5Wzp7_0),.din(w_dff_A_WMIFTPsb4_0),.clk(gclk));
	jdff dff_A_mKcd5Wzp7_0(.dout(w_dff_A_Znl8z9bx8_0),.din(w_dff_A_mKcd5Wzp7_0),.clk(gclk));
	jdff dff_A_Znl8z9bx8_0(.dout(w_dff_A_ure21g7j4_0),.din(w_dff_A_Znl8z9bx8_0),.clk(gclk));
	jdff dff_A_ure21g7j4_0(.dout(w_dff_A_eaLZXhEP2_0),.din(w_dff_A_ure21g7j4_0),.clk(gclk));
	jdff dff_A_eaLZXhEP2_0(.dout(w_dff_A_wyt5FgrK6_0),.din(w_dff_A_eaLZXhEP2_0),.clk(gclk));
	jdff dff_A_wyt5FgrK6_0(.dout(w_dff_A_dFcjsN7R2_0),.din(w_dff_A_wyt5FgrK6_0),.clk(gclk));
	jdff dff_A_dFcjsN7R2_0(.dout(w_dff_A_WjliDwrF1_0),.din(w_dff_A_dFcjsN7R2_0),.clk(gclk));
	jdff dff_A_WjliDwrF1_0(.dout(w_dff_A_Yz1i94GP0_0),.din(w_dff_A_WjliDwrF1_0),.clk(gclk));
	jdff dff_A_Yz1i94GP0_0(.dout(w_dff_A_KCOoc4MH6_0),.din(w_dff_A_Yz1i94GP0_0),.clk(gclk));
	jdff dff_A_KCOoc4MH6_0(.dout(w_dff_A_a42OPxXh5_0),.din(w_dff_A_KCOoc4MH6_0),.clk(gclk));
	jdff dff_A_a42OPxXh5_0(.dout(w_dff_A_S39VlzLt6_0),.din(w_dff_A_a42OPxXh5_0),.clk(gclk));
	jdff dff_A_S39VlzLt6_0(.dout(w_dff_A_uWsDV42Q3_0),.din(w_dff_A_S39VlzLt6_0),.clk(gclk));
	jdff dff_A_uWsDV42Q3_0(.dout(w_dff_A_5csQeihD0_0),.din(w_dff_A_uWsDV42Q3_0),.clk(gclk));
	jdff dff_A_5csQeihD0_0(.dout(w_dff_A_qxYRl1AQ1_0),.din(w_dff_A_5csQeihD0_0),.clk(gclk));
	jdff dff_A_qxYRl1AQ1_0(.dout(G544),.din(w_dff_A_qxYRl1AQ1_0),.clk(gclk));
	jdff dff_A_DLdvL5Ht9_1(.dout(w_dff_A_HOcIIMqs8_0),.din(w_dff_A_DLdvL5Ht9_1),.clk(gclk));
	jdff dff_A_HOcIIMqs8_0(.dout(w_dff_A_hoznheuJ8_0),.din(w_dff_A_HOcIIMqs8_0),.clk(gclk));
	jdff dff_A_hoznheuJ8_0(.dout(w_dff_A_rAYN32AO2_0),.din(w_dff_A_hoznheuJ8_0),.clk(gclk));
	jdff dff_A_rAYN32AO2_0(.dout(w_dff_A_rLEFmK6y2_0),.din(w_dff_A_rAYN32AO2_0),.clk(gclk));
	jdff dff_A_rLEFmK6y2_0(.dout(w_dff_A_L6XdCxsM8_0),.din(w_dff_A_rLEFmK6y2_0),.clk(gclk));
	jdff dff_A_L6XdCxsM8_0(.dout(w_dff_A_bWjUG67T1_0),.din(w_dff_A_L6XdCxsM8_0),.clk(gclk));
	jdff dff_A_bWjUG67T1_0(.dout(w_dff_A_O5nDktmS3_0),.din(w_dff_A_bWjUG67T1_0),.clk(gclk));
	jdff dff_A_O5nDktmS3_0(.dout(w_dff_A_FLNitFLc8_0),.din(w_dff_A_O5nDktmS3_0),.clk(gclk));
	jdff dff_A_FLNitFLc8_0(.dout(w_dff_A_tMsHjJkH2_0),.din(w_dff_A_FLNitFLc8_0),.clk(gclk));
	jdff dff_A_tMsHjJkH2_0(.dout(w_dff_A_UUhXu5p53_0),.din(w_dff_A_tMsHjJkH2_0),.clk(gclk));
	jdff dff_A_UUhXu5p53_0(.dout(w_dff_A_2XVEdEIp7_0),.din(w_dff_A_UUhXu5p53_0),.clk(gclk));
	jdff dff_A_2XVEdEIp7_0(.dout(w_dff_A_EpM0sfpu3_0),.din(w_dff_A_2XVEdEIp7_0),.clk(gclk));
	jdff dff_A_EpM0sfpu3_0(.dout(w_dff_A_z2ub1JVL2_0),.din(w_dff_A_EpM0sfpu3_0),.clk(gclk));
	jdff dff_A_z2ub1JVL2_0(.dout(w_dff_A_xjb6HRGR7_0),.din(w_dff_A_z2ub1JVL2_0),.clk(gclk));
	jdff dff_A_xjb6HRGR7_0(.dout(w_dff_A_jngDomR09_0),.din(w_dff_A_xjb6HRGR7_0),.clk(gclk));
	jdff dff_A_jngDomR09_0(.dout(w_dff_A_K9nYleKo0_0),.din(w_dff_A_jngDomR09_0),.clk(gclk));
	jdff dff_A_K9nYleKo0_0(.dout(w_dff_A_YgD4JF749_0),.din(w_dff_A_K9nYleKo0_0),.clk(gclk));
	jdff dff_A_YgD4JF749_0(.dout(w_dff_A_PatGGNCK5_0),.din(w_dff_A_YgD4JF749_0),.clk(gclk));
	jdff dff_A_PatGGNCK5_0(.dout(w_dff_A_dsW7JR7S4_0),.din(w_dff_A_PatGGNCK5_0),.clk(gclk));
	jdff dff_A_dsW7JR7S4_0(.dout(w_dff_A_jAR6E5a07_0),.din(w_dff_A_dsW7JR7S4_0),.clk(gclk));
	jdff dff_A_jAR6E5a07_0(.dout(w_dff_A_bVnPyNSV0_0),.din(w_dff_A_jAR6E5a07_0),.clk(gclk));
	jdff dff_A_bVnPyNSV0_0(.dout(w_dff_A_hwVmDXjr0_0),.din(w_dff_A_bVnPyNSV0_0),.clk(gclk));
	jdff dff_A_hwVmDXjr0_0(.dout(w_dff_A_Kzan7UU56_0),.din(w_dff_A_hwVmDXjr0_0),.clk(gclk));
	jdff dff_A_Kzan7UU56_0(.dout(w_dff_A_yF40Rt5Y4_0),.din(w_dff_A_Kzan7UU56_0),.clk(gclk));
	jdff dff_A_yF40Rt5Y4_0(.dout(w_dff_A_DDAFCUvJ3_0),.din(w_dff_A_yF40Rt5Y4_0),.clk(gclk));
	jdff dff_A_DDAFCUvJ3_0(.dout(w_dff_A_xB6wulfQ6_0),.din(w_dff_A_DDAFCUvJ3_0),.clk(gclk));
	jdff dff_A_xB6wulfQ6_0(.dout(w_dff_A_cNjKZeet2_0),.din(w_dff_A_xB6wulfQ6_0),.clk(gclk));
	jdff dff_A_cNjKZeet2_0(.dout(w_dff_A_28m52jwX9_0),.din(w_dff_A_cNjKZeet2_0),.clk(gclk));
	jdff dff_A_28m52jwX9_0(.dout(w_dff_A_9CZbkAR68_0),.din(w_dff_A_28m52jwX9_0),.clk(gclk));
	jdff dff_A_9CZbkAR68_0(.dout(w_dff_A_qDRc3Jw05_0),.din(w_dff_A_9CZbkAR68_0),.clk(gclk));
	jdff dff_A_qDRc3Jw05_0(.dout(w_dff_A_hxum9Leg2_0),.din(w_dff_A_qDRc3Jw05_0),.clk(gclk));
	jdff dff_A_hxum9Leg2_0(.dout(w_dff_A_CF9t3HuT2_0),.din(w_dff_A_hxum9Leg2_0),.clk(gclk));
	jdff dff_A_CF9t3HuT2_0(.dout(w_dff_A_ceVtjhnF2_0),.din(w_dff_A_CF9t3HuT2_0),.clk(gclk));
	jdff dff_A_ceVtjhnF2_0(.dout(w_dff_A_K4LptOkN3_0),.din(w_dff_A_ceVtjhnF2_0),.clk(gclk));
	jdff dff_A_K4LptOkN3_0(.dout(w_dff_A_U4hyG6aO5_0),.din(w_dff_A_K4LptOkN3_0),.clk(gclk));
	jdff dff_A_U4hyG6aO5_0(.dout(w_dff_A_ImkWfIsC8_0),.din(w_dff_A_U4hyG6aO5_0),.clk(gclk));
	jdff dff_A_ImkWfIsC8_0(.dout(w_dff_A_n0NYp1dL5_0),.din(w_dff_A_ImkWfIsC8_0),.clk(gclk));
	jdff dff_A_n0NYp1dL5_0(.dout(w_dff_A_b9rPRZxf7_0),.din(w_dff_A_n0NYp1dL5_0),.clk(gclk));
	jdff dff_A_b9rPRZxf7_0(.dout(G540),.din(w_dff_A_b9rPRZxf7_0),.clk(gclk));
	jdff dff_A_EW0imUD51_1(.dout(w_dff_A_26C0lEin4_0),.din(w_dff_A_EW0imUD51_1),.clk(gclk));
	jdff dff_A_26C0lEin4_0(.dout(w_dff_A_wINPRdya4_0),.din(w_dff_A_26C0lEin4_0),.clk(gclk));
	jdff dff_A_wINPRdya4_0(.dout(w_dff_A_pXTcFp8K9_0),.din(w_dff_A_wINPRdya4_0),.clk(gclk));
	jdff dff_A_pXTcFp8K9_0(.dout(w_dff_A_t3T7prDM5_0),.din(w_dff_A_pXTcFp8K9_0),.clk(gclk));
	jdff dff_A_t3T7prDM5_0(.dout(w_dff_A_eBpafFru6_0),.din(w_dff_A_t3T7prDM5_0),.clk(gclk));
	jdff dff_A_eBpafFru6_0(.dout(w_dff_A_oryNXrsh3_0),.din(w_dff_A_eBpafFru6_0),.clk(gclk));
	jdff dff_A_oryNXrsh3_0(.dout(w_dff_A_pSLTGfiz8_0),.din(w_dff_A_oryNXrsh3_0),.clk(gclk));
	jdff dff_A_pSLTGfiz8_0(.dout(w_dff_A_tPV5bS8u1_0),.din(w_dff_A_pSLTGfiz8_0),.clk(gclk));
	jdff dff_A_tPV5bS8u1_0(.dout(w_dff_A_GeGU1QUC8_0),.din(w_dff_A_tPV5bS8u1_0),.clk(gclk));
	jdff dff_A_GeGU1QUC8_0(.dout(w_dff_A_XiUMFY6i1_0),.din(w_dff_A_GeGU1QUC8_0),.clk(gclk));
	jdff dff_A_XiUMFY6i1_0(.dout(w_dff_A_w99GgYdx4_0),.din(w_dff_A_XiUMFY6i1_0),.clk(gclk));
	jdff dff_A_w99GgYdx4_0(.dout(w_dff_A_s7QlhHlg1_0),.din(w_dff_A_w99GgYdx4_0),.clk(gclk));
	jdff dff_A_s7QlhHlg1_0(.dout(w_dff_A_Etx7XtMV4_0),.din(w_dff_A_s7QlhHlg1_0),.clk(gclk));
	jdff dff_A_Etx7XtMV4_0(.dout(w_dff_A_lbbHW5266_0),.din(w_dff_A_Etx7XtMV4_0),.clk(gclk));
	jdff dff_A_lbbHW5266_0(.dout(w_dff_A_sKzts2hu5_0),.din(w_dff_A_lbbHW5266_0),.clk(gclk));
	jdff dff_A_sKzts2hu5_0(.dout(w_dff_A_wqyYimta8_0),.din(w_dff_A_sKzts2hu5_0),.clk(gclk));
	jdff dff_A_wqyYimta8_0(.dout(w_dff_A_uU8jEQhe4_0),.din(w_dff_A_wqyYimta8_0),.clk(gclk));
	jdff dff_A_uU8jEQhe4_0(.dout(w_dff_A_YYva5GVY8_0),.din(w_dff_A_uU8jEQhe4_0),.clk(gclk));
	jdff dff_A_YYva5GVY8_0(.dout(w_dff_A_94xw8laE5_0),.din(w_dff_A_YYva5GVY8_0),.clk(gclk));
	jdff dff_A_94xw8laE5_0(.dout(w_dff_A_dILC9Khq9_0),.din(w_dff_A_94xw8laE5_0),.clk(gclk));
	jdff dff_A_dILC9Khq9_0(.dout(w_dff_A_2qdXm90B8_0),.din(w_dff_A_dILC9Khq9_0),.clk(gclk));
	jdff dff_A_2qdXm90B8_0(.dout(w_dff_A_q5P21ugw6_0),.din(w_dff_A_2qdXm90B8_0),.clk(gclk));
	jdff dff_A_q5P21ugw6_0(.dout(w_dff_A_3TlxiIuo9_0),.din(w_dff_A_q5P21ugw6_0),.clk(gclk));
	jdff dff_A_3TlxiIuo9_0(.dout(w_dff_A_01JH3J1W4_0),.din(w_dff_A_3TlxiIuo9_0),.clk(gclk));
	jdff dff_A_01JH3J1W4_0(.dout(w_dff_A_Ril6aFfp9_0),.din(w_dff_A_01JH3J1W4_0),.clk(gclk));
	jdff dff_A_Ril6aFfp9_0(.dout(w_dff_A_FrqJ7RtD0_0),.din(w_dff_A_Ril6aFfp9_0),.clk(gclk));
	jdff dff_A_FrqJ7RtD0_0(.dout(w_dff_A_b8kAt2EB8_0),.din(w_dff_A_FrqJ7RtD0_0),.clk(gclk));
	jdff dff_A_b8kAt2EB8_0(.dout(w_dff_A_eatSQTXx9_0),.din(w_dff_A_b8kAt2EB8_0),.clk(gclk));
	jdff dff_A_eatSQTXx9_0(.dout(w_dff_A_lZiGRDVi9_0),.din(w_dff_A_eatSQTXx9_0),.clk(gclk));
	jdff dff_A_lZiGRDVi9_0(.dout(w_dff_A_PKa4odit5_0),.din(w_dff_A_lZiGRDVi9_0),.clk(gclk));
	jdff dff_A_PKa4odit5_0(.dout(w_dff_A_hzjcbEMe3_0),.din(w_dff_A_PKa4odit5_0),.clk(gclk));
	jdff dff_A_hzjcbEMe3_0(.dout(w_dff_A_JUIwAcP90_0),.din(w_dff_A_hzjcbEMe3_0),.clk(gclk));
	jdff dff_A_JUIwAcP90_0(.dout(w_dff_A_7Zx8ASuy4_0),.din(w_dff_A_JUIwAcP90_0),.clk(gclk));
	jdff dff_A_7Zx8ASuy4_0(.dout(w_dff_A_vAl48w8K5_0),.din(w_dff_A_7Zx8ASuy4_0),.clk(gclk));
	jdff dff_A_vAl48w8K5_0(.dout(w_dff_A_KV5L78DF2_0),.din(w_dff_A_vAl48w8K5_0),.clk(gclk));
	jdff dff_A_KV5L78DF2_0(.dout(w_dff_A_NbQIdvFX0_0),.din(w_dff_A_KV5L78DF2_0),.clk(gclk));
	jdff dff_A_NbQIdvFX0_0(.dout(w_dff_A_jANELNGQ5_0),.din(w_dff_A_NbQIdvFX0_0),.clk(gclk));
	jdff dff_A_jANELNGQ5_0(.dout(w_dff_A_Wg2Zu0QT2_0),.din(w_dff_A_jANELNGQ5_0),.clk(gclk));
	jdff dff_A_Wg2Zu0QT2_0(.dout(G538),.din(w_dff_A_Wg2Zu0QT2_0),.clk(gclk));
	jdff dff_A_pZScGDyA2_1(.dout(w_dff_A_Dz0znsbc8_0),.din(w_dff_A_pZScGDyA2_1),.clk(gclk));
	jdff dff_A_Dz0znsbc8_0(.dout(w_dff_A_LJveWNLP7_0),.din(w_dff_A_Dz0znsbc8_0),.clk(gclk));
	jdff dff_A_LJveWNLP7_0(.dout(w_dff_A_hYlLDHVy5_0),.din(w_dff_A_LJveWNLP7_0),.clk(gclk));
	jdff dff_A_hYlLDHVy5_0(.dout(w_dff_A_oWA8x1w36_0),.din(w_dff_A_hYlLDHVy5_0),.clk(gclk));
	jdff dff_A_oWA8x1w36_0(.dout(w_dff_A_4hhUBxVE4_0),.din(w_dff_A_oWA8x1w36_0),.clk(gclk));
	jdff dff_A_4hhUBxVE4_0(.dout(w_dff_A_Sfop3p7p8_0),.din(w_dff_A_4hhUBxVE4_0),.clk(gclk));
	jdff dff_A_Sfop3p7p8_0(.dout(w_dff_A_PUMgXenJ7_0),.din(w_dff_A_Sfop3p7p8_0),.clk(gclk));
	jdff dff_A_PUMgXenJ7_0(.dout(w_dff_A_uc13hQny4_0),.din(w_dff_A_PUMgXenJ7_0),.clk(gclk));
	jdff dff_A_uc13hQny4_0(.dout(w_dff_A_toIw3Va90_0),.din(w_dff_A_uc13hQny4_0),.clk(gclk));
	jdff dff_A_toIw3Va90_0(.dout(w_dff_A_OK1tV9WE5_0),.din(w_dff_A_toIw3Va90_0),.clk(gclk));
	jdff dff_A_OK1tV9WE5_0(.dout(w_dff_A_e6k42ZkM0_0),.din(w_dff_A_OK1tV9WE5_0),.clk(gclk));
	jdff dff_A_e6k42ZkM0_0(.dout(w_dff_A_1uZx7O7X2_0),.din(w_dff_A_e6k42ZkM0_0),.clk(gclk));
	jdff dff_A_1uZx7O7X2_0(.dout(w_dff_A_SWTDTC4A3_0),.din(w_dff_A_1uZx7O7X2_0),.clk(gclk));
	jdff dff_A_SWTDTC4A3_0(.dout(w_dff_A_ATjbpP5w8_0),.din(w_dff_A_SWTDTC4A3_0),.clk(gclk));
	jdff dff_A_ATjbpP5w8_0(.dout(w_dff_A_F7bHCY530_0),.din(w_dff_A_ATjbpP5w8_0),.clk(gclk));
	jdff dff_A_F7bHCY530_0(.dout(w_dff_A_Bw9tKLlx7_0),.din(w_dff_A_F7bHCY530_0),.clk(gclk));
	jdff dff_A_Bw9tKLlx7_0(.dout(w_dff_A_5aPjWhOc5_0),.din(w_dff_A_Bw9tKLlx7_0),.clk(gclk));
	jdff dff_A_5aPjWhOc5_0(.dout(w_dff_A_OgSL8DjQ5_0),.din(w_dff_A_5aPjWhOc5_0),.clk(gclk));
	jdff dff_A_OgSL8DjQ5_0(.dout(w_dff_A_7phPNwun4_0),.din(w_dff_A_OgSL8DjQ5_0),.clk(gclk));
	jdff dff_A_7phPNwun4_0(.dout(w_dff_A_Gboaby8G3_0),.din(w_dff_A_7phPNwun4_0),.clk(gclk));
	jdff dff_A_Gboaby8G3_0(.dout(w_dff_A_RTNloDsB1_0),.din(w_dff_A_Gboaby8G3_0),.clk(gclk));
	jdff dff_A_RTNloDsB1_0(.dout(w_dff_A_mZPJaOnL3_0),.din(w_dff_A_RTNloDsB1_0),.clk(gclk));
	jdff dff_A_mZPJaOnL3_0(.dout(w_dff_A_cb0gjv0B3_0),.din(w_dff_A_mZPJaOnL3_0),.clk(gclk));
	jdff dff_A_cb0gjv0B3_0(.dout(w_dff_A_srQ33LFz4_0),.din(w_dff_A_cb0gjv0B3_0),.clk(gclk));
	jdff dff_A_srQ33LFz4_0(.dout(w_dff_A_UAaU5ua07_0),.din(w_dff_A_srQ33LFz4_0),.clk(gclk));
	jdff dff_A_UAaU5ua07_0(.dout(w_dff_A_SESMrgmB8_0),.din(w_dff_A_UAaU5ua07_0),.clk(gclk));
	jdff dff_A_SESMrgmB8_0(.dout(w_dff_A_ttbdKH5X0_0),.din(w_dff_A_SESMrgmB8_0),.clk(gclk));
	jdff dff_A_ttbdKH5X0_0(.dout(w_dff_A_w0xWYzyw2_0),.din(w_dff_A_ttbdKH5X0_0),.clk(gclk));
	jdff dff_A_w0xWYzyw2_0(.dout(w_dff_A_OuQnam1G8_0),.din(w_dff_A_w0xWYzyw2_0),.clk(gclk));
	jdff dff_A_OuQnam1G8_0(.dout(w_dff_A_rzB2tTdl4_0),.din(w_dff_A_OuQnam1G8_0),.clk(gclk));
	jdff dff_A_rzB2tTdl4_0(.dout(w_dff_A_74XDc4Gf3_0),.din(w_dff_A_rzB2tTdl4_0),.clk(gclk));
	jdff dff_A_74XDc4Gf3_0(.dout(w_dff_A_Hysq3mT26_0),.din(w_dff_A_74XDc4Gf3_0),.clk(gclk));
	jdff dff_A_Hysq3mT26_0(.dout(w_dff_A_x2js2btP5_0),.din(w_dff_A_Hysq3mT26_0),.clk(gclk));
	jdff dff_A_x2js2btP5_0(.dout(w_dff_A_8qxLEd5G3_0),.din(w_dff_A_x2js2btP5_0),.clk(gclk));
	jdff dff_A_8qxLEd5G3_0(.dout(w_dff_A_GoKdhjaH3_0),.din(w_dff_A_8qxLEd5G3_0),.clk(gclk));
	jdff dff_A_GoKdhjaH3_0(.dout(w_dff_A_xid1jguN1_0),.din(w_dff_A_GoKdhjaH3_0),.clk(gclk));
	jdff dff_A_xid1jguN1_0(.dout(w_dff_A_nvwqbOaQ0_0),.din(w_dff_A_xid1jguN1_0),.clk(gclk));
	jdff dff_A_nvwqbOaQ0_0(.dout(w_dff_A_uAzFVU012_0),.din(w_dff_A_nvwqbOaQ0_0),.clk(gclk));
	jdff dff_A_uAzFVU012_0(.dout(G536),.din(w_dff_A_uAzFVU012_0),.clk(gclk));
	jdff dff_A_s9CBI2X99_1(.dout(w_dff_A_5j4X6org3_0),.din(w_dff_A_s9CBI2X99_1),.clk(gclk));
	jdff dff_A_5j4X6org3_0(.dout(w_dff_A_o8iTZWdY2_0),.din(w_dff_A_5j4X6org3_0),.clk(gclk));
	jdff dff_A_o8iTZWdY2_0(.dout(w_dff_A_P4vQ4pzD5_0),.din(w_dff_A_o8iTZWdY2_0),.clk(gclk));
	jdff dff_A_P4vQ4pzD5_0(.dout(w_dff_A_unbKZawH9_0),.din(w_dff_A_P4vQ4pzD5_0),.clk(gclk));
	jdff dff_A_unbKZawH9_0(.dout(w_dff_A_35C307ns7_0),.din(w_dff_A_unbKZawH9_0),.clk(gclk));
	jdff dff_A_35C307ns7_0(.dout(w_dff_A_tV1Kezob9_0),.din(w_dff_A_35C307ns7_0),.clk(gclk));
	jdff dff_A_tV1Kezob9_0(.dout(w_dff_A_REkXp1r70_0),.din(w_dff_A_tV1Kezob9_0),.clk(gclk));
	jdff dff_A_REkXp1r70_0(.dout(w_dff_A_WUrqD82e6_0),.din(w_dff_A_REkXp1r70_0),.clk(gclk));
	jdff dff_A_WUrqD82e6_0(.dout(w_dff_A_5x2nP9jM6_0),.din(w_dff_A_WUrqD82e6_0),.clk(gclk));
	jdff dff_A_5x2nP9jM6_0(.dout(w_dff_A_GzdYYtnu4_0),.din(w_dff_A_5x2nP9jM6_0),.clk(gclk));
	jdff dff_A_GzdYYtnu4_0(.dout(w_dff_A_M8ltJ3DN2_0),.din(w_dff_A_GzdYYtnu4_0),.clk(gclk));
	jdff dff_A_M8ltJ3DN2_0(.dout(w_dff_A_YAhXaJ6b0_0),.din(w_dff_A_M8ltJ3DN2_0),.clk(gclk));
	jdff dff_A_YAhXaJ6b0_0(.dout(w_dff_A_586ElPPZ2_0),.din(w_dff_A_YAhXaJ6b0_0),.clk(gclk));
	jdff dff_A_586ElPPZ2_0(.dout(w_dff_A_rS5yQATm5_0),.din(w_dff_A_586ElPPZ2_0),.clk(gclk));
	jdff dff_A_rS5yQATm5_0(.dout(w_dff_A_yI3DnthI3_0),.din(w_dff_A_rS5yQATm5_0),.clk(gclk));
	jdff dff_A_yI3DnthI3_0(.dout(w_dff_A_0OP8pJvZ1_0),.din(w_dff_A_yI3DnthI3_0),.clk(gclk));
	jdff dff_A_0OP8pJvZ1_0(.dout(w_dff_A_m5xsyH0s3_0),.din(w_dff_A_0OP8pJvZ1_0),.clk(gclk));
	jdff dff_A_m5xsyH0s3_0(.dout(w_dff_A_B2gofKCl5_0),.din(w_dff_A_m5xsyH0s3_0),.clk(gclk));
	jdff dff_A_B2gofKCl5_0(.dout(w_dff_A_H6WoT1RM1_0),.din(w_dff_A_B2gofKCl5_0),.clk(gclk));
	jdff dff_A_H6WoT1RM1_0(.dout(w_dff_A_LvF4yQfq3_0),.din(w_dff_A_H6WoT1RM1_0),.clk(gclk));
	jdff dff_A_LvF4yQfq3_0(.dout(w_dff_A_nE6UP5G59_0),.din(w_dff_A_LvF4yQfq3_0),.clk(gclk));
	jdff dff_A_nE6UP5G59_0(.dout(w_dff_A_APzV3JU79_0),.din(w_dff_A_nE6UP5G59_0),.clk(gclk));
	jdff dff_A_APzV3JU79_0(.dout(w_dff_A_FdlJiHep2_0),.din(w_dff_A_APzV3JU79_0),.clk(gclk));
	jdff dff_A_FdlJiHep2_0(.dout(w_dff_A_sumutRLf2_0),.din(w_dff_A_FdlJiHep2_0),.clk(gclk));
	jdff dff_A_sumutRLf2_0(.dout(w_dff_A_Fmc8i1Op4_0),.din(w_dff_A_sumutRLf2_0),.clk(gclk));
	jdff dff_A_Fmc8i1Op4_0(.dout(w_dff_A_saZHOdSU0_0),.din(w_dff_A_Fmc8i1Op4_0),.clk(gclk));
	jdff dff_A_saZHOdSU0_0(.dout(w_dff_A_3GP0EtA17_0),.din(w_dff_A_saZHOdSU0_0),.clk(gclk));
	jdff dff_A_3GP0EtA17_0(.dout(w_dff_A_4GEYyXez1_0),.din(w_dff_A_3GP0EtA17_0),.clk(gclk));
	jdff dff_A_4GEYyXez1_0(.dout(w_dff_A_VxlFqlQU1_0),.din(w_dff_A_4GEYyXez1_0),.clk(gclk));
	jdff dff_A_VxlFqlQU1_0(.dout(w_dff_A_AUPmesxs4_0),.din(w_dff_A_VxlFqlQU1_0),.clk(gclk));
	jdff dff_A_AUPmesxs4_0(.dout(w_dff_A_8xehiPFf6_0),.din(w_dff_A_AUPmesxs4_0),.clk(gclk));
	jdff dff_A_8xehiPFf6_0(.dout(w_dff_A_zWkRpF5C4_0),.din(w_dff_A_8xehiPFf6_0),.clk(gclk));
	jdff dff_A_zWkRpF5C4_0(.dout(w_dff_A_LM15TwUm5_0),.din(w_dff_A_zWkRpF5C4_0),.clk(gclk));
	jdff dff_A_LM15TwUm5_0(.dout(w_dff_A_YVNYLe6J0_0),.din(w_dff_A_LM15TwUm5_0),.clk(gclk));
	jdff dff_A_YVNYLe6J0_0(.dout(w_dff_A_ijOsg7Oa3_0),.din(w_dff_A_YVNYLe6J0_0),.clk(gclk));
	jdff dff_A_ijOsg7Oa3_0(.dout(w_dff_A_EXZmuuH19_0),.din(w_dff_A_ijOsg7Oa3_0),.clk(gclk));
	jdff dff_A_EXZmuuH19_0(.dout(w_dff_A_3zZ4H4rX1_0),.din(w_dff_A_EXZmuuH19_0),.clk(gclk));
	jdff dff_A_3zZ4H4rX1_0(.dout(w_dff_A_FmHOqaXh5_0),.din(w_dff_A_3zZ4H4rX1_0),.clk(gclk));
	jdff dff_A_FmHOqaXh5_0(.dout(G534),.din(w_dff_A_FmHOqaXh5_0),.clk(gclk));
	jdff dff_A_ltJWpPGm4_1(.dout(w_dff_A_bTj4dEHH2_0),.din(w_dff_A_ltJWpPGm4_1),.clk(gclk));
	jdff dff_A_bTj4dEHH2_0(.dout(w_dff_A_n8ApaKVc7_0),.din(w_dff_A_bTj4dEHH2_0),.clk(gclk));
	jdff dff_A_n8ApaKVc7_0(.dout(w_dff_A_KcfK5MyF3_0),.din(w_dff_A_n8ApaKVc7_0),.clk(gclk));
	jdff dff_A_KcfK5MyF3_0(.dout(w_dff_A_pE7lSduZ5_0),.din(w_dff_A_KcfK5MyF3_0),.clk(gclk));
	jdff dff_A_pE7lSduZ5_0(.dout(w_dff_A_YiQbfKdg3_0),.din(w_dff_A_pE7lSduZ5_0),.clk(gclk));
	jdff dff_A_YiQbfKdg3_0(.dout(w_dff_A_D69IDZIi1_0),.din(w_dff_A_YiQbfKdg3_0),.clk(gclk));
	jdff dff_A_D69IDZIi1_0(.dout(w_dff_A_yRF65uNC9_0),.din(w_dff_A_D69IDZIi1_0),.clk(gclk));
	jdff dff_A_yRF65uNC9_0(.dout(w_dff_A_YjkzyKuc2_0),.din(w_dff_A_yRF65uNC9_0),.clk(gclk));
	jdff dff_A_YjkzyKuc2_0(.dout(w_dff_A_TWTwWK5n6_0),.din(w_dff_A_YjkzyKuc2_0),.clk(gclk));
	jdff dff_A_TWTwWK5n6_0(.dout(w_dff_A_yPgFgPSA9_0),.din(w_dff_A_TWTwWK5n6_0),.clk(gclk));
	jdff dff_A_yPgFgPSA9_0(.dout(w_dff_A_sGQUdmmi7_0),.din(w_dff_A_yPgFgPSA9_0),.clk(gclk));
	jdff dff_A_sGQUdmmi7_0(.dout(w_dff_A_i6TZp9aW1_0),.din(w_dff_A_sGQUdmmi7_0),.clk(gclk));
	jdff dff_A_i6TZp9aW1_0(.dout(w_dff_A_N7DxbTFP1_0),.din(w_dff_A_i6TZp9aW1_0),.clk(gclk));
	jdff dff_A_N7DxbTFP1_0(.dout(w_dff_A_PP9eikLr5_0),.din(w_dff_A_N7DxbTFP1_0),.clk(gclk));
	jdff dff_A_PP9eikLr5_0(.dout(w_dff_A_VLGLq12v6_0),.din(w_dff_A_PP9eikLr5_0),.clk(gclk));
	jdff dff_A_VLGLq12v6_0(.dout(w_dff_A_Wu7GTIuA1_0),.din(w_dff_A_VLGLq12v6_0),.clk(gclk));
	jdff dff_A_Wu7GTIuA1_0(.dout(w_dff_A_EY5H5PSt2_0),.din(w_dff_A_Wu7GTIuA1_0),.clk(gclk));
	jdff dff_A_EY5H5PSt2_0(.dout(w_dff_A_VTdLg4rc3_0),.din(w_dff_A_EY5H5PSt2_0),.clk(gclk));
	jdff dff_A_VTdLg4rc3_0(.dout(w_dff_A_ZSDcuK9b9_0),.din(w_dff_A_VTdLg4rc3_0),.clk(gclk));
	jdff dff_A_ZSDcuK9b9_0(.dout(w_dff_A_hMNeXxaf3_0),.din(w_dff_A_ZSDcuK9b9_0),.clk(gclk));
	jdff dff_A_hMNeXxaf3_0(.dout(w_dff_A_Yvj76dXK0_0),.din(w_dff_A_hMNeXxaf3_0),.clk(gclk));
	jdff dff_A_Yvj76dXK0_0(.dout(w_dff_A_Oxxn2wMM0_0),.din(w_dff_A_Yvj76dXK0_0),.clk(gclk));
	jdff dff_A_Oxxn2wMM0_0(.dout(w_dff_A_73939TPZ4_0),.din(w_dff_A_Oxxn2wMM0_0),.clk(gclk));
	jdff dff_A_73939TPZ4_0(.dout(w_dff_A_cCQA6j7L3_0),.din(w_dff_A_73939TPZ4_0),.clk(gclk));
	jdff dff_A_cCQA6j7L3_0(.dout(w_dff_A_PF9gHu5I0_0),.din(w_dff_A_cCQA6j7L3_0),.clk(gclk));
	jdff dff_A_PF9gHu5I0_0(.dout(w_dff_A_PjWrK1Ch8_0),.din(w_dff_A_PF9gHu5I0_0),.clk(gclk));
	jdff dff_A_PjWrK1Ch8_0(.dout(w_dff_A_bz0hL5Dy8_0),.din(w_dff_A_PjWrK1Ch8_0),.clk(gclk));
	jdff dff_A_bz0hL5Dy8_0(.dout(w_dff_A_PF4f4Foc7_0),.din(w_dff_A_bz0hL5Dy8_0),.clk(gclk));
	jdff dff_A_PF4f4Foc7_0(.dout(w_dff_A_TmwLJyQp7_0),.din(w_dff_A_PF4f4Foc7_0),.clk(gclk));
	jdff dff_A_TmwLJyQp7_0(.dout(w_dff_A_nJBGiABp0_0),.din(w_dff_A_TmwLJyQp7_0),.clk(gclk));
	jdff dff_A_nJBGiABp0_0(.dout(w_dff_A_orQpsPhc2_0),.din(w_dff_A_nJBGiABp0_0),.clk(gclk));
	jdff dff_A_orQpsPhc2_0(.dout(w_dff_A_7A4MWDON8_0),.din(w_dff_A_orQpsPhc2_0),.clk(gclk));
	jdff dff_A_7A4MWDON8_0(.dout(w_dff_A_vbzK9DWS0_0),.din(w_dff_A_7A4MWDON8_0),.clk(gclk));
	jdff dff_A_vbzK9DWS0_0(.dout(w_dff_A_SrlVGlhG1_0),.din(w_dff_A_vbzK9DWS0_0),.clk(gclk));
	jdff dff_A_SrlVGlhG1_0(.dout(w_dff_A_6cxfcSvs8_0),.din(w_dff_A_SrlVGlhG1_0),.clk(gclk));
	jdff dff_A_6cxfcSvs8_0(.dout(w_dff_A_hGP8F4OX5_0),.din(w_dff_A_6cxfcSvs8_0),.clk(gclk));
	jdff dff_A_hGP8F4OX5_0(.dout(w_dff_A_i6mFKTzI7_0),.din(w_dff_A_hGP8F4OX5_0),.clk(gclk));
	jdff dff_A_i6mFKTzI7_0(.dout(w_dff_A_KDNPJ6ir4_0),.din(w_dff_A_i6mFKTzI7_0),.clk(gclk));
	jdff dff_A_KDNPJ6ir4_0(.dout(G532),.din(w_dff_A_KDNPJ6ir4_0),.clk(gclk));
	jdff dff_A_YJS1iCK09_1(.dout(w_dff_A_TbVdD3vB2_0),.din(w_dff_A_YJS1iCK09_1),.clk(gclk));
	jdff dff_A_TbVdD3vB2_0(.dout(w_dff_A_NnG0DdCZ7_0),.din(w_dff_A_TbVdD3vB2_0),.clk(gclk));
	jdff dff_A_NnG0DdCZ7_0(.dout(w_dff_A_0Mw1IltL6_0),.din(w_dff_A_NnG0DdCZ7_0),.clk(gclk));
	jdff dff_A_0Mw1IltL6_0(.dout(w_dff_A_KMqhhc703_0),.din(w_dff_A_0Mw1IltL6_0),.clk(gclk));
	jdff dff_A_KMqhhc703_0(.dout(w_dff_A_UgpTv6zH6_0),.din(w_dff_A_KMqhhc703_0),.clk(gclk));
	jdff dff_A_UgpTv6zH6_0(.dout(w_dff_A_gagAgT4D0_0),.din(w_dff_A_UgpTv6zH6_0),.clk(gclk));
	jdff dff_A_gagAgT4D0_0(.dout(w_dff_A_X9OInrxT8_0),.din(w_dff_A_gagAgT4D0_0),.clk(gclk));
	jdff dff_A_X9OInrxT8_0(.dout(w_dff_A_edachBqU8_0),.din(w_dff_A_X9OInrxT8_0),.clk(gclk));
	jdff dff_A_edachBqU8_0(.dout(w_dff_A_o8L9tTTP2_0),.din(w_dff_A_edachBqU8_0),.clk(gclk));
	jdff dff_A_o8L9tTTP2_0(.dout(w_dff_A_t5yS1FMO9_0),.din(w_dff_A_o8L9tTTP2_0),.clk(gclk));
	jdff dff_A_t5yS1FMO9_0(.dout(w_dff_A_2QeghzNY7_0),.din(w_dff_A_t5yS1FMO9_0),.clk(gclk));
	jdff dff_A_2QeghzNY7_0(.dout(w_dff_A_uiJ2ECX90_0),.din(w_dff_A_2QeghzNY7_0),.clk(gclk));
	jdff dff_A_uiJ2ECX90_0(.dout(w_dff_A_ZESKld5F3_0),.din(w_dff_A_uiJ2ECX90_0),.clk(gclk));
	jdff dff_A_ZESKld5F3_0(.dout(w_dff_A_qddnKWYm6_0),.din(w_dff_A_ZESKld5F3_0),.clk(gclk));
	jdff dff_A_qddnKWYm6_0(.dout(w_dff_A_QmZJafKr2_0),.din(w_dff_A_qddnKWYm6_0),.clk(gclk));
	jdff dff_A_QmZJafKr2_0(.dout(w_dff_A_Ia459EA71_0),.din(w_dff_A_QmZJafKr2_0),.clk(gclk));
	jdff dff_A_Ia459EA71_0(.dout(w_dff_A_P4GwI2Vz9_0),.din(w_dff_A_Ia459EA71_0),.clk(gclk));
	jdff dff_A_P4GwI2Vz9_0(.dout(w_dff_A_8dHBC7Oa4_0),.din(w_dff_A_P4GwI2Vz9_0),.clk(gclk));
	jdff dff_A_8dHBC7Oa4_0(.dout(w_dff_A_1CPyePqK3_0),.din(w_dff_A_8dHBC7Oa4_0),.clk(gclk));
	jdff dff_A_1CPyePqK3_0(.dout(w_dff_A_XVkRIzdC1_0),.din(w_dff_A_1CPyePqK3_0),.clk(gclk));
	jdff dff_A_XVkRIzdC1_0(.dout(w_dff_A_17zQs4O20_0),.din(w_dff_A_XVkRIzdC1_0),.clk(gclk));
	jdff dff_A_17zQs4O20_0(.dout(w_dff_A_2ih7ywQW7_0),.din(w_dff_A_17zQs4O20_0),.clk(gclk));
	jdff dff_A_2ih7ywQW7_0(.dout(w_dff_A_3VKPvNBR8_0),.din(w_dff_A_2ih7ywQW7_0),.clk(gclk));
	jdff dff_A_3VKPvNBR8_0(.dout(w_dff_A_wJWYmI1s0_0),.din(w_dff_A_3VKPvNBR8_0),.clk(gclk));
	jdff dff_A_wJWYmI1s0_0(.dout(w_dff_A_46ZLSEbS5_0),.din(w_dff_A_wJWYmI1s0_0),.clk(gclk));
	jdff dff_A_46ZLSEbS5_0(.dout(w_dff_A_ejOkQggK5_0),.din(w_dff_A_46ZLSEbS5_0),.clk(gclk));
	jdff dff_A_ejOkQggK5_0(.dout(w_dff_A_S9o3y3cQ1_0),.din(w_dff_A_ejOkQggK5_0),.clk(gclk));
	jdff dff_A_S9o3y3cQ1_0(.dout(w_dff_A_jO09T9Oj6_0),.din(w_dff_A_S9o3y3cQ1_0),.clk(gclk));
	jdff dff_A_jO09T9Oj6_0(.dout(w_dff_A_s1PEjzWx4_0),.din(w_dff_A_jO09T9Oj6_0),.clk(gclk));
	jdff dff_A_s1PEjzWx4_0(.dout(w_dff_A_J4QPgZ4j4_0),.din(w_dff_A_s1PEjzWx4_0),.clk(gclk));
	jdff dff_A_J4QPgZ4j4_0(.dout(w_dff_A_UyQeu1gk3_0),.din(w_dff_A_J4QPgZ4j4_0),.clk(gclk));
	jdff dff_A_UyQeu1gk3_0(.dout(w_dff_A_jf9T34HT1_0),.din(w_dff_A_UyQeu1gk3_0),.clk(gclk));
	jdff dff_A_jf9T34HT1_0(.dout(w_dff_A_0lHXl7NV9_0),.din(w_dff_A_jf9T34HT1_0),.clk(gclk));
	jdff dff_A_0lHXl7NV9_0(.dout(w_dff_A_EV38FxhT5_0),.din(w_dff_A_0lHXl7NV9_0),.clk(gclk));
	jdff dff_A_EV38FxhT5_0(.dout(w_dff_A_PKVQcffY0_0),.din(w_dff_A_EV38FxhT5_0),.clk(gclk));
	jdff dff_A_PKVQcffY0_0(.dout(w_dff_A_8hyZE7070_0),.din(w_dff_A_PKVQcffY0_0),.clk(gclk));
	jdff dff_A_8hyZE7070_0(.dout(w_dff_A_0FAgAEJO9_0),.din(w_dff_A_8hyZE7070_0),.clk(gclk));
	jdff dff_A_0FAgAEJO9_0(.dout(w_dff_A_SnNak6mp8_0),.din(w_dff_A_0FAgAEJO9_0),.clk(gclk));
	jdff dff_A_SnNak6mp8_0(.dout(G530),.din(w_dff_A_SnNak6mp8_0),.clk(gclk));
	jdff dff_A_ThUKi2cH2_1(.dout(w_dff_A_xn8OdA137_0),.din(w_dff_A_ThUKi2cH2_1),.clk(gclk));
	jdff dff_A_xn8OdA137_0(.dout(w_dff_A_VX6DQ02v2_0),.din(w_dff_A_xn8OdA137_0),.clk(gclk));
	jdff dff_A_VX6DQ02v2_0(.dout(w_dff_A_qQFbfMUI1_0),.din(w_dff_A_VX6DQ02v2_0),.clk(gclk));
	jdff dff_A_qQFbfMUI1_0(.dout(w_dff_A_SZZlzdoY1_0),.din(w_dff_A_qQFbfMUI1_0),.clk(gclk));
	jdff dff_A_SZZlzdoY1_0(.dout(w_dff_A_9x1ZqXLj1_0),.din(w_dff_A_SZZlzdoY1_0),.clk(gclk));
	jdff dff_A_9x1ZqXLj1_0(.dout(w_dff_A_lZ8gwEzV6_0),.din(w_dff_A_9x1ZqXLj1_0),.clk(gclk));
	jdff dff_A_lZ8gwEzV6_0(.dout(w_dff_A_TTy78zse9_0),.din(w_dff_A_lZ8gwEzV6_0),.clk(gclk));
	jdff dff_A_TTy78zse9_0(.dout(w_dff_A_dkYbxvAD5_0),.din(w_dff_A_TTy78zse9_0),.clk(gclk));
	jdff dff_A_dkYbxvAD5_0(.dout(w_dff_A_rVubgCGZ7_0),.din(w_dff_A_dkYbxvAD5_0),.clk(gclk));
	jdff dff_A_rVubgCGZ7_0(.dout(w_dff_A_u0KJr7cm1_0),.din(w_dff_A_rVubgCGZ7_0),.clk(gclk));
	jdff dff_A_u0KJr7cm1_0(.dout(w_dff_A_iHkEg4030_0),.din(w_dff_A_u0KJr7cm1_0),.clk(gclk));
	jdff dff_A_iHkEg4030_0(.dout(w_dff_A_67zJikhZ5_0),.din(w_dff_A_iHkEg4030_0),.clk(gclk));
	jdff dff_A_67zJikhZ5_0(.dout(w_dff_A_ARQmbsby9_0),.din(w_dff_A_67zJikhZ5_0),.clk(gclk));
	jdff dff_A_ARQmbsby9_0(.dout(w_dff_A_SvRG6qyz2_0),.din(w_dff_A_ARQmbsby9_0),.clk(gclk));
	jdff dff_A_SvRG6qyz2_0(.dout(w_dff_A_hS4mnYRb5_0),.din(w_dff_A_SvRG6qyz2_0),.clk(gclk));
	jdff dff_A_hS4mnYRb5_0(.dout(w_dff_A_UmqymFCp1_0),.din(w_dff_A_hS4mnYRb5_0),.clk(gclk));
	jdff dff_A_UmqymFCp1_0(.dout(w_dff_A_uCk6lHbm7_0),.din(w_dff_A_UmqymFCp1_0),.clk(gclk));
	jdff dff_A_uCk6lHbm7_0(.dout(w_dff_A_OR48rN5f0_0),.din(w_dff_A_uCk6lHbm7_0),.clk(gclk));
	jdff dff_A_OR48rN5f0_0(.dout(w_dff_A_9RxGd0mk4_0),.din(w_dff_A_OR48rN5f0_0),.clk(gclk));
	jdff dff_A_9RxGd0mk4_0(.dout(w_dff_A_0t1bdfl26_0),.din(w_dff_A_9RxGd0mk4_0),.clk(gclk));
	jdff dff_A_0t1bdfl26_0(.dout(w_dff_A_VhCp261p1_0),.din(w_dff_A_0t1bdfl26_0),.clk(gclk));
	jdff dff_A_VhCp261p1_0(.dout(w_dff_A_ILBL7SRY2_0),.din(w_dff_A_VhCp261p1_0),.clk(gclk));
	jdff dff_A_ILBL7SRY2_0(.dout(w_dff_A_j3mpOVkK7_0),.din(w_dff_A_ILBL7SRY2_0),.clk(gclk));
	jdff dff_A_j3mpOVkK7_0(.dout(w_dff_A_2AhICZnV6_0),.din(w_dff_A_j3mpOVkK7_0),.clk(gclk));
	jdff dff_A_2AhICZnV6_0(.dout(w_dff_A_Xqm8grg42_0),.din(w_dff_A_2AhICZnV6_0),.clk(gclk));
	jdff dff_A_Xqm8grg42_0(.dout(w_dff_A_byw5h8b02_0),.din(w_dff_A_Xqm8grg42_0),.clk(gclk));
	jdff dff_A_byw5h8b02_0(.dout(w_dff_A_ftFp8D6W9_0),.din(w_dff_A_byw5h8b02_0),.clk(gclk));
	jdff dff_A_ftFp8D6W9_0(.dout(w_dff_A_j2sNVIHr0_0),.din(w_dff_A_ftFp8D6W9_0),.clk(gclk));
	jdff dff_A_j2sNVIHr0_0(.dout(w_dff_A_8nDB3CRG2_0),.din(w_dff_A_j2sNVIHr0_0),.clk(gclk));
	jdff dff_A_8nDB3CRG2_0(.dout(w_dff_A_B5AJLaOR1_0),.din(w_dff_A_8nDB3CRG2_0),.clk(gclk));
	jdff dff_A_B5AJLaOR1_0(.dout(w_dff_A_nZcpkXBO8_0),.din(w_dff_A_B5AJLaOR1_0),.clk(gclk));
	jdff dff_A_nZcpkXBO8_0(.dout(w_dff_A_5U2Bz5y88_0),.din(w_dff_A_nZcpkXBO8_0),.clk(gclk));
	jdff dff_A_5U2Bz5y88_0(.dout(w_dff_A_uEbCVBHr1_0),.din(w_dff_A_5U2Bz5y88_0),.clk(gclk));
	jdff dff_A_uEbCVBHr1_0(.dout(w_dff_A_oQb8kAjb1_0),.din(w_dff_A_uEbCVBHr1_0),.clk(gclk));
	jdff dff_A_oQb8kAjb1_0(.dout(w_dff_A_IywEnK069_0),.din(w_dff_A_oQb8kAjb1_0),.clk(gclk));
	jdff dff_A_IywEnK069_0(.dout(w_dff_A_vEQNVOj77_0),.din(w_dff_A_IywEnK069_0),.clk(gclk));
	jdff dff_A_vEQNVOj77_0(.dout(w_dff_A_pRi1a1yi5_0),.din(w_dff_A_vEQNVOj77_0),.clk(gclk));
	jdff dff_A_pRi1a1yi5_0(.dout(w_dff_A_27Rgy5BW4_0),.din(w_dff_A_pRi1a1yi5_0),.clk(gclk));
	jdff dff_A_27Rgy5BW4_0(.dout(G528),.din(w_dff_A_27Rgy5BW4_0),.clk(gclk));
	jdff dff_A_7DWNk9T28_1(.dout(w_dff_A_GPbwSp8Y7_0),.din(w_dff_A_7DWNk9T28_1),.clk(gclk));
	jdff dff_A_GPbwSp8Y7_0(.dout(w_dff_A_MS3QaBnO0_0),.din(w_dff_A_GPbwSp8Y7_0),.clk(gclk));
	jdff dff_A_MS3QaBnO0_0(.dout(w_dff_A_RCPFmIum0_0),.din(w_dff_A_MS3QaBnO0_0),.clk(gclk));
	jdff dff_A_RCPFmIum0_0(.dout(w_dff_A_neqVBslu4_0),.din(w_dff_A_RCPFmIum0_0),.clk(gclk));
	jdff dff_A_neqVBslu4_0(.dout(w_dff_A_KmsC0oP25_0),.din(w_dff_A_neqVBslu4_0),.clk(gclk));
	jdff dff_A_KmsC0oP25_0(.dout(w_dff_A_MILeSvMh8_0),.din(w_dff_A_KmsC0oP25_0),.clk(gclk));
	jdff dff_A_MILeSvMh8_0(.dout(w_dff_A_KOgqUn8M5_0),.din(w_dff_A_MILeSvMh8_0),.clk(gclk));
	jdff dff_A_KOgqUn8M5_0(.dout(w_dff_A_h9b3Mp9F5_0),.din(w_dff_A_KOgqUn8M5_0),.clk(gclk));
	jdff dff_A_h9b3Mp9F5_0(.dout(w_dff_A_eDz3EFhw6_0),.din(w_dff_A_h9b3Mp9F5_0),.clk(gclk));
	jdff dff_A_eDz3EFhw6_0(.dout(w_dff_A_quOz00uA6_0),.din(w_dff_A_eDz3EFhw6_0),.clk(gclk));
	jdff dff_A_quOz00uA6_0(.dout(w_dff_A_nBPxCYg98_0),.din(w_dff_A_quOz00uA6_0),.clk(gclk));
	jdff dff_A_nBPxCYg98_0(.dout(w_dff_A_3t2382n48_0),.din(w_dff_A_nBPxCYg98_0),.clk(gclk));
	jdff dff_A_3t2382n48_0(.dout(w_dff_A_QvNZENNn7_0),.din(w_dff_A_3t2382n48_0),.clk(gclk));
	jdff dff_A_QvNZENNn7_0(.dout(w_dff_A_2AnsEprB6_0),.din(w_dff_A_QvNZENNn7_0),.clk(gclk));
	jdff dff_A_2AnsEprB6_0(.dout(w_dff_A_ZHgUQeHx9_0),.din(w_dff_A_2AnsEprB6_0),.clk(gclk));
	jdff dff_A_ZHgUQeHx9_0(.dout(w_dff_A_nRGZjNJJ2_0),.din(w_dff_A_ZHgUQeHx9_0),.clk(gclk));
	jdff dff_A_nRGZjNJJ2_0(.dout(w_dff_A_oOCp26wR0_0),.din(w_dff_A_nRGZjNJJ2_0),.clk(gclk));
	jdff dff_A_oOCp26wR0_0(.dout(w_dff_A_jAfaHDjI4_0),.din(w_dff_A_oOCp26wR0_0),.clk(gclk));
	jdff dff_A_jAfaHDjI4_0(.dout(w_dff_A_92NsBwqc2_0),.din(w_dff_A_jAfaHDjI4_0),.clk(gclk));
	jdff dff_A_92NsBwqc2_0(.dout(w_dff_A_D6IxUAoF9_0),.din(w_dff_A_92NsBwqc2_0),.clk(gclk));
	jdff dff_A_D6IxUAoF9_0(.dout(w_dff_A_VBz9XKmS4_0),.din(w_dff_A_D6IxUAoF9_0),.clk(gclk));
	jdff dff_A_VBz9XKmS4_0(.dout(w_dff_A_1YgUQNqL8_0),.din(w_dff_A_VBz9XKmS4_0),.clk(gclk));
	jdff dff_A_1YgUQNqL8_0(.dout(w_dff_A_S6Jrppwh8_0),.din(w_dff_A_1YgUQNqL8_0),.clk(gclk));
	jdff dff_A_S6Jrppwh8_0(.dout(w_dff_A_qHubb2Kl7_0),.din(w_dff_A_S6Jrppwh8_0),.clk(gclk));
	jdff dff_A_qHubb2Kl7_0(.dout(w_dff_A_5yPzmDu28_0),.din(w_dff_A_qHubb2Kl7_0),.clk(gclk));
	jdff dff_A_5yPzmDu28_0(.dout(w_dff_A_po4c7hv07_0),.din(w_dff_A_5yPzmDu28_0),.clk(gclk));
	jdff dff_A_po4c7hv07_0(.dout(w_dff_A_zpz9j1RA2_0),.din(w_dff_A_po4c7hv07_0),.clk(gclk));
	jdff dff_A_zpz9j1RA2_0(.dout(w_dff_A_jumjBDQd2_0),.din(w_dff_A_zpz9j1RA2_0),.clk(gclk));
	jdff dff_A_jumjBDQd2_0(.dout(w_dff_A_L8x3EYEC8_0),.din(w_dff_A_jumjBDQd2_0),.clk(gclk));
	jdff dff_A_L8x3EYEC8_0(.dout(w_dff_A_XFamfHR42_0),.din(w_dff_A_L8x3EYEC8_0),.clk(gclk));
	jdff dff_A_XFamfHR42_0(.dout(w_dff_A_gLD2oU346_0),.din(w_dff_A_XFamfHR42_0),.clk(gclk));
	jdff dff_A_gLD2oU346_0(.dout(w_dff_A_R8nDrZIW9_0),.din(w_dff_A_gLD2oU346_0),.clk(gclk));
	jdff dff_A_R8nDrZIW9_0(.dout(w_dff_A_020cK1fd5_0),.din(w_dff_A_R8nDrZIW9_0),.clk(gclk));
	jdff dff_A_020cK1fd5_0(.dout(w_dff_A_qRr5YlwW2_0),.din(w_dff_A_020cK1fd5_0),.clk(gclk));
	jdff dff_A_qRr5YlwW2_0(.dout(w_dff_A_yHEuMzV22_0),.din(w_dff_A_qRr5YlwW2_0),.clk(gclk));
	jdff dff_A_yHEuMzV22_0(.dout(w_dff_A_miszG4F57_0),.din(w_dff_A_yHEuMzV22_0),.clk(gclk));
	jdff dff_A_miszG4F57_0(.dout(w_dff_A_iZWM93os3_0),.din(w_dff_A_miszG4F57_0),.clk(gclk));
	jdff dff_A_iZWM93os3_0(.dout(w_dff_A_lXXplaG52_0),.din(w_dff_A_iZWM93os3_0),.clk(gclk));
	jdff dff_A_lXXplaG52_0(.dout(G526),.din(w_dff_A_lXXplaG52_0),.clk(gclk));
	jdff dff_A_KWb9btUV8_1(.dout(w_dff_A_7wQgQEAD2_0),.din(w_dff_A_KWb9btUV8_1),.clk(gclk));
	jdff dff_A_7wQgQEAD2_0(.dout(w_dff_A_1QoJXjGR3_0),.din(w_dff_A_7wQgQEAD2_0),.clk(gclk));
	jdff dff_A_1QoJXjGR3_0(.dout(w_dff_A_QFdvQS6w0_0),.din(w_dff_A_1QoJXjGR3_0),.clk(gclk));
	jdff dff_A_QFdvQS6w0_0(.dout(w_dff_A_A9KPtago5_0),.din(w_dff_A_QFdvQS6w0_0),.clk(gclk));
	jdff dff_A_A9KPtago5_0(.dout(w_dff_A_WdZgDvQ91_0),.din(w_dff_A_A9KPtago5_0),.clk(gclk));
	jdff dff_A_WdZgDvQ91_0(.dout(w_dff_A_Ok5dBrgs0_0),.din(w_dff_A_WdZgDvQ91_0),.clk(gclk));
	jdff dff_A_Ok5dBrgs0_0(.dout(w_dff_A_f2s49wTY3_0),.din(w_dff_A_Ok5dBrgs0_0),.clk(gclk));
	jdff dff_A_f2s49wTY3_0(.dout(w_dff_A_pOfHl5DV2_0),.din(w_dff_A_f2s49wTY3_0),.clk(gclk));
	jdff dff_A_pOfHl5DV2_0(.dout(w_dff_A_T4dIaOIi1_0),.din(w_dff_A_pOfHl5DV2_0),.clk(gclk));
	jdff dff_A_T4dIaOIi1_0(.dout(w_dff_A_FTgag51p5_0),.din(w_dff_A_T4dIaOIi1_0),.clk(gclk));
	jdff dff_A_FTgag51p5_0(.dout(w_dff_A_czAU8MEn8_0),.din(w_dff_A_FTgag51p5_0),.clk(gclk));
	jdff dff_A_czAU8MEn8_0(.dout(w_dff_A_I7yfueF96_0),.din(w_dff_A_czAU8MEn8_0),.clk(gclk));
	jdff dff_A_I7yfueF96_0(.dout(w_dff_A_fdwEG1Nz3_0),.din(w_dff_A_I7yfueF96_0),.clk(gclk));
	jdff dff_A_fdwEG1Nz3_0(.dout(w_dff_A_ZniZFP1Y8_0),.din(w_dff_A_fdwEG1Nz3_0),.clk(gclk));
	jdff dff_A_ZniZFP1Y8_0(.dout(w_dff_A_23MY2xiG1_0),.din(w_dff_A_ZniZFP1Y8_0),.clk(gclk));
	jdff dff_A_23MY2xiG1_0(.dout(w_dff_A_UpeCYdxG6_0),.din(w_dff_A_23MY2xiG1_0),.clk(gclk));
	jdff dff_A_UpeCYdxG6_0(.dout(w_dff_A_WyfAiTCP8_0),.din(w_dff_A_UpeCYdxG6_0),.clk(gclk));
	jdff dff_A_WyfAiTCP8_0(.dout(w_dff_A_ElcTUQB91_0),.din(w_dff_A_WyfAiTCP8_0),.clk(gclk));
	jdff dff_A_ElcTUQB91_0(.dout(w_dff_A_EDpJjPvG1_0),.din(w_dff_A_ElcTUQB91_0),.clk(gclk));
	jdff dff_A_EDpJjPvG1_0(.dout(w_dff_A_AkCpCpk23_0),.din(w_dff_A_EDpJjPvG1_0),.clk(gclk));
	jdff dff_A_AkCpCpk23_0(.dout(w_dff_A_sImYZN0Z7_0),.din(w_dff_A_AkCpCpk23_0),.clk(gclk));
	jdff dff_A_sImYZN0Z7_0(.dout(w_dff_A_Dcmsywqt3_0),.din(w_dff_A_sImYZN0Z7_0),.clk(gclk));
	jdff dff_A_Dcmsywqt3_0(.dout(w_dff_A_G17aN4Ui6_0),.din(w_dff_A_Dcmsywqt3_0),.clk(gclk));
	jdff dff_A_G17aN4Ui6_0(.dout(w_dff_A_ihS8N92j6_0),.din(w_dff_A_G17aN4Ui6_0),.clk(gclk));
	jdff dff_A_ihS8N92j6_0(.dout(w_dff_A_chl4Yehu0_0),.din(w_dff_A_ihS8N92j6_0),.clk(gclk));
	jdff dff_A_chl4Yehu0_0(.dout(w_dff_A_g5guW00w0_0),.din(w_dff_A_chl4Yehu0_0),.clk(gclk));
	jdff dff_A_g5guW00w0_0(.dout(w_dff_A_PCZMgcec4_0),.din(w_dff_A_g5guW00w0_0),.clk(gclk));
	jdff dff_A_PCZMgcec4_0(.dout(w_dff_A_CyN3oALh9_0),.din(w_dff_A_PCZMgcec4_0),.clk(gclk));
	jdff dff_A_CyN3oALh9_0(.dout(w_dff_A_NuqozF7E7_0),.din(w_dff_A_CyN3oALh9_0),.clk(gclk));
	jdff dff_A_NuqozF7E7_0(.dout(w_dff_A_1IEEYlq61_0),.din(w_dff_A_NuqozF7E7_0),.clk(gclk));
	jdff dff_A_1IEEYlq61_0(.dout(w_dff_A_jGiIuj499_0),.din(w_dff_A_1IEEYlq61_0),.clk(gclk));
	jdff dff_A_jGiIuj499_0(.dout(w_dff_A_bGbD4Y8e4_0),.din(w_dff_A_jGiIuj499_0),.clk(gclk));
	jdff dff_A_bGbD4Y8e4_0(.dout(w_dff_A_pREiaToH1_0),.din(w_dff_A_bGbD4Y8e4_0),.clk(gclk));
	jdff dff_A_pREiaToH1_0(.dout(w_dff_A_9fqtvgvi1_0),.din(w_dff_A_pREiaToH1_0),.clk(gclk));
	jdff dff_A_9fqtvgvi1_0(.dout(w_dff_A_k6cdTKzc3_0),.din(w_dff_A_9fqtvgvi1_0),.clk(gclk));
	jdff dff_A_k6cdTKzc3_0(.dout(w_dff_A_4MMsdCtT3_0),.din(w_dff_A_k6cdTKzc3_0),.clk(gclk));
	jdff dff_A_4MMsdCtT3_0(.dout(w_dff_A_kDXVf9032_0),.din(w_dff_A_4MMsdCtT3_0),.clk(gclk));
	jdff dff_A_kDXVf9032_0(.dout(w_dff_A_oCouwUys8_0),.din(w_dff_A_kDXVf9032_0),.clk(gclk));
	jdff dff_A_oCouwUys8_0(.dout(G524),.din(w_dff_A_oCouwUys8_0),.clk(gclk));
	jdff dff_A_Ecw3XE0C8_1(.dout(w_dff_A_JxtG2gM51_0),.din(w_dff_A_Ecw3XE0C8_1),.clk(gclk));
	jdff dff_A_JxtG2gM51_0(.dout(w_dff_A_w9givJGQ5_0),.din(w_dff_A_JxtG2gM51_0),.clk(gclk));
	jdff dff_A_w9givJGQ5_0(.dout(w_dff_A_BX5t45CH8_0),.din(w_dff_A_w9givJGQ5_0),.clk(gclk));
	jdff dff_A_BX5t45CH8_0(.dout(w_dff_A_eAeQP5g77_0),.din(w_dff_A_BX5t45CH8_0),.clk(gclk));
	jdff dff_A_eAeQP5g77_0(.dout(w_dff_A_dkTfI9qz8_0),.din(w_dff_A_eAeQP5g77_0),.clk(gclk));
	jdff dff_A_dkTfI9qz8_0(.dout(w_dff_A_y4j5juJP0_0),.din(w_dff_A_dkTfI9qz8_0),.clk(gclk));
	jdff dff_A_y4j5juJP0_0(.dout(w_dff_A_6D3O5RuW5_0),.din(w_dff_A_y4j5juJP0_0),.clk(gclk));
	jdff dff_A_6D3O5RuW5_0(.dout(w_dff_A_8zl4laL25_0),.din(w_dff_A_6D3O5RuW5_0),.clk(gclk));
	jdff dff_A_8zl4laL25_0(.dout(w_dff_A_F9zbjyzh8_0),.din(w_dff_A_8zl4laL25_0),.clk(gclk));
	jdff dff_A_F9zbjyzh8_0(.dout(w_dff_A_fRURxQSj2_0),.din(w_dff_A_F9zbjyzh8_0),.clk(gclk));
	jdff dff_A_fRURxQSj2_0(.dout(w_dff_A_ZcNOHpNk4_0),.din(w_dff_A_fRURxQSj2_0),.clk(gclk));
	jdff dff_A_ZcNOHpNk4_0(.dout(w_dff_A_Pyr9ZYRo9_0),.din(w_dff_A_ZcNOHpNk4_0),.clk(gclk));
	jdff dff_A_Pyr9ZYRo9_0(.dout(w_dff_A_hvojzIHa4_0),.din(w_dff_A_Pyr9ZYRo9_0),.clk(gclk));
	jdff dff_A_hvojzIHa4_0(.dout(w_dff_A_E8yhJQnZ7_0),.din(w_dff_A_hvojzIHa4_0),.clk(gclk));
	jdff dff_A_E8yhJQnZ7_0(.dout(w_dff_A_8GVBXo291_0),.din(w_dff_A_E8yhJQnZ7_0),.clk(gclk));
	jdff dff_A_8GVBXo291_0(.dout(w_dff_A_9lKYjnjk7_0),.din(w_dff_A_8GVBXo291_0),.clk(gclk));
	jdff dff_A_9lKYjnjk7_0(.dout(w_dff_A_cmNluERk6_0),.din(w_dff_A_9lKYjnjk7_0),.clk(gclk));
	jdff dff_A_cmNluERk6_0(.dout(w_dff_A_CZQDbA8H0_0),.din(w_dff_A_cmNluERk6_0),.clk(gclk));
	jdff dff_A_CZQDbA8H0_0(.dout(w_dff_A_wQK9nt550_0),.din(w_dff_A_CZQDbA8H0_0),.clk(gclk));
	jdff dff_A_wQK9nt550_0(.dout(w_dff_A_G9kc5lVR6_0),.din(w_dff_A_wQK9nt550_0),.clk(gclk));
	jdff dff_A_G9kc5lVR6_0(.dout(w_dff_A_Augx0A7H8_0),.din(w_dff_A_G9kc5lVR6_0),.clk(gclk));
	jdff dff_A_Augx0A7H8_0(.dout(w_dff_A_MsGYMzO90_0),.din(w_dff_A_Augx0A7H8_0),.clk(gclk));
	jdff dff_A_MsGYMzO90_0(.dout(w_dff_A_rzFpPzJV4_0),.din(w_dff_A_MsGYMzO90_0),.clk(gclk));
	jdff dff_A_rzFpPzJV4_0(.dout(w_dff_A_E9msK8wW2_0),.din(w_dff_A_rzFpPzJV4_0),.clk(gclk));
	jdff dff_A_E9msK8wW2_0(.dout(w_dff_A_r2Lmlu2r1_0),.din(w_dff_A_E9msK8wW2_0),.clk(gclk));
	jdff dff_A_r2Lmlu2r1_0(.dout(w_dff_A_V6c6oLjl9_0),.din(w_dff_A_r2Lmlu2r1_0),.clk(gclk));
	jdff dff_A_V6c6oLjl9_0(.dout(w_dff_A_pCm67LpO3_0),.din(w_dff_A_V6c6oLjl9_0),.clk(gclk));
	jdff dff_A_pCm67LpO3_0(.dout(w_dff_A_wznbd0EH2_0),.din(w_dff_A_pCm67LpO3_0),.clk(gclk));
	jdff dff_A_wznbd0EH2_0(.dout(w_dff_A_9z0AByg69_0),.din(w_dff_A_wznbd0EH2_0),.clk(gclk));
	jdff dff_A_9z0AByg69_0(.dout(w_dff_A_gEiuKOGj2_0),.din(w_dff_A_9z0AByg69_0),.clk(gclk));
	jdff dff_A_gEiuKOGj2_0(.dout(w_dff_A_xArsL7LR1_0),.din(w_dff_A_gEiuKOGj2_0),.clk(gclk));
	jdff dff_A_xArsL7LR1_0(.dout(w_dff_A_p6iOJAju7_0),.din(w_dff_A_xArsL7LR1_0),.clk(gclk));
	jdff dff_A_p6iOJAju7_0(.dout(w_dff_A_tadBGjSV2_0),.din(w_dff_A_p6iOJAju7_0),.clk(gclk));
	jdff dff_A_tadBGjSV2_0(.dout(w_dff_A_A14g1eR75_0),.din(w_dff_A_tadBGjSV2_0),.clk(gclk));
	jdff dff_A_A14g1eR75_0(.dout(w_dff_A_3BrMdQ0f5_0),.din(w_dff_A_A14g1eR75_0),.clk(gclk));
	jdff dff_A_3BrMdQ0f5_0(.dout(w_dff_A_XzfZhxu66_0),.din(w_dff_A_3BrMdQ0f5_0),.clk(gclk));
	jdff dff_A_XzfZhxu66_0(.dout(w_dff_A_uxlMMV2T6_0),.din(w_dff_A_XzfZhxu66_0),.clk(gclk));
	jdff dff_A_uxlMMV2T6_0(.dout(G279),.din(w_dff_A_uxlMMV2T6_0),.clk(gclk));
	jdff dff_A_mkapjFNr2_1(.dout(w_dff_A_gseXjABl7_0),.din(w_dff_A_mkapjFNr2_1),.clk(gclk));
	jdff dff_A_gseXjABl7_0(.dout(w_dff_A_VSopTJoF1_0),.din(w_dff_A_gseXjABl7_0),.clk(gclk));
	jdff dff_A_VSopTJoF1_0(.dout(w_dff_A_M1BkhQtZ6_0),.din(w_dff_A_VSopTJoF1_0),.clk(gclk));
	jdff dff_A_M1BkhQtZ6_0(.dout(w_dff_A_5PH3PAnc6_0),.din(w_dff_A_M1BkhQtZ6_0),.clk(gclk));
	jdff dff_A_5PH3PAnc6_0(.dout(w_dff_A_5St6i9pA1_0),.din(w_dff_A_5PH3PAnc6_0),.clk(gclk));
	jdff dff_A_5St6i9pA1_0(.dout(w_dff_A_DaujxEGc1_0),.din(w_dff_A_5St6i9pA1_0),.clk(gclk));
	jdff dff_A_DaujxEGc1_0(.dout(w_dff_A_OeMst2Un4_0),.din(w_dff_A_DaujxEGc1_0),.clk(gclk));
	jdff dff_A_OeMst2Un4_0(.dout(w_dff_A_HAbOU5VZ0_0),.din(w_dff_A_OeMst2Un4_0),.clk(gclk));
	jdff dff_A_HAbOU5VZ0_0(.dout(w_dff_A_zZBKXntg1_0),.din(w_dff_A_HAbOU5VZ0_0),.clk(gclk));
	jdff dff_A_zZBKXntg1_0(.dout(w_dff_A_u9PKfo3T1_0),.din(w_dff_A_zZBKXntg1_0),.clk(gclk));
	jdff dff_A_u9PKfo3T1_0(.dout(w_dff_A_p9LCjROE3_0),.din(w_dff_A_u9PKfo3T1_0),.clk(gclk));
	jdff dff_A_p9LCjROE3_0(.dout(w_dff_A_9c6bRCCB5_0),.din(w_dff_A_p9LCjROE3_0),.clk(gclk));
	jdff dff_A_9c6bRCCB5_0(.dout(w_dff_A_62APR6QZ6_0),.din(w_dff_A_9c6bRCCB5_0),.clk(gclk));
	jdff dff_A_62APR6QZ6_0(.dout(w_dff_A_MGYQNllt8_0),.din(w_dff_A_62APR6QZ6_0),.clk(gclk));
	jdff dff_A_MGYQNllt8_0(.dout(w_dff_A_QL6RY0b14_0),.din(w_dff_A_MGYQNllt8_0),.clk(gclk));
	jdff dff_A_QL6RY0b14_0(.dout(w_dff_A_mMvxT7Yz4_0),.din(w_dff_A_QL6RY0b14_0),.clk(gclk));
	jdff dff_A_mMvxT7Yz4_0(.dout(w_dff_A_CwAxFP3j3_0),.din(w_dff_A_mMvxT7Yz4_0),.clk(gclk));
	jdff dff_A_CwAxFP3j3_0(.dout(w_dff_A_jmiroCuE7_0),.din(w_dff_A_CwAxFP3j3_0),.clk(gclk));
	jdff dff_A_jmiroCuE7_0(.dout(w_dff_A_eEITPnr53_0),.din(w_dff_A_jmiroCuE7_0),.clk(gclk));
	jdff dff_A_eEITPnr53_0(.dout(w_dff_A_DVJWp4ud6_0),.din(w_dff_A_eEITPnr53_0),.clk(gclk));
	jdff dff_A_DVJWp4ud6_0(.dout(w_dff_A_XpqYFIWo5_0),.din(w_dff_A_DVJWp4ud6_0),.clk(gclk));
	jdff dff_A_XpqYFIWo5_0(.dout(w_dff_A_g3P4FDHU6_0),.din(w_dff_A_XpqYFIWo5_0),.clk(gclk));
	jdff dff_A_g3P4FDHU6_0(.dout(w_dff_A_Zl2UCqnZ8_0),.din(w_dff_A_g3P4FDHU6_0),.clk(gclk));
	jdff dff_A_Zl2UCqnZ8_0(.dout(w_dff_A_ExnCMEin5_0),.din(w_dff_A_Zl2UCqnZ8_0),.clk(gclk));
	jdff dff_A_ExnCMEin5_0(.dout(w_dff_A_MbZyLN2u2_0),.din(w_dff_A_ExnCMEin5_0),.clk(gclk));
	jdff dff_A_MbZyLN2u2_0(.dout(w_dff_A_OZJ01zsz1_0),.din(w_dff_A_MbZyLN2u2_0),.clk(gclk));
	jdff dff_A_OZJ01zsz1_0(.dout(w_dff_A_MQ7WdUvN5_0),.din(w_dff_A_OZJ01zsz1_0),.clk(gclk));
	jdff dff_A_MQ7WdUvN5_0(.dout(w_dff_A_yAiHocCZ2_0),.din(w_dff_A_MQ7WdUvN5_0),.clk(gclk));
	jdff dff_A_yAiHocCZ2_0(.dout(w_dff_A_JCq70if10_0),.din(w_dff_A_yAiHocCZ2_0),.clk(gclk));
	jdff dff_A_JCq70if10_0(.dout(w_dff_A_wLat4gce2_0),.din(w_dff_A_JCq70if10_0),.clk(gclk));
	jdff dff_A_wLat4gce2_0(.dout(w_dff_A_Dsfqz4gA9_0),.din(w_dff_A_wLat4gce2_0),.clk(gclk));
	jdff dff_A_Dsfqz4gA9_0(.dout(w_dff_A_0JEkb5Ut9_0),.din(w_dff_A_Dsfqz4gA9_0),.clk(gclk));
	jdff dff_A_0JEkb5Ut9_0(.dout(w_dff_A_COggvmzL5_0),.din(w_dff_A_0JEkb5Ut9_0),.clk(gclk));
	jdff dff_A_COggvmzL5_0(.dout(w_dff_A_Ap4Dv5kD4_0),.din(w_dff_A_COggvmzL5_0),.clk(gclk));
	jdff dff_A_Ap4Dv5kD4_0(.dout(w_dff_A_RBEDV1Rf6_0),.din(w_dff_A_Ap4Dv5kD4_0),.clk(gclk));
	jdff dff_A_RBEDV1Rf6_0(.dout(w_dff_A_KQ4WqkKx5_0),.din(w_dff_A_RBEDV1Rf6_0),.clk(gclk));
	jdff dff_A_KQ4WqkKx5_0(.dout(w_dff_A_F62O6jpF7_0),.din(w_dff_A_KQ4WqkKx5_0),.clk(gclk));
	jdff dff_A_F62O6jpF7_0(.dout(w_dff_A_SAgjieT26_0),.din(w_dff_A_F62O6jpF7_0),.clk(gclk));
	jdff dff_A_SAgjieT26_0(.dout(G436),.din(w_dff_A_SAgjieT26_0),.clk(gclk));
	jdff dff_A_JNSQA5WW0_1(.dout(w_dff_A_sZ2Ye7S04_0),.din(w_dff_A_JNSQA5WW0_1),.clk(gclk));
	jdff dff_A_sZ2Ye7S04_0(.dout(w_dff_A_p9J2VSBu8_0),.din(w_dff_A_sZ2Ye7S04_0),.clk(gclk));
	jdff dff_A_p9J2VSBu8_0(.dout(w_dff_A_fCUDzCgx7_0),.din(w_dff_A_p9J2VSBu8_0),.clk(gclk));
	jdff dff_A_fCUDzCgx7_0(.dout(w_dff_A_UxmXelcD8_0),.din(w_dff_A_fCUDzCgx7_0),.clk(gclk));
	jdff dff_A_UxmXelcD8_0(.dout(w_dff_A_dd5dwjNi9_0),.din(w_dff_A_UxmXelcD8_0),.clk(gclk));
	jdff dff_A_dd5dwjNi9_0(.dout(w_dff_A_IJyDPoxj6_0),.din(w_dff_A_dd5dwjNi9_0),.clk(gclk));
	jdff dff_A_IJyDPoxj6_0(.dout(w_dff_A_Ukr7kAib5_0),.din(w_dff_A_IJyDPoxj6_0),.clk(gclk));
	jdff dff_A_Ukr7kAib5_0(.dout(w_dff_A_t0MR3e8e7_0),.din(w_dff_A_Ukr7kAib5_0),.clk(gclk));
	jdff dff_A_t0MR3e8e7_0(.dout(w_dff_A_mZb1Kx5i2_0),.din(w_dff_A_t0MR3e8e7_0),.clk(gclk));
	jdff dff_A_mZb1Kx5i2_0(.dout(w_dff_A_sbK9BLBZ5_0),.din(w_dff_A_mZb1Kx5i2_0),.clk(gclk));
	jdff dff_A_sbK9BLBZ5_0(.dout(w_dff_A_I68zm5vB6_0),.din(w_dff_A_sbK9BLBZ5_0),.clk(gclk));
	jdff dff_A_I68zm5vB6_0(.dout(w_dff_A_Zso0yqaY5_0),.din(w_dff_A_I68zm5vB6_0),.clk(gclk));
	jdff dff_A_Zso0yqaY5_0(.dout(w_dff_A_CSt4kDh24_0),.din(w_dff_A_Zso0yqaY5_0),.clk(gclk));
	jdff dff_A_CSt4kDh24_0(.dout(w_dff_A_uC9RWX2K2_0),.din(w_dff_A_CSt4kDh24_0),.clk(gclk));
	jdff dff_A_uC9RWX2K2_0(.dout(w_dff_A_Pc6eUPN04_0),.din(w_dff_A_uC9RWX2K2_0),.clk(gclk));
	jdff dff_A_Pc6eUPN04_0(.dout(w_dff_A_tUeVAjnK3_0),.din(w_dff_A_Pc6eUPN04_0),.clk(gclk));
	jdff dff_A_tUeVAjnK3_0(.dout(w_dff_A_1MuqX2YZ2_0),.din(w_dff_A_tUeVAjnK3_0),.clk(gclk));
	jdff dff_A_1MuqX2YZ2_0(.dout(w_dff_A_twvCwRQT9_0),.din(w_dff_A_1MuqX2YZ2_0),.clk(gclk));
	jdff dff_A_twvCwRQT9_0(.dout(w_dff_A_7x8xuhKI4_0),.din(w_dff_A_twvCwRQT9_0),.clk(gclk));
	jdff dff_A_7x8xuhKI4_0(.dout(w_dff_A_ewI8G7jQ8_0),.din(w_dff_A_7x8xuhKI4_0),.clk(gclk));
	jdff dff_A_ewI8G7jQ8_0(.dout(w_dff_A_ktRMidhS3_0),.din(w_dff_A_ewI8G7jQ8_0),.clk(gclk));
	jdff dff_A_ktRMidhS3_0(.dout(w_dff_A_rERIW63D6_0),.din(w_dff_A_ktRMidhS3_0),.clk(gclk));
	jdff dff_A_rERIW63D6_0(.dout(w_dff_A_Y6T4ICtY3_0),.din(w_dff_A_rERIW63D6_0),.clk(gclk));
	jdff dff_A_Y6T4ICtY3_0(.dout(w_dff_A_1TIdyplS2_0),.din(w_dff_A_Y6T4ICtY3_0),.clk(gclk));
	jdff dff_A_1TIdyplS2_0(.dout(w_dff_A_4rFqcHvh3_0),.din(w_dff_A_1TIdyplS2_0),.clk(gclk));
	jdff dff_A_4rFqcHvh3_0(.dout(w_dff_A_0f0qnMpj7_0),.din(w_dff_A_4rFqcHvh3_0),.clk(gclk));
	jdff dff_A_0f0qnMpj7_0(.dout(w_dff_A_79ZePbnR8_0),.din(w_dff_A_0f0qnMpj7_0),.clk(gclk));
	jdff dff_A_79ZePbnR8_0(.dout(w_dff_A_g5sNgMBQ3_0),.din(w_dff_A_79ZePbnR8_0),.clk(gclk));
	jdff dff_A_g5sNgMBQ3_0(.dout(w_dff_A_6jAGtIOk9_0),.din(w_dff_A_g5sNgMBQ3_0),.clk(gclk));
	jdff dff_A_6jAGtIOk9_0(.dout(w_dff_A_vSpJVBrE1_0),.din(w_dff_A_6jAGtIOk9_0),.clk(gclk));
	jdff dff_A_vSpJVBrE1_0(.dout(w_dff_A_mYbgiXqX8_0),.din(w_dff_A_vSpJVBrE1_0),.clk(gclk));
	jdff dff_A_mYbgiXqX8_0(.dout(w_dff_A_bEvidwvA1_0),.din(w_dff_A_mYbgiXqX8_0),.clk(gclk));
	jdff dff_A_bEvidwvA1_0(.dout(w_dff_A_46ntLdMS0_0),.din(w_dff_A_bEvidwvA1_0),.clk(gclk));
	jdff dff_A_46ntLdMS0_0(.dout(w_dff_A_V98IpRcV3_0),.din(w_dff_A_46ntLdMS0_0),.clk(gclk));
	jdff dff_A_V98IpRcV3_0(.dout(w_dff_A_a57WLguh3_0),.din(w_dff_A_V98IpRcV3_0),.clk(gclk));
	jdff dff_A_a57WLguh3_0(.dout(w_dff_A_qWkNnZEb1_0),.din(w_dff_A_a57WLguh3_0),.clk(gclk));
	jdff dff_A_qWkNnZEb1_0(.dout(w_dff_A_zzpcdWs51_0),.din(w_dff_A_qWkNnZEb1_0),.clk(gclk));
	jdff dff_A_zzpcdWs51_0(.dout(w_dff_A_bK1yUz2T7_0),.din(w_dff_A_zzpcdWs51_0),.clk(gclk));
	jdff dff_A_bK1yUz2T7_0(.dout(G478),.din(w_dff_A_bK1yUz2T7_0),.clk(gclk));
	jdff dff_A_UcGMKMoa0_1(.dout(w_dff_A_Jx3pVlHg4_0),.din(w_dff_A_UcGMKMoa0_1),.clk(gclk));
	jdff dff_A_Jx3pVlHg4_0(.dout(w_dff_A_EoD5PMn01_0),.din(w_dff_A_Jx3pVlHg4_0),.clk(gclk));
	jdff dff_A_EoD5PMn01_0(.dout(w_dff_A_zJgKbrJK3_0),.din(w_dff_A_EoD5PMn01_0),.clk(gclk));
	jdff dff_A_zJgKbrJK3_0(.dout(w_dff_A_SXVwpqOM7_0),.din(w_dff_A_zJgKbrJK3_0),.clk(gclk));
	jdff dff_A_SXVwpqOM7_0(.dout(w_dff_A_0AU0VOUP1_0),.din(w_dff_A_SXVwpqOM7_0),.clk(gclk));
	jdff dff_A_0AU0VOUP1_0(.dout(w_dff_A_5jMvbd6v9_0),.din(w_dff_A_0AU0VOUP1_0),.clk(gclk));
	jdff dff_A_5jMvbd6v9_0(.dout(w_dff_A_oJQSa3TH1_0),.din(w_dff_A_5jMvbd6v9_0),.clk(gclk));
	jdff dff_A_oJQSa3TH1_0(.dout(w_dff_A_JEC6AGJ29_0),.din(w_dff_A_oJQSa3TH1_0),.clk(gclk));
	jdff dff_A_JEC6AGJ29_0(.dout(w_dff_A_4risWdAi4_0),.din(w_dff_A_JEC6AGJ29_0),.clk(gclk));
	jdff dff_A_4risWdAi4_0(.dout(w_dff_A_p7yvjMcI6_0),.din(w_dff_A_4risWdAi4_0),.clk(gclk));
	jdff dff_A_p7yvjMcI6_0(.dout(w_dff_A_QxRaRArh5_0),.din(w_dff_A_p7yvjMcI6_0),.clk(gclk));
	jdff dff_A_QxRaRArh5_0(.dout(w_dff_A_1MaeLNCf7_0),.din(w_dff_A_QxRaRArh5_0),.clk(gclk));
	jdff dff_A_1MaeLNCf7_0(.dout(w_dff_A_hJV1y4ok9_0),.din(w_dff_A_1MaeLNCf7_0),.clk(gclk));
	jdff dff_A_hJV1y4ok9_0(.dout(w_dff_A_Bpyenhtu7_0),.din(w_dff_A_hJV1y4ok9_0),.clk(gclk));
	jdff dff_A_Bpyenhtu7_0(.dout(w_dff_A_bMwFIHxA3_0),.din(w_dff_A_Bpyenhtu7_0),.clk(gclk));
	jdff dff_A_bMwFIHxA3_0(.dout(w_dff_A_7L91PiaT8_0),.din(w_dff_A_bMwFIHxA3_0),.clk(gclk));
	jdff dff_A_7L91PiaT8_0(.dout(w_dff_A_ZHMStFjQ9_0),.din(w_dff_A_7L91PiaT8_0),.clk(gclk));
	jdff dff_A_ZHMStFjQ9_0(.dout(w_dff_A_HiyQfKje3_0),.din(w_dff_A_ZHMStFjQ9_0),.clk(gclk));
	jdff dff_A_HiyQfKje3_0(.dout(w_dff_A_t08A0Wh90_0),.din(w_dff_A_HiyQfKje3_0),.clk(gclk));
	jdff dff_A_t08A0Wh90_0(.dout(w_dff_A_yYxBmyyI7_0),.din(w_dff_A_t08A0Wh90_0),.clk(gclk));
	jdff dff_A_yYxBmyyI7_0(.dout(w_dff_A_uHsWKiTq6_0),.din(w_dff_A_yYxBmyyI7_0),.clk(gclk));
	jdff dff_A_uHsWKiTq6_0(.dout(w_dff_A_COmVAiYt6_0),.din(w_dff_A_uHsWKiTq6_0),.clk(gclk));
	jdff dff_A_COmVAiYt6_0(.dout(w_dff_A_OB4xrie35_0),.din(w_dff_A_COmVAiYt6_0),.clk(gclk));
	jdff dff_A_OB4xrie35_0(.dout(w_dff_A_4cazQZu34_0),.din(w_dff_A_OB4xrie35_0),.clk(gclk));
	jdff dff_A_4cazQZu34_0(.dout(w_dff_A_Azxin5gJ9_0),.din(w_dff_A_4cazQZu34_0),.clk(gclk));
	jdff dff_A_Azxin5gJ9_0(.dout(w_dff_A_uNKUOqjj9_0),.din(w_dff_A_Azxin5gJ9_0),.clk(gclk));
	jdff dff_A_uNKUOqjj9_0(.dout(w_dff_A_nUDK1cDz3_0),.din(w_dff_A_uNKUOqjj9_0),.clk(gclk));
	jdff dff_A_nUDK1cDz3_0(.dout(w_dff_A_YKtJb5iH1_0),.din(w_dff_A_nUDK1cDz3_0),.clk(gclk));
	jdff dff_A_YKtJb5iH1_0(.dout(w_dff_A_AB1fkHal0_0),.din(w_dff_A_YKtJb5iH1_0),.clk(gclk));
	jdff dff_A_AB1fkHal0_0(.dout(w_dff_A_YJKu4n7R1_0),.din(w_dff_A_AB1fkHal0_0),.clk(gclk));
	jdff dff_A_YJKu4n7R1_0(.dout(w_dff_A_JQOtpg7T5_0),.din(w_dff_A_YJKu4n7R1_0),.clk(gclk));
	jdff dff_A_JQOtpg7T5_0(.dout(w_dff_A_2l7LCQqd5_0),.din(w_dff_A_JQOtpg7T5_0),.clk(gclk));
	jdff dff_A_2l7LCQqd5_0(.dout(w_dff_A_xLawbqg44_0),.din(w_dff_A_2l7LCQqd5_0),.clk(gclk));
	jdff dff_A_xLawbqg44_0(.dout(w_dff_A_TI0CfsI76_0),.din(w_dff_A_xLawbqg44_0),.clk(gclk));
	jdff dff_A_TI0CfsI76_0(.dout(w_dff_A_TyRnyetE3_0),.din(w_dff_A_TI0CfsI76_0),.clk(gclk));
	jdff dff_A_TyRnyetE3_0(.dout(w_dff_A_EjvaFcqK0_0),.din(w_dff_A_TyRnyetE3_0),.clk(gclk));
	jdff dff_A_EjvaFcqK0_0(.dout(w_dff_A_RImng3S02_0),.din(w_dff_A_EjvaFcqK0_0),.clk(gclk));
	jdff dff_A_RImng3S02_0(.dout(w_dff_A_0zcSSwgI6_0),.din(w_dff_A_RImng3S02_0),.clk(gclk));
	jdff dff_A_0zcSSwgI6_0(.dout(G522),.din(w_dff_A_0zcSSwgI6_0),.clk(gclk));
	jdff dff_A_l29pao1a2_2(.dout(w_dff_A_vpHsIN2M8_0),.din(w_dff_A_l29pao1a2_2),.clk(gclk));
	jdff dff_A_vpHsIN2M8_0(.dout(w_dff_A_twkstNKm7_0),.din(w_dff_A_vpHsIN2M8_0),.clk(gclk));
	jdff dff_A_twkstNKm7_0(.dout(w_dff_A_o8UYQHkv5_0),.din(w_dff_A_twkstNKm7_0),.clk(gclk));
	jdff dff_A_o8UYQHkv5_0(.dout(w_dff_A_Z72aivL71_0),.din(w_dff_A_o8UYQHkv5_0),.clk(gclk));
	jdff dff_A_Z72aivL71_0(.dout(w_dff_A_VR5xCiLY6_0),.din(w_dff_A_Z72aivL71_0),.clk(gclk));
	jdff dff_A_VR5xCiLY6_0(.dout(w_dff_A_puoj0En35_0),.din(w_dff_A_VR5xCiLY6_0),.clk(gclk));
	jdff dff_A_puoj0En35_0(.dout(w_dff_A_ftHEnxS79_0),.din(w_dff_A_puoj0En35_0),.clk(gclk));
	jdff dff_A_ftHEnxS79_0(.dout(w_dff_A_CW0krvaF6_0),.din(w_dff_A_ftHEnxS79_0),.clk(gclk));
	jdff dff_A_CW0krvaF6_0(.dout(w_dff_A_trhOOQNj2_0),.din(w_dff_A_CW0krvaF6_0),.clk(gclk));
	jdff dff_A_trhOOQNj2_0(.dout(w_dff_A_onFXXuws4_0),.din(w_dff_A_trhOOQNj2_0),.clk(gclk));
	jdff dff_A_onFXXuws4_0(.dout(w_dff_A_cvvdYd0z6_0),.din(w_dff_A_onFXXuws4_0),.clk(gclk));
	jdff dff_A_cvvdYd0z6_0(.dout(w_dff_A_qDjEyS7M6_0),.din(w_dff_A_cvvdYd0z6_0),.clk(gclk));
	jdff dff_A_qDjEyS7M6_0(.dout(w_dff_A_qHCHfUXE1_0),.din(w_dff_A_qDjEyS7M6_0),.clk(gclk));
	jdff dff_A_qHCHfUXE1_0(.dout(w_dff_A_RhaAMeBP5_0),.din(w_dff_A_qHCHfUXE1_0),.clk(gclk));
	jdff dff_A_RhaAMeBP5_0(.dout(w_dff_A_MbwJ5eIo9_0),.din(w_dff_A_RhaAMeBP5_0),.clk(gclk));
	jdff dff_A_MbwJ5eIo9_0(.dout(w_dff_A_r595fPhb1_0),.din(w_dff_A_MbwJ5eIo9_0),.clk(gclk));
	jdff dff_A_r595fPhb1_0(.dout(w_dff_A_aODRENxC7_0),.din(w_dff_A_r595fPhb1_0),.clk(gclk));
	jdff dff_A_aODRENxC7_0(.dout(w_dff_A_Y3mPe2o84_0),.din(w_dff_A_aODRENxC7_0),.clk(gclk));
	jdff dff_A_Y3mPe2o84_0(.dout(w_dff_A_LKkzhW2h4_0),.din(w_dff_A_Y3mPe2o84_0),.clk(gclk));
	jdff dff_A_LKkzhW2h4_0(.dout(w_dff_A_O1Uh8qCm5_0),.din(w_dff_A_LKkzhW2h4_0),.clk(gclk));
	jdff dff_A_O1Uh8qCm5_0(.dout(w_dff_A_IMhJg36c7_0),.din(w_dff_A_O1Uh8qCm5_0),.clk(gclk));
	jdff dff_A_IMhJg36c7_0(.dout(w_dff_A_NS5V6sgc8_0),.din(w_dff_A_IMhJg36c7_0),.clk(gclk));
	jdff dff_A_NS5V6sgc8_0(.dout(w_dff_A_ip84immA1_0),.din(w_dff_A_NS5V6sgc8_0),.clk(gclk));
	jdff dff_A_ip84immA1_0(.dout(w_dff_A_1ua8GXzo3_0),.din(w_dff_A_ip84immA1_0),.clk(gclk));
	jdff dff_A_1ua8GXzo3_0(.dout(w_dff_A_mVzlf2gk4_0),.din(w_dff_A_1ua8GXzo3_0),.clk(gclk));
	jdff dff_A_mVzlf2gk4_0(.dout(w_dff_A_eI88lScm7_0),.din(w_dff_A_mVzlf2gk4_0),.clk(gclk));
	jdff dff_A_eI88lScm7_0(.dout(w_dff_A_w4tfmbqf3_0),.din(w_dff_A_eI88lScm7_0),.clk(gclk));
	jdff dff_A_w4tfmbqf3_0(.dout(w_dff_A_TtIABepv9_0),.din(w_dff_A_w4tfmbqf3_0),.clk(gclk));
	jdff dff_A_TtIABepv9_0(.dout(w_dff_A_EJj0UGy71_0),.din(w_dff_A_TtIABepv9_0),.clk(gclk));
	jdff dff_A_EJj0UGy71_0(.dout(w_dff_A_ZCSFIX2b7_0),.din(w_dff_A_EJj0UGy71_0),.clk(gclk));
	jdff dff_A_ZCSFIX2b7_0(.dout(w_dff_A_xPWT8kjR8_0),.din(w_dff_A_ZCSFIX2b7_0),.clk(gclk));
	jdff dff_A_xPWT8kjR8_0(.dout(w_dff_A_IlJbGYVQ9_0),.din(w_dff_A_xPWT8kjR8_0),.clk(gclk));
	jdff dff_A_IlJbGYVQ9_0(.dout(w_dff_A_7mNEW4CC9_0),.din(w_dff_A_IlJbGYVQ9_0),.clk(gclk));
	jdff dff_A_7mNEW4CC9_0(.dout(w_dff_A_II3vq1OJ0_0),.din(w_dff_A_7mNEW4CC9_0),.clk(gclk));
	jdff dff_A_II3vq1OJ0_0(.dout(w_dff_A_KOVwRCJu8_0),.din(w_dff_A_II3vq1OJ0_0),.clk(gclk));
	jdff dff_A_KOVwRCJu8_0(.dout(w_dff_A_SeCEcx126_0),.din(w_dff_A_KOVwRCJu8_0),.clk(gclk));
	jdff dff_A_SeCEcx126_0(.dout(w_dff_A_fskGHtJ71_0),.din(w_dff_A_SeCEcx126_0),.clk(gclk));
	jdff dff_A_fskGHtJ71_0(.dout(G402),.din(w_dff_A_fskGHtJ71_0),.clk(gclk));
	jdff dff_A_f9BvEB0p2_1(.dout(w_dff_A_QmFN9ecY0_0),.din(w_dff_A_f9BvEB0p2_1),.clk(gclk));
	jdff dff_A_QmFN9ecY0_0(.dout(w_dff_A_ABvL59jj2_0),.din(w_dff_A_QmFN9ecY0_0),.clk(gclk));
	jdff dff_A_ABvL59jj2_0(.dout(w_dff_A_2Q5aWDyp0_0),.din(w_dff_A_ABvL59jj2_0),.clk(gclk));
	jdff dff_A_2Q5aWDyp0_0(.dout(w_dff_A_G2h1cVhs3_0),.din(w_dff_A_2Q5aWDyp0_0),.clk(gclk));
	jdff dff_A_G2h1cVhs3_0(.dout(w_dff_A_9x4m3eGD3_0),.din(w_dff_A_G2h1cVhs3_0),.clk(gclk));
	jdff dff_A_9x4m3eGD3_0(.dout(w_dff_A_QTuckQAp2_0),.din(w_dff_A_9x4m3eGD3_0),.clk(gclk));
	jdff dff_A_QTuckQAp2_0(.dout(w_dff_A_ChHE3GpA4_0),.din(w_dff_A_QTuckQAp2_0),.clk(gclk));
	jdff dff_A_ChHE3GpA4_0(.dout(w_dff_A_uL8ms4jz8_0),.din(w_dff_A_ChHE3GpA4_0),.clk(gclk));
	jdff dff_A_uL8ms4jz8_0(.dout(w_dff_A_rz2Tsc6i4_0),.din(w_dff_A_uL8ms4jz8_0),.clk(gclk));
	jdff dff_A_rz2Tsc6i4_0(.dout(w_dff_A_4s3dByA95_0),.din(w_dff_A_rz2Tsc6i4_0),.clk(gclk));
	jdff dff_A_4s3dByA95_0(.dout(w_dff_A_04nuj0MO6_0),.din(w_dff_A_4s3dByA95_0),.clk(gclk));
	jdff dff_A_04nuj0MO6_0(.dout(w_dff_A_lq2F7Xmy0_0),.din(w_dff_A_04nuj0MO6_0),.clk(gclk));
	jdff dff_A_lq2F7Xmy0_0(.dout(w_dff_A_hayGb6pg4_0),.din(w_dff_A_lq2F7Xmy0_0),.clk(gclk));
	jdff dff_A_hayGb6pg4_0(.dout(w_dff_A_sGDSKULh9_0),.din(w_dff_A_hayGb6pg4_0),.clk(gclk));
	jdff dff_A_sGDSKULh9_0(.dout(w_dff_A_N6ev3BFD3_0),.din(w_dff_A_sGDSKULh9_0),.clk(gclk));
	jdff dff_A_N6ev3BFD3_0(.dout(w_dff_A_8Oaw93Af3_0),.din(w_dff_A_N6ev3BFD3_0),.clk(gclk));
	jdff dff_A_8Oaw93Af3_0(.dout(w_dff_A_S4oO2WE52_0),.din(w_dff_A_8Oaw93Af3_0),.clk(gclk));
	jdff dff_A_S4oO2WE52_0(.dout(w_dff_A_vdtiLAcA9_0),.din(w_dff_A_S4oO2WE52_0),.clk(gclk));
	jdff dff_A_vdtiLAcA9_0(.dout(w_dff_A_OLhZKdKE8_0),.din(w_dff_A_vdtiLAcA9_0),.clk(gclk));
	jdff dff_A_OLhZKdKE8_0(.dout(w_dff_A_jnYdKqCs7_0),.din(w_dff_A_OLhZKdKE8_0),.clk(gclk));
	jdff dff_A_jnYdKqCs7_0(.dout(w_dff_A_skrNjDKt5_0),.din(w_dff_A_jnYdKqCs7_0),.clk(gclk));
	jdff dff_A_skrNjDKt5_0(.dout(w_dff_A_PcC3T0l90_0),.din(w_dff_A_skrNjDKt5_0),.clk(gclk));
	jdff dff_A_PcC3T0l90_0(.dout(w_dff_A_eHZ51nIy2_0),.din(w_dff_A_PcC3T0l90_0),.clk(gclk));
	jdff dff_A_eHZ51nIy2_0(.dout(w_dff_A_e7UtXRq43_0),.din(w_dff_A_eHZ51nIy2_0),.clk(gclk));
	jdff dff_A_e7UtXRq43_0(.dout(w_dff_A_B5iqlsxA6_0),.din(w_dff_A_e7UtXRq43_0),.clk(gclk));
	jdff dff_A_B5iqlsxA6_0(.dout(w_dff_A_UCla0D5N8_0),.din(w_dff_A_B5iqlsxA6_0),.clk(gclk));
	jdff dff_A_UCla0D5N8_0(.dout(w_dff_A_AVUd1WYq7_0),.din(w_dff_A_UCla0D5N8_0),.clk(gclk));
	jdff dff_A_AVUd1WYq7_0(.dout(w_dff_A_sWaSxgmF6_0),.din(w_dff_A_AVUd1WYq7_0),.clk(gclk));
	jdff dff_A_sWaSxgmF6_0(.dout(w_dff_A_JshhyMeG4_0),.din(w_dff_A_sWaSxgmF6_0),.clk(gclk));
	jdff dff_A_JshhyMeG4_0(.dout(w_dff_A_WPCzSxIp7_0),.din(w_dff_A_JshhyMeG4_0),.clk(gclk));
	jdff dff_A_WPCzSxIp7_0(.dout(w_dff_A_fRz2Ewyi3_0),.din(w_dff_A_WPCzSxIp7_0),.clk(gclk));
	jdff dff_A_fRz2Ewyi3_0(.dout(w_dff_A_nNAPGyfd0_0),.din(w_dff_A_fRz2Ewyi3_0),.clk(gclk));
	jdff dff_A_nNAPGyfd0_0(.dout(w_dff_A_n9nueMw50_0),.din(w_dff_A_nNAPGyfd0_0),.clk(gclk));
	jdff dff_A_n9nueMw50_0(.dout(w_dff_A_q3x932343_0),.din(w_dff_A_n9nueMw50_0),.clk(gclk));
	jdff dff_A_q3x932343_0(.dout(w_dff_A_mGOYjGEC3_0),.din(w_dff_A_q3x932343_0),.clk(gclk));
	jdff dff_A_mGOYjGEC3_0(.dout(G404),.din(w_dff_A_mGOYjGEC3_0),.clk(gclk));
	jdff dff_A_cVJigQ0M0_1(.dout(w_dff_A_UUcobrs82_0),.din(w_dff_A_cVJigQ0M0_1),.clk(gclk));
	jdff dff_A_UUcobrs82_0(.dout(w_dff_A_DK6Wrpyk9_0),.din(w_dff_A_UUcobrs82_0),.clk(gclk));
	jdff dff_A_DK6Wrpyk9_0(.dout(w_dff_A_7G9uf8QO5_0),.din(w_dff_A_DK6Wrpyk9_0),.clk(gclk));
	jdff dff_A_7G9uf8QO5_0(.dout(w_dff_A_nkDNo1se6_0),.din(w_dff_A_7G9uf8QO5_0),.clk(gclk));
	jdff dff_A_nkDNo1se6_0(.dout(w_dff_A_h81KICLp8_0),.din(w_dff_A_nkDNo1se6_0),.clk(gclk));
	jdff dff_A_h81KICLp8_0(.dout(w_dff_A_nioisLAD5_0),.din(w_dff_A_h81KICLp8_0),.clk(gclk));
	jdff dff_A_nioisLAD5_0(.dout(w_dff_A_LJlZtDij9_0),.din(w_dff_A_nioisLAD5_0),.clk(gclk));
	jdff dff_A_LJlZtDij9_0(.dout(w_dff_A_813iFHv09_0),.din(w_dff_A_LJlZtDij9_0),.clk(gclk));
	jdff dff_A_813iFHv09_0(.dout(w_dff_A_axJ7XbcL9_0),.din(w_dff_A_813iFHv09_0),.clk(gclk));
	jdff dff_A_axJ7XbcL9_0(.dout(w_dff_A_0oRzjyim8_0),.din(w_dff_A_axJ7XbcL9_0),.clk(gclk));
	jdff dff_A_0oRzjyim8_0(.dout(w_dff_A_Vdx44zb02_0),.din(w_dff_A_0oRzjyim8_0),.clk(gclk));
	jdff dff_A_Vdx44zb02_0(.dout(w_dff_A_nMldML9W4_0),.din(w_dff_A_Vdx44zb02_0),.clk(gclk));
	jdff dff_A_nMldML9W4_0(.dout(w_dff_A_kc4iEzfq2_0),.din(w_dff_A_nMldML9W4_0),.clk(gclk));
	jdff dff_A_kc4iEzfq2_0(.dout(w_dff_A_HeU802GO1_0),.din(w_dff_A_kc4iEzfq2_0),.clk(gclk));
	jdff dff_A_HeU802GO1_0(.dout(w_dff_A_xoKHy0wl1_0),.din(w_dff_A_HeU802GO1_0),.clk(gclk));
	jdff dff_A_xoKHy0wl1_0(.dout(w_dff_A_jneBexU33_0),.din(w_dff_A_xoKHy0wl1_0),.clk(gclk));
	jdff dff_A_jneBexU33_0(.dout(w_dff_A_DZpTgcTD7_0),.din(w_dff_A_jneBexU33_0),.clk(gclk));
	jdff dff_A_DZpTgcTD7_0(.dout(w_dff_A_kaSynU7e8_0),.din(w_dff_A_DZpTgcTD7_0),.clk(gclk));
	jdff dff_A_kaSynU7e8_0(.dout(w_dff_A_AzYZCCN58_0),.din(w_dff_A_kaSynU7e8_0),.clk(gclk));
	jdff dff_A_AzYZCCN58_0(.dout(w_dff_A_GlViQ2a47_0),.din(w_dff_A_AzYZCCN58_0),.clk(gclk));
	jdff dff_A_GlViQ2a47_0(.dout(w_dff_A_DDb3mBxp7_0),.din(w_dff_A_GlViQ2a47_0),.clk(gclk));
	jdff dff_A_DDb3mBxp7_0(.dout(w_dff_A_IWg0Q6zc7_0),.din(w_dff_A_DDb3mBxp7_0),.clk(gclk));
	jdff dff_A_IWg0Q6zc7_0(.dout(w_dff_A_NafJUaX61_0),.din(w_dff_A_IWg0Q6zc7_0),.clk(gclk));
	jdff dff_A_NafJUaX61_0(.dout(w_dff_A_MuXb125O4_0),.din(w_dff_A_NafJUaX61_0),.clk(gclk));
	jdff dff_A_MuXb125O4_0(.dout(w_dff_A_w8SPfYI32_0),.din(w_dff_A_MuXb125O4_0),.clk(gclk));
	jdff dff_A_w8SPfYI32_0(.dout(w_dff_A_ctGLWZTc9_0),.din(w_dff_A_w8SPfYI32_0),.clk(gclk));
	jdff dff_A_ctGLWZTc9_0(.dout(w_dff_A_RMUWSGP52_0),.din(w_dff_A_ctGLWZTc9_0),.clk(gclk));
	jdff dff_A_RMUWSGP52_0(.dout(w_dff_A_9tM1MDuc0_0),.din(w_dff_A_RMUWSGP52_0),.clk(gclk));
	jdff dff_A_9tM1MDuc0_0(.dout(w_dff_A_A7nEpr661_0),.din(w_dff_A_9tM1MDuc0_0),.clk(gclk));
	jdff dff_A_A7nEpr661_0(.dout(w_dff_A_VHpXnndZ9_0),.din(w_dff_A_A7nEpr661_0),.clk(gclk));
	jdff dff_A_VHpXnndZ9_0(.dout(w_dff_A_ooj0XJgm7_0),.din(w_dff_A_VHpXnndZ9_0),.clk(gclk));
	jdff dff_A_ooj0XJgm7_0(.dout(w_dff_A_vCu00N991_0),.din(w_dff_A_ooj0XJgm7_0),.clk(gclk));
	jdff dff_A_vCu00N991_0(.dout(w_dff_A_HlqCQLAY6_0),.din(w_dff_A_vCu00N991_0),.clk(gclk));
	jdff dff_A_HlqCQLAY6_0(.dout(w_dff_A_rg1a1AVl8_0),.din(w_dff_A_HlqCQLAY6_0),.clk(gclk));
	jdff dff_A_rg1a1AVl8_0(.dout(w_dff_A_7zVj4Qf74_0),.din(w_dff_A_rg1a1AVl8_0),.clk(gclk));
	jdff dff_A_7zVj4Qf74_0(.dout(G406),.din(w_dff_A_7zVj4Qf74_0),.clk(gclk));
	jdff dff_A_uXZKF6Yh3_1(.dout(w_dff_A_QAPZCd5D5_0),.din(w_dff_A_uXZKF6Yh3_1),.clk(gclk));
	jdff dff_A_QAPZCd5D5_0(.dout(w_dff_A_wGjYtbn99_0),.din(w_dff_A_QAPZCd5D5_0),.clk(gclk));
	jdff dff_A_wGjYtbn99_0(.dout(w_dff_A_p4seJZne1_0),.din(w_dff_A_wGjYtbn99_0),.clk(gclk));
	jdff dff_A_p4seJZne1_0(.dout(w_dff_A_dzeNiATj5_0),.din(w_dff_A_p4seJZne1_0),.clk(gclk));
	jdff dff_A_dzeNiATj5_0(.dout(w_dff_A_NzNxO6yS0_0),.din(w_dff_A_dzeNiATj5_0),.clk(gclk));
	jdff dff_A_NzNxO6yS0_0(.dout(w_dff_A_ABdOXtSb4_0),.din(w_dff_A_NzNxO6yS0_0),.clk(gclk));
	jdff dff_A_ABdOXtSb4_0(.dout(w_dff_A_BE4Jz0VU6_0),.din(w_dff_A_ABdOXtSb4_0),.clk(gclk));
	jdff dff_A_BE4Jz0VU6_0(.dout(w_dff_A_hpHsj7jz7_0),.din(w_dff_A_BE4Jz0VU6_0),.clk(gclk));
	jdff dff_A_hpHsj7jz7_0(.dout(w_dff_A_6NEzPVXR5_0),.din(w_dff_A_hpHsj7jz7_0),.clk(gclk));
	jdff dff_A_6NEzPVXR5_0(.dout(w_dff_A_UFzQSGYo5_0),.din(w_dff_A_6NEzPVXR5_0),.clk(gclk));
	jdff dff_A_UFzQSGYo5_0(.dout(w_dff_A_CzELws3Q1_0),.din(w_dff_A_UFzQSGYo5_0),.clk(gclk));
	jdff dff_A_CzELws3Q1_0(.dout(w_dff_A_lu92C5VG8_0),.din(w_dff_A_CzELws3Q1_0),.clk(gclk));
	jdff dff_A_lu92C5VG8_0(.dout(w_dff_A_fVmzrn5z1_0),.din(w_dff_A_lu92C5VG8_0),.clk(gclk));
	jdff dff_A_fVmzrn5z1_0(.dout(w_dff_A_FjVfwBkm4_0),.din(w_dff_A_fVmzrn5z1_0),.clk(gclk));
	jdff dff_A_FjVfwBkm4_0(.dout(w_dff_A_2CaVv1wK5_0),.din(w_dff_A_FjVfwBkm4_0),.clk(gclk));
	jdff dff_A_2CaVv1wK5_0(.dout(w_dff_A_jTZG1E9T2_0),.din(w_dff_A_2CaVv1wK5_0),.clk(gclk));
	jdff dff_A_jTZG1E9T2_0(.dout(w_dff_A_LgsP8qEz8_0),.din(w_dff_A_jTZG1E9T2_0),.clk(gclk));
	jdff dff_A_LgsP8qEz8_0(.dout(w_dff_A_cPj50RB71_0),.din(w_dff_A_LgsP8qEz8_0),.clk(gclk));
	jdff dff_A_cPj50RB71_0(.dout(w_dff_A_9BFB27r18_0),.din(w_dff_A_cPj50RB71_0),.clk(gclk));
	jdff dff_A_9BFB27r18_0(.dout(w_dff_A_pMPG5zP03_0),.din(w_dff_A_9BFB27r18_0),.clk(gclk));
	jdff dff_A_pMPG5zP03_0(.dout(w_dff_A_XaLre3FV2_0),.din(w_dff_A_pMPG5zP03_0),.clk(gclk));
	jdff dff_A_XaLre3FV2_0(.dout(w_dff_A_6Ei26ZAL3_0),.din(w_dff_A_XaLre3FV2_0),.clk(gclk));
	jdff dff_A_6Ei26ZAL3_0(.dout(w_dff_A_cKqrvQBg8_0),.din(w_dff_A_6Ei26ZAL3_0),.clk(gclk));
	jdff dff_A_cKqrvQBg8_0(.dout(w_dff_A_HJRmcQFq0_0),.din(w_dff_A_cKqrvQBg8_0),.clk(gclk));
	jdff dff_A_HJRmcQFq0_0(.dout(w_dff_A_FQcqCSdl9_0),.din(w_dff_A_HJRmcQFq0_0),.clk(gclk));
	jdff dff_A_FQcqCSdl9_0(.dout(w_dff_A_OvIeQQXb0_0),.din(w_dff_A_FQcqCSdl9_0),.clk(gclk));
	jdff dff_A_OvIeQQXb0_0(.dout(w_dff_A_qXxicUeF3_0),.din(w_dff_A_OvIeQQXb0_0),.clk(gclk));
	jdff dff_A_qXxicUeF3_0(.dout(w_dff_A_ms99laM27_0),.din(w_dff_A_qXxicUeF3_0),.clk(gclk));
	jdff dff_A_ms99laM27_0(.dout(w_dff_A_OjMdN8nn0_0),.din(w_dff_A_ms99laM27_0),.clk(gclk));
	jdff dff_A_OjMdN8nn0_0(.dout(w_dff_A_SSDbt0Ut6_0),.din(w_dff_A_OjMdN8nn0_0),.clk(gclk));
	jdff dff_A_SSDbt0Ut6_0(.dout(w_dff_A_gZ5rN5JU7_0),.din(w_dff_A_SSDbt0Ut6_0),.clk(gclk));
	jdff dff_A_gZ5rN5JU7_0(.dout(w_dff_A_1KAVeFYD7_0),.din(w_dff_A_gZ5rN5JU7_0),.clk(gclk));
	jdff dff_A_1KAVeFYD7_0(.dout(w_dff_A_oG7cPQNU3_0),.din(w_dff_A_1KAVeFYD7_0),.clk(gclk));
	jdff dff_A_oG7cPQNU3_0(.dout(w_dff_A_A0RuoFMe1_0),.din(w_dff_A_oG7cPQNU3_0),.clk(gclk));
	jdff dff_A_A0RuoFMe1_0(.dout(w_dff_A_SzsJbbxU2_0),.din(w_dff_A_A0RuoFMe1_0),.clk(gclk));
	jdff dff_A_SzsJbbxU2_0(.dout(G408),.din(w_dff_A_SzsJbbxU2_0),.clk(gclk));
	jdff dff_A_vLRVPHpJ9_1(.dout(w_dff_A_pETu6NWu8_0),.din(w_dff_A_vLRVPHpJ9_1),.clk(gclk));
	jdff dff_A_pETu6NWu8_0(.dout(w_dff_A_0q4VzV568_0),.din(w_dff_A_pETu6NWu8_0),.clk(gclk));
	jdff dff_A_0q4VzV568_0(.dout(w_dff_A_LCWWeUNO3_0),.din(w_dff_A_0q4VzV568_0),.clk(gclk));
	jdff dff_A_LCWWeUNO3_0(.dout(w_dff_A_x6jMIy466_0),.din(w_dff_A_LCWWeUNO3_0),.clk(gclk));
	jdff dff_A_x6jMIy466_0(.dout(w_dff_A_fKMs039R1_0),.din(w_dff_A_x6jMIy466_0),.clk(gclk));
	jdff dff_A_fKMs039R1_0(.dout(w_dff_A_ZtjpM78x7_0),.din(w_dff_A_fKMs039R1_0),.clk(gclk));
	jdff dff_A_ZtjpM78x7_0(.dout(w_dff_A_l4xmYpXr7_0),.din(w_dff_A_ZtjpM78x7_0),.clk(gclk));
	jdff dff_A_l4xmYpXr7_0(.dout(w_dff_A_90B53fqI6_0),.din(w_dff_A_l4xmYpXr7_0),.clk(gclk));
	jdff dff_A_90B53fqI6_0(.dout(w_dff_A_VorGZjvp6_0),.din(w_dff_A_90B53fqI6_0),.clk(gclk));
	jdff dff_A_VorGZjvp6_0(.dout(w_dff_A_MF5KCvsH8_0),.din(w_dff_A_VorGZjvp6_0),.clk(gclk));
	jdff dff_A_MF5KCvsH8_0(.dout(w_dff_A_3KFt32vo5_0),.din(w_dff_A_MF5KCvsH8_0),.clk(gclk));
	jdff dff_A_3KFt32vo5_0(.dout(w_dff_A_Bygal0ww1_0),.din(w_dff_A_3KFt32vo5_0),.clk(gclk));
	jdff dff_A_Bygal0ww1_0(.dout(w_dff_A_OLmDZgpm8_0),.din(w_dff_A_Bygal0ww1_0),.clk(gclk));
	jdff dff_A_OLmDZgpm8_0(.dout(w_dff_A_WFWLv4Ef7_0),.din(w_dff_A_OLmDZgpm8_0),.clk(gclk));
	jdff dff_A_WFWLv4Ef7_0(.dout(w_dff_A_yCfeM25i3_0),.din(w_dff_A_WFWLv4Ef7_0),.clk(gclk));
	jdff dff_A_yCfeM25i3_0(.dout(w_dff_A_RafLgjDR8_0),.din(w_dff_A_yCfeM25i3_0),.clk(gclk));
	jdff dff_A_RafLgjDR8_0(.dout(w_dff_A_VngPkwI53_0),.din(w_dff_A_RafLgjDR8_0),.clk(gclk));
	jdff dff_A_VngPkwI53_0(.dout(w_dff_A_vsN2pBpa8_0),.din(w_dff_A_VngPkwI53_0),.clk(gclk));
	jdff dff_A_vsN2pBpa8_0(.dout(w_dff_A_8nALCqNr5_0),.din(w_dff_A_vsN2pBpa8_0),.clk(gclk));
	jdff dff_A_8nALCqNr5_0(.dout(w_dff_A_bUTpaOBi0_0),.din(w_dff_A_8nALCqNr5_0),.clk(gclk));
	jdff dff_A_bUTpaOBi0_0(.dout(w_dff_A_jBOyfPDn4_0),.din(w_dff_A_bUTpaOBi0_0),.clk(gclk));
	jdff dff_A_jBOyfPDn4_0(.dout(w_dff_A_LvD3dYgc2_0),.din(w_dff_A_jBOyfPDn4_0),.clk(gclk));
	jdff dff_A_LvD3dYgc2_0(.dout(w_dff_A_ze9uco4J0_0),.din(w_dff_A_LvD3dYgc2_0),.clk(gclk));
	jdff dff_A_ze9uco4J0_0(.dout(w_dff_A_1mImsz3t5_0),.din(w_dff_A_ze9uco4J0_0),.clk(gclk));
	jdff dff_A_1mImsz3t5_0(.dout(w_dff_A_zdcSQLJZ4_0),.din(w_dff_A_1mImsz3t5_0),.clk(gclk));
	jdff dff_A_zdcSQLJZ4_0(.dout(w_dff_A_CSmIodxh4_0),.din(w_dff_A_zdcSQLJZ4_0),.clk(gclk));
	jdff dff_A_CSmIodxh4_0(.dout(w_dff_A_QauGlLGA8_0),.din(w_dff_A_CSmIodxh4_0),.clk(gclk));
	jdff dff_A_QauGlLGA8_0(.dout(w_dff_A_ajnPqiCO0_0),.din(w_dff_A_QauGlLGA8_0),.clk(gclk));
	jdff dff_A_ajnPqiCO0_0(.dout(w_dff_A_VGbi1yME3_0),.din(w_dff_A_ajnPqiCO0_0),.clk(gclk));
	jdff dff_A_VGbi1yME3_0(.dout(w_dff_A_JNv0kTSU6_0),.din(w_dff_A_VGbi1yME3_0),.clk(gclk));
	jdff dff_A_JNv0kTSU6_0(.dout(w_dff_A_larRg07u8_0),.din(w_dff_A_JNv0kTSU6_0),.clk(gclk));
	jdff dff_A_larRg07u8_0(.dout(w_dff_A_CBsy12Sx9_0),.din(w_dff_A_larRg07u8_0),.clk(gclk));
	jdff dff_A_CBsy12Sx9_0(.dout(w_dff_A_Txxc89Ca1_0),.din(w_dff_A_CBsy12Sx9_0),.clk(gclk));
	jdff dff_A_Txxc89Ca1_0(.dout(w_dff_A_ZeCSr41v6_0),.din(w_dff_A_Txxc89Ca1_0),.clk(gclk));
	jdff dff_A_ZeCSr41v6_0(.dout(w_dff_A_BviXlD0x7_0),.din(w_dff_A_ZeCSr41v6_0),.clk(gclk));
	jdff dff_A_BviXlD0x7_0(.dout(G410),.din(w_dff_A_BviXlD0x7_0),.clk(gclk));
	jdff dff_A_UmRpndW02_1(.dout(w_dff_A_g6aYWzKz7_0),.din(w_dff_A_UmRpndW02_1),.clk(gclk));
	jdff dff_A_g6aYWzKz7_0(.dout(w_dff_A_iNeR9I6u7_0),.din(w_dff_A_g6aYWzKz7_0),.clk(gclk));
	jdff dff_A_iNeR9I6u7_0(.dout(w_dff_A_SgN08v1v3_0),.din(w_dff_A_iNeR9I6u7_0),.clk(gclk));
	jdff dff_A_SgN08v1v3_0(.dout(w_dff_A_rINHG92u2_0),.din(w_dff_A_SgN08v1v3_0),.clk(gclk));
	jdff dff_A_rINHG92u2_0(.dout(w_dff_A_lNY9aq9L3_0),.din(w_dff_A_rINHG92u2_0),.clk(gclk));
	jdff dff_A_lNY9aq9L3_0(.dout(w_dff_A_PU6oLifR3_0),.din(w_dff_A_lNY9aq9L3_0),.clk(gclk));
	jdff dff_A_PU6oLifR3_0(.dout(w_dff_A_PplyFSli5_0),.din(w_dff_A_PU6oLifR3_0),.clk(gclk));
	jdff dff_A_PplyFSli5_0(.dout(w_dff_A_7Ie371jD9_0),.din(w_dff_A_PplyFSli5_0),.clk(gclk));
	jdff dff_A_7Ie371jD9_0(.dout(w_dff_A_tQiVhEhr4_0),.din(w_dff_A_7Ie371jD9_0),.clk(gclk));
	jdff dff_A_tQiVhEhr4_0(.dout(w_dff_A_ECIM6ThG5_0),.din(w_dff_A_tQiVhEhr4_0),.clk(gclk));
	jdff dff_A_ECIM6ThG5_0(.dout(w_dff_A_lxKSkcwZ0_0),.din(w_dff_A_ECIM6ThG5_0),.clk(gclk));
	jdff dff_A_lxKSkcwZ0_0(.dout(w_dff_A_7idhb0VO5_0),.din(w_dff_A_lxKSkcwZ0_0),.clk(gclk));
	jdff dff_A_7idhb0VO5_0(.dout(w_dff_A_CYtfvawb0_0),.din(w_dff_A_7idhb0VO5_0),.clk(gclk));
	jdff dff_A_CYtfvawb0_0(.dout(w_dff_A_dC8Rr2P03_0),.din(w_dff_A_CYtfvawb0_0),.clk(gclk));
	jdff dff_A_dC8Rr2P03_0(.dout(w_dff_A_7QABMPlQ5_0),.din(w_dff_A_dC8Rr2P03_0),.clk(gclk));
	jdff dff_A_7QABMPlQ5_0(.dout(w_dff_A_36BMpCoG5_0),.din(w_dff_A_7QABMPlQ5_0),.clk(gclk));
	jdff dff_A_36BMpCoG5_0(.dout(w_dff_A_s1jtSIvt7_0),.din(w_dff_A_36BMpCoG5_0),.clk(gclk));
	jdff dff_A_s1jtSIvt7_0(.dout(w_dff_A_gnEyxGXA9_0),.din(w_dff_A_s1jtSIvt7_0),.clk(gclk));
	jdff dff_A_gnEyxGXA9_0(.dout(w_dff_A_4mUNCGDX5_0),.din(w_dff_A_gnEyxGXA9_0),.clk(gclk));
	jdff dff_A_4mUNCGDX5_0(.dout(w_dff_A_EerkGR6q7_0),.din(w_dff_A_4mUNCGDX5_0),.clk(gclk));
	jdff dff_A_EerkGR6q7_0(.dout(w_dff_A_jKNmD0wk7_0),.din(w_dff_A_EerkGR6q7_0),.clk(gclk));
	jdff dff_A_jKNmD0wk7_0(.dout(w_dff_A_cFHSo8kd3_0),.din(w_dff_A_jKNmD0wk7_0),.clk(gclk));
	jdff dff_A_cFHSo8kd3_0(.dout(w_dff_A_5hlrKPv12_0),.din(w_dff_A_cFHSo8kd3_0),.clk(gclk));
	jdff dff_A_5hlrKPv12_0(.dout(w_dff_A_HzBBmX0l4_0),.din(w_dff_A_5hlrKPv12_0),.clk(gclk));
	jdff dff_A_HzBBmX0l4_0(.dout(w_dff_A_P24sqcHi5_0),.din(w_dff_A_HzBBmX0l4_0),.clk(gclk));
	jdff dff_A_P24sqcHi5_0(.dout(w_dff_A_GtbN2OiQ3_0),.din(w_dff_A_P24sqcHi5_0),.clk(gclk));
	jdff dff_A_GtbN2OiQ3_0(.dout(w_dff_A_AVkXWHZx7_0),.din(w_dff_A_GtbN2OiQ3_0),.clk(gclk));
	jdff dff_A_AVkXWHZx7_0(.dout(w_dff_A_156IjwjA0_0),.din(w_dff_A_AVkXWHZx7_0),.clk(gclk));
	jdff dff_A_156IjwjA0_0(.dout(w_dff_A_13QnXjkB8_0),.din(w_dff_A_156IjwjA0_0),.clk(gclk));
	jdff dff_A_13QnXjkB8_0(.dout(w_dff_A_0D7KPyRq7_0),.din(w_dff_A_13QnXjkB8_0),.clk(gclk));
	jdff dff_A_0D7KPyRq7_0(.dout(w_dff_A_8JSeBPHl2_0),.din(w_dff_A_0D7KPyRq7_0),.clk(gclk));
	jdff dff_A_8JSeBPHl2_0(.dout(w_dff_A_Jkjwe1l57_0),.din(w_dff_A_8JSeBPHl2_0),.clk(gclk));
	jdff dff_A_Jkjwe1l57_0(.dout(w_dff_A_yOBfpf2J7_0),.din(w_dff_A_Jkjwe1l57_0),.clk(gclk));
	jdff dff_A_yOBfpf2J7_0(.dout(w_dff_A_8zlEVCJZ9_0),.din(w_dff_A_yOBfpf2J7_0),.clk(gclk));
	jdff dff_A_8zlEVCJZ9_0(.dout(w_dff_A_XZm1WecU4_0),.din(w_dff_A_8zlEVCJZ9_0),.clk(gclk));
	jdff dff_A_XZm1WecU4_0(.dout(w_dff_A_wXxqaB6A9_0),.din(w_dff_A_XZm1WecU4_0),.clk(gclk));
	jdff dff_A_wXxqaB6A9_0(.dout(w_dff_A_AtyoT8ZO0_0),.din(w_dff_A_wXxqaB6A9_0),.clk(gclk));
	jdff dff_A_AtyoT8ZO0_0(.dout(w_dff_A_olSL7hVn3_0),.din(w_dff_A_AtyoT8ZO0_0),.clk(gclk));
	jdff dff_A_olSL7hVn3_0(.dout(G432),.din(w_dff_A_olSL7hVn3_0),.clk(gclk));
	jdff dff_A_GvhcWMRm2_1(.dout(w_dff_A_8Nfw95BS7_0),.din(w_dff_A_GvhcWMRm2_1),.clk(gclk));
	jdff dff_A_8Nfw95BS7_0(.dout(w_dff_A_sYlMZort9_0),.din(w_dff_A_8Nfw95BS7_0),.clk(gclk));
	jdff dff_A_sYlMZort9_0(.dout(w_dff_A_LPUJtTLt0_0),.din(w_dff_A_sYlMZort9_0),.clk(gclk));
	jdff dff_A_LPUJtTLt0_0(.dout(w_dff_A_Mu5BzN2u8_0),.din(w_dff_A_LPUJtTLt0_0),.clk(gclk));
	jdff dff_A_Mu5BzN2u8_0(.dout(w_dff_A_8znLl8dS8_0),.din(w_dff_A_Mu5BzN2u8_0),.clk(gclk));
	jdff dff_A_8znLl8dS8_0(.dout(w_dff_A_HZ15V9MR7_0),.din(w_dff_A_8znLl8dS8_0),.clk(gclk));
	jdff dff_A_HZ15V9MR7_0(.dout(w_dff_A_HXvb78Tb1_0),.din(w_dff_A_HZ15V9MR7_0),.clk(gclk));
	jdff dff_A_HXvb78Tb1_0(.dout(w_dff_A_NhK5mDNZ6_0),.din(w_dff_A_HXvb78Tb1_0),.clk(gclk));
	jdff dff_A_NhK5mDNZ6_0(.dout(w_dff_A_7LhMwXib8_0),.din(w_dff_A_NhK5mDNZ6_0),.clk(gclk));
	jdff dff_A_7LhMwXib8_0(.dout(w_dff_A_69w0CmSt1_0),.din(w_dff_A_7LhMwXib8_0),.clk(gclk));
	jdff dff_A_69w0CmSt1_0(.dout(w_dff_A_0qmWonwJ3_0),.din(w_dff_A_69w0CmSt1_0),.clk(gclk));
	jdff dff_A_0qmWonwJ3_0(.dout(w_dff_A_asimPkSb1_0),.din(w_dff_A_0qmWonwJ3_0),.clk(gclk));
	jdff dff_A_asimPkSb1_0(.dout(w_dff_A_4eGrZ8K15_0),.din(w_dff_A_asimPkSb1_0),.clk(gclk));
	jdff dff_A_4eGrZ8K15_0(.dout(w_dff_A_8QLY8DaK4_0),.din(w_dff_A_4eGrZ8K15_0),.clk(gclk));
	jdff dff_A_8QLY8DaK4_0(.dout(w_dff_A_EF3nEqlO5_0),.din(w_dff_A_8QLY8DaK4_0),.clk(gclk));
	jdff dff_A_EF3nEqlO5_0(.dout(w_dff_A_IqDXQpKH1_0),.din(w_dff_A_EF3nEqlO5_0),.clk(gclk));
	jdff dff_A_IqDXQpKH1_0(.dout(w_dff_A_GIZWvFyN2_0),.din(w_dff_A_IqDXQpKH1_0),.clk(gclk));
	jdff dff_A_GIZWvFyN2_0(.dout(w_dff_A_HV7wdW6r1_0),.din(w_dff_A_GIZWvFyN2_0),.clk(gclk));
	jdff dff_A_HV7wdW6r1_0(.dout(w_dff_A_X6gXpop32_0),.din(w_dff_A_HV7wdW6r1_0),.clk(gclk));
	jdff dff_A_X6gXpop32_0(.dout(w_dff_A_d0h6NpRa9_0),.din(w_dff_A_X6gXpop32_0),.clk(gclk));
	jdff dff_A_d0h6NpRa9_0(.dout(w_dff_A_RDD70BOP3_0),.din(w_dff_A_d0h6NpRa9_0),.clk(gclk));
	jdff dff_A_RDD70BOP3_0(.dout(w_dff_A_bHDwJCfG7_0),.din(w_dff_A_RDD70BOP3_0),.clk(gclk));
	jdff dff_A_bHDwJCfG7_0(.dout(w_dff_A_YN49zphR2_0),.din(w_dff_A_bHDwJCfG7_0),.clk(gclk));
	jdff dff_A_YN49zphR2_0(.dout(w_dff_A_ch18PvVw0_0),.din(w_dff_A_YN49zphR2_0),.clk(gclk));
	jdff dff_A_ch18PvVw0_0(.dout(w_dff_A_YowinJjM0_0),.din(w_dff_A_ch18PvVw0_0),.clk(gclk));
	jdff dff_A_YowinJjM0_0(.dout(w_dff_A_nifW53gz9_0),.din(w_dff_A_YowinJjM0_0),.clk(gclk));
	jdff dff_A_nifW53gz9_0(.dout(w_dff_A_pzh1n70A3_0),.din(w_dff_A_nifW53gz9_0),.clk(gclk));
	jdff dff_A_pzh1n70A3_0(.dout(w_dff_A_MfXwBtvq8_0),.din(w_dff_A_pzh1n70A3_0),.clk(gclk));
	jdff dff_A_MfXwBtvq8_0(.dout(w_dff_A_teoyOoBm3_0),.din(w_dff_A_MfXwBtvq8_0),.clk(gclk));
	jdff dff_A_teoyOoBm3_0(.dout(w_dff_A_RF3bfCx54_0),.din(w_dff_A_teoyOoBm3_0),.clk(gclk));
	jdff dff_A_RF3bfCx54_0(.dout(w_dff_A_N9sllnDa5_0),.din(w_dff_A_RF3bfCx54_0),.clk(gclk));
	jdff dff_A_N9sllnDa5_0(.dout(w_dff_A_z4GtcDGJ2_0),.din(w_dff_A_N9sllnDa5_0),.clk(gclk));
	jdff dff_A_z4GtcDGJ2_0(.dout(w_dff_A_3iHvKG7B1_0),.din(w_dff_A_z4GtcDGJ2_0),.clk(gclk));
	jdff dff_A_3iHvKG7B1_0(.dout(w_dff_A_4k6m9DqR5_0),.din(w_dff_A_3iHvKG7B1_0),.clk(gclk));
	jdff dff_A_4k6m9DqR5_0(.dout(w_dff_A_B1CqK4mr5_0),.din(w_dff_A_4k6m9DqR5_0),.clk(gclk));
	jdff dff_A_B1CqK4mr5_0(.dout(w_dff_A_ebVxtHs96_0),.din(w_dff_A_B1CqK4mr5_0),.clk(gclk));
	jdff dff_A_ebVxtHs96_0(.dout(w_dff_A_StI7oTcp7_0),.din(w_dff_A_ebVxtHs96_0),.clk(gclk));
	jdff dff_A_StI7oTcp7_0(.dout(w_dff_A_u4outPN43_0),.din(w_dff_A_StI7oTcp7_0),.clk(gclk));
	jdff dff_A_u4outPN43_0(.dout(G446),.din(w_dff_A_u4outPN43_0),.clk(gclk));
	jdff dff_A_shAXd2VJ7_2(.dout(w_dff_A_sBOX5pMf4_0),.din(w_dff_A_shAXd2VJ7_2),.clk(gclk));
	jdff dff_A_sBOX5pMf4_0(.dout(w_dff_A_d8gA6SAU7_0),.din(w_dff_A_sBOX5pMf4_0),.clk(gclk));
	jdff dff_A_d8gA6SAU7_0(.dout(w_dff_A_POQLqnuM1_0),.din(w_dff_A_d8gA6SAU7_0),.clk(gclk));
	jdff dff_A_POQLqnuM1_0(.dout(w_dff_A_eSQrbb492_0),.din(w_dff_A_POQLqnuM1_0),.clk(gclk));
	jdff dff_A_eSQrbb492_0(.dout(w_dff_A_8Ea9HJjE5_0),.din(w_dff_A_eSQrbb492_0),.clk(gclk));
	jdff dff_A_8Ea9HJjE5_0(.dout(w_dff_A_Yixjxbt06_0),.din(w_dff_A_8Ea9HJjE5_0),.clk(gclk));
	jdff dff_A_Yixjxbt06_0(.dout(w_dff_A_vXgtixgr3_0),.din(w_dff_A_Yixjxbt06_0),.clk(gclk));
	jdff dff_A_vXgtixgr3_0(.dout(w_dff_A_psz6UQtf2_0),.din(w_dff_A_vXgtixgr3_0),.clk(gclk));
	jdff dff_A_psz6UQtf2_0(.dout(w_dff_A_4tNNQwRC4_0),.din(w_dff_A_psz6UQtf2_0),.clk(gclk));
	jdff dff_A_4tNNQwRC4_0(.dout(w_dff_A_qhHSbbHM5_0),.din(w_dff_A_4tNNQwRC4_0),.clk(gclk));
	jdff dff_A_qhHSbbHM5_0(.dout(w_dff_A_wFFAiIgn5_0),.din(w_dff_A_qhHSbbHM5_0),.clk(gclk));
	jdff dff_A_wFFAiIgn5_0(.dout(w_dff_A_axaXoooe0_0),.din(w_dff_A_wFFAiIgn5_0),.clk(gclk));
	jdff dff_A_axaXoooe0_0(.dout(w_dff_A_AmH0nBOK3_0),.din(w_dff_A_axaXoooe0_0),.clk(gclk));
	jdff dff_A_AmH0nBOK3_0(.dout(w_dff_A_mj3N1yxe0_0),.din(w_dff_A_AmH0nBOK3_0),.clk(gclk));
	jdff dff_A_mj3N1yxe0_0(.dout(w_dff_A_cyfgnMUv7_0),.din(w_dff_A_mj3N1yxe0_0),.clk(gclk));
	jdff dff_A_cyfgnMUv7_0(.dout(w_dff_A_ZptR4TQq8_0),.din(w_dff_A_cyfgnMUv7_0),.clk(gclk));
	jdff dff_A_ZptR4TQq8_0(.dout(w_dff_A_ZK6uJmzb0_0),.din(w_dff_A_ZptR4TQq8_0),.clk(gclk));
	jdff dff_A_ZK6uJmzb0_0(.dout(w_dff_A_VZSmSLFH6_0),.din(w_dff_A_ZK6uJmzb0_0),.clk(gclk));
	jdff dff_A_VZSmSLFH6_0(.dout(w_dff_A_GmlhfgGs2_0),.din(w_dff_A_VZSmSLFH6_0),.clk(gclk));
	jdff dff_A_GmlhfgGs2_0(.dout(w_dff_A_87i4wdCQ9_0),.din(w_dff_A_GmlhfgGs2_0),.clk(gclk));
	jdff dff_A_87i4wdCQ9_0(.dout(w_dff_A_5jRbM2bp8_0),.din(w_dff_A_87i4wdCQ9_0),.clk(gclk));
	jdff dff_A_5jRbM2bp8_0(.dout(w_dff_A_kv8hPPfP8_0),.din(w_dff_A_5jRbM2bp8_0),.clk(gclk));
	jdff dff_A_kv8hPPfP8_0(.dout(w_dff_A_CHkdAiIW0_0),.din(w_dff_A_kv8hPPfP8_0),.clk(gclk));
	jdff dff_A_CHkdAiIW0_0(.dout(w_dff_A_BzQBSkrh8_0),.din(w_dff_A_CHkdAiIW0_0),.clk(gclk));
	jdff dff_A_BzQBSkrh8_0(.dout(w_dff_A_lKYiOSZv8_0),.din(w_dff_A_BzQBSkrh8_0),.clk(gclk));
	jdff dff_A_lKYiOSZv8_0(.dout(w_dff_A_rB1y8qcf4_0),.din(w_dff_A_lKYiOSZv8_0),.clk(gclk));
	jdff dff_A_rB1y8qcf4_0(.dout(w_dff_A_5jWupdvD4_0),.din(w_dff_A_rB1y8qcf4_0),.clk(gclk));
	jdff dff_A_5jWupdvD4_0(.dout(w_dff_A_557gGvBh8_0),.din(w_dff_A_5jWupdvD4_0),.clk(gclk));
	jdff dff_A_557gGvBh8_0(.dout(w_dff_A_GhHtLrJ53_0),.din(w_dff_A_557gGvBh8_0),.clk(gclk));
	jdff dff_A_GhHtLrJ53_0(.dout(w_dff_A_F8mbicrI9_0),.din(w_dff_A_GhHtLrJ53_0),.clk(gclk));
	jdff dff_A_F8mbicrI9_0(.dout(w_dff_A_6USjyokI4_0),.din(w_dff_A_F8mbicrI9_0),.clk(gclk));
	jdff dff_A_6USjyokI4_0(.dout(w_dff_A_jLUQKHfc6_0),.din(w_dff_A_6USjyokI4_0),.clk(gclk));
	jdff dff_A_jLUQKHfc6_0(.dout(w_dff_A_L5JoTiLQ0_0),.din(w_dff_A_jLUQKHfc6_0),.clk(gclk));
	jdff dff_A_L5JoTiLQ0_0(.dout(w_dff_A_uFMOIDk74_0),.din(w_dff_A_L5JoTiLQ0_0),.clk(gclk));
	jdff dff_A_uFMOIDk74_0(.dout(w_dff_A_TD9z5fXV5_0),.din(w_dff_A_uFMOIDk74_0),.clk(gclk));
	jdff dff_A_TD9z5fXV5_0(.dout(w_dff_A_gOSHElLu0_0),.din(w_dff_A_TD9z5fXV5_0),.clk(gclk));
	jdff dff_A_gOSHElLu0_0(.dout(G284),.din(w_dff_A_gOSHElLu0_0),.clk(gclk));
	jdff dff_A_80dpXEcR8_1(.dout(w_dff_A_QtRn1iNZ1_0),.din(w_dff_A_80dpXEcR8_1),.clk(gclk));
	jdff dff_A_QtRn1iNZ1_0(.dout(w_dff_A_6f9MzD7l5_0),.din(w_dff_A_QtRn1iNZ1_0),.clk(gclk));
	jdff dff_A_6f9MzD7l5_0(.dout(w_dff_A_pyRvFWsR5_0),.din(w_dff_A_6f9MzD7l5_0),.clk(gclk));
	jdff dff_A_pyRvFWsR5_0(.dout(w_dff_A_iVauyqfL4_0),.din(w_dff_A_pyRvFWsR5_0),.clk(gclk));
	jdff dff_A_iVauyqfL4_0(.dout(w_dff_A_ivkVRNC56_0),.din(w_dff_A_iVauyqfL4_0),.clk(gclk));
	jdff dff_A_ivkVRNC56_0(.dout(w_dff_A_UlF54cb87_0),.din(w_dff_A_ivkVRNC56_0),.clk(gclk));
	jdff dff_A_UlF54cb87_0(.dout(w_dff_A_tkhvg9TS1_0),.din(w_dff_A_UlF54cb87_0),.clk(gclk));
	jdff dff_A_tkhvg9TS1_0(.dout(w_dff_A_10xolld75_0),.din(w_dff_A_tkhvg9TS1_0),.clk(gclk));
	jdff dff_A_10xolld75_0(.dout(w_dff_A_EVz7tDW14_0),.din(w_dff_A_10xolld75_0),.clk(gclk));
	jdff dff_A_EVz7tDW14_0(.dout(w_dff_A_iax3o9Jk5_0),.din(w_dff_A_EVz7tDW14_0),.clk(gclk));
	jdff dff_A_iax3o9Jk5_0(.dout(w_dff_A_ULKJWwH77_0),.din(w_dff_A_iax3o9Jk5_0),.clk(gclk));
	jdff dff_A_ULKJWwH77_0(.dout(w_dff_A_nrke1Mab4_0),.din(w_dff_A_ULKJWwH77_0),.clk(gclk));
	jdff dff_A_nrke1Mab4_0(.dout(w_dff_A_9oXUnIOz7_0),.din(w_dff_A_nrke1Mab4_0),.clk(gclk));
	jdff dff_A_9oXUnIOz7_0(.dout(w_dff_A_8LNW5BtM0_0),.din(w_dff_A_9oXUnIOz7_0),.clk(gclk));
	jdff dff_A_8LNW5BtM0_0(.dout(w_dff_A_TK7FDZtd3_0),.din(w_dff_A_8LNW5BtM0_0),.clk(gclk));
	jdff dff_A_TK7FDZtd3_0(.dout(w_dff_A_nNm2M1T17_0),.din(w_dff_A_TK7FDZtd3_0),.clk(gclk));
	jdff dff_A_nNm2M1T17_0(.dout(w_dff_A_ikf2zKF11_0),.din(w_dff_A_nNm2M1T17_0),.clk(gclk));
	jdff dff_A_ikf2zKF11_0(.dout(w_dff_A_VFjj4J008_0),.din(w_dff_A_ikf2zKF11_0),.clk(gclk));
	jdff dff_A_VFjj4J008_0(.dout(w_dff_A_Uhod3cOY3_0),.din(w_dff_A_VFjj4J008_0),.clk(gclk));
	jdff dff_A_Uhod3cOY3_0(.dout(w_dff_A_zpKaUDB92_0),.din(w_dff_A_Uhod3cOY3_0),.clk(gclk));
	jdff dff_A_zpKaUDB92_0(.dout(w_dff_A_LGuYaKgw8_0),.din(w_dff_A_zpKaUDB92_0),.clk(gclk));
	jdff dff_A_LGuYaKgw8_0(.dout(w_dff_A_UlWOZn0M5_0),.din(w_dff_A_LGuYaKgw8_0),.clk(gclk));
	jdff dff_A_UlWOZn0M5_0(.dout(w_dff_A_hIFWfd6U2_0),.din(w_dff_A_UlWOZn0M5_0),.clk(gclk));
	jdff dff_A_hIFWfd6U2_0(.dout(w_dff_A_WBICRSrf0_0),.din(w_dff_A_hIFWfd6U2_0),.clk(gclk));
	jdff dff_A_WBICRSrf0_0(.dout(w_dff_A_MlfVKyUe7_0),.din(w_dff_A_WBICRSrf0_0),.clk(gclk));
	jdff dff_A_MlfVKyUe7_0(.dout(w_dff_A_O1RgAoCZ5_0),.din(w_dff_A_MlfVKyUe7_0),.clk(gclk));
	jdff dff_A_O1RgAoCZ5_0(.dout(w_dff_A_9t05lWiJ1_0),.din(w_dff_A_O1RgAoCZ5_0),.clk(gclk));
	jdff dff_A_9t05lWiJ1_0(.dout(w_dff_A_8e3Ab73a8_0),.din(w_dff_A_9t05lWiJ1_0),.clk(gclk));
	jdff dff_A_8e3Ab73a8_0(.dout(w_dff_A_IOr5R2l06_0),.din(w_dff_A_8e3Ab73a8_0),.clk(gclk));
	jdff dff_A_IOr5R2l06_0(.dout(w_dff_A_OhjlDZ687_0),.din(w_dff_A_IOr5R2l06_0),.clk(gclk));
	jdff dff_A_OhjlDZ687_0(.dout(w_dff_A_PVC1HXKf8_0),.din(w_dff_A_OhjlDZ687_0),.clk(gclk));
	jdff dff_A_PVC1HXKf8_0(.dout(w_dff_A_BhGFb2IV8_0),.din(w_dff_A_PVC1HXKf8_0),.clk(gclk));
	jdff dff_A_BhGFb2IV8_0(.dout(w_dff_A_BeLrqKEh3_0),.din(w_dff_A_BhGFb2IV8_0),.clk(gclk));
	jdff dff_A_BeLrqKEh3_0(.dout(w_dff_A_3DQjD6g93_0),.din(w_dff_A_BeLrqKEh3_0),.clk(gclk));
	jdff dff_A_3DQjD6g93_0(.dout(w_dff_A_9Uq65EFi0_0),.din(w_dff_A_3DQjD6g93_0),.clk(gclk));
	jdff dff_A_9Uq65EFi0_0(.dout(w_dff_A_AniK33Dp4_0),.din(w_dff_A_9Uq65EFi0_0),.clk(gclk));
	jdff dff_A_AniK33Dp4_0(.dout(w_dff_A_gJN29yv56_0),.din(w_dff_A_AniK33Dp4_0),.clk(gclk));
	jdff dff_A_gJN29yv56_0(.dout(G286),.din(w_dff_A_gJN29yv56_0),.clk(gclk));
	jdff dff_A_2ffOjGSw0_2(.dout(w_dff_A_lZwHf6R40_0),.din(w_dff_A_2ffOjGSw0_2),.clk(gclk));
	jdff dff_A_lZwHf6R40_0(.dout(w_dff_A_y4g9cm1v4_0),.din(w_dff_A_lZwHf6R40_0),.clk(gclk));
	jdff dff_A_y4g9cm1v4_0(.dout(w_dff_A_pvsCAZDH1_0),.din(w_dff_A_y4g9cm1v4_0),.clk(gclk));
	jdff dff_A_pvsCAZDH1_0(.dout(w_dff_A_SBvcXEsb3_0),.din(w_dff_A_pvsCAZDH1_0),.clk(gclk));
	jdff dff_A_SBvcXEsb3_0(.dout(w_dff_A_KeUUZKkh9_0),.din(w_dff_A_SBvcXEsb3_0),.clk(gclk));
	jdff dff_A_KeUUZKkh9_0(.dout(w_dff_A_D0XsJf9x0_0),.din(w_dff_A_KeUUZKkh9_0),.clk(gclk));
	jdff dff_A_D0XsJf9x0_0(.dout(w_dff_A_LO9zKj3B5_0),.din(w_dff_A_D0XsJf9x0_0),.clk(gclk));
	jdff dff_A_LO9zKj3B5_0(.dout(w_dff_A_RsJhGyoV5_0),.din(w_dff_A_LO9zKj3B5_0),.clk(gclk));
	jdff dff_A_RsJhGyoV5_0(.dout(w_dff_A_9DeQYJjo2_0),.din(w_dff_A_RsJhGyoV5_0),.clk(gclk));
	jdff dff_A_9DeQYJjo2_0(.dout(w_dff_A_B2c7gVPS9_0),.din(w_dff_A_9DeQYJjo2_0),.clk(gclk));
	jdff dff_A_B2c7gVPS9_0(.dout(w_dff_A_UrI4DLaB7_0),.din(w_dff_A_B2c7gVPS9_0),.clk(gclk));
	jdff dff_A_UrI4DLaB7_0(.dout(w_dff_A_Z5WxMyim5_0),.din(w_dff_A_UrI4DLaB7_0),.clk(gclk));
	jdff dff_A_Z5WxMyim5_0(.dout(w_dff_A_zQC6m5t67_0),.din(w_dff_A_Z5WxMyim5_0),.clk(gclk));
	jdff dff_A_zQC6m5t67_0(.dout(w_dff_A_fgLj68N53_0),.din(w_dff_A_zQC6m5t67_0),.clk(gclk));
	jdff dff_A_fgLj68N53_0(.dout(w_dff_A_qbGJPf7C7_0),.din(w_dff_A_fgLj68N53_0),.clk(gclk));
	jdff dff_A_qbGJPf7C7_0(.dout(w_dff_A_SpMBQ90i0_0),.din(w_dff_A_qbGJPf7C7_0),.clk(gclk));
	jdff dff_A_SpMBQ90i0_0(.dout(w_dff_A_w6PG7JqV9_0),.din(w_dff_A_SpMBQ90i0_0),.clk(gclk));
	jdff dff_A_w6PG7JqV9_0(.dout(w_dff_A_rUAgz0BP6_0),.din(w_dff_A_w6PG7JqV9_0),.clk(gclk));
	jdff dff_A_rUAgz0BP6_0(.dout(w_dff_A_lTS3vKVH0_0),.din(w_dff_A_rUAgz0BP6_0),.clk(gclk));
	jdff dff_A_lTS3vKVH0_0(.dout(w_dff_A_A5gke3At5_0),.din(w_dff_A_lTS3vKVH0_0),.clk(gclk));
	jdff dff_A_A5gke3At5_0(.dout(w_dff_A_ZtR7t5VX8_0),.din(w_dff_A_A5gke3At5_0),.clk(gclk));
	jdff dff_A_ZtR7t5VX8_0(.dout(w_dff_A_ZDWOUPiC8_0),.din(w_dff_A_ZtR7t5VX8_0),.clk(gclk));
	jdff dff_A_ZDWOUPiC8_0(.dout(w_dff_A_hoafLdX80_0),.din(w_dff_A_ZDWOUPiC8_0),.clk(gclk));
	jdff dff_A_hoafLdX80_0(.dout(w_dff_A_5racRmi43_0),.din(w_dff_A_hoafLdX80_0),.clk(gclk));
	jdff dff_A_5racRmi43_0(.dout(w_dff_A_ijAeR4rh3_0),.din(w_dff_A_5racRmi43_0),.clk(gclk));
	jdff dff_A_ijAeR4rh3_0(.dout(w_dff_A_ImcgR7xm9_0),.din(w_dff_A_ijAeR4rh3_0),.clk(gclk));
	jdff dff_A_ImcgR7xm9_0(.dout(w_dff_A_Sd58F3UK2_0),.din(w_dff_A_ImcgR7xm9_0),.clk(gclk));
	jdff dff_A_Sd58F3UK2_0(.dout(w_dff_A_cQ8qT2dE3_0),.din(w_dff_A_Sd58F3UK2_0),.clk(gclk));
	jdff dff_A_cQ8qT2dE3_0(.dout(w_dff_A_G3kR2pin3_0),.din(w_dff_A_cQ8qT2dE3_0),.clk(gclk));
	jdff dff_A_G3kR2pin3_0(.dout(w_dff_A_E4NHioB47_0),.din(w_dff_A_G3kR2pin3_0),.clk(gclk));
	jdff dff_A_E4NHioB47_0(.dout(w_dff_A_CptaiCnM7_0),.din(w_dff_A_E4NHioB47_0),.clk(gclk));
	jdff dff_A_CptaiCnM7_0(.dout(w_dff_A_9TQb8tTY9_0),.din(w_dff_A_CptaiCnM7_0),.clk(gclk));
	jdff dff_A_9TQb8tTY9_0(.dout(w_dff_A_tyy4Ebdq7_0),.din(w_dff_A_9TQb8tTY9_0),.clk(gclk));
	jdff dff_A_tyy4Ebdq7_0(.dout(w_dff_A_xxyNTzB67_0),.din(w_dff_A_tyy4Ebdq7_0),.clk(gclk));
	jdff dff_A_xxyNTzB67_0(.dout(w_dff_A_BJDi9gcw9_0),.din(w_dff_A_xxyNTzB67_0),.clk(gclk));
	jdff dff_A_BJDi9gcw9_0(.dout(w_dff_A_I9mtoSGP1_0),.din(w_dff_A_BJDi9gcw9_0),.clk(gclk));
	jdff dff_A_I9mtoSGP1_0(.dout(G289),.din(w_dff_A_I9mtoSGP1_0),.clk(gclk));
	jdff dff_A_5CWJDb799_2(.dout(w_dff_A_gBIXloda6_0),.din(w_dff_A_5CWJDb799_2),.clk(gclk));
	jdff dff_A_gBIXloda6_0(.dout(w_dff_A_lmqIViUF0_0),.din(w_dff_A_gBIXloda6_0),.clk(gclk));
	jdff dff_A_lmqIViUF0_0(.dout(w_dff_A_JSXejjHQ0_0),.din(w_dff_A_lmqIViUF0_0),.clk(gclk));
	jdff dff_A_JSXejjHQ0_0(.dout(w_dff_A_d7GRBcPd6_0),.din(w_dff_A_JSXejjHQ0_0),.clk(gclk));
	jdff dff_A_d7GRBcPd6_0(.dout(w_dff_A_lHw19Lfd9_0),.din(w_dff_A_d7GRBcPd6_0),.clk(gclk));
	jdff dff_A_lHw19Lfd9_0(.dout(w_dff_A_1enBGeNJ6_0),.din(w_dff_A_lHw19Lfd9_0),.clk(gclk));
	jdff dff_A_1enBGeNJ6_0(.dout(w_dff_A_T9eJqdRv8_0),.din(w_dff_A_1enBGeNJ6_0),.clk(gclk));
	jdff dff_A_T9eJqdRv8_0(.dout(w_dff_A_RvoX3PVw5_0),.din(w_dff_A_T9eJqdRv8_0),.clk(gclk));
	jdff dff_A_RvoX3PVw5_0(.dout(w_dff_A_sAWPyZ7B9_0),.din(w_dff_A_RvoX3PVw5_0),.clk(gclk));
	jdff dff_A_sAWPyZ7B9_0(.dout(w_dff_A_6bQx5k2h2_0),.din(w_dff_A_sAWPyZ7B9_0),.clk(gclk));
	jdff dff_A_6bQx5k2h2_0(.dout(w_dff_A_MIMuAJRc2_0),.din(w_dff_A_6bQx5k2h2_0),.clk(gclk));
	jdff dff_A_MIMuAJRc2_0(.dout(w_dff_A_G7bHtZWK7_0),.din(w_dff_A_MIMuAJRc2_0),.clk(gclk));
	jdff dff_A_G7bHtZWK7_0(.dout(w_dff_A_VI3Fp35F9_0),.din(w_dff_A_G7bHtZWK7_0),.clk(gclk));
	jdff dff_A_VI3Fp35F9_0(.dout(w_dff_A_bk9s3Rj58_0),.din(w_dff_A_VI3Fp35F9_0),.clk(gclk));
	jdff dff_A_bk9s3Rj58_0(.dout(w_dff_A_JWuAjjag5_0),.din(w_dff_A_bk9s3Rj58_0),.clk(gclk));
	jdff dff_A_JWuAjjag5_0(.dout(w_dff_A_TXvXQldr2_0),.din(w_dff_A_JWuAjjag5_0),.clk(gclk));
	jdff dff_A_TXvXQldr2_0(.dout(w_dff_A_fwdvcNeG0_0),.din(w_dff_A_TXvXQldr2_0),.clk(gclk));
	jdff dff_A_fwdvcNeG0_0(.dout(w_dff_A_yAH4vpjM2_0),.din(w_dff_A_fwdvcNeG0_0),.clk(gclk));
	jdff dff_A_yAH4vpjM2_0(.dout(w_dff_A_wMQptCx18_0),.din(w_dff_A_yAH4vpjM2_0),.clk(gclk));
	jdff dff_A_wMQptCx18_0(.dout(w_dff_A_amkVk9Oq1_0),.din(w_dff_A_wMQptCx18_0),.clk(gclk));
	jdff dff_A_amkVk9Oq1_0(.dout(w_dff_A_j40ug4rP7_0),.din(w_dff_A_amkVk9Oq1_0),.clk(gclk));
	jdff dff_A_j40ug4rP7_0(.dout(w_dff_A_MBybOkkQ0_0),.din(w_dff_A_j40ug4rP7_0),.clk(gclk));
	jdff dff_A_MBybOkkQ0_0(.dout(w_dff_A_v7DppBZp6_0),.din(w_dff_A_MBybOkkQ0_0),.clk(gclk));
	jdff dff_A_v7DppBZp6_0(.dout(w_dff_A_Zb9ekEIH1_0),.din(w_dff_A_v7DppBZp6_0),.clk(gclk));
	jdff dff_A_Zb9ekEIH1_0(.dout(w_dff_A_v48GulAq7_0),.din(w_dff_A_Zb9ekEIH1_0),.clk(gclk));
	jdff dff_A_v48GulAq7_0(.dout(w_dff_A_vteSKWGg3_0),.din(w_dff_A_v48GulAq7_0),.clk(gclk));
	jdff dff_A_vteSKWGg3_0(.dout(w_dff_A_TTWLxi272_0),.din(w_dff_A_vteSKWGg3_0),.clk(gclk));
	jdff dff_A_TTWLxi272_0(.dout(w_dff_A_wRXPZGqq9_0),.din(w_dff_A_TTWLxi272_0),.clk(gclk));
	jdff dff_A_wRXPZGqq9_0(.dout(w_dff_A_hYG6VFTD3_0),.din(w_dff_A_wRXPZGqq9_0),.clk(gclk));
	jdff dff_A_hYG6VFTD3_0(.dout(w_dff_A_6UpMiI3Z2_0),.din(w_dff_A_hYG6VFTD3_0),.clk(gclk));
	jdff dff_A_6UpMiI3Z2_0(.dout(w_dff_A_pCuZM0lV5_0),.din(w_dff_A_6UpMiI3Z2_0),.clk(gclk));
	jdff dff_A_pCuZM0lV5_0(.dout(w_dff_A_rKqX1lhP6_0),.din(w_dff_A_pCuZM0lV5_0),.clk(gclk));
	jdff dff_A_rKqX1lhP6_0(.dout(w_dff_A_4scZZCVe2_0),.din(w_dff_A_rKqX1lhP6_0),.clk(gclk));
	jdff dff_A_4scZZCVe2_0(.dout(w_dff_A_KuyJyPJT5_0),.din(w_dff_A_4scZZCVe2_0),.clk(gclk));
	jdff dff_A_KuyJyPJT5_0(.dout(w_dff_A_NYKCgtdD7_0),.din(w_dff_A_KuyJyPJT5_0),.clk(gclk));
	jdff dff_A_NYKCgtdD7_0(.dout(G292),.din(w_dff_A_NYKCgtdD7_0),.clk(gclk));
	jdff dff_A_5UJxVmwi0_1(.dout(w_dff_A_b2XBNgqA6_0),.din(w_dff_A_5UJxVmwi0_1),.clk(gclk));
	jdff dff_A_b2XBNgqA6_0(.dout(w_dff_A_eEgdHU7Q1_0),.din(w_dff_A_b2XBNgqA6_0),.clk(gclk));
	jdff dff_A_eEgdHU7Q1_0(.dout(w_dff_A_OPwWvTME9_0),.din(w_dff_A_eEgdHU7Q1_0),.clk(gclk));
	jdff dff_A_OPwWvTME9_0(.dout(w_dff_A_XxpWVlXX4_0),.din(w_dff_A_OPwWvTME9_0),.clk(gclk));
	jdff dff_A_XxpWVlXX4_0(.dout(w_dff_A_M4ISSJIz9_0),.din(w_dff_A_XxpWVlXX4_0),.clk(gclk));
	jdff dff_A_M4ISSJIz9_0(.dout(w_dff_A_sR6jGFbd4_0),.din(w_dff_A_M4ISSJIz9_0),.clk(gclk));
	jdff dff_A_sR6jGFbd4_0(.dout(w_dff_A_F7t6vG9k5_0),.din(w_dff_A_sR6jGFbd4_0),.clk(gclk));
	jdff dff_A_F7t6vG9k5_0(.dout(w_dff_A_YTEGXAvm4_0),.din(w_dff_A_F7t6vG9k5_0),.clk(gclk));
	jdff dff_A_YTEGXAvm4_0(.dout(w_dff_A_qluAPOsF2_0),.din(w_dff_A_YTEGXAvm4_0),.clk(gclk));
	jdff dff_A_qluAPOsF2_0(.dout(w_dff_A_HA1Jo9N09_0),.din(w_dff_A_qluAPOsF2_0),.clk(gclk));
	jdff dff_A_HA1Jo9N09_0(.dout(w_dff_A_R1xys3UN0_0),.din(w_dff_A_HA1Jo9N09_0),.clk(gclk));
	jdff dff_A_R1xys3UN0_0(.dout(w_dff_A_YuGT2vLL5_0),.din(w_dff_A_R1xys3UN0_0),.clk(gclk));
	jdff dff_A_YuGT2vLL5_0(.dout(w_dff_A_yhE1oluh6_0),.din(w_dff_A_YuGT2vLL5_0),.clk(gclk));
	jdff dff_A_yhE1oluh6_0(.dout(w_dff_A_57palikL4_0),.din(w_dff_A_yhE1oluh6_0),.clk(gclk));
	jdff dff_A_57palikL4_0(.dout(w_dff_A_nRMANwxx1_0),.din(w_dff_A_57palikL4_0),.clk(gclk));
	jdff dff_A_nRMANwxx1_0(.dout(w_dff_A_Ci6ruBFk3_0),.din(w_dff_A_nRMANwxx1_0),.clk(gclk));
	jdff dff_A_Ci6ruBFk3_0(.dout(w_dff_A_wI9VE5U23_0),.din(w_dff_A_Ci6ruBFk3_0),.clk(gclk));
	jdff dff_A_wI9VE5U23_0(.dout(w_dff_A_UOulhVea0_0),.din(w_dff_A_wI9VE5U23_0),.clk(gclk));
	jdff dff_A_UOulhVea0_0(.dout(w_dff_A_KfzX7r6E1_0),.din(w_dff_A_UOulhVea0_0),.clk(gclk));
	jdff dff_A_KfzX7r6E1_0(.dout(w_dff_A_zitRS7j84_0),.din(w_dff_A_KfzX7r6E1_0),.clk(gclk));
	jdff dff_A_zitRS7j84_0(.dout(w_dff_A_m58o1jfZ3_0),.din(w_dff_A_zitRS7j84_0),.clk(gclk));
	jdff dff_A_m58o1jfZ3_0(.dout(w_dff_A_oTpXEnrE9_0),.din(w_dff_A_m58o1jfZ3_0),.clk(gclk));
	jdff dff_A_oTpXEnrE9_0(.dout(w_dff_A_ve2dmMk57_0),.din(w_dff_A_oTpXEnrE9_0),.clk(gclk));
	jdff dff_A_ve2dmMk57_0(.dout(w_dff_A_CFovSXlD4_0),.din(w_dff_A_ve2dmMk57_0),.clk(gclk));
	jdff dff_A_CFovSXlD4_0(.dout(w_dff_A_63Jd9I6I5_0),.din(w_dff_A_CFovSXlD4_0),.clk(gclk));
	jdff dff_A_63Jd9I6I5_0(.dout(w_dff_A_72UBYXcW8_0),.din(w_dff_A_63Jd9I6I5_0),.clk(gclk));
	jdff dff_A_72UBYXcW8_0(.dout(w_dff_A_VMcvQswL1_0),.din(w_dff_A_72UBYXcW8_0),.clk(gclk));
	jdff dff_A_VMcvQswL1_0(.dout(w_dff_A_gIB7J3tz4_0),.din(w_dff_A_VMcvQswL1_0),.clk(gclk));
	jdff dff_A_gIB7J3tz4_0(.dout(w_dff_A_pUXQxgje3_0),.din(w_dff_A_gIB7J3tz4_0),.clk(gclk));
	jdff dff_A_pUXQxgje3_0(.dout(w_dff_A_aVMdw0M67_0),.din(w_dff_A_pUXQxgje3_0),.clk(gclk));
	jdff dff_A_aVMdw0M67_0(.dout(w_dff_A_rYW2m9Lx6_0),.din(w_dff_A_aVMdw0M67_0),.clk(gclk));
	jdff dff_A_rYW2m9Lx6_0(.dout(w_dff_A_5SGfGcPQ0_0),.din(w_dff_A_rYW2m9Lx6_0),.clk(gclk));
	jdff dff_A_5SGfGcPQ0_0(.dout(w_dff_A_Brk5I6Kr5_0),.din(w_dff_A_5SGfGcPQ0_0),.clk(gclk));
	jdff dff_A_Brk5I6Kr5_0(.dout(w_dff_A_cChG1fMn0_0),.din(w_dff_A_Brk5I6Kr5_0),.clk(gclk));
	jdff dff_A_cChG1fMn0_0(.dout(w_dff_A_z1L8L5Ah3_0),.din(w_dff_A_cChG1fMn0_0),.clk(gclk));
	jdff dff_A_z1L8L5Ah3_0(.dout(w_dff_A_THGPqgYF5_0),.din(w_dff_A_z1L8L5Ah3_0),.clk(gclk));
	jdff dff_A_THGPqgYF5_0(.dout(w_dff_A_UkS5GTox6_0),.din(w_dff_A_THGPqgYF5_0),.clk(gclk));
	jdff dff_A_UkS5GTox6_0(.dout(G341),.din(w_dff_A_UkS5GTox6_0),.clk(gclk));
	jdff dff_A_LYTWwnQT3_2(.dout(w_dff_A_rOhaXiQu9_0),.din(w_dff_A_LYTWwnQT3_2),.clk(gclk));
	jdff dff_A_rOhaXiQu9_0(.dout(w_dff_A_qSnjebqh5_0),.din(w_dff_A_rOhaXiQu9_0),.clk(gclk));
	jdff dff_A_qSnjebqh5_0(.dout(w_dff_A_axO0PiAe0_0),.din(w_dff_A_qSnjebqh5_0),.clk(gclk));
	jdff dff_A_axO0PiAe0_0(.dout(w_dff_A_qag10fA49_0),.din(w_dff_A_axO0PiAe0_0),.clk(gclk));
	jdff dff_A_qag10fA49_0(.dout(w_dff_A_Jfcy6ivk8_0),.din(w_dff_A_qag10fA49_0),.clk(gclk));
	jdff dff_A_Jfcy6ivk8_0(.dout(w_dff_A_e9npHuAR1_0),.din(w_dff_A_Jfcy6ivk8_0),.clk(gclk));
	jdff dff_A_e9npHuAR1_0(.dout(w_dff_A_M4OBSOlH5_0),.din(w_dff_A_e9npHuAR1_0),.clk(gclk));
	jdff dff_A_M4OBSOlH5_0(.dout(w_dff_A_sp0YFyoC1_0),.din(w_dff_A_M4OBSOlH5_0),.clk(gclk));
	jdff dff_A_sp0YFyoC1_0(.dout(w_dff_A_npVOn1jy5_0),.din(w_dff_A_sp0YFyoC1_0),.clk(gclk));
	jdff dff_A_npVOn1jy5_0(.dout(w_dff_A_RzB7xMFP5_0),.din(w_dff_A_npVOn1jy5_0),.clk(gclk));
	jdff dff_A_RzB7xMFP5_0(.dout(w_dff_A_kS9mjGrh5_0),.din(w_dff_A_RzB7xMFP5_0),.clk(gclk));
	jdff dff_A_kS9mjGrh5_0(.dout(w_dff_A_UWfax2q97_0),.din(w_dff_A_kS9mjGrh5_0),.clk(gclk));
	jdff dff_A_UWfax2q97_0(.dout(w_dff_A_PZlZX5CP8_0),.din(w_dff_A_UWfax2q97_0),.clk(gclk));
	jdff dff_A_PZlZX5CP8_0(.dout(w_dff_A_6k2aV4Wv5_0),.din(w_dff_A_PZlZX5CP8_0),.clk(gclk));
	jdff dff_A_6k2aV4Wv5_0(.dout(w_dff_A_x7H4R5ju3_0),.din(w_dff_A_6k2aV4Wv5_0),.clk(gclk));
	jdff dff_A_x7H4R5ju3_0(.dout(w_dff_A_JWp8zvp55_0),.din(w_dff_A_x7H4R5ju3_0),.clk(gclk));
	jdff dff_A_JWp8zvp55_0(.dout(w_dff_A_U4U6aH6s4_0),.din(w_dff_A_JWp8zvp55_0),.clk(gclk));
	jdff dff_A_U4U6aH6s4_0(.dout(w_dff_A_4ZuLP4ev6_0),.din(w_dff_A_U4U6aH6s4_0),.clk(gclk));
	jdff dff_A_4ZuLP4ev6_0(.dout(w_dff_A_1OYAlXSC9_0),.din(w_dff_A_4ZuLP4ev6_0),.clk(gclk));
	jdff dff_A_1OYAlXSC9_0(.dout(w_dff_A_7RyYZd4j5_0),.din(w_dff_A_1OYAlXSC9_0),.clk(gclk));
	jdff dff_A_7RyYZd4j5_0(.dout(w_dff_A_7CBFCoj75_0),.din(w_dff_A_7RyYZd4j5_0),.clk(gclk));
	jdff dff_A_7CBFCoj75_0(.dout(w_dff_A_xtSKDinO3_0),.din(w_dff_A_7CBFCoj75_0),.clk(gclk));
	jdff dff_A_xtSKDinO3_0(.dout(w_dff_A_YBmOpkG23_0),.din(w_dff_A_xtSKDinO3_0),.clk(gclk));
	jdff dff_A_YBmOpkG23_0(.dout(w_dff_A_njEXYHq94_0),.din(w_dff_A_YBmOpkG23_0),.clk(gclk));
	jdff dff_A_njEXYHq94_0(.dout(w_dff_A_l9zCHjn00_0),.din(w_dff_A_njEXYHq94_0),.clk(gclk));
	jdff dff_A_l9zCHjn00_0(.dout(w_dff_A_y6mXuzjy1_0),.din(w_dff_A_l9zCHjn00_0),.clk(gclk));
	jdff dff_A_y6mXuzjy1_0(.dout(w_dff_A_SqhIIYuN3_0),.din(w_dff_A_y6mXuzjy1_0),.clk(gclk));
	jdff dff_A_SqhIIYuN3_0(.dout(w_dff_A_Fy68E4ri0_0),.din(w_dff_A_SqhIIYuN3_0),.clk(gclk));
	jdff dff_A_Fy68E4ri0_0(.dout(w_dff_A_MMhPxFZC5_0),.din(w_dff_A_Fy68E4ri0_0),.clk(gclk));
	jdff dff_A_MMhPxFZC5_0(.dout(w_dff_A_5ICq8oAh5_0),.din(w_dff_A_MMhPxFZC5_0),.clk(gclk));
	jdff dff_A_5ICq8oAh5_0(.dout(w_dff_A_cSWnvPqz8_0),.din(w_dff_A_5ICq8oAh5_0),.clk(gclk));
	jdff dff_A_cSWnvPqz8_0(.dout(w_dff_A_tTnXYDlF1_0),.din(w_dff_A_cSWnvPqz8_0),.clk(gclk));
	jdff dff_A_tTnXYDlF1_0(.dout(w_dff_A_AxbIMWhd7_0),.din(w_dff_A_tTnXYDlF1_0),.clk(gclk));
	jdff dff_A_AxbIMWhd7_0(.dout(w_dff_A_JtGuUzYo4_0),.din(w_dff_A_AxbIMWhd7_0),.clk(gclk));
	jdff dff_A_JtGuUzYo4_0(.dout(w_dff_A_XXnkcJya1_0),.din(w_dff_A_JtGuUzYo4_0),.clk(gclk));
	jdff dff_A_XXnkcJya1_0(.dout(G281),.din(w_dff_A_XXnkcJya1_0),.clk(gclk));
	jdff dff_A_v6D1FION8_1(.dout(w_dff_A_WXnqrcDo0_0),.din(w_dff_A_v6D1FION8_1),.clk(gclk));
	jdff dff_A_WXnqrcDo0_0(.dout(w_dff_A_h4wWoAuY3_0),.din(w_dff_A_WXnqrcDo0_0),.clk(gclk));
	jdff dff_A_h4wWoAuY3_0(.dout(w_dff_A_J2Y6GuVK3_0),.din(w_dff_A_h4wWoAuY3_0),.clk(gclk));
	jdff dff_A_J2Y6GuVK3_0(.dout(w_dff_A_GrZzI1TX9_0),.din(w_dff_A_J2Y6GuVK3_0),.clk(gclk));
	jdff dff_A_GrZzI1TX9_0(.dout(w_dff_A_oAmrXrWR6_0),.din(w_dff_A_GrZzI1TX9_0),.clk(gclk));
	jdff dff_A_oAmrXrWR6_0(.dout(w_dff_A_vz6SqLEs1_0),.din(w_dff_A_oAmrXrWR6_0),.clk(gclk));
	jdff dff_A_vz6SqLEs1_0(.dout(w_dff_A_riF2gTTT2_0),.din(w_dff_A_vz6SqLEs1_0),.clk(gclk));
	jdff dff_A_riF2gTTT2_0(.dout(w_dff_A_txUkHtJJ7_0),.din(w_dff_A_riF2gTTT2_0),.clk(gclk));
	jdff dff_A_txUkHtJJ7_0(.dout(w_dff_A_tfPqtxZD4_0),.din(w_dff_A_txUkHtJJ7_0),.clk(gclk));
	jdff dff_A_tfPqtxZD4_0(.dout(w_dff_A_GqLnxeAP1_0),.din(w_dff_A_tfPqtxZD4_0),.clk(gclk));
	jdff dff_A_GqLnxeAP1_0(.dout(w_dff_A_a3qliUqZ3_0),.din(w_dff_A_GqLnxeAP1_0),.clk(gclk));
	jdff dff_A_a3qliUqZ3_0(.dout(w_dff_A_YsXibD2e5_0),.din(w_dff_A_a3qliUqZ3_0),.clk(gclk));
	jdff dff_A_YsXibD2e5_0(.dout(w_dff_A_jxRaui4Z3_0),.din(w_dff_A_YsXibD2e5_0),.clk(gclk));
	jdff dff_A_jxRaui4Z3_0(.dout(w_dff_A_UXIeOfXk5_0),.din(w_dff_A_jxRaui4Z3_0),.clk(gclk));
	jdff dff_A_UXIeOfXk5_0(.dout(w_dff_A_QXgHYmff0_0),.din(w_dff_A_UXIeOfXk5_0),.clk(gclk));
	jdff dff_A_QXgHYmff0_0(.dout(w_dff_A_HchAHDuA6_0),.din(w_dff_A_QXgHYmff0_0),.clk(gclk));
	jdff dff_A_HchAHDuA6_0(.dout(w_dff_A_FiyQ8NZB0_0),.din(w_dff_A_HchAHDuA6_0),.clk(gclk));
	jdff dff_A_FiyQ8NZB0_0(.dout(w_dff_A_85hrb3iP2_0),.din(w_dff_A_FiyQ8NZB0_0),.clk(gclk));
	jdff dff_A_85hrb3iP2_0(.dout(w_dff_A_9tsud5Bl6_0),.din(w_dff_A_85hrb3iP2_0),.clk(gclk));
	jdff dff_A_9tsud5Bl6_0(.dout(w_dff_A_wZehHiKb2_0),.din(w_dff_A_9tsud5Bl6_0),.clk(gclk));
	jdff dff_A_wZehHiKb2_0(.dout(w_dff_A_1Oqsl1bb5_0),.din(w_dff_A_wZehHiKb2_0),.clk(gclk));
	jdff dff_A_1Oqsl1bb5_0(.dout(w_dff_A_oflB3tYa7_0),.din(w_dff_A_1Oqsl1bb5_0),.clk(gclk));
	jdff dff_A_oflB3tYa7_0(.dout(w_dff_A_asaIc2GR5_0),.din(w_dff_A_oflB3tYa7_0),.clk(gclk));
	jdff dff_A_asaIc2GR5_0(.dout(w_dff_A_6tFU48pa8_0),.din(w_dff_A_asaIc2GR5_0),.clk(gclk));
	jdff dff_A_6tFU48pa8_0(.dout(w_dff_A_A77uKbXu1_0),.din(w_dff_A_6tFU48pa8_0),.clk(gclk));
	jdff dff_A_A77uKbXu1_0(.dout(w_dff_A_uplEs2uz3_0),.din(w_dff_A_A77uKbXu1_0),.clk(gclk));
	jdff dff_A_uplEs2uz3_0(.dout(w_dff_A_l7IEkgS81_0),.din(w_dff_A_uplEs2uz3_0),.clk(gclk));
	jdff dff_A_l7IEkgS81_0(.dout(w_dff_A_HHM2aAnN1_0),.din(w_dff_A_l7IEkgS81_0),.clk(gclk));
	jdff dff_A_HHM2aAnN1_0(.dout(w_dff_A_K3LEQtDj6_0),.din(w_dff_A_HHM2aAnN1_0),.clk(gclk));
	jdff dff_A_K3LEQtDj6_0(.dout(w_dff_A_bk1vyzJA0_0),.din(w_dff_A_K3LEQtDj6_0),.clk(gclk));
	jdff dff_A_bk1vyzJA0_0(.dout(w_dff_A_ZthzvxHl9_0),.din(w_dff_A_bk1vyzJA0_0),.clk(gclk));
	jdff dff_A_ZthzvxHl9_0(.dout(w_dff_A_pIUJ1OB06_0),.din(w_dff_A_ZthzvxHl9_0),.clk(gclk));
	jdff dff_A_pIUJ1OB06_0(.dout(w_dff_A_5zKAxaVt0_0),.din(w_dff_A_pIUJ1OB06_0),.clk(gclk));
	jdff dff_A_5zKAxaVt0_0(.dout(w_dff_A_1OuSgU3z5_0),.din(w_dff_A_5zKAxaVt0_0),.clk(gclk));
	jdff dff_A_1OuSgU3z5_0(.dout(w_dff_A_FD6u7nH66_0),.din(w_dff_A_1OuSgU3z5_0),.clk(gclk));
	jdff dff_A_FD6u7nH66_0(.dout(w_dff_A_VmfczGuC8_0),.din(w_dff_A_FD6u7nH66_0),.clk(gclk));
	jdff dff_A_VmfczGuC8_0(.dout(w_dff_A_6j1uDAKw2_0),.din(w_dff_A_VmfczGuC8_0),.clk(gclk));
	jdff dff_A_6j1uDAKw2_0(.dout(w_dff_A_yULD7g5r5_0),.din(w_dff_A_6j1uDAKw2_0),.clk(gclk));
	jdff dff_A_yULD7g5r5_0(.dout(G453),.din(w_dff_A_yULD7g5r5_0),.clk(gclk));
	jdff dff_A_6JNnbqa23_2(.dout(w_dff_A_TgSBmCTr9_0),.din(w_dff_A_6JNnbqa23_2),.clk(gclk));
	jdff dff_A_TgSBmCTr9_0(.dout(w_dff_A_nsEkwB1u2_0),.din(w_dff_A_TgSBmCTr9_0),.clk(gclk));
	jdff dff_A_nsEkwB1u2_0(.dout(w_dff_A_xENo23u41_0),.din(w_dff_A_nsEkwB1u2_0),.clk(gclk));
	jdff dff_A_xENo23u41_0(.dout(w_dff_A_J1Wq44AT9_0),.din(w_dff_A_xENo23u41_0),.clk(gclk));
	jdff dff_A_J1Wq44AT9_0(.dout(w_dff_A_WwNDomRU8_0),.din(w_dff_A_J1Wq44AT9_0),.clk(gclk));
	jdff dff_A_WwNDomRU8_0(.dout(w_dff_A_MZuE6uKN3_0),.din(w_dff_A_WwNDomRU8_0),.clk(gclk));
	jdff dff_A_MZuE6uKN3_0(.dout(w_dff_A_uDcMwWqz3_0),.din(w_dff_A_MZuE6uKN3_0),.clk(gclk));
	jdff dff_A_uDcMwWqz3_0(.dout(w_dff_A_jnpnw1D61_0),.din(w_dff_A_uDcMwWqz3_0),.clk(gclk));
	jdff dff_A_jnpnw1D61_0(.dout(w_dff_A_tJ1NdhgQ2_0),.din(w_dff_A_jnpnw1D61_0),.clk(gclk));
	jdff dff_A_tJ1NdhgQ2_0(.dout(w_dff_A_iyNZ2jFh6_0),.din(w_dff_A_tJ1NdhgQ2_0),.clk(gclk));
	jdff dff_A_iyNZ2jFh6_0(.dout(w_dff_A_lbjLwgey2_0),.din(w_dff_A_iyNZ2jFh6_0),.clk(gclk));
	jdff dff_A_lbjLwgey2_0(.dout(w_dff_A_UMBV82v74_0),.din(w_dff_A_lbjLwgey2_0),.clk(gclk));
	jdff dff_A_UMBV82v74_0(.dout(w_dff_A_mboFH9Xs4_0),.din(w_dff_A_UMBV82v74_0),.clk(gclk));
	jdff dff_A_mboFH9Xs4_0(.dout(w_dff_A_NU65Fn1J5_0),.din(w_dff_A_mboFH9Xs4_0),.clk(gclk));
	jdff dff_A_NU65Fn1J5_0(.dout(w_dff_A_evzEM4tN1_0),.din(w_dff_A_NU65Fn1J5_0),.clk(gclk));
	jdff dff_A_evzEM4tN1_0(.dout(w_dff_A_UbO1NeX40_0),.din(w_dff_A_evzEM4tN1_0),.clk(gclk));
	jdff dff_A_UbO1NeX40_0(.dout(w_dff_A_UmRaH5YV2_0),.din(w_dff_A_UbO1NeX40_0),.clk(gclk));
	jdff dff_A_UmRaH5YV2_0(.dout(w_dff_A_njncPKZm2_0),.din(w_dff_A_UmRaH5YV2_0),.clk(gclk));
	jdff dff_A_njncPKZm2_0(.dout(w_dff_A_RcIDBfhq2_0),.din(w_dff_A_njncPKZm2_0),.clk(gclk));
	jdff dff_A_RcIDBfhq2_0(.dout(w_dff_A_64X2WlhV8_0),.din(w_dff_A_RcIDBfhq2_0),.clk(gclk));
	jdff dff_A_64X2WlhV8_0(.dout(w_dff_A_j9qVIGQX3_0),.din(w_dff_A_64X2WlhV8_0),.clk(gclk));
	jdff dff_A_j9qVIGQX3_0(.dout(w_dff_A_y4Cspc1X9_0),.din(w_dff_A_j9qVIGQX3_0),.clk(gclk));
	jdff dff_A_y4Cspc1X9_0(.dout(w_dff_A_bi8BWD2L9_0),.din(w_dff_A_y4Cspc1X9_0),.clk(gclk));
	jdff dff_A_bi8BWD2L9_0(.dout(w_dff_A_tpnaq9my9_0),.din(w_dff_A_bi8BWD2L9_0),.clk(gclk));
	jdff dff_A_tpnaq9my9_0(.dout(w_dff_A_uXa5h7pz6_0),.din(w_dff_A_tpnaq9my9_0),.clk(gclk));
	jdff dff_A_uXa5h7pz6_0(.dout(w_dff_A_byOiI9Mn9_0),.din(w_dff_A_uXa5h7pz6_0),.clk(gclk));
	jdff dff_A_byOiI9Mn9_0(.dout(w_dff_A_rCz93Nd91_0),.din(w_dff_A_byOiI9Mn9_0),.clk(gclk));
	jdff dff_A_rCz93Nd91_0(.dout(w_dff_A_JJJQY4Cb6_0),.din(w_dff_A_rCz93Nd91_0),.clk(gclk));
	jdff dff_A_JJJQY4Cb6_0(.dout(w_dff_A_0LPf6fYh5_0),.din(w_dff_A_JJJQY4Cb6_0),.clk(gclk));
	jdff dff_A_0LPf6fYh5_0(.dout(w_dff_A_hrYBhWcf5_0),.din(w_dff_A_0LPf6fYh5_0),.clk(gclk));
	jdff dff_A_hrYBhWcf5_0(.dout(w_dff_A_qrCIzEHB0_0),.din(w_dff_A_hrYBhWcf5_0),.clk(gclk));
	jdff dff_A_qrCIzEHB0_0(.dout(w_dff_A_uIzUog2C5_0),.din(w_dff_A_qrCIzEHB0_0),.clk(gclk));
	jdff dff_A_uIzUog2C5_0(.dout(w_dff_A_Da6qkFV23_0),.din(w_dff_A_uIzUog2C5_0),.clk(gclk));
	jdff dff_A_Da6qkFV23_0(.dout(w_dff_A_2BUrEj0k5_0),.din(w_dff_A_Da6qkFV23_0),.clk(gclk));
	jdff dff_A_2BUrEj0k5_0(.dout(w_dff_A_75b2Pduh5_0),.din(w_dff_A_2BUrEj0k5_0),.clk(gclk));
	jdff dff_A_75b2Pduh5_0(.dout(w_dff_A_YFaS9lDM2_0),.din(w_dff_A_75b2Pduh5_0),.clk(gclk));
	jdff dff_A_YFaS9lDM2_0(.dout(w_dff_A_nnznEvcV8_0),.din(w_dff_A_YFaS9lDM2_0),.clk(gclk));
	jdff dff_A_nnznEvcV8_0(.dout(G278),.din(w_dff_A_nnznEvcV8_0),.clk(gclk));
	jdff dff_A_JUhLnoel6_2(.dout(w_dff_A_YIPQoqhU6_0),.din(w_dff_A_JUhLnoel6_2),.clk(gclk));
	jdff dff_A_YIPQoqhU6_0(.dout(w_dff_A_xU9CMkso1_0),.din(w_dff_A_YIPQoqhU6_0),.clk(gclk));
	jdff dff_A_xU9CMkso1_0(.dout(w_dff_A_fWTD6whD3_0),.din(w_dff_A_xU9CMkso1_0),.clk(gclk));
	jdff dff_A_fWTD6whD3_0(.dout(w_dff_A_WwJWWjDG7_0),.din(w_dff_A_fWTD6whD3_0),.clk(gclk));
	jdff dff_A_WwJWWjDG7_0(.dout(w_dff_A_WUQ9TBw92_0),.din(w_dff_A_WwJWWjDG7_0),.clk(gclk));
	jdff dff_A_WUQ9TBw92_0(.dout(w_dff_A_Rmjp52Px5_0),.din(w_dff_A_WUQ9TBw92_0),.clk(gclk));
	jdff dff_A_Rmjp52Px5_0(.dout(w_dff_A_7HILhU292_0),.din(w_dff_A_Rmjp52Px5_0),.clk(gclk));
	jdff dff_A_7HILhU292_0(.dout(w_dff_A_pB5TzMQF2_0),.din(w_dff_A_7HILhU292_0),.clk(gclk));
	jdff dff_A_pB5TzMQF2_0(.dout(w_dff_A_5WNYiVIZ8_0),.din(w_dff_A_pB5TzMQF2_0),.clk(gclk));
	jdff dff_A_5WNYiVIZ8_0(.dout(w_dff_A_r269STCO2_0),.din(w_dff_A_5WNYiVIZ8_0),.clk(gclk));
	jdff dff_A_r269STCO2_0(.dout(w_dff_A_t7zpBKCr2_0),.din(w_dff_A_r269STCO2_0),.clk(gclk));
	jdff dff_A_t7zpBKCr2_0(.dout(w_dff_A_c8nFuvde7_0),.din(w_dff_A_t7zpBKCr2_0),.clk(gclk));
	jdff dff_A_c8nFuvde7_0(.dout(w_dff_A_steTrupJ0_0),.din(w_dff_A_c8nFuvde7_0),.clk(gclk));
	jdff dff_A_steTrupJ0_0(.dout(w_dff_A_sHvWjVfY7_0),.din(w_dff_A_steTrupJ0_0),.clk(gclk));
	jdff dff_A_sHvWjVfY7_0(.dout(w_dff_A_3qGhr6OA7_0),.din(w_dff_A_sHvWjVfY7_0),.clk(gclk));
	jdff dff_A_3qGhr6OA7_0(.dout(w_dff_A_L2wcn2YN5_0),.din(w_dff_A_3qGhr6OA7_0),.clk(gclk));
	jdff dff_A_L2wcn2YN5_0(.dout(w_dff_A_S7Ay9VY61_0),.din(w_dff_A_L2wcn2YN5_0),.clk(gclk));
	jdff dff_A_S7Ay9VY61_0(.dout(w_dff_A_HFCc6Y289_0),.din(w_dff_A_S7Ay9VY61_0),.clk(gclk));
	jdff dff_A_HFCc6Y289_0(.dout(w_dff_A_vz9gJvBL0_0),.din(w_dff_A_HFCc6Y289_0),.clk(gclk));
	jdff dff_A_vz9gJvBL0_0(.dout(w_dff_A_OgeEnrSc8_0),.din(w_dff_A_vz9gJvBL0_0),.clk(gclk));
	jdff dff_A_OgeEnrSc8_0(.dout(w_dff_A_DhQvmmJb6_0),.din(w_dff_A_OgeEnrSc8_0),.clk(gclk));
	jdff dff_A_DhQvmmJb6_0(.dout(w_dff_A_yWxvpk0L9_0),.din(w_dff_A_DhQvmmJb6_0),.clk(gclk));
	jdff dff_A_yWxvpk0L9_0(.dout(w_dff_A_LeDvghwO5_0),.din(w_dff_A_yWxvpk0L9_0),.clk(gclk));
	jdff dff_A_LeDvghwO5_0(.dout(w_dff_A_uAscGIOG7_0),.din(w_dff_A_LeDvghwO5_0),.clk(gclk));
	jdff dff_A_uAscGIOG7_0(.dout(w_dff_A_2fGdQq3H6_0),.din(w_dff_A_uAscGIOG7_0),.clk(gclk));
	jdff dff_A_2fGdQq3H6_0(.dout(w_dff_A_OOpz2K8o9_0),.din(w_dff_A_2fGdQq3H6_0),.clk(gclk));
	jdff dff_A_OOpz2K8o9_0(.dout(w_dff_A_IsIB4EQA3_0),.din(w_dff_A_OOpz2K8o9_0),.clk(gclk));
	jdff dff_A_IsIB4EQA3_0(.dout(w_dff_A_8Ch04RuM5_0),.din(w_dff_A_IsIB4EQA3_0),.clk(gclk));
	jdff dff_A_8Ch04RuM5_0(.dout(w_dff_A_HffPPdwN1_0),.din(w_dff_A_8Ch04RuM5_0),.clk(gclk));
	jdff dff_A_HffPPdwN1_0(.dout(w_dff_A_U6TSY54Z8_0),.din(w_dff_A_HffPPdwN1_0),.clk(gclk));
	jdff dff_A_U6TSY54Z8_0(.dout(w_dff_A_wp0QpJAL5_0),.din(w_dff_A_U6TSY54Z8_0),.clk(gclk));
	jdff dff_A_wp0QpJAL5_0(.dout(w_dff_A_UzUYjMgM6_0),.din(w_dff_A_wp0QpJAL5_0),.clk(gclk));
	jdff dff_A_UzUYjMgM6_0(.dout(G373),.din(w_dff_A_UzUYjMgM6_0),.clk(gclk));
	jdff dff_A_WgdesOxS6_2(.dout(w_dff_A_0MAjtAZX9_0),.din(w_dff_A_WgdesOxS6_2),.clk(gclk));
	jdff dff_A_0MAjtAZX9_0(.dout(w_dff_A_XnWGpai63_0),.din(w_dff_A_0MAjtAZX9_0),.clk(gclk));
	jdff dff_A_XnWGpai63_0(.dout(w_dff_A_uPiXm35k8_0),.din(w_dff_A_XnWGpai63_0),.clk(gclk));
	jdff dff_A_uPiXm35k8_0(.dout(w_dff_A_Jpk3n4926_0),.din(w_dff_A_uPiXm35k8_0),.clk(gclk));
	jdff dff_A_Jpk3n4926_0(.dout(w_dff_A_MiuRKQMd9_0),.din(w_dff_A_Jpk3n4926_0),.clk(gclk));
	jdff dff_A_MiuRKQMd9_0(.dout(w_dff_A_h8e3CzGx6_0),.din(w_dff_A_MiuRKQMd9_0),.clk(gclk));
	jdff dff_A_h8e3CzGx6_0(.dout(w_dff_A_JjFLABj79_0),.din(w_dff_A_h8e3CzGx6_0),.clk(gclk));
	jdff dff_A_JjFLABj79_0(.dout(w_dff_A_iGD8WHOb0_0),.din(w_dff_A_JjFLABj79_0),.clk(gclk));
	jdff dff_A_iGD8WHOb0_0(.dout(w_dff_A_4rCrF3xX4_0),.din(w_dff_A_iGD8WHOb0_0),.clk(gclk));
	jdff dff_A_4rCrF3xX4_0(.dout(w_dff_A_6dZOUxLq7_0),.din(w_dff_A_4rCrF3xX4_0),.clk(gclk));
	jdff dff_A_6dZOUxLq7_0(.dout(G258),.din(w_dff_A_6dZOUxLq7_0),.clk(gclk));
	jdff dff_A_gVGYXbAZ9_2(.dout(w_dff_A_NqrjpIF95_0),.din(w_dff_A_gVGYXbAZ9_2),.clk(gclk));
	jdff dff_A_NqrjpIF95_0(.dout(w_dff_A_HNivIQsl8_0),.din(w_dff_A_NqrjpIF95_0),.clk(gclk));
	jdff dff_A_HNivIQsl8_0(.dout(w_dff_A_QY9Wrn8O2_0),.din(w_dff_A_HNivIQsl8_0),.clk(gclk));
	jdff dff_A_QY9Wrn8O2_0(.dout(w_dff_A_TuTty8EX9_0),.din(w_dff_A_QY9Wrn8O2_0),.clk(gclk));
	jdff dff_A_TuTty8EX9_0(.dout(w_dff_A_LX2u7u419_0),.din(w_dff_A_TuTty8EX9_0),.clk(gclk));
	jdff dff_A_LX2u7u419_0(.dout(w_dff_A_yAKUWmNi4_0),.din(w_dff_A_LX2u7u419_0),.clk(gclk));
	jdff dff_A_yAKUWmNi4_0(.dout(w_dff_A_7HlLi65N3_0),.din(w_dff_A_yAKUWmNi4_0),.clk(gclk));
	jdff dff_A_7HlLi65N3_0(.dout(w_dff_A_qsajmEeY3_0),.din(w_dff_A_7HlLi65N3_0),.clk(gclk));
	jdff dff_A_qsajmEeY3_0(.dout(w_dff_A_J8pd6cwc7_0),.din(w_dff_A_qsajmEeY3_0),.clk(gclk));
	jdff dff_A_J8pd6cwc7_0(.dout(w_dff_A_52ewoE7D6_0),.din(w_dff_A_J8pd6cwc7_0),.clk(gclk));
	jdff dff_A_52ewoE7D6_0(.dout(G264),.din(w_dff_A_52ewoE7D6_0),.clk(gclk));
	jdff dff_A_hPnAfq4F4_2(.dout(w_dff_A_iNwMUUHK5_0),.din(w_dff_A_hPnAfq4F4_2),.clk(gclk));
	jdff dff_A_iNwMUUHK5_0(.dout(w_dff_A_PFOM2LhJ2_0),.din(w_dff_A_iNwMUUHK5_0),.clk(gclk));
	jdff dff_A_PFOM2LhJ2_0(.dout(w_dff_A_nWiicRqs2_0),.din(w_dff_A_PFOM2LhJ2_0),.clk(gclk));
	jdff dff_A_nWiicRqs2_0(.dout(w_dff_A_rnXX74dU7_0),.din(w_dff_A_nWiicRqs2_0),.clk(gclk));
	jdff dff_A_rnXX74dU7_0(.dout(w_dff_A_a49ATBdq9_0),.din(w_dff_A_rnXX74dU7_0),.clk(gclk));
	jdff dff_A_a49ATBdq9_0(.dout(w_dff_A_xbkIkvNl6_0),.din(w_dff_A_a49ATBdq9_0),.clk(gclk));
	jdff dff_A_xbkIkvNl6_0(.dout(w_dff_A_APefuJA21_0),.din(w_dff_A_xbkIkvNl6_0),.clk(gclk));
	jdff dff_A_APefuJA21_0(.dout(w_dff_A_r4f54s5A3_0),.din(w_dff_A_APefuJA21_0),.clk(gclk));
	jdff dff_A_r4f54s5A3_0(.dout(w_dff_A_heXjPChd8_0),.din(w_dff_A_r4f54s5A3_0),.clk(gclk));
	jdff dff_A_heXjPChd8_0(.dout(w_dff_A_Vz7q3ErZ5_0),.din(w_dff_A_heXjPChd8_0),.clk(gclk));
	jdff dff_A_Vz7q3ErZ5_0(.dout(w_dff_A_1OtQR8rD3_0),.din(w_dff_A_Vz7q3ErZ5_0),.clk(gclk));
	jdff dff_A_1OtQR8rD3_0(.dout(w_dff_A_MIaF2AKB6_0),.din(w_dff_A_1OtQR8rD3_0),.clk(gclk));
	jdff dff_A_MIaF2AKB6_0(.dout(w_dff_A_nGmhZ0yO2_0),.din(w_dff_A_MIaF2AKB6_0),.clk(gclk));
	jdff dff_A_nGmhZ0yO2_0(.dout(w_dff_A_EdCsBd2c5_0),.din(w_dff_A_nGmhZ0yO2_0),.clk(gclk));
	jdff dff_A_EdCsBd2c5_0(.dout(w_dff_A_T4b63vDR7_0),.din(w_dff_A_EdCsBd2c5_0),.clk(gclk));
	jdff dff_A_T4b63vDR7_0(.dout(w_dff_A_A1kwbq6i9_0),.din(w_dff_A_T4b63vDR7_0),.clk(gclk));
	jdff dff_A_A1kwbq6i9_0(.dout(w_dff_A_QY6wIL7V5_0),.din(w_dff_A_A1kwbq6i9_0),.clk(gclk));
	jdff dff_A_QY6wIL7V5_0(.dout(w_dff_A_oyuiGHus1_0),.din(w_dff_A_QY6wIL7V5_0),.clk(gclk));
	jdff dff_A_oyuiGHus1_0(.dout(w_dff_A_FoXPssr27_0),.din(w_dff_A_oyuiGHus1_0),.clk(gclk));
	jdff dff_A_FoXPssr27_0(.dout(w_dff_A_L2IfLhs72_0),.din(w_dff_A_FoXPssr27_0),.clk(gclk));
	jdff dff_A_L2IfLhs72_0(.dout(w_dff_A_chT3XV4f0_0),.din(w_dff_A_L2IfLhs72_0),.clk(gclk));
	jdff dff_A_chT3XV4f0_0(.dout(w_dff_A_fumqalSS2_0),.din(w_dff_A_chT3XV4f0_0),.clk(gclk));
	jdff dff_A_fumqalSS2_0(.dout(w_dff_A_2nnZdTm25_0),.din(w_dff_A_fumqalSS2_0),.clk(gclk));
	jdff dff_A_2nnZdTm25_0(.dout(w_dff_A_2wIBugvy5_0),.din(w_dff_A_2nnZdTm25_0),.clk(gclk));
	jdff dff_A_2wIBugvy5_0(.dout(G388),.din(w_dff_A_2wIBugvy5_0),.clk(gclk));
	jdff dff_A_gTjHNFqz8_2(.dout(w_dff_A_WKNUtcIs5_0),.din(w_dff_A_gTjHNFqz8_2),.clk(gclk));
	jdff dff_A_WKNUtcIs5_0(.dout(w_dff_A_rbcDPmp47_0),.din(w_dff_A_WKNUtcIs5_0),.clk(gclk));
	jdff dff_A_rbcDPmp47_0(.dout(w_dff_A_Wn738bAv0_0),.din(w_dff_A_rbcDPmp47_0),.clk(gclk));
	jdff dff_A_Wn738bAv0_0(.dout(w_dff_A_tevt4oG43_0),.din(w_dff_A_Wn738bAv0_0),.clk(gclk));
	jdff dff_A_tevt4oG43_0(.dout(w_dff_A_gMkcfKNc5_0),.din(w_dff_A_tevt4oG43_0),.clk(gclk));
	jdff dff_A_gMkcfKNc5_0(.dout(w_dff_A_hA6kEm0g5_0),.din(w_dff_A_gMkcfKNc5_0),.clk(gclk));
	jdff dff_A_hA6kEm0g5_0(.dout(w_dff_A_n20VkMtD0_0),.din(w_dff_A_hA6kEm0g5_0),.clk(gclk));
	jdff dff_A_n20VkMtD0_0(.dout(w_dff_A_HeVyyHWm8_0),.din(w_dff_A_n20VkMtD0_0),.clk(gclk));
	jdff dff_A_HeVyyHWm8_0(.dout(w_dff_A_OEhLT8dJ8_0),.din(w_dff_A_HeVyyHWm8_0),.clk(gclk));
	jdff dff_A_OEhLT8dJ8_0(.dout(w_dff_A_QxwFQzQX8_0),.din(w_dff_A_OEhLT8dJ8_0),.clk(gclk));
	jdff dff_A_QxwFQzQX8_0(.dout(w_dff_A_u5vFU4tv9_0),.din(w_dff_A_QxwFQzQX8_0),.clk(gclk));
	jdff dff_A_u5vFU4tv9_0(.dout(w_dff_A_LiReZLmP4_0),.din(w_dff_A_u5vFU4tv9_0),.clk(gclk));
	jdff dff_A_LiReZLmP4_0(.dout(w_dff_A_Vlzubrbv1_0),.din(w_dff_A_LiReZLmP4_0),.clk(gclk));
	jdff dff_A_Vlzubrbv1_0(.dout(w_dff_A_h0zZEJrs3_0),.din(w_dff_A_Vlzubrbv1_0),.clk(gclk));
	jdff dff_A_h0zZEJrs3_0(.dout(w_dff_A_7VuxU29p2_0),.din(w_dff_A_h0zZEJrs3_0),.clk(gclk));
	jdff dff_A_7VuxU29p2_0(.dout(w_dff_A_lKhtrzhY2_0),.din(w_dff_A_7VuxU29p2_0),.clk(gclk));
	jdff dff_A_lKhtrzhY2_0(.dout(w_dff_A_TmBXw6hR3_0),.din(w_dff_A_lKhtrzhY2_0),.clk(gclk));
	jdff dff_A_TmBXw6hR3_0(.dout(w_dff_A_peZAriNm4_0),.din(w_dff_A_TmBXw6hR3_0),.clk(gclk));
	jdff dff_A_peZAriNm4_0(.dout(w_dff_A_xZMnHIwy8_0),.din(w_dff_A_peZAriNm4_0),.clk(gclk));
	jdff dff_A_xZMnHIwy8_0(.dout(w_dff_A_4uGXzQWa7_0),.din(w_dff_A_xZMnHIwy8_0),.clk(gclk));
	jdff dff_A_4uGXzQWa7_0(.dout(w_dff_A_Wyp9HWKV7_0),.din(w_dff_A_4uGXzQWa7_0),.clk(gclk));
	jdff dff_A_Wyp9HWKV7_0(.dout(w_dff_A_MAcM2TRw3_0),.din(w_dff_A_Wyp9HWKV7_0),.clk(gclk));
	jdff dff_A_MAcM2TRw3_0(.dout(w_dff_A_lwhkvxhm6_0),.din(w_dff_A_MAcM2TRw3_0),.clk(gclk));
	jdff dff_A_lwhkvxhm6_0(.dout(w_dff_A_5wo7rnwH5_0),.din(w_dff_A_lwhkvxhm6_0),.clk(gclk));
	jdff dff_A_5wo7rnwH5_0(.dout(w_dff_A_CYQWdov97_0),.din(w_dff_A_5wo7rnwH5_0),.clk(gclk));
	jdff dff_A_CYQWdov97_0(.dout(w_dff_A_z7yc9I0i3_0),.din(w_dff_A_CYQWdov97_0),.clk(gclk));
	jdff dff_A_z7yc9I0i3_0(.dout(G391),.din(w_dff_A_z7yc9I0i3_0),.clk(gclk));
	jdff dff_A_5B1bkyF47_2(.dout(w_dff_A_Ttn95e517_0),.din(w_dff_A_5B1bkyF47_2),.clk(gclk));
	jdff dff_A_Ttn95e517_0(.dout(w_dff_A_8t703pIG5_0),.din(w_dff_A_Ttn95e517_0),.clk(gclk));
	jdff dff_A_8t703pIG5_0(.dout(w_dff_A_qUGBXbCV2_0),.din(w_dff_A_8t703pIG5_0),.clk(gclk));
	jdff dff_A_qUGBXbCV2_0(.dout(w_dff_A_L8C51wfk8_0),.din(w_dff_A_qUGBXbCV2_0),.clk(gclk));
	jdff dff_A_L8C51wfk8_0(.dout(w_dff_A_sJCoUQNH1_0),.din(w_dff_A_L8C51wfk8_0),.clk(gclk));
	jdff dff_A_sJCoUQNH1_0(.dout(w_dff_A_GmKIpH9Y4_0),.din(w_dff_A_sJCoUQNH1_0),.clk(gclk));
	jdff dff_A_GmKIpH9Y4_0(.dout(w_dff_A_rNfIFAE02_0),.din(w_dff_A_GmKIpH9Y4_0),.clk(gclk));
	jdff dff_A_rNfIFAE02_0(.dout(w_dff_A_4f4qySzM1_0),.din(w_dff_A_rNfIFAE02_0),.clk(gclk));
	jdff dff_A_4f4qySzM1_0(.dout(w_dff_A_3ncSnTUK7_0),.din(w_dff_A_4f4qySzM1_0),.clk(gclk));
	jdff dff_A_3ncSnTUK7_0(.dout(w_dff_A_2eEKXkb91_0),.din(w_dff_A_3ncSnTUK7_0),.clk(gclk));
	jdff dff_A_2eEKXkb91_0(.dout(w_dff_A_MyHPrs2b8_0),.din(w_dff_A_2eEKXkb91_0),.clk(gclk));
	jdff dff_A_MyHPrs2b8_0(.dout(w_dff_A_5VaeJNyz4_0),.din(w_dff_A_MyHPrs2b8_0),.clk(gclk));
	jdff dff_A_5VaeJNyz4_0(.dout(w_dff_A_h2PRlNUO8_0),.din(w_dff_A_5VaeJNyz4_0),.clk(gclk));
	jdff dff_A_h2PRlNUO8_0(.dout(w_dff_A_LUECO1XC8_0),.din(w_dff_A_h2PRlNUO8_0),.clk(gclk));
	jdff dff_A_LUECO1XC8_0(.dout(w_dff_A_vnvenVbj8_0),.din(w_dff_A_LUECO1XC8_0),.clk(gclk));
	jdff dff_A_vnvenVbj8_0(.dout(w_dff_A_qhYYZH6r5_0),.din(w_dff_A_vnvenVbj8_0),.clk(gclk));
	jdff dff_A_qhYYZH6r5_0(.dout(w_dff_A_nT7D9dZC8_0),.din(w_dff_A_qhYYZH6r5_0),.clk(gclk));
	jdff dff_A_nT7D9dZC8_0(.dout(w_dff_A_EX1eb4ry4_0),.din(w_dff_A_nT7D9dZC8_0),.clk(gclk));
	jdff dff_A_EX1eb4ry4_0(.dout(w_dff_A_lk9Gz33w6_0),.din(w_dff_A_EX1eb4ry4_0),.clk(gclk));
	jdff dff_A_lk9Gz33w6_0(.dout(w_dff_A_RcZ9vyPH6_0),.din(w_dff_A_lk9Gz33w6_0),.clk(gclk));
	jdff dff_A_RcZ9vyPH6_0(.dout(w_dff_A_5XM4gxYI7_0),.din(w_dff_A_RcZ9vyPH6_0),.clk(gclk));
	jdff dff_A_5XM4gxYI7_0(.dout(w_dff_A_nj0FVd7u8_0),.din(w_dff_A_5XM4gxYI7_0),.clk(gclk));
	jdff dff_A_nj0FVd7u8_0(.dout(w_dff_A_UFeAFPWr9_0),.din(w_dff_A_nj0FVd7u8_0),.clk(gclk));
	jdff dff_A_UFeAFPWr9_0(.dout(w_dff_A_B9QL6Qe05_0),.din(w_dff_A_UFeAFPWr9_0),.clk(gclk));
	jdff dff_A_B9QL6Qe05_0(.dout(w_dff_A_ped9jlaL8_0),.din(w_dff_A_B9QL6Qe05_0),.clk(gclk));
	jdff dff_A_ped9jlaL8_0(.dout(w_dff_A_IokUSfhx5_0),.din(w_dff_A_ped9jlaL8_0),.clk(gclk));
	jdff dff_A_IokUSfhx5_0(.dout(w_dff_A_b6l6bhqQ5_0),.din(w_dff_A_IokUSfhx5_0),.clk(gclk));
	jdff dff_A_b6l6bhqQ5_0(.dout(w_dff_A_gIFno2YV5_0),.din(w_dff_A_b6l6bhqQ5_0),.clk(gclk));
	jdff dff_A_gIFno2YV5_0(.dout(w_dff_A_zTDeMC165_0),.din(w_dff_A_gIFno2YV5_0),.clk(gclk));
	jdff dff_A_zTDeMC165_0(.dout(G394),.din(w_dff_A_zTDeMC165_0),.clk(gclk));
	jdff dff_A_fpenTOu76_2(.dout(w_dff_A_cwWDxqXY1_0),.din(w_dff_A_fpenTOu76_2),.clk(gclk));
	jdff dff_A_cwWDxqXY1_0(.dout(w_dff_A_CAivFeWN1_0),.din(w_dff_A_cwWDxqXY1_0),.clk(gclk));
	jdff dff_A_CAivFeWN1_0(.dout(w_dff_A_5BBLyt4O1_0),.din(w_dff_A_CAivFeWN1_0),.clk(gclk));
	jdff dff_A_5BBLyt4O1_0(.dout(w_dff_A_PuUG3zsC7_0),.din(w_dff_A_5BBLyt4O1_0),.clk(gclk));
	jdff dff_A_PuUG3zsC7_0(.dout(w_dff_A_LscEx0BE1_0),.din(w_dff_A_PuUG3zsC7_0),.clk(gclk));
	jdff dff_A_LscEx0BE1_0(.dout(w_dff_A_7GqgwZiS1_0),.din(w_dff_A_LscEx0BE1_0),.clk(gclk));
	jdff dff_A_7GqgwZiS1_0(.dout(w_dff_A_v8dGGnxG1_0),.din(w_dff_A_7GqgwZiS1_0),.clk(gclk));
	jdff dff_A_v8dGGnxG1_0(.dout(w_dff_A_6jUbPnNn8_0),.din(w_dff_A_v8dGGnxG1_0),.clk(gclk));
	jdff dff_A_6jUbPnNn8_0(.dout(w_dff_A_jWCE1zxJ0_0),.din(w_dff_A_6jUbPnNn8_0),.clk(gclk));
	jdff dff_A_jWCE1zxJ0_0(.dout(w_dff_A_djldMywr3_0),.din(w_dff_A_jWCE1zxJ0_0),.clk(gclk));
	jdff dff_A_djldMywr3_0(.dout(w_dff_A_H2nKMvgE4_0),.din(w_dff_A_djldMywr3_0),.clk(gclk));
	jdff dff_A_H2nKMvgE4_0(.dout(w_dff_A_5eLdNyu16_0),.din(w_dff_A_H2nKMvgE4_0),.clk(gclk));
	jdff dff_A_5eLdNyu16_0(.dout(w_dff_A_DLAr7g077_0),.din(w_dff_A_5eLdNyu16_0),.clk(gclk));
	jdff dff_A_DLAr7g077_0(.dout(w_dff_A_HlNsc1Mn2_0),.din(w_dff_A_DLAr7g077_0),.clk(gclk));
	jdff dff_A_HlNsc1Mn2_0(.dout(w_dff_A_CA924rQb5_0),.din(w_dff_A_HlNsc1Mn2_0),.clk(gclk));
	jdff dff_A_CA924rQb5_0(.dout(w_dff_A_IhlIqXHJ2_0),.din(w_dff_A_CA924rQb5_0),.clk(gclk));
	jdff dff_A_IhlIqXHJ2_0(.dout(w_dff_A_GtW6pevU5_0),.din(w_dff_A_IhlIqXHJ2_0),.clk(gclk));
	jdff dff_A_GtW6pevU5_0(.dout(w_dff_A_AT9S9VJt0_0),.din(w_dff_A_GtW6pevU5_0),.clk(gclk));
	jdff dff_A_AT9S9VJt0_0(.dout(w_dff_A_wKFIr6Cp0_0),.din(w_dff_A_AT9S9VJt0_0),.clk(gclk));
	jdff dff_A_wKFIr6Cp0_0(.dout(w_dff_A_dDURwMH97_0),.din(w_dff_A_wKFIr6Cp0_0),.clk(gclk));
	jdff dff_A_dDURwMH97_0(.dout(w_dff_A_2RcdRk0R1_0),.din(w_dff_A_dDURwMH97_0),.clk(gclk));
	jdff dff_A_2RcdRk0R1_0(.dout(w_dff_A_uR8sQkJh2_0),.din(w_dff_A_2RcdRk0R1_0),.clk(gclk));
	jdff dff_A_uR8sQkJh2_0(.dout(w_dff_A_aVhbpkvT9_0),.din(w_dff_A_uR8sQkJh2_0),.clk(gclk));
	jdff dff_A_aVhbpkvT9_0(.dout(w_dff_A_tGUeM6AL7_0),.din(w_dff_A_aVhbpkvT9_0),.clk(gclk));
	jdff dff_A_tGUeM6AL7_0(.dout(w_dff_A_JGTVUj4L7_0),.din(w_dff_A_tGUeM6AL7_0),.clk(gclk));
	jdff dff_A_JGTVUj4L7_0(.dout(w_dff_A_5YcxzyGN2_0),.din(w_dff_A_JGTVUj4L7_0),.clk(gclk));
	jdff dff_A_5YcxzyGN2_0(.dout(w_dff_A_MNdxUWzQ8_0),.din(w_dff_A_5YcxzyGN2_0),.clk(gclk));
	jdff dff_A_MNdxUWzQ8_0(.dout(w_dff_A_yF8MwC7r1_0),.din(w_dff_A_MNdxUWzQ8_0),.clk(gclk));
	jdff dff_A_yF8MwC7r1_0(.dout(w_dff_A_AMEMdVHP1_0),.din(w_dff_A_yF8MwC7r1_0),.clk(gclk));
	jdff dff_A_AMEMdVHP1_0(.dout(w_dff_A_ttfj0vH04_0),.din(w_dff_A_AMEMdVHP1_0),.clk(gclk));
	jdff dff_A_ttfj0vH04_0(.dout(G397),.din(w_dff_A_ttfj0vH04_0),.clk(gclk));
	jdff dff_A_TNQcEwwd4_2(.dout(w_dff_A_RRZKL7iL4_0),.din(w_dff_A_TNQcEwwd4_2),.clk(gclk));
	jdff dff_A_RRZKL7iL4_0(.dout(w_dff_A_3P5NaF2r5_0),.din(w_dff_A_RRZKL7iL4_0),.clk(gclk));
	jdff dff_A_3P5NaF2r5_0(.dout(w_dff_A_YonoLV990_0),.din(w_dff_A_3P5NaF2r5_0),.clk(gclk));
	jdff dff_A_YonoLV990_0(.dout(w_dff_A_oHh0BOtM0_0),.din(w_dff_A_YonoLV990_0),.clk(gclk));
	jdff dff_A_oHh0BOtM0_0(.dout(w_dff_A_3nrLiEVZ3_0),.din(w_dff_A_oHh0BOtM0_0),.clk(gclk));
	jdff dff_A_3nrLiEVZ3_0(.dout(w_dff_A_RIjcep6Q8_0),.din(w_dff_A_3nrLiEVZ3_0),.clk(gclk));
	jdff dff_A_RIjcep6Q8_0(.dout(w_dff_A_g23pRVwW7_0),.din(w_dff_A_RIjcep6Q8_0),.clk(gclk));
	jdff dff_A_g23pRVwW7_0(.dout(w_dff_A_neoHDwvD0_0),.din(w_dff_A_g23pRVwW7_0),.clk(gclk));
	jdff dff_A_neoHDwvD0_0(.dout(w_dff_A_ZISIHtAJ1_0),.din(w_dff_A_neoHDwvD0_0),.clk(gclk));
	jdff dff_A_ZISIHtAJ1_0(.dout(w_dff_A_qlxHZB3k5_0),.din(w_dff_A_ZISIHtAJ1_0),.clk(gclk));
	jdff dff_A_qlxHZB3k5_0(.dout(w_dff_A_nLYwuqj32_0),.din(w_dff_A_qlxHZB3k5_0),.clk(gclk));
	jdff dff_A_nLYwuqj32_0(.dout(w_dff_A_qSlaXN8l8_0),.din(w_dff_A_nLYwuqj32_0),.clk(gclk));
	jdff dff_A_qSlaXN8l8_0(.dout(w_dff_A_itfXPfYC3_0),.din(w_dff_A_qSlaXN8l8_0),.clk(gclk));
	jdff dff_A_itfXPfYC3_0(.dout(w_dff_A_vwKU9xyl8_0),.din(w_dff_A_itfXPfYC3_0),.clk(gclk));
	jdff dff_A_vwKU9xyl8_0(.dout(w_dff_A_1DnrtLmJ0_0),.din(w_dff_A_vwKU9xyl8_0),.clk(gclk));
	jdff dff_A_1DnrtLmJ0_0(.dout(w_dff_A_HZeatMJE7_0),.din(w_dff_A_1DnrtLmJ0_0),.clk(gclk));
	jdff dff_A_HZeatMJE7_0(.dout(w_dff_A_4xjDzBpk8_0),.din(w_dff_A_HZeatMJE7_0),.clk(gclk));
	jdff dff_A_4xjDzBpk8_0(.dout(w_dff_A_Wfi1tSMF9_0),.din(w_dff_A_4xjDzBpk8_0),.clk(gclk));
	jdff dff_A_Wfi1tSMF9_0(.dout(w_dff_A_4arLJuD57_0),.din(w_dff_A_Wfi1tSMF9_0),.clk(gclk));
	jdff dff_A_4arLJuD57_0(.dout(G376),.din(w_dff_A_4arLJuD57_0),.clk(gclk));
	jdff dff_A_RCtQWRw62_2(.dout(w_dff_A_wcCPGPVJ7_0),.din(w_dff_A_RCtQWRw62_2),.clk(gclk));
	jdff dff_A_wcCPGPVJ7_0(.dout(w_dff_A_YvBnnsTX1_0),.din(w_dff_A_wcCPGPVJ7_0),.clk(gclk));
	jdff dff_A_YvBnnsTX1_0(.dout(w_dff_A_2S5E8xlm4_0),.din(w_dff_A_YvBnnsTX1_0),.clk(gclk));
	jdff dff_A_2S5E8xlm4_0(.dout(w_dff_A_F3SD8t3w8_0),.din(w_dff_A_2S5E8xlm4_0),.clk(gclk));
	jdff dff_A_F3SD8t3w8_0(.dout(w_dff_A_CozWiyfC4_0),.din(w_dff_A_F3SD8t3w8_0),.clk(gclk));
	jdff dff_A_CozWiyfC4_0(.dout(w_dff_A_pkWkkBzf1_0),.din(w_dff_A_CozWiyfC4_0),.clk(gclk));
	jdff dff_A_pkWkkBzf1_0(.dout(w_dff_A_ROpv3ED38_0),.din(w_dff_A_pkWkkBzf1_0),.clk(gclk));
	jdff dff_A_ROpv3ED38_0(.dout(w_dff_A_9gQuaPxf8_0),.din(w_dff_A_ROpv3ED38_0),.clk(gclk));
	jdff dff_A_9gQuaPxf8_0(.dout(w_dff_A_LH8pqbTX2_0),.din(w_dff_A_9gQuaPxf8_0),.clk(gclk));
	jdff dff_A_LH8pqbTX2_0(.dout(w_dff_A_x10gWTsH5_0),.din(w_dff_A_LH8pqbTX2_0),.clk(gclk));
	jdff dff_A_x10gWTsH5_0(.dout(w_dff_A_TxYwJokZ6_0),.din(w_dff_A_x10gWTsH5_0),.clk(gclk));
	jdff dff_A_TxYwJokZ6_0(.dout(w_dff_A_cN0aZ28w5_0),.din(w_dff_A_TxYwJokZ6_0),.clk(gclk));
	jdff dff_A_cN0aZ28w5_0(.dout(w_dff_A_s8ahpQih9_0),.din(w_dff_A_cN0aZ28w5_0),.clk(gclk));
	jdff dff_A_s8ahpQih9_0(.dout(w_dff_A_qs21yKio3_0),.din(w_dff_A_s8ahpQih9_0),.clk(gclk));
	jdff dff_A_qs21yKio3_0(.dout(w_dff_A_6o22pCvI9_0),.din(w_dff_A_qs21yKio3_0),.clk(gclk));
	jdff dff_A_6o22pCvI9_0(.dout(w_dff_A_pEagct3R1_0),.din(w_dff_A_6o22pCvI9_0),.clk(gclk));
	jdff dff_A_pEagct3R1_0(.dout(w_dff_A_ItHBpcHd1_0),.din(w_dff_A_pEagct3R1_0),.clk(gclk));
	jdff dff_A_ItHBpcHd1_0(.dout(w_dff_A_hR0gFTZn6_0),.din(w_dff_A_ItHBpcHd1_0),.clk(gclk));
	jdff dff_A_hR0gFTZn6_0(.dout(w_dff_A_VP3xdPTV0_0),.din(w_dff_A_hR0gFTZn6_0),.clk(gclk));
	jdff dff_A_VP3xdPTV0_0(.dout(w_dff_A_pqvkgzNJ8_0),.din(w_dff_A_VP3xdPTV0_0),.clk(gclk));
	jdff dff_A_pqvkgzNJ8_0(.dout(w_dff_A_WPg6b8Tt1_0),.din(w_dff_A_pqvkgzNJ8_0),.clk(gclk));
	jdff dff_A_WPg6b8Tt1_0(.dout(G379),.din(w_dff_A_WPg6b8Tt1_0),.clk(gclk));
	jdff dff_A_OwLg3vyW3_2(.dout(w_dff_A_fvxalksz5_0),.din(w_dff_A_OwLg3vyW3_2),.clk(gclk));
	jdff dff_A_fvxalksz5_0(.dout(w_dff_A_rC8rH8iX2_0),.din(w_dff_A_fvxalksz5_0),.clk(gclk));
	jdff dff_A_rC8rH8iX2_0(.dout(w_dff_A_srhtw1sZ8_0),.din(w_dff_A_rC8rH8iX2_0),.clk(gclk));
	jdff dff_A_srhtw1sZ8_0(.dout(w_dff_A_D8D7JTuH6_0),.din(w_dff_A_srhtw1sZ8_0),.clk(gclk));
	jdff dff_A_D8D7JTuH6_0(.dout(w_dff_A_BeNOCHJK7_0),.din(w_dff_A_D8D7JTuH6_0),.clk(gclk));
	jdff dff_A_BeNOCHJK7_0(.dout(w_dff_A_y8Nwq1Ec0_0),.din(w_dff_A_BeNOCHJK7_0),.clk(gclk));
	jdff dff_A_y8Nwq1Ec0_0(.dout(w_dff_A_vu1tZF2J9_0),.din(w_dff_A_y8Nwq1Ec0_0),.clk(gclk));
	jdff dff_A_vu1tZF2J9_0(.dout(w_dff_A_1hAiqw6U1_0),.din(w_dff_A_vu1tZF2J9_0),.clk(gclk));
	jdff dff_A_1hAiqw6U1_0(.dout(w_dff_A_wTmaZm8A1_0),.din(w_dff_A_1hAiqw6U1_0),.clk(gclk));
	jdff dff_A_wTmaZm8A1_0(.dout(w_dff_A_qoAP9IPY5_0),.din(w_dff_A_wTmaZm8A1_0),.clk(gclk));
	jdff dff_A_qoAP9IPY5_0(.dout(w_dff_A_Vn4DOyHy3_0),.din(w_dff_A_qoAP9IPY5_0),.clk(gclk));
	jdff dff_A_Vn4DOyHy3_0(.dout(w_dff_A_BkJWTfI02_0),.din(w_dff_A_Vn4DOyHy3_0),.clk(gclk));
	jdff dff_A_BkJWTfI02_0(.dout(w_dff_A_JoP7uMAJ8_0),.din(w_dff_A_BkJWTfI02_0),.clk(gclk));
	jdff dff_A_JoP7uMAJ8_0(.dout(w_dff_A_Eo61JeLz8_0),.din(w_dff_A_JoP7uMAJ8_0),.clk(gclk));
	jdff dff_A_Eo61JeLz8_0(.dout(w_dff_A_h2gs3CPy0_0),.din(w_dff_A_Eo61JeLz8_0),.clk(gclk));
	jdff dff_A_h2gs3CPy0_0(.dout(w_dff_A_3hektXhU1_0),.din(w_dff_A_h2gs3CPy0_0),.clk(gclk));
	jdff dff_A_3hektXhU1_0(.dout(w_dff_A_8z8TXkf17_0),.din(w_dff_A_3hektXhU1_0),.clk(gclk));
	jdff dff_A_8z8TXkf17_0(.dout(w_dff_A_b83fJIyn8_0),.din(w_dff_A_8z8TXkf17_0),.clk(gclk));
	jdff dff_A_b83fJIyn8_0(.dout(w_dff_A_SeBPHW0r9_0),.din(w_dff_A_b83fJIyn8_0),.clk(gclk));
	jdff dff_A_SeBPHW0r9_0(.dout(w_dff_A_ksVtyhS00_0),.din(w_dff_A_SeBPHW0r9_0),.clk(gclk));
	jdff dff_A_ksVtyhS00_0(.dout(w_dff_A_4eq7X4Hm1_0),.din(w_dff_A_ksVtyhS00_0),.clk(gclk));
	jdff dff_A_4eq7X4Hm1_0(.dout(G382),.din(w_dff_A_4eq7X4Hm1_0),.clk(gclk));
	jdff dff_A_BjAxq4mU0_2(.dout(w_dff_A_AlaYxrBK0_0),.din(w_dff_A_BjAxq4mU0_2),.clk(gclk));
	jdff dff_A_AlaYxrBK0_0(.dout(w_dff_A_8Np7gqqZ4_0),.din(w_dff_A_AlaYxrBK0_0),.clk(gclk));
	jdff dff_A_8Np7gqqZ4_0(.dout(w_dff_A_FjVQ1N0P3_0),.din(w_dff_A_8Np7gqqZ4_0),.clk(gclk));
	jdff dff_A_FjVQ1N0P3_0(.dout(w_dff_A_YizKHwPR9_0),.din(w_dff_A_FjVQ1N0P3_0),.clk(gclk));
	jdff dff_A_YizKHwPR9_0(.dout(w_dff_A_wMP8YfKD9_0),.din(w_dff_A_YizKHwPR9_0),.clk(gclk));
	jdff dff_A_wMP8YfKD9_0(.dout(w_dff_A_ktN8mmT99_0),.din(w_dff_A_wMP8YfKD9_0),.clk(gclk));
	jdff dff_A_ktN8mmT99_0(.dout(w_dff_A_JtAFwv1D8_0),.din(w_dff_A_ktN8mmT99_0),.clk(gclk));
	jdff dff_A_JtAFwv1D8_0(.dout(w_dff_A_GBlqMzBr5_0),.din(w_dff_A_JtAFwv1D8_0),.clk(gclk));
	jdff dff_A_GBlqMzBr5_0(.dout(w_dff_A_IV9sS5hg3_0),.din(w_dff_A_GBlqMzBr5_0),.clk(gclk));
	jdff dff_A_IV9sS5hg3_0(.dout(w_dff_A_tkCW5NPm9_0),.din(w_dff_A_IV9sS5hg3_0),.clk(gclk));
	jdff dff_A_tkCW5NPm9_0(.dout(w_dff_A_yYfyuP0p9_0),.din(w_dff_A_tkCW5NPm9_0),.clk(gclk));
	jdff dff_A_yYfyuP0p9_0(.dout(w_dff_A_JcOduGcL3_0),.din(w_dff_A_yYfyuP0p9_0),.clk(gclk));
	jdff dff_A_JcOduGcL3_0(.dout(w_dff_A_GqbmMOa65_0),.din(w_dff_A_JcOduGcL3_0),.clk(gclk));
	jdff dff_A_GqbmMOa65_0(.dout(w_dff_A_UW2H3DRS7_0),.din(w_dff_A_GqbmMOa65_0),.clk(gclk));
	jdff dff_A_UW2H3DRS7_0(.dout(w_dff_A_30Z7lW6x8_0),.din(w_dff_A_UW2H3DRS7_0),.clk(gclk));
	jdff dff_A_30Z7lW6x8_0(.dout(w_dff_A_e1uFaW1d9_0),.din(w_dff_A_30Z7lW6x8_0),.clk(gclk));
	jdff dff_A_e1uFaW1d9_0(.dout(w_dff_A_Yz3OiWn37_0),.din(w_dff_A_e1uFaW1d9_0),.clk(gclk));
	jdff dff_A_Yz3OiWn37_0(.dout(w_dff_A_AlUDMGWd7_0),.din(w_dff_A_Yz3OiWn37_0),.clk(gclk));
	jdff dff_A_AlUDMGWd7_0(.dout(w_dff_A_Ml85E7gs4_0),.din(w_dff_A_AlUDMGWd7_0),.clk(gclk));
	jdff dff_A_Ml85E7gs4_0(.dout(w_dff_A_rT4QnQEg1_0),.din(w_dff_A_Ml85E7gs4_0),.clk(gclk));
	jdff dff_A_rT4QnQEg1_0(.dout(w_dff_A_aUq1rw834_0),.din(w_dff_A_rT4QnQEg1_0),.clk(gclk));
	jdff dff_A_aUq1rw834_0(.dout(w_dff_A_08KUKXUt9_0),.din(w_dff_A_aUq1rw834_0),.clk(gclk));
	jdff dff_A_08KUKXUt9_0(.dout(w_dff_A_7nAMY1rS0_0),.din(w_dff_A_08KUKXUt9_0),.clk(gclk));
	jdff dff_A_7nAMY1rS0_0(.dout(G385),.din(w_dff_A_7nAMY1rS0_0),.clk(gclk));
	jdff dff_A_2m0EwwEg5_1(.dout(w_dff_A_I79e2AdF7_0),.din(w_dff_A_2m0EwwEg5_1),.clk(gclk));
	jdff dff_A_I79e2AdF7_0(.dout(w_dff_A_6GkCo1DY6_0),.din(w_dff_A_I79e2AdF7_0),.clk(gclk));
	jdff dff_A_6GkCo1DY6_0(.dout(w_dff_A_Lzey1E5Q1_0),.din(w_dff_A_6GkCo1DY6_0),.clk(gclk));
	jdff dff_A_Lzey1E5Q1_0(.dout(w_dff_A_vCziq13r3_0),.din(w_dff_A_Lzey1E5Q1_0),.clk(gclk));
	jdff dff_A_vCziq13r3_0(.dout(w_dff_A_GyxDS2LV9_0),.din(w_dff_A_vCziq13r3_0),.clk(gclk));
	jdff dff_A_GyxDS2LV9_0(.dout(w_dff_A_zjVysDTQ8_0),.din(w_dff_A_GyxDS2LV9_0),.clk(gclk));
	jdff dff_A_zjVysDTQ8_0(.dout(w_dff_A_kvqK0fIk0_0),.din(w_dff_A_zjVysDTQ8_0),.clk(gclk));
	jdff dff_A_kvqK0fIk0_0(.dout(w_dff_A_cugCo0mY1_0),.din(w_dff_A_kvqK0fIk0_0),.clk(gclk));
	jdff dff_A_cugCo0mY1_0(.dout(w_dff_A_yswv97vH4_0),.din(w_dff_A_cugCo0mY1_0),.clk(gclk));
	jdff dff_A_yswv97vH4_0(.dout(w_dff_A_OTfUuAtz5_0),.din(w_dff_A_yswv97vH4_0),.clk(gclk));
	jdff dff_A_OTfUuAtz5_0(.dout(w_dff_A_znDqZmWn2_0),.din(w_dff_A_OTfUuAtz5_0),.clk(gclk));
	jdff dff_A_znDqZmWn2_0(.dout(w_dff_A_AnYQczUh4_0),.din(w_dff_A_znDqZmWn2_0),.clk(gclk));
	jdff dff_A_AnYQczUh4_0(.dout(w_dff_A_21UXCDvQ8_0),.din(w_dff_A_AnYQczUh4_0),.clk(gclk));
	jdff dff_A_21UXCDvQ8_0(.dout(w_dff_A_2JPM1RxN1_0),.din(w_dff_A_21UXCDvQ8_0),.clk(gclk));
	jdff dff_A_2JPM1RxN1_0(.dout(w_dff_A_EPkzaIMr8_0),.din(w_dff_A_2JPM1RxN1_0),.clk(gclk));
	jdff dff_A_EPkzaIMr8_0(.dout(w_dff_A_3Zt31WK36_0),.din(w_dff_A_EPkzaIMr8_0),.clk(gclk));
	jdff dff_A_3Zt31WK36_0(.dout(w_dff_A_PY7L3h4w1_0),.din(w_dff_A_3Zt31WK36_0),.clk(gclk));
	jdff dff_A_PY7L3h4w1_0(.dout(w_dff_A_JT2Qq6Wb8_0),.din(w_dff_A_PY7L3h4w1_0),.clk(gclk));
	jdff dff_A_JT2Qq6Wb8_0(.dout(w_dff_A_UeYTx0wR9_0),.din(w_dff_A_JT2Qq6Wb8_0),.clk(gclk));
	jdff dff_A_UeYTx0wR9_0(.dout(w_dff_A_619BqzGV5_0),.din(w_dff_A_UeYTx0wR9_0),.clk(gclk));
	jdff dff_A_619BqzGV5_0(.dout(w_dff_A_jSmQNULw3_0),.din(w_dff_A_619BqzGV5_0),.clk(gclk));
	jdff dff_A_jSmQNULw3_0(.dout(w_dff_A_B36V9xMd3_0),.din(w_dff_A_jSmQNULw3_0),.clk(gclk));
	jdff dff_A_B36V9xMd3_0(.dout(w_dff_A_hSejvORY1_0),.din(w_dff_A_B36V9xMd3_0),.clk(gclk));
	jdff dff_A_hSejvORY1_0(.dout(w_dff_A_mRNqj3FC6_0),.din(w_dff_A_hSejvORY1_0),.clk(gclk));
	jdff dff_A_mRNqj3FC6_0(.dout(w_dff_A_WTjy3ssg7_0),.din(w_dff_A_mRNqj3FC6_0),.clk(gclk));
	jdff dff_A_WTjy3ssg7_0(.dout(w_dff_A_3zbxlb3T1_0),.din(w_dff_A_WTjy3ssg7_0),.clk(gclk));
	jdff dff_A_3zbxlb3T1_0(.dout(w_dff_A_ktr9uM4W4_0),.din(w_dff_A_3zbxlb3T1_0),.clk(gclk));
	jdff dff_A_ktr9uM4W4_0(.dout(G412),.din(w_dff_A_ktr9uM4W4_0),.clk(gclk));
	jdff dff_A_67FtK3pA2_1(.dout(w_dff_A_9dgE1jca0_0),.din(w_dff_A_67FtK3pA2_1),.clk(gclk));
	jdff dff_A_9dgE1jca0_0(.dout(w_dff_A_EP3B2JAi3_0),.din(w_dff_A_9dgE1jca0_0),.clk(gclk));
	jdff dff_A_EP3B2JAi3_0(.dout(w_dff_A_73V960tj1_0),.din(w_dff_A_EP3B2JAi3_0),.clk(gclk));
	jdff dff_A_73V960tj1_0(.dout(w_dff_A_9E9W0fdr0_0),.din(w_dff_A_73V960tj1_0),.clk(gclk));
	jdff dff_A_9E9W0fdr0_0(.dout(w_dff_A_D1dyQpxn2_0),.din(w_dff_A_9E9W0fdr0_0),.clk(gclk));
	jdff dff_A_D1dyQpxn2_0(.dout(w_dff_A_GXm1967f7_0),.din(w_dff_A_D1dyQpxn2_0),.clk(gclk));
	jdff dff_A_GXm1967f7_0(.dout(w_dff_A_XfvMSRI60_0),.din(w_dff_A_GXm1967f7_0),.clk(gclk));
	jdff dff_A_XfvMSRI60_0(.dout(w_dff_A_LEh3Tolj0_0),.din(w_dff_A_XfvMSRI60_0),.clk(gclk));
	jdff dff_A_LEh3Tolj0_0(.dout(w_dff_A_8dce071Y0_0),.din(w_dff_A_LEh3Tolj0_0),.clk(gclk));
	jdff dff_A_8dce071Y0_0(.dout(w_dff_A_bh23YbnF9_0),.din(w_dff_A_8dce071Y0_0),.clk(gclk));
	jdff dff_A_bh23YbnF9_0(.dout(w_dff_A_Sx3YBwK79_0),.din(w_dff_A_bh23YbnF9_0),.clk(gclk));
	jdff dff_A_Sx3YBwK79_0(.dout(w_dff_A_TMjMIq1m6_0),.din(w_dff_A_Sx3YBwK79_0),.clk(gclk));
	jdff dff_A_TMjMIq1m6_0(.dout(w_dff_A_fDoeD3mO3_0),.din(w_dff_A_TMjMIq1m6_0),.clk(gclk));
	jdff dff_A_fDoeD3mO3_0(.dout(w_dff_A_BrM7y7Wq4_0),.din(w_dff_A_fDoeD3mO3_0),.clk(gclk));
	jdff dff_A_BrM7y7Wq4_0(.dout(w_dff_A_MyPP7GLA4_0),.din(w_dff_A_BrM7y7Wq4_0),.clk(gclk));
	jdff dff_A_MyPP7GLA4_0(.dout(w_dff_A_5QZCV04S1_0),.din(w_dff_A_MyPP7GLA4_0),.clk(gclk));
	jdff dff_A_5QZCV04S1_0(.dout(w_dff_A_szl0iRQX2_0),.din(w_dff_A_5QZCV04S1_0),.clk(gclk));
	jdff dff_A_szl0iRQX2_0(.dout(w_dff_A_PpeJRPJC2_0),.din(w_dff_A_szl0iRQX2_0),.clk(gclk));
	jdff dff_A_PpeJRPJC2_0(.dout(w_dff_A_alQXCNca7_0),.din(w_dff_A_PpeJRPJC2_0),.clk(gclk));
	jdff dff_A_alQXCNca7_0(.dout(w_dff_A_qpNJ4XxK8_0),.din(w_dff_A_alQXCNca7_0),.clk(gclk));
	jdff dff_A_qpNJ4XxK8_0(.dout(w_dff_A_iltF4K2b2_0),.din(w_dff_A_qpNJ4XxK8_0),.clk(gclk));
	jdff dff_A_iltF4K2b2_0(.dout(w_dff_A_PGClOh0e2_0),.din(w_dff_A_iltF4K2b2_0),.clk(gclk));
	jdff dff_A_PGClOh0e2_0(.dout(w_dff_A_QXLh2RUm6_0),.din(w_dff_A_PGClOh0e2_0),.clk(gclk));
	jdff dff_A_QXLh2RUm6_0(.dout(w_dff_A_Y1iaUumO9_0),.din(w_dff_A_QXLh2RUm6_0),.clk(gclk));
	jdff dff_A_Y1iaUumO9_0(.dout(w_dff_A_JNrj9jQy8_0),.din(w_dff_A_Y1iaUumO9_0),.clk(gclk));
	jdff dff_A_JNrj9jQy8_0(.dout(w_dff_A_tvKswgPv6_0),.din(w_dff_A_JNrj9jQy8_0),.clk(gclk));
	jdff dff_A_tvKswgPv6_0(.dout(w_dff_A_wyNujQAN6_0),.din(w_dff_A_tvKswgPv6_0),.clk(gclk));
	jdff dff_A_wyNujQAN6_0(.dout(w_dff_A_gUc6hg5Q3_0),.din(w_dff_A_wyNujQAN6_0),.clk(gclk));
	jdff dff_A_gUc6hg5Q3_0(.dout(w_dff_A_Prsmcg8I7_0),.din(w_dff_A_gUc6hg5Q3_0),.clk(gclk));
	jdff dff_A_Prsmcg8I7_0(.dout(G414),.din(w_dff_A_Prsmcg8I7_0),.clk(gclk));
	jdff dff_A_uaKJXgnV6_1(.dout(w_dff_A_h5JBuQF76_0),.din(w_dff_A_uaKJXgnV6_1),.clk(gclk));
	jdff dff_A_h5JBuQF76_0(.dout(w_dff_A_2ZJ62Hke8_0),.din(w_dff_A_h5JBuQF76_0),.clk(gclk));
	jdff dff_A_2ZJ62Hke8_0(.dout(w_dff_A_ZNUX4UNg4_0),.din(w_dff_A_2ZJ62Hke8_0),.clk(gclk));
	jdff dff_A_ZNUX4UNg4_0(.dout(w_dff_A_WIkNu8zs2_0),.din(w_dff_A_ZNUX4UNg4_0),.clk(gclk));
	jdff dff_A_WIkNu8zs2_0(.dout(w_dff_A_rS9ARH322_0),.din(w_dff_A_WIkNu8zs2_0),.clk(gclk));
	jdff dff_A_rS9ARH322_0(.dout(w_dff_A_i0Hh5bi44_0),.din(w_dff_A_rS9ARH322_0),.clk(gclk));
	jdff dff_A_i0Hh5bi44_0(.dout(w_dff_A_3I0MAEwU7_0),.din(w_dff_A_i0Hh5bi44_0),.clk(gclk));
	jdff dff_A_3I0MAEwU7_0(.dout(w_dff_A_LwMR0Vku3_0),.din(w_dff_A_3I0MAEwU7_0),.clk(gclk));
	jdff dff_A_LwMR0Vku3_0(.dout(w_dff_A_P2s9Y6sz8_0),.din(w_dff_A_LwMR0Vku3_0),.clk(gclk));
	jdff dff_A_P2s9Y6sz8_0(.dout(w_dff_A_iWZ45yAQ5_0),.din(w_dff_A_P2s9Y6sz8_0),.clk(gclk));
	jdff dff_A_iWZ45yAQ5_0(.dout(w_dff_A_uTKPxXnP2_0),.din(w_dff_A_iWZ45yAQ5_0),.clk(gclk));
	jdff dff_A_uTKPxXnP2_0(.dout(w_dff_A_EkrwcEyk3_0),.din(w_dff_A_uTKPxXnP2_0),.clk(gclk));
	jdff dff_A_EkrwcEyk3_0(.dout(w_dff_A_K5yjHLD10_0),.din(w_dff_A_EkrwcEyk3_0),.clk(gclk));
	jdff dff_A_K5yjHLD10_0(.dout(w_dff_A_WJi3thGz1_0),.din(w_dff_A_K5yjHLD10_0),.clk(gclk));
	jdff dff_A_WJi3thGz1_0(.dout(w_dff_A_uxlGiOiS8_0),.din(w_dff_A_WJi3thGz1_0),.clk(gclk));
	jdff dff_A_uxlGiOiS8_0(.dout(w_dff_A_hUpOauQa6_0),.din(w_dff_A_uxlGiOiS8_0),.clk(gclk));
	jdff dff_A_hUpOauQa6_0(.dout(w_dff_A_PiMq0HRz4_0),.din(w_dff_A_hUpOauQa6_0),.clk(gclk));
	jdff dff_A_PiMq0HRz4_0(.dout(w_dff_A_ignETw157_0),.din(w_dff_A_PiMq0HRz4_0),.clk(gclk));
	jdff dff_A_ignETw157_0(.dout(w_dff_A_sJCbjRRJ7_0),.din(w_dff_A_ignETw157_0),.clk(gclk));
	jdff dff_A_sJCbjRRJ7_0(.dout(w_dff_A_hsKkG99B8_0),.din(w_dff_A_sJCbjRRJ7_0),.clk(gclk));
	jdff dff_A_hsKkG99B8_0(.dout(w_dff_A_iDVVtPbT9_0),.din(w_dff_A_hsKkG99B8_0),.clk(gclk));
	jdff dff_A_iDVVtPbT9_0(.dout(w_dff_A_LHAjMOk64_0),.din(w_dff_A_iDVVtPbT9_0),.clk(gclk));
	jdff dff_A_LHAjMOk64_0(.dout(w_dff_A_VIofv5Dt7_0),.din(w_dff_A_LHAjMOk64_0),.clk(gclk));
	jdff dff_A_VIofv5Dt7_0(.dout(w_dff_A_ZaDQpY7l0_0),.din(w_dff_A_VIofv5Dt7_0),.clk(gclk));
	jdff dff_A_ZaDQpY7l0_0(.dout(w_dff_A_6bOOtbGN8_0),.din(w_dff_A_ZaDQpY7l0_0),.clk(gclk));
	jdff dff_A_6bOOtbGN8_0(.dout(w_dff_A_pMyue93u8_0),.din(w_dff_A_6bOOtbGN8_0),.clk(gclk));
	jdff dff_A_pMyue93u8_0(.dout(w_dff_A_AerFbYG80_0),.din(w_dff_A_pMyue93u8_0),.clk(gclk));
	jdff dff_A_AerFbYG80_0(.dout(w_dff_A_4Eh9CV0b4_0),.din(w_dff_A_AerFbYG80_0),.clk(gclk));
	jdff dff_A_4Eh9CV0b4_0(.dout(G416),.din(w_dff_A_4Eh9CV0b4_0),.clk(gclk));
	jdff dff_A_82ekGnhb0_2(.dout(w_dff_A_mKWthDho3_0),.din(w_dff_A_82ekGnhb0_2),.clk(gclk));
	jdff dff_A_mKWthDho3_0(.dout(w_dff_A_FsWRfJGQ1_0),.din(w_dff_A_mKWthDho3_0),.clk(gclk));
	jdff dff_A_FsWRfJGQ1_0(.dout(w_dff_A_GLDRUKkP5_0),.din(w_dff_A_FsWRfJGQ1_0),.clk(gclk));
	jdff dff_A_GLDRUKkP5_0(.dout(w_dff_A_mMq5Lym85_0),.din(w_dff_A_GLDRUKkP5_0),.clk(gclk));
	jdff dff_A_mMq5Lym85_0(.dout(w_dff_A_jigFhaxh6_0),.din(w_dff_A_mMq5Lym85_0),.clk(gclk));
	jdff dff_A_jigFhaxh6_0(.dout(w_dff_A_f8nkZmKJ0_0),.din(w_dff_A_jigFhaxh6_0),.clk(gclk));
	jdff dff_A_f8nkZmKJ0_0(.dout(w_dff_A_UsT9TBU19_0),.din(w_dff_A_f8nkZmKJ0_0),.clk(gclk));
	jdff dff_A_UsT9TBU19_0(.dout(w_dff_A_3HsUEeS55_0),.din(w_dff_A_UsT9TBU19_0),.clk(gclk));
	jdff dff_A_3HsUEeS55_0(.dout(w_dff_A_UMuR8MuL9_0),.din(w_dff_A_3HsUEeS55_0),.clk(gclk));
	jdff dff_A_UMuR8MuL9_0(.dout(w_dff_A_pO8AZ6KA9_0),.din(w_dff_A_UMuR8MuL9_0),.clk(gclk));
	jdff dff_A_pO8AZ6KA9_0(.dout(G249),.din(w_dff_A_pO8AZ6KA9_0),.clk(gclk));
	jdff dff_A_ZJcOyy2e3_2(.dout(w_dff_A_COdxG20V3_0),.din(w_dff_A_ZJcOyy2e3_2),.clk(gclk));
	jdff dff_A_COdxG20V3_0(.dout(w_dff_A_143LnfCB1_0),.din(w_dff_A_COdxG20V3_0),.clk(gclk));
	jdff dff_A_143LnfCB1_0(.dout(w_dff_A_GkHFLnsU3_0),.din(w_dff_A_143LnfCB1_0),.clk(gclk));
	jdff dff_A_GkHFLnsU3_0(.dout(w_dff_A_5KTqZrHY2_0),.din(w_dff_A_GkHFLnsU3_0),.clk(gclk));
	jdff dff_A_5KTqZrHY2_0(.dout(w_dff_A_jc0uY5c56_0),.din(w_dff_A_5KTqZrHY2_0),.clk(gclk));
	jdff dff_A_jc0uY5c56_0(.dout(w_dff_A_dCB0pl8P9_0),.din(w_dff_A_jc0uY5c56_0),.clk(gclk));
	jdff dff_A_dCB0pl8P9_0(.dout(w_dff_A_Xza456590_0),.din(w_dff_A_dCB0pl8P9_0),.clk(gclk));
	jdff dff_A_Xza456590_0(.dout(w_dff_A_QxziYi5t2_0),.din(w_dff_A_Xza456590_0),.clk(gclk));
	jdff dff_A_QxziYi5t2_0(.dout(w_dff_A_yn8UVNzb7_0),.din(w_dff_A_QxziYi5t2_0),.clk(gclk));
	jdff dff_A_yn8UVNzb7_0(.dout(w_dff_A_2F7OlOpe4_0),.din(w_dff_A_yn8UVNzb7_0),.clk(gclk));
	jdff dff_A_2F7OlOpe4_0(.dout(G295),.din(w_dff_A_2F7OlOpe4_0),.clk(gclk));
	jdff dff_A_fhIVqjCk4_2(.dout(w_dff_A_NchF0ExF4_0),.din(w_dff_A_fhIVqjCk4_2),.clk(gclk));
	jdff dff_A_NchF0ExF4_0(.dout(w_dff_A_MF4fZL7G0_0),.din(w_dff_A_NchF0ExF4_0),.clk(gclk));
	jdff dff_A_MF4fZL7G0_0(.dout(w_dff_A_WEzBVKBl6_0),.din(w_dff_A_MF4fZL7G0_0),.clk(gclk));
	jdff dff_A_WEzBVKBl6_0(.dout(G324),.din(w_dff_A_WEzBVKBl6_0),.clk(gclk));
	jdff dff_A_V1fSan9U2_1(.dout(w_dff_A_Ns3mTjbj3_0),.din(w_dff_A_V1fSan9U2_1),.clk(gclk));
	jdff dff_A_Ns3mTjbj3_0(.dout(w_dff_A_bvZgs5WK5_0),.din(w_dff_A_Ns3mTjbj3_0),.clk(gclk));
	jdff dff_A_bvZgs5WK5_0(.dout(w_dff_A_wIVhEDTH4_0),.din(w_dff_A_bvZgs5WK5_0),.clk(gclk));
	jdff dff_A_wIVhEDTH4_0(.dout(w_dff_A_WyUpv4VO2_0),.din(w_dff_A_wIVhEDTH4_0),.clk(gclk));
	jdff dff_A_WyUpv4VO2_0(.dout(w_dff_A_8yYfWPyb3_0),.din(w_dff_A_WyUpv4VO2_0),.clk(gclk));
	jdff dff_A_8yYfWPyb3_0(.dout(w_dff_A_8LWQXudB1_0),.din(w_dff_A_8yYfWPyb3_0),.clk(gclk));
	jdff dff_A_8LWQXudB1_0(.dout(w_dff_A_L4X1tgIA8_0),.din(w_dff_A_8LWQXudB1_0),.clk(gclk));
	jdff dff_A_L4X1tgIA8_0(.dout(w_dff_A_1LZTMBJY8_0),.din(w_dff_A_L4X1tgIA8_0),.clk(gclk));
	jdff dff_A_1LZTMBJY8_0(.dout(w_dff_A_TxdXcCOk2_0),.din(w_dff_A_1LZTMBJY8_0),.clk(gclk));
	jdff dff_A_TxdXcCOk2_0(.dout(w_dff_A_on29UYq85_0),.din(w_dff_A_TxdXcCOk2_0),.clk(gclk));
	jdff dff_A_on29UYq85_0(.dout(w_dff_A_2IKsu5tu1_0),.din(w_dff_A_on29UYq85_0),.clk(gclk));
	jdff dff_A_2IKsu5tu1_0(.dout(w_dff_A_JCARljA63_0),.din(w_dff_A_2IKsu5tu1_0),.clk(gclk));
	jdff dff_A_JCARljA63_0(.dout(w_dff_A_W2uEw8W79_0),.din(w_dff_A_JCARljA63_0),.clk(gclk));
	jdff dff_A_W2uEw8W79_0(.dout(w_dff_A_5ijsCaKo7_0),.din(w_dff_A_W2uEw8W79_0),.clk(gclk));
	jdff dff_A_5ijsCaKo7_0(.dout(w_dff_A_yVOnFs1x9_0),.din(w_dff_A_5ijsCaKo7_0),.clk(gclk));
	jdff dff_A_yVOnFs1x9_0(.dout(w_dff_A_eoMt9YBF5_0),.din(w_dff_A_yVOnFs1x9_0),.clk(gclk));
	jdff dff_A_eoMt9YBF5_0(.dout(w_dff_A_62aXicn74_0),.din(w_dff_A_eoMt9YBF5_0),.clk(gclk));
	jdff dff_A_62aXicn74_0(.dout(w_dff_A_3y16qGmv6_0),.din(w_dff_A_62aXicn74_0),.clk(gclk));
	jdff dff_A_3y16qGmv6_0(.dout(w_dff_A_lBVvOCYB5_0),.din(w_dff_A_3y16qGmv6_0),.clk(gclk));
	jdff dff_A_lBVvOCYB5_0(.dout(w_dff_A_MXthOtod9_0),.din(w_dff_A_lBVvOCYB5_0),.clk(gclk));
	jdff dff_A_MXthOtod9_0(.dout(G252),.din(w_dff_A_MXthOtod9_0),.clk(gclk));
	jdff dff_A_GCOhVMYb7_2(.dout(w_dff_A_N3V3GSHY4_0),.din(w_dff_A_GCOhVMYb7_2),.clk(gclk));
	jdff dff_A_N3V3GSHY4_0(.dout(w_dff_A_WheD8US29_0),.din(w_dff_A_N3V3GSHY4_0),.clk(gclk));
	jdff dff_A_WheD8US29_0(.dout(w_dff_A_mzqW7H6v3_0),.din(w_dff_A_WheD8US29_0),.clk(gclk));
	jdff dff_A_mzqW7H6v3_0(.dout(w_dff_A_fn9tgkcG9_0),.din(w_dff_A_mzqW7H6v3_0),.clk(gclk));
	jdff dff_A_fn9tgkcG9_0(.dout(w_dff_A_OoLH6zQG7_0),.din(w_dff_A_fn9tgkcG9_0),.clk(gclk));
	jdff dff_A_OoLH6zQG7_0(.dout(G310),.din(w_dff_A_OoLH6zQG7_0),.clk(gclk));
	jdff dff_A_bWmbwUsV7_2(.dout(w_dff_A_fEr1VKOp6_0),.din(w_dff_A_bWmbwUsV7_2),.clk(gclk));
	jdff dff_A_fEr1VKOp6_0(.dout(w_dff_A_XgVXNhuH4_0),.din(w_dff_A_fEr1VKOp6_0),.clk(gclk));
	jdff dff_A_XgVXNhuH4_0(.dout(w_dff_A_QMRmzlLC3_0),.din(w_dff_A_XgVXNhuH4_0),.clk(gclk));
	jdff dff_A_QMRmzlLC3_0(.dout(w_dff_A_LTETGmhr2_0),.din(w_dff_A_QMRmzlLC3_0),.clk(gclk));
	jdff dff_A_LTETGmhr2_0(.dout(G313),.din(w_dff_A_LTETGmhr2_0),.clk(gclk));
	jdff dff_A_Zs4DPBih4_2(.dout(w_dff_A_7yna31FM6_0),.din(w_dff_A_Zs4DPBih4_2),.clk(gclk));
	jdff dff_A_7yna31FM6_0(.dout(w_dff_A_Epkq8GxI7_0),.din(w_dff_A_7yna31FM6_0),.clk(gclk));
	jdff dff_A_Epkq8GxI7_0(.dout(w_dff_A_j3fxXw7N2_0),.din(w_dff_A_Epkq8GxI7_0),.clk(gclk));
	jdff dff_A_j3fxXw7N2_0(.dout(w_dff_A_mNPRPVNR2_0),.din(w_dff_A_j3fxXw7N2_0),.clk(gclk));
	jdff dff_A_mNPRPVNR2_0(.dout(w_dff_A_d3U8Z1yA2_0),.din(w_dff_A_mNPRPVNR2_0),.clk(gclk));
	jdff dff_A_d3U8Z1yA2_0(.dout(w_dff_A_8O4ZoJvT0_0),.din(w_dff_A_d3U8Z1yA2_0),.clk(gclk));
	jdff dff_A_8O4ZoJvT0_0(.dout(w_dff_A_b15N8rKA5_0),.din(w_dff_A_8O4ZoJvT0_0),.clk(gclk));
	jdff dff_A_b15N8rKA5_0(.dout(w_dff_A_uF1Aix0e0_0),.din(w_dff_A_b15N8rKA5_0),.clk(gclk));
	jdff dff_A_uF1Aix0e0_0(.dout(G316),.din(w_dff_A_uF1Aix0e0_0),.clk(gclk));
	jdff dff_A_A2Ayl1W59_2(.dout(w_dff_A_6QfHv3ah8_0),.din(w_dff_A_A2Ayl1W59_2),.clk(gclk));
	jdff dff_A_6QfHv3ah8_0(.dout(w_dff_A_t4yerWQ56_0),.din(w_dff_A_6QfHv3ah8_0),.clk(gclk));
	jdff dff_A_t4yerWQ56_0(.dout(w_dff_A_k8SIRAVT3_0),.din(w_dff_A_t4yerWQ56_0),.clk(gclk));
	jdff dff_A_k8SIRAVT3_0(.dout(w_dff_A_mWHsMMDK2_0),.din(w_dff_A_k8SIRAVT3_0),.clk(gclk));
	jdff dff_A_mWHsMMDK2_0(.dout(w_dff_A_B914WQtK6_0),.din(w_dff_A_mWHsMMDK2_0),.clk(gclk));
	jdff dff_A_B914WQtK6_0(.dout(w_dff_A_Thea6Efg8_0),.din(w_dff_A_B914WQtK6_0),.clk(gclk));
	jdff dff_A_Thea6Efg8_0(.dout(w_dff_A_9GdNTB9o9_0),.din(w_dff_A_Thea6Efg8_0),.clk(gclk));
	jdff dff_A_9GdNTB9o9_0(.dout(w_dff_A_JEMRoawf2_0),.din(w_dff_A_9GdNTB9o9_0),.clk(gclk));
	jdff dff_A_JEMRoawf2_0(.dout(G319),.din(w_dff_A_JEMRoawf2_0),.clk(gclk));
	jdff dff_A_Di2h08h34_2(.dout(w_dff_A_cGtTuxfP2_0),.din(w_dff_A_Di2h08h34_2),.clk(gclk));
	jdff dff_A_cGtTuxfP2_0(.dout(G327),.din(w_dff_A_cGtTuxfP2_0),.clk(gclk));
	jdff dff_A_mrhQvpES1_2(.dout(w_dff_A_zDkIfLAq2_0),.din(w_dff_A_mrhQvpES1_2),.clk(gclk));
	jdff dff_A_zDkIfLAq2_0(.dout(G330),.din(w_dff_A_zDkIfLAq2_0),.clk(gclk));
	jdff dff_A_iQ4quPVT4_2(.dout(w_dff_A_awmdFMC91_0),.din(w_dff_A_iQ4quPVT4_2),.clk(gclk));
	jdff dff_A_awmdFMC91_0(.dout(G336),.din(w_dff_A_awmdFMC91_0),.clk(gclk));
	jdff dff_A_bYZjOR4l8_2(.dout(w_dff_A_Sg8h2GHg4_0),.din(w_dff_A_bYZjOR4l8_2),.clk(gclk));
	jdff dff_A_Sg8h2GHg4_0(.dout(w_dff_A_xodhc1gd3_0),.din(w_dff_A_Sg8h2GHg4_0),.clk(gclk));
	jdff dff_A_xodhc1gd3_0(.dout(w_dff_A_zhCzkvGB9_0),.din(w_dff_A_xodhc1gd3_0),.clk(gclk));
	jdff dff_A_zhCzkvGB9_0(.dout(w_dff_A_4Rt6owKt7_0),.din(w_dff_A_zhCzkvGB9_0),.clk(gclk));
	jdff dff_A_4Rt6owKt7_0(.dout(w_dff_A_v9kVG2yQ4_0),.din(w_dff_A_4Rt6owKt7_0),.clk(gclk));
	jdff dff_A_v9kVG2yQ4_0(.dout(w_dff_A_XgARWpSg8_0),.din(w_dff_A_v9kVG2yQ4_0),.clk(gclk));
	jdff dff_A_XgARWpSg8_0(.dout(w_dff_A_YMDJDxIo4_0),.din(w_dff_A_XgARWpSg8_0),.clk(gclk));
	jdff dff_A_YMDJDxIo4_0(.dout(w_dff_A_0mQReEc72_0),.din(w_dff_A_YMDJDxIo4_0),.clk(gclk));
	jdff dff_A_0mQReEc72_0(.dout(w_dff_A_9SM2rFlR4_0),.din(w_dff_A_0mQReEc72_0),.clk(gclk));
	jdff dff_A_9SM2rFlR4_0(.dout(w_dff_A_QWXKn5Ug5_0),.din(w_dff_A_9SM2rFlR4_0),.clk(gclk));
	jdff dff_A_QWXKn5Ug5_0(.dout(w_dff_A_s8pf0N6O3_0),.din(w_dff_A_QWXKn5Ug5_0),.clk(gclk));
	jdff dff_A_s8pf0N6O3_0(.dout(w_dff_A_DRWXHmrG5_0),.din(w_dff_A_s8pf0N6O3_0),.clk(gclk));
	jdff dff_A_DRWXHmrG5_0(.dout(w_dff_A_2lVtROAw7_0),.din(w_dff_A_DRWXHmrG5_0),.clk(gclk));
	jdff dff_A_2lVtROAw7_0(.dout(w_dff_A_ut142qF65_0),.din(w_dff_A_2lVtROAw7_0),.clk(gclk));
	jdff dff_A_ut142qF65_0(.dout(w_dff_A_Kf58cNfz8_0),.din(w_dff_A_ut142qF65_0),.clk(gclk));
	jdff dff_A_Kf58cNfz8_0(.dout(w_dff_A_aPeUoKoA8_0),.din(w_dff_A_Kf58cNfz8_0),.clk(gclk));
	jdff dff_A_aPeUoKoA8_0(.dout(w_dff_A_SEuCHR110_0),.din(w_dff_A_aPeUoKoA8_0),.clk(gclk));
	jdff dff_A_SEuCHR110_0(.dout(w_dff_A_0APREGL63_0),.din(w_dff_A_SEuCHR110_0),.clk(gclk));
	jdff dff_A_0APREGL63_0(.dout(w_dff_A_4unxHd6X7_0),.din(w_dff_A_0APREGL63_0),.clk(gclk));
	jdff dff_A_4unxHd6X7_0(.dout(w_dff_A_fpSu00BN5_0),.din(w_dff_A_4unxHd6X7_0),.clk(gclk));
	jdff dff_A_fpSu00BN5_0(.dout(w_dff_A_VsyDl8U20_0),.din(w_dff_A_fpSu00BN5_0),.clk(gclk));
	jdff dff_A_VsyDl8U20_0(.dout(w_dff_A_aMAuTsPq4_0),.din(w_dff_A_VsyDl8U20_0),.clk(gclk));
	jdff dff_A_aMAuTsPq4_0(.dout(w_dff_A_pU2kcv4h2_0),.din(w_dff_A_aMAuTsPq4_0),.clk(gclk));
	jdff dff_A_pU2kcv4h2_0(.dout(w_dff_A_HbeBnZqG9_0),.din(w_dff_A_pU2kcv4h2_0),.clk(gclk));
	jdff dff_A_HbeBnZqG9_0(.dout(G418),.din(w_dff_A_HbeBnZqG9_0),.clk(gclk));
	jdff dff_A_xYcOwCKE4_2(.dout(w_dff_A_lp4BZ3Ra3_0),.din(w_dff_A_xYcOwCKE4_2),.clk(gclk));
	jdff dff_A_lp4BZ3Ra3_0(.dout(w_dff_A_MNWCFF3m6_0),.din(w_dff_A_lp4BZ3Ra3_0),.clk(gclk));
	jdff dff_A_MNWCFF3m6_0(.dout(w_dff_A_S8kL1AYv6_0),.din(w_dff_A_MNWCFF3m6_0),.clk(gclk));
	jdff dff_A_S8kL1AYv6_0(.dout(w_dff_A_9QEweryx9_0),.din(w_dff_A_S8kL1AYv6_0),.clk(gclk));
	jdff dff_A_9QEweryx9_0(.dout(w_dff_A_cWJs2vos8_0),.din(w_dff_A_9QEweryx9_0),.clk(gclk));
	jdff dff_A_cWJs2vos8_0(.dout(G298),.din(w_dff_A_cWJs2vos8_0),.clk(gclk));
	jdff dff_A_DKHFtTxw2_2(.dout(w_dff_A_GYaUbAuZ3_0),.din(w_dff_A_DKHFtTxw2_2),.clk(gclk));
	jdff dff_A_GYaUbAuZ3_0(.dout(w_dff_A_5z2Rx1GY8_0),.din(w_dff_A_GYaUbAuZ3_0),.clk(gclk));
	jdff dff_A_5z2Rx1GY8_0(.dout(w_dff_A_v62LrHl38_0),.din(w_dff_A_5z2Rx1GY8_0),.clk(gclk));
	jdff dff_A_v62LrHl38_0(.dout(w_dff_A_o6GMIi889_0),.din(w_dff_A_v62LrHl38_0),.clk(gclk));
	jdff dff_A_o6GMIi889_0(.dout(w_dff_A_FFhDPAqN4_0),.din(w_dff_A_o6GMIi889_0),.clk(gclk));
	jdff dff_A_FFhDPAqN4_0(.dout(G301),.din(w_dff_A_FFhDPAqN4_0),.clk(gclk));
	jdff dff_A_xHBLP3f76_2(.dout(w_dff_A_AcBhlfou6_0),.din(w_dff_A_xHBLP3f76_2),.clk(gclk));
	jdff dff_A_AcBhlfou6_0(.dout(w_dff_A_ftPGgdGO7_0),.din(w_dff_A_AcBhlfou6_0),.clk(gclk));
	jdff dff_A_ftPGgdGO7_0(.dout(w_dff_A_Vd1u5Ds90_0),.din(w_dff_A_ftPGgdGO7_0),.clk(gclk));
	jdff dff_A_Vd1u5Ds90_0(.dout(w_dff_A_WUj3Bhz24_0),.din(w_dff_A_Vd1u5Ds90_0),.clk(gclk));
	jdff dff_A_WUj3Bhz24_0(.dout(w_dff_A_5FgrVi0f7_0),.din(w_dff_A_WUj3Bhz24_0),.clk(gclk));
	jdff dff_A_5FgrVi0f7_0(.dout(G304),.din(w_dff_A_5FgrVi0f7_0),.clk(gclk));
	jdff dff_A_kmbXyAx51_2(.dout(w_dff_A_6Xe8z1hJ0_0),.din(w_dff_A_kmbXyAx51_2),.clk(gclk));
	jdff dff_A_6Xe8z1hJ0_0(.dout(w_dff_A_k7mUY3ae4_0),.din(w_dff_A_6Xe8z1hJ0_0),.clk(gclk));
	jdff dff_A_k7mUY3ae4_0(.dout(w_dff_A_gyjqWEac6_0),.din(w_dff_A_k7mUY3ae4_0),.clk(gclk));
	jdff dff_A_gyjqWEac6_0(.dout(w_dff_A_n2xGXPLM7_0),.din(w_dff_A_gyjqWEac6_0),.clk(gclk));
	jdff dff_A_n2xGXPLM7_0(.dout(w_dff_A_RAwpjRFA3_0),.din(w_dff_A_n2xGXPLM7_0),.clk(gclk));
	jdff dff_A_RAwpjRFA3_0(.dout(w_dff_A_KCAQtB6M2_0),.din(w_dff_A_RAwpjRFA3_0),.clk(gclk));
	jdff dff_A_KCAQtB6M2_0(.dout(w_dff_A_CNeCHZog3_0),.din(w_dff_A_KCAQtB6M2_0),.clk(gclk));
	jdff dff_A_CNeCHZog3_0(.dout(G307),.din(w_dff_A_CNeCHZog3_0),.clk(gclk));
	jdff dff_A_g9igXi8t2_2(.dout(w_dff_A_QWF5MNSI7_0),.din(w_dff_A_g9igXi8t2_2),.clk(gclk));
	jdff dff_A_QWF5MNSI7_0(.dout(w_dff_A_JiJS0Jb39_0),.din(w_dff_A_QWF5MNSI7_0),.clk(gclk));
	jdff dff_A_JiJS0Jb39_0(.dout(w_dff_A_QvmVZT986_0),.din(w_dff_A_JiJS0Jb39_0),.clk(gclk));
	jdff dff_A_QvmVZT986_0(.dout(w_dff_A_YT14wwP74_0),.din(w_dff_A_QvmVZT986_0),.clk(gclk));
	jdff dff_A_YT14wwP74_0(.dout(w_dff_A_reEqvgj73_0),.din(w_dff_A_YT14wwP74_0),.clk(gclk));
	jdff dff_A_reEqvgj73_0(.dout(w_dff_A_4lwNbUNa5_0),.din(w_dff_A_reEqvgj73_0),.clk(gclk));
	jdff dff_A_4lwNbUNa5_0(.dout(w_dff_A_7YGOf3Tg3_0),.din(w_dff_A_4lwNbUNa5_0),.clk(gclk));
	jdff dff_A_7YGOf3Tg3_0(.dout(w_dff_A_Q3YppFAk3_0),.din(w_dff_A_7YGOf3Tg3_0),.clk(gclk));
	jdff dff_A_Q3YppFAk3_0(.dout(w_dff_A_guZB8wGF9_0),.din(w_dff_A_Q3YppFAk3_0),.clk(gclk));
	jdff dff_A_guZB8wGF9_0(.dout(w_dff_A_22TNwHTZ8_0),.din(w_dff_A_guZB8wGF9_0),.clk(gclk));
	jdff dff_A_22TNwHTZ8_0(.dout(w_dff_A_dz8hkwqB1_0),.din(w_dff_A_22TNwHTZ8_0),.clk(gclk));
	jdff dff_A_dz8hkwqB1_0(.dout(w_dff_A_mDA0UIXU1_0),.din(w_dff_A_dz8hkwqB1_0),.clk(gclk));
	jdff dff_A_mDA0UIXU1_0(.dout(w_dff_A_OrLuNpyR6_0),.din(w_dff_A_mDA0UIXU1_0),.clk(gclk));
	jdff dff_A_OrLuNpyR6_0(.dout(w_dff_A_7PDWFlxK6_0),.din(w_dff_A_OrLuNpyR6_0),.clk(gclk));
	jdff dff_A_7PDWFlxK6_0(.dout(w_dff_A_sizJU5Kv2_0),.din(w_dff_A_7PDWFlxK6_0),.clk(gclk));
	jdff dff_A_sizJU5Kv2_0(.dout(w_dff_A_w8OodaHw7_0),.din(w_dff_A_sizJU5Kv2_0),.clk(gclk));
	jdff dff_A_w8OodaHw7_0(.dout(w_dff_A_bNDGyu6c7_0),.din(w_dff_A_w8OodaHw7_0),.clk(gclk));
	jdff dff_A_bNDGyu6c7_0(.dout(w_dff_A_TGOisIUX3_0),.din(w_dff_A_bNDGyu6c7_0),.clk(gclk));
	jdff dff_A_TGOisIUX3_0(.dout(w_dff_A_CsRxIJfP3_0),.din(w_dff_A_TGOisIUX3_0),.clk(gclk));
	jdff dff_A_CsRxIJfP3_0(.dout(G344),.din(w_dff_A_CsRxIJfP3_0),.clk(gclk));
	jdff dff_A_DGJTufCb5_2(.dout(w_dff_A_4jJHDijp6_0),.din(w_dff_A_DGJTufCb5_2),.clk(gclk));
	jdff dff_A_4jJHDijp6_0(.dout(G419),.din(w_dff_A_4jJHDijp6_0),.clk(gclk));
	jdff dff_A_RDG8Zhod6_2(.dout(w_dff_A_7lbDtceC0_0),.din(w_dff_A_RDG8Zhod6_2),.clk(gclk));
	jdff dff_A_7lbDtceC0_0(.dout(G471),.din(w_dff_A_7lbDtceC0_0),.clk(gclk));
	jdff dff_A_Snttc1Yu1_2(.dout(w_dff_A_j4qyzTbw6_0),.din(w_dff_A_Snttc1Yu1_2),.clk(gclk));
	jdff dff_A_j4qyzTbw6_0(.dout(w_dff_A_zInl2alh1_0),.din(w_dff_A_j4qyzTbw6_0),.clk(gclk));
	jdff dff_A_zInl2alh1_0(.dout(w_dff_A_t3ajAGXb6_0),.din(w_dff_A_zInl2alh1_0),.clk(gclk));
	jdff dff_A_t3ajAGXb6_0(.dout(w_dff_A_2MmhuD854_0),.din(w_dff_A_t3ajAGXb6_0),.clk(gclk));
	jdff dff_A_2MmhuD854_0(.dout(w_dff_A_WSPM8UuE1_0),.din(w_dff_A_2MmhuD854_0),.clk(gclk));
	jdff dff_A_WSPM8UuE1_0(.dout(w_dff_A_ffCIwah64_0),.din(w_dff_A_WSPM8UuE1_0),.clk(gclk));
	jdff dff_A_ffCIwah64_0(.dout(w_dff_A_M1ogNM1q4_0),.din(w_dff_A_ffCIwah64_0),.clk(gclk));
	jdff dff_A_M1ogNM1q4_0(.dout(w_dff_A_wvPK4jcW6_0),.din(w_dff_A_M1ogNM1q4_0),.clk(gclk));
	jdff dff_A_wvPK4jcW6_0(.dout(w_dff_A_Ay7YtLpr7_0),.din(w_dff_A_wvPK4jcW6_0),.clk(gclk));
	jdff dff_A_Ay7YtLpr7_0(.dout(w_dff_A_n09qDzQp9_0),.din(w_dff_A_Ay7YtLpr7_0),.clk(gclk));
	jdff dff_A_n09qDzQp9_0(.dout(w_dff_A_cFBNnqgR7_0),.din(w_dff_A_n09qDzQp9_0),.clk(gclk));
	jdff dff_A_cFBNnqgR7_0(.dout(w_dff_A_BqNKQ9v92_0),.din(w_dff_A_cFBNnqgR7_0),.clk(gclk));
	jdff dff_A_BqNKQ9v92_0(.dout(w_dff_A_NTodMKiG3_0),.din(w_dff_A_BqNKQ9v92_0),.clk(gclk));
	jdff dff_A_NTodMKiG3_0(.dout(w_dff_A_PP7ucWkp5_0),.din(w_dff_A_NTodMKiG3_0),.clk(gclk));
	jdff dff_A_PP7ucWkp5_0(.dout(w_dff_A_1ZcJDa6n1_0),.din(w_dff_A_PP7ucWkp5_0),.clk(gclk));
	jdff dff_A_1ZcJDa6n1_0(.dout(w_dff_A_8bC3HfEN8_0),.din(w_dff_A_1ZcJDa6n1_0),.clk(gclk));
	jdff dff_A_8bC3HfEN8_0(.dout(w_dff_A_iJoqc8sB5_0),.din(w_dff_A_8bC3HfEN8_0),.clk(gclk));
	jdff dff_A_iJoqc8sB5_0(.dout(G359),.din(w_dff_A_iJoqc8sB5_0),.clk(gclk));
	jdff dff_A_T4PMdRc97_2(.dout(w_dff_A_TKO326SN7_0),.din(w_dff_A_T4PMdRc97_2),.clk(gclk));
	jdff dff_A_TKO326SN7_0(.dout(w_dff_A_PKXtIPsC3_0),.din(w_dff_A_TKO326SN7_0),.clk(gclk));
	jdff dff_A_PKXtIPsC3_0(.dout(w_dff_A_UMRMhsY89_0),.din(w_dff_A_PKXtIPsC3_0),.clk(gclk));
	jdff dff_A_UMRMhsY89_0(.dout(w_dff_A_Yh1FBwUM8_0),.din(w_dff_A_UMRMhsY89_0),.clk(gclk));
	jdff dff_A_Yh1FBwUM8_0(.dout(w_dff_A_Z3HXBjD97_0),.din(w_dff_A_Yh1FBwUM8_0),.clk(gclk));
	jdff dff_A_Z3HXBjD97_0(.dout(w_dff_A_vDcxGj9e0_0),.din(w_dff_A_Z3HXBjD97_0),.clk(gclk));
	jdff dff_A_vDcxGj9e0_0(.dout(w_dff_A_KTcEJu3D9_0),.din(w_dff_A_vDcxGj9e0_0),.clk(gclk));
	jdff dff_A_KTcEJu3D9_0(.dout(w_dff_A_iDMvqfhM1_0),.din(w_dff_A_KTcEJu3D9_0),.clk(gclk));
	jdff dff_A_iDMvqfhM1_0(.dout(w_dff_A_k7cGj2179_0),.din(w_dff_A_iDMvqfhM1_0),.clk(gclk));
	jdff dff_A_k7cGj2179_0(.dout(w_dff_A_dRvmNNQ72_0),.din(w_dff_A_k7cGj2179_0),.clk(gclk));
	jdff dff_A_dRvmNNQ72_0(.dout(w_dff_A_YJfnu9sG4_0),.din(w_dff_A_dRvmNNQ72_0),.clk(gclk));
	jdff dff_A_YJfnu9sG4_0(.dout(w_dff_A_R1B35dN19_0),.din(w_dff_A_YJfnu9sG4_0),.clk(gclk));
	jdff dff_A_R1B35dN19_0(.dout(w_dff_A_Abow7xoR7_0),.din(w_dff_A_R1B35dN19_0),.clk(gclk));
	jdff dff_A_Abow7xoR7_0(.dout(w_dff_A_qP62sMNU0_0),.din(w_dff_A_Abow7xoR7_0),.clk(gclk));
	jdff dff_A_qP62sMNU0_0(.dout(w_dff_A_iy0AUKON6_0),.din(w_dff_A_qP62sMNU0_0),.clk(gclk));
	jdff dff_A_iy0AUKON6_0(.dout(w_dff_A_LXYKvGO26_0),.din(w_dff_A_iy0AUKON6_0),.clk(gclk));
	jdff dff_A_LXYKvGO26_0(.dout(w_dff_A_zt3cnxgn0_0),.din(w_dff_A_LXYKvGO26_0),.clk(gclk));
	jdff dff_A_zt3cnxgn0_0(.dout(G362),.din(w_dff_A_zt3cnxgn0_0),.clk(gclk));
	jdff dff_A_B7P868BX1_2(.dout(w_dff_A_twqNrC4O3_0),.din(w_dff_A_B7P868BX1_2),.clk(gclk));
	jdff dff_A_twqNrC4O3_0(.dout(w_dff_A_r2E4A33R4_0),.din(w_dff_A_twqNrC4O3_0),.clk(gclk));
	jdff dff_A_r2E4A33R4_0(.dout(w_dff_A_eimFmXYt7_0),.din(w_dff_A_r2E4A33R4_0),.clk(gclk));
	jdff dff_A_eimFmXYt7_0(.dout(w_dff_A_VKBRRyAn1_0),.din(w_dff_A_eimFmXYt7_0),.clk(gclk));
	jdff dff_A_VKBRRyAn1_0(.dout(w_dff_A_puVLSrGL2_0),.din(w_dff_A_VKBRRyAn1_0),.clk(gclk));
	jdff dff_A_puVLSrGL2_0(.dout(w_dff_A_z9J559Ir9_0),.din(w_dff_A_puVLSrGL2_0),.clk(gclk));
	jdff dff_A_z9J559Ir9_0(.dout(w_dff_A_2Rw37lrH3_0),.din(w_dff_A_z9J559Ir9_0),.clk(gclk));
	jdff dff_A_2Rw37lrH3_0(.dout(w_dff_A_ATgClKxn7_0),.din(w_dff_A_2Rw37lrH3_0),.clk(gclk));
	jdff dff_A_ATgClKxn7_0(.dout(w_dff_A_yzPcVvkx7_0),.din(w_dff_A_ATgClKxn7_0),.clk(gclk));
	jdff dff_A_yzPcVvkx7_0(.dout(w_dff_A_RvmMBtZn8_0),.din(w_dff_A_yzPcVvkx7_0),.clk(gclk));
	jdff dff_A_RvmMBtZn8_0(.dout(w_dff_A_YXZXptmH8_0),.din(w_dff_A_RvmMBtZn8_0),.clk(gclk));
	jdff dff_A_YXZXptmH8_0(.dout(w_dff_A_qXK4AFGg4_0),.din(w_dff_A_YXZXptmH8_0),.clk(gclk));
	jdff dff_A_qXK4AFGg4_0(.dout(w_dff_A_UJlvFUtW7_0),.din(w_dff_A_qXK4AFGg4_0),.clk(gclk));
	jdff dff_A_UJlvFUtW7_0(.dout(w_dff_A_MSYfMvN65_0),.din(w_dff_A_UJlvFUtW7_0),.clk(gclk));
	jdff dff_A_MSYfMvN65_0(.dout(w_dff_A_d14eUvhp3_0),.din(w_dff_A_MSYfMvN65_0),.clk(gclk));
	jdff dff_A_d14eUvhp3_0(.dout(w_dff_A_2PjQjbGr0_0),.din(w_dff_A_d14eUvhp3_0),.clk(gclk));
	jdff dff_A_2PjQjbGr0_0(.dout(w_dff_A_JRksjT0Y4_0),.din(w_dff_A_2PjQjbGr0_0),.clk(gclk));
	jdff dff_A_JRksjT0Y4_0(.dout(G365),.din(w_dff_A_JRksjT0Y4_0),.clk(gclk));
	jdff dff_A_eHl8FGiB3_2(.dout(w_dff_A_ymbhNT8k6_0),.din(w_dff_A_eHl8FGiB3_2),.clk(gclk));
	jdff dff_A_ymbhNT8k6_0(.dout(w_dff_A_mGxwTEWz5_0),.din(w_dff_A_ymbhNT8k6_0),.clk(gclk));
	jdff dff_A_mGxwTEWz5_0(.dout(w_dff_A_9CU3jchR9_0),.din(w_dff_A_mGxwTEWz5_0),.clk(gclk));
	jdff dff_A_9CU3jchR9_0(.dout(w_dff_A_pClrmOfj1_0),.din(w_dff_A_9CU3jchR9_0),.clk(gclk));
	jdff dff_A_pClrmOfj1_0(.dout(w_dff_A_KUfJE5t25_0),.din(w_dff_A_pClrmOfj1_0),.clk(gclk));
	jdff dff_A_KUfJE5t25_0(.dout(w_dff_A_sfMyqbEA3_0),.din(w_dff_A_KUfJE5t25_0),.clk(gclk));
	jdff dff_A_sfMyqbEA3_0(.dout(w_dff_A_hr863h1V0_0),.din(w_dff_A_sfMyqbEA3_0),.clk(gclk));
	jdff dff_A_hr863h1V0_0(.dout(w_dff_A_6owKjLva0_0),.din(w_dff_A_hr863h1V0_0),.clk(gclk));
	jdff dff_A_6owKjLva0_0(.dout(w_dff_A_86LP1u9I2_0),.din(w_dff_A_6owKjLva0_0),.clk(gclk));
	jdff dff_A_86LP1u9I2_0(.dout(w_dff_A_qmNOK5M19_0),.din(w_dff_A_86LP1u9I2_0),.clk(gclk));
	jdff dff_A_qmNOK5M19_0(.dout(w_dff_A_kYOh8TQN1_0),.din(w_dff_A_qmNOK5M19_0),.clk(gclk));
	jdff dff_A_kYOh8TQN1_0(.dout(w_dff_A_3V49KIAp6_0),.din(w_dff_A_kYOh8TQN1_0),.clk(gclk));
	jdff dff_A_3V49KIAp6_0(.dout(w_dff_A_OFiyNJQp4_0),.din(w_dff_A_3V49KIAp6_0),.clk(gclk));
	jdff dff_A_OFiyNJQp4_0(.dout(w_dff_A_x1IFlwdf7_0),.din(w_dff_A_OFiyNJQp4_0),.clk(gclk));
	jdff dff_A_x1IFlwdf7_0(.dout(w_dff_A_9Qe4mkAm0_0),.din(w_dff_A_x1IFlwdf7_0),.clk(gclk));
	jdff dff_A_9Qe4mkAm0_0(.dout(w_dff_A_SAGprpq54_0),.din(w_dff_A_9Qe4mkAm0_0),.clk(gclk));
	jdff dff_A_SAGprpq54_0(.dout(w_dff_A_CTqnyzxH1_0),.din(w_dff_A_SAGprpq54_0),.clk(gclk));
	jdff dff_A_CTqnyzxH1_0(.dout(G368),.din(w_dff_A_CTqnyzxH1_0),.clk(gclk));
	jdff dff_A_5mhHFufl9_2(.dout(w_dff_A_19WJnn0R1_0),.din(w_dff_A_5mhHFufl9_2),.clk(gclk));
	jdff dff_A_19WJnn0R1_0(.dout(w_dff_A_duRybRl99_0),.din(w_dff_A_19WJnn0R1_0),.clk(gclk));
	jdff dff_A_duRybRl99_0(.dout(w_dff_A_SLFzaVaZ8_0),.din(w_dff_A_duRybRl99_0),.clk(gclk));
	jdff dff_A_SLFzaVaZ8_0(.dout(w_dff_A_aZmbzrCo5_0),.din(w_dff_A_SLFzaVaZ8_0),.clk(gclk));
	jdff dff_A_aZmbzrCo5_0(.dout(w_dff_A_LJOtiIoB9_0),.din(w_dff_A_aZmbzrCo5_0),.clk(gclk));
	jdff dff_A_LJOtiIoB9_0(.dout(w_dff_A_GgEsdxbu5_0),.din(w_dff_A_LJOtiIoB9_0),.clk(gclk));
	jdff dff_A_GgEsdxbu5_0(.dout(w_dff_A_BiWMoxcW3_0),.din(w_dff_A_GgEsdxbu5_0),.clk(gclk));
	jdff dff_A_BiWMoxcW3_0(.dout(w_dff_A_l5BLak9X0_0),.din(w_dff_A_BiWMoxcW3_0),.clk(gclk));
	jdff dff_A_l5BLak9X0_0(.dout(w_dff_A_XIjrMCKd7_0),.din(w_dff_A_l5BLak9X0_0),.clk(gclk));
	jdff dff_A_XIjrMCKd7_0(.dout(w_dff_A_4OEcOAsP4_0),.din(w_dff_A_XIjrMCKd7_0),.clk(gclk));
	jdff dff_A_4OEcOAsP4_0(.dout(w_dff_A_tSCJWxxE3_0),.din(w_dff_A_4OEcOAsP4_0),.clk(gclk));
	jdff dff_A_tSCJWxxE3_0(.dout(w_dff_A_Yj5j4oGV8_0),.din(w_dff_A_tSCJWxxE3_0),.clk(gclk));
	jdff dff_A_Yj5j4oGV8_0(.dout(G347),.din(w_dff_A_Yj5j4oGV8_0),.clk(gclk));
	jdff dff_A_xY7oVWid9_2(.dout(w_dff_A_H7Bpe8DN4_0),.din(w_dff_A_xY7oVWid9_2),.clk(gclk));
	jdff dff_A_H7Bpe8DN4_0(.dout(w_dff_A_0aNFDEvN2_0),.din(w_dff_A_H7Bpe8DN4_0),.clk(gclk));
	jdff dff_A_0aNFDEvN2_0(.dout(w_dff_A_KFanRTyL6_0),.din(w_dff_A_0aNFDEvN2_0),.clk(gclk));
	jdff dff_A_KFanRTyL6_0(.dout(w_dff_A_yNWv5jkV2_0),.din(w_dff_A_KFanRTyL6_0),.clk(gclk));
	jdff dff_A_yNWv5jkV2_0(.dout(w_dff_A_hieiPy7B8_0),.din(w_dff_A_yNWv5jkV2_0),.clk(gclk));
	jdff dff_A_hieiPy7B8_0(.dout(w_dff_A_D2G9Ea7L4_0),.din(w_dff_A_hieiPy7B8_0),.clk(gclk));
	jdff dff_A_D2G9Ea7L4_0(.dout(w_dff_A_oykV85p26_0),.din(w_dff_A_D2G9Ea7L4_0),.clk(gclk));
	jdff dff_A_oykV85p26_0(.dout(w_dff_A_Lm3IZnW65_0),.din(w_dff_A_oykV85p26_0),.clk(gclk));
	jdff dff_A_Lm3IZnW65_0(.dout(w_dff_A_g0i1D3m36_0),.din(w_dff_A_Lm3IZnW65_0),.clk(gclk));
	jdff dff_A_g0i1D3m36_0(.dout(w_dff_A_eUYqKwrW7_0),.din(w_dff_A_g0i1D3m36_0),.clk(gclk));
	jdff dff_A_eUYqKwrW7_0(.dout(w_dff_A_6YL5nnzd4_0),.din(w_dff_A_eUYqKwrW7_0),.clk(gclk));
	jdff dff_A_6YL5nnzd4_0(.dout(w_dff_A_pimnF4Yg8_0),.din(w_dff_A_6YL5nnzd4_0),.clk(gclk));
	jdff dff_A_pimnF4Yg8_0(.dout(w_dff_A_WzTSYKqK5_0),.din(w_dff_A_pimnF4Yg8_0),.clk(gclk));
	jdff dff_A_WzTSYKqK5_0(.dout(G350),.din(w_dff_A_WzTSYKqK5_0),.clk(gclk));
	jdff dff_A_fHXgdtt22_2(.dout(w_dff_A_gTNWBnM93_0),.din(w_dff_A_fHXgdtt22_2),.clk(gclk));
	jdff dff_A_gTNWBnM93_0(.dout(w_dff_A_TdsFmoIP6_0),.din(w_dff_A_gTNWBnM93_0),.clk(gclk));
	jdff dff_A_TdsFmoIP6_0(.dout(w_dff_A_gAUiuOrl9_0),.din(w_dff_A_TdsFmoIP6_0),.clk(gclk));
	jdff dff_A_gAUiuOrl9_0(.dout(w_dff_A_Muibnq176_0),.din(w_dff_A_gAUiuOrl9_0),.clk(gclk));
	jdff dff_A_Muibnq176_0(.dout(w_dff_A_oVp5WkuG8_0),.din(w_dff_A_Muibnq176_0),.clk(gclk));
	jdff dff_A_oVp5WkuG8_0(.dout(w_dff_A_xtkFZcCD1_0),.din(w_dff_A_oVp5WkuG8_0),.clk(gclk));
	jdff dff_A_xtkFZcCD1_0(.dout(w_dff_A_qQDQ2b2E7_0),.din(w_dff_A_xtkFZcCD1_0),.clk(gclk));
	jdff dff_A_qQDQ2b2E7_0(.dout(w_dff_A_qJXakTve7_0),.din(w_dff_A_qQDQ2b2E7_0),.clk(gclk));
	jdff dff_A_qJXakTve7_0(.dout(w_dff_A_WlpHqxfu4_0),.din(w_dff_A_qJXakTve7_0),.clk(gclk));
	jdff dff_A_WlpHqxfu4_0(.dout(w_dff_A_ybmJz2dY0_0),.din(w_dff_A_WlpHqxfu4_0),.clk(gclk));
	jdff dff_A_ybmJz2dY0_0(.dout(w_dff_A_4uaK6ABo8_0),.din(w_dff_A_ybmJz2dY0_0),.clk(gclk));
	jdff dff_A_4uaK6ABo8_0(.dout(w_dff_A_Q2BsnpJv6_0),.din(w_dff_A_4uaK6ABo8_0),.clk(gclk));
	jdff dff_A_Q2BsnpJv6_0(.dout(w_dff_A_YEAUu2gz1_0),.din(w_dff_A_Q2BsnpJv6_0),.clk(gclk));
	jdff dff_A_YEAUu2gz1_0(.dout(w_dff_A_xXTSCJ4S6_0),.din(w_dff_A_YEAUu2gz1_0),.clk(gclk));
	jdff dff_A_xXTSCJ4S6_0(.dout(w_dff_A_VECBTTSw6_0),.din(w_dff_A_xXTSCJ4S6_0),.clk(gclk));
	jdff dff_A_VECBTTSw6_0(.dout(G353),.din(w_dff_A_VECBTTSw6_0),.clk(gclk));
	jdff dff_A_DuDkDjYi5_2(.dout(w_dff_A_dDB7qp5P3_0),.din(w_dff_A_DuDkDjYi5_2),.clk(gclk));
	jdff dff_A_dDB7qp5P3_0(.dout(w_dff_A_ujPwQOr92_0),.din(w_dff_A_dDB7qp5P3_0),.clk(gclk));
	jdff dff_A_ujPwQOr92_0(.dout(w_dff_A_uv51KXtt9_0),.din(w_dff_A_ujPwQOr92_0),.clk(gclk));
	jdff dff_A_uv51KXtt9_0(.dout(w_dff_A_8SNbUtTT7_0),.din(w_dff_A_uv51KXtt9_0),.clk(gclk));
	jdff dff_A_8SNbUtTT7_0(.dout(w_dff_A_VDkiLel90_0),.din(w_dff_A_8SNbUtTT7_0),.clk(gclk));
	jdff dff_A_VDkiLel90_0(.dout(w_dff_A_Xq16iuJx4_0),.din(w_dff_A_VDkiLel90_0),.clk(gclk));
	jdff dff_A_Xq16iuJx4_0(.dout(w_dff_A_EmpRYlBd5_0),.din(w_dff_A_Xq16iuJx4_0),.clk(gclk));
	jdff dff_A_EmpRYlBd5_0(.dout(w_dff_A_zQ4WrqJF6_0),.din(w_dff_A_EmpRYlBd5_0),.clk(gclk));
	jdff dff_A_zQ4WrqJF6_0(.dout(w_dff_A_TaBkhPJf7_0),.din(w_dff_A_zQ4WrqJF6_0),.clk(gclk));
	jdff dff_A_TaBkhPJf7_0(.dout(w_dff_A_Xnsx3GZd2_0),.din(w_dff_A_TaBkhPJf7_0),.clk(gclk));
	jdff dff_A_Xnsx3GZd2_0(.dout(w_dff_A_qPoyoRLT4_0),.din(w_dff_A_Xnsx3GZd2_0),.clk(gclk));
	jdff dff_A_qPoyoRLT4_0(.dout(w_dff_A_7PqEaO3n3_0),.din(w_dff_A_qPoyoRLT4_0),.clk(gclk));
	jdff dff_A_7PqEaO3n3_0(.dout(w_dff_A_WYwLRXyU9_0),.din(w_dff_A_7PqEaO3n3_0),.clk(gclk));
	jdff dff_A_WYwLRXyU9_0(.dout(w_dff_A_LxYwAEA64_0),.din(w_dff_A_WYwLRXyU9_0),.clk(gclk));
	jdff dff_A_LxYwAEA64_0(.dout(w_dff_A_TAKFhnAa9_0),.din(w_dff_A_LxYwAEA64_0),.clk(gclk));
	jdff dff_A_TAKFhnAa9_0(.dout(w_dff_A_NVjqnmDu3_0),.din(w_dff_A_TAKFhnAa9_0),.clk(gclk));
	jdff dff_A_NVjqnmDu3_0(.dout(w_dff_A_xgoaf3wx5_0),.din(w_dff_A_NVjqnmDu3_0),.clk(gclk));
	jdff dff_A_xgoaf3wx5_0(.dout(G356),.din(w_dff_A_xgoaf3wx5_0),.clk(gclk));
	jdff dff_A_jSAFT7W59_2(.dout(w_dff_A_ithHaM9Q9_0),.din(w_dff_A_jSAFT7W59_2),.clk(gclk));
	jdff dff_A_ithHaM9Q9_0(.dout(w_dff_A_v6w6Ftd80_0),.din(w_dff_A_ithHaM9Q9_0),.clk(gclk));
	jdff dff_A_v6w6Ftd80_0(.dout(w_dff_A_Vl2GIAja8_0),.din(w_dff_A_v6w6Ftd80_0),.clk(gclk));
	jdff dff_A_Vl2GIAja8_0(.dout(w_dff_A_Cmblx7ZX3_0),.din(w_dff_A_Vl2GIAja8_0),.clk(gclk));
	jdff dff_A_Cmblx7ZX3_0(.dout(w_dff_A_t9rU1ift3_0),.din(w_dff_A_Cmblx7ZX3_0),.clk(gclk));
	jdff dff_A_t9rU1ift3_0(.dout(G321),.din(w_dff_A_t9rU1ift3_0),.clk(gclk));
	jdff dff_A_ViLkVnO16_2(.dout(G338),.din(w_dff_A_ViLkVnO16_2),.clk(gclk));
	jdff dff_A_zgLAj29Z1_2(.dout(w_dff_A_8Py4PAuS1_0),.din(w_dff_A_zgLAj29Z1_2),.clk(gclk));
	jdff dff_A_8Py4PAuS1_0(.dout(w_dff_A_i0vAyBVg6_0),.din(w_dff_A_8Py4PAuS1_0),.clk(gclk));
	jdff dff_A_i0vAyBVg6_0(.dout(w_dff_A_LbjnRCS27_0),.din(w_dff_A_i0vAyBVg6_0),.clk(gclk));
	jdff dff_A_LbjnRCS27_0(.dout(w_dff_A_n8oqx6re5_0),.din(w_dff_A_LbjnRCS27_0),.clk(gclk));
	jdff dff_A_n8oqx6re5_0(.dout(w_dff_A_00ppykpA8_0),.din(w_dff_A_n8oqx6re5_0),.clk(gclk));
	jdff dff_A_00ppykpA8_0(.dout(w_dff_A_kaB0RiT85_0),.din(w_dff_A_00ppykpA8_0),.clk(gclk));
	jdff dff_A_kaB0RiT85_0(.dout(w_dff_A_rcSvvZI04_0),.din(w_dff_A_kaB0RiT85_0),.clk(gclk));
	jdff dff_A_rcSvvZI04_0(.dout(w_dff_A_GfgDLexN6_0),.din(w_dff_A_rcSvvZI04_0),.clk(gclk));
	jdff dff_A_GfgDLexN6_0(.dout(w_dff_A_OWNeayUu7_0),.din(w_dff_A_GfgDLexN6_0),.clk(gclk));
	jdff dff_A_OWNeayUu7_0(.dout(w_dff_A_bquQDG432_0),.din(w_dff_A_OWNeayUu7_0),.clk(gclk));
	jdff dff_A_bquQDG432_0(.dout(w_dff_A_kOGCfB0W4_0),.din(w_dff_A_bquQDG432_0),.clk(gclk));
	jdff dff_A_kOGCfB0W4_0(.dout(w_dff_A_xkYPtzHz6_0),.din(w_dff_A_kOGCfB0W4_0),.clk(gclk));
	jdff dff_A_xkYPtzHz6_0(.dout(w_dff_A_I849F7qj0_0),.din(w_dff_A_xkYPtzHz6_0),.clk(gclk));
	jdff dff_A_I849F7qj0_0(.dout(w_dff_A_jfGPZSUK9_0),.din(w_dff_A_I849F7qj0_0),.clk(gclk));
	jdff dff_A_jfGPZSUK9_0(.dout(w_dff_A_EJgYPLe23_0),.din(w_dff_A_jfGPZSUK9_0),.clk(gclk));
	jdff dff_A_EJgYPLe23_0(.dout(w_dff_A_tx596gK83_0),.din(w_dff_A_EJgYPLe23_0),.clk(gclk));
	jdff dff_A_tx596gK83_0(.dout(G370),.din(w_dff_A_tx596gK83_0),.clk(gclk));
	jdff dff_A_h2dOt8HR5_2(.dout(w_dff_A_hqGjitwK4_0),.din(w_dff_A_h2dOt8HR5_2),.clk(gclk));
	jdff dff_A_hqGjitwK4_0(.dout(w_dff_A_jjcjwSm05_0),.din(w_dff_A_hqGjitwK4_0),.clk(gclk));
	jdff dff_A_jjcjwSm05_0(.dout(w_dff_A_F75Ogi0B6_0),.din(w_dff_A_jjcjwSm05_0),.clk(gclk));
	jdff dff_A_F75Ogi0B6_0(.dout(w_dff_A_FU5Di0Jo4_0),.din(w_dff_A_F75Ogi0B6_0),.clk(gclk));
	jdff dff_A_FU5Di0Jo4_0(.dout(w_dff_A_sOfyeLFc0_0),.din(w_dff_A_FU5Di0Jo4_0),.clk(gclk));
	jdff dff_A_sOfyeLFc0_0(.dout(w_dff_A_4JhhMymf1_0),.din(w_dff_A_sOfyeLFc0_0),.clk(gclk));
	jdff dff_A_4JhhMymf1_0(.dout(w_dff_A_Y3P78nY31_0),.din(w_dff_A_4JhhMymf1_0),.clk(gclk));
	jdff dff_A_Y3P78nY31_0(.dout(w_dff_A_aNI955nh5_0),.din(w_dff_A_Y3P78nY31_0),.clk(gclk));
	jdff dff_A_aNI955nh5_0(.dout(w_dff_A_aU3f0mlL2_0),.din(w_dff_A_aNI955nh5_0),.clk(gclk));
	jdff dff_A_aU3f0mlL2_0(.dout(w_dff_A_n6MTmMDB2_0),.din(w_dff_A_aU3f0mlL2_0),.clk(gclk));
	jdff dff_A_n6MTmMDB2_0(.dout(w_dff_A_YGVnJeVP7_0),.din(w_dff_A_n6MTmMDB2_0),.clk(gclk));
	jdff dff_A_YGVnJeVP7_0(.dout(w_dff_A_MYi7ROnW9_0),.din(w_dff_A_YGVnJeVP7_0),.clk(gclk));
	jdff dff_A_MYi7ROnW9_0(.dout(w_dff_A_EIJTCDdr0_0),.din(w_dff_A_MYi7ROnW9_0),.clk(gclk));
	jdff dff_A_EIJTCDdr0_0(.dout(w_dff_A_n1wO9CLk5_0),.din(w_dff_A_EIJTCDdr0_0),.clk(gclk));
	jdff dff_A_n1wO9CLk5_0(.dout(w_dff_A_hRfp8CU42_0),.din(w_dff_A_n1wO9CLk5_0),.clk(gclk));
	jdff dff_A_hRfp8CU42_0(.dout(w_dff_A_YlkdBaCC6_0),.din(w_dff_A_hRfp8CU42_0),.clk(gclk));
	jdff dff_A_YlkdBaCC6_0(.dout(w_dff_A_uxLl9poC2_0),.din(w_dff_A_YlkdBaCC6_0),.clk(gclk));
	jdff dff_A_uxLl9poC2_0(.dout(w_dff_A_MmJRikpF7_0),.din(w_dff_A_uxLl9poC2_0),.clk(gclk));
	jdff dff_A_MmJRikpF7_0(.dout(w_dff_A_X5aQ5GJ57_0),.din(w_dff_A_MmJRikpF7_0),.clk(gclk));
	jdff dff_A_X5aQ5GJ57_0(.dout(w_dff_A_vRhT0YsU5_0),.din(w_dff_A_X5aQ5GJ57_0),.clk(gclk));
	jdff dff_A_vRhT0YsU5_0(.dout(G399),.din(w_dff_A_vRhT0YsU5_0),.clk(gclk));
endmodule

