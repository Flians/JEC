/*
gf_c499:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jdff: 477
	jand: 69
	jor: 2

Summary:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jdff: 477
	jand: 69
	jor: 2

The maximum logic level gap of any gate:
	gf_c499: 11
*/

module gf_c499(gclk, Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr, God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10, God11, God12, God13, God14, God15, God16, God17, God18, God19, God20, God21, God22, God23, God24, God25, God26, God27, God28, God29, God30, God31);
	input gclk;
	input Gid0;
	input Gid1;
	input Gid2;
	input Gid3;
	input Gid4;
	input Gid5;
	input Gid6;
	input Gid7;
	input Gid8;
	input Gid9;
	input Gid10;
	input Gid11;
	input Gid12;
	input Gid13;
	input Gid14;
	input Gid15;
	input Gid16;
	input Gid17;
	input Gid18;
	input Gid19;
	input Gid20;
	input Gid21;
	input Gid22;
	input Gid23;
	input Gid24;
	input Gid25;
	input Gid26;
	input Gid27;
	input Gid28;
	input Gid29;
	input Gid30;
	input Gid31;
	input Gic0;
	input Gic1;
	input Gic2;
	input Gic3;
	input Gic4;
	input Gic5;
	input Gic6;
	input Gic7;
	input Gr;
	output God0;
	output God1;
	output God2;
	output God3;
	output God4;
	output God5;
	output God6;
	output God7;
	output God8;
	output God9;
	output God10;
	output God11;
	output God12;
	output God13;
	output God14;
	output God15;
	output God16;
	output God17;
	output God18;
	output God19;
	output God20;
	output God21;
	output God22;
	output God23;
	output God24;
	output God25;
	output God26;
	output God27;
	output God28;
	output God29;
	output God30;
	output God31;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n180;
	wire n182;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n208;
	wire n210;
	wire n212;
	wire n214;
	wire n215;
	wire n217;
	wire n219;
	wire n221;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n236;
	wire n238;
	wire n240;
	wire n242;
	wire n243;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n257;
	wire n259;
	wire n261;
	wire n263;
	wire n264;
	wire n266;
	wire n268;
	wire n270;
	wire [2:0] w_Gid0_0;
	wire [2:0] w_Gid1_0;
	wire [2:0] w_Gid2_0;
	wire [2:0] w_Gid3_0;
	wire [2:0] w_Gid4_0;
	wire [2:0] w_Gid5_0;
	wire [2:0] w_Gid6_0;
	wire [2:0] w_Gid7_0;
	wire [2:0] w_Gid8_0;
	wire [2:0] w_Gid9_0;
	wire [2:0] w_Gid10_0;
	wire [2:0] w_Gid11_0;
	wire [2:0] w_Gid12_0;
	wire [2:0] w_Gid13_0;
	wire [2:0] w_Gid14_0;
	wire [2:0] w_Gid15_0;
	wire [2:0] w_Gid16_0;
	wire [2:0] w_Gid17_0;
	wire [2:0] w_Gid18_0;
	wire [2:0] w_Gid19_0;
	wire [2:0] w_Gid20_0;
	wire [2:0] w_Gid21_0;
	wire [2:0] w_Gid22_0;
	wire [2:0] w_Gid23_0;
	wire [2:0] w_Gid24_0;
	wire [2:0] w_Gid25_0;
	wire [2:0] w_Gid26_0;
	wire [2:0] w_Gid27_0;
	wire [2:0] w_Gid28_0;
	wire [2:0] w_Gid29_0;
	wire [2:0] w_Gid30_0;
	wire [2:0] w_Gid31_0;
	wire [2:0] w_Gr_0;
	wire [2:0] w_Gr_1;
	wire [2:0] w_Gr_2;
	wire [1:0] w_Gr_3;
	wire [1:0] w_n75_0;
	wire [1:0] w_n76_0;
	wire [1:0] w_n80_0;
	wire [1:0] w_n83_0;
	wire [1:0] w_n84_0;
	wire [2:0] w_n85_0;
	wire [2:0] w_n85_1;
	wire [1:0] w_n85_2;
	wire [1:0] w_n88_0;
	wire [1:0] w_n89_0;
	wire [1:0] w_n94_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n110_0;
	wire [2:0] w_n112_0;
	wire [2:0] w_n112_1;
	wire [2:0] w_n112_2;
	wire [1:0] w_n113_0;
	wire [1:0] w_n116_0;
	wire [1:0] w_n117_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n124_0;
	wire [1:0] w_n125_0;
	wire [2:0] w_n126_0;
	wire [2:0] w_n126_1;
	wire [1:0] w_n126_2;
	wire [1:0] w_n128_0;
	wire [1:0] w_n134_0;
	wire [1:0] w_n135_0;
	wire [1:0] w_n136_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n143_0;
	wire [2:0] w_n147_0;
	wire [2:0] w_n147_1;
	wire [1:0] w_n147_2;
	wire [2:0] w_n149_0;
	wire [2:0] w_n149_1;
	wire [1:0] w_n149_2;
	wire [1:0] w_n153_0;
	wire [1:0] w_n156_0;
	wire [2:0] w_n159_0;
	wire [2:0] w_n166_0;
	wire [2:0] w_n166_1;
	wire [2:0] w_n166_2;
	wire [1:0] w_n169_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n173_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n175_0;
	wire [2:0] w_n177_0;
	wire [1:0] w_n177_1;
	wire [2:0] w_n187_0;
	wire [2:0] w_n187_1;
	wire [1:0] w_n187_2;
	wire [1:0] w_n188_0;
	wire [1:0] w_n190_0;
	wire [2:0] w_n191_0;
	wire [1:0] w_n191_1;
	wire [1:0] w_n200_0;
	wire [2:0] w_n202_0;
	wire [2:0] w_n202_1;
	wire [1:0] w_n202_2;
	wire [1:0] w_n203_0;
	wire [2:0] w_n205_0;
	wire [1:0] w_n205_1;
	wire [2:0] w_n214_0;
	wire [1:0] w_n214_1;
	wire [1:0] w_n223_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n233_0;
	wire [1:0] w_n233_1;
	wire [1:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [1:0] w_n243_1;
	wire [1:0] w_n253_0;
	wire [2:0] w_n254_0;
	wire [1:0] w_n254_1;
	wire [2:0] w_n263_0;
	wire [1:0] w_n263_1;
	wire w_dff_A_aDdyPWb38_0;
	wire w_dff_B_rcJR4sP54_2;
	wire w_dff_B_QzVgACRg1_2;
	wire w_dff_A_6GE9eT2e6_1;
	wire w_dff_B_Bv2Pjeql0_2;
	wire w_dff_B_PvPK2uh24_2;
	wire w_dff_B_U6YQwxGQ5_2;
	wire w_dff_B_u6YsHwn04_2;
	wire w_dff_B_K1qUrywU9_0;
	wire w_dff_A_vYm9ffK76_0;
	wire w_dff_A_8m7vKhDh8_0;
	wire w_dff_A_jTKP7wBN4_0;
	wire w_dff_A_rdAhtn6n6_0;
	wire w_dff_A_BpR7RP2O6_0;
	wire w_dff_A_IaMk4a494_0;
	wire w_dff_A_tz9wkayk6_0;
	wire w_dff_A_8CAR0Ip75_0;
	wire w_dff_A_nA7QdfNz7_0;
	wire w_dff_A_zKRcJdAD1_0;
	wire w_dff_A_0QEC5RPS1_0;
	wire w_dff_A_rNaUt7z90_0;
	wire w_dff_A_oWVKbCJm2_0;
	wire w_dff_A_njpK3b4y3_0;
	wire w_dff_A_Yz4tRNK61_0;
	wire w_dff_A_MXWJnoX17_0;
	wire w_dff_A_4XJDLIu03_0;
	wire w_dff_A_gz9d8heg8_0;
	wire w_dff_A_xlqmfJVf2_0;
	wire w_dff_A_AcoMs2LU8_0;
	wire w_dff_B_aFKaFGhu2_1;
	wire w_dff_B_eq9fE1rP2_1;
	wire w_dff_B_ZnGIKCip6_1;
	wire w_dff_A_Lcf74BXH1_0;
	wire w_dff_A_yQRXNvKO5_0;
	wire w_dff_A_GNcnHxCq3_0;
	wire w_dff_A_kTdAH3H60_0;
	wire w_dff_A_ItvWWmwT7_0;
	wire w_dff_B_Ae8t9VTK3_2;
	wire w_dff_B_dfkZpVnf5_2;
	wire w_dff_B_HHc0DKmb7_2;
	wire w_dff_B_1bGkhgnf2_2;
	wire w_dff_A_y8WsmTur5_0;
	wire w_dff_A_B6YCX7mG2_0;
	wire w_dff_A_2feKF3Zk2_0;
	wire w_dff_A_FK9RJOmj1_0;
	wire w_dff_A_Pwr49xPF5_0;
	wire w_dff_B_hESeV1NC0_1;
	wire w_dff_B_LSyfilou3_1;
	wire w_dff_B_rl6k19680_1;
	wire w_dff_A_dRHQyIA50_1;
	wire w_dff_A_66PxB4UL7_0;
	wire w_dff_A_fBWtJRhz3_0;
	wire w_dff_A_zuwmcgl61_0;
	wire w_dff_A_ZCoSJqDL0_0;
	wire w_dff_A_HPvauYvh8_0;
	wire w_dff_A_cxvYa9bb2_0;
	wire w_dff_A_NDutoFw33_2;
	wire w_dff_A_e1EDB06P4_2;
	wire w_dff_A_4IkPgO2g2_2;
	wire w_dff_A_ZzQbgp3B2_2;
	wire w_dff_A_ksU8C2KW5_2;
	wire w_dff_A_gCAR8UGY4_2;
	wire w_dff_A_ykLkWruT0_0;
	wire w_dff_A_QOKelfPT2_0;
	wire w_dff_A_JyJpomq77_0;
	wire w_dff_A_2i641phh3_0;
	wire w_dff_A_YPAYDX9B4_0;
	wire w_dff_A_jiBeYxFr6_0;
	wire w_dff_A_wddZOLmr2_0;
	wire w_dff_A_vQpDA4Vz2_0;
	wire w_dff_A_7REOox3M7_2;
	wire w_dff_A_EJ3WYniq1_2;
	wire w_dff_A_qqG1XOGj3_2;
	wire w_dff_A_Mwo6TomW6_2;
	wire w_dff_A_yYXSBgGe6_2;
	wire w_dff_A_ohv5oZ1X2_2;
	wire w_dff_B_Wmn3ofzU8_0;
	wire w_dff_A_BlxLJbn71_1;
	wire w_dff_A_DI3JYTHQ3_0;
	wire w_dff_A_Hm5n4ftz9_0;
	wire w_dff_A_ipGqDGh94_0;
	wire w_dff_A_8HehDjDy2_0;
	wire w_dff_A_O9Bze4Dq9_0;
	wire w_dff_A_HCBrWaSp5_0;
	wire w_dff_A_x0x1Am6P9_2;
	wire w_dff_A_cSpIwoL75_2;
	wire w_dff_A_j6NDuhV37_2;
	wire w_dff_A_nhBJw5ZR7_2;
	wire w_dff_A_uGMXUnrz9_2;
	wire w_dff_A_XhUlaSPc8_2;
	wire w_dff_A_QKvtC1f67_0;
	wire w_dff_A_mneKHFDU5_0;
	wire w_dff_A_4kVdwhdl2_0;
	wire w_dff_A_sDuJvpTu9_0;
	wire w_dff_A_e4GOGSkB8_0;
	wire w_dff_A_HFfemwmf6_0;
	wire w_dff_A_KBcOM4Jl7_0;
	wire w_dff_A_shjmP9hR0_0;
	wire w_dff_A_ZBVWvipt1_0;
	wire w_dff_A_FFGOan2N3_0;
	wire w_dff_A_PrYQ8vk06_2;
	wire w_dff_A_HspB0UhW9_2;
	wire w_dff_A_Y6koNCAW7_2;
	wire w_dff_A_5bUNF2l39_2;
	wire w_dff_A_MRD4AoNy9_2;
	wire w_dff_A_uzwkQZ2I5_2;
	wire w_dff_B_u4RzZMEj3_0;
	wire w_dff_A_JE9A9tqp1_0;
	wire w_dff_A_v3ut1IpA9_0;
	wire w_dff_A_CwaotxFj9_0;
	wire w_dff_A_JATZXH7W9_0;
	wire w_dff_A_KkUIyz2i2_0;
	wire w_dff_A_QSOiowHf1_1;
	wire w_dff_A_BFwUrL8z7_0;
	wire w_dff_A_zXBYBGc16_0;
	wire w_dff_A_iFM7iU6v1_0;
	wire w_dff_A_Hxu5YBEq6_0;
	wire w_dff_A_kx1wugWw2_0;
	wire w_dff_A_VvM6vgff7_0;
	wire w_dff_A_r58lH3V02_0;
	wire w_dff_A_wCD0Yq4R2_0;
	wire w_dff_A_UDu7eOFq7_0;
	wire w_dff_A_z1gSDu4R5_0;
	wire w_dff_A_TPnZuobl3_0;
	wire w_dff_A_GQByEKuD8_0;
	wire w_dff_A_jbxrsE4h6_0;
	wire w_dff_A_xMBmPMU74_0;
	wire w_dff_A_4xZOwaeg3_0;
	wire w_dff_A_lJ1zL3Ms5_0;
	wire w_dff_A_9CVvwYn06_0;
	wire w_dff_A_KRopvc4R2_0;
	wire w_dff_A_M4plUTxg3_0;
	wire w_dff_A_P5oWNlu53_0;
	wire w_dff_A_i01bXCXd8_0;
	wire w_dff_A_P9mIro7b7_0;
	wire w_dff_A_Bz7PX8Da4_0;
	wire w_dff_A_AqmayLVM3_0;
	wire w_dff_A_FCqsPleW6_0;
	wire w_dff_A_HoLhvVbY8_0;
	wire w_dff_A_sM694yDn0_0;
	wire w_dff_A_oAfJG4058_0;
	wire w_dff_A_vPyibuVt2_0;
	wire w_dff_A_4gDemzTZ7_0;
	wire w_dff_A_wAzpbYQS3_0;
	wire w_dff_A_bFF7kmy35_0;
	wire w_dff_A_8NOL1TLa2_0;
	wire w_dff_A_NPj9osNJ3_0;
	wire w_dff_A_XzXrlRO07_0;
	wire w_dff_A_yzRbYqvA2_0;
	wire w_dff_A_YnV5BC8T0_0;
	wire w_dff_A_Wln0iari3_0;
	wire w_dff_A_iQnEU6171_0;
	wire w_dff_A_Klm57AT37_0;
	wire w_dff_A_nRbvuv8M9_1;
	wire w_dff_A_hAVEAOku5_0;
	wire w_dff_A_GvIgEcnP9_0;
	wire w_dff_A_Te3X00v68_0;
	wire w_dff_A_q5Yf0Vyz3_0;
	wire w_dff_A_8DPc9Uzb7_0;
	wire w_dff_A_wUv7iXPn9_0;
	wire w_dff_A_9ubRGCaK3_0;
	wire w_dff_A_HABd7t814_0;
	wire w_dff_A_x9baV45f4_0;
	wire w_dff_A_1r2cNNVA0_0;
	wire w_dff_A_vb3rHJys2_0;
	wire w_dff_A_pOuc5m0H8_0;
	wire w_dff_A_CtZl4NmD8_0;
	wire w_dff_A_D6MRQnTe2_0;
	wire w_dff_A_6Tt91TuU1_0;
	wire w_dff_A_xqW3bDJy5_0;
	wire w_dff_A_KtOsEIdM1_0;
	wire w_dff_A_FcfR02qE9_0;
	wire w_dff_A_uam4Mvpt2_0;
	wire w_dff_A_SMk4Rzs98_0;
	wire w_dff_A_6p8rAL8X3_0;
	wire w_dff_A_qBIYq7za9_0;
	wire w_dff_A_8LMXLivq2_0;
	wire w_dff_A_BFZ4Gl6V7_0;
	wire w_dff_A_RYeFefF50_0;
	wire w_dff_A_wtKv9GSC0_0;
	wire w_dff_A_XoTgZfTW8_0;
	wire w_dff_A_N1Saaqg35_0;
	wire w_dff_A_gu1ax10V9_0;
	wire w_dff_A_9wkS9wKr2_0;
	wire w_dff_A_ducNOe8L5_0;
	wire w_dff_A_7D9VR66J9_0;
	wire w_dff_A_8WQZR0Lo2_0;
	wire w_dff_A_hzTifEEj1_0;
	wire w_dff_A_kk0O9RQQ1_0;
	wire w_dff_A_IiNwgC7z6_0;
	wire w_dff_A_ayfZBSiF5_0;
	wire w_dff_A_zCH76v066_0;
	wire w_dff_A_skjfGmJy5_0;
	wire w_dff_A_lLJru4AI4_0;
	wire w_dff_B_i2QgCSY68_2;
	wire w_dff_B_nLoB99Yf0_2;
	wire w_dff_B_5jl0f5es0_2;
	wire w_dff_B_d6TFRYE03_2;
	wire w_dff_A_UgUr8UBQ2_0;
	wire w_dff_A_9vHPGOCY0_0;
	wire w_dff_A_TVdCrnvH6_0;
	wire w_dff_A_mLuBbqSX2_0;
	wire w_dff_A_6RpvnYwd5_0;
	wire w_dff_A_8GFgmSi75_0;
	wire w_dff_A_uAOKY6xX6_0;
	wire w_dff_A_tVccIOZq0_0;
	wire w_dff_A_i68Mpp0q3_0;
	wire w_dff_A_5pI5wIum6_0;
	wire w_dff_A_fhfL7ZNh2_0;
	wire w_dff_A_QtYcn6H17_0;
	wire w_dff_A_N5MTlNjS2_0;
	wire w_dff_A_j8fZ2d6n1_0;
	wire w_dff_A_8RceGFPk9_0;
	wire w_dff_A_Azv9j80w7_0;
	wire w_dff_A_ws4PACSk6_0;
	wire w_dff_A_5PSOEEr27_0;
	wire w_dff_A_g93EImtD5_0;
	wire w_dff_A_0SJj0lBu8_0;
	wire w_dff_A_HNuj0yP36_0;
	wire w_dff_A_zJqql4ae2_0;
	wire w_dff_A_oon9BExA8_0;
	wire w_dff_A_kABiU4ks4_0;
	wire w_dff_A_qzAnkGuX6_0;
	wire w_dff_A_t9UoYn2L6_0;
	wire w_dff_A_yLqZb8ab4_0;
	wire w_dff_A_f1RmbKaB7_0;
	wire w_dff_A_fJL16Qb31_0;
	wire w_dff_A_LyMrNUTW1_0;
	wire w_dff_A_Rn5TqlOD3_0;
	wire w_dff_A_UWXZGQUD1_0;
	wire w_dff_A_KtrV4DP85_0;
	wire w_dff_A_tRHN7J6B8_0;
	wire w_dff_A_EiyU3HGR1_0;
	wire w_dff_A_EWmpaWPZ1_0;
	wire w_dff_A_CNgnRqxO1_0;
	wire w_dff_A_UOdM8lSR2_0;
	wire w_dff_A_rOeqALvP1_0;
	wire w_dff_A_wYS3BdfW6_0;
	wire w_dff_A_qFWcYLoC7_0;
	wire w_dff_A_JmEtiWwd6_0;
	wire w_dff_A_GmVmhRdX0_0;
	wire w_dff_A_WJUEV0YA2_0;
	wire w_dff_A_maGIHF550_0;
	wire w_dff_A_rBrydVzj8_0;
	wire w_dff_A_Yi4eIttP4_0;
	wire w_dff_A_Ab6nBgXj9_0;
	wire w_dff_A_Z9o0sFDI8_0;
	wire w_dff_A_GZgjHeOx8_0;
	wire w_dff_A_kZnL2V1h6_0;
	wire w_dff_A_lGMmi9g90_0;
	wire w_dff_A_BAqnZPKJ8_0;
	wire w_dff_A_vJQWoq4r7_0;
	wire w_dff_A_hQvNw3Qa3_0;
	wire w_dff_A_fsyqxTHM3_0;
	wire w_dff_A_PH0OJDwd1_0;
	wire w_dff_A_k7y2Wtrb7_0;
	wire w_dff_A_nnFGBZ531_0;
	wire w_dff_A_R9sJ7BM73_0;
	wire w_dff_A_nqcVuyQD6_0;
	wire w_dff_A_DJEzk7og9_0;
	wire w_dff_A_F8Vfn9dx4_0;
	wire w_dff_A_WKlTuUQc7_0;
	wire w_dff_A_QMdbRlZh5_0;
	wire w_dff_A_drsbM2rL6_0;
	wire w_dff_A_APMNqhGG7_0;
	wire w_dff_A_UJlRumnJ0_0;
	wire w_dff_A_X69MC0nZ4_0;
	wire w_dff_A_Zu7sxXR45_0;
	wire w_dff_A_7xihvIPF0_0;
	wire w_dff_A_ALfTx6m19_0;
	wire w_dff_A_culgjWxi5_0;
	wire w_dff_A_Pr0Wo26f8_0;
	wire w_dff_A_BCldgjlb5_0;
	wire w_dff_A_zFSxSAr91_0;
	wire w_dff_A_qOe9KJQn9_0;
	wire w_dff_A_mlIfPHH50_0;
	wire w_dff_A_gEQ2B0xt9_0;
	wire w_dff_A_vWwtNhQM4_0;
	wire w_dff_A_qWKTROdI5_0;
	wire w_dff_A_eu05rmxx8_0;
	wire w_dff_A_T2YkXJPR8_0;
	wire w_dff_A_VQhWYieE2_0;
	wire w_dff_A_9ma5OEpZ6_0;
	wire w_dff_A_8BagOsUg4_0;
	wire w_dff_A_HMtBuOwS0_0;
	wire w_dff_A_3k77Rm1d7_0;
	wire w_dff_A_Rt1Zs4yD5_0;
	wire w_dff_A_R6hLT1gF6_0;
	wire w_dff_A_Ee2OX39E3_0;
	wire w_dff_A_pMjxcQUz9_0;
	wire w_dff_A_JH6rEZM93_0;
	wire w_dff_A_Ccze5qj86_0;
	wire w_dff_A_LX3bRr914_0;
	wire w_dff_A_I8rUbnB55_0;
	wire w_dff_A_hJqy3NvD0_0;
	wire w_dff_A_LmhYSz0f9_0;
	wire w_dff_A_8M1roRHN0_0;
	wire w_dff_A_ER1JIcbh4_0;
	wire w_dff_A_zEsPKpjQ5_0;
	wire w_dff_A_XhjLBntL7_0;
	wire w_dff_A_mL1eZsne1_0;
	wire w_dff_A_vA3dOAXc9_0;
	wire w_dff_A_kbDH5LK66_0;
	wire w_dff_A_1uTknrlB2_0;
	wire w_dff_A_JDtv5Dbc7_0;
	wire w_dff_A_hAJX8MYo6_0;
	wire w_dff_A_SkR9i0C66_0;
	wire w_dff_A_nLTRSfP39_0;
	wire w_dff_A_IZAKN65i9_0;
	wire w_dff_A_fU09Vo9m5_0;
	wire w_dff_A_IKH5coRy4_0;
	wire w_dff_A_mNK3ulU47_0;
	wire w_dff_A_c2ZlCHke9_0;
	wire w_dff_A_AXj4PQA77_0;
	wire w_dff_A_bDJzTEBM7_0;
	wire w_dff_A_VCEw40Ni6_0;
	wire w_dff_A_4XYts8Ih4_0;
	wire w_dff_A_OiQ4UZXn2_0;
	wire w_dff_A_GEQXTNG92_0;
	wire w_dff_A_TrJ5Ua3e6_0;
	wire w_dff_A_gi3HS6BD6_0;
	wire w_dff_A_i8cqEZ3d1_0;
	wire w_dff_A_y7p6YtTU9_0;
	wire w_dff_A_Gbttuphg8_0;
	wire w_dff_A_Da0CxEfd3_0;
	wire w_dff_A_KCBCdx4k0_0;
	wire w_dff_A_TQHmocMZ4_0;
	wire w_dff_A_BNTmMqoF1_0;
	wire w_dff_A_54N0ugNR8_0;
	wire w_dff_A_YiYD7WbE9_0;
	wire w_dff_A_NkiZxHnA9_0;
	wire w_dff_A_UsLC33ks8_0;
	wire w_dff_A_XXhkhR7c0_0;
	wire w_dff_A_7qIiETBN5_0;
	wire w_dff_A_yCSWFzxC4_0;
	wire w_dff_A_z0xVy3rQ8_0;
	wire w_dff_A_Fl31Y6cF4_0;
	wire w_dff_A_XBN8ZKPt8_0;
	wire w_dff_A_hZtC0qdE5_0;
	wire w_dff_A_qTZFW09T6_0;
	wire w_dff_A_WYgKLuSK9_0;
	wire w_dff_A_ipJAZuyO5_0;
	wire w_dff_A_Shhlcgov3_0;
	wire w_dff_A_8BknCDYj9_0;
	wire w_dff_A_bfr27rka7_0;
	wire w_dff_A_t2CEq2bh9_0;
	wire w_dff_A_xqUB5j9J1_0;
	wire w_dff_A_60zMKwgT3_0;
	wire w_dff_A_FYOqB6Jq1_0;
	wire w_dff_A_PuMsEJvb8_0;
	wire w_dff_A_vupwB64w1_0;
	wire w_dff_A_vn5rWJvX4_0;
	wire w_dff_A_L7uZj2Jn7_0;
	wire w_dff_A_lG6GjrXS9_0;
	wire w_dff_A_7gIX5W2F1_0;
	wire w_dff_A_40U1t4ak5_0;
	wire w_dff_A_yaObO7Ng2_0;
	wire w_dff_A_D0kKTEau4_0;
	wire w_dff_A_gQzXy2BT0_0;
	wire w_dff_A_JuY88UlQ3_0;
	wire w_dff_A_e7s5LfX73_0;
	wire w_dff_A_9kS1c7it8_0;
	wire w_dff_A_E4hNQIqu8_0;
	wire w_dff_A_QPhhcsxM2_0;
	wire w_dff_A_CBl3IIGX8_0;
	wire w_dff_A_pBg22DGl9_0;
	wire w_dff_A_xmyBsTe45_0;
	wire w_dff_A_T4A39mOC7_0;
	wire w_dff_A_ySQpeBkw8_0;
	wire w_dff_A_xEK5MWRf0_0;
	wire w_dff_A_xbrBFJZR3_0;
	wire w_dff_A_DnccThX34_0;
	wire w_dff_A_Rp9G3c4u3_0;
	wire w_dff_A_EBBf7ufV7_0;
	wire w_dff_A_mTG1dvKJ5_0;
	wire w_dff_A_wVx6AIv85_0;
	wire w_dff_A_FK2uUZDw2_0;
	wire w_dff_A_X95GqGPh5_0;
	wire w_dff_A_iNpbyG9T4_0;
	wire w_dff_A_d1OKbcRq4_0;
	wire w_dff_A_E28qXkd37_0;
	wire w_dff_A_Ubj9B6lp2_0;
	wire w_dff_A_OWywckru0_0;
	wire w_dff_A_X5Pwss0z4_0;
	wire w_dff_A_lCN1uvi33_0;
	wire w_dff_A_V5zIibt05_0;
	wire w_dff_A_QhE8VnNu5_0;
	wire w_dff_A_QVH7nSfG6_0;
	wire w_dff_A_WGwoBsqf6_0;
	wire w_dff_A_m0p89FOw6_0;
	wire w_dff_A_uUIN0ozZ2_0;
	wire w_dff_A_SdPtLtkQ1_0;
	wire w_dff_A_XW0H1AoH0_0;
	wire w_dff_A_QMFA5xbD2_0;
	wire w_dff_A_ZZGI2iuE9_0;
	wire w_dff_A_xZ34f1IN0_0;
	wire w_dff_A_WvYyWxzg7_0;
	wire w_dff_A_m0X0DNV68_0;
	wire w_dff_A_BJiU8Dli1_0;
	wire w_dff_A_HgPP4Jc56_0;
	wire w_dff_A_NxDc3Nsk1_0;
	wire w_dff_A_oIdN7jbs0_0;
	wire w_dff_A_kXAsLSNA0_0;
	wire w_dff_A_44Qqi6fu9_0;
	wire w_dff_A_MdgH81Vo4_0;
	wire w_dff_A_TUXxjpHt8_0;
	wire w_dff_A_T3JgPuRN1_0;
	wire w_dff_A_6Ut0vQrG8_0;
	wire w_dff_A_kpB5NQOi3_0;
	wire w_dff_A_KB8rMTdo9_0;
	wire w_dff_A_npAutbBS9_0;
	wire w_dff_A_TA17G0Iy6_0;
	wire w_dff_A_1NjX9CGf4_0;
	wire w_dff_A_rEfNOk1Z8_0;
	wire w_dff_A_Wfivb2Fg1_0;
	wire w_dff_A_dDbXMIj37_0;
	wire w_dff_A_ieHKHVNB2_0;
	wire w_dff_A_I3AI6Ynl2_0;
	wire w_dff_A_1NfHusSD0_0;
	wire w_dff_A_GXEKt2T89_0;
	wire w_dff_A_bLcg0G0I9_0;
	wire w_dff_A_jXpx4bnO2_0;
	wire w_dff_A_1nL2d3l84_0;
	wire w_dff_A_DXADtZmy9_0;
	wire w_dff_A_IUELqlgn3_0;
	wire w_dff_A_78fXIHfE7_0;
	wire w_dff_A_WBG4S1Ro9_0;
	wire w_dff_A_azHUBSfr1_0;
	wire w_dff_A_OvFkGplN9_0;
	wire w_dff_A_pjxyb87j2_0;
	wire w_dff_A_9dhgkiV36_0;
	wire w_dff_A_uSrkTRLw1_0;
	wire w_dff_A_KTtfpoyp0_0;
	wire w_dff_A_6uFoeYcl2_0;
	wire w_dff_A_Mad77qnx2_0;
	wire w_dff_A_fu0y72oP4_0;
	wire w_dff_A_WrbW5WG71_0;
	wire w_dff_A_zYdL2D6e2_0;
	wire w_dff_A_C0FtiK1q2_0;
	wire w_dff_A_xZbhjjVs0_0;
	wire w_dff_A_xEvsVRYM8_0;
	wire w_dff_A_6cnefFmO1_0;
	wire w_dff_A_dqvs45f62_0;
	wire w_dff_A_tSlxDHv67_0;
	wire w_dff_A_4hMMClrs5_0;
	wire w_dff_A_BC7Rpd9W8_0;
	wire w_dff_A_y0DY56H69_0;
	wire w_dff_A_Osg1ps4M8_0;
	wire w_dff_A_su0c3OnU2_0;
	wire w_dff_A_ErCKavnX3_0;
	wire w_dff_A_R0VntRor0_0;
	wire w_dff_A_5kiC1pva1_0;
	wire w_dff_A_fYFzoGo40_0;
	wire w_dff_A_krNofpEG7_0;
	wire w_dff_A_AjSCsUfW6_0;
	wire w_dff_A_6HlXHswn6_0;
	wire w_dff_A_vpL9BUYb6_0;
	wire w_dff_A_yZj45uEo2_0;
	wire w_dff_A_pDS8zIsB7_0;
	wire w_dff_A_aBvtiYMn9_0;
	wire w_dff_A_iJKwPfTv6_0;
	wire w_dff_A_PMYQK5Tj0_2;
	wire w_dff_A_5M6o6Ub95_2;
	wire w_dff_A_34PC55qj0_2;
	wire w_dff_A_VTAVybd45_2;
	wire w_dff_A_Fwn0Ij8d6_2;
	wire w_dff_A_n7m9VX7F7_2;
	wire w_dff_A_PYCXl0ap5_2;
	wire w_dff_A_XgvbmHBM3_2;
	wire w_dff_A_SsQEgfrU1_2;
	wire w_dff_A_P1nnemrt1_2;
	wire w_dff_A_YC1eikXb3_2;
	wire w_dff_A_gri3Jqev7_2;
	wire w_dff_A_wRRP0kLL9_2;
	wire w_dff_A_4nkykmME2_2;
	wire w_dff_A_UxhabKGn3_2;
	wire w_dff_A_7GIr0kJS3_2;
	jxor g000(.dina(w_Gid12_0[2]),.dinb(w_Gid8_0[2]),.dout(n73),.clk(gclk));
	jxor g001(.dina(w_Gid4_0[2]),.dinb(w_Gid0_0[2]),.dout(n74),.clk(gclk));
	jxor g002(.dina(n74),.dinb(n73),.dout(n75),.clk(gclk));
	jand g003(.dina(w_Gr_3[1]),.dinb(Gic0),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_n76_0[1]),.dinb(w_n75_0[1]),.dout(n77),.clk(gclk));
	jxor g005(.dina(w_Gid19_0[2]),.dinb(w_Gid18_0[2]),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_Gid17_0[2]),.dinb(w_Gid16_0[2]),.dout(n79),.clk(gclk));
	jxor g007(.dina(n79),.dinb(n78),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_Gid23_0[2]),.dinb(w_Gid22_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(w_Gid21_0[2]),.dinb(w_Gid20_0[2]),.dout(n82),.clk(gclk));
	jxor g010(.dina(n82),.dinb(n81),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_n83_0[1]),.dinb(w_n80_0[1]),.dout(n84),.clk(gclk));
	jxor g012(.dina(w_n84_0[1]),.dinb(n77),.dout(n85),.clk(gclk));
	jxor g013(.dina(w_Gid31_0[2]),.dinb(w_Gid27_0[2]),.dout(n86),.clk(gclk));
	jxor g014(.dina(w_Gid23_0[1]),.dinb(w_Gid19_0[1]),.dout(n87),.clk(gclk));
	jxor g015(.dina(n87),.dinb(n86),.dout(n88),.clk(gclk));
	jand g016(.dina(w_Gr_3[0]),.dinb(Gic7),.dout(n89),.clk(gclk));
	jnot g017(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jxor g018(.dina(n90),.dinb(w_n88_0[1]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_Gid7_0[2]),.dinb(w_Gid6_0[2]),.dout(n92),.clk(gclk));
	jxor g020(.dina(w_Gid5_0[2]),.dinb(w_Gid4_0[1]),.dout(n93),.clk(gclk));
	jxor g021(.dina(n93),.dinb(n92),.dout(n94),.clk(gclk));
	jxor g022(.dina(w_Gid15_0[2]),.dinb(w_Gid14_0[2]),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_Gid13_0[2]),.dinb(w_Gid12_0[1]),.dout(n96),.clk(gclk));
	jxor g024(.dina(n96),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_n97_0[1]),.dinb(w_n94_0[1]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_n98_0[1]),.dinb(n91),.dout(n99),.clk(gclk));
	jxor g027(.dina(w_Gid30_0[2]),.dinb(w_Gid26_0[2]),.dout(n100),.clk(gclk));
	jxor g028(.dina(w_Gid22_0[1]),.dinb(w_Gid18_0[1]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n100),.dout(n102),.clk(gclk));
	jand g030(.dina(w_Gr_2[2]),.dinb(Gic6),.dout(n103),.clk(gclk));
	jxor g031(.dina(w_dff_B_Wmn3ofzU8_0),.dinb(n102),.dout(n104),.clk(gclk));
	jxor g032(.dina(w_Gid3_0[2]),.dinb(w_Gid2_0[2]),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_Gid1_0[2]),.dinb(w_Gid0_0[1]),.dout(n106),.clk(gclk));
	jxor g034(.dina(n106),.dinb(n105),.dout(n107),.clk(gclk));
	jxor g035(.dina(w_Gid11_0[2]),.dinb(w_Gid10_0[2]),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_Gid9_0[2]),.dinb(w_Gid8_0[1]),.dout(n109),.clk(gclk));
	jxor g037(.dina(n109),.dinb(n108),.dout(n110),.clk(gclk));
	jxor g038(.dina(w_n110_0[1]),.dinb(w_n107_0[1]),.dout(n111),.clk(gclk));
	jxor g039(.dina(n111),.dinb(n104),.dout(n112),.clk(gclk));
	jand g040(.dina(w_n112_2[2]),.dinb(w_n99_0[1]),.dout(n113),.clk(gclk));
	jxor g041(.dina(w_Gid13_0[1]),.dinb(w_Gid9_0[1]),.dout(n114),.clk(gclk));
	jxor g042(.dina(w_Gid5_0[1]),.dinb(w_Gid1_0[1]),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jand g044(.dina(w_Gr_2[1]),.dinb(Gic1),.dout(n117),.clk(gclk));
	jxor g045(.dina(w_n117_0[1]),.dinb(w_n116_0[1]),.dout(n118),.clk(gclk));
	jxor g046(.dina(w_Gid31_0[1]),.dinb(w_Gid30_0[1]),.dout(n119),.clk(gclk));
	jxor g047(.dina(w_Gid29_0[2]),.dinb(w_Gid28_0[2]),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(n119),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_Gid27_0[1]),.dinb(w_Gid26_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_Gid25_0[2]),.dinb(w_Gid24_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(w_n124_0[2]),.dinb(w_n121_0[2]),.dout(n125),.clk(gclk));
	jxor g053(.dina(w_n125_0[1]),.dinb(n118),.dout(n126),.clk(gclk));
	jxor g054(.dina(w_n126_2[1]),.dinb(w_n85_2[1]),.dout(n127),.clk(gclk));
	jand g055(.dina(w_Gr_2[0]),.dinb(Gic3),.dout(n128),.clk(gclk));
	jnot g056(.din(w_n128_0[1]),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(w_n121_0[1]),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_Gid15_0[1]),.dinb(w_Gid11_0[1]),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_Gid7_0[1]),.dinb(w_Gid3_0[1]),.dout(n132),.clk(gclk));
	jxor g060(.dina(n132),.dinb(n131),.dout(n133),.clk(gclk));
	jxor g061(.dina(n133),.dinb(w_n83_0[0]),.dout(n134),.clk(gclk));
	jxor g062(.dina(w_n134_0[1]),.dinb(n130),.dout(n135),.clk(gclk));
	jand g063(.dina(w_Gr_1[2]),.dinb(Gic2),.dout(n136),.clk(gclk));
	jnot g064(.din(w_n136_0[1]),.dout(n137),.clk(gclk));
	jxor g065(.dina(n137),.dinb(w_n124_0[1]),.dout(n138),.clk(gclk));
	jxor g066(.dina(w_Gid14_0[1]),.dinb(w_Gid10_0[1]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_Gid6_0[1]),.dinb(w_Gid2_0[1]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g069(.dina(n141),.dinb(w_n80_0[0]),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_n142_0[1]),.dinb(n138),.dout(n143),.clk(gclk));
	jand g071(.dina(w_n143_0[1]),.dinb(w_n135_0[1]),.dout(n144),.clk(gclk));
	jand g072(.dina(n144),.dinb(n127),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_n128_0[0]),.dinb(w_n121_0[0]),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_n134_0[0]),.dinb(n146),.dout(n147),.clk(gclk));
	jxor g075(.dina(w_n136_0[0]),.dinb(w_n124_0[0]),.dout(n148),.clk(gclk));
	jxor g076(.dina(w_n142_0[0]),.dinb(n148),.dout(n149),.clk(gclk));
	jxor g077(.dina(w_n149_2[1]),.dinb(w_n147_2[1]),.dout(n150),.clk(gclk));
	jnot g078(.din(w_n76_0[0]),.dout(n151),.clk(gclk));
	jxor g079(.dina(n151),.dinb(w_n75_0[0]),.dout(n152),.clk(gclk));
	jxor g080(.dina(w_n84_0[0]),.dinb(n152),.dout(n153),.clk(gclk));
	jnot g081(.din(w_n117_0[0]),.dout(n154),.clk(gclk));
	jxor g082(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_n125_0[0]),.dinb(n155),.dout(n156),.clk(gclk));
	jand g084(.dina(w_n156_0[1]),.dinb(w_n153_0[1]),.dout(n157),.clk(gclk));
	jand g085(.dina(n157),.dinb(n150),.dout(n158),.clk(gclk));
	jor g086(.dina(n158),.dinb(n145),.dout(n159),.clk(gclk));
	jxor g087(.dina(w_Gid28_0[1]),.dinb(w_Gid24_0[1]),.dout(n160),.clk(gclk));
	jxor g088(.dina(w_Gid20_0[1]),.dinb(w_Gid16_0[1]),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(n160),.dout(n162),.clk(gclk));
	jand g090(.dina(w_Gr_1[1]),.dinb(Gic4),.dout(n163),.clk(gclk));
	jxor g091(.dina(w_dff_B_u4RzZMEj3_0),.dinb(n162),.dout(n164),.clk(gclk));
	jxor g092(.dina(w_n107_0[0]),.dinb(w_n94_0[0]),.dout(n165),.clk(gclk));
	jxor g093(.dina(n165),.dinb(n164),.dout(n166),.clk(gclk));
	jxor g094(.dina(w_Gid29_0[1]),.dinb(w_Gid25_0[1]),.dout(n167),.clk(gclk));
	jxor g095(.dina(w_Gid21_0[1]),.dinb(w_Gid17_0[1]),.dout(n168),.clk(gclk));
	jxor g096(.dina(n168),.dinb(n167),.dout(n169),.clk(gclk));
	jand g097(.dina(w_Gr_1[0]),.dinb(Gic5),.dout(n170),.clk(gclk));
	jnot g098(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jxor g099(.dina(n171),.dinb(w_n169_0[1]),.dout(n172),.clk(gclk));
	jxor g100(.dina(w_n110_0[0]),.dinb(w_n97_0[0]),.dout(n173),.clk(gclk));
	jxor g101(.dina(w_n173_0[1]),.dinb(n172),.dout(n174),.clk(gclk));
	jand g102(.dina(w_n174_0[1]),.dinb(w_n166_2[2]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_0[1]),.dinb(w_n159_0[2]),.dout(n176),.clk(gclk));
	jand g104(.dina(n176),.dinb(w_n113_0[1]),.dout(n177),.clk(gclk));
	jand g105(.dina(w_n177_1[1]),.dinb(w_n85_2[0]),.dout(n178),.clk(gclk));
	jxor g106(.dina(n178),.dinb(w_Gid0_0[0]),.dout(w_dff_A_PMYQK5Tj0_2),.clk(gclk));
	jand g107(.dina(w_n177_1[0]),.dinb(w_n126_2[0]),.dout(n180),.clk(gclk));
	jxor g108(.dina(n180),.dinb(w_Gid1_0[0]),.dout(w_dff_A_5M6o6Ub95_2),.clk(gclk));
	jand g109(.dina(w_n177_0[2]),.dinb(w_n149_2[0]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_Gid2_0[0]),.dout(w_dff_A_34PC55qj0_2),.clk(gclk));
	jand g111(.dina(w_n177_0[1]),.dinb(w_n147_2[0]),.dout(n184),.clk(gclk));
	jxor g112(.dina(n184),.dinb(w_Gid3_0[0]),.dout(w_dff_A_VTAVybd45_2),.clk(gclk));
	jxor g113(.dina(w_n89_0[0]),.dinb(w_n88_0[0]),.dout(n186),.clk(gclk));
	jxor g114(.dina(w_n98_0[0]),.dinb(n186),.dout(n187),.clk(gclk));
	jnot g115(.din(w_n112_2[1]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n188_0[1]),.dinb(w_n187_2[1]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_dff_B_K1qUrywU9_0),.dinb(w_n159_0[1]),.dout(n190),.clk(gclk));
	jand g118(.dina(w_n190_0[1]),.dinb(w_n175_0[0]),.dout(n191),.clk(gclk));
	jand g119(.dina(w_n191_1[1]),.dinb(w_n85_1[2]),.dout(n192),.clk(gclk));
	jxor g120(.dina(n192),.dinb(w_Gid4_0[0]),.dout(w_dff_A_Fwn0Ij8d6_2),.clk(gclk));
	jand g121(.dina(w_n191_1[0]),.dinb(w_n126_1[2]),.dout(n194),.clk(gclk));
	jxor g122(.dina(n194),.dinb(w_Gid5_0[0]),.dout(w_dff_A_n7m9VX7F7_2),.clk(gclk));
	jand g123(.dina(w_n191_0[2]),.dinb(w_n149_1[2]),.dout(n196),.clk(gclk));
	jxor g124(.dina(n196),.dinb(w_Gid6_0[0]),.dout(w_dff_A_PYCXl0ap5_2),.clk(gclk));
	jand g125(.dina(w_n191_0[1]),.dinb(w_n147_1[2]),.dout(n198),.clk(gclk));
	jxor g126(.dina(n198),.dinb(w_Gid7_0[0]),.dout(w_dff_A_XgvbmHBM3_2),.clk(gclk));
	jnot g127(.din(w_n166_2[1]),.dout(n200),.clk(gclk));
	jxor g128(.dina(w_n170_0[0]),.dinb(w_n169_0[0]),.dout(n201),.clk(gclk));
	jxor g129(.dina(w_n173_0[0]),.dinb(n201),.dout(n202),.clk(gclk));
	jand g130(.dina(w_n202_2[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jand g131(.dina(w_n159_0[0]),.dinb(w_n113_0[0]),.dout(n204),.clk(gclk));
	jand g132(.dina(n204),.dinb(w_n203_0[1]),.dout(n205),.clk(gclk));
	jand g133(.dina(w_n205_1[1]),.dinb(w_n85_1[1]),.dout(n206),.clk(gclk));
	jxor g134(.dina(n206),.dinb(w_Gid8_0[0]),.dout(w_dff_A_SsQEgfrU1_2),.clk(gclk));
	jand g135(.dina(w_n205_1[0]),.dinb(w_n126_1[1]),.dout(n208),.clk(gclk));
	jxor g136(.dina(n208),.dinb(w_Gid9_0[0]),.dout(w_dff_A_P1nnemrt1_2),.clk(gclk));
	jand g137(.dina(w_n205_0[2]),.dinb(w_n149_1[1]),.dout(n210),.clk(gclk));
	jxor g138(.dina(n210),.dinb(w_Gid10_0[0]),.dout(w_dff_A_YC1eikXb3_2),.clk(gclk));
	jand g139(.dina(w_n205_0[1]),.dinb(w_n147_1[1]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_Gid11_0[0]),.dout(w_dff_A_gri3Jqev7_2),.clk(gclk));
	jand g141(.dina(w_n203_0[0]),.dinb(w_n190_0[0]),.dout(n214),.clk(gclk));
	jand g142(.dina(w_n214_1[1]),.dinb(w_n85_1[0]),.dout(n215),.clk(gclk));
	jxor g143(.dina(n215),.dinb(w_Gid12_0[0]),.dout(w_dff_A_wRRP0kLL9_2),.clk(gclk));
	jand g144(.dina(w_n214_1[0]),.dinb(w_n126_1[0]),.dout(n217),.clk(gclk));
	jxor g145(.dina(n217),.dinb(w_Gid13_0[0]),.dout(w_dff_A_4nkykmME2_2),.clk(gclk));
	jand g146(.dina(w_n214_0[2]),.dinb(w_n149_1[0]),.dout(n219),.clk(gclk));
	jxor g147(.dina(n219),.dinb(w_Gid14_0[0]),.dout(w_dff_A_UxhabKGn3_2),.clk(gclk));
	jand g148(.dina(w_n214_0[1]),.dinb(w_n147_1[0]),.dout(n221),.clk(gclk));
	jxor g149(.dina(n221),.dinb(w_Gid15_0[0]),.dout(w_dff_A_7GIr0kJS3_2),.clk(gclk));
	jand g150(.dina(w_n149_0[2]),.dinb(w_n135_0[0]),.dout(n223),.clk(gclk));
	jand g151(.dina(w_n156_0[0]),.dinb(w_n85_0[2]),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n112_2[0]),.dinb(w_n187_2[0]),.dout(n225),.clk(gclk));
	jand g153(.dina(n225),.dinb(w_n174_0[0]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(w_n200_0[0]),.dout(n227),.clk(gclk));
	jxor g155(.dina(w_n202_2[0]),.dinb(w_n166_2[0]),.dout(n228),.clk(gclk));
	jand g156(.dina(n228),.dinb(w_n99_0[0]),.dout(n229),.clk(gclk));
	jand g157(.dina(n229),.dinb(w_n188_0[0]),.dout(n230),.clk(gclk));
	jor g158(.dina(n230),.dinb(n227),.dout(n231),.clk(gclk));
	jand g159(.dina(w_n231_0[1]),.dinb(w_dff_B_ZnGIKCip6_1),.dout(n232),.clk(gclk));
	jand g160(.dina(w_n232_0[1]),.dinb(w_n223_0[1]),.dout(n233),.clk(gclk));
	jand g161(.dina(w_n233_1[1]),.dinb(w_n166_1[2]),.dout(n234),.clk(gclk));
	jxor g162(.dina(n234),.dinb(w_Gid16_0[0]),.dout(God16),.clk(gclk));
	jand g163(.dina(w_n233_1[0]),.dinb(w_n202_1[2]),.dout(n236),.clk(gclk));
	jxor g164(.dina(n236),.dinb(w_Gid17_0[0]),.dout(God17),.clk(gclk));
	jand g165(.dina(w_n233_0[2]),.dinb(w_n112_1[2]),.dout(n238),.clk(gclk));
	jxor g166(.dina(n238),.dinb(w_Gid18_0[0]),.dout(God18),.clk(gclk));
	jand g167(.dina(w_n233_0[1]),.dinb(w_n187_1[2]),.dout(n240),.clk(gclk));
	jxor g168(.dina(n240),.dinb(w_Gid19_0[0]),.dout(God19),.clk(gclk));
	jand g169(.dina(w_n143_0[0]),.dinb(w_n147_0[2]),.dout(n242),.clk(gclk));
	jand g170(.dina(w_n232_0[0]),.dinb(w_n242_0[1]),.dout(n243),.clk(gclk));
	jand g171(.dina(w_n243_1[1]),.dinb(w_n166_1[1]),.dout(n244),.clk(gclk));
	jxor g172(.dina(n244),.dinb(w_Gid20_0[0]),.dout(God20),.clk(gclk));
	jand g173(.dina(w_n243_1[0]),.dinb(w_n202_1[1]),.dout(n246),.clk(gclk));
	jxor g174(.dina(n246),.dinb(w_Gid21_0[0]),.dout(God21),.clk(gclk));
	jand g175(.dina(w_n243_0[2]),.dinb(w_n112_1[1]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_Gid22_0[0]),.dout(God22),.clk(gclk));
	jand g177(.dina(w_n243_0[1]),.dinb(w_n187_1[1]),.dout(n250),.clk(gclk));
	jxor g178(.dina(n250),.dinb(w_Gid23_0[0]),.dout(God23),.clk(gclk));
	jand g179(.dina(w_n126_0[2]),.dinb(w_n153_0[0]),.dout(n252),.clk(gclk));
	jand g180(.dina(w_n231_0[0]),.dinb(w_dff_B_rl6k19680_1),.dout(n253),.clk(gclk));
	jand g181(.dina(w_n253_0[1]),.dinb(w_n223_0[0]),.dout(n254),.clk(gclk));
	jand g182(.dina(w_n254_1[1]),.dinb(w_n166_1[0]),.dout(n255),.clk(gclk));
	jxor g183(.dina(n255),.dinb(w_Gid24_0[0]),.dout(God24),.clk(gclk));
	jand g184(.dina(w_n254_1[0]),.dinb(w_n202_1[0]),.dout(n257),.clk(gclk));
	jxor g185(.dina(n257),.dinb(w_Gid25_0[0]),.dout(God25),.clk(gclk));
	jand g186(.dina(w_n254_0[2]),.dinb(w_n112_1[0]),.dout(n259),.clk(gclk));
	jxor g187(.dina(n259),.dinb(w_Gid26_0[0]),.dout(God26),.clk(gclk));
	jand g188(.dina(w_n254_0[1]),.dinb(w_n187_1[0]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_Gid27_0[0]),.dout(God27),.clk(gclk));
	jand g190(.dina(w_n253_0[0]),.dinb(w_n242_0[0]),.dout(n263),.clk(gclk));
	jand g191(.dina(w_n263_1[1]),.dinb(w_n166_0[2]),.dout(n264),.clk(gclk));
	jxor g192(.dina(n264),.dinb(w_Gid28_0[0]),.dout(God28),.clk(gclk));
	jand g193(.dina(w_n263_1[0]),.dinb(w_n202_0[2]),.dout(n266),.clk(gclk));
	jxor g194(.dina(n266),.dinb(w_Gid29_0[0]),.dout(God29),.clk(gclk));
	jand g195(.dina(w_n263_0[2]),.dinb(w_n112_0[2]),.dout(n268),.clk(gclk));
	jxor g196(.dina(n268),.dinb(w_Gid30_0[0]),.dout(God30),.clk(gclk));
	jand g197(.dina(w_n263_0[1]),.dinb(w_n187_0[2]),.dout(n270),.clk(gclk));
	jxor g198(.dina(n270),.dinb(w_Gid31_0[0]),.dout(God31),.clk(gclk));
	jspl3 jspl3_w_Gid0_0(.douta(w_dff_A_SMk4Rzs98_0),.doutb(w_Gid0_0[1]),.doutc(w_Gid0_0[2]),.din(Gid0));
	jspl3 jspl3_w_Gid1_0(.douta(w_dff_A_P5oWNlu53_0),.doutb(w_Gid1_0[1]),.doutc(w_Gid1_0[2]),.din(Gid1));
	jspl3 jspl3_w_Gid2_0(.douta(w_dff_A_0SJj0lBu8_0),.doutb(w_Gid2_0[1]),.doutc(w_Gid2_0[2]),.din(Gid2));
	jspl3 jspl3_w_Gid3_0(.douta(w_dff_A_vn5rWJvX4_0),.doutb(w_Gid3_0[1]),.doutc(w_Gid3_0[2]),.din(Gid3));
	jspl3 jspl3_w_Gid4_0(.douta(w_dff_A_1r2cNNVA0_0),.doutb(w_Gid4_0[1]),.doutc(w_Gid4_0[2]),.din(Gid4));
	jspl3 jspl3_w_Gid5_0(.douta(w_dff_A_z1gSDu4R5_0),.doutb(w_Gid5_0[1]),.doutc(w_Gid5_0[2]),.din(Gid5));
	jspl3 jspl3_w_Gid6_0(.douta(w_dff_A_5pI5wIum6_0),.doutb(w_Gid6_0[1]),.doutc(w_Gid6_0[2]),.din(Gid6));
	jspl3 jspl3_w_Gid7_0(.douta(w_dff_A_ipJAZuyO5_0),.doutb(w_Gid7_0[1]),.doutc(w_Gid7_0[2]),.din(Gid7));
	jspl3 jspl3_w_Gid8_0(.douta(w_dff_A_lLJru4AI4_0),.doutb(w_Gid8_0[1]),.doutc(w_Gid8_0[2]),.din(Gid8));
	jspl3 jspl3_w_Gid9_0(.douta(w_dff_A_Klm57AT37_0),.doutb(w_Gid9_0[1]),.doutc(w_Gid9_0[2]),.din(Gid9));
	jspl3 jspl3_w_Gid10_0(.douta(w_dff_A_wYS3BdfW6_0),.doutb(w_Gid10_0[1]),.doutc(w_Gid10_0[2]),.din(Gid10));
	jspl3 jspl3_w_Gid11_0(.douta(w_dff_A_DnccThX34_0),.doutb(w_Gid11_0[1]),.doutc(w_Gid11_0[2]),.din(Gid11));
	jspl3 jspl3_w_Gid12_0(.douta(w_dff_A_9wkS9wKr2_0),.doutb(w_Gid12_0[1]),.doutc(w_Gid12_0[2]),.din(Gid12));
	jspl3 jspl3_w_Gid13_0(.douta(w_dff_A_4gDemzTZ7_0),.doutb(w_Gid13_0[1]),.doutc(w_Gid13_0[2]),.din(Gid13));
	jspl3 jspl3_w_Gid14_0(.douta(w_dff_A_LyMrNUTW1_0),.doutb(w_Gid14_0[1]),.doutc(w_Gid14_0[2]),.din(Gid14));
	jspl3 jspl3_w_Gid15_0(.douta(w_dff_A_9kS1c7it8_0),.doutb(w_Gid15_0[1]),.doutc(w_Gid15_0[2]),.din(Gid15));
	jspl3 jspl3_w_Gid16_0(.douta(w_dff_A_DJEzk7og9_0),.doutb(w_Gid16_0[1]),.doutc(w_Gid16_0[2]),.din(Gid16));
	jspl3 jspl3_w_Gid17_0(.douta(w_dff_A_kZnL2V1h6_0),.doutb(w_Gid17_0[1]),.doutc(w_Gid17_0[2]),.din(Gid17));
	jspl3 jspl3_w_Gid18_0(.douta(w_dff_A_VQhWYieE2_0),.doutb(w_Gid18_0[1]),.doutc(w_Gid18_0[2]),.din(Gid18));
	jspl3 jspl3_w_Gid19_0(.douta(w_dff_A_culgjWxi5_0),.doutb(w_Gid19_0[1]),.doutc(w_Gid19_0[2]),.din(Gid19));
	jspl3 jspl3_w_Gid20_0(.douta(w_dff_A_QMFA5xbD2_0),.doutb(w_Gid20_0[1]),.doutc(w_Gid20_0[2]),.din(Gid20));
	jspl3 jspl3_w_Gid21_0(.douta(w_dff_A_OWywckru0_0),.doutb(w_Gid21_0[1]),.doutc(w_Gid21_0[2]),.din(Gid21));
	jspl3 jspl3_w_Gid22_0(.douta(w_dff_A_dDbXMIj37_0),.doutb(w_Gid22_0[1]),.doutc(w_Gid22_0[2]),.din(Gid22));
	jspl3 jspl3_w_Gid23_0(.douta(w_dff_A_MdgH81Vo4_0),.doutb(w_Gid23_0[1]),.doutc(w_Gid23_0[2]),.din(Gid23));
	jspl3 jspl3_w_Gid24_0(.douta(w_dff_A_JDtv5Dbc7_0),.doutb(w_Gid24_0[1]),.doutc(w_Gid24_0[2]),.din(Gid24));
	jspl3 jspl3_w_Gid25_0(.douta(w_dff_A_I8rUbnB55_0),.doutb(w_Gid25_0[1]),.doutc(w_Gid25_0[2]),.din(Gid25));
	jspl3 jspl3_w_Gid26_0(.douta(w_dff_A_TQHmocMZ4_0),.doutb(w_Gid26_0[1]),.doutc(w_Gid26_0[2]),.din(Gid26));
	jspl3 jspl3_w_Gid27_0(.douta(w_dff_A_VCEw40Ni6_0),.doutb(w_Gid27_0[1]),.doutc(w_Gid27_0[2]),.din(Gid27));
	jspl3 jspl3_w_Gid28_0(.douta(w_dff_A_C0FtiK1q2_0),.doutb(w_Gid28_0[1]),.doutc(w_Gid28_0[2]),.din(Gid28));
	jspl3 jspl3_w_Gid29_0(.douta(w_dff_A_azHUBSfr1_0),.doutb(w_Gid29_0[1]),.doutc(w_Gid29_0[2]),.din(Gid29));
	jspl3 jspl3_w_Gid30_0(.douta(w_dff_A_iJKwPfTv6_0),.doutb(w_Gid30_0[1]),.doutc(w_Gid30_0[2]),.din(Gid30));
	jspl3 jspl3_w_Gid31_0(.douta(w_dff_A_ErCKavnX3_0),.doutb(w_Gid31_0[1]),.doutc(w_Gid31_0[2]),.din(Gid31));
	jspl3 jspl3_w_Gr_0(.douta(w_Gr_0[0]),.doutb(w_Gr_0[1]),.doutc(w_Gr_0[2]),.din(Gr));
	jspl3 jspl3_w_Gr_1(.douta(w_Gr_1[0]),.doutb(w_Gr_1[1]),.doutc(w_Gr_1[2]),.din(w_Gr_0[0]));
	jspl3 jspl3_w_Gr_2(.douta(w_Gr_2[0]),.doutb(w_Gr_2[1]),.doutc(w_Gr_2[2]),.din(w_Gr_0[1]));
	jspl jspl_w_Gr_3(.douta(w_Gr_3[0]),.doutb(w_Gr_3[1]),.din(w_Gr_0[2]));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_dff_A_nRbvuv8M9_1),.din(n76));
	jspl jspl_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_ItvWWmwT7_0),.doutb(w_n85_0[1]),.doutc(w_n85_0[2]),.din(n85));
	jspl3 jspl3_w_n85_1(.douta(w_n85_1[0]),.doutb(w_n85_1[1]),.doutc(w_n85_1[2]),.din(w_n85_0[0]));
	jspl jspl_w_n85_2(.douta(w_dff_A_AcoMs2LU8_0),.doutb(w_n85_2[1]),.din(w_n85_0[1]));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n89_0(.douta(w_dff_A_QKvtC1f67_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_dff_A_ykLkWruT0_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_vQpDA4Vz2_0),.doutb(w_n112_0[1]),.doutc(w_dff_A_ohv5oZ1X2_2),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_dff_A_6GE9eT2e6_1),.din(w_dff_B_PvPK2uh24_2));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.din(n116));
	jspl jspl_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_QSOiowHf1_1),.din(n117));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.doutc(w_n124_0[2]),.din(n124));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_KkUIyz2i2_0),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl3 jspl3_w_n126_1(.douta(w_n126_1[0]),.doutb(w_n126_1[1]),.doutc(w_n126_1[2]),.din(w_n126_0[0]));
	jspl jspl_w_n126_2(.douta(w_dff_A_Yz4tRNK61_0),.doutb(w_n126_2[1]),.din(w_n126_0[1]));
	jspl jspl_w_n128_0(.douta(w_dff_A_ieHKHVNB2_0),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n134_0(.douta(w_n134_0[0]),.doutb(w_n134_0[1]),.din(n134));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n136_0(.douta(w_dff_A_9ma5OEpZ6_0),.doutb(w_n136_0[1]),.din(n136));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl3 jspl3_w_n147_0(.douta(w_dff_A_UsLC33ks8_0),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n147_1(.douta(w_n147_1[0]),.doutb(w_n147_1[1]),.doutc(w_n147_1[2]),.din(w_n147_0[0]));
	jspl jspl_w_n147_2(.douta(w_dff_A_zKRcJdAD1_0),.doutb(w_n147_2[1]),.din(w_n147_0[1]));
	jspl3 jspl3_w_n149_0(.douta(w_dff_A_Pwr49xPF5_0),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_n149_1[1]),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_BpR7RP2O6_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl jspl_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.din(n153));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl3 jspl3_w_n166_0(.douta(w_dff_A_FFGOan2N3_0),.doutb(w_n166_0[1]),.doutc(w_dff_A_uzwkQZ2I5_2),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.doutc(w_n166_1[2]),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_n166_2[2]),.din(w_n166_0[1]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_dff_A_4kVdwhdl2_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl jspl_w_n174_0(.douta(w_dff_A_mneKHFDU5_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_dff_A_aDdyPWb38_0),.doutb(w_n175_0[1]),.din(w_dff_B_QzVgACRg1_2));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl jspl_w_n177_1(.douta(w_n177_1[0]),.doutb(w_n177_1[1]),.din(w_n177_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_dff_A_HCBrWaSp5_0),.doutb(w_n187_0[1]),.doutc(w_dff_A_XhUlaSPc8_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_n187_1[0]),.doutb(w_n187_1[1]),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n187_2(.douta(w_n187_2[0]),.doutb(w_dff_A_BlxLJbn71_1),.din(w_n187_0[1]));
	jspl jspl_w_n188_0(.douta(w_dff_A_QOKelfPT2_0),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n191_1(.douta(w_n191_1[0]),.doutb(w_n191_1[1]),.din(w_n191_0[0]));
	jspl jspl_w_n200_0(.douta(w_dff_A_sDuJvpTu9_0),.doutb(w_n200_0[1]),.din(n200));
	jspl3 jspl3_w_n202_0(.douta(w_dff_A_cxvYa9bb2_0),.doutb(w_n202_0[1]),.doutc(w_dff_A_gCAR8UGY4_2),.din(n202));
	jspl3 jspl3_w_n202_1(.douta(w_n202_1[0]),.doutb(w_n202_1[1]),.doutc(w_n202_1[2]),.din(w_n202_0[0]));
	jspl jspl_w_n202_2(.douta(w_n202_2[0]),.doutb(w_dff_A_dRHQyIA50_1),.din(w_n202_0[1]));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(w_dff_B_u6YsHwn04_2));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(n205));
	jspl jspl_w_n205_1(.douta(w_n205_1[0]),.doutb(w_n205_1[1]),.din(w_n205_0[0]));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl jspl_w_n214_1(.douta(w_n214_1[0]),.doutb(w_n214_1[1]),.din(w_n214_0[0]));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.din(w_dff_B_1bGkhgnf2_2));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(w_dff_B_d6TFRYE03_2));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n243_1(.douta(w_n243_1[0]),.doutb(w_n243_1[1]),.din(w_n243_0[0]));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.doutc(w_n263_0[2]),.din(n263));
	jspl jspl_w_n263_1(.douta(w_n263_1[0]),.doutb(w_n263_1[1]),.din(w_n263_0[0]));
	jdff dff_A_aDdyPWb38_0(.dout(w_n175_0[0]),.din(w_dff_A_aDdyPWb38_0),.clk(gclk));
	jdff dff_B_rcJR4sP54_2(.din(n175),.dout(w_dff_B_rcJR4sP54_2),.clk(gclk));
	jdff dff_B_QzVgACRg1_2(.din(w_dff_B_rcJR4sP54_2),.dout(w_dff_B_QzVgACRg1_2),.clk(gclk));
	jdff dff_A_6GE9eT2e6_1(.dout(w_n113_0[1]),.din(w_dff_A_6GE9eT2e6_1),.clk(gclk));
	jdff dff_B_Bv2Pjeql0_2(.din(n113),.dout(w_dff_B_Bv2Pjeql0_2),.clk(gclk));
	jdff dff_B_PvPK2uh24_2(.din(w_dff_B_Bv2Pjeql0_2),.dout(w_dff_B_PvPK2uh24_2),.clk(gclk));
	jdff dff_B_U6YQwxGQ5_2(.din(n203),.dout(w_dff_B_U6YQwxGQ5_2),.clk(gclk));
	jdff dff_B_u6YsHwn04_2(.din(w_dff_B_U6YQwxGQ5_2),.dout(w_dff_B_u6YsHwn04_2),.clk(gclk));
	jdff dff_B_K1qUrywU9_0(.din(n189),.dout(w_dff_B_K1qUrywU9_0),.clk(gclk));
	jdff dff_A_vYm9ffK76_0(.dout(w_n149_2[0]),.din(w_dff_A_vYm9ffK76_0),.clk(gclk));
	jdff dff_A_8m7vKhDh8_0(.dout(w_dff_A_vYm9ffK76_0),.din(w_dff_A_8m7vKhDh8_0),.clk(gclk));
	jdff dff_A_jTKP7wBN4_0(.dout(w_dff_A_8m7vKhDh8_0),.din(w_dff_A_jTKP7wBN4_0),.clk(gclk));
	jdff dff_A_rdAhtn6n6_0(.dout(w_dff_A_jTKP7wBN4_0),.din(w_dff_A_rdAhtn6n6_0),.clk(gclk));
	jdff dff_A_BpR7RP2O6_0(.dout(w_dff_A_rdAhtn6n6_0),.din(w_dff_A_BpR7RP2O6_0),.clk(gclk));
	jdff dff_A_IaMk4a494_0(.dout(w_n147_2[0]),.din(w_dff_A_IaMk4a494_0),.clk(gclk));
	jdff dff_A_tz9wkayk6_0(.dout(w_dff_A_IaMk4a494_0),.din(w_dff_A_tz9wkayk6_0),.clk(gclk));
	jdff dff_A_8CAR0Ip75_0(.dout(w_dff_A_tz9wkayk6_0),.din(w_dff_A_8CAR0Ip75_0),.clk(gclk));
	jdff dff_A_nA7QdfNz7_0(.dout(w_dff_A_8CAR0Ip75_0),.din(w_dff_A_nA7QdfNz7_0),.clk(gclk));
	jdff dff_A_zKRcJdAD1_0(.dout(w_dff_A_nA7QdfNz7_0),.din(w_dff_A_zKRcJdAD1_0),.clk(gclk));
	jdff dff_A_0QEC5RPS1_0(.dout(w_n126_2[0]),.din(w_dff_A_0QEC5RPS1_0),.clk(gclk));
	jdff dff_A_rNaUt7z90_0(.dout(w_dff_A_0QEC5RPS1_0),.din(w_dff_A_rNaUt7z90_0),.clk(gclk));
	jdff dff_A_oWVKbCJm2_0(.dout(w_dff_A_rNaUt7z90_0),.din(w_dff_A_oWVKbCJm2_0),.clk(gclk));
	jdff dff_A_njpK3b4y3_0(.dout(w_dff_A_oWVKbCJm2_0),.din(w_dff_A_njpK3b4y3_0),.clk(gclk));
	jdff dff_A_Yz4tRNK61_0(.dout(w_dff_A_njpK3b4y3_0),.din(w_dff_A_Yz4tRNK61_0),.clk(gclk));
	jdff dff_A_MXWJnoX17_0(.dout(w_n85_2[0]),.din(w_dff_A_MXWJnoX17_0),.clk(gclk));
	jdff dff_A_4XJDLIu03_0(.dout(w_dff_A_MXWJnoX17_0),.din(w_dff_A_4XJDLIu03_0),.clk(gclk));
	jdff dff_A_gz9d8heg8_0(.dout(w_dff_A_4XJDLIu03_0),.din(w_dff_A_gz9d8heg8_0),.clk(gclk));
	jdff dff_A_xlqmfJVf2_0(.dout(w_dff_A_gz9d8heg8_0),.din(w_dff_A_xlqmfJVf2_0),.clk(gclk));
	jdff dff_A_AcoMs2LU8_0(.dout(w_dff_A_xlqmfJVf2_0),.din(w_dff_A_AcoMs2LU8_0),.clk(gclk));
	jdff dff_B_aFKaFGhu2_1(.din(n224),.dout(w_dff_B_aFKaFGhu2_1),.clk(gclk));
	jdff dff_B_eq9fE1rP2_1(.din(w_dff_B_aFKaFGhu2_1),.dout(w_dff_B_eq9fE1rP2_1),.clk(gclk));
	jdff dff_B_ZnGIKCip6_1(.din(w_dff_B_eq9fE1rP2_1),.dout(w_dff_B_ZnGIKCip6_1),.clk(gclk));
	jdff dff_A_Lcf74BXH1_0(.dout(w_n85_0[0]),.din(w_dff_A_Lcf74BXH1_0),.clk(gclk));
	jdff dff_A_yQRXNvKO5_0(.dout(w_dff_A_Lcf74BXH1_0),.din(w_dff_A_yQRXNvKO5_0),.clk(gclk));
	jdff dff_A_GNcnHxCq3_0(.dout(w_dff_A_yQRXNvKO5_0),.din(w_dff_A_GNcnHxCq3_0),.clk(gclk));
	jdff dff_A_kTdAH3H60_0(.dout(w_dff_A_GNcnHxCq3_0),.din(w_dff_A_kTdAH3H60_0),.clk(gclk));
	jdff dff_A_ItvWWmwT7_0(.dout(w_dff_A_kTdAH3H60_0),.din(w_dff_A_ItvWWmwT7_0),.clk(gclk));
	jdff dff_B_Ae8t9VTK3_2(.din(n223),.dout(w_dff_B_Ae8t9VTK3_2),.clk(gclk));
	jdff dff_B_dfkZpVnf5_2(.din(w_dff_B_Ae8t9VTK3_2),.dout(w_dff_B_dfkZpVnf5_2),.clk(gclk));
	jdff dff_B_HHc0DKmb7_2(.din(w_dff_B_dfkZpVnf5_2),.dout(w_dff_B_HHc0DKmb7_2),.clk(gclk));
	jdff dff_B_1bGkhgnf2_2(.din(w_dff_B_HHc0DKmb7_2),.dout(w_dff_B_1bGkhgnf2_2),.clk(gclk));
	jdff dff_A_y8WsmTur5_0(.dout(w_n149_0[0]),.din(w_dff_A_y8WsmTur5_0),.clk(gclk));
	jdff dff_A_B6YCX7mG2_0(.dout(w_dff_A_y8WsmTur5_0),.din(w_dff_A_B6YCX7mG2_0),.clk(gclk));
	jdff dff_A_2feKF3Zk2_0(.dout(w_dff_A_B6YCX7mG2_0),.din(w_dff_A_2feKF3Zk2_0),.clk(gclk));
	jdff dff_A_FK9RJOmj1_0(.dout(w_dff_A_2feKF3Zk2_0),.din(w_dff_A_FK9RJOmj1_0),.clk(gclk));
	jdff dff_A_Pwr49xPF5_0(.dout(w_dff_A_FK9RJOmj1_0),.din(w_dff_A_Pwr49xPF5_0),.clk(gclk));
	jdff dff_B_hESeV1NC0_1(.din(n252),.dout(w_dff_B_hESeV1NC0_1),.clk(gclk));
	jdff dff_B_LSyfilou3_1(.din(w_dff_B_hESeV1NC0_1),.dout(w_dff_B_LSyfilou3_1),.clk(gclk));
	jdff dff_B_rl6k19680_1(.din(w_dff_B_LSyfilou3_1),.dout(w_dff_B_rl6k19680_1),.clk(gclk));
	jdff dff_A_dRHQyIA50_1(.dout(w_n202_2[1]),.din(w_dff_A_dRHQyIA50_1),.clk(gclk));
	jdff dff_A_66PxB4UL7_0(.dout(w_n202_0[0]),.din(w_dff_A_66PxB4UL7_0),.clk(gclk));
	jdff dff_A_fBWtJRhz3_0(.dout(w_dff_A_66PxB4UL7_0),.din(w_dff_A_fBWtJRhz3_0),.clk(gclk));
	jdff dff_A_zuwmcgl61_0(.dout(w_dff_A_fBWtJRhz3_0),.din(w_dff_A_zuwmcgl61_0),.clk(gclk));
	jdff dff_A_ZCoSJqDL0_0(.dout(w_dff_A_zuwmcgl61_0),.din(w_dff_A_ZCoSJqDL0_0),.clk(gclk));
	jdff dff_A_HPvauYvh8_0(.dout(w_dff_A_ZCoSJqDL0_0),.din(w_dff_A_HPvauYvh8_0),.clk(gclk));
	jdff dff_A_cxvYa9bb2_0(.dout(w_dff_A_HPvauYvh8_0),.din(w_dff_A_cxvYa9bb2_0),.clk(gclk));
	jdff dff_A_NDutoFw33_2(.dout(w_n202_0[2]),.din(w_dff_A_NDutoFw33_2),.clk(gclk));
	jdff dff_A_e1EDB06P4_2(.dout(w_dff_A_NDutoFw33_2),.din(w_dff_A_e1EDB06P4_2),.clk(gclk));
	jdff dff_A_4IkPgO2g2_2(.dout(w_dff_A_e1EDB06P4_2),.din(w_dff_A_4IkPgO2g2_2),.clk(gclk));
	jdff dff_A_ZzQbgp3B2_2(.dout(w_dff_A_4IkPgO2g2_2),.din(w_dff_A_ZzQbgp3B2_2),.clk(gclk));
	jdff dff_A_ksU8C2KW5_2(.dout(w_dff_A_ZzQbgp3B2_2),.din(w_dff_A_ksU8C2KW5_2),.clk(gclk));
	jdff dff_A_gCAR8UGY4_2(.dout(w_dff_A_ksU8C2KW5_2),.din(w_dff_A_gCAR8UGY4_2),.clk(gclk));
	jdff dff_A_ykLkWruT0_0(.dout(w_n99_0[0]),.din(w_dff_A_ykLkWruT0_0),.clk(gclk));
	jdff dff_A_QOKelfPT2_0(.dout(w_n188_0[0]),.din(w_dff_A_QOKelfPT2_0),.clk(gclk));
	jdff dff_A_JyJpomq77_0(.dout(w_n112_0[0]),.din(w_dff_A_JyJpomq77_0),.clk(gclk));
	jdff dff_A_2i641phh3_0(.dout(w_dff_A_JyJpomq77_0),.din(w_dff_A_2i641phh3_0),.clk(gclk));
	jdff dff_A_YPAYDX9B4_0(.dout(w_dff_A_2i641phh3_0),.din(w_dff_A_YPAYDX9B4_0),.clk(gclk));
	jdff dff_A_jiBeYxFr6_0(.dout(w_dff_A_YPAYDX9B4_0),.din(w_dff_A_jiBeYxFr6_0),.clk(gclk));
	jdff dff_A_wddZOLmr2_0(.dout(w_dff_A_jiBeYxFr6_0),.din(w_dff_A_wddZOLmr2_0),.clk(gclk));
	jdff dff_A_vQpDA4Vz2_0(.dout(w_dff_A_wddZOLmr2_0),.din(w_dff_A_vQpDA4Vz2_0),.clk(gclk));
	jdff dff_A_7REOox3M7_2(.dout(w_n112_0[2]),.din(w_dff_A_7REOox3M7_2),.clk(gclk));
	jdff dff_A_EJ3WYniq1_2(.dout(w_dff_A_7REOox3M7_2),.din(w_dff_A_EJ3WYniq1_2),.clk(gclk));
	jdff dff_A_qqG1XOGj3_2(.dout(w_dff_A_EJ3WYniq1_2),.din(w_dff_A_qqG1XOGj3_2),.clk(gclk));
	jdff dff_A_Mwo6TomW6_2(.dout(w_dff_A_qqG1XOGj3_2),.din(w_dff_A_Mwo6TomW6_2),.clk(gclk));
	jdff dff_A_yYXSBgGe6_2(.dout(w_dff_A_Mwo6TomW6_2),.din(w_dff_A_yYXSBgGe6_2),.clk(gclk));
	jdff dff_A_ohv5oZ1X2_2(.dout(w_dff_A_yYXSBgGe6_2),.din(w_dff_A_ohv5oZ1X2_2),.clk(gclk));
	jdff dff_B_Wmn3ofzU8_0(.din(n103),.dout(w_dff_B_Wmn3ofzU8_0),.clk(gclk));
	jdff dff_A_BlxLJbn71_1(.dout(w_n187_2[1]),.din(w_dff_A_BlxLJbn71_1),.clk(gclk));
	jdff dff_A_DI3JYTHQ3_0(.dout(w_n187_0[0]),.din(w_dff_A_DI3JYTHQ3_0),.clk(gclk));
	jdff dff_A_Hm5n4ftz9_0(.dout(w_dff_A_DI3JYTHQ3_0),.din(w_dff_A_Hm5n4ftz9_0),.clk(gclk));
	jdff dff_A_ipGqDGh94_0(.dout(w_dff_A_Hm5n4ftz9_0),.din(w_dff_A_ipGqDGh94_0),.clk(gclk));
	jdff dff_A_8HehDjDy2_0(.dout(w_dff_A_ipGqDGh94_0),.din(w_dff_A_8HehDjDy2_0),.clk(gclk));
	jdff dff_A_O9Bze4Dq9_0(.dout(w_dff_A_8HehDjDy2_0),.din(w_dff_A_O9Bze4Dq9_0),.clk(gclk));
	jdff dff_A_HCBrWaSp5_0(.dout(w_dff_A_O9Bze4Dq9_0),.din(w_dff_A_HCBrWaSp5_0),.clk(gclk));
	jdff dff_A_x0x1Am6P9_2(.dout(w_n187_0[2]),.din(w_dff_A_x0x1Am6P9_2),.clk(gclk));
	jdff dff_A_cSpIwoL75_2(.dout(w_dff_A_x0x1Am6P9_2),.din(w_dff_A_cSpIwoL75_2),.clk(gclk));
	jdff dff_A_j6NDuhV37_2(.dout(w_dff_A_cSpIwoL75_2),.din(w_dff_A_j6NDuhV37_2),.clk(gclk));
	jdff dff_A_nhBJw5ZR7_2(.dout(w_dff_A_j6NDuhV37_2),.din(w_dff_A_nhBJw5ZR7_2),.clk(gclk));
	jdff dff_A_uGMXUnrz9_2(.dout(w_dff_A_nhBJw5ZR7_2),.din(w_dff_A_uGMXUnrz9_2),.clk(gclk));
	jdff dff_A_XhUlaSPc8_2(.dout(w_dff_A_uGMXUnrz9_2),.din(w_dff_A_XhUlaSPc8_2),.clk(gclk));
	jdff dff_A_QKvtC1f67_0(.dout(w_n89_0[0]),.din(w_dff_A_QKvtC1f67_0),.clk(gclk));
	jdff dff_A_mneKHFDU5_0(.dout(w_n174_0[0]),.din(w_dff_A_mneKHFDU5_0),.clk(gclk));
	jdff dff_A_4kVdwhdl2_0(.dout(w_n170_0[0]),.din(w_dff_A_4kVdwhdl2_0),.clk(gclk));
	jdff dff_A_sDuJvpTu9_0(.dout(w_n200_0[0]),.din(w_dff_A_sDuJvpTu9_0),.clk(gclk));
	jdff dff_A_e4GOGSkB8_0(.dout(w_n166_0[0]),.din(w_dff_A_e4GOGSkB8_0),.clk(gclk));
	jdff dff_A_HFfemwmf6_0(.dout(w_dff_A_e4GOGSkB8_0),.din(w_dff_A_HFfemwmf6_0),.clk(gclk));
	jdff dff_A_KBcOM4Jl7_0(.dout(w_dff_A_HFfemwmf6_0),.din(w_dff_A_KBcOM4Jl7_0),.clk(gclk));
	jdff dff_A_shjmP9hR0_0(.dout(w_dff_A_KBcOM4Jl7_0),.din(w_dff_A_shjmP9hR0_0),.clk(gclk));
	jdff dff_A_ZBVWvipt1_0(.dout(w_dff_A_shjmP9hR0_0),.din(w_dff_A_ZBVWvipt1_0),.clk(gclk));
	jdff dff_A_FFGOan2N3_0(.dout(w_dff_A_ZBVWvipt1_0),.din(w_dff_A_FFGOan2N3_0),.clk(gclk));
	jdff dff_A_PrYQ8vk06_2(.dout(w_n166_0[2]),.din(w_dff_A_PrYQ8vk06_2),.clk(gclk));
	jdff dff_A_HspB0UhW9_2(.dout(w_dff_A_PrYQ8vk06_2),.din(w_dff_A_HspB0UhW9_2),.clk(gclk));
	jdff dff_A_Y6koNCAW7_2(.dout(w_dff_A_HspB0UhW9_2),.din(w_dff_A_Y6koNCAW7_2),.clk(gclk));
	jdff dff_A_5bUNF2l39_2(.dout(w_dff_A_Y6koNCAW7_2),.din(w_dff_A_5bUNF2l39_2),.clk(gclk));
	jdff dff_A_MRD4AoNy9_2(.dout(w_dff_A_5bUNF2l39_2),.din(w_dff_A_MRD4AoNy9_2),.clk(gclk));
	jdff dff_A_uzwkQZ2I5_2(.dout(w_dff_A_MRD4AoNy9_2),.din(w_dff_A_uzwkQZ2I5_2),.clk(gclk));
	jdff dff_B_u4RzZMEj3_0(.din(n163),.dout(w_dff_B_u4RzZMEj3_0),.clk(gclk));
	jdff dff_A_JE9A9tqp1_0(.dout(w_n126_0[0]),.din(w_dff_A_JE9A9tqp1_0),.clk(gclk));
	jdff dff_A_v3ut1IpA9_0(.dout(w_dff_A_JE9A9tqp1_0),.din(w_dff_A_v3ut1IpA9_0),.clk(gclk));
	jdff dff_A_CwaotxFj9_0(.dout(w_dff_A_v3ut1IpA9_0),.din(w_dff_A_CwaotxFj9_0),.clk(gclk));
	jdff dff_A_JATZXH7W9_0(.dout(w_dff_A_CwaotxFj9_0),.din(w_dff_A_JATZXH7W9_0),.clk(gclk));
	jdff dff_A_KkUIyz2i2_0(.dout(w_dff_A_JATZXH7W9_0),.din(w_dff_A_KkUIyz2i2_0),.clk(gclk));
	jdff dff_A_QSOiowHf1_1(.dout(w_n117_0[1]),.din(w_dff_A_QSOiowHf1_1),.clk(gclk));
	jdff dff_A_BFwUrL8z7_0(.dout(w_Gid5_0[0]),.din(w_dff_A_BFwUrL8z7_0),.clk(gclk));
	jdff dff_A_zXBYBGc16_0(.dout(w_dff_A_BFwUrL8z7_0),.din(w_dff_A_zXBYBGc16_0),.clk(gclk));
	jdff dff_A_iFM7iU6v1_0(.dout(w_dff_A_zXBYBGc16_0),.din(w_dff_A_iFM7iU6v1_0),.clk(gclk));
	jdff dff_A_Hxu5YBEq6_0(.dout(w_dff_A_iFM7iU6v1_0),.din(w_dff_A_Hxu5YBEq6_0),.clk(gclk));
	jdff dff_A_kx1wugWw2_0(.dout(w_dff_A_Hxu5YBEq6_0),.din(w_dff_A_kx1wugWw2_0),.clk(gclk));
	jdff dff_A_VvM6vgff7_0(.dout(w_dff_A_kx1wugWw2_0),.din(w_dff_A_VvM6vgff7_0),.clk(gclk));
	jdff dff_A_r58lH3V02_0(.dout(w_dff_A_VvM6vgff7_0),.din(w_dff_A_r58lH3V02_0),.clk(gclk));
	jdff dff_A_wCD0Yq4R2_0(.dout(w_dff_A_r58lH3V02_0),.din(w_dff_A_wCD0Yq4R2_0),.clk(gclk));
	jdff dff_A_UDu7eOFq7_0(.dout(w_dff_A_wCD0Yq4R2_0),.din(w_dff_A_UDu7eOFq7_0),.clk(gclk));
	jdff dff_A_z1gSDu4R5_0(.dout(w_dff_A_UDu7eOFq7_0),.din(w_dff_A_z1gSDu4R5_0),.clk(gclk));
	jdff dff_A_TPnZuobl3_0(.dout(w_Gid1_0[0]),.din(w_dff_A_TPnZuobl3_0),.clk(gclk));
	jdff dff_A_GQByEKuD8_0(.dout(w_dff_A_TPnZuobl3_0),.din(w_dff_A_GQByEKuD8_0),.clk(gclk));
	jdff dff_A_jbxrsE4h6_0(.dout(w_dff_A_GQByEKuD8_0),.din(w_dff_A_jbxrsE4h6_0),.clk(gclk));
	jdff dff_A_xMBmPMU74_0(.dout(w_dff_A_jbxrsE4h6_0),.din(w_dff_A_xMBmPMU74_0),.clk(gclk));
	jdff dff_A_4xZOwaeg3_0(.dout(w_dff_A_xMBmPMU74_0),.din(w_dff_A_4xZOwaeg3_0),.clk(gclk));
	jdff dff_A_lJ1zL3Ms5_0(.dout(w_dff_A_4xZOwaeg3_0),.din(w_dff_A_lJ1zL3Ms5_0),.clk(gclk));
	jdff dff_A_9CVvwYn06_0(.dout(w_dff_A_lJ1zL3Ms5_0),.din(w_dff_A_9CVvwYn06_0),.clk(gclk));
	jdff dff_A_KRopvc4R2_0(.dout(w_dff_A_9CVvwYn06_0),.din(w_dff_A_KRopvc4R2_0),.clk(gclk));
	jdff dff_A_M4plUTxg3_0(.dout(w_dff_A_KRopvc4R2_0),.din(w_dff_A_M4plUTxg3_0),.clk(gclk));
	jdff dff_A_P5oWNlu53_0(.dout(w_dff_A_M4plUTxg3_0),.din(w_dff_A_P5oWNlu53_0),.clk(gclk));
	jdff dff_A_i01bXCXd8_0(.dout(w_Gid13_0[0]),.din(w_dff_A_i01bXCXd8_0),.clk(gclk));
	jdff dff_A_P9mIro7b7_0(.dout(w_dff_A_i01bXCXd8_0),.din(w_dff_A_P9mIro7b7_0),.clk(gclk));
	jdff dff_A_Bz7PX8Da4_0(.dout(w_dff_A_P9mIro7b7_0),.din(w_dff_A_Bz7PX8Da4_0),.clk(gclk));
	jdff dff_A_AqmayLVM3_0(.dout(w_dff_A_Bz7PX8Da4_0),.din(w_dff_A_AqmayLVM3_0),.clk(gclk));
	jdff dff_A_FCqsPleW6_0(.dout(w_dff_A_AqmayLVM3_0),.din(w_dff_A_FCqsPleW6_0),.clk(gclk));
	jdff dff_A_HoLhvVbY8_0(.dout(w_dff_A_FCqsPleW6_0),.din(w_dff_A_HoLhvVbY8_0),.clk(gclk));
	jdff dff_A_sM694yDn0_0(.dout(w_dff_A_HoLhvVbY8_0),.din(w_dff_A_sM694yDn0_0),.clk(gclk));
	jdff dff_A_oAfJG4058_0(.dout(w_dff_A_sM694yDn0_0),.din(w_dff_A_oAfJG4058_0),.clk(gclk));
	jdff dff_A_vPyibuVt2_0(.dout(w_dff_A_oAfJG4058_0),.din(w_dff_A_vPyibuVt2_0),.clk(gclk));
	jdff dff_A_4gDemzTZ7_0(.dout(w_dff_A_vPyibuVt2_0),.din(w_dff_A_4gDemzTZ7_0),.clk(gclk));
	jdff dff_A_wAzpbYQS3_0(.dout(w_Gid9_0[0]),.din(w_dff_A_wAzpbYQS3_0),.clk(gclk));
	jdff dff_A_bFF7kmy35_0(.dout(w_dff_A_wAzpbYQS3_0),.din(w_dff_A_bFF7kmy35_0),.clk(gclk));
	jdff dff_A_8NOL1TLa2_0(.dout(w_dff_A_bFF7kmy35_0),.din(w_dff_A_8NOL1TLa2_0),.clk(gclk));
	jdff dff_A_NPj9osNJ3_0(.dout(w_dff_A_8NOL1TLa2_0),.din(w_dff_A_NPj9osNJ3_0),.clk(gclk));
	jdff dff_A_XzXrlRO07_0(.dout(w_dff_A_NPj9osNJ3_0),.din(w_dff_A_XzXrlRO07_0),.clk(gclk));
	jdff dff_A_yzRbYqvA2_0(.dout(w_dff_A_XzXrlRO07_0),.din(w_dff_A_yzRbYqvA2_0),.clk(gclk));
	jdff dff_A_YnV5BC8T0_0(.dout(w_dff_A_yzRbYqvA2_0),.din(w_dff_A_YnV5BC8T0_0),.clk(gclk));
	jdff dff_A_Wln0iari3_0(.dout(w_dff_A_YnV5BC8T0_0),.din(w_dff_A_Wln0iari3_0),.clk(gclk));
	jdff dff_A_iQnEU6171_0(.dout(w_dff_A_Wln0iari3_0),.din(w_dff_A_iQnEU6171_0),.clk(gclk));
	jdff dff_A_Klm57AT37_0(.dout(w_dff_A_iQnEU6171_0),.din(w_dff_A_Klm57AT37_0),.clk(gclk));
	jdff dff_A_nRbvuv8M9_1(.dout(w_n76_0[1]),.din(w_dff_A_nRbvuv8M9_1),.clk(gclk));
	jdff dff_A_hAVEAOku5_0(.dout(w_Gid4_0[0]),.din(w_dff_A_hAVEAOku5_0),.clk(gclk));
	jdff dff_A_GvIgEcnP9_0(.dout(w_dff_A_hAVEAOku5_0),.din(w_dff_A_GvIgEcnP9_0),.clk(gclk));
	jdff dff_A_Te3X00v68_0(.dout(w_dff_A_GvIgEcnP9_0),.din(w_dff_A_Te3X00v68_0),.clk(gclk));
	jdff dff_A_q5Yf0Vyz3_0(.dout(w_dff_A_Te3X00v68_0),.din(w_dff_A_q5Yf0Vyz3_0),.clk(gclk));
	jdff dff_A_8DPc9Uzb7_0(.dout(w_dff_A_q5Yf0Vyz3_0),.din(w_dff_A_8DPc9Uzb7_0),.clk(gclk));
	jdff dff_A_wUv7iXPn9_0(.dout(w_dff_A_8DPc9Uzb7_0),.din(w_dff_A_wUv7iXPn9_0),.clk(gclk));
	jdff dff_A_9ubRGCaK3_0(.dout(w_dff_A_wUv7iXPn9_0),.din(w_dff_A_9ubRGCaK3_0),.clk(gclk));
	jdff dff_A_HABd7t814_0(.dout(w_dff_A_9ubRGCaK3_0),.din(w_dff_A_HABd7t814_0),.clk(gclk));
	jdff dff_A_x9baV45f4_0(.dout(w_dff_A_HABd7t814_0),.din(w_dff_A_x9baV45f4_0),.clk(gclk));
	jdff dff_A_1r2cNNVA0_0(.dout(w_dff_A_x9baV45f4_0),.din(w_dff_A_1r2cNNVA0_0),.clk(gclk));
	jdff dff_A_vb3rHJys2_0(.dout(w_Gid0_0[0]),.din(w_dff_A_vb3rHJys2_0),.clk(gclk));
	jdff dff_A_pOuc5m0H8_0(.dout(w_dff_A_vb3rHJys2_0),.din(w_dff_A_pOuc5m0H8_0),.clk(gclk));
	jdff dff_A_CtZl4NmD8_0(.dout(w_dff_A_pOuc5m0H8_0),.din(w_dff_A_CtZl4NmD8_0),.clk(gclk));
	jdff dff_A_D6MRQnTe2_0(.dout(w_dff_A_CtZl4NmD8_0),.din(w_dff_A_D6MRQnTe2_0),.clk(gclk));
	jdff dff_A_6Tt91TuU1_0(.dout(w_dff_A_D6MRQnTe2_0),.din(w_dff_A_6Tt91TuU1_0),.clk(gclk));
	jdff dff_A_xqW3bDJy5_0(.dout(w_dff_A_6Tt91TuU1_0),.din(w_dff_A_xqW3bDJy5_0),.clk(gclk));
	jdff dff_A_KtOsEIdM1_0(.dout(w_dff_A_xqW3bDJy5_0),.din(w_dff_A_KtOsEIdM1_0),.clk(gclk));
	jdff dff_A_FcfR02qE9_0(.dout(w_dff_A_KtOsEIdM1_0),.din(w_dff_A_FcfR02qE9_0),.clk(gclk));
	jdff dff_A_uam4Mvpt2_0(.dout(w_dff_A_FcfR02qE9_0),.din(w_dff_A_uam4Mvpt2_0),.clk(gclk));
	jdff dff_A_SMk4Rzs98_0(.dout(w_dff_A_uam4Mvpt2_0),.din(w_dff_A_SMk4Rzs98_0),.clk(gclk));
	jdff dff_A_6p8rAL8X3_0(.dout(w_Gid12_0[0]),.din(w_dff_A_6p8rAL8X3_0),.clk(gclk));
	jdff dff_A_qBIYq7za9_0(.dout(w_dff_A_6p8rAL8X3_0),.din(w_dff_A_qBIYq7za9_0),.clk(gclk));
	jdff dff_A_8LMXLivq2_0(.dout(w_dff_A_qBIYq7za9_0),.din(w_dff_A_8LMXLivq2_0),.clk(gclk));
	jdff dff_A_BFZ4Gl6V7_0(.dout(w_dff_A_8LMXLivq2_0),.din(w_dff_A_BFZ4Gl6V7_0),.clk(gclk));
	jdff dff_A_RYeFefF50_0(.dout(w_dff_A_BFZ4Gl6V7_0),.din(w_dff_A_RYeFefF50_0),.clk(gclk));
	jdff dff_A_wtKv9GSC0_0(.dout(w_dff_A_RYeFefF50_0),.din(w_dff_A_wtKv9GSC0_0),.clk(gclk));
	jdff dff_A_XoTgZfTW8_0(.dout(w_dff_A_wtKv9GSC0_0),.din(w_dff_A_XoTgZfTW8_0),.clk(gclk));
	jdff dff_A_N1Saaqg35_0(.dout(w_dff_A_XoTgZfTW8_0),.din(w_dff_A_N1Saaqg35_0),.clk(gclk));
	jdff dff_A_gu1ax10V9_0(.dout(w_dff_A_N1Saaqg35_0),.din(w_dff_A_gu1ax10V9_0),.clk(gclk));
	jdff dff_A_9wkS9wKr2_0(.dout(w_dff_A_gu1ax10V9_0),.din(w_dff_A_9wkS9wKr2_0),.clk(gclk));
	jdff dff_A_ducNOe8L5_0(.dout(w_Gid8_0[0]),.din(w_dff_A_ducNOe8L5_0),.clk(gclk));
	jdff dff_A_7D9VR66J9_0(.dout(w_dff_A_ducNOe8L5_0),.din(w_dff_A_7D9VR66J9_0),.clk(gclk));
	jdff dff_A_8WQZR0Lo2_0(.dout(w_dff_A_7D9VR66J9_0),.din(w_dff_A_8WQZR0Lo2_0),.clk(gclk));
	jdff dff_A_hzTifEEj1_0(.dout(w_dff_A_8WQZR0Lo2_0),.din(w_dff_A_hzTifEEj1_0),.clk(gclk));
	jdff dff_A_kk0O9RQQ1_0(.dout(w_dff_A_hzTifEEj1_0),.din(w_dff_A_kk0O9RQQ1_0),.clk(gclk));
	jdff dff_A_IiNwgC7z6_0(.dout(w_dff_A_kk0O9RQQ1_0),.din(w_dff_A_IiNwgC7z6_0),.clk(gclk));
	jdff dff_A_ayfZBSiF5_0(.dout(w_dff_A_IiNwgC7z6_0),.din(w_dff_A_ayfZBSiF5_0),.clk(gclk));
	jdff dff_A_zCH76v066_0(.dout(w_dff_A_ayfZBSiF5_0),.din(w_dff_A_zCH76v066_0),.clk(gclk));
	jdff dff_A_skjfGmJy5_0(.dout(w_dff_A_zCH76v066_0),.din(w_dff_A_skjfGmJy5_0),.clk(gclk));
	jdff dff_A_lLJru4AI4_0(.dout(w_dff_A_skjfGmJy5_0),.din(w_dff_A_lLJru4AI4_0),.clk(gclk));
	jdff dff_B_i2QgCSY68_2(.din(n242),.dout(w_dff_B_i2QgCSY68_2),.clk(gclk));
	jdff dff_B_nLoB99Yf0_2(.din(w_dff_B_i2QgCSY68_2),.dout(w_dff_B_nLoB99Yf0_2),.clk(gclk));
	jdff dff_B_5jl0f5es0_2(.din(w_dff_B_nLoB99Yf0_2),.dout(w_dff_B_5jl0f5es0_2),.clk(gclk));
	jdff dff_B_d6TFRYE03_2(.din(w_dff_B_5jl0f5es0_2),.dout(w_dff_B_d6TFRYE03_2),.clk(gclk));
	jdff dff_A_UgUr8UBQ2_0(.dout(w_Gid6_0[0]),.din(w_dff_A_UgUr8UBQ2_0),.clk(gclk));
	jdff dff_A_9vHPGOCY0_0(.dout(w_dff_A_UgUr8UBQ2_0),.din(w_dff_A_9vHPGOCY0_0),.clk(gclk));
	jdff dff_A_TVdCrnvH6_0(.dout(w_dff_A_9vHPGOCY0_0),.din(w_dff_A_TVdCrnvH6_0),.clk(gclk));
	jdff dff_A_mLuBbqSX2_0(.dout(w_dff_A_TVdCrnvH6_0),.din(w_dff_A_mLuBbqSX2_0),.clk(gclk));
	jdff dff_A_6RpvnYwd5_0(.dout(w_dff_A_mLuBbqSX2_0),.din(w_dff_A_6RpvnYwd5_0),.clk(gclk));
	jdff dff_A_8GFgmSi75_0(.dout(w_dff_A_6RpvnYwd5_0),.din(w_dff_A_8GFgmSi75_0),.clk(gclk));
	jdff dff_A_uAOKY6xX6_0(.dout(w_dff_A_8GFgmSi75_0),.din(w_dff_A_uAOKY6xX6_0),.clk(gclk));
	jdff dff_A_tVccIOZq0_0(.dout(w_dff_A_uAOKY6xX6_0),.din(w_dff_A_tVccIOZq0_0),.clk(gclk));
	jdff dff_A_i68Mpp0q3_0(.dout(w_dff_A_tVccIOZq0_0),.din(w_dff_A_i68Mpp0q3_0),.clk(gclk));
	jdff dff_A_5pI5wIum6_0(.dout(w_dff_A_i68Mpp0q3_0),.din(w_dff_A_5pI5wIum6_0),.clk(gclk));
	jdff dff_A_fhfL7ZNh2_0(.dout(w_Gid2_0[0]),.din(w_dff_A_fhfL7ZNh2_0),.clk(gclk));
	jdff dff_A_QtYcn6H17_0(.dout(w_dff_A_fhfL7ZNh2_0),.din(w_dff_A_QtYcn6H17_0),.clk(gclk));
	jdff dff_A_N5MTlNjS2_0(.dout(w_dff_A_QtYcn6H17_0),.din(w_dff_A_N5MTlNjS2_0),.clk(gclk));
	jdff dff_A_j8fZ2d6n1_0(.dout(w_dff_A_N5MTlNjS2_0),.din(w_dff_A_j8fZ2d6n1_0),.clk(gclk));
	jdff dff_A_8RceGFPk9_0(.dout(w_dff_A_j8fZ2d6n1_0),.din(w_dff_A_8RceGFPk9_0),.clk(gclk));
	jdff dff_A_Azv9j80w7_0(.dout(w_dff_A_8RceGFPk9_0),.din(w_dff_A_Azv9j80w7_0),.clk(gclk));
	jdff dff_A_ws4PACSk6_0(.dout(w_dff_A_Azv9j80w7_0),.din(w_dff_A_ws4PACSk6_0),.clk(gclk));
	jdff dff_A_5PSOEEr27_0(.dout(w_dff_A_ws4PACSk6_0),.din(w_dff_A_5PSOEEr27_0),.clk(gclk));
	jdff dff_A_g93EImtD5_0(.dout(w_dff_A_5PSOEEr27_0),.din(w_dff_A_g93EImtD5_0),.clk(gclk));
	jdff dff_A_0SJj0lBu8_0(.dout(w_dff_A_g93EImtD5_0),.din(w_dff_A_0SJj0lBu8_0),.clk(gclk));
	jdff dff_A_HNuj0yP36_0(.dout(w_Gid14_0[0]),.din(w_dff_A_HNuj0yP36_0),.clk(gclk));
	jdff dff_A_zJqql4ae2_0(.dout(w_dff_A_HNuj0yP36_0),.din(w_dff_A_zJqql4ae2_0),.clk(gclk));
	jdff dff_A_oon9BExA8_0(.dout(w_dff_A_zJqql4ae2_0),.din(w_dff_A_oon9BExA8_0),.clk(gclk));
	jdff dff_A_kABiU4ks4_0(.dout(w_dff_A_oon9BExA8_0),.din(w_dff_A_kABiU4ks4_0),.clk(gclk));
	jdff dff_A_qzAnkGuX6_0(.dout(w_dff_A_kABiU4ks4_0),.din(w_dff_A_qzAnkGuX6_0),.clk(gclk));
	jdff dff_A_t9UoYn2L6_0(.dout(w_dff_A_qzAnkGuX6_0),.din(w_dff_A_t9UoYn2L6_0),.clk(gclk));
	jdff dff_A_yLqZb8ab4_0(.dout(w_dff_A_t9UoYn2L6_0),.din(w_dff_A_yLqZb8ab4_0),.clk(gclk));
	jdff dff_A_f1RmbKaB7_0(.dout(w_dff_A_yLqZb8ab4_0),.din(w_dff_A_f1RmbKaB7_0),.clk(gclk));
	jdff dff_A_fJL16Qb31_0(.dout(w_dff_A_f1RmbKaB7_0),.din(w_dff_A_fJL16Qb31_0),.clk(gclk));
	jdff dff_A_LyMrNUTW1_0(.dout(w_dff_A_fJL16Qb31_0),.din(w_dff_A_LyMrNUTW1_0),.clk(gclk));
	jdff dff_A_Rn5TqlOD3_0(.dout(w_Gid10_0[0]),.din(w_dff_A_Rn5TqlOD3_0),.clk(gclk));
	jdff dff_A_UWXZGQUD1_0(.dout(w_dff_A_Rn5TqlOD3_0),.din(w_dff_A_UWXZGQUD1_0),.clk(gclk));
	jdff dff_A_KtrV4DP85_0(.dout(w_dff_A_UWXZGQUD1_0),.din(w_dff_A_KtrV4DP85_0),.clk(gclk));
	jdff dff_A_tRHN7J6B8_0(.dout(w_dff_A_KtrV4DP85_0),.din(w_dff_A_tRHN7J6B8_0),.clk(gclk));
	jdff dff_A_EiyU3HGR1_0(.dout(w_dff_A_tRHN7J6B8_0),.din(w_dff_A_EiyU3HGR1_0),.clk(gclk));
	jdff dff_A_EWmpaWPZ1_0(.dout(w_dff_A_EiyU3HGR1_0),.din(w_dff_A_EWmpaWPZ1_0),.clk(gclk));
	jdff dff_A_CNgnRqxO1_0(.dout(w_dff_A_EWmpaWPZ1_0),.din(w_dff_A_CNgnRqxO1_0),.clk(gclk));
	jdff dff_A_UOdM8lSR2_0(.dout(w_dff_A_CNgnRqxO1_0),.din(w_dff_A_UOdM8lSR2_0),.clk(gclk));
	jdff dff_A_rOeqALvP1_0(.dout(w_dff_A_UOdM8lSR2_0),.din(w_dff_A_rOeqALvP1_0),.clk(gclk));
	jdff dff_A_wYS3BdfW6_0(.dout(w_dff_A_rOeqALvP1_0),.din(w_dff_A_wYS3BdfW6_0),.clk(gclk));
	jdff dff_A_qFWcYLoC7_0(.dout(w_Gid17_0[0]),.din(w_dff_A_qFWcYLoC7_0),.clk(gclk));
	jdff dff_A_JmEtiWwd6_0(.dout(w_dff_A_qFWcYLoC7_0),.din(w_dff_A_JmEtiWwd6_0),.clk(gclk));
	jdff dff_A_GmVmhRdX0_0(.dout(w_dff_A_JmEtiWwd6_0),.din(w_dff_A_GmVmhRdX0_0),.clk(gclk));
	jdff dff_A_WJUEV0YA2_0(.dout(w_dff_A_GmVmhRdX0_0),.din(w_dff_A_WJUEV0YA2_0),.clk(gclk));
	jdff dff_A_maGIHF550_0(.dout(w_dff_A_WJUEV0YA2_0),.din(w_dff_A_maGIHF550_0),.clk(gclk));
	jdff dff_A_rBrydVzj8_0(.dout(w_dff_A_maGIHF550_0),.din(w_dff_A_rBrydVzj8_0),.clk(gclk));
	jdff dff_A_Yi4eIttP4_0(.dout(w_dff_A_rBrydVzj8_0),.din(w_dff_A_Yi4eIttP4_0),.clk(gclk));
	jdff dff_A_Ab6nBgXj9_0(.dout(w_dff_A_Yi4eIttP4_0),.din(w_dff_A_Ab6nBgXj9_0),.clk(gclk));
	jdff dff_A_Z9o0sFDI8_0(.dout(w_dff_A_Ab6nBgXj9_0),.din(w_dff_A_Z9o0sFDI8_0),.clk(gclk));
	jdff dff_A_GZgjHeOx8_0(.dout(w_dff_A_Z9o0sFDI8_0),.din(w_dff_A_GZgjHeOx8_0),.clk(gclk));
	jdff dff_A_kZnL2V1h6_0(.dout(w_dff_A_GZgjHeOx8_0),.din(w_dff_A_kZnL2V1h6_0),.clk(gclk));
	jdff dff_A_lGMmi9g90_0(.dout(w_Gid16_0[0]),.din(w_dff_A_lGMmi9g90_0),.clk(gclk));
	jdff dff_A_BAqnZPKJ8_0(.dout(w_dff_A_lGMmi9g90_0),.din(w_dff_A_BAqnZPKJ8_0),.clk(gclk));
	jdff dff_A_vJQWoq4r7_0(.dout(w_dff_A_BAqnZPKJ8_0),.din(w_dff_A_vJQWoq4r7_0),.clk(gclk));
	jdff dff_A_hQvNw3Qa3_0(.dout(w_dff_A_vJQWoq4r7_0),.din(w_dff_A_hQvNw3Qa3_0),.clk(gclk));
	jdff dff_A_fsyqxTHM3_0(.dout(w_dff_A_hQvNw3Qa3_0),.din(w_dff_A_fsyqxTHM3_0),.clk(gclk));
	jdff dff_A_PH0OJDwd1_0(.dout(w_dff_A_fsyqxTHM3_0),.din(w_dff_A_PH0OJDwd1_0),.clk(gclk));
	jdff dff_A_k7y2Wtrb7_0(.dout(w_dff_A_PH0OJDwd1_0),.din(w_dff_A_k7y2Wtrb7_0),.clk(gclk));
	jdff dff_A_nnFGBZ531_0(.dout(w_dff_A_k7y2Wtrb7_0),.din(w_dff_A_nnFGBZ531_0),.clk(gclk));
	jdff dff_A_R9sJ7BM73_0(.dout(w_dff_A_nnFGBZ531_0),.din(w_dff_A_R9sJ7BM73_0),.clk(gclk));
	jdff dff_A_nqcVuyQD6_0(.dout(w_dff_A_R9sJ7BM73_0),.din(w_dff_A_nqcVuyQD6_0),.clk(gclk));
	jdff dff_A_DJEzk7og9_0(.dout(w_dff_A_nqcVuyQD6_0),.din(w_dff_A_DJEzk7og9_0),.clk(gclk));
	jdff dff_A_F8Vfn9dx4_0(.dout(w_Gid19_0[0]),.din(w_dff_A_F8Vfn9dx4_0),.clk(gclk));
	jdff dff_A_WKlTuUQc7_0(.dout(w_dff_A_F8Vfn9dx4_0),.din(w_dff_A_WKlTuUQc7_0),.clk(gclk));
	jdff dff_A_QMdbRlZh5_0(.dout(w_dff_A_WKlTuUQc7_0),.din(w_dff_A_QMdbRlZh5_0),.clk(gclk));
	jdff dff_A_drsbM2rL6_0(.dout(w_dff_A_QMdbRlZh5_0),.din(w_dff_A_drsbM2rL6_0),.clk(gclk));
	jdff dff_A_APMNqhGG7_0(.dout(w_dff_A_drsbM2rL6_0),.din(w_dff_A_APMNqhGG7_0),.clk(gclk));
	jdff dff_A_UJlRumnJ0_0(.dout(w_dff_A_APMNqhGG7_0),.din(w_dff_A_UJlRumnJ0_0),.clk(gclk));
	jdff dff_A_X69MC0nZ4_0(.dout(w_dff_A_UJlRumnJ0_0),.din(w_dff_A_X69MC0nZ4_0),.clk(gclk));
	jdff dff_A_Zu7sxXR45_0(.dout(w_dff_A_X69MC0nZ4_0),.din(w_dff_A_Zu7sxXR45_0),.clk(gclk));
	jdff dff_A_7xihvIPF0_0(.dout(w_dff_A_Zu7sxXR45_0),.din(w_dff_A_7xihvIPF0_0),.clk(gclk));
	jdff dff_A_ALfTx6m19_0(.dout(w_dff_A_7xihvIPF0_0),.din(w_dff_A_ALfTx6m19_0),.clk(gclk));
	jdff dff_A_culgjWxi5_0(.dout(w_dff_A_ALfTx6m19_0),.din(w_dff_A_culgjWxi5_0),.clk(gclk));
	jdff dff_A_Pr0Wo26f8_0(.dout(w_Gid18_0[0]),.din(w_dff_A_Pr0Wo26f8_0),.clk(gclk));
	jdff dff_A_BCldgjlb5_0(.dout(w_dff_A_Pr0Wo26f8_0),.din(w_dff_A_BCldgjlb5_0),.clk(gclk));
	jdff dff_A_zFSxSAr91_0(.dout(w_dff_A_BCldgjlb5_0),.din(w_dff_A_zFSxSAr91_0),.clk(gclk));
	jdff dff_A_qOe9KJQn9_0(.dout(w_dff_A_zFSxSAr91_0),.din(w_dff_A_qOe9KJQn9_0),.clk(gclk));
	jdff dff_A_mlIfPHH50_0(.dout(w_dff_A_qOe9KJQn9_0),.din(w_dff_A_mlIfPHH50_0),.clk(gclk));
	jdff dff_A_gEQ2B0xt9_0(.dout(w_dff_A_mlIfPHH50_0),.din(w_dff_A_gEQ2B0xt9_0),.clk(gclk));
	jdff dff_A_vWwtNhQM4_0(.dout(w_dff_A_gEQ2B0xt9_0),.din(w_dff_A_vWwtNhQM4_0),.clk(gclk));
	jdff dff_A_qWKTROdI5_0(.dout(w_dff_A_vWwtNhQM4_0),.din(w_dff_A_qWKTROdI5_0),.clk(gclk));
	jdff dff_A_eu05rmxx8_0(.dout(w_dff_A_qWKTROdI5_0),.din(w_dff_A_eu05rmxx8_0),.clk(gclk));
	jdff dff_A_T2YkXJPR8_0(.dout(w_dff_A_eu05rmxx8_0),.din(w_dff_A_T2YkXJPR8_0),.clk(gclk));
	jdff dff_A_VQhWYieE2_0(.dout(w_dff_A_T2YkXJPR8_0),.din(w_dff_A_VQhWYieE2_0),.clk(gclk));
	jdff dff_A_9ma5OEpZ6_0(.dout(w_n136_0[0]),.din(w_dff_A_9ma5OEpZ6_0),.clk(gclk));
	jdff dff_A_8BagOsUg4_0(.dout(w_Gid25_0[0]),.din(w_dff_A_8BagOsUg4_0),.clk(gclk));
	jdff dff_A_HMtBuOwS0_0(.dout(w_dff_A_8BagOsUg4_0),.din(w_dff_A_HMtBuOwS0_0),.clk(gclk));
	jdff dff_A_3k77Rm1d7_0(.dout(w_dff_A_HMtBuOwS0_0),.din(w_dff_A_3k77Rm1d7_0),.clk(gclk));
	jdff dff_A_Rt1Zs4yD5_0(.dout(w_dff_A_3k77Rm1d7_0),.din(w_dff_A_Rt1Zs4yD5_0),.clk(gclk));
	jdff dff_A_R6hLT1gF6_0(.dout(w_dff_A_Rt1Zs4yD5_0),.din(w_dff_A_R6hLT1gF6_0),.clk(gclk));
	jdff dff_A_Ee2OX39E3_0(.dout(w_dff_A_R6hLT1gF6_0),.din(w_dff_A_Ee2OX39E3_0),.clk(gclk));
	jdff dff_A_pMjxcQUz9_0(.dout(w_dff_A_Ee2OX39E3_0),.din(w_dff_A_pMjxcQUz9_0),.clk(gclk));
	jdff dff_A_JH6rEZM93_0(.dout(w_dff_A_pMjxcQUz9_0),.din(w_dff_A_JH6rEZM93_0),.clk(gclk));
	jdff dff_A_Ccze5qj86_0(.dout(w_dff_A_JH6rEZM93_0),.din(w_dff_A_Ccze5qj86_0),.clk(gclk));
	jdff dff_A_LX3bRr914_0(.dout(w_dff_A_Ccze5qj86_0),.din(w_dff_A_LX3bRr914_0),.clk(gclk));
	jdff dff_A_I8rUbnB55_0(.dout(w_dff_A_LX3bRr914_0),.din(w_dff_A_I8rUbnB55_0),.clk(gclk));
	jdff dff_A_hJqy3NvD0_0(.dout(w_Gid24_0[0]),.din(w_dff_A_hJqy3NvD0_0),.clk(gclk));
	jdff dff_A_LmhYSz0f9_0(.dout(w_dff_A_hJqy3NvD0_0),.din(w_dff_A_LmhYSz0f9_0),.clk(gclk));
	jdff dff_A_8M1roRHN0_0(.dout(w_dff_A_LmhYSz0f9_0),.din(w_dff_A_8M1roRHN0_0),.clk(gclk));
	jdff dff_A_ER1JIcbh4_0(.dout(w_dff_A_8M1roRHN0_0),.din(w_dff_A_ER1JIcbh4_0),.clk(gclk));
	jdff dff_A_zEsPKpjQ5_0(.dout(w_dff_A_ER1JIcbh4_0),.din(w_dff_A_zEsPKpjQ5_0),.clk(gclk));
	jdff dff_A_XhjLBntL7_0(.dout(w_dff_A_zEsPKpjQ5_0),.din(w_dff_A_XhjLBntL7_0),.clk(gclk));
	jdff dff_A_mL1eZsne1_0(.dout(w_dff_A_XhjLBntL7_0),.din(w_dff_A_mL1eZsne1_0),.clk(gclk));
	jdff dff_A_vA3dOAXc9_0(.dout(w_dff_A_mL1eZsne1_0),.din(w_dff_A_vA3dOAXc9_0),.clk(gclk));
	jdff dff_A_kbDH5LK66_0(.dout(w_dff_A_vA3dOAXc9_0),.din(w_dff_A_kbDH5LK66_0),.clk(gclk));
	jdff dff_A_1uTknrlB2_0(.dout(w_dff_A_kbDH5LK66_0),.din(w_dff_A_1uTknrlB2_0),.clk(gclk));
	jdff dff_A_JDtv5Dbc7_0(.dout(w_dff_A_1uTknrlB2_0),.din(w_dff_A_JDtv5Dbc7_0),.clk(gclk));
	jdff dff_A_hAJX8MYo6_0(.dout(w_Gid27_0[0]),.din(w_dff_A_hAJX8MYo6_0),.clk(gclk));
	jdff dff_A_SkR9i0C66_0(.dout(w_dff_A_hAJX8MYo6_0),.din(w_dff_A_SkR9i0C66_0),.clk(gclk));
	jdff dff_A_nLTRSfP39_0(.dout(w_dff_A_SkR9i0C66_0),.din(w_dff_A_nLTRSfP39_0),.clk(gclk));
	jdff dff_A_IZAKN65i9_0(.dout(w_dff_A_nLTRSfP39_0),.din(w_dff_A_IZAKN65i9_0),.clk(gclk));
	jdff dff_A_fU09Vo9m5_0(.dout(w_dff_A_IZAKN65i9_0),.din(w_dff_A_fU09Vo9m5_0),.clk(gclk));
	jdff dff_A_IKH5coRy4_0(.dout(w_dff_A_fU09Vo9m5_0),.din(w_dff_A_IKH5coRy4_0),.clk(gclk));
	jdff dff_A_mNK3ulU47_0(.dout(w_dff_A_IKH5coRy4_0),.din(w_dff_A_mNK3ulU47_0),.clk(gclk));
	jdff dff_A_c2ZlCHke9_0(.dout(w_dff_A_mNK3ulU47_0),.din(w_dff_A_c2ZlCHke9_0),.clk(gclk));
	jdff dff_A_AXj4PQA77_0(.dout(w_dff_A_c2ZlCHke9_0),.din(w_dff_A_AXj4PQA77_0),.clk(gclk));
	jdff dff_A_bDJzTEBM7_0(.dout(w_dff_A_AXj4PQA77_0),.din(w_dff_A_bDJzTEBM7_0),.clk(gclk));
	jdff dff_A_VCEw40Ni6_0(.dout(w_dff_A_bDJzTEBM7_0),.din(w_dff_A_VCEw40Ni6_0),.clk(gclk));
	jdff dff_A_4XYts8Ih4_0(.dout(w_Gid26_0[0]),.din(w_dff_A_4XYts8Ih4_0),.clk(gclk));
	jdff dff_A_OiQ4UZXn2_0(.dout(w_dff_A_4XYts8Ih4_0),.din(w_dff_A_OiQ4UZXn2_0),.clk(gclk));
	jdff dff_A_GEQXTNG92_0(.dout(w_dff_A_OiQ4UZXn2_0),.din(w_dff_A_GEQXTNG92_0),.clk(gclk));
	jdff dff_A_TrJ5Ua3e6_0(.dout(w_dff_A_GEQXTNG92_0),.din(w_dff_A_TrJ5Ua3e6_0),.clk(gclk));
	jdff dff_A_gi3HS6BD6_0(.dout(w_dff_A_TrJ5Ua3e6_0),.din(w_dff_A_gi3HS6BD6_0),.clk(gclk));
	jdff dff_A_i8cqEZ3d1_0(.dout(w_dff_A_gi3HS6BD6_0),.din(w_dff_A_i8cqEZ3d1_0),.clk(gclk));
	jdff dff_A_y7p6YtTU9_0(.dout(w_dff_A_i8cqEZ3d1_0),.din(w_dff_A_y7p6YtTU9_0),.clk(gclk));
	jdff dff_A_Gbttuphg8_0(.dout(w_dff_A_y7p6YtTU9_0),.din(w_dff_A_Gbttuphg8_0),.clk(gclk));
	jdff dff_A_Da0CxEfd3_0(.dout(w_dff_A_Gbttuphg8_0),.din(w_dff_A_Da0CxEfd3_0),.clk(gclk));
	jdff dff_A_KCBCdx4k0_0(.dout(w_dff_A_Da0CxEfd3_0),.din(w_dff_A_KCBCdx4k0_0),.clk(gclk));
	jdff dff_A_TQHmocMZ4_0(.dout(w_dff_A_KCBCdx4k0_0),.din(w_dff_A_TQHmocMZ4_0),.clk(gclk));
	jdff dff_A_BNTmMqoF1_0(.dout(w_n147_0[0]),.din(w_dff_A_BNTmMqoF1_0),.clk(gclk));
	jdff dff_A_54N0ugNR8_0(.dout(w_dff_A_BNTmMqoF1_0),.din(w_dff_A_54N0ugNR8_0),.clk(gclk));
	jdff dff_A_YiYD7WbE9_0(.dout(w_dff_A_54N0ugNR8_0),.din(w_dff_A_YiYD7WbE9_0),.clk(gclk));
	jdff dff_A_NkiZxHnA9_0(.dout(w_dff_A_YiYD7WbE9_0),.din(w_dff_A_NkiZxHnA9_0),.clk(gclk));
	jdff dff_A_UsLC33ks8_0(.dout(w_dff_A_NkiZxHnA9_0),.din(w_dff_A_UsLC33ks8_0),.clk(gclk));
	jdff dff_A_XXhkhR7c0_0(.dout(w_Gid7_0[0]),.din(w_dff_A_XXhkhR7c0_0),.clk(gclk));
	jdff dff_A_7qIiETBN5_0(.dout(w_dff_A_XXhkhR7c0_0),.din(w_dff_A_7qIiETBN5_0),.clk(gclk));
	jdff dff_A_yCSWFzxC4_0(.dout(w_dff_A_7qIiETBN5_0),.din(w_dff_A_yCSWFzxC4_0),.clk(gclk));
	jdff dff_A_z0xVy3rQ8_0(.dout(w_dff_A_yCSWFzxC4_0),.din(w_dff_A_z0xVy3rQ8_0),.clk(gclk));
	jdff dff_A_Fl31Y6cF4_0(.dout(w_dff_A_z0xVy3rQ8_0),.din(w_dff_A_Fl31Y6cF4_0),.clk(gclk));
	jdff dff_A_XBN8ZKPt8_0(.dout(w_dff_A_Fl31Y6cF4_0),.din(w_dff_A_XBN8ZKPt8_0),.clk(gclk));
	jdff dff_A_hZtC0qdE5_0(.dout(w_dff_A_XBN8ZKPt8_0),.din(w_dff_A_hZtC0qdE5_0),.clk(gclk));
	jdff dff_A_qTZFW09T6_0(.dout(w_dff_A_hZtC0qdE5_0),.din(w_dff_A_qTZFW09T6_0),.clk(gclk));
	jdff dff_A_WYgKLuSK9_0(.dout(w_dff_A_qTZFW09T6_0),.din(w_dff_A_WYgKLuSK9_0),.clk(gclk));
	jdff dff_A_ipJAZuyO5_0(.dout(w_dff_A_WYgKLuSK9_0),.din(w_dff_A_ipJAZuyO5_0),.clk(gclk));
	jdff dff_A_Shhlcgov3_0(.dout(w_Gid3_0[0]),.din(w_dff_A_Shhlcgov3_0),.clk(gclk));
	jdff dff_A_8BknCDYj9_0(.dout(w_dff_A_Shhlcgov3_0),.din(w_dff_A_8BknCDYj9_0),.clk(gclk));
	jdff dff_A_bfr27rka7_0(.dout(w_dff_A_8BknCDYj9_0),.din(w_dff_A_bfr27rka7_0),.clk(gclk));
	jdff dff_A_t2CEq2bh9_0(.dout(w_dff_A_bfr27rka7_0),.din(w_dff_A_t2CEq2bh9_0),.clk(gclk));
	jdff dff_A_xqUB5j9J1_0(.dout(w_dff_A_t2CEq2bh9_0),.din(w_dff_A_xqUB5j9J1_0),.clk(gclk));
	jdff dff_A_60zMKwgT3_0(.dout(w_dff_A_xqUB5j9J1_0),.din(w_dff_A_60zMKwgT3_0),.clk(gclk));
	jdff dff_A_FYOqB6Jq1_0(.dout(w_dff_A_60zMKwgT3_0),.din(w_dff_A_FYOqB6Jq1_0),.clk(gclk));
	jdff dff_A_PuMsEJvb8_0(.dout(w_dff_A_FYOqB6Jq1_0),.din(w_dff_A_PuMsEJvb8_0),.clk(gclk));
	jdff dff_A_vupwB64w1_0(.dout(w_dff_A_PuMsEJvb8_0),.din(w_dff_A_vupwB64w1_0),.clk(gclk));
	jdff dff_A_vn5rWJvX4_0(.dout(w_dff_A_vupwB64w1_0),.din(w_dff_A_vn5rWJvX4_0),.clk(gclk));
	jdff dff_A_L7uZj2Jn7_0(.dout(w_Gid15_0[0]),.din(w_dff_A_L7uZj2Jn7_0),.clk(gclk));
	jdff dff_A_lG6GjrXS9_0(.dout(w_dff_A_L7uZj2Jn7_0),.din(w_dff_A_lG6GjrXS9_0),.clk(gclk));
	jdff dff_A_7gIX5W2F1_0(.dout(w_dff_A_lG6GjrXS9_0),.din(w_dff_A_7gIX5W2F1_0),.clk(gclk));
	jdff dff_A_40U1t4ak5_0(.dout(w_dff_A_7gIX5W2F1_0),.din(w_dff_A_40U1t4ak5_0),.clk(gclk));
	jdff dff_A_yaObO7Ng2_0(.dout(w_dff_A_40U1t4ak5_0),.din(w_dff_A_yaObO7Ng2_0),.clk(gclk));
	jdff dff_A_D0kKTEau4_0(.dout(w_dff_A_yaObO7Ng2_0),.din(w_dff_A_D0kKTEau4_0),.clk(gclk));
	jdff dff_A_gQzXy2BT0_0(.dout(w_dff_A_D0kKTEau4_0),.din(w_dff_A_gQzXy2BT0_0),.clk(gclk));
	jdff dff_A_JuY88UlQ3_0(.dout(w_dff_A_gQzXy2BT0_0),.din(w_dff_A_JuY88UlQ3_0),.clk(gclk));
	jdff dff_A_e7s5LfX73_0(.dout(w_dff_A_JuY88UlQ3_0),.din(w_dff_A_e7s5LfX73_0),.clk(gclk));
	jdff dff_A_9kS1c7it8_0(.dout(w_dff_A_e7s5LfX73_0),.din(w_dff_A_9kS1c7it8_0),.clk(gclk));
	jdff dff_A_E4hNQIqu8_0(.dout(w_Gid11_0[0]),.din(w_dff_A_E4hNQIqu8_0),.clk(gclk));
	jdff dff_A_QPhhcsxM2_0(.dout(w_dff_A_E4hNQIqu8_0),.din(w_dff_A_QPhhcsxM2_0),.clk(gclk));
	jdff dff_A_CBl3IIGX8_0(.dout(w_dff_A_QPhhcsxM2_0),.din(w_dff_A_CBl3IIGX8_0),.clk(gclk));
	jdff dff_A_pBg22DGl9_0(.dout(w_dff_A_CBl3IIGX8_0),.din(w_dff_A_pBg22DGl9_0),.clk(gclk));
	jdff dff_A_xmyBsTe45_0(.dout(w_dff_A_pBg22DGl9_0),.din(w_dff_A_xmyBsTe45_0),.clk(gclk));
	jdff dff_A_T4A39mOC7_0(.dout(w_dff_A_xmyBsTe45_0),.din(w_dff_A_T4A39mOC7_0),.clk(gclk));
	jdff dff_A_ySQpeBkw8_0(.dout(w_dff_A_T4A39mOC7_0),.din(w_dff_A_ySQpeBkw8_0),.clk(gclk));
	jdff dff_A_xEK5MWRf0_0(.dout(w_dff_A_ySQpeBkw8_0),.din(w_dff_A_xEK5MWRf0_0),.clk(gclk));
	jdff dff_A_xbrBFJZR3_0(.dout(w_dff_A_xEK5MWRf0_0),.din(w_dff_A_xbrBFJZR3_0),.clk(gclk));
	jdff dff_A_DnccThX34_0(.dout(w_dff_A_xbrBFJZR3_0),.din(w_dff_A_DnccThX34_0),.clk(gclk));
	jdff dff_A_Rp9G3c4u3_0(.dout(w_Gid21_0[0]),.din(w_dff_A_Rp9G3c4u3_0),.clk(gclk));
	jdff dff_A_EBBf7ufV7_0(.dout(w_dff_A_Rp9G3c4u3_0),.din(w_dff_A_EBBf7ufV7_0),.clk(gclk));
	jdff dff_A_mTG1dvKJ5_0(.dout(w_dff_A_EBBf7ufV7_0),.din(w_dff_A_mTG1dvKJ5_0),.clk(gclk));
	jdff dff_A_wVx6AIv85_0(.dout(w_dff_A_mTG1dvKJ5_0),.din(w_dff_A_wVx6AIv85_0),.clk(gclk));
	jdff dff_A_FK2uUZDw2_0(.dout(w_dff_A_wVx6AIv85_0),.din(w_dff_A_FK2uUZDw2_0),.clk(gclk));
	jdff dff_A_X95GqGPh5_0(.dout(w_dff_A_FK2uUZDw2_0),.din(w_dff_A_X95GqGPh5_0),.clk(gclk));
	jdff dff_A_iNpbyG9T4_0(.dout(w_dff_A_X95GqGPh5_0),.din(w_dff_A_iNpbyG9T4_0),.clk(gclk));
	jdff dff_A_d1OKbcRq4_0(.dout(w_dff_A_iNpbyG9T4_0),.din(w_dff_A_d1OKbcRq4_0),.clk(gclk));
	jdff dff_A_E28qXkd37_0(.dout(w_dff_A_d1OKbcRq4_0),.din(w_dff_A_E28qXkd37_0),.clk(gclk));
	jdff dff_A_Ubj9B6lp2_0(.dout(w_dff_A_E28qXkd37_0),.din(w_dff_A_Ubj9B6lp2_0),.clk(gclk));
	jdff dff_A_OWywckru0_0(.dout(w_dff_A_Ubj9B6lp2_0),.din(w_dff_A_OWywckru0_0),.clk(gclk));
	jdff dff_A_X5Pwss0z4_0(.dout(w_Gid20_0[0]),.din(w_dff_A_X5Pwss0z4_0),.clk(gclk));
	jdff dff_A_lCN1uvi33_0(.dout(w_dff_A_X5Pwss0z4_0),.din(w_dff_A_lCN1uvi33_0),.clk(gclk));
	jdff dff_A_V5zIibt05_0(.dout(w_dff_A_lCN1uvi33_0),.din(w_dff_A_V5zIibt05_0),.clk(gclk));
	jdff dff_A_QhE8VnNu5_0(.dout(w_dff_A_V5zIibt05_0),.din(w_dff_A_QhE8VnNu5_0),.clk(gclk));
	jdff dff_A_QVH7nSfG6_0(.dout(w_dff_A_QhE8VnNu5_0),.din(w_dff_A_QVH7nSfG6_0),.clk(gclk));
	jdff dff_A_WGwoBsqf6_0(.dout(w_dff_A_QVH7nSfG6_0),.din(w_dff_A_WGwoBsqf6_0),.clk(gclk));
	jdff dff_A_m0p89FOw6_0(.dout(w_dff_A_WGwoBsqf6_0),.din(w_dff_A_m0p89FOw6_0),.clk(gclk));
	jdff dff_A_uUIN0ozZ2_0(.dout(w_dff_A_m0p89FOw6_0),.din(w_dff_A_uUIN0ozZ2_0),.clk(gclk));
	jdff dff_A_SdPtLtkQ1_0(.dout(w_dff_A_uUIN0ozZ2_0),.din(w_dff_A_SdPtLtkQ1_0),.clk(gclk));
	jdff dff_A_XW0H1AoH0_0(.dout(w_dff_A_SdPtLtkQ1_0),.din(w_dff_A_XW0H1AoH0_0),.clk(gclk));
	jdff dff_A_QMFA5xbD2_0(.dout(w_dff_A_XW0H1AoH0_0),.din(w_dff_A_QMFA5xbD2_0),.clk(gclk));
	jdff dff_A_ZZGI2iuE9_0(.dout(w_Gid23_0[0]),.din(w_dff_A_ZZGI2iuE9_0),.clk(gclk));
	jdff dff_A_xZ34f1IN0_0(.dout(w_dff_A_ZZGI2iuE9_0),.din(w_dff_A_xZ34f1IN0_0),.clk(gclk));
	jdff dff_A_WvYyWxzg7_0(.dout(w_dff_A_xZ34f1IN0_0),.din(w_dff_A_WvYyWxzg7_0),.clk(gclk));
	jdff dff_A_m0X0DNV68_0(.dout(w_dff_A_WvYyWxzg7_0),.din(w_dff_A_m0X0DNV68_0),.clk(gclk));
	jdff dff_A_BJiU8Dli1_0(.dout(w_dff_A_m0X0DNV68_0),.din(w_dff_A_BJiU8Dli1_0),.clk(gclk));
	jdff dff_A_HgPP4Jc56_0(.dout(w_dff_A_BJiU8Dli1_0),.din(w_dff_A_HgPP4Jc56_0),.clk(gclk));
	jdff dff_A_NxDc3Nsk1_0(.dout(w_dff_A_HgPP4Jc56_0),.din(w_dff_A_NxDc3Nsk1_0),.clk(gclk));
	jdff dff_A_oIdN7jbs0_0(.dout(w_dff_A_NxDc3Nsk1_0),.din(w_dff_A_oIdN7jbs0_0),.clk(gclk));
	jdff dff_A_kXAsLSNA0_0(.dout(w_dff_A_oIdN7jbs0_0),.din(w_dff_A_kXAsLSNA0_0),.clk(gclk));
	jdff dff_A_44Qqi6fu9_0(.dout(w_dff_A_kXAsLSNA0_0),.din(w_dff_A_44Qqi6fu9_0),.clk(gclk));
	jdff dff_A_MdgH81Vo4_0(.dout(w_dff_A_44Qqi6fu9_0),.din(w_dff_A_MdgH81Vo4_0),.clk(gclk));
	jdff dff_A_TUXxjpHt8_0(.dout(w_Gid22_0[0]),.din(w_dff_A_TUXxjpHt8_0),.clk(gclk));
	jdff dff_A_T3JgPuRN1_0(.dout(w_dff_A_TUXxjpHt8_0),.din(w_dff_A_T3JgPuRN1_0),.clk(gclk));
	jdff dff_A_6Ut0vQrG8_0(.dout(w_dff_A_T3JgPuRN1_0),.din(w_dff_A_6Ut0vQrG8_0),.clk(gclk));
	jdff dff_A_kpB5NQOi3_0(.dout(w_dff_A_6Ut0vQrG8_0),.din(w_dff_A_kpB5NQOi3_0),.clk(gclk));
	jdff dff_A_KB8rMTdo9_0(.dout(w_dff_A_kpB5NQOi3_0),.din(w_dff_A_KB8rMTdo9_0),.clk(gclk));
	jdff dff_A_npAutbBS9_0(.dout(w_dff_A_KB8rMTdo9_0),.din(w_dff_A_npAutbBS9_0),.clk(gclk));
	jdff dff_A_TA17G0Iy6_0(.dout(w_dff_A_npAutbBS9_0),.din(w_dff_A_TA17G0Iy6_0),.clk(gclk));
	jdff dff_A_1NjX9CGf4_0(.dout(w_dff_A_TA17G0Iy6_0),.din(w_dff_A_1NjX9CGf4_0),.clk(gclk));
	jdff dff_A_rEfNOk1Z8_0(.dout(w_dff_A_1NjX9CGf4_0),.din(w_dff_A_rEfNOk1Z8_0),.clk(gclk));
	jdff dff_A_Wfivb2Fg1_0(.dout(w_dff_A_rEfNOk1Z8_0),.din(w_dff_A_Wfivb2Fg1_0),.clk(gclk));
	jdff dff_A_dDbXMIj37_0(.dout(w_dff_A_Wfivb2Fg1_0),.din(w_dff_A_dDbXMIj37_0),.clk(gclk));
	jdff dff_A_ieHKHVNB2_0(.dout(w_n128_0[0]),.din(w_dff_A_ieHKHVNB2_0),.clk(gclk));
	jdff dff_A_I3AI6Ynl2_0(.dout(w_Gid29_0[0]),.din(w_dff_A_I3AI6Ynl2_0),.clk(gclk));
	jdff dff_A_1NfHusSD0_0(.dout(w_dff_A_I3AI6Ynl2_0),.din(w_dff_A_1NfHusSD0_0),.clk(gclk));
	jdff dff_A_GXEKt2T89_0(.dout(w_dff_A_1NfHusSD0_0),.din(w_dff_A_GXEKt2T89_0),.clk(gclk));
	jdff dff_A_bLcg0G0I9_0(.dout(w_dff_A_GXEKt2T89_0),.din(w_dff_A_bLcg0G0I9_0),.clk(gclk));
	jdff dff_A_jXpx4bnO2_0(.dout(w_dff_A_bLcg0G0I9_0),.din(w_dff_A_jXpx4bnO2_0),.clk(gclk));
	jdff dff_A_1nL2d3l84_0(.dout(w_dff_A_jXpx4bnO2_0),.din(w_dff_A_1nL2d3l84_0),.clk(gclk));
	jdff dff_A_DXADtZmy9_0(.dout(w_dff_A_1nL2d3l84_0),.din(w_dff_A_DXADtZmy9_0),.clk(gclk));
	jdff dff_A_IUELqlgn3_0(.dout(w_dff_A_DXADtZmy9_0),.din(w_dff_A_IUELqlgn3_0),.clk(gclk));
	jdff dff_A_78fXIHfE7_0(.dout(w_dff_A_IUELqlgn3_0),.din(w_dff_A_78fXIHfE7_0),.clk(gclk));
	jdff dff_A_WBG4S1Ro9_0(.dout(w_dff_A_78fXIHfE7_0),.din(w_dff_A_WBG4S1Ro9_0),.clk(gclk));
	jdff dff_A_azHUBSfr1_0(.dout(w_dff_A_WBG4S1Ro9_0),.din(w_dff_A_azHUBSfr1_0),.clk(gclk));
	jdff dff_A_OvFkGplN9_0(.dout(w_Gid28_0[0]),.din(w_dff_A_OvFkGplN9_0),.clk(gclk));
	jdff dff_A_pjxyb87j2_0(.dout(w_dff_A_OvFkGplN9_0),.din(w_dff_A_pjxyb87j2_0),.clk(gclk));
	jdff dff_A_9dhgkiV36_0(.dout(w_dff_A_pjxyb87j2_0),.din(w_dff_A_9dhgkiV36_0),.clk(gclk));
	jdff dff_A_uSrkTRLw1_0(.dout(w_dff_A_9dhgkiV36_0),.din(w_dff_A_uSrkTRLw1_0),.clk(gclk));
	jdff dff_A_KTtfpoyp0_0(.dout(w_dff_A_uSrkTRLw1_0),.din(w_dff_A_KTtfpoyp0_0),.clk(gclk));
	jdff dff_A_6uFoeYcl2_0(.dout(w_dff_A_KTtfpoyp0_0),.din(w_dff_A_6uFoeYcl2_0),.clk(gclk));
	jdff dff_A_Mad77qnx2_0(.dout(w_dff_A_6uFoeYcl2_0),.din(w_dff_A_Mad77qnx2_0),.clk(gclk));
	jdff dff_A_fu0y72oP4_0(.dout(w_dff_A_Mad77qnx2_0),.din(w_dff_A_fu0y72oP4_0),.clk(gclk));
	jdff dff_A_WrbW5WG71_0(.dout(w_dff_A_fu0y72oP4_0),.din(w_dff_A_WrbW5WG71_0),.clk(gclk));
	jdff dff_A_zYdL2D6e2_0(.dout(w_dff_A_WrbW5WG71_0),.din(w_dff_A_zYdL2D6e2_0),.clk(gclk));
	jdff dff_A_C0FtiK1q2_0(.dout(w_dff_A_zYdL2D6e2_0),.din(w_dff_A_C0FtiK1q2_0),.clk(gclk));
	jdff dff_A_xZbhjjVs0_0(.dout(w_Gid31_0[0]),.din(w_dff_A_xZbhjjVs0_0),.clk(gclk));
	jdff dff_A_xEvsVRYM8_0(.dout(w_dff_A_xZbhjjVs0_0),.din(w_dff_A_xEvsVRYM8_0),.clk(gclk));
	jdff dff_A_6cnefFmO1_0(.dout(w_dff_A_xEvsVRYM8_0),.din(w_dff_A_6cnefFmO1_0),.clk(gclk));
	jdff dff_A_dqvs45f62_0(.dout(w_dff_A_6cnefFmO1_0),.din(w_dff_A_dqvs45f62_0),.clk(gclk));
	jdff dff_A_tSlxDHv67_0(.dout(w_dff_A_dqvs45f62_0),.din(w_dff_A_tSlxDHv67_0),.clk(gclk));
	jdff dff_A_4hMMClrs5_0(.dout(w_dff_A_tSlxDHv67_0),.din(w_dff_A_4hMMClrs5_0),.clk(gclk));
	jdff dff_A_BC7Rpd9W8_0(.dout(w_dff_A_4hMMClrs5_0),.din(w_dff_A_BC7Rpd9W8_0),.clk(gclk));
	jdff dff_A_y0DY56H69_0(.dout(w_dff_A_BC7Rpd9W8_0),.din(w_dff_A_y0DY56H69_0),.clk(gclk));
	jdff dff_A_Osg1ps4M8_0(.dout(w_dff_A_y0DY56H69_0),.din(w_dff_A_Osg1ps4M8_0),.clk(gclk));
	jdff dff_A_su0c3OnU2_0(.dout(w_dff_A_Osg1ps4M8_0),.din(w_dff_A_su0c3OnU2_0),.clk(gclk));
	jdff dff_A_ErCKavnX3_0(.dout(w_dff_A_su0c3OnU2_0),.din(w_dff_A_ErCKavnX3_0),.clk(gclk));
	jdff dff_A_R0VntRor0_0(.dout(w_Gid30_0[0]),.din(w_dff_A_R0VntRor0_0),.clk(gclk));
	jdff dff_A_5kiC1pva1_0(.dout(w_dff_A_R0VntRor0_0),.din(w_dff_A_5kiC1pva1_0),.clk(gclk));
	jdff dff_A_fYFzoGo40_0(.dout(w_dff_A_5kiC1pva1_0),.din(w_dff_A_fYFzoGo40_0),.clk(gclk));
	jdff dff_A_krNofpEG7_0(.dout(w_dff_A_fYFzoGo40_0),.din(w_dff_A_krNofpEG7_0),.clk(gclk));
	jdff dff_A_AjSCsUfW6_0(.dout(w_dff_A_krNofpEG7_0),.din(w_dff_A_AjSCsUfW6_0),.clk(gclk));
	jdff dff_A_6HlXHswn6_0(.dout(w_dff_A_AjSCsUfW6_0),.din(w_dff_A_6HlXHswn6_0),.clk(gclk));
	jdff dff_A_vpL9BUYb6_0(.dout(w_dff_A_6HlXHswn6_0),.din(w_dff_A_vpL9BUYb6_0),.clk(gclk));
	jdff dff_A_yZj45uEo2_0(.dout(w_dff_A_vpL9BUYb6_0),.din(w_dff_A_yZj45uEo2_0),.clk(gclk));
	jdff dff_A_pDS8zIsB7_0(.dout(w_dff_A_yZj45uEo2_0),.din(w_dff_A_pDS8zIsB7_0),.clk(gclk));
	jdff dff_A_aBvtiYMn9_0(.dout(w_dff_A_pDS8zIsB7_0),.din(w_dff_A_aBvtiYMn9_0),.clk(gclk));
	jdff dff_A_iJKwPfTv6_0(.dout(w_dff_A_aBvtiYMn9_0),.din(w_dff_A_iJKwPfTv6_0),.clk(gclk));
	jdff dff_A_PMYQK5Tj0_2(.dout(God0),.din(w_dff_A_PMYQK5Tj0_2),.clk(gclk));
	jdff dff_A_5M6o6Ub95_2(.dout(God1),.din(w_dff_A_5M6o6Ub95_2),.clk(gclk));
	jdff dff_A_34PC55qj0_2(.dout(God2),.din(w_dff_A_34PC55qj0_2),.clk(gclk));
	jdff dff_A_VTAVybd45_2(.dout(God3),.din(w_dff_A_VTAVybd45_2),.clk(gclk));
	jdff dff_A_Fwn0Ij8d6_2(.dout(God4),.din(w_dff_A_Fwn0Ij8d6_2),.clk(gclk));
	jdff dff_A_n7m9VX7F7_2(.dout(God5),.din(w_dff_A_n7m9VX7F7_2),.clk(gclk));
	jdff dff_A_PYCXl0ap5_2(.dout(God6),.din(w_dff_A_PYCXl0ap5_2),.clk(gclk));
	jdff dff_A_XgvbmHBM3_2(.dout(God7),.din(w_dff_A_XgvbmHBM3_2),.clk(gclk));
	jdff dff_A_SsQEgfrU1_2(.dout(God8),.din(w_dff_A_SsQEgfrU1_2),.clk(gclk));
	jdff dff_A_P1nnemrt1_2(.dout(God9),.din(w_dff_A_P1nnemrt1_2),.clk(gclk));
	jdff dff_A_YC1eikXb3_2(.dout(God10),.din(w_dff_A_YC1eikXb3_2),.clk(gclk));
	jdff dff_A_gri3Jqev7_2(.dout(God11),.din(w_dff_A_gri3Jqev7_2),.clk(gclk));
	jdff dff_A_wRRP0kLL9_2(.dout(God12),.din(w_dff_A_wRRP0kLL9_2),.clk(gclk));
	jdff dff_A_4nkykmME2_2(.dout(God13),.din(w_dff_A_4nkykmME2_2),.clk(gclk));
	jdff dff_A_UxhabKGn3_2(.dout(God14),.din(w_dff_A_UxhabKGn3_2),.clk(gclk));
	jdff dff_A_7GIr0kJS3_2(.dout(God15),.din(w_dff_A_7GIr0kJS3_2),.clk(gclk));
endmodule

