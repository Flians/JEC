/*

c1908:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 1045
	jand: 128
	jor: 102

Summary:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 1045
	jand: 128
	jor: 102
*/

module c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n202;
	wire n204;
	wire n205;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n222;
	wire n224;
	wire n225;
	wire n226;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire[2:0] w_G101_0;
	wire[2:0] w_G104_0;
	wire[2:0] w_G107_0;
	wire[2:0] w_G110_0;
	wire[1:0] w_G110_1;
	wire[1:0] w_G113_0;
	wire[2:0] w_G116_0;
	wire[2:0] w_G119_0;
	wire[2:0] w_G122_0;
	wire[1:0] w_G122_1;
	wire[2:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[1:0] w_G128_1;
	wire[1:0] w_G131_0;
	wire[2:0] w_G134_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G140_0;
	wire[2:0] w_G143_0;
	wire[1:0] w_G143_1;
	wire[2:0] w_G146_0;
	wire[2:0] w_G210_0;
	wire[1:0] w_G214_0;
	wire[2:0] w_G217_0;
	wire[1:0] w_G221_0;
	wire[1:0] w_G224_0;
	wire[1:0] w_G227_0;
	wire[2:0] w_G234_0;
	wire[2:0] w_G237_0;
	wire[2:0] w_G469_0;
	wire[1:0] w_G472_0;
	wire[2:0] w_G475_0;
	wire[2:0] w_G478_0;
	wire[2:0] w_G902_0;
	wire[2:0] w_G902_1;
	wire[2:0] w_G902_2;
	wire[2:0] w_G902_3;
	wire[2:0] w_G952_0;
	wire[2:0] w_G953_0;
	wire[2:0] w_G953_1;
	wire[1:0] w_n59_0;
	wire[2:0] w_n60_0;
	wire[2:0] w_n61_0;
	wire[2:0] w_n61_1;
	wire[2:0] w_n61_2;
	wire[2:0] w_n61_3;
	wire[1:0] w_n62_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n68_0;
	wire[2:0] w_n70_0;
	wire[2:0] w_n70_1;
	wire[2:0] w_n70_2;
	wire[1:0] w_n70_3;
	wire[1:0] w_n71_0;
	wire[1:0] w_n73_0;
	wire[2:0] w_n74_0;
	wire[1:0] w_n74_1;
	wire[1:0] w_n77_0;
	wire[1:0] w_n79_0;
	wire[2:0] w_n81_0;
	wire[1:0] w_n82_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[2:0] w_n90_0;
	wire[2:0] w_n92_0;
	wire[2:0] w_n92_1;
	wire[2:0] w_n93_0;
	wire[1:0] w_n94_0;
	wire[2:0] w_n95_0;
	wire[2:0] w_n96_0;
	wire[1:0] w_n97_0;
	wire[1:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[2:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n109_0;
	wire[2:0] w_n110_0;
	wire[2:0] w_n112_0;
	wire[1:0] w_n112_1;
	wire[2:0] w_n117_0;
	wire[1:0] w_n118_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[2:0] w_n121_0;
	wire[1:0] w_n121_1;
	wire[1:0] w_n122_0;
	wire[2:0] w_n130_0;
	wire[1:0] w_n131_0;
	wire[2:0] w_n132_0;
	wire[2:0] w_n141_0;
	wire[1:0] w_n142_0;
	wire[2:0] w_n143_0;
	wire[1:0] w_n143_1;
	wire[2:0] w_n144_0;
	wire[2:0] w_n144_1;
	wire[1:0] w_n145_0;
	wire[1:0] w_n146_0;
	wire[1:0] w_n147_0;
	wire[2:0] w_n151_0;
	wire[1:0] w_n152_0;
	wire[2:0] w_n153_0;
	wire[2:0] w_n154_0;
	wire[1:0] w_n154_1;
	wire[2:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[2:0] w_n158_0;
	wire[1:0] w_n158_1;
	wire[2:0] w_n159_0;
	wire[1:0] w_n159_1;
	wire[1:0] w_n160_0;
	wire[2:0] w_n161_0;
	wire[1:0] w_n162_0;
	wire[2:0] w_n163_0;
	wire[1:0] w_n164_0;
	wire[2:0] w_n166_0;
	wire[1:0] w_n166_1;
	wire[1:0] w_n167_0;
	wire[2:0] w_n168_0;
	wire[1:0] w_n169_0;
	wire[1:0] w_n172_0;
	wire[2:0] w_n174_0;
	wire[1:0] w_n174_1;
	wire[1:0] w_n175_0;
	wire[1:0] w_n177_0;
	wire[2:0] w_n179_0;
	wire[1:0] w_n180_0;
	wire[2:0] w_n181_0;
	wire[2:0] w_n183_0;
	wire[2:0] w_n184_0;
	wire[1:0] w_n184_1;
	wire[2:0] w_n185_0;
	wire[1:0] w_n186_0;
	wire[2:0] w_n188_0;
	wire[1:0] w_n189_0;
	wire[1:0] w_n190_0;
	wire[2:0] w_n192_0;
	wire[1:0] w_n193_0;
	wire[2:0] w_n196_0;
	wire[2:0] w_n197_0;
	wire[1:0] w_n197_1;
	wire[2:0] w_n198_0;
	wire[1:0] w_n198_1;
	wire[1:0] w_n199_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n202_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n212_0;
	wire[1:0] w_n213_0;
	wire[2:0] w_n216_0;
	wire[2:0] w_n217_0;
	wire[2:0] w_n218_0;
	wire[1:0] w_n218_1;
	wire[1:0] w_n219_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n222_0;
	wire[1:0] w_n226_0;
	wire[1:0] w_n228_0;
	wire[2:0] w_n244_0;
	wire[2:0] w_n244_1;
	wire[2:0] w_n244_2;
	wire[1:0] w_n252_0;
	wire[2:0] w_n253_0;
	wire[2:0] w_n254_0;
	wire[1:0] w_n254_1;
	wire[2:0] w_n273_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n275_0;
	wire[2:0] w_n276_0;
	wire[1:0] w_n276_1;
	wire[1:0] w_n277_0;
	wire[1:0] w_n278_0;
	wire[1:0] w_n280_0;
	wire[2:0] w_n281_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n286_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n289_0;
	wire[2:0] w_n290_0;
	wire[1:0] w_n291_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n309_0;
	wire[2:0] w_n311_0;
	wire[2:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n318_0;
	wire[1:0] w_n325_0;
	wire[1:0] w_n334_0;
	wire[2:0] w_n335_0;
	wire[2:0] w_n335_1;
	wire[1:0] w_n335_2;
	wire[1:0] w_n336_0;
	wire[2:0] w_n340_0;
	wire[2:0] w_n340_1;
	wire[1:0] w_n340_2;
	wire[1:0] w_n346_0;
	wire[1:0] w_n355_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n395_0;
	wire w_dff_B_87bOp2Dn6_0;
	wire w_dff_B_7EPSNGhf3_0;
	wire w_dff_B_n8utcfpF5_0;
	wire w_dff_B_UPSYHjBa0_0;
	wire w_dff_B_RmygajzI7_0;
	wire w_dff_B_xfuKnVey6_0;
	wire w_dff_B_WqfXkezP9_0;
	wire w_dff_B_NXzlyw5l3_0;
	wire w_dff_B_efvta5zN5_1;
	wire w_dff_B_RRIAtJGU4_1;
	wire w_dff_B_SCWmaTYi6_0;
	wire w_dff_B_oeV6Bnr73_0;
	wire w_dff_A_w1LRiMgX4_1;
	wire w_dff_B_ffzbGroE8_2;
	wire w_dff_B_oE9QYs901_2;
	wire w_dff_B_HchSND1N3_0;
	wire w_dff_B_NQnUtYsK0_0;
	wire w_dff_B_2rVMevCL3_1;
	wire w_dff_B_JrWMiEAL9_1;
	wire w_dff_B_CdeKqlzU0_1;
	wire w_dff_B_6UeguRop8_1;
	wire w_dff_B_gbDAL4yQ9_1;
	wire w_dff_B_8YIKaS3Q4_1;
	wire w_dff_B_Ltn759w28_1;
	wire w_dff_B_5MO2mbjK0_1;
	wire w_dff_B_mRxGlBQw8_1;
	wire w_dff_B_0EoOZv3n9_1;
	wire w_dff_B_jtQwMBmn6_1;
	wire w_dff_B_gnaP1tmM2_1;
	wire w_dff_B_6nTKUK5i8_0;
	wire w_dff_B_3XEJPL3B0_0;
	wire w_dff_B_ZQxSm2Hy8_0;
	wire w_dff_B_TgTPCfoI8_0;
	wire w_dff_B_yaPhb7sG4_0;
	wire w_dff_B_QQY9Zqxy4_0;
	wire w_dff_B_MQqHOlKA4_0;
	wire w_dff_B_TEzwHQ728_0;
	wire w_dff_B_Bwi442li8_0;
	wire w_dff_B_PrAKKe2k3_0;
	wire w_dff_B_s46XYIaT3_0;
	wire w_dff_B_QGb7rWg47_0;
	wire w_dff_B_VRCL3miz9_0;
	wire w_dff_B_tCazLvko6_0;
	wire w_dff_A_PLb05sP82_0;
	wire w_dff_A_VwyzMuxh0_0;
	wire w_dff_A_AP0J3wpp0_0;
	wire w_dff_A_VBce0eM76_0;
	wire w_dff_A_iL4p3XwZ7_0;
	wire w_dff_A_8B8EmH428_0;
	wire w_dff_A_xZrc1hw80_0;
	wire w_dff_A_lDlFOIXc2_0;
	wire w_dff_A_da4Fr2co1_0;
	wire w_dff_A_A7DPSFRy2_0;
	wire w_dff_A_VxuOEcPy6_0;
	wire w_dff_A_eclfmUr33_0;
	wire w_dff_A_2CLhYjZW0_0;
	wire w_dff_A_k57PodTn7_0;
	wire w_dff_A_tnTHw7G86_0;
	wire w_dff_B_EMJWFZeT6_1;
	wire w_dff_B_0Lm1mm1f4_1;
	wire w_dff_B_9olJ5uMv3_1;
	wire w_dff_B_5B6R03Jt6_1;
	wire w_dff_B_Gxzs4Bdx9_1;
	wire w_dff_B_sW2URFvA7_1;
	wire w_dff_B_ZCuoqVvF1_1;
	wire w_dff_B_bUGtMhTw1_1;
	wire w_dff_B_k14CYDZ95_1;
	wire w_dff_B_dQFnZUCt6_1;
	wire w_dff_B_WgABFuDi2_1;
	wire w_dff_B_kPV2oe9U6_1;
	wire w_dff_B_hS2AizXh1_0;
	wire w_dff_B_QDQ36sKV7_0;
	wire w_dff_B_N9jgM4oF5_0;
	wire w_dff_B_6IOFgYHm9_0;
	wire w_dff_B_oNTF7GxA0_0;
	wire w_dff_B_3eb7y8xu1_0;
	wire w_dff_B_uqEmhBw49_0;
	wire w_dff_B_VYR1kyWC0_0;
	wire w_dff_B_kIhGJ28b7_0;
	wire w_dff_B_cpqG3vRd2_0;
	wire w_dff_B_C3wiqR8Y3_0;
	wire w_dff_B_LH6297VJ0_0;
	wire w_dff_B_Flx2KE5N8_0;
	wire w_dff_B_xtRc2aEM8_0;
	wire w_dff_A_9xGKUnYC8_0;
	wire w_dff_A_FWOljebP4_0;
	wire w_dff_A_kzXMQSPo7_0;
	wire w_dff_A_e0SIynSB3_0;
	wire w_dff_A_jzaYJtxw4_0;
	wire w_dff_A_xoj7Wjnk8_0;
	wire w_dff_A_rF1peoG50_0;
	wire w_dff_A_WSoTL0gh4_0;
	wire w_dff_A_uPBe1R1J3_0;
	wire w_dff_A_erVE1r2B7_0;
	wire w_dff_A_dE7RRdtE9_0;
	wire w_dff_A_KjJuUzWy9_0;
	wire w_dff_A_NH0SwtXT7_0;
	wire w_dff_A_FmyFiHIR5_0;
	wire w_dff_A_qFbPGn452_0;
	wire w_dff_B_FJJWjWYM7_1;
	wire w_dff_B_k8MqHn3t9_1;
	wire w_dff_B_zwnjIeiK8_1;
	wire w_dff_B_JqS2EPZr7_1;
	wire w_dff_B_5Yzj6bd25_1;
	wire w_dff_B_IRVWZmf29_1;
	wire w_dff_B_aHmAifBI7_1;
	wire w_dff_B_CXKRjkup3_1;
	wire w_dff_B_1XDmuVL00_1;
	wire w_dff_B_NXvphe786_1;
	wire w_dff_B_RFLLM3IV4_1;
	wire w_dff_B_YbF1Pfnz5_1;
	wire w_dff_B_vpfRtk9D0_0;
	wire w_dff_B_o0rhkiDo3_0;
	wire w_dff_B_gwqHUlfu5_0;
	wire w_dff_B_wCo0NCMB2_0;
	wire w_dff_B_jie2EpRX0_0;
	wire w_dff_B_dKYklQW12_0;
	wire w_dff_B_GHXsExDM4_0;
	wire w_dff_B_lE7cFnSs2_0;
	wire w_dff_B_6kwKJZot7_0;
	wire w_dff_B_8EaBU1Eg0_0;
	wire w_dff_B_iq1igln77_0;
	wire w_dff_B_wTMFt1eP9_0;
	wire w_dff_B_E3S5Ybt36_0;
	wire w_dff_B_CDFvh2JA5_0;
	wire w_dff_A_vLkHJ5s99_0;
	wire w_dff_A_Wz3c9hGM8_0;
	wire w_dff_A_XTYGtVyz8_0;
	wire w_dff_A_Rb7KIZkO4_0;
	wire w_dff_A_untx1rbH5_0;
	wire w_dff_A_i1BstMmA3_0;
	wire w_dff_A_P7pfCRud0_0;
	wire w_dff_A_yDVYZKAu3_0;
	wire w_dff_A_T8moYjYn7_0;
	wire w_dff_A_10vTaxdQ8_0;
	wire w_dff_A_ETervw5G5_0;
	wire w_dff_A_YmfehQHz7_0;
	wire w_dff_A_D363rGBi5_0;
	wire w_dff_A_VtVtXx9l5_0;
	wire w_dff_A_BaKcvWCA8_0;
	wire w_dff_B_kb1An8e37_1;
	wire w_dff_B_hnW3HoZl2_1;
	wire w_dff_B_kuaDvfmG2_1;
	wire w_dff_B_YmBqXeyF8_1;
	wire w_dff_B_PHYeC3ry8_1;
	wire w_dff_B_DlHf5knJ6_1;
	wire w_dff_B_s6W44nz43_1;
	wire w_dff_B_yTE4MABn3_1;
	wire w_dff_B_dekRpRMT9_1;
	wire w_dff_B_EhMBCw9K8_1;
	wire w_dff_B_4uSkO2d68_1;
	wire w_dff_B_uNXQ2yTB4_1;
	wire w_dff_B_0Hjd63n28_0;
	wire w_dff_B_hlq442934_0;
	wire w_dff_B_OTEDu9Q83_0;
	wire w_dff_B_EpMVBOMw2_0;
	wire w_dff_B_79oD9aer7_0;
	wire w_dff_B_JGQBD7BZ4_0;
	wire w_dff_B_C12t8k9v5_0;
	wire w_dff_B_oPsM1g8r3_0;
	wire w_dff_B_qmNqaiHI0_0;
	wire w_dff_B_WhlBGXK76_0;
	wire w_dff_B_G4UFy2um8_0;
	wire w_dff_B_PYidTrXO6_0;
	wire w_dff_B_75LSLCq09_0;
	wire w_dff_B_QxbYTAa80_0;
	wire w_dff_A_aiSCGz7O5_0;
	wire w_dff_A_VgYQpamO8_0;
	wire w_dff_A_3FtZ9Gmg3_0;
	wire w_dff_A_EtZfJLHb2_0;
	wire w_dff_A_ReleY0UH9_0;
	wire w_dff_A_Mqyqz53w0_0;
	wire w_dff_A_Ilcp6WiR8_0;
	wire w_dff_A_nVdmpPMU2_0;
	wire w_dff_A_mVvD6MKm1_0;
	wire w_dff_A_n0hF5aWI9_0;
	wire w_dff_A_hlbiBiCn7_0;
	wire w_dff_A_Lbvojlos8_0;
	wire w_dff_A_PpZJM5409_0;
	wire w_dff_A_cSwTILFg5_0;
	wire w_dff_A_bYMbuxKl5_0;
	wire w_dff_B_3rFXgPFh9_1;
	wire w_dff_B_0LY0pZrb6_0;
	wire w_dff_B_ROZDpAaR2_0;
	wire w_dff_B_F01UjAOe8_0;
	wire w_dff_B_ZwaM6reX6_0;
	wire w_dff_B_kXQ6hvyY7_0;
	wire w_dff_B_vvTWKtXD0_0;
	wire w_dff_B_KbPhcMyl3_0;
	wire w_dff_B_gwMoCEKh4_0;
	wire w_dff_B_JJ2FDzwg5_0;
	wire w_dff_B_XrPFzcc91_0;
	wire w_dff_B_QTyRJJdr1_0;
	wire w_dff_B_cPtKHVpI7_0;
	wire w_dff_B_ZPZysFsS6_0;
	wire w_dff_B_r9UUnYqn5_0;
	wire w_dff_A_UlZV1zJ91_1;
	wire w_dff_A_5WXqnS2S7_1;
	wire w_dff_A_9mB84Hqz8_1;
	wire w_dff_A_rp5j1TAM3_1;
	wire w_dff_A_eDYiX4ky7_1;
	wire w_dff_A_NNnaF8UE5_1;
	wire w_dff_A_1VjhMmOB9_1;
	wire w_dff_A_Yc4LdnPn0_1;
	wire w_dff_A_Yzc98HWj1_1;
	wire w_dff_A_7xlSI9do8_1;
	wire w_dff_A_6IxUmO6m5_1;
	wire w_dff_A_SmnZ541m5_1;
	wire w_dff_A_7FwV4aLd3_1;
	wire w_dff_A_a1RD86qw0_1;
	wire w_dff_A_D8Wqng4N3_1;
	wire w_dff_B_Dbri4POt1_1;
	wire w_dff_B_Q7tqGaGw2_1;
	wire w_dff_B_xN5SDyhd0_1;
	wire w_dff_B_gOpwTTqT0_1;
	wire w_dff_B_hXY9ravn1_1;
	wire w_dff_B_AmhuZh2S3_1;
	wire w_dff_B_NhPVS65S6_1;
	wire w_dff_B_nhObHOLc5_1;
	wire w_dff_B_JvCZmWV14_1;
	wire w_dff_B_nHFJlcOV4_1;
	wire w_dff_B_IVn7fjfZ9_1;
	wire w_dff_B_I6gRvqVv4_1;
	wire w_dff_B_ko09xkuE4_1;
	wire w_dff_B_pBnm7llM9_1;
	wire w_dff_B_xmqYbzs75_1;
	wire w_dff_B_bNzKWLox1_0;
	wire w_dff_B_EbHeg9E11_0;
	wire w_dff_B_MATPjOp15_0;
	wire w_dff_B_nRgoqobJ7_0;
	wire w_dff_B_uOBEpA8d6_0;
	wire w_dff_B_pMFW7uyy6_0;
	wire w_dff_B_QGtF6uyi2_0;
	wire w_dff_B_1iYajag89_0;
	wire w_dff_B_xfUySCc40_0;
	wire w_dff_B_Ssv97t0V0_0;
	wire w_dff_B_yXH21rMx8_0;
	wire w_dff_B_WCNOHD9j6_0;
	wire w_dff_B_EDuWhzQ47_0;
	wire w_dff_B_L3uD0Hyc4_0;
	wire w_dff_B_FuQFQQAz1_0;
	wire w_dff_B_3BVc73Hu4_0;
	wire w_dff_B_ls4aoIiI5_0;
	wire w_dff_B_y831cesS0_0;
	wire w_dff_B_tK02ByYW3_0;
	wire w_dff_B_cupCJfLT3_0;
	wire w_dff_B_XHdNCY1C0_0;
	wire w_dff_B_a43oumxU9_0;
	wire w_dff_B_81GGm6a58_0;
	wire w_dff_B_8D8R4uzi7_0;
	wire w_dff_B_Wxwyns1d6_0;
	wire w_dff_B_i2ZLgkmr8_1;
	wire w_dff_B_8j7wOmlc8_1;
	wire w_dff_B_6LORq5xz3_0;
	wire w_dff_B_TugF7XTs1_0;
	wire w_dff_B_vmoqKux69_0;
	wire w_dff_B_j9CgkoDt0_0;
	wire w_dff_B_cUjSGt0f8_0;
	wire w_dff_B_6Oq4KqUR5_0;
	wire w_dff_B_UuKCp4g08_0;
	wire w_dff_B_yPMVfwtr6_0;
	wire w_dff_B_3JxjyQcm6_0;
	wire w_dff_B_9latNVrB7_0;
	wire w_dff_B_J81RkvBt1_0;
	wire w_dff_B_hWJJgJB85_0;
	wire w_dff_B_3QYbYrbm0_0;
	wire w_dff_B_FlWjvmng7_1;
	wire w_dff_B_XkZapgF37_0;
	wire w_dff_A_qOvmg9cl6_0;
	wire w_dff_A_vH4ZGHON8_0;
	wire w_dff_A_ZagKAg6M8_2;
	wire w_dff_A_M7YcBVR91_2;
	wire w_dff_A_hGQAbzib8_0;
	wire w_dff_A_j8MwRq0V6_2;
	wire w_dff_B_irItOaNe5_3;
	wire w_dff_B_KIiYPtj29_0;
	wire w_dff_A_FQT5dyl84_0;
	wire w_dff_A_ZVxorm683_2;
	wire w_dff_A_Hafs6tmu3_2;
	wire w_dff_A_dBmESVvk1_0;
	wire w_dff_A_SkE9QDgu5_0;
	wire w_dff_A_xphs99ls2_1;
	wire w_dff_A_hsnnmuCv1_1;
	wire w_dff_A_pkz4VgKi7_0;
	wire w_dff_A_U7V0YSX17_2;
	wire w_dff_B_MkLyWnOY7_3;
	wire w_dff_A_Z0sc88C71_0;
	wire w_dff_A_LS0OlbDu1_0;
	wire w_dff_A_ezwITuSn2_1;
	wire w_dff_A_k8eG48ky1_1;
	wire w_dff_A_QpL5amcm0_2;
	wire w_dff_A_xZt7LRzF2_2;
	wire w_dff_A_GnX2E4J12_2;
	wire w_dff_B_m8neVkhE9_3;
	wire w_dff_A_XWqpTgAq9_1;
	wire w_dff_A_EWvyHitg1_1;
	wire w_dff_A_ZACxQElf1_1;
	wire w_dff_A_l9XTGDeg8_1;
	wire w_dff_A_npN2hmbO2_2;
	wire w_dff_A_2FZx9MYs5_2;
	wire w_dff_A_l35YzkKC2_2;
	wire w_dff_A_fHH7YDY19_2;
	wire w_dff_B_pLektpro5_3;
	wire w_dff_B_H8ARiGba5_3;
	wire w_dff_B_6yfJjcJB8_3;
	wire w_dff_B_9H8gVqG19_3;
	wire w_dff_B_ompYDYwR9_3;
	wire w_dff_B_MUwemsSK1_3;
	wire w_dff_B_DTKlaCO11_3;
	wire w_dff_B_rN5AlINv4_3;
	wire w_dff_B_IWPAWgS61_3;
	wire w_dff_B_9d9lGbvZ4_3;
	wire w_dff_B_flcQQ9b53_3;
	wire w_dff_B_dj9wFQAO7_3;
	wire w_dff_B_9i4j02lf4_3;
	wire w_dff_B_swvHy0uK6_3;
	wire w_dff_B_7JHBBpwe3_3;
	wire w_dff_B_zDweCeiP0_3;
	wire w_dff_B_pG1xOg5Q9_1;
	wire w_dff_B_g28bMA9v8_1;
	wire w_dff_B_hllqSuK67_1;
	wire w_dff_B_g7eQvssc8_1;
	wire w_dff_B_tls9DdDw4_1;
	wire w_dff_B_OLaJSHoj9_1;
	wire w_dff_B_nysGo9QM1_1;
	wire w_dff_B_r86hjLOJ8_1;
	wire w_dff_B_iYKnZW357_1;
	wire w_dff_B_dFZsLN1Y7_1;
	wire w_dff_B_MRxDTQWd2_1;
	wire w_dff_B_dEAPrYKo2_0;
	wire w_dff_B_w2JDPKYv3_0;
	wire w_dff_B_VGT2LlO66_0;
	wire w_dff_B_yQodEHlx0_0;
	wire w_dff_B_KPuWEk0j7_0;
	wire w_dff_B_bbrLuMRc2_0;
	wire w_dff_B_X306fpbu2_0;
	wire w_dff_B_GGY02Drb7_0;
	wire w_dff_B_Oie8pYVk4_0;
	wire w_dff_B_NYJln6Np0_0;
	wire w_dff_B_1StzCjHM6_0;
	wire w_dff_B_rkG1HUsr8_0;
	wire w_dff_B_EQJPGoen2_0;
	wire w_dff_B_cXxrWteb3_0;
	wire w_dff_A_NIax9h3X6_0;
	wire w_dff_A_iKKKJ23l9_0;
	wire w_dff_A_xlTmhS4j5_0;
	wire w_dff_A_IXviYaWx1_0;
	wire w_dff_A_kTeVdeRX4_0;
	wire w_dff_A_SE7hUOsb9_0;
	wire w_dff_A_swHCo9AP2_0;
	wire w_dff_A_Vrwm4S622_0;
	wire w_dff_A_gbnZpzJY2_0;
	wire w_dff_A_M7iHoaWE9_0;
	wire w_dff_A_GYTrGeeS0_0;
	wire w_dff_A_q4Y4a0Yf6_0;
	wire w_dff_A_8hE18YhF3_0;
	wire w_dff_A_kyDYNBv42_0;
	wire w_dff_A_j9yRjunC8_0;
	wire w_dff_B_48Z0yb8N8_0;
	wire w_dff_B_Z1qjeC8T8_0;
	wire w_dff_A_TcrzHSSq9_1;
	wire w_dff_A_TmET4rrF7_1;
	wire w_dff_B_DjmXnYWK5_2;
	wire w_dff_A_8FL7BuWU7_1;
	wire w_dff_A_PmJZcSWs4_1;
	wire w_dff_A_RaitYgNH5_2;
	wire w_dff_A_Mzvb4cNp0_2;
	wire w_dff_B_M7qw6BmR9_3;
	wire w_dff_B_pOEkBLmB1_3;
	wire w_dff_A_zxpVdtJC4_0;
	wire w_dff_A_S0gXY9FI0_1;
	wire w_dff_B_NvAM7Nba6_3;
	wire w_dff_A_B1jwbQ744_1;
	wire w_dff_A_VmapFO1s6_2;
	wire w_dff_B_raYUAsUH5_3;
	wire w_dff_A_bALUpook7_0;
	wire w_dff_A_GLbWVTBc5_0;
	wire w_dff_A_724vyw0z0_0;
	wire w_dff_A_6xpSDlhg7_1;
	wire w_dff_A_v9IRINiZ2_1;
	wire w_dff_A_QPbox9xq7_1;
	wire w_dff_B_CKUBDPhr6_0;
	wire w_dff_B_vaIuTYF12_1;
	wire w_dff_B_PSFF9oYg4_0;
	wire w_dff_A_jiVXwrw15_1;
	wire w_dff_A_DPVzRc6d1_0;
	wire w_dff_B_TEqAAgl68_3;
	wire w_dff_A_xVKWZllH7_0;
	wire w_dff_A_FlTTx5ZE9_0;
	wire w_dff_B_owlxZTpc5_3;
	wire w_dff_A_zc2exPZ20_0;
	wire w_dff_A_mNchYbv10_0;
	wire w_dff_A_OFRntSuX5_2;
	wire w_dff_A_uma05frZ8_2;
	wire w_dff_B_rjIpW8xh5_2;
	wire w_dff_A_rmQXyUD25_1;
	wire w_dff_A_LI1M4O6h8_1;
	wire w_dff_A_qBFBJK5w9_2;
	wire w_dff_A_RUEtXAqY8_2;
	wire w_dff_B_Qp1ZNaVn8_1;
	wire w_dff_B_LM6CR5XI4_1;
	wire w_dff_B_HvLhY8AC0_1;
	wire w_dff_B_5Joslp8J0_1;
	wire w_dff_B_c9ZLC9CU5_1;
	wire w_dff_A_7J0PynwU1_0;
	wire w_dff_A_mAI8a6530_0;
	wire w_dff_A_VYcFzFhk6_0;
	wire w_dff_A_XWYVQCkV9_0;
	wire w_dff_A_pF8YWz8c8_0;
	wire w_dff_A_Exlr2Eoo1_0;
	wire w_dff_A_BYVIeeHr4_0;
	wire w_dff_A_vjDNgY8s5_0;
	wire w_dff_A_YlonpCgY7_0;
	wire w_dff_A_TCZ09ifv2_0;
	wire w_dff_A_IrqCsY0U8_0;
	wire w_dff_A_juWZbGN95_1;
	wire w_dff_B_bEywQSYi2_3;
	wire w_dff_B_bdT2QtA68_2;
	wire w_dff_A_Tz13o3B98_1;
	wire w_dff_A_GoMmkFZB3_1;
	wire w_dff_A_LD3Dv2xE4_2;
	wire w_dff_A_5TdxSzju1_2;
	wire w_dff_B_5bAE8v1W6_1;
	wire w_dff_B_yBRMCjK85_1;
	wire w_dff_B_8L2iblMT8_1;
	wire w_dff_B_zqYjqX8i2_1;
	wire w_dff_B_0iPv6gzG1_1;
	wire w_dff_A_rEBYjwos2_0;
	wire w_dff_A_7e25JeQW8_0;
	wire w_dff_A_Bbeih4ml6_0;
	wire w_dff_A_05gUz8eC3_0;
	wire w_dff_A_bH7EHXLC5_0;
	wire w_dff_A_X13iLN897_0;
	wire w_dff_A_uiojGWRL6_0;
	wire w_dff_A_JjRXqtp87_0;
	wire w_dff_A_7x6m75oJ1_0;
	wire w_dff_A_DExDTuAx1_0;
	wire w_dff_A_mk4gPCmd3_0;
	wire w_dff_A_rGr1XINl7_0;
	wire w_dff_B_jnzZwyXB6_1;
	wire w_dff_B_L8QKAwC11_1;
	wire w_dff_A_53JJPNRr4_1;
	wire w_dff_A_o3uS6aLv0_1;
	wire w_dff_A_DM8gqVOJ3_1;
	wire w_dff_A_l6FC1KZH0_1;
	wire w_dff_A_I28831662_1;
	wire w_dff_A_OxoHZ5Ps2_1;
	wire w_dff_A_LQhley7s3_0;
	wire w_dff_A_nnlDv0iF6_0;
	wire w_dff_A_UYoiRhCm8_0;
	wire w_dff_A_GN3tzEEp0_0;
	wire w_dff_A_DMDHVcJa9_0;
	wire w_dff_A_Uk705U1L4_0;
	wire w_dff_A_hTrlKjcn8_0;
	wire w_dff_A_ibCtApuJ3_0;
	wire w_dff_A_32W4jJMI8_0;
	wire w_dff_A_x0jYfg461_0;
	wire w_dff_A_25ba2pdN7_0;
	wire w_dff_A_VM9zdHHW2_0;
	wire w_dff_B_bdvoMKgx8_1;
	wire w_dff_B_t0UNrw4Z3_1;
	wire w_dff_B_IEDcSjra0_1;
	wire w_dff_B_fzf9OgLb8_0;
	wire w_dff_A_CtGg71EJ0_1;
	wire w_dff_A_wXDaLGka3_1;
	wire w_dff_A_p6SYAq3i8_1;
	wire w_dff_A_EeA4weBH6_1;
	wire w_dff_A_A1OTIQDY1_1;
	wire w_dff_A_HidJcISd9_1;
	wire w_dff_B_cI1V1wQt5_3;
	wire w_dff_B_TII2KWyq0_3;
	wire w_dff_A_VM14KFsj4_0;
	wire w_dff_A_pt6Y1sLI2_0;
	wire w_dff_A_7y0MB23R2_0;
	wire w_dff_A_Da3mUR3W3_1;
	wire w_dff_A_GVKFDLUy0_1;
	wire w_dff_A_rICxkPtJ8_1;
	wire w_dff_B_1zEFzQYj5_1;
	wire w_dff_A_hupSypvR0_0;
	wire w_dff_A_9hQcCyMw8_1;
	wire w_dff_A_Yp6jucyo8_1;
	wire w_dff_A_VX7vXtxt6_1;
	wire w_dff_A_6DZDx5TQ8_1;
	wire w_dff_A_NrfbGgaG0_1;
	wire w_dff_A_XrWe4vcE5_1;
	wire w_dff_A_8voFaRrL2_1;
	wire w_dff_A_YuDYZB8u6_1;
	wire w_dff_A_11mm1uNl8_1;
	wire w_dff_A_AtNUKxE55_1;
	wire w_dff_A_IbXovPq23_1;
	wire w_dff_A_Tfcn9HTa0_1;
	wire w_dff_A_ZMW53MW68_1;
	wire w_dff_A_Vjc72R8L5_1;
	wire w_dff_A_1vw4cqIS8_1;
	wire w_dff_A_SUlDxw8x9_1;
	wire w_dff_A_r5d4qCrU5_1;
	wire w_dff_A_fWz20p4R0_1;
	wire w_dff_A_7Us8wD3e1_1;
	wire w_dff_A_U131JysR2_1;
	wire w_dff_A_saO30qQ77_1;
	wire w_dff_A_DmHOwzrL9_1;
	wire w_dff_A_IoiwkHxL6_1;
	wire w_dff_A_pNwj3ERr8_1;
	wire w_dff_A_pv0B8K8e8_1;
	wire w_dff_A_wWPGREJB6_1;
	wire w_dff_A_tcPEUmQq8_1;
	wire w_dff_B_23RAqRpQ9_3;
	wire w_dff_B_7Y2DWtMV5_1;
	wire w_dff_A_9iLFHuQA5_2;
	wire w_dff_A_IAxImSs79_1;
	wire w_dff_A_6LwPzpr78_1;
	wire w_dff_A_QeIaXzPy7_2;
	wire w_dff_A_j7Zy7O2B8_2;
	wire w_dff_A_CvDs9rKb2_1;
	wire w_dff_A_0p0bzACN2_1;
	wire w_dff_A_cMFhgO2J9_1;
	wire w_dff_A_NTcFWbYE3_1;
	wire w_dff_A_HvS80Czb7_1;
	wire w_dff_A_j5LbCEsr0_1;
	wire w_dff_B_3HrIOuAs7_2;
	wire w_dff_B_gSd8pB4c1_2;
	wire w_dff_B_n1oB1xGr7_2;
	wire w_dff_B_AJ4NIPbd6_2;
	wire w_dff_A_B7k92NuB0_1;
	wire w_dff_A_zl8609TL1_1;
	wire w_dff_A_gAP7lnGJ9_2;
	wire w_dff_A_QFYNjmhw9_2;
	wire w_dff_A_0FYkV1dJ2_2;
	wire w_dff_A_L5vz5Btl7_0;
	wire w_dff_A_01SBQoWa6_0;
	wire w_dff_A_gE7Nowti9_0;
	wire w_dff_A_zBOTKbEV6_0;
	wire w_dff_A_iHmhUX007_0;
	wire w_dff_A_6HqoROxp0_0;
	wire w_dff_A_klwCKbVv7_0;
	wire w_dff_A_Cnsov7UN0_0;
	wire w_dff_A_KoiLVggi2_0;
	wire w_dff_A_i59WwYfY7_0;
	wire w_dff_B_vGQlEkZ78_1;
	wire w_dff_B_Bw6YcVAi9_1;
	wire w_dff_B_MBQeGfwG0_1;
	wire w_dff_B_iV8nUqg47_0;
	wire w_dff_B_NNq6FVvX2_0;
	wire w_dff_B_BelyrYIz1_0;
	wire w_dff_A_fFZrmiXs5_2;
	wire w_dff_A_AmL7gSWu2_2;
	wire w_dff_A_rUkWVoqt7_2;
	wire w_dff_A_honyHz3o2_2;
	wire w_dff_A_rQXRt57y5_0;
	wire w_dff_A_UIGrPf6h3_0;
	wire w_dff_A_NRjXV6Yh0_0;
	wire w_dff_A_814i3DzR1_0;
	wire w_dff_A_qM7cLgsS9_0;
	wire w_dff_A_IQMPX2U20_0;
	wire w_dff_A_YeUhj9EY4_0;
	wire w_dff_A_tjj0vqVn2_0;
	wire w_dff_A_PyS38Hry9_0;
	wire w_dff_A_W8ddvjR15_2;
	wire w_dff_A_iRp9Pgqu7_2;
	wire w_dff_A_6Stgew7U1_2;
	wire w_dff_A_zWlwC2Ou2_2;
	wire w_dff_A_aK5RmE8l4_0;
	wire w_dff_B_Noibk2AT2_3;
	wire w_dff_B_wO5IPQdQ4_1;
	wire w_dff_B_DoqiWlGc8_1;
	wire w_dff_B_054wAfNi9_1;
	wire w_dff_B_YiO9UU9a3_1;
	wire w_dff_B_IDrOGnTz9_1;
	wire w_dff_A_g1zixX7E3_0;
	wire w_dff_A_tpkSHp4F4_0;
	wire w_dff_A_vXyxFrkh0_0;
	wire w_dff_A_EHajfGsu6_0;
	wire w_dff_A_AUESdjAj7_0;
	wire w_dff_A_ehIEWmHZ3_0;
	wire w_dff_A_2g9Q7j5z3_0;
	wire w_dff_A_B7KGnKDP7_0;
	wire w_dff_A_smkwssbt8_0;
	wire w_dff_A_mfNqk30O9_0;
	wire w_dff_A_j87yRcQF3_0;
	wire w_dff_A_VzVx22lW7_0;
	wire w_dff_B_eKKvfRZ89_1;
	wire w_dff_B_eXj6DoYl4_1;
	wire w_dff_B_cFSZjj0a2_2;
	wire w_dff_A_leZGNIq02_0;
	wire w_dff_A_1PN84TZ54_0;
	wire w_dff_A_FzLgC7cX9_0;
	wire w_dff_A_4gt6HTaA9_0;
	wire w_dff_A_AnPH0Xfn5_0;
	wire w_dff_A_aVzZ3h7f1_0;
	wire w_dff_A_CFJD27Pf8_0;
	wire w_dff_A_0CqJW5CV4_0;
	wire w_dff_A_VrUYHfgX8_0;
	wire w_dff_A_w2N3Q8iA4_0;
	wire w_dff_A_CmjkHV433_0;
	wire w_dff_A_YVDvWf2Z5_0;
	wire w_dff_A_kYbTGiMo9_2;
	wire w_dff_A_oZdnrC5n2_2;
	wire w_dff_A_Ih4YruBg6_2;
	wire w_dff_A_QMRJReU24_2;
	wire w_dff_A_J7KElagk8_2;
	wire w_dff_A_kUKg9n2E9_2;
	wire w_dff_B_DmgtZOLf4_2;
	wire w_dff_B_7kQIQ15r4_2;
	wire w_dff_B_IxfoKFtQ6_2;
	wire w_dff_A_EdUnV6IY8_0;
	wire w_dff_A_u3i1uTpQ7_0;
	wire w_dff_A_dcsRzTbO3_0;
	wire w_dff_A_QhbAil4O7_0;
	wire w_dff_B_rah6lkTt0_1;
	wire w_dff_A_3Rl7pbnY6_0;
	wire w_dff_A_redLIpgw6_0;
	wire w_dff_A_WkPdH8WO6_0;
	wire w_dff_A_60j5QT485_0;
	wire w_dff_A_ggVshsIh6_1;
	wire w_dff_A_89kZRE0r3_2;
	wire w_dff_A_2roPytqy0_1;
	wire w_dff_A_yCpBk0Y09_1;
	wire w_dff_A_sv65aGNS4_1;
	wire w_dff_B_UGeduBdz0_1;
	wire w_dff_B_CkLetjez8_1;
	wire w_dff_B_kUSsOW6B4_1;
	wire w_dff_A_ZHkqUpbp4_0;
	wire w_dff_A_4k2uxTUi5_0;
	wire w_dff_A_Hc370YHl1_0;
	wire w_dff_A_KgxHdDWL2_0;
	wire w_dff_A_JZJ5cXPt2_0;
	wire w_dff_A_dTumLa988_0;
	wire w_dff_A_EvNMH0Mw6_0;
	wire w_dff_A_b34TpyAV9_0;
	wire w_dff_A_E3sWM7kP7_0;
	wire w_dff_A_f7xTYwhE4_0;
	wire w_dff_A_hdnF33qb9_0;
	wire w_dff_A_g1ORjDxT3_0;
	wire w_dff_B_FO9vK7AP2_1;
	wire w_dff_A_PnlwhtQw8_0;
	wire w_dff_A_JZ5m6VnO8_0;
	wire w_dff_A_WGfH91Yx6_0;
	wire w_dff_A_xGpjIgIh5_0;
	wire w_dff_A_zKsRrzPj3_0;
	wire w_dff_A_WDVkUHBz1_0;
	wire w_dff_A_pi9Y8krL5_0;
	wire w_dff_A_486T9eco4_0;
	wire w_dff_A_aqGOVTYM0_0;
	wire w_dff_A_P29qcHQQ6_0;
	wire w_dff_A_ArXJfFfX1_0;
	wire w_dff_A_ZQxUeYFV5_0;
	wire w_dff_A_Yo8kznD37_1;
	wire w_dff_A_nAprNfw33_1;
	wire w_dff_B_Cs8bBDdu8_2;
	wire w_dff_A_ISIF9isV8_0;
	wire w_dff_A_aIhkJofu7_0;
	wire w_dff_A_lNHD9F7Q7_0;
	wire w_dff_A_SECMuhex4_0;
	wire w_dff_A_hNNPIpT05_0;
	wire w_dff_A_A4c9U7eH1_0;
	wire w_dff_A_C4HrPy779_0;
	wire w_dff_A_EngtZWI63_0;
	wire w_dff_A_guHP7NST5_0;
	wire w_dff_A_jh3iVW3D0_0;
	wire w_dff_A_ATqskvdz9_0;
	wire w_dff_A_hCN9fHM94_0;
	wire w_dff_A_wN0Zf4xK3_0;
	wire w_dff_B_dnr6vzjO6_1;
	wire w_dff_A_MDB8iETe1_0;
	wire w_dff_A_ksRPY3xq2_0;
	wire w_dff_A_hWjPEOkq3_0;
	wire w_dff_A_xpQzUwJK8_0;
	wire w_dff_A_h3pQ6Ceu2_0;
	wire w_dff_A_APAWADrK7_0;
	wire w_dff_A_y1czvHnx1_0;
	wire w_dff_A_NO4oX8BS0_0;
	wire w_dff_A_lahtR6aK2_0;
	wire w_dff_A_OjVz81K20_0;
	wire w_dff_A_ix3vRjwt2_0;
	wire w_dff_A_II0a2sMc3_0;
	wire w_dff_A_o5GIHIjc2_0;
	wire w_dff_A_yMyujAxK1_0;
	wire w_dff_A_eouqoC498_0;
	wire w_dff_A_DyTSIePs4_0;
	wire w_dff_A_gZPj3fv32_0;
	wire w_dff_A_dxVpsDi56_0;
	wire w_dff_A_fi8J9VmA6_0;
	wire w_dff_A_o7Kn8B2X4_0;
	wire w_dff_A_z5woJNMy4_0;
	wire w_dff_A_TWFjMZ5A5_0;
	wire w_dff_A_7wFpHwdV9_0;
	wire w_dff_A_JUN6cAtx4_0;
	wire w_dff_A_p2qQeJRt6_1;
	wire w_dff_A_L3g0NJor4_1;
	wire w_dff_A_Ddh5DIGQ4_1;
	wire w_dff_A_k3DB6E8w3_1;
	wire w_dff_A_v1JzMh499_1;
	wire w_dff_A_r1xBo5yf9_1;
	wire w_dff_A_X5HSDzXy6_1;
	wire w_dff_A_AMZjBZ5Q2_1;
	wire w_dff_A_kKuEV2AB0_1;
	wire w_dff_A_BVnIvebr8_1;
	wire w_dff_A_YVVRTht70_1;
	wire w_dff_A_wobpuE6y1_1;
	wire w_dff_A_2Z629HSC4_1;
	wire w_dff_A_SIogjVJG3_1;
	wire w_dff_A_w6arXA8v7_1;
	wire w_dff_A_Ec8Ld3O35_2;
	wire w_dff_A_y6kskGDT1_1;
	wire w_dff_A_YUUqTcvI8_1;
	wire w_dff_A_eKSMDSod0_1;
	wire w_dff_A_MJweIFhr8_1;
	wire w_dff_A_aclXEIyw0_1;
	wire w_dff_A_BRAQ6cGg2_1;
	wire w_dff_A_THMf1PB55_1;
	wire w_dff_A_ZWW6Y2wf2_1;
	wire w_dff_A_lVBgeQoh8_1;
	wire w_dff_A_9rMQASy27_1;
	wire w_dff_A_x4qXe0lD9_1;
	wire w_dff_A_j1Zh2E308_1;
	wire w_dff_A_mh9vj8Iq4_1;
	wire w_dff_A_xdJPCwPR5_1;
	wire w_dff_A_nyPTpRkc4_1;
	wire w_dff_A_QmhLiQbM1_1;
	wire w_dff_A_DssgHyMX5_1;
	wire w_dff_A_XuI57YRK1_1;
	wire w_dff_A_FWBCGhG24_1;
	wire w_dff_A_KmRdp1rA2_1;
	wire w_dff_A_t4wq9cUJ4_1;
	wire w_dff_A_iqaD8r9z4_1;
	wire w_dff_A_lgzrQ1LR2_1;
	wire w_dff_A_9tvp1E123_1;
	wire w_dff_A_VhmM6P478_1;
	wire w_dff_A_snbUpo1Z0_0;
	wire w_dff_A_D50ukLQQ6_0;
	wire w_dff_A_g6rrSMku3_0;
	wire w_dff_A_Hj9aZnJU9_0;
	wire w_dff_A_pp7OSwDu3_0;
	wire w_dff_A_LIv5uAeB7_1;
	wire w_dff_A_Tg4ZrqNW5_1;
	wire w_dff_A_nCCG4xHc5_1;
	wire w_dff_A_oqHOa6lF5_1;
	wire w_dff_A_5I2AiDSb2_1;
	wire w_dff_A_UFa8GZ8p3_2;
	wire w_dff_A_xiag4azV4_2;
	wire w_dff_A_qjYLtkfG3_2;
	wire w_dff_A_nDJp6hBW3_2;
	wire w_dff_A_paufcRPd3_2;
	wire w_dff_A_4i9eyJnQ9_2;
	wire w_dff_A_QRdg40aF4_2;
	wire w_dff_A_WHE8BckL9_1;
	wire w_dff_A_CWymT7yq3_0;
	wire w_dff_A_bO0UbUXO9_0;
	wire w_dff_A_RaerdxAK0_0;
	wire w_dff_A_rjQlVEfz9_0;
	wire w_dff_A_90p0szhD7_0;
	wire w_dff_A_HNI1iM831_0;
	wire w_dff_A_Hh7OsBkk2_0;
	wire w_dff_A_9F4TfS4E5_0;
	wire w_dff_A_OoH6eD4R6_0;
	wire w_dff_A_bZCrDLAh8_0;
	wire w_dff_A_O49NUb3s5_0;
	wire w_dff_A_MCYmCCnC0_0;
	wire w_dff_A_h0Dffoh04_0;
	wire w_dff_A_8nKWwOI41_0;
	wire w_dff_A_NSKguIuh7_0;
	wire w_dff_A_4naNH1m66_0;
	wire w_dff_A_4vTOr4r51_0;
	wire w_dff_A_aeqoslnv0_0;
	wire w_dff_A_qhB5ACh29_0;
	wire w_dff_A_rIfMH1le8_0;
	wire w_dff_A_QTILc4YB6_0;
	wire w_dff_A_brTqkjB06_0;
	wire w_dff_A_w6mxQNlP6_0;
	wire w_dff_A_N8483xR91_0;
	wire w_dff_A_cB1mUdX04_1;
	wire w_dff_A_SEF5qUbG5_1;
	wire w_dff_A_mwoS1c6A6_1;
	wire w_dff_A_rGZpNTE14_1;
	wire w_dff_A_lY0cgKZ79_1;
	wire w_dff_A_sTKLxUYb7_1;
	wire w_dff_A_rmas8ajd6_1;
	wire w_dff_A_qVDZP92s6_1;
	wire w_dff_A_TJTqvTeT9_1;
	wire w_dff_A_dNVObq0U6_1;
	wire w_dff_A_3dbCYNXb1_1;
	wire w_dff_A_1alljOBI3_1;
	wire w_dff_A_8nD2dtlC4_1;
	wire w_dff_A_CUgDdtaZ2_1;
	wire w_dff_A_v8bqlD7a2_1;
	wire w_dff_A_3a2JHqZY5_2;
	wire w_dff_A_VhO82LPz1_2;
	wire w_dff_A_0YJ11Z8j2_2;
	wire w_dff_A_bZeC2siw3_2;
	wire w_dff_A_XlG72CDe4_2;
	wire w_dff_A_7mUSggM42_2;
	wire w_dff_A_2AgwEJ7B3_2;
	wire w_dff_A_VgXDAfB17_2;
	wire w_dff_A_CIoGP6cw2_2;
	wire w_dff_A_NXFnoskI5_2;
	wire w_dff_A_moeBF56a3_2;
	wire w_dff_A_oEcTbdz11_2;
	wire w_dff_A_JhRr7uuN4_2;
	wire w_dff_A_GcbRdbm23_2;
	wire w_dff_A_5XAaL6JI8_2;
	wire w_dff_A_o71ohj0b8_1;
	wire w_dff_A_ZTUYCujP4_0;
	wire w_dff_A_iCXY3wNZ1_0;
	wire w_dff_A_wPhlVCtG5_0;
	wire w_dff_A_jig1QCiK7_0;
	wire w_dff_A_gL8JFqHC1_0;
	wire w_dff_A_mn71MHuM9_0;
	wire w_dff_A_F5iUrl6o0_0;
	wire w_dff_A_EkrmMm8i8_0;
	wire w_dff_A_vMimOC1k9_0;
	wire w_dff_A_KL0o4pkr0_0;
	wire w_dff_A_BD31Yy7l0_0;
	wire w_dff_A_qpCYztlw5_2;
	wire w_dff_B_Kjj8zeKW6_3;
	wire w_dff_A_03eJseTV7_1;
	wire w_dff_A_RFfJsU3L2_0;
	wire w_dff_A_NmQBxOPY0_0;
	wire w_dff_A_DvTUDHWg5_0;
	wire w_dff_A_DZ3kNWmy3_0;
	wire w_dff_A_bBe5pjPZ5_0;
	wire w_dff_A_0HeKcJ4V4_0;
	wire w_dff_A_aPPxyjUa3_0;
	wire w_dff_A_RaAq9WJD3_0;
	wire w_dff_A_JThiMuv48_0;
	wire w_dff_A_hp8YCXT01_0;
	wire w_dff_A_o068Pd0r7_0;
	wire w_dff_A_dwW8yMJR4_0;
	wire w_dff_A_fBT6QHjD8_0;
	wire w_dff_A_r6ZIXBe10_0;
	wire w_dff_A_RQkaPbBk4_0;
	wire w_dff_A_ZoSmQTxH3_0;
	wire w_dff_A_VCVnypZW6_0;
	wire w_dff_A_8Bo9Hc4X8_0;
	wire w_dff_A_uUoghMSM2_0;
	wire w_dff_A_qjS0guJK4_0;
	wire w_dff_A_Z6StphLR2_0;
	wire w_dff_A_FUBdNWPA0_0;
	wire w_dff_A_kJRBKz5K4_0;
	wire w_dff_A_ZkCocvNM8_0;
	wire w_dff_A_JB0yltDU4_0;
	wire w_dff_A_Hih7WZBh5_0;
	wire w_dff_A_z6WDJsky7_0;
	wire w_dff_A_r0EMzGvt8_0;
	wire w_dff_A_oHVSIxFd0_0;
	wire w_dff_A_vMm4ViDN6_0;
	wire w_dff_A_vHkAoap27_0;
	wire w_dff_A_yqD3fYIL6_0;
	wire w_dff_A_LlRkeM6N6_0;
	wire w_dff_A_AiDsZfnE9_0;
	wire w_dff_A_4cC0n8LY6_0;
	wire w_dff_A_J8lUbPxx5_0;
	wire w_dff_B_6gfZuDbi7_1;
	wire w_dff_A_9eFwGtyh4_0;
	wire w_dff_A_hdwgpgnO3_0;
	wire w_dff_A_596yo6Vi2_0;
	wire w_dff_A_j4x7Z8LB3_0;
	wire w_dff_A_VQFfDJ7K8_0;
	wire w_dff_A_mAbMNXvs3_0;
	wire w_dff_A_TmJVRVwT5_0;
	wire w_dff_A_Ja1R6rpZ0_0;
	wire w_dff_A_nszDdtmS8_0;
	wire w_dff_A_XL1cAoy86_0;
	wire w_dff_A_PivG70kI5_0;
	wire w_dff_A_jSIN758f0_0;
	wire w_dff_A_PLIYJFqk0_1;
	wire w_dff_A_48NzCRVX1_1;
	wire w_dff_A_4eB1vzSh6_1;
	wire w_dff_A_lJ9so47W8_1;
	wire w_dff_A_2Ij2tSQU3_1;
	wire w_dff_A_dnWcQex08_1;
	wire w_dff_A_Iux8xokn0_1;
	wire w_dff_A_Xa1wW3WC9_1;
	wire w_dff_A_Ma8atjKv5_1;
	wire w_dff_A_oVoRhqSM1_1;
	wire w_dff_A_SsHMTVMO1_1;
	wire w_dff_A_OabsjFqx3_1;
	wire w_dff_A_ew04d99e6_2;
	wire w_dff_A_LRvXUAPF7_0;
	wire w_dff_A_P4TUrj3J0_1;
	wire w_dff_A_VFoEQOwg3_1;
	wire w_dff_A_zb5LOJgW4_1;
	wire w_dff_A_7wRUYp1D7_1;
	wire w_dff_A_FpzwSYq85_1;
	wire w_dff_A_2ozmdymg6_1;
	wire w_dff_A_bunV11Jf6_1;
	wire w_dff_A_vMUNhKiV5_1;
	wire w_dff_A_GjTl6uMF1_1;
	wire w_dff_A_WV88DE9N7_1;
	wire w_dff_A_VLLucF106_1;
	wire w_dff_A_kQaYuDZR3_1;
	wire w_dff_A_KXZGKMQm0_1;
	wire w_dff_A_HWVpkStF9_0;
	wire w_dff_A_lEJQRov87_0;
	wire w_dff_A_GpyikO766_0;
	wire w_dff_A_r1sFdeFC2_0;
	wire w_dff_A_8GxpfENN9_0;
	wire w_dff_A_NMVIQQEQ4_0;
	wire w_dff_A_81lGVsSg0_0;
	wire w_dff_A_zV6syvDI7_0;
	wire w_dff_A_b4A1Gu0B7_0;
	wire w_dff_A_RIbDXy913_0;
	wire w_dff_A_4w2dD41U6_0;
	wire w_dff_A_UxdBwvIm7_0;
	wire w_dff_A_e4gkRgac2_0;
	wire w_dff_A_0kABJPeN4_0;
	wire w_dff_A_fPyMpqqX8_0;
	wire w_dff_A_xssdjAiS9_0;
	wire w_dff_A_r7vOCYgc2_0;
	wire w_dff_A_lH6Tg2A75_0;
	wire w_dff_A_IE0wfjbX8_0;
	wire w_dff_A_AFQ64MTR9_0;
	wire w_dff_A_gyiGt1BC9_0;
	wire w_dff_A_VALhBbBd9_0;
	wire w_dff_A_YExgF0Dl7_0;
	wire w_dff_A_dxOoY1ou1_2;
	wire w_dff_A_Sb2aoAom9_2;
	wire w_dff_B_CjQz1sfH8_3;
	wire w_dff_A_t8lApJZ77_0;
	wire w_dff_A_xWUoS5Qy4_0;
	wire w_dff_A_GO0x0GVu1_0;
	wire w_dff_A_MlhHHKkS4_0;
	wire w_dff_A_et69PjZh9_0;
	wire w_dff_A_LEhKMlEW4_0;
	wire w_dff_A_yfkd2Jae4_0;
	wire w_dff_A_GHHk1Mfc7_0;
	wire w_dff_A_hGHzXt5B3_0;
	wire w_dff_A_ZNmJ56nX8_0;
	wire w_dff_A_WTVSMNBA4_0;
	wire w_dff_A_3yL4B5kd1_0;
	wire w_dff_A_ORIxZwkf0_2;
	wire w_dff_A_ycqjFhlk7_0;
	wire w_dff_A_MpiUFeaL3_0;
	wire w_dff_A_pOjbguua1_0;
	wire w_dff_A_tXrCSyVW4_0;
	wire w_dff_A_dHWsy6DF0_0;
	wire w_dff_A_VI5jphLn7_0;
	wire w_dff_A_bKM2r4hu9_2;
	wire w_dff_A_WV8ToBqA8_0;
	wire w_dff_A_fmigtWPK1_0;
	wire w_dff_A_SSNbB8xX0_0;
	wire w_dff_A_MgTCBivD9_0;
	wire w_dff_A_DqRhxA1J7_0;
	wire w_dff_A_jKIa7hMH7_0;
	wire w_dff_A_V5YicqZf1_2;
	wire w_dff_A_eRsXNH8k3_0;
	wire w_dff_A_QagbEwuI0_0;
	wire w_dff_A_nUuyKVi23_0;
	wire w_dff_A_Pq1YFTcR4_0;
	wire w_dff_A_WfsOKEuB5_0;
	wire w_dff_A_mzd5uUs53_0;
	wire w_dff_A_Z87hynQv1_2;
	wire w_dff_A_LPJYAfXf5_0;
	wire w_dff_A_3AWSMHqz1_0;
	wire w_dff_A_OSD9DhOH8_0;
	wire w_dff_A_dDXVwRUp2_0;
	wire w_dff_A_XUJijzqz7_0;
	wire w_dff_A_u5TTwT6p4_0;
	wire w_dff_A_FSygimdF5_2;
	wire w_dff_A_QDNmg8Tt6_0;
	wire w_dff_A_A6W6S7Mx7_0;
	wire w_dff_A_PMweFv0y1_0;
	wire w_dff_A_HhOoxF5I6_0;
	wire w_dff_A_Spf1me6F2_0;
	wire w_dff_A_BW4y78P94_0;
	wire w_dff_A_RZoms0eR5_2;
	wire w_dff_A_YZJptP9c8_0;
	wire w_dff_A_lVVxvWyr1_0;
	wire w_dff_A_7sneRSUN9_0;
	wire w_dff_A_vVhtA5lP9_0;
	wire w_dff_A_T9bLOFgY9_0;
	wire w_dff_A_CcrjtClQ3_0;
	wire w_dff_A_NQySwvJu6_2;
	wire w_dff_A_p55143YZ7_0;
	wire w_dff_A_IDYeaL2B4_0;
	wire w_dff_A_7dEOFYhG3_0;
	wire w_dff_A_H9lozehi6_0;
	wire w_dff_A_mQYWtEAA9_0;
	wire w_dff_A_bcjyiXsn8_0;
	wire w_dff_A_TQOLLgwC9_2;
	wire w_dff_A_pmEkwUVb2_0;
	wire w_dff_A_9aFBBIwN7_0;
	wire w_dff_A_POutuJXy3_0;
	wire w_dff_A_M7NiAXy27_0;
	wire w_dff_A_9FGCjAMl1_0;
	wire w_dff_A_3iU71VsT9_0;
	wire w_dff_A_5Ycg22Kv1_2;
	wire w_dff_A_qIqGPx9B2_0;
	wire w_dff_A_AXvst8434_0;
	wire w_dff_A_ZGdw4PWF5_0;
	wire w_dff_A_YI3b27bo9_0;
	wire w_dff_A_vcZyp59v1_0;
	wire w_dff_A_mwCnbsbj3_0;
	wire w_dff_A_lzIT8M3g4_2;
	wire w_dff_A_rfh8kOMA4_0;
	wire w_dff_A_CYnUaVIB6_0;
	wire w_dff_A_7Pa96jhw6_0;
	wire w_dff_A_sEGMMIQM9_0;
	wire w_dff_A_VHQRqxOg6_0;
	wire w_dff_A_Sj71KOIq9_0;
	wire w_dff_A_uvUXLcwz5_2;
	wire w_dff_A_iRljTdW81_0;
	wire w_dff_A_JxUgbM0U2_0;
	wire w_dff_A_Z5XN34oW7_0;
	wire w_dff_A_io1Mu50u3_0;
	wire w_dff_A_4YK3SS4q2_0;
	wire w_dff_A_LLu33uYp7_0;
	wire w_dff_A_P2cnVXRN3_2;
	wire w_dff_A_XxmygrCQ4_0;
	wire w_dff_A_q5q0f57m1_0;
	wire w_dff_A_nbWLKJ4h0_0;
	wire w_dff_A_hbjlsx3U7_0;
	wire w_dff_A_BmdcwmAi6_0;
	wire w_dff_A_9UcKii0l6_0;
	wire w_dff_A_AZ2yvGcJ3_2;
	wire w_dff_A_vAuxRXTY8_0;
	wire w_dff_A_FBZA62DK0_0;
	wire w_dff_A_5VW6dXCi3_0;
	wire w_dff_A_lMWWcJgq9_0;
	wire w_dff_A_KBalGWIV8_0;
	wire w_dff_A_RuziirYU4_0;
	wire w_dff_A_h1KbCkLi7_2;
	wire w_dff_A_csfwnwYU8_0;
	wire w_dff_A_IAoeHS3R0_0;
	wire w_dff_A_dyyzbw0S6_0;
	wire w_dff_A_4lSJi6Dc8_0;
	wire w_dff_A_nKg3xQLb8_0;
	wire w_dff_A_6Jvh7HyU0_0;
	wire w_dff_A_FiQj09nF1_2;
	wire w_dff_A_jdMXLw3G7_0;
	wire w_dff_A_ig4vAVge4_0;
	wire w_dff_A_yJtbTHFj1_0;
	wire w_dff_A_1zMHCGuL5_0;
	wire w_dff_A_bORZuoLS6_0;
	wire w_dff_A_6BPlr4yS6_0;
	wire w_dff_A_WA84vgUW7_2;
	wire w_dff_A_jPhWAmZk1_0;
	wire w_dff_A_XPGCH2QZ1_0;
	wire w_dff_A_pGX9e0om2_0;
	wire w_dff_A_Wti0b0ev4_0;
	wire w_dff_A_UMJhHJEx7_0;
	wire w_dff_A_YNLFgSwq3_0;
	wire w_dff_A_sQC4fYt42_2;
	wire w_dff_A_V1e0H1oc8_2;
	wire w_dff_A_uG0hByNW5_2;
	wire w_dff_A_2ICqsIVK0_0;
	jnot g000(.din(w_G146_0[2]),.dout(n58),.clk(gclk));
	jxor g001(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n59),.clk(gclk));
	jxor g002(.dina(w_n59_0[1]),.dinb(n58),.dout(n60),.clk(gclk));
	jnot g003(.din(w_G953_1[2]),.dout(n61),.clk(gclk));
	jand g004(.dina(w_n61_3[2]),.dinb(w_G234_0[2]),.dout(n62),.clk(gclk));
	jand g005(.dina(w_n62_0[1]),.dinb(w_G221_0[1]),.dout(n63),.clk(gclk));
	jxor g006(.dina(n63),.dinb(w_G137_0[2]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_G128_1[1]),.dinb(w_G119_0[2]),.dout(n65),.clk(gclk));
	jxor g008(.dina(w_dff_B_BelyrYIz1_0),.dinb(n64),.dout(n66),.clk(gclk));
	jxor g009(.dina(n66),.dinb(w_G110_1[1]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_n67_0[1]),.dinb(w_n60_0[2]),.dout(n68),.clk(gclk));
	jor g011(.dina(w_n68_0[1]),.dinb(w_G902_3[2]),.dout(n69),.clk(gclk));
	jnot g012(.din(w_G902_3[1]),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_3[1]),.dinb(w_G234_0[1]),.dout(n71),.clk(gclk));
	jnot g014(.din(w_n71_0[1]),.dout(n72),.clk(gclk));
	jand g015(.dina(n72),.dinb(w_G217_0[2]),.dout(n73),.clk(gclk));
	jxor g016(.dina(w_n73_0[1]),.dinb(n69),.dout(n74),.clk(gclk));
	jnot g017(.din(w_G134_0[2]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_G137_0[1]),.dinb(n75),.dout(n76),.clk(gclk));
	jnot g019(.din(w_G131_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_G146_0[1]),.dinb(w_G143_1[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(n78),.dinb(w_G128_1[0]),.dout(n79),.clk(gclk));
	jxor g022(.dina(w_n79_0[1]),.dinb(w_n77_0[1]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_dff_B_6gfZuDbi7_1),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[1]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(w_n82_0[1]),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_1[1]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[2]),.dinb(w_n70_3[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(n91),.dinb(w_G472_0[1]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[2]),.dinb(w_n74_1[1]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[0]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_0[2]),.dout(n96),.clk(gclk));
	jand g039(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n97),.clk(gclk));
	jnot g040(.din(w_G110_1[0]),.dout(n98),.clk(gclk));
	jxor g041(.dina(w_G122_1[1]),.dinb(n98),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n100),.clk(gclk));
	jxor g043(.dina(n100),.dinb(w_G101_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_n101_0[1]),.dinb(w_n84_0[0]),.dout(n102),.clk(gclk));
	jxor g045(.dina(n102),.dinb(w_dff_B_dnr6vzjO6_1),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n61_3[1]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n79_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(w_dff_B_FO9vK7AP2_1),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n103_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[2]),.dinb(w_n70_2[2]),.dout(n108),.clk(gclk));
	jxor g051(.dina(w_n108_0[1]),.dinb(w_n97_0[1]),.dout(n109),.clk(gclk));
	jand g052(.dina(w_n109_0[1]),.dinb(w_n96_0[2]),.dout(n110),.clk(gclk));
	jnot g053(.din(w_G221_0[0]),.dout(n111),.clk(gclk));
	jor g054(.dina(w_n71_0[0]),.dinb(w_dff_B_rah6lkTt0_1),.dout(n112),.clk(gclk));
	jxor g055(.dina(w_G140_0[1]),.dinb(w_G110_0[2]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n61_3[0]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(n114),.dinb(w_n101_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(w_dff_B_eXj6DoYl4_1),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n81_0[1]),.dout(n117),.clk(gclk));
	jand g060(.dina(w_n117_0[2]),.dinb(w_n70_2[1]),.dout(n118),.clk(gclk));
	jxor g061(.dina(w_n118_0[1]),.dinb(w_G469_0[2]),.dout(n119),.clk(gclk));
	jand g062(.dina(w_n119_0[1]),.dinb(w_n112_1[1]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n110_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_1[1]),.dinb(w_n93_0[2]),.dout(n122),.clk(gclk));
	jnot g065(.din(w_G478_0[2]),.dout(n123),.clk(gclk));
	jxor g066(.dina(w_G143_1[0]),.dinb(w_G128_0[2]),.dout(n124),.clk(gclk));
	jand g067(.dina(w_n62_0[0]),.dinb(w_G217_0[1]),.dout(n125),.clk(gclk));
	jxor g068(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n126),.clk(gclk));
	jxor g069(.dina(w_G134_0[1]),.dinb(w_G107_0[1]),.dout(n127),.clk(gclk));
	jxor g070(.dina(n127),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g071(.dina(w_dff_B_fzf9OgLb8_0),.dinb(n125),.dout(n129),.clk(gclk));
	jxor g072(.dina(n129),.dinb(w_dff_B_IEDcSjra0_1),.dout(n130),.clk(gclk));
	jand g073(.dina(w_n130_0[2]),.dinb(w_n70_2[0]),.dout(n131),.clk(gclk));
	jxor g074(.dina(w_n131_0[1]),.dinb(w_dff_B_c9ZLC9CU5_1),.dout(n132),.clk(gclk));
	jnot g075(.din(w_G475_0[2]),.dout(n133),.clk(gclk));
	jxor g076(.dina(w_G143_0[2]),.dinb(w_n77_0[0]),.dout(n134),.clk(gclk));
	jxor g077(.dina(w_G122_0[2]),.dinb(w_n82_0[0]),.dout(n135),.clk(gclk));
	jxor g078(.dina(n135),.dinb(w_G104_0[1]),.dout(n136),.clk(gclk));
	jnot g079(.din(w_G214_0[0]),.dout(n137),.clk(gclk));
	jor g080(.dina(w_n86_0[0]),.dinb(n137),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(w_n60_0[1]),.dout(n139),.clk(gclk));
	jxor g082(.dina(n139),.dinb(n136),.dout(n140),.clk(gclk));
	jxor g083(.dina(n140),.dinb(w_dff_B_L8QKAwC11_1),.dout(n141),.clk(gclk));
	jand g084(.dina(w_n141_0[2]),.dinb(w_n70_1[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_n142_0[1]),.dinb(w_dff_B_0iPv6gzG1_1),.dout(n143),.clk(gclk));
	jand g086(.dina(w_n143_1[1]),.dinb(w_n132_0[2]),.dout(n144),.clk(gclk));
	jor g087(.dina(w_n61_2[2]),.dinb(w_dff_B_7Y2DWtMV5_1),.dout(n145),.clk(gclk));
	jand g088(.dina(w_G237_0[0]),.dinb(w_G234_0[0]),.dout(n146),.clk(gclk));
	jor g089(.dina(w_n146_0[1]),.dinb(w_n70_1[1]),.dout(n147),.clk(gclk));
	jor g090(.dina(w_n147_0[1]),.dinb(w_n145_0[1]),.dout(n148),.clk(gclk));
	jnot g091(.din(w_n146_0[0]),.dout(n149),.clk(gclk));
	jand g092(.dina(w_n61_2[1]),.dinb(w_G952_0[2]),.dout(n150),.clk(gclk));
	jand g093(.dina(n150),.dinb(n149),.dout(n151),.clk(gclk));
	jnot g094(.din(w_n151_0[2]),.dout(n152),.clk(gclk));
	jand g095(.dina(w_n152_0[1]),.dinb(w_dff_B_1zEFzQYj5_1),.dout(n153),.clk(gclk));
	jnot g096(.din(w_n153_0[2]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n144_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[2]),.dinb(w_n122_0[1]),.dout(n156),.clk(gclk));
	jxor g099(.dina(w_n156_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_ORIxZwkf0_2),.clk(gclk));
	jnot g100(.din(w_n92_1[1]),.dout(n158),.clk(gclk));
	jand g101(.dina(w_n158_1[1]),.dinb(w_n74_1[0]),.dout(n159),.clk(gclk));
	jand g102(.dina(w_n159_1[1]),.dinb(w_n121_1[0]),.dout(n160),.clk(gclk));
	jxor g103(.dina(w_n142_0[0]),.dinb(w_G475_0[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_0[2]),.dinb(w_n132_0[1]),.dout(n162),.clk(gclk));
	jand g105(.dina(w_n162_0[1]),.dinb(w_n154_1[0]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_0[2]),.dinb(w_n160_0[1]),.dout(n164),.clk(gclk));
	jxor g107(.dina(w_n164_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_bKM2r4hu9_2),.clk(gclk));
	jxor g108(.dina(w_n131_0[0]),.dinb(w_G478_0[1]),.dout(n166),.clk(gclk));
	jand g109(.dina(w_n143_1[0]),.dinb(w_n166_1[1]),.dout(n167),.clk(gclk));
	jand g110(.dina(w_n167_0[1]),.dinb(w_n154_0[2]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n168_0[2]),.dinb(w_n160_0[0]),.dout(n169),.clk(gclk));
	jxor g112(.dina(w_n169_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_V5YicqZf1_2),.clk(gclk));
	jnot g113(.din(w_n60_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n67_0[0]),.dinb(w_dff_B_MBQeGfwG0_1),.dout(n172),.clk(gclk));
	jand g115(.dina(w_n172_0[1]),.dinb(w_n70_1[0]),.dout(n173),.clk(gclk));
	jxor g116(.dina(w_n73_0[0]),.dinb(n173),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n158_1[0]),.dinb(w_n174_1[1]),.dout(n175),.clk(gclk));
	jand g118(.dina(w_n175_0[1]),.dinb(w_n155_0[1]),.dout(n176),.clk(gclk));
	jand g119(.dina(n176),.dinb(w_n121_0[2]),.dout(n177),.clk(gclk));
	jxor g120(.dina(w_n177_0[1]),.dinb(w_G110_0[1]),.dout(w_dff_A_Z87hynQv1_2),.clk(gclk));
	jand g121(.dina(w_n92_1[0]),.dinb(w_n174_1[0]),.dout(n179),.clk(gclk));
	jand g122(.dina(w_n179_0[2]),.dinb(w_n121_0[1]),.dout(n180),.clk(gclk));
	jor g123(.dina(w_n61_2[0]),.dinb(w_dff_B_vaIuTYF12_1),.dout(n181),.clk(gclk));
	jor g124(.dina(w_n181_0[2]),.dinb(w_n147_0[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(w_dff_B_CKUBDPhr6_0),.dinb(w_n152_0[0]),.dout(n183),.clk(gclk));
	jnot g126(.din(w_n183_0[2]),.dout(n184),.clk(gclk));
	jand g127(.dina(w_n184_1[1]),.dinb(w_n167_0[0]),.dout(n185),.clk(gclk));
	jand g128(.dina(w_n185_0[2]),.dinb(w_n180_0[1]),.dout(n186),.clk(gclk));
	jxor g129(.dina(w_n186_0[1]),.dinb(w_G128_0[1]),.dout(w_dff_A_FSygimdF5_2),.clk(gclk));
	jand g130(.dina(w_n161_0[1]),.dinb(w_n166_1[0]),.dout(n188),.clk(gclk));
	jand g131(.dina(w_n188_0[2]),.dinb(w_n184_1[0]),.dout(n189),.clk(gclk));
	jand g132(.dina(w_n189_0[1]),.dinb(w_n122_0[0]),.dout(n190),.clk(gclk));
	jxor g133(.dina(w_n190_0[1]),.dinb(w_G143_0[1]),.dout(w_dff_A_RZoms0eR5_2),.clk(gclk));
	jand g134(.dina(w_n184_0[2]),.dinb(w_n162_0[0]),.dout(n192),.clk(gclk));
	jand g135(.dina(w_n192_0[2]),.dinb(w_n180_0[0]),.dout(n193),.clk(gclk));
	jxor g136(.dina(w_n193_0[1]),.dinb(w_G146_0[0]),.dout(w_dff_A_NQySwvJu6_2),.clk(gclk));
	jnot g137(.din(w_G469_0[1]),.dout(n195),.clk(gclk));
	jxor g138(.dina(w_n118_0[0]),.dinb(w_dff_B_IDrOGnTz9_1),.dout(n196),.clk(gclk));
	jand g139(.dina(w_n196_0[2]),.dinb(w_n112_1[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n110_0[1]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_1[1]),.dinb(w_n93_0[1]),.dout(n199),.clk(gclk));
	jand g142(.dina(w_n199_0[1]),.dinb(w_n163_0[1]),.dout(n200),.clk(gclk));
	jxor g143(.dina(w_n200_0[1]),.dinb(w_G113_0[0]),.dout(w_dff_A_TQOLLgwC9_2),.clk(gclk));
	jand g144(.dina(w_n199_0[0]),.dinb(w_n168_0[1]),.dout(n202),.clk(gclk));
	jxor g145(.dina(w_n202_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_5Ycg22Kv1_2),.clk(gclk));
	jand g146(.dina(w_n198_1[0]),.dinb(w_n179_0[1]),.dout(n204),.clk(gclk));
	jand g147(.dina(n204),.dinb(w_n155_0[0]),.dout(n205),.clk(gclk));
	jxor g148(.dina(w_n205_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_lzIT8M3g4_2),.clk(gclk));
	jand g149(.dina(w_n197_1[0]),.dinb(w_n159_1[0]),.dout(n207),.clk(gclk));
	jand g150(.dina(w_n154_0[1]),.dinb(w_n110_0[0]),.dout(n208),.clk(gclk));
	jand g151(.dina(n208),.dinb(w_n188_0[1]),.dout(n209),.clk(gclk));
	jand g152(.dina(w_dff_B_KIiYPtj29_0),.dinb(w_n207_0[1]),.dout(n210),.clk(gclk));
	jxor g153(.dina(w_n210_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_uvUXLcwz5_2),.clk(gclk));
	jand g154(.dina(w_n192_0[1]),.dinb(w_n175_0[0]),.dout(n212),.clk(gclk));
	jand g155(.dina(w_n212_0[1]),.dinb(w_n198_0[2]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_n213_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_P2cnVXRN3_2),.clk(gclk));
	jnot g157(.din(w_n97_0[0]),.dout(n215),.clk(gclk));
	jxor g158(.dina(w_n108_0[0]),.dinb(w_dff_B_kUSsOW6B4_1),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_0[2]),.dinb(w_n96_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[2]),.dinb(w_n120_0[0]),.dout(n218),.clk(gclk));
	jand g161(.dina(w_n218_1[1]),.dinb(w_n93_0[0]),.dout(n219),.clk(gclk));
	jand g162(.dina(w_n219_0[1]),.dinb(w_n192_0[0]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_AZ2yvGcJ3_2),.clk(gclk));
	jand g164(.dina(w_n219_0[0]),.dinb(w_n185_0[1]),.dout(n222),.clk(gclk));
	jxor g165(.dina(w_n222_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_h1KbCkLi7_2),.clk(gclk));
	jand g166(.dina(w_n184_0[1]),.dinb(w_n144_1[1]),.dout(n224),.clk(gclk));
	jand g167(.dina(w_dff_B_XkZapgF37_0),.dinb(w_n179_0[0]),.dout(n225),.clk(gclk));
	jand g168(.dina(n225),.dinb(w_n218_1[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_FiQj09nF1_2),.clk(gclk));
	jand g170(.dina(w_n218_0[2]),.dinb(w_n212_0[0]),.dout(n228),.clk(gclk));
	jxor g171(.dina(w_n228_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_WA84vgUW7_2),.clk(gclk));
	jor g172(.dina(w_n177_0[0]),.dinb(w_n169_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n202_0[0]),.dinb(w_n164_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(n230),.dout(n232),.clk(gclk));
	jor g175(.dina(w_n205_0[0]),.dinb(w_n156_0[0]),.dout(n233),.clk(gclk));
	jor g176(.dina(w_n210_0[0]),.dinb(w_n200_0[0]),.dout(n234),.clk(gclk));
	jor g177(.dina(n234),.dinb(n233),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(n232),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n193_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n222_0[0]),.dinb(w_n186_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jor g182(.dina(w_n228_0[0]),.dinb(w_n190_0[0]),.dout(n240),.clk(gclk));
	jor g183(.dina(w_n226_0[0]),.dinb(w_n213_0[0]),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n240),.dout(n242),.clk(gclk));
	jor g185(.dina(n242),.dinb(n239),.dout(n243),.clk(gclk));
	jor g186(.dina(n243),.dinb(n236),.dout(n244),.clk(gclk));
	jor g187(.dina(w_n218_0[1]),.dinb(w_n198_0[1]),.dout(n245),.clk(gclk));
	jand g188(.dina(n245),.dinb(w_n144_1[0]),.dout(n246),.clk(gclk));
	jand g189(.dina(w_n217_0[1]),.dinb(w_n197_0[2]),.dout(n247),.clk(gclk));
	jxor g190(.dina(w_n143_0[2]),.dinb(w_n132_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(w_dff_B_NQnUtYsK0_0),.dinb(n247),.dout(n249),.clk(gclk));
	jor g192(.dina(w_dff_B_HchSND1N3_0),.dinb(n246),.dout(n250),.clk(gclk));
	jand g193(.dina(n250),.dinb(w_n159_0[2]),.dout(n251),.clk(gclk));
	jand g194(.dina(w_n217_0[0]),.dinb(w_n144_0[2]),.dout(n252),.clk(gclk));
	jor g195(.dina(w_n92_0[2]),.dinb(w_n174_0[2]),.dout(n253),.clk(gclk));
	jor g196(.dina(w_n158_0[2]),.dinb(w_n74_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(w_n197_0[1]),.dinb(w_n254_1[1]),.dout(n255),.clk(gclk));
	jand g198(.dina(n255),.dinb(w_n253_0[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_n252_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(n257),.dinb(n251),.dout(n258),.clk(gclk));
	jand g201(.dina(n258),.dinb(w_n151_0[1]),.dout(n259),.clk(gclk));
	jxor g202(.dina(w_n112_0[2]),.dinb(w_n96_0[0]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n151_0[0]),.dout(n261),.clk(gclk));
	jand g204(.dina(w_dff_B_oeV6Bnr73_0),.dinb(w_n196_0[1]),.dout(n262),.clk(gclk));
	jand g205(.dina(n262),.dinb(w_n216_0[1]),.dout(n263),.clk(gclk));
	jand g206(.dina(w_n159_0[1]),.dinb(w_n144_0[1]),.dout(n264),.clk(gclk));
	jand g207(.dina(n264),.dinb(w_dff_B_RRIAtJGU4_1),.dout(n265),.clk(gclk));
	jor g208(.dina(w_dff_B_NXzlyw5l3_0),.dinb(n259),.dout(n266),.clk(gclk));
	jor g209(.dina(n266),.dinb(w_n244_2[2]),.dout(n267),.clk(gclk));
	jand g210(.dina(n267),.dinb(w_G952_0[1]),.dout(n268),.clk(gclk));
	jand g211(.dina(w_n252_0[0]),.dinb(w_n207_0[0]),.dout(n269),.clk(gclk));
	jor g212(.dina(n269),.dinb(w_G953_1[0]),.dout(n270),.clk(gclk));
	jor g213(.dina(w_dff_B_RmygajzI7_0),.dinb(n268),.dout(w_dff_A_sQC4fYt42_2),.clk(gclk));
	jnot g214(.din(w_n107_0[1]),.dout(n272),.clk(gclk));
	jor g215(.dina(w_n216_0[0]),.dinb(w_n95_0[1]),.dout(n273),.clk(gclk));
	jnot g216(.din(w_n112_0[1]),.dout(n274),.clk(gclk));
	jor g217(.dina(w_n196_0[0]),.dinb(w_n274_0[1]),.dout(n275),.clk(gclk));
	jor g218(.dina(w_n275_0[1]),.dinb(w_n273_0[2]),.dout(n276),.clk(gclk));
	jor g219(.dina(w_n253_0[1]),.dinb(w_n276_1[1]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n168_0[0]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n278_0[1]),.dinb(w_n277_0[1]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n161_0[0]),.dinb(w_n166_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n153_0[1]),.dinb(w_n280_0[1]),.dout(n281),.clk(gclk));
	jor g224(.dina(w_n92_0[1]),.dinb(w_n74_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_0[1]),.dinb(w_n281_0[2]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n276_1[0]),.dout(n284),.clk(gclk));
	jand g227(.dina(n284),.dinb(n279),.dout(n285),.clk(gclk));
	jnot g228(.din(w_n163_0[0]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n277_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n158_0[1]),.dinb(w_n174_0[1]),.dout(n288),.clk(gclk));
	jor g231(.dina(w_n119_0[0]),.dinb(w_n274_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(w_n289_0[1]),.dinb(w_n273_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n290_0[2]),.dinb(w_n288_0[2]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n291_0[1]),.dinb(w_n278_0[0]),.dout(n292),.clk(gclk));
	jand g235(.dina(n292),.dinb(n287),.dout(n293),.clk(gclk));
	jand g236(.dina(n293),.dinb(n285),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n276_0[2]),.dinb(w_n288_0[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n281_0[1]),.dinb(w_n295_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(w_n290_0[1]),.dinb(w_n254_1[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(n297),.dinb(w_n281_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n296),.dout(n299),.clk(gclk));
	jor g242(.dina(w_n291_0[0]),.dinb(w_n286_0[0]),.dout(n300),.clk(gclk));
	jor g243(.dina(w_n289_0[0]),.dinb(w_n253_0[0]),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n188_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n153_0[0]),.dinb(w_n273_0[0]),.dout(n303),.clk(gclk));
	jor g246(.dina(n303),.dinb(n302),.dout(n304),.clk(gclk));
	jor g247(.dina(w_dff_B_PSFF9oYg4_0),.dinb(n301),.dout(n305),.clk(gclk));
	jand g248(.dina(n305),.dinb(n300),.dout(n306),.clk(gclk));
	jand g249(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jand g250(.dina(n307),.dinb(n294),.dout(n308),.clk(gclk));
	jor g251(.dina(w_n254_0[2]),.dinb(w_n276_0[1]),.dout(n309),.clk(gclk));
	jor g252(.dina(w_n143_0[1]),.dinb(w_n166_0[1]),.dout(n310),.clk(gclk));
	jor g253(.dina(w_n183_0[1]),.dinb(n310),.dout(n311),.clk(gclk));
	jor g254(.dina(w_n311_0[2]),.dinb(w_n309_0[1]),.dout(n312),.clk(gclk));
	jor g255(.dina(w_n109_0[0]),.dinb(w_n95_0[0]),.dout(n313),.clk(gclk));
	jor g256(.dina(n313),.dinb(w_n275_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n314_0[2]),.dinb(w_n288_0[0]),.dout(n315),.clk(gclk));
	jor g258(.dina(w_n315_0[1]),.dinb(w_n311_0[1]),.dout(n316),.clk(gclk));
	jand g259(.dina(n316),.dinb(n312),.dout(n317),.clk(gclk));
	jnot g260(.din(w_n185_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(w_n318_0[1]),.dinb(w_n309_0[0]),.dout(n319),.clk(gclk));
	jor g262(.dina(w_n315_0[0]),.dinb(w_n318_0[0]),.dout(n320),.clk(gclk));
	jand g263(.dina(n320),.dinb(n319),.dout(n321),.clk(gclk));
	jand g264(.dina(n321),.dinb(n317),.dout(n322),.clk(gclk));
	jnot g265(.din(w_n189_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(w_dff_B_Z1qjeC8T8_0),.dinb(w_n295_0[0]),.dout(n324),.clk(gclk));
	jor g267(.dina(w_n311_0[0]),.dinb(w_n282_0[0]),.dout(n325),.clk(gclk));
	jor g268(.dina(w_n314_0[1]),.dinb(w_n325_0[1]),.dout(n326),.clk(gclk));
	jand g269(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n325_0[0]),.dinb(w_n290_0[0]),.dout(n328),.clk(gclk));
	jor g271(.dina(w_n183_0[0]),.dinb(w_n280_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(w_dff_B_48Z0yb8N8_0),.dinb(w_n254_0[1]),.dout(n330),.clk(gclk));
	jor g273(.dina(n330),.dinb(w_n314_0[0]),.dout(n331),.clk(gclk));
	jand g274(.dina(n331),.dinb(n328),.dout(n332),.clk(gclk));
	jand g275(.dina(n332),.dinb(n327),.dout(n333),.clk(gclk));
	jand g276(.dina(n333),.dinb(n322),.dout(n334),.clk(gclk));
	jand g277(.dina(w_n334_0[1]),.dinb(w_n308_0[1]),.dout(n335),.clk(gclk));
	jand g278(.dina(w_G902_2[2]),.dinb(w_G210_0[0]),.dout(n336),.clk(gclk));
	jnot g279(.din(w_n336_0[1]),.dout(n337),.clk(gclk));
	jor g280(.dina(w_dff_B_tCazLvko6_0),.dinb(w_n335_2[1]),.dout(n338),.clk(gclk));
	jor g281(.dina(n338),.dinb(w_dff_B_gnaP1tmM2_1),.dout(n339),.clk(gclk));
	jor g282(.dina(w_n61_1[2]),.dinb(w_G952_0[0]),.dout(n340),.clk(gclk));
	jand g283(.dina(w_n336_0[0]),.dinb(w_n244_2[1]),.dout(n341),.clk(gclk));
	jor g284(.dina(n341),.dinb(w_n107_0[0]),.dout(n342),.clk(gclk));
	jand g285(.dina(n342),.dinb(w_n340_2[1]),.dout(n343),.clk(gclk));
	jand g286(.dina(n343),.dinb(w_dff_B_2rVMevCL3_1),.dout(G51),.clk(gclk));
	jnot g287(.din(w_n117_0[1]),.dout(n345),.clk(gclk));
	jand g288(.dina(w_G902_2[1]),.dinb(w_G469_0[0]),.dout(n346),.clk(gclk));
	jnot g289(.din(w_n346_0[1]),.dout(n347),.clk(gclk));
	jor g290(.dina(w_dff_B_xtRc2aEM8_0),.dinb(w_n335_2[0]),.dout(n348),.clk(gclk));
	jor g291(.dina(n348),.dinb(w_dff_B_kPV2oe9U6_1),.dout(n349),.clk(gclk));
	jand g292(.dina(w_n346_0[0]),.dinb(w_n244_2[0]),.dout(n350),.clk(gclk));
	jor g293(.dina(n350),.dinb(w_n117_0[0]),.dout(n351),.clk(gclk));
	jand g294(.dina(n351),.dinb(w_n340_2[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_dff_B_EMJWFZeT6_1),.dout(G54),.clk(gclk));
	jnot g296(.din(w_n141_0[1]),.dout(n354),.clk(gclk));
	jand g297(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n355),.clk(gclk));
	jnot g298(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jor g299(.dina(w_dff_B_CDFvh2JA5_0),.dinb(w_n335_1[2]),.dout(n357),.clk(gclk));
	jor g300(.dina(n357),.dinb(w_dff_B_YbF1Pfnz5_1),.dout(n358),.clk(gclk));
	jand g301(.dina(w_n355_0[0]),.dinb(w_n244_1[2]),.dout(n359),.clk(gclk));
	jor g302(.dina(n359),.dinb(w_n141_0[0]),.dout(n360),.clk(gclk));
	jand g303(.dina(n360),.dinb(w_n340_1[2]),.dout(n361),.clk(gclk));
	jand g304(.dina(n361),.dinb(w_dff_B_FJJWjWYM7_1),.dout(G60),.clk(gclk));
	jnot g305(.din(w_n130_0[1]),.dout(n363),.clk(gclk));
	jand g306(.dina(w_G902_1[2]),.dinb(w_G478_0[0]),.dout(n364),.clk(gclk));
	jnot g307(.din(w_n364_0[1]),.dout(n365),.clk(gclk));
	jor g308(.dina(w_dff_B_QxbYTAa80_0),.dinb(w_n335_1[1]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(w_dff_B_uNXQ2yTB4_1),.dout(n367),.clk(gclk));
	jand g310(.dina(w_n364_0[0]),.dinb(w_n244_1[1]),.dout(n368),.clk(gclk));
	jor g311(.dina(n368),.dinb(w_n130_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(n369),.dinb(w_n340_1[1]),.dout(n370),.clk(gclk));
	jand g313(.dina(n370),.dinb(w_dff_B_kb1An8e37_1),.dout(G63),.clk(gclk));
	jand g314(.dina(w_G902_1[1]),.dinb(w_G217_0[0]),.dout(n372),.clk(gclk));
	jand g315(.dina(w_n372_0[1]),.dinb(w_n244_1[0]),.dout(n373),.clk(gclk));
	jor g316(.dina(n373),.dinb(w_n172_0[0]),.dout(n374),.clk(gclk));
	jnot g317(.din(w_n372_0[0]),.dout(n375),.clk(gclk));
	jor g318(.dina(w_dff_B_r9UUnYqn5_0),.dinb(w_n335_1[0]),.dout(n376),.clk(gclk));
	jor g319(.dina(n376),.dinb(w_n68_0[0]),.dout(n377),.clk(gclk));
	jand g320(.dina(n377),.dinb(w_n340_1[0]),.dout(n378),.clk(gclk));
	jand g321(.dina(n378),.dinb(w_dff_B_3rFXgPFh9_1),.dout(G66),.clk(gclk));
	jnot g322(.din(w_n145_0[0]),.dout(n380),.clk(gclk));
	jor g323(.dina(w_n308_0[0]),.dinb(w_G953_0[2]),.dout(n381),.clk(gclk));
	jor g324(.dina(w_n61_1[1]),.dinb(w_G224_0[0]),.dout(n382),.clk(gclk));
	jand g325(.dina(w_dff_B_L3uD0Hyc4_0),.dinb(n381),.dout(n383),.clk(gclk));
	jxor g326(.dina(n383),.dinb(w_n103_0[0]),.dout(n384),.clk(gclk));
	jor g327(.dina(n384),.dinb(w_dff_B_xmqYbzs75_1),.dout(w_dff_A_V1e0H1oc8_2),.clk(gclk));
	jor g328(.dina(w_n334_0[0]),.dinb(w_G953_0[1]),.dout(n386),.clk(gclk));
	jor g329(.dina(w_n61_1[0]),.dinb(w_G227_0[0]),.dout(n387),.clk(gclk));
	jand g330(.dina(n387),.dinb(w_n181_0[1]),.dout(n388),.clk(gclk));
	jand g331(.dina(w_dff_B_3QYbYrbm0_0),.dinb(n386),.dout(n389),.clk(gclk));
	jnot g332(.din(w_n181_0[0]),.dout(n390),.clk(gclk));
	jxor g333(.dina(w_n81_0[0]),.dinb(w_n59_0[0]),.dout(n391),.clk(gclk));
	jor g334(.dina(n391),.dinb(w_dff_B_8j7wOmlc8_1),.dout(n392),.clk(gclk));
	jxor g335(.dina(w_dff_B_Wxwyns1d6_0),.dinb(n389),.dout(w_dff_A_uG0hByNW5_2),.clk(gclk));
	jnot g336(.din(w_n90_0[1]),.dout(n394),.clk(gclk));
	jand g337(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n395),.clk(gclk));
	jnot g338(.din(w_n395_0[1]),.dout(n396),.clk(gclk));
	jor g339(.dina(w_dff_B_cXxrWteb3_0),.dinb(w_n335_0[2]),.dout(n397),.clk(gclk));
	jor g340(.dina(n397),.dinb(w_dff_B_MRxDTQWd2_1),.dout(n398),.clk(gclk));
	jand g341(.dina(w_n395_0[0]),.dinb(w_n244_0[2]),.dout(n399),.clk(gclk));
	jor g342(.dina(n399),.dinb(w_n90_0[0]),.dout(n400),.clk(gclk));
	jand g343(.dina(n400),.dinb(w_n340_0[2]),.dout(n401),.clk(gclk));
	jand g344(.dina(n401),.dinb(w_dff_B_FlWjvmng7_1),.dout(G57),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_BD31Yy7l0_0),.doutb(w_G101_0[1]),.doutc(w_dff_A_qpCYztlw5_2),.din(w_dff_B_Kjj8zeKW6_3));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_JUN6cAtx4_0),.doutb(w_dff_A_L3g0NJor4_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_II0a2sMc3_0),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_G110_0[0]),.doutb(w_dff_A_DssgHyMX5_1),.doutc(w_G110_0[2]),.din(G110));
	jspl jspl_w_G110_1(.douta(w_G110_1[0]),.doutb(w_dff_A_aclXEIyw0_1),.din(w_G110_0[0]));
	jspl jspl_w_G113_0(.douta(w_dff_A_J8lUbPxx5_0),.doutb(w_G113_0[1]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_ZkCocvNM8_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_dwW8yMJR4_0),.doutb(w_G119_0[1]),.doutc(w_G119_0[2]),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_w6arXA8v7_1),.doutc(w_dff_A_Ec8Ld3O35_2),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_dff_A_Ddh5DIGQ4_1),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_ZQxUeYFV5_0),.doutb(w_dff_A_nAprNfw33_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_dff_A_kQaYuDZR3_1),.doutc(w_G128_0[2]),.din(G128));
	jspl jspl_w_G128_1(.douta(w_dff_A_LRvXUAPF7_0),.doutb(w_G128_1[1]),.din(w_G128_0[0]));
	jspl jspl_w_G131_0(.douta(w_dff_A_UxdBwvIm7_0),.doutb(w_G131_0[1]),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_3yL4B5kd1_0),.doutb(w_G134_0[1]),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_YExgF0Dl7_0),.doutb(w_G137_0[1]),.doutc(w_dff_A_Sb2aoAom9_2),.din(w_dff_B_CjQz1sfH8_3));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_YVDvWf2Z5_0),.doutb(w_G140_0[1]),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_dff_A_OabsjFqx3_1),.doutc(w_dff_A_ew04d99e6_2),.din(G143));
	jspl jspl_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.din(w_G143_0[0]));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_jSIN758f0_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(G146));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_dff_A_o71ohj0b8_1),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_dff_A_WHE8BckL9_1),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_G217_0[0]),.doutb(w_dff_A_zl8609TL1_1),.doutc(w_dff_A_0FYkV1dJ2_2),.din(G217));
	jspl jspl_w_G221_0(.douta(w_G221_0[0]),.doutb(w_dff_A_yCpBk0Y09_1),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_G224_0[1]),.din(w_dff_B_Cs8bBDdu8_2));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_G227_0[1]),.din(w_dff_B_cFSZjj0a2_2));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_dff_A_ggVshsIh6_1),.doutc(w_dff_A_89kZRE0r3_2),.din(G234));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_G469_0[0]),.doutb(w_G469_0[1]),.doutc(w_dff_A_kUKg9n2E9_2),.din(G469));
	jspl jspl_w_G472_0(.douta(w_G472_0[0]),.doutb(w_dff_A_j5LbCEsr0_1),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_OxoHZ5Ps2_1),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_G478_0[0]),.doutb(w_dff_A_HidJcISd9_1),.doutc(w_G478_0[2]),.din(G478));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_G902_1[1]),.doutc(w_G902_1[2]),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_G902_2[1]),.doutc(w_G902_2[2]),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_G902_3[0]),.doutb(w_G902_3[1]),.doutc(w_dff_A_QRdg40aF4_2),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_dff_A_tcPEUmQq8_1),.doutc(w_G952_0[2]),.din(w_dff_B_23RAqRpQ9_3));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_dff_A_v8bqlD7a2_1),.doutc(w_dff_A_5XAaL6JI8_2),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_N8483xR91_0),.doutb(w_G953_1[1]),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_n59_0(.douta(w_dff_A_NRjXV6Yh0_0),.doutb(w_n59_0[1]),.din(n59));
	jspl3 jspl3_w_n60_0(.douta(w_n60_0[0]),.doutb(w_n60_0[1]),.doutc(w_dff_A_honyHz3o2_2),.din(n60));
	jspl3 jspl3_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.doutc(w_n61_0[2]),.din(n61));
	jspl3 jspl3_w_n61_1(.douta(w_n61_1[0]),.doutb(w_n61_1[1]),.doutc(w_n61_1[2]),.din(w_n61_0[0]));
	jspl3 jspl3_w_n61_2(.douta(w_n61_2[0]),.doutb(w_n61_2[1]),.doutc(w_n61_2[2]),.din(w_n61_0[1]));
	jspl3 jspl3_w_n61_3(.douta(w_n61_3[0]),.doutb(w_n61_3[1]),.doutc(w_n61_3[2]),.din(w_n61_0[2]));
	jspl jspl_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n68_0(.douta(w_dff_A_TCZ09ifv2_0),.doutb(w_n68_0[1]),.din(n68));
	jspl3 jspl3_w_n70_0(.douta(w_n70_0[0]),.doutb(w_dff_A_t4wq9cUJ4_1),.doutc(w_n70_0[2]),.din(n70));
	jspl3 jspl3_w_n70_1(.douta(w_dff_A_PyS38Hry9_0),.doutb(w_n70_1[1]),.doutc(w_dff_A_zWlwC2Ou2_2),.din(w_n70_0[0]));
	jspl3 jspl3_w_n70_2(.douta(w_n70_2[0]),.doutb(w_n70_2[1]),.doutc(w_n70_2[2]),.din(w_n70_0[1]));
	jspl jspl_w_n70_3(.douta(w_dff_A_60j5QT485_0),.doutb(w_n70_3[1]),.din(w_n70_0[2]));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(w_dff_B_AJ4NIPbd6_2));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_dff_A_KXZGKMQm0_1),.din(n77));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl jspl_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_03eJseTV7_1),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n90_0(.douta(w_dff_A_MCYmCCnC0_0),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_dff_A_6LwPzpr78_1),.doutc(w_dff_A_j7Zy7O2B8_2),.din(n92));
	jspl3 jspl3_w_n92_1(.douta(w_dff_A_mNchYbv10_0),.doutb(w_n92_1[1]),.doutc(w_dff_A_uma05frZ8_2),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_dff_A_pp7OSwDu3_0),.doutb(w_dff_A_5I2AiDSb2_1),.doutc(w_n95_0[2]),.din(n95));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_l9XTGDeg8_1),.doutc(w_dff_A_fHH7YDY19_2),.din(n96));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_dff_A_VhmM6P478_1),.din(n97));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_dff_A_wN0Zf4xK3_0),.doutb(w_n103_0[1]),.din(n103));
	jspl3 jspl3_w_n107_0(.douta(w_dff_A_g1ORjDxT3_0),.doutb(w_n107_0[1]),.doutc(w_n107_0[2]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.doutc(w_n110_0[2]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_QhbAil4O7_0),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_dff_A_VzVx22lW7_0),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_dff_A_GnX2E4J12_2),.din(w_dff_B_m8neVkhE9_3));
	jspl jspl_w_n121_1(.douta(w_n121_1[0]),.doutb(w_n121_1[1]),.din(w_n121_0[0]));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_VM9zdHHW2_0),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n141_0(.douta(w_dff_A_rGr1XINl7_0),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl jspl_w_n143_1(.douta(w_n143_1[0]),.doutb(w_n143_1[1]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_dff_A_k8eG48ky1_1),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_dff_A_LS0OlbDu1_0),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl3 jspl3_w_n151_0(.douta(w_dff_A_hupSypvR0_0),.doutb(w_dff_A_IbXovPq23_1),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_dff_A_7y0MB23R2_0),.doutb(w_dff_A_rICxkPtJ8_1),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(w_dff_B_TII2KWyq0_3));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_dff_A_pkz4VgKi7_0),.doutb(w_n155_0[1]),.doutc(w_dff_A_U7V0YSX17_2),.din(w_dff_B_MkLyWnOY7_3));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.doutc(w_n158_0[2]),.din(w_dff_B_owlxZTpc5_3));
	jspl jspl_w_n158_1(.douta(w_n158_1[0]),.doutb(w_n158_1[1]),.din(w_n158_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_dff_A_xZt7LRzF2_2),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_dff_A_LI1M4O6h8_1),.doutc(w_dff_A_RUEtXAqY8_2),.din(n163));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl jspl_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.din(w_n166_0[0]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_dff_A_GoMmkFZB3_1),.doutc(w_dff_A_5TdxSzju1_2),.din(n168));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n172_0(.douta(w_dff_A_i59WwYfY7_0),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.doutc(w_n174_0[2]),.din(n174));
	jspl jspl_w_n174_1(.douta(w_n174_1[0]),.doutb(w_n174_1[1]),.din(w_n174_0[0]));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.doutc(w_n179_0[2]),.din(n179));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n183_0(.douta(w_dff_A_724vyw0z0_0),.doutb(w_dff_A_QPbox9xq7_1),.doutc(w_n183_0[2]),.din(n183));
	jspl3 jspl3_w_n184_0(.douta(w_n184_0[0]),.doutb(w_n184_0[1]),.doutc(w_n184_0[2]),.din(w_dff_B_pOEkBLmB1_3));
	jspl jspl_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_dff_A_PmJZcSWs4_1),.doutc(w_dff_A_Mzvb4cNp0_2),.din(n185));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl3 jspl3_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_jiVXwrw15_1),.doutc(w_n188_0[2]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_dff_A_TmET4rrF7_1),.din(n189));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_dff_A_hGQAbzib8_0),.doutb(w_n192_0[1]),.doutc(w_dff_A_j8MwRq0V6_2),.din(w_dff_B_irItOaNe5_3));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl3 jspl3_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(n196));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_dff_A_hsnnmuCv1_1),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_dff_A_SkE9QDgu5_0),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_dff_A_FQT5dyl84_0),.doutb(w_n198_0[1]),.doutc(w_dff_A_Hafs6tmu3_2),.din(n198));
	jspl jspl_w_n198_1(.douta(w_n198_1[0]),.doutb(w_n198_1[1]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_dff_A_sv65aGNS4_1),.doutc(w_n216_0[2]),.din(n216));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl3 jspl3_w_n218_0(.douta(w_dff_A_vH4ZGHON8_0),.doutb(w_n218_0[1]),.doutc(w_dff_A_M7YcBVR91_2),.din(n218));
	jspl jspl_w_n218_1(.douta(w_dff_A_qOvmg9cl6_0),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl3 jspl3_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.doutc(w_n244_0[2]),.din(n244));
	jspl3 jspl3_w_n244_1(.douta(w_n244_1[0]),.doutb(w_n244_1[1]),.doutc(w_n244_1[2]),.din(w_n244_0[0]));
	jspl3 jspl3_w_n244_2(.douta(w_n244_2[0]),.doutb(w_n244_2[1]),.doutc(w_n244_2[2]),.din(w_n244_0[1]));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_w1LRiMgX4_1),.din(w_dff_B_oE9QYs901_2));
	jspl3 jspl3_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.doutc(w_dff_A_9iLFHuQA5_2),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_IxfoKFtQ6_2));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_n276_0[2]),.din(w_dff_B_Noibk2AT2_3));
	jspl jspl_w_n276_1(.douta(w_dff_A_aK5RmE8l4_0),.doutb(w_n276_1[1]),.din(w_n276_0[0]));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(w_dff_B_bdT2QtA68_2));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n281_0(.douta(w_dff_A_IrqCsY0U8_0),.doutb(w_dff_A_juWZbGN95_1),.doutc(w_n281_0[2]),.din(w_dff_B_bEywQSYi2_3));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(w_dff_B_rjIpW8xh5_2));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n289_0(.douta(w_dff_A_FlTTx5ZE9_0),.doutb(w_n289_0[1]),.din(n289));
	jspl3 jspl3_w_n290_0(.douta(w_dff_A_DPVzRc6d1_0),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(w_dff_B_TEqAAgl68_3));
	jspl jspl_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.din(n291));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_dff_A_B1jwbQ744_1),.doutc(w_dff_A_VmapFO1s6_2),.din(w_dff_B_raYUAsUH5_3));
	jspl3 jspl3_w_n314_0(.douta(w_dff_A_zxpVdtJC4_0),.doutb(w_dff_A_S0gXY9FI0_1),.doutc(w_n314_0[2]),.din(w_dff_B_NvAM7Nba6_3));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(w_dff_B_DjmXnYWK5_2));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.doutc(w_n335_1[2]),.din(w_n335_0[0]));
	jspl jspl_w_n335_2(.douta(w_n335_2[0]),.doutb(w_n335_2[1]),.din(w_n335_0[1]));
	jspl jspl_w_n336_0(.douta(w_dff_A_tnTHw7G86_0),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.doutc(w_n340_0[2]),.din(w_dff_B_zDweCeiP0_3));
	jspl3 jspl3_w_n340_1(.douta(w_n340_1[0]),.doutb(w_n340_1[1]),.doutc(w_n340_1[2]),.din(w_n340_0[0]));
	jspl jspl_w_n340_2(.douta(w_n340_2[0]),.doutb(w_n340_2[1]),.din(w_n340_0[1]));
	jspl jspl_w_n346_0(.douta(w_dff_A_qFbPGn452_0),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n355_0(.douta(w_dff_A_BaKcvWCA8_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n364_0(.douta(w_dff_A_bYMbuxKl5_0),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_D8Wqng4N3_1),.din(n372));
	jspl jspl_w_n395_0(.douta(w_dff_A_j9yRjunC8_0),.doutb(w_n395_0[1]),.din(n395));
	jdff dff_B_87bOp2Dn6_0(.din(n270),.dout(w_dff_B_87bOp2Dn6_0),.clk(gclk));
	jdff dff_B_7EPSNGhf3_0(.din(w_dff_B_87bOp2Dn6_0),.dout(w_dff_B_7EPSNGhf3_0),.clk(gclk));
	jdff dff_B_n8utcfpF5_0(.din(w_dff_B_7EPSNGhf3_0),.dout(w_dff_B_n8utcfpF5_0),.clk(gclk));
	jdff dff_B_UPSYHjBa0_0(.din(w_dff_B_n8utcfpF5_0),.dout(w_dff_B_UPSYHjBa0_0),.clk(gclk));
	jdff dff_B_RmygajzI7_0(.din(w_dff_B_UPSYHjBa0_0),.dout(w_dff_B_RmygajzI7_0),.clk(gclk));
	jdff dff_B_xfuKnVey6_0(.din(n265),.dout(w_dff_B_xfuKnVey6_0),.clk(gclk));
	jdff dff_B_WqfXkezP9_0(.din(w_dff_B_xfuKnVey6_0),.dout(w_dff_B_WqfXkezP9_0),.clk(gclk));
	jdff dff_B_NXzlyw5l3_0(.din(w_dff_B_WqfXkezP9_0),.dout(w_dff_B_NXzlyw5l3_0),.clk(gclk));
	jdff dff_B_efvta5zN5_1(.din(n263),.dout(w_dff_B_efvta5zN5_1),.clk(gclk));
	jdff dff_B_RRIAtJGU4_1(.din(w_dff_B_efvta5zN5_1),.dout(w_dff_B_RRIAtJGU4_1),.clk(gclk));
	jdff dff_B_SCWmaTYi6_0(.din(n261),.dout(w_dff_B_SCWmaTYi6_0),.clk(gclk));
	jdff dff_B_oeV6Bnr73_0(.din(w_dff_B_SCWmaTYi6_0),.dout(w_dff_B_oeV6Bnr73_0),.clk(gclk));
	jdff dff_A_w1LRiMgX4_1(.dout(w_n252_0[1]),.din(w_dff_A_w1LRiMgX4_1),.clk(gclk));
	jdff dff_B_ffzbGroE8_2(.din(n252),.dout(w_dff_B_ffzbGroE8_2),.clk(gclk));
	jdff dff_B_oE9QYs901_2(.din(w_dff_B_ffzbGroE8_2),.dout(w_dff_B_oE9QYs901_2),.clk(gclk));
	jdff dff_B_HchSND1N3_0(.din(n249),.dout(w_dff_B_HchSND1N3_0),.clk(gclk));
	jdff dff_B_NQnUtYsK0_0(.din(n248),.dout(w_dff_B_NQnUtYsK0_0),.clk(gclk));
	jdff dff_B_2rVMevCL3_1(.din(n339),.dout(w_dff_B_2rVMevCL3_1),.clk(gclk));
	jdff dff_B_JrWMiEAL9_1(.din(n272),.dout(w_dff_B_JrWMiEAL9_1),.clk(gclk));
	jdff dff_B_CdeKqlzU0_1(.din(w_dff_B_JrWMiEAL9_1),.dout(w_dff_B_CdeKqlzU0_1),.clk(gclk));
	jdff dff_B_6UeguRop8_1(.din(w_dff_B_CdeKqlzU0_1),.dout(w_dff_B_6UeguRop8_1),.clk(gclk));
	jdff dff_B_gbDAL4yQ9_1(.din(w_dff_B_6UeguRop8_1),.dout(w_dff_B_gbDAL4yQ9_1),.clk(gclk));
	jdff dff_B_8YIKaS3Q4_1(.din(w_dff_B_gbDAL4yQ9_1),.dout(w_dff_B_8YIKaS3Q4_1),.clk(gclk));
	jdff dff_B_Ltn759w28_1(.din(w_dff_B_8YIKaS3Q4_1),.dout(w_dff_B_Ltn759w28_1),.clk(gclk));
	jdff dff_B_5MO2mbjK0_1(.din(w_dff_B_Ltn759w28_1),.dout(w_dff_B_5MO2mbjK0_1),.clk(gclk));
	jdff dff_B_mRxGlBQw8_1(.din(w_dff_B_5MO2mbjK0_1),.dout(w_dff_B_mRxGlBQw8_1),.clk(gclk));
	jdff dff_B_0EoOZv3n9_1(.din(w_dff_B_mRxGlBQw8_1),.dout(w_dff_B_0EoOZv3n9_1),.clk(gclk));
	jdff dff_B_jtQwMBmn6_1(.din(w_dff_B_0EoOZv3n9_1),.dout(w_dff_B_jtQwMBmn6_1),.clk(gclk));
	jdff dff_B_gnaP1tmM2_1(.din(w_dff_B_jtQwMBmn6_1),.dout(w_dff_B_gnaP1tmM2_1),.clk(gclk));
	jdff dff_B_6nTKUK5i8_0(.din(n337),.dout(w_dff_B_6nTKUK5i8_0),.clk(gclk));
	jdff dff_B_3XEJPL3B0_0(.din(w_dff_B_6nTKUK5i8_0),.dout(w_dff_B_3XEJPL3B0_0),.clk(gclk));
	jdff dff_B_ZQxSm2Hy8_0(.din(w_dff_B_3XEJPL3B0_0),.dout(w_dff_B_ZQxSm2Hy8_0),.clk(gclk));
	jdff dff_B_TgTPCfoI8_0(.din(w_dff_B_ZQxSm2Hy8_0),.dout(w_dff_B_TgTPCfoI8_0),.clk(gclk));
	jdff dff_B_yaPhb7sG4_0(.din(w_dff_B_TgTPCfoI8_0),.dout(w_dff_B_yaPhb7sG4_0),.clk(gclk));
	jdff dff_B_QQY9Zqxy4_0(.din(w_dff_B_yaPhb7sG4_0),.dout(w_dff_B_QQY9Zqxy4_0),.clk(gclk));
	jdff dff_B_MQqHOlKA4_0(.din(w_dff_B_QQY9Zqxy4_0),.dout(w_dff_B_MQqHOlKA4_0),.clk(gclk));
	jdff dff_B_TEzwHQ728_0(.din(w_dff_B_MQqHOlKA4_0),.dout(w_dff_B_TEzwHQ728_0),.clk(gclk));
	jdff dff_B_Bwi442li8_0(.din(w_dff_B_TEzwHQ728_0),.dout(w_dff_B_Bwi442li8_0),.clk(gclk));
	jdff dff_B_PrAKKe2k3_0(.din(w_dff_B_Bwi442li8_0),.dout(w_dff_B_PrAKKe2k3_0),.clk(gclk));
	jdff dff_B_s46XYIaT3_0(.din(w_dff_B_PrAKKe2k3_0),.dout(w_dff_B_s46XYIaT3_0),.clk(gclk));
	jdff dff_B_QGb7rWg47_0(.din(w_dff_B_s46XYIaT3_0),.dout(w_dff_B_QGb7rWg47_0),.clk(gclk));
	jdff dff_B_VRCL3miz9_0(.din(w_dff_B_QGb7rWg47_0),.dout(w_dff_B_VRCL3miz9_0),.clk(gclk));
	jdff dff_B_tCazLvko6_0(.din(w_dff_B_VRCL3miz9_0),.dout(w_dff_B_tCazLvko6_0),.clk(gclk));
	jdff dff_A_PLb05sP82_0(.dout(w_n336_0[0]),.din(w_dff_A_PLb05sP82_0),.clk(gclk));
	jdff dff_A_VwyzMuxh0_0(.dout(w_dff_A_PLb05sP82_0),.din(w_dff_A_VwyzMuxh0_0),.clk(gclk));
	jdff dff_A_AP0J3wpp0_0(.dout(w_dff_A_VwyzMuxh0_0),.din(w_dff_A_AP0J3wpp0_0),.clk(gclk));
	jdff dff_A_VBce0eM76_0(.dout(w_dff_A_AP0J3wpp0_0),.din(w_dff_A_VBce0eM76_0),.clk(gclk));
	jdff dff_A_iL4p3XwZ7_0(.dout(w_dff_A_VBce0eM76_0),.din(w_dff_A_iL4p3XwZ7_0),.clk(gclk));
	jdff dff_A_8B8EmH428_0(.dout(w_dff_A_iL4p3XwZ7_0),.din(w_dff_A_8B8EmH428_0),.clk(gclk));
	jdff dff_A_xZrc1hw80_0(.dout(w_dff_A_8B8EmH428_0),.din(w_dff_A_xZrc1hw80_0),.clk(gclk));
	jdff dff_A_lDlFOIXc2_0(.dout(w_dff_A_xZrc1hw80_0),.din(w_dff_A_lDlFOIXc2_0),.clk(gclk));
	jdff dff_A_da4Fr2co1_0(.dout(w_dff_A_lDlFOIXc2_0),.din(w_dff_A_da4Fr2co1_0),.clk(gclk));
	jdff dff_A_A7DPSFRy2_0(.dout(w_dff_A_da4Fr2co1_0),.din(w_dff_A_A7DPSFRy2_0),.clk(gclk));
	jdff dff_A_VxuOEcPy6_0(.dout(w_dff_A_A7DPSFRy2_0),.din(w_dff_A_VxuOEcPy6_0),.clk(gclk));
	jdff dff_A_eclfmUr33_0(.dout(w_dff_A_VxuOEcPy6_0),.din(w_dff_A_eclfmUr33_0),.clk(gclk));
	jdff dff_A_2CLhYjZW0_0(.dout(w_dff_A_eclfmUr33_0),.din(w_dff_A_2CLhYjZW0_0),.clk(gclk));
	jdff dff_A_k57PodTn7_0(.dout(w_dff_A_2CLhYjZW0_0),.din(w_dff_A_k57PodTn7_0),.clk(gclk));
	jdff dff_A_tnTHw7G86_0(.dout(w_dff_A_k57PodTn7_0),.din(w_dff_A_tnTHw7G86_0),.clk(gclk));
	jdff dff_B_EMJWFZeT6_1(.din(n349),.dout(w_dff_B_EMJWFZeT6_1),.clk(gclk));
	jdff dff_B_0Lm1mm1f4_1(.din(n345),.dout(w_dff_B_0Lm1mm1f4_1),.clk(gclk));
	jdff dff_B_9olJ5uMv3_1(.din(w_dff_B_0Lm1mm1f4_1),.dout(w_dff_B_9olJ5uMv3_1),.clk(gclk));
	jdff dff_B_5B6R03Jt6_1(.din(w_dff_B_9olJ5uMv3_1),.dout(w_dff_B_5B6R03Jt6_1),.clk(gclk));
	jdff dff_B_Gxzs4Bdx9_1(.din(w_dff_B_5B6R03Jt6_1),.dout(w_dff_B_Gxzs4Bdx9_1),.clk(gclk));
	jdff dff_B_sW2URFvA7_1(.din(w_dff_B_Gxzs4Bdx9_1),.dout(w_dff_B_sW2URFvA7_1),.clk(gclk));
	jdff dff_B_ZCuoqVvF1_1(.din(w_dff_B_sW2URFvA7_1),.dout(w_dff_B_ZCuoqVvF1_1),.clk(gclk));
	jdff dff_B_bUGtMhTw1_1(.din(w_dff_B_ZCuoqVvF1_1),.dout(w_dff_B_bUGtMhTw1_1),.clk(gclk));
	jdff dff_B_k14CYDZ95_1(.din(w_dff_B_bUGtMhTw1_1),.dout(w_dff_B_k14CYDZ95_1),.clk(gclk));
	jdff dff_B_dQFnZUCt6_1(.din(w_dff_B_k14CYDZ95_1),.dout(w_dff_B_dQFnZUCt6_1),.clk(gclk));
	jdff dff_B_WgABFuDi2_1(.din(w_dff_B_dQFnZUCt6_1),.dout(w_dff_B_WgABFuDi2_1),.clk(gclk));
	jdff dff_B_kPV2oe9U6_1(.din(w_dff_B_WgABFuDi2_1),.dout(w_dff_B_kPV2oe9U6_1),.clk(gclk));
	jdff dff_B_hS2AizXh1_0(.din(n347),.dout(w_dff_B_hS2AizXh1_0),.clk(gclk));
	jdff dff_B_QDQ36sKV7_0(.din(w_dff_B_hS2AizXh1_0),.dout(w_dff_B_QDQ36sKV7_0),.clk(gclk));
	jdff dff_B_N9jgM4oF5_0(.din(w_dff_B_QDQ36sKV7_0),.dout(w_dff_B_N9jgM4oF5_0),.clk(gclk));
	jdff dff_B_6IOFgYHm9_0(.din(w_dff_B_N9jgM4oF5_0),.dout(w_dff_B_6IOFgYHm9_0),.clk(gclk));
	jdff dff_B_oNTF7GxA0_0(.din(w_dff_B_6IOFgYHm9_0),.dout(w_dff_B_oNTF7GxA0_0),.clk(gclk));
	jdff dff_B_3eb7y8xu1_0(.din(w_dff_B_oNTF7GxA0_0),.dout(w_dff_B_3eb7y8xu1_0),.clk(gclk));
	jdff dff_B_uqEmhBw49_0(.din(w_dff_B_3eb7y8xu1_0),.dout(w_dff_B_uqEmhBw49_0),.clk(gclk));
	jdff dff_B_VYR1kyWC0_0(.din(w_dff_B_uqEmhBw49_0),.dout(w_dff_B_VYR1kyWC0_0),.clk(gclk));
	jdff dff_B_kIhGJ28b7_0(.din(w_dff_B_VYR1kyWC0_0),.dout(w_dff_B_kIhGJ28b7_0),.clk(gclk));
	jdff dff_B_cpqG3vRd2_0(.din(w_dff_B_kIhGJ28b7_0),.dout(w_dff_B_cpqG3vRd2_0),.clk(gclk));
	jdff dff_B_C3wiqR8Y3_0(.din(w_dff_B_cpqG3vRd2_0),.dout(w_dff_B_C3wiqR8Y3_0),.clk(gclk));
	jdff dff_B_LH6297VJ0_0(.din(w_dff_B_C3wiqR8Y3_0),.dout(w_dff_B_LH6297VJ0_0),.clk(gclk));
	jdff dff_B_Flx2KE5N8_0(.din(w_dff_B_LH6297VJ0_0),.dout(w_dff_B_Flx2KE5N8_0),.clk(gclk));
	jdff dff_B_xtRc2aEM8_0(.din(w_dff_B_Flx2KE5N8_0),.dout(w_dff_B_xtRc2aEM8_0),.clk(gclk));
	jdff dff_A_9xGKUnYC8_0(.dout(w_n346_0[0]),.din(w_dff_A_9xGKUnYC8_0),.clk(gclk));
	jdff dff_A_FWOljebP4_0(.dout(w_dff_A_9xGKUnYC8_0),.din(w_dff_A_FWOljebP4_0),.clk(gclk));
	jdff dff_A_kzXMQSPo7_0(.dout(w_dff_A_FWOljebP4_0),.din(w_dff_A_kzXMQSPo7_0),.clk(gclk));
	jdff dff_A_e0SIynSB3_0(.dout(w_dff_A_kzXMQSPo7_0),.din(w_dff_A_e0SIynSB3_0),.clk(gclk));
	jdff dff_A_jzaYJtxw4_0(.dout(w_dff_A_e0SIynSB3_0),.din(w_dff_A_jzaYJtxw4_0),.clk(gclk));
	jdff dff_A_xoj7Wjnk8_0(.dout(w_dff_A_jzaYJtxw4_0),.din(w_dff_A_xoj7Wjnk8_0),.clk(gclk));
	jdff dff_A_rF1peoG50_0(.dout(w_dff_A_xoj7Wjnk8_0),.din(w_dff_A_rF1peoG50_0),.clk(gclk));
	jdff dff_A_WSoTL0gh4_0(.dout(w_dff_A_rF1peoG50_0),.din(w_dff_A_WSoTL0gh4_0),.clk(gclk));
	jdff dff_A_uPBe1R1J3_0(.dout(w_dff_A_WSoTL0gh4_0),.din(w_dff_A_uPBe1R1J3_0),.clk(gclk));
	jdff dff_A_erVE1r2B7_0(.dout(w_dff_A_uPBe1R1J3_0),.din(w_dff_A_erVE1r2B7_0),.clk(gclk));
	jdff dff_A_dE7RRdtE9_0(.dout(w_dff_A_erVE1r2B7_0),.din(w_dff_A_dE7RRdtE9_0),.clk(gclk));
	jdff dff_A_KjJuUzWy9_0(.dout(w_dff_A_dE7RRdtE9_0),.din(w_dff_A_KjJuUzWy9_0),.clk(gclk));
	jdff dff_A_NH0SwtXT7_0(.dout(w_dff_A_KjJuUzWy9_0),.din(w_dff_A_NH0SwtXT7_0),.clk(gclk));
	jdff dff_A_FmyFiHIR5_0(.dout(w_dff_A_NH0SwtXT7_0),.din(w_dff_A_FmyFiHIR5_0),.clk(gclk));
	jdff dff_A_qFbPGn452_0(.dout(w_dff_A_FmyFiHIR5_0),.din(w_dff_A_qFbPGn452_0),.clk(gclk));
	jdff dff_B_FJJWjWYM7_1(.din(n358),.dout(w_dff_B_FJJWjWYM7_1),.clk(gclk));
	jdff dff_B_k8MqHn3t9_1(.din(n354),.dout(w_dff_B_k8MqHn3t9_1),.clk(gclk));
	jdff dff_B_zwnjIeiK8_1(.din(w_dff_B_k8MqHn3t9_1),.dout(w_dff_B_zwnjIeiK8_1),.clk(gclk));
	jdff dff_B_JqS2EPZr7_1(.din(w_dff_B_zwnjIeiK8_1),.dout(w_dff_B_JqS2EPZr7_1),.clk(gclk));
	jdff dff_B_5Yzj6bd25_1(.din(w_dff_B_JqS2EPZr7_1),.dout(w_dff_B_5Yzj6bd25_1),.clk(gclk));
	jdff dff_B_IRVWZmf29_1(.din(w_dff_B_5Yzj6bd25_1),.dout(w_dff_B_IRVWZmf29_1),.clk(gclk));
	jdff dff_B_aHmAifBI7_1(.din(w_dff_B_IRVWZmf29_1),.dout(w_dff_B_aHmAifBI7_1),.clk(gclk));
	jdff dff_B_CXKRjkup3_1(.din(w_dff_B_aHmAifBI7_1),.dout(w_dff_B_CXKRjkup3_1),.clk(gclk));
	jdff dff_B_1XDmuVL00_1(.din(w_dff_B_CXKRjkup3_1),.dout(w_dff_B_1XDmuVL00_1),.clk(gclk));
	jdff dff_B_NXvphe786_1(.din(w_dff_B_1XDmuVL00_1),.dout(w_dff_B_NXvphe786_1),.clk(gclk));
	jdff dff_B_RFLLM3IV4_1(.din(w_dff_B_NXvphe786_1),.dout(w_dff_B_RFLLM3IV4_1),.clk(gclk));
	jdff dff_B_YbF1Pfnz5_1(.din(w_dff_B_RFLLM3IV4_1),.dout(w_dff_B_YbF1Pfnz5_1),.clk(gclk));
	jdff dff_B_vpfRtk9D0_0(.din(n356),.dout(w_dff_B_vpfRtk9D0_0),.clk(gclk));
	jdff dff_B_o0rhkiDo3_0(.din(w_dff_B_vpfRtk9D0_0),.dout(w_dff_B_o0rhkiDo3_0),.clk(gclk));
	jdff dff_B_gwqHUlfu5_0(.din(w_dff_B_o0rhkiDo3_0),.dout(w_dff_B_gwqHUlfu5_0),.clk(gclk));
	jdff dff_B_wCo0NCMB2_0(.din(w_dff_B_gwqHUlfu5_0),.dout(w_dff_B_wCo0NCMB2_0),.clk(gclk));
	jdff dff_B_jie2EpRX0_0(.din(w_dff_B_wCo0NCMB2_0),.dout(w_dff_B_jie2EpRX0_0),.clk(gclk));
	jdff dff_B_dKYklQW12_0(.din(w_dff_B_jie2EpRX0_0),.dout(w_dff_B_dKYklQW12_0),.clk(gclk));
	jdff dff_B_GHXsExDM4_0(.din(w_dff_B_dKYklQW12_0),.dout(w_dff_B_GHXsExDM4_0),.clk(gclk));
	jdff dff_B_lE7cFnSs2_0(.din(w_dff_B_GHXsExDM4_0),.dout(w_dff_B_lE7cFnSs2_0),.clk(gclk));
	jdff dff_B_6kwKJZot7_0(.din(w_dff_B_lE7cFnSs2_0),.dout(w_dff_B_6kwKJZot7_0),.clk(gclk));
	jdff dff_B_8EaBU1Eg0_0(.din(w_dff_B_6kwKJZot7_0),.dout(w_dff_B_8EaBU1Eg0_0),.clk(gclk));
	jdff dff_B_iq1igln77_0(.din(w_dff_B_8EaBU1Eg0_0),.dout(w_dff_B_iq1igln77_0),.clk(gclk));
	jdff dff_B_wTMFt1eP9_0(.din(w_dff_B_iq1igln77_0),.dout(w_dff_B_wTMFt1eP9_0),.clk(gclk));
	jdff dff_B_E3S5Ybt36_0(.din(w_dff_B_wTMFt1eP9_0),.dout(w_dff_B_E3S5Ybt36_0),.clk(gclk));
	jdff dff_B_CDFvh2JA5_0(.din(w_dff_B_E3S5Ybt36_0),.dout(w_dff_B_CDFvh2JA5_0),.clk(gclk));
	jdff dff_A_vLkHJ5s99_0(.dout(w_n355_0[0]),.din(w_dff_A_vLkHJ5s99_0),.clk(gclk));
	jdff dff_A_Wz3c9hGM8_0(.dout(w_dff_A_vLkHJ5s99_0),.din(w_dff_A_Wz3c9hGM8_0),.clk(gclk));
	jdff dff_A_XTYGtVyz8_0(.dout(w_dff_A_Wz3c9hGM8_0),.din(w_dff_A_XTYGtVyz8_0),.clk(gclk));
	jdff dff_A_Rb7KIZkO4_0(.dout(w_dff_A_XTYGtVyz8_0),.din(w_dff_A_Rb7KIZkO4_0),.clk(gclk));
	jdff dff_A_untx1rbH5_0(.dout(w_dff_A_Rb7KIZkO4_0),.din(w_dff_A_untx1rbH5_0),.clk(gclk));
	jdff dff_A_i1BstMmA3_0(.dout(w_dff_A_untx1rbH5_0),.din(w_dff_A_i1BstMmA3_0),.clk(gclk));
	jdff dff_A_P7pfCRud0_0(.dout(w_dff_A_i1BstMmA3_0),.din(w_dff_A_P7pfCRud0_0),.clk(gclk));
	jdff dff_A_yDVYZKAu3_0(.dout(w_dff_A_P7pfCRud0_0),.din(w_dff_A_yDVYZKAu3_0),.clk(gclk));
	jdff dff_A_T8moYjYn7_0(.dout(w_dff_A_yDVYZKAu3_0),.din(w_dff_A_T8moYjYn7_0),.clk(gclk));
	jdff dff_A_10vTaxdQ8_0(.dout(w_dff_A_T8moYjYn7_0),.din(w_dff_A_10vTaxdQ8_0),.clk(gclk));
	jdff dff_A_ETervw5G5_0(.dout(w_dff_A_10vTaxdQ8_0),.din(w_dff_A_ETervw5G5_0),.clk(gclk));
	jdff dff_A_YmfehQHz7_0(.dout(w_dff_A_ETervw5G5_0),.din(w_dff_A_YmfehQHz7_0),.clk(gclk));
	jdff dff_A_D363rGBi5_0(.dout(w_dff_A_YmfehQHz7_0),.din(w_dff_A_D363rGBi5_0),.clk(gclk));
	jdff dff_A_VtVtXx9l5_0(.dout(w_dff_A_D363rGBi5_0),.din(w_dff_A_VtVtXx9l5_0),.clk(gclk));
	jdff dff_A_BaKcvWCA8_0(.dout(w_dff_A_VtVtXx9l5_0),.din(w_dff_A_BaKcvWCA8_0),.clk(gclk));
	jdff dff_B_kb1An8e37_1(.din(n367),.dout(w_dff_B_kb1An8e37_1),.clk(gclk));
	jdff dff_B_hnW3HoZl2_1(.din(n363),.dout(w_dff_B_hnW3HoZl2_1),.clk(gclk));
	jdff dff_B_kuaDvfmG2_1(.din(w_dff_B_hnW3HoZl2_1),.dout(w_dff_B_kuaDvfmG2_1),.clk(gclk));
	jdff dff_B_YmBqXeyF8_1(.din(w_dff_B_kuaDvfmG2_1),.dout(w_dff_B_YmBqXeyF8_1),.clk(gclk));
	jdff dff_B_PHYeC3ry8_1(.din(w_dff_B_YmBqXeyF8_1),.dout(w_dff_B_PHYeC3ry8_1),.clk(gclk));
	jdff dff_B_DlHf5knJ6_1(.din(w_dff_B_PHYeC3ry8_1),.dout(w_dff_B_DlHf5knJ6_1),.clk(gclk));
	jdff dff_B_s6W44nz43_1(.din(w_dff_B_DlHf5knJ6_1),.dout(w_dff_B_s6W44nz43_1),.clk(gclk));
	jdff dff_B_yTE4MABn3_1(.din(w_dff_B_s6W44nz43_1),.dout(w_dff_B_yTE4MABn3_1),.clk(gclk));
	jdff dff_B_dekRpRMT9_1(.din(w_dff_B_yTE4MABn3_1),.dout(w_dff_B_dekRpRMT9_1),.clk(gclk));
	jdff dff_B_EhMBCw9K8_1(.din(w_dff_B_dekRpRMT9_1),.dout(w_dff_B_EhMBCw9K8_1),.clk(gclk));
	jdff dff_B_4uSkO2d68_1(.din(w_dff_B_EhMBCw9K8_1),.dout(w_dff_B_4uSkO2d68_1),.clk(gclk));
	jdff dff_B_uNXQ2yTB4_1(.din(w_dff_B_4uSkO2d68_1),.dout(w_dff_B_uNXQ2yTB4_1),.clk(gclk));
	jdff dff_B_0Hjd63n28_0(.din(n365),.dout(w_dff_B_0Hjd63n28_0),.clk(gclk));
	jdff dff_B_hlq442934_0(.din(w_dff_B_0Hjd63n28_0),.dout(w_dff_B_hlq442934_0),.clk(gclk));
	jdff dff_B_OTEDu9Q83_0(.din(w_dff_B_hlq442934_0),.dout(w_dff_B_OTEDu9Q83_0),.clk(gclk));
	jdff dff_B_EpMVBOMw2_0(.din(w_dff_B_OTEDu9Q83_0),.dout(w_dff_B_EpMVBOMw2_0),.clk(gclk));
	jdff dff_B_79oD9aer7_0(.din(w_dff_B_EpMVBOMw2_0),.dout(w_dff_B_79oD9aer7_0),.clk(gclk));
	jdff dff_B_JGQBD7BZ4_0(.din(w_dff_B_79oD9aer7_0),.dout(w_dff_B_JGQBD7BZ4_0),.clk(gclk));
	jdff dff_B_C12t8k9v5_0(.din(w_dff_B_JGQBD7BZ4_0),.dout(w_dff_B_C12t8k9v5_0),.clk(gclk));
	jdff dff_B_oPsM1g8r3_0(.din(w_dff_B_C12t8k9v5_0),.dout(w_dff_B_oPsM1g8r3_0),.clk(gclk));
	jdff dff_B_qmNqaiHI0_0(.din(w_dff_B_oPsM1g8r3_0),.dout(w_dff_B_qmNqaiHI0_0),.clk(gclk));
	jdff dff_B_WhlBGXK76_0(.din(w_dff_B_qmNqaiHI0_0),.dout(w_dff_B_WhlBGXK76_0),.clk(gclk));
	jdff dff_B_G4UFy2um8_0(.din(w_dff_B_WhlBGXK76_0),.dout(w_dff_B_G4UFy2um8_0),.clk(gclk));
	jdff dff_B_PYidTrXO6_0(.din(w_dff_B_G4UFy2um8_0),.dout(w_dff_B_PYidTrXO6_0),.clk(gclk));
	jdff dff_B_75LSLCq09_0(.din(w_dff_B_PYidTrXO6_0),.dout(w_dff_B_75LSLCq09_0),.clk(gclk));
	jdff dff_B_QxbYTAa80_0(.din(w_dff_B_75LSLCq09_0),.dout(w_dff_B_QxbYTAa80_0),.clk(gclk));
	jdff dff_A_aiSCGz7O5_0(.dout(w_n364_0[0]),.din(w_dff_A_aiSCGz7O5_0),.clk(gclk));
	jdff dff_A_VgYQpamO8_0(.dout(w_dff_A_aiSCGz7O5_0),.din(w_dff_A_VgYQpamO8_0),.clk(gclk));
	jdff dff_A_3FtZ9Gmg3_0(.dout(w_dff_A_VgYQpamO8_0),.din(w_dff_A_3FtZ9Gmg3_0),.clk(gclk));
	jdff dff_A_EtZfJLHb2_0(.dout(w_dff_A_3FtZ9Gmg3_0),.din(w_dff_A_EtZfJLHb2_0),.clk(gclk));
	jdff dff_A_ReleY0UH9_0(.dout(w_dff_A_EtZfJLHb2_0),.din(w_dff_A_ReleY0UH9_0),.clk(gclk));
	jdff dff_A_Mqyqz53w0_0(.dout(w_dff_A_ReleY0UH9_0),.din(w_dff_A_Mqyqz53w0_0),.clk(gclk));
	jdff dff_A_Ilcp6WiR8_0(.dout(w_dff_A_Mqyqz53w0_0),.din(w_dff_A_Ilcp6WiR8_0),.clk(gclk));
	jdff dff_A_nVdmpPMU2_0(.dout(w_dff_A_Ilcp6WiR8_0),.din(w_dff_A_nVdmpPMU2_0),.clk(gclk));
	jdff dff_A_mVvD6MKm1_0(.dout(w_dff_A_nVdmpPMU2_0),.din(w_dff_A_mVvD6MKm1_0),.clk(gclk));
	jdff dff_A_n0hF5aWI9_0(.dout(w_dff_A_mVvD6MKm1_0),.din(w_dff_A_n0hF5aWI9_0),.clk(gclk));
	jdff dff_A_hlbiBiCn7_0(.dout(w_dff_A_n0hF5aWI9_0),.din(w_dff_A_hlbiBiCn7_0),.clk(gclk));
	jdff dff_A_Lbvojlos8_0(.dout(w_dff_A_hlbiBiCn7_0),.din(w_dff_A_Lbvojlos8_0),.clk(gclk));
	jdff dff_A_PpZJM5409_0(.dout(w_dff_A_Lbvojlos8_0),.din(w_dff_A_PpZJM5409_0),.clk(gclk));
	jdff dff_A_cSwTILFg5_0(.dout(w_dff_A_PpZJM5409_0),.din(w_dff_A_cSwTILFg5_0),.clk(gclk));
	jdff dff_A_bYMbuxKl5_0(.dout(w_dff_A_cSwTILFg5_0),.din(w_dff_A_bYMbuxKl5_0),.clk(gclk));
	jdff dff_B_3rFXgPFh9_1(.din(n374),.dout(w_dff_B_3rFXgPFh9_1),.clk(gclk));
	jdff dff_B_0LY0pZrb6_0(.din(n375),.dout(w_dff_B_0LY0pZrb6_0),.clk(gclk));
	jdff dff_B_ROZDpAaR2_0(.din(w_dff_B_0LY0pZrb6_0),.dout(w_dff_B_ROZDpAaR2_0),.clk(gclk));
	jdff dff_B_F01UjAOe8_0(.din(w_dff_B_ROZDpAaR2_0),.dout(w_dff_B_F01UjAOe8_0),.clk(gclk));
	jdff dff_B_ZwaM6reX6_0(.din(w_dff_B_F01UjAOe8_0),.dout(w_dff_B_ZwaM6reX6_0),.clk(gclk));
	jdff dff_B_kXQ6hvyY7_0(.din(w_dff_B_ZwaM6reX6_0),.dout(w_dff_B_kXQ6hvyY7_0),.clk(gclk));
	jdff dff_B_vvTWKtXD0_0(.din(w_dff_B_kXQ6hvyY7_0),.dout(w_dff_B_vvTWKtXD0_0),.clk(gclk));
	jdff dff_B_KbPhcMyl3_0(.din(w_dff_B_vvTWKtXD0_0),.dout(w_dff_B_KbPhcMyl3_0),.clk(gclk));
	jdff dff_B_gwMoCEKh4_0(.din(w_dff_B_KbPhcMyl3_0),.dout(w_dff_B_gwMoCEKh4_0),.clk(gclk));
	jdff dff_B_JJ2FDzwg5_0(.din(w_dff_B_gwMoCEKh4_0),.dout(w_dff_B_JJ2FDzwg5_0),.clk(gclk));
	jdff dff_B_XrPFzcc91_0(.din(w_dff_B_JJ2FDzwg5_0),.dout(w_dff_B_XrPFzcc91_0),.clk(gclk));
	jdff dff_B_QTyRJJdr1_0(.din(w_dff_B_XrPFzcc91_0),.dout(w_dff_B_QTyRJJdr1_0),.clk(gclk));
	jdff dff_B_cPtKHVpI7_0(.din(w_dff_B_QTyRJJdr1_0),.dout(w_dff_B_cPtKHVpI7_0),.clk(gclk));
	jdff dff_B_ZPZysFsS6_0(.din(w_dff_B_cPtKHVpI7_0),.dout(w_dff_B_ZPZysFsS6_0),.clk(gclk));
	jdff dff_B_r9UUnYqn5_0(.din(w_dff_B_ZPZysFsS6_0),.dout(w_dff_B_r9UUnYqn5_0),.clk(gclk));
	jdff dff_A_UlZV1zJ91_1(.dout(w_n372_0[1]),.din(w_dff_A_UlZV1zJ91_1),.clk(gclk));
	jdff dff_A_5WXqnS2S7_1(.dout(w_dff_A_UlZV1zJ91_1),.din(w_dff_A_5WXqnS2S7_1),.clk(gclk));
	jdff dff_A_9mB84Hqz8_1(.dout(w_dff_A_5WXqnS2S7_1),.din(w_dff_A_9mB84Hqz8_1),.clk(gclk));
	jdff dff_A_rp5j1TAM3_1(.dout(w_dff_A_9mB84Hqz8_1),.din(w_dff_A_rp5j1TAM3_1),.clk(gclk));
	jdff dff_A_eDYiX4ky7_1(.dout(w_dff_A_rp5j1TAM3_1),.din(w_dff_A_eDYiX4ky7_1),.clk(gclk));
	jdff dff_A_NNnaF8UE5_1(.dout(w_dff_A_eDYiX4ky7_1),.din(w_dff_A_NNnaF8UE5_1),.clk(gclk));
	jdff dff_A_1VjhMmOB9_1(.dout(w_dff_A_NNnaF8UE5_1),.din(w_dff_A_1VjhMmOB9_1),.clk(gclk));
	jdff dff_A_Yc4LdnPn0_1(.dout(w_dff_A_1VjhMmOB9_1),.din(w_dff_A_Yc4LdnPn0_1),.clk(gclk));
	jdff dff_A_Yzc98HWj1_1(.dout(w_dff_A_Yc4LdnPn0_1),.din(w_dff_A_Yzc98HWj1_1),.clk(gclk));
	jdff dff_A_7xlSI9do8_1(.dout(w_dff_A_Yzc98HWj1_1),.din(w_dff_A_7xlSI9do8_1),.clk(gclk));
	jdff dff_A_6IxUmO6m5_1(.dout(w_dff_A_7xlSI9do8_1),.din(w_dff_A_6IxUmO6m5_1),.clk(gclk));
	jdff dff_A_SmnZ541m5_1(.dout(w_dff_A_6IxUmO6m5_1),.din(w_dff_A_SmnZ541m5_1),.clk(gclk));
	jdff dff_A_7FwV4aLd3_1(.dout(w_dff_A_SmnZ541m5_1),.din(w_dff_A_7FwV4aLd3_1),.clk(gclk));
	jdff dff_A_a1RD86qw0_1(.dout(w_dff_A_7FwV4aLd3_1),.din(w_dff_A_a1RD86qw0_1),.clk(gclk));
	jdff dff_A_D8Wqng4N3_1(.dout(w_dff_A_a1RD86qw0_1),.din(w_dff_A_D8Wqng4N3_1),.clk(gclk));
	jdff dff_B_Dbri4POt1_1(.din(n380),.dout(w_dff_B_Dbri4POt1_1),.clk(gclk));
	jdff dff_B_Q7tqGaGw2_1(.din(w_dff_B_Dbri4POt1_1),.dout(w_dff_B_Q7tqGaGw2_1),.clk(gclk));
	jdff dff_B_xN5SDyhd0_1(.din(w_dff_B_Q7tqGaGw2_1),.dout(w_dff_B_xN5SDyhd0_1),.clk(gclk));
	jdff dff_B_gOpwTTqT0_1(.din(w_dff_B_xN5SDyhd0_1),.dout(w_dff_B_gOpwTTqT0_1),.clk(gclk));
	jdff dff_B_hXY9ravn1_1(.din(w_dff_B_gOpwTTqT0_1),.dout(w_dff_B_hXY9ravn1_1),.clk(gclk));
	jdff dff_B_AmhuZh2S3_1(.din(w_dff_B_hXY9ravn1_1),.dout(w_dff_B_AmhuZh2S3_1),.clk(gclk));
	jdff dff_B_NhPVS65S6_1(.din(w_dff_B_AmhuZh2S3_1),.dout(w_dff_B_NhPVS65S6_1),.clk(gclk));
	jdff dff_B_nhObHOLc5_1(.din(w_dff_B_NhPVS65S6_1),.dout(w_dff_B_nhObHOLc5_1),.clk(gclk));
	jdff dff_B_JvCZmWV14_1(.din(w_dff_B_nhObHOLc5_1),.dout(w_dff_B_JvCZmWV14_1),.clk(gclk));
	jdff dff_B_nHFJlcOV4_1(.din(w_dff_B_JvCZmWV14_1),.dout(w_dff_B_nHFJlcOV4_1),.clk(gclk));
	jdff dff_B_IVn7fjfZ9_1(.din(w_dff_B_nHFJlcOV4_1),.dout(w_dff_B_IVn7fjfZ9_1),.clk(gclk));
	jdff dff_B_I6gRvqVv4_1(.din(w_dff_B_IVn7fjfZ9_1),.dout(w_dff_B_I6gRvqVv4_1),.clk(gclk));
	jdff dff_B_ko09xkuE4_1(.din(w_dff_B_I6gRvqVv4_1),.dout(w_dff_B_ko09xkuE4_1),.clk(gclk));
	jdff dff_B_pBnm7llM9_1(.din(w_dff_B_ko09xkuE4_1),.dout(w_dff_B_pBnm7llM9_1),.clk(gclk));
	jdff dff_B_xmqYbzs75_1(.din(w_dff_B_pBnm7llM9_1),.dout(w_dff_B_xmqYbzs75_1),.clk(gclk));
	jdff dff_B_bNzKWLox1_0(.din(n382),.dout(w_dff_B_bNzKWLox1_0),.clk(gclk));
	jdff dff_B_EbHeg9E11_0(.din(w_dff_B_bNzKWLox1_0),.dout(w_dff_B_EbHeg9E11_0),.clk(gclk));
	jdff dff_B_MATPjOp15_0(.din(w_dff_B_EbHeg9E11_0),.dout(w_dff_B_MATPjOp15_0),.clk(gclk));
	jdff dff_B_nRgoqobJ7_0(.din(w_dff_B_MATPjOp15_0),.dout(w_dff_B_nRgoqobJ7_0),.clk(gclk));
	jdff dff_B_uOBEpA8d6_0(.din(w_dff_B_nRgoqobJ7_0),.dout(w_dff_B_uOBEpA8d6_0),.clk(gclk));
	jdff dff_B_pMFW7uyy6_0(.din(w_dff_B_uOBEpA8d6_0),.dout(w_dff_B_pMFW7uyy6_0),.clk(gclk));
	jdff dff_B_QGtF6uyi2_0(.din(w_dff_B_pMFW7uyy6_0),.dout(w_dff_B_QGtF6uyi2_0),.clk(gclk));
	jdff dff_B_1iYajag89_0(.din(w_dff_B_QGtF6uyi2_0),.dout(w_dff_B_1iYajag89_0),.clk(gclk));
	jdff dff_B_xfUySCc40_0(.din(w_dff_B_1iYajag89_0),.dout(w_dff_B_xfUySCc40_0),.clk(gclk));
	jdff dff_B_Ssv97t0V0_0(.din(w_dff_B_xfUySCc40_0),.dout(w_dff_B_Ssv97t0V0_0),.clk(gclk));
	jdff dff_B_yXH21rMx8_0(.din(w_dff_B_Ssv97t0V0_0),.dout(w_dff_B_yXH21rMx8_0),.clk(gclk));
	jdff dff_B_WCNOHD9j6_0(.din(w_dff_B_yXH21rMx8_0),.dout(w_dff_B_WCNOHD9j6_0),.clk(gclk));
	jdff dff_B_EDuWhzQ47_0(.din(w_dff_B_WCNOHD9j6_0),.dout(w_dff_B_EDuWhzQ47_0),.clk(gclk));
	jdff dff_B_L3uD0Hyc4_0(.din(w_dff_B_EDuWhzQ47_0),.dout(w_dff_B_L3uD0Hyc4_0),.clk(gclk));
	jdff dff_B_FuQFQQAz1_0(.din(n392),.dout(w_dff_B_FuQFQQAz1_0),.clk(gclk));
	jdff dff_B_3BVc73Hu4_0(.din(w_dff_B_FuQFQQAz1_0),.dout(w_dff_B_3BVc73Hu4_0),.clk(gclk));
	jdff dff_B_ls4aoIiI5_0(.din(w_dff_B_3BVc73Hu4_0),.dout(w_dff_B_ls4aoIiI5_0),.clk(gclk));
	jdff dff_B_y831cesS0_0(.din(w_dff_B_ls4aoIiI5_0),.dout(w_dff_B_y831cesS0_0),.clk(gclk));
	jdff dff_B_tK02ByYW3_0(.din(w_dff_B_y831cesS0_0),.dout(w_dff_B_tK02ByYW3_0),.clk(gclk));
	jdff dff_B_cupCJfLT3_0(.din(w_dff_B_tK02ByYW3_0),.dout(w_dff_B_cupCJfLT3_0),.clk(gclk));
	jdff dff_B_XHdNCY1C0_0(.din(w_dff_B_cupCJfLT3_0),.dout(w_dff_B_XHdNCY1C0_0),.clk(gclk));
	jdff dff_B_a43oumxU9_0(.din(w_dff_B_XHdNCY1C0_0),.dout(w_dff_B_a43oumxU9_0),.clk(gclk));
	jdff dff_B_81GGm6a58_0(.din(w_dff_B_a43oumxU9_0),.dout(w_dff_B_81GGm6a58_0),.clk(gclk));
	jdff dff_B_8D8R4uzi7_0(.din(w_dff_B_81GGm6a58_0),.dout(w_dff_B_8D8R4uzi7_0),.clk(gclk));
	jdff dff_B_Wxwyns1d6_0(.din(w_dff_B_8D8R4uzi7_0),.dout(w_dff_B_Wxwyns1d6_0),.clk(gclk));
	jdff dff_B_i2ZLgkmr8_1(.din(n390),.dout(w_dff_B_i2ZLgkmr8_1),.clk(gclk));
	jdff dff_B_8j7wOmlc8_1(.din(w_dff_B_i2ZLgkmr8_1),.dout(w_dff_B_8j7wOmlc8_1),.clk(gclk));
	jdff dff_B_6LORq5xz3_0(.din(n388),.dout(w_dff_B_6LORq5xz3_0),.clk(gclk));
	jdff dff_B_TugF7XTs1_0(.din(w_dff_B_6LORq5xz3_0),.dout(w_dff_B_TugF7XTs1_0),.clk(gclk));
	jdff dff_B_vmoqKux69_0(.din(w_dff_B_TugF7XTs1_0),.dout(w_dff_B_vmoqKux69_0),.clk(gclk));
	jdff dff_B_j9CgkoDt0_0(.din(w_dff_B_vmoqKux69_0),.dout(w_dff_B_j9CgkoDt0_0),.clk(gclk));
	jdff dff_B_cUjSGt0f8_0(.din(w_dff_B_j9CgkoDt0_0),.dout(w_dff_B_cUjSGt0f8_0),.clk(gclk));
	jdff dff_B_6Oq4KqUR5_0(.din(w_dff_B_cUjSGt0f8_0),.dout(w_dff_B_6Oq4KqUR5_0),.clk(gclk));
	jdff dff_B_UuKCp4g08_0(.din(w_dff_B_6Oq4KqUR5_0),.dout(w_dff_B_UuKCp4g08_0),.clk(gclk));
	jdff dff_B_yPMVfwtr6_0(.din(w_dff_B_UuKCp4g08_0),.dout(w_dff_B_yPMVfwtr6_0),.clk(gclk));
	jdff dff_B_3JxjyQcm6_0(.din(w_dff_B_yPMVfwtr6_0),.dout(w_dff_B_3JxjyQcm6_0),.clk(gclk));
	jdff dff_B_9latNVrB7_0(.din(w_dff_B_3JxjyQcm6_0),.dout(w_dff_B_9latNVrB7_0),.clk(gclk));
	jdff dff_B_J81RkvBt1_0(.din(w_dff_B_9latNVrB7_0),.dout(w_dff_B_J81RkvBt1_0),.clk(gclk));
	jdff dff_B_hWJJgJB85_0(.din(w_dff_B_J81RkvBt1_0),.dout(w_dff_B_hWJJgJB85_0),.clk(gclk));
	jdff dff_B_3QYbYrbm0_0(.din(w_dff_B_hWJJgJB85_0),.dout(w_dff_B_3QYbYrbm0_0),.clk(gclk));
	jdff dff_B_FlWjvmng7_1(.din(n398),.dout(w_dff_B_FlWjvmng7_1),.clk(gclk));
	jdff dff_B_XkZapgF37_0(.din(n224),.dout(w_dff_B_XkZapgF37_0),.clk(gclk));
	jdff dff_A_qOvmg9cl6_0(.dout(w_n218_1[0]),.din(w_dff_A_qOvmg9cl6_0),.clk(gclk));
	jdff dff_A_vH4ZGHON8_0(.dout(w_n218_0[0]),.din(w_dff_A_vH4ZGHON8_0),.clk(gclk));
	jdff dff_A_ZagKAg6M8_2(.dout(w_n218_0[2]),.din(w_dff_A_ZagKAg6M8_2),.clk(gclk));
	jdff dff_A_M7YcBVR91_2(.dout(w_dff_A_ZagKAg6M8_2),.din(w_dff_A_M7YcBVR91_2),.clk(gclk));
	jdff dff_A_hGQAbzib8_0(.dout(w_n192_0[0]),.din(w_dff_A_hGQAbzib8_0),.clk(gclk));
	jdff dff_A_j8MwRq0V6_2(.dout(w_n192_0[2]),.din(w_dff_A_j8MwRq0V6_2),.clk(gclk));
	jdff dff_B_irItOaNe5_3(.din(n192),.dout(w_dff_B_irItOaNe5_3),.clk(gclk));
	jdff dff_B_KIiYPtj29_0(.din(n209),.dout(w_dff_B_KIiYPtj29_0),.clk(gclk));
	jdff dff_A_FQT5dyl84_0(.dout(w_n198_0[0]),.din(w_dff_A_FQT5dyl84_0),.clk(gclk));
	jdff dff_A_ZVxorm683_2(.dout(w_n198_0[2]),.din(w_dff_A_ZVxorm683_2),.clk(gclk));
	jdff dff_A_Hafs6tmu3_2(.dout(w_dff_A_ZVxorm683_2),.din(w_dff_A_Hafs6tmu3_2),.clk(gclk));
	jdff dff_A_dBmESVvk1_0(.dout(w_n197_1[0]),.din(w_dff_A_dBmESVvk1_0),.clk(gclk));
	jdff dff_A_SkE9QDgu5_0(.dout(w_dff_A_dBmESVvk1_0),.din(w_dff_A_SkE9QDgu5_0),.clk(gclk));
	jdff dff_A_xphs99ls2_1(.dout(w_n197_0[1]),.din(w_dff_A_xphs99ls2_1),.clk(gclk));
	jdff dff_A_hsnnmuCv1_1(.dout(w_dff_A_xphs99ls2_1),.din(w_dff_A_hsnnmuCv1_1),.clk(gclk));
	jdff dff_A_pkz4VgKi7_0(.dout(w_n155_0[0]),.din(w_dff_A_pkz4VgKi7_0),.clk(gclk));
	jdff dff_A_U7V0YSX17_2(.dout(w_n155_0[2]),.din(w_dff_A_U7V0YSX17_2),.clk(gclk));
	jdff dff_B_MkLyWnOY7_3(.din(n155),.dout(w_dff_B_MkLyWnOY7_3),.clk(gclk));
	jdff dff_A_Z0sc88C71_0(.dout(w_n144_1[0]),.din(w_dff_A_Z0sc88C71_0),.clk(gclk));
	jdff dff_A_LS0OlbDu1_0(.dout(w_dff_A_Z0sc88C71_0),.din(w_dff_A_LS0OlbDu1_0),.clk(gclk));
	jdff dff_A_ezwITuSn2_1(.dout(w_n144_0[1]),.din(w_dff_A_ezwITuSn2_1),.clk(gclk));
	jdff dff_A_k8eG48ky1_1(.dout(w_dff_A_ezwITuSn2_1),.din(w_dff_A_k8eG48ky1_1),.clk(gclk));
	jdff dff_A_QpL5amcm0_2(.dout(w_n159_0[2]),.din(w_dff_A_QpL5amcm0_2),.clk(gclk));
	jdff dff_A_xZt7LRzF2_2(.dout(w_dff_A_QpL5amcm0_2),.din(w_dff_A_xZt7LRzF2_2),.clk(gclk));
	jdff dff_A_GnX2E4J12_2(.dout(w_n121_0[2]),.din(w_dff_A_GnX2E4J12_2),.clk(gclk));
	jdff dff_B_m8neVkhE9_3(.din(n121),.dout(w_dff_B_m8neVkhE9_3),.clk(gclk));
	jdff dff_A_XWqpTgAq9_1(.dout(w_n96_0[1]),.din(w_dff_A_XWqpTgAq9_1),.clk(gclk));
	jdff dff_A_EWvyHitg1_1(.dout(w_dff_A_XWqpTgAq9_1),.din(w_dff_A_EWvyHitg1_1),.clk(gclk));
	jdff dff_A_ZACxQElf1_1(.dout(w_dff_A_EWvyHitg1_1),.din(w_dff_A_ZACxQElf1_1),.clk(gclk));
	jdff dff_A_l9XTGDeg8_1(.dout(w_dff_A_ZACxQElf1_1),.din(w_dff_A_l9XTGDeg8_1),.clk(gclk));
	jdff dff_A_npN2hmbO2_2(.dout(w_n96_0[2]),.din(w_dff_A_npN2hmbO2_2),.clk(gclk));
	jdff dff_A_2FZx9MYs5_2(.dout(w_dff_A_npN2hmbO2_2),.din(w_dff_A_2FZx9MYs5_2),.clk(gclk));
	jdff dff_A_l35YzkKC2_2(.dout(w_dff_A_2FZx9MYs5_2),.din(w_dff_A_l35YzkKC2_2),.clk(gclk));
	jdff dff_A_fHH7YDY19_2(.dout(w_dff_A_l35YzkKC2_2),.din(w_dff_A_fHH7YDY19_2),.clk(gclk));
	jdff dff_B_pLektpro5_3(.din(n340),.dout(w_dff_B_pLektpro5_3),.clk(gclk));
	jdff dff_B_H8ARiGba5_3(.din(w_dff_B_pLektpro5_3),.dout(w_dff_B_H8ARiGba5_3),.clk(gclk));
	jdff dff_B_6yfJjcJB8_3(.din(w_dff_B_H8ARiGba5_3),.dout(w_dff_B_6yfJjcJB8_3),.clk(gclk));
	jdff dff_B_9H8gVqG19_3(.din(w_dff_B_6yfJjcJB8_3),.dout(w_dff_B_9H8gVqG19_3),.clk(gclk));
	jdff dff_B_ompYDYwR9_3(.din(w_dff_B_9H8gVqG19_3),.dout(w_dff_B_ompYDYwR9_3),.clk(gclk));
	jdff dff_B_MUwemsSK1_3(.din(w_dff_B_ompYDYwR9_3),.dout(w_dff_B_MUwemsSK1_3),.clk(gclk));
	jdff dff_B_DTKlaCO11_3(.din(w_dff_B_MUwemsSK1_3),.dout(w_dff_B_DTKlaCO11_3),.clk(gclk));
	jdff dff_B_rN5AlINv4_3(.din(w_dff_B_DTKlaCO11_3),.dout(w_dff_B_rN5AlINv4_3),.clk(gclk));
	jdff dff_B_IWPAWgS61_3(.din(w_dff_B_rN5AlINv4_3),.dout(w_dff_B_IWPAWgS61_3),.clk(gclk));
	jdff dff_B_9d9lGbvZ4_3(.din(w_dff_B_IWPAWgS61_3),.dout(w_dff_B_9d9lGbvZ4_3),.clk(gclk));
	jdff dff_B_flcQQ9b53_3(.din(w_dff_B_9d9lGbvZ4_3),.dout(w_dff_B_flcQQ9b53_3),.clk(gclk));
	jdff dff_B_dj9wFQAO7_3(.din(w_dff_B_flcQQ9b53_3),.dout(w_dff_B_dj9wFQAO7_3),.clk(gclk));
	jdff dff_B_9i4j02lf4_3(.din(w_dff_B_dj9wFQAO7_3),.dout(w_dff_B_9i4j02lf4_3),.clk(gclk));
	jdff dff_B_swvHy0uK6_3(.din(w_dff_B_9i4j02lf4_3),.dout(w_dff_B_swvHy0uK6_3),.clk(gclk));
	jdff dff_B_7JHBBpwe3_3(.din(w_dff_B_swvHy0uK6_3),.dout(w_dff_B_7JHBBpwe3_3),.clk(gclk));
	jdff dff_B_zDweCeiP0_3(.din(w_dff_B_7JHBBpwe3_3),.dout(w_dff_B_zDweCeiP0_3),.clk(gclk));
	jdff dff_B_pG1xOg5Q9_1(.din(n394),.dout(w_dff_B_pG1xOg5Q9_1),.clk(gclk));
	jdff dff_B_g28bMA9v8_1(.din(w_dff_B_pG1xOg5Q9_1),.dout(w_dff_B_g28bMA9v8_1),.clk(gclk));
	jdff dff_B_hllqSuK67_1(.din(w_dff_B_g28bMA9v8_1),.dout(w_dff_B_hllqSuK67_1),.clk(gclk));
	jdff dff_B_g7eQvssc8_1(.din(w_dff_B_hllqSuK67_1),.dout(w_dff_B_g7eQvssc8_1),.clk(gclk));
	jdff dff_B_tls9DdDw4_1(.din(w_dff_B_g7eQvssc8_1),.dout(w_dff_B_tls9DdDw4_1),.clk(gclk));
	jdff dff_B_OLaJSHoj9_1(.din(w_dff_B_tls9DdDw4_1),.dout(w_dff_B_OLaJSHoj9_1),.clk(gclk));
	jdff dff_B_nysGo9QM1_1(.din(w_dff_B_OLaJSHoj9_1),.dout(w_dff_B_nysGo9QM1_1),.clk(gclk));
	jdff dff_B_r86hjLOJ8_1(.din(w_dff_B_nysGo9QM1_1),.dout(w_dff_B_r86hjLOJ8_1),.clk(gclk));
	jdff dff_B_iYKnZW357_1(.din(w_dff_B_r86hjLOJ8_1),.dout(w_dff_B_iYKnZW357_1),.clk(gclk));
	jdff dff_B_dFZsLN1Y7_1(.din(w_dff_B_iYKnZW357_1),.dout(w_dff_B_dFZsLN1Y7_1),.clk(gclk));
	jdff dff_B_MRxDTQWd2_1(.din(w_dff_B_dFZsLN1Y7_1),.dout(w_dff_B_MRxDTQWd2_1),.clk(gclk));
	jdff dff_B_dEAPrYKo2_0(.din(n396),.dout(w_dff_B_dEAPrYKo2_0),.clk(gclk));
	jdff dff_B_w2JDPKYv3_0(.din(w_dff_B_dEAPrYKo2_0),.dout(w_dff_B_w2JDPKYv3_0),.clk(gclk));
	jdff dff_B_VGT2LlO66_0(.din(w_dff_B_w2JDPKYv3_0),.dout(w_dff_B_VGT2LlO66_0),.clk(gclk));
	jdff dff_B_yQodEHlx0_0(.din(w_dff_B_VGT2LlO66_0),.dout(w_dff_B_yQodEHlx0_0),.clk(gclk));
	jdff dff_B_KPuWEk0j7_0(.din(w_dff_B_yQodEHlx0_0),.dout(w_dff_B_KPuWEk0j7_0),.clk(gclk));
	jdff dff_B_bbrLuMRc2_0(.din(w_dff_B_KPuWEk0j7_0),.dout(w_dff_B_bbrLuMRc2_0),.clk(gclk));
	jdff dff_B_X306fpbu2_0(.din(w_dff_B_bbrLuMRc2_0),.dout(w_dff_B_X306fpbu2_0),.clk(gclk));
	jdff dff_B_GGY02Drb7_0(.din(w_dff_B_X306fpbu2_0),.dout(w_dff_B_GGY02Drb7_0),.clk(gclk));
	jdff dff_B_Oie8pYVk4_0(.din(w_dff_B_GGY02Drb7_0),.dout(w_dff_B_Oie8pYVk4_0),.clk(gclk));
	jdff dff_B_NYJln6Np0_0(.din(w_dff_B_Oie8pYVk4_0),.dout(w_dff_B_NYJln6Np0_0),.clk(gclk));
	jdff dff_B_1StzCjHM6_0(.din(w_dff_B_NYJln6Np0_0),.dout(w_dff_B_1StzCjHM6_0),.clk(gclk));
	jdff dff_B_rkG1HUsr8_0(.din(w_dff_B_1StzCjHM6_0),.dout(w_dff_B_rkG1HUsr8_0),.clk(gclk));
	jdff dff_B_EQJPGoen2_0(.din(w_dff_B_rkG1HUsr8_0),.dout(w_dff_B_EQJPGoen2_0),.clk(gclk));
	jdff dff_B_cXxrWteb3_0(.din(w_dff_B_EQJPGoen2_0),.dout(w_dff_B_cXxrWteb3_0),.clk(gclk));
	jdff dff_A_NIax9h3X6_0(.dout(w_n395_0[0]),.din(w_dff_A_NIax9h3X6_0),.clk(gclk));
	jdff dff_A_iKKKJ23l9_0(.dout(w_dff_A_NIax9h3X6_0),.din(w_dff_A_iKKKJ23l9_0),.clk(gclk));
	jdff dff_A_xlTmhS4j5_0(.dout(w_dff_A_iKKKJ23l9_0),.din(w_dff_A_xlTmhS4j5_0),.clk(gclk));
	jdff dff_A_IXviYaWx1_0(.dout(w_dff_A_xlTmhS4j5_0),.din(w_dff_A_IXviYaWx1_0),.clk(gclk));
	jdff dff_A_kTeVdeRX4_0(.dout(w_dff_A_IXviYaWx1_0),.din(w_dff_A_kTeVdeRX4_0),.clk(gclk));
	jdff dff_A_SE7hUOsb9_0(.dout(w_dff_A_kTeVdeRX4_0),.din(w_dff_A_SE7hUOsb9_0),.clk(gclk));
	jdff dff_A_swHCo9AP2_0(.dout(w_dff_A_SE7hUOsb9_0),.din(w_dff_A_swHCo9AP2_0),.clk(gclk));
	jdff dff_A_Vrwm4S622_0(.dout(w_dff_A_swHCo9AP2_0),.din(w_dff_A_Vrwm4S622_0),.clk(gclk));
	jdff dff_A_gbnZpzJY2_0(.dout(w_dff_A_Vrwm4S622_0),.din(w_dff_A_gbnZpzJY2_0),.clk(gclk));
	jdff dff_A_M7iHoaWE9_0(.dout(w_dff_A_gbnZpzJY2_0),.din(w_dff_A_M7iHoaWE9_0),.clk(gclk));
	jdff dff_A_GYTrGeeS0_0(.dout(w_dff_A_M7iHoaWE9_0),.din(w_dff_A_GYTrGeeS0_0),.clk(gclk));
	jdff dff_A_q4Y4a0Yf6_0(.dout(w_dff_A_GYTrGeeS0_0),.din(w_dff_A_q4Y4a0Yf6_0),.clk(gclk));
	jdff dff_A_8hE18YhF3_0(.dout(w_dff_A_q4Y4a0Yf6_0),.din(w_dff_A_8hE18YhF3_0),.clk(gclk));
	jdff dff_A_kyDYNBv42_0(.dout(w_dff_A_8hE18YhF3_0),.din(w_dff_A_kyDYNBv42_0),.clk(gclk));
	jdff dff_A_j9yRjunC8_0(.dout(w_dff_A_kyDYNBv42_0),.din(w_dff_A_j9yRjunC8_0),.clk(gclk));
	jdff dff_B_48Z0yb8N8_0(.din(n329),.dout(w_dff_B_48Z0yb8N8_0),.clk(gclk));
	jdff dff_B_Z1qjeC8T8_0(.din(n323),.dout(w_dff_B_Z1qjeC8T8_0),.clk(gclk));
	jdff dff_A_TcrzHSSq9_1(.dout(w_n189_0[1]),.din(w_dff_A_TcrzHSSq9_1),.clk(gclk));
	jdff dff_A_TmET4rrF7_1(.dout(w_dff_A_TcrzHSSq9_1),.din(w_dff_A_TmET4rrF7_1),.clk(gclk));
	jdff dff_B_DjmXnYWK5_2(.din(n318),.dout(w_dff_B_DjmXnYWK5_2),.clk(gclk));
	jdff dff_A_8FL7BuWU7_1(.dout(w_n185_0[1]),.din(w_dff_A_8FL7BuWU7_1),.clk(gclk));
	jdff dff_A_PmJZcSWs4_1(.dout(w_dff_A_8FL7BuWU7_1),.din(w_dff_A_PmJZcSWs4_1),.clk(gclk));
	jdff dff_A_RaitYgNH5_2(.dout(w_n185_0[2]),.din(w_dff_A_RaitYgNH5_2),.clk(gclk));
	jdff dff_A_Mzvb4cNp0_2(.dout(w_dff_A_RaitYgNH5_2),.din(w_dff_A_Mzvb4cNp0_2),.clk(gclk));
	jdff dff_B_M7qw6BmR9_3(.din(n184),.dout(w_dff_B_M7qw6BmR9_3),.clk(gclk));
	jdff dff_B_pOEkBLmB1_3(.din(w_dff_B_M7qw6BmR9_3),.dout(w_dff_B_pOEkBLmB1_3),.clk(gclk));
	jdff dff_A_zxpVdtJC4_0(.dout(w_n314_0[0]),.din(w_dff_A_zxpVdtJC4_0),.clk(gclk));
	jdff dff_A_S0gXY9FI0_1(.dout(w_n314_0[1]),.din(w_dff_A_S0gXY9FI0_1),.clk(gclk));
	jdff dff_B_NvAM7Nba6_3(.din(n314),.dout(w_dff_B_NvAM7Nba6_3),.clk(gclk));
	jdff dff_A_B1jwbQ744_1(.dout(w_n311_0[1]),.din(w_dff_A_B1jwbQ744_1),.clk(gclk));
	jdff dff_A_VmapFO1s6_2(.dout(w_n311_0[2]),.din(w_dff_A_VmapFO1s6_2),.clk(gclk));
	jdff dff_B_raYUAsUH5_3(.din(n311),.dout(w_dff_B_raYUAsUH5_3),.clk(gclk));
	jdff dff_A_bALUpook7_0(.dout(w_n183_0[0]),.din(w_dff_A_bALUpook7_0),.clk(gclk));
	jdff dff_A_GLbWVTBc5_0(.dout(w_dff_A_bALUpook7_0),.din(w_dff_A_GLbWVTBc5_0),.clk(gclk));
	jdff dff_A_724vyw0z0_0(.dout(w_dff_A_GLbWVTBc5_0),.din(w_dff_A_724vyw0z0_0),.clk(gclk));
	jdff dff_A_6xpSDlhg7_1(.dout(w_n183_0[1]),.din(w_dff_A_6xpSDlhg7_1),.clk(gclk));
	jdff dff_A_v9IRINiZ2_1(.dout(w_dff_A_6xpSDlhg7_1),.din(w_dff_A_v9IRINiZ2_1),.clk(gclk));
	jdff dff_A_QPbox9xq7_1(.dout(w_dff_A_v9IRINiZ2_1),.din(w_dff_A_QPbox9xq7_1),.clk(gclk));
	jdff dff_B_CKUBDPhr6_0(.din(n182),.dout(w_dff_B_CKUBDPhr6_0),.clk(gclk));
	jdff dff_B_vaIuTYF12_1(.din(G900),.dout(w_dff_B_vaIuTYF12_1),.clk(gclk));
	jdff dff_B_PSFF9oYg4_0(.din(n304),.dout(w_dff_B_PSFF9oYg4_0),.clk(gclk));
	jdff dff_A_jiVXwrw15_1(.dout(w_n188_0[1]),.din(w_dff_A_jiVXwrw15_1),.clk(gclk));
	jdff dff_A_DPVzRc6d1_0(.dout(w_n290_0[0]),.din(w_dff_A_DPVzRc6d1_0),.clk(gclk));
	jdff dff_B_TEqAAgl68_3(.din(n290),.dout(w_dff_B_TEqAAgl68_3),.clk(gclk));
	jdff dff_A_xVKWZllH7_0(.dout(w_n289_0[0]),.din(w_dff_A_xVKWZllH7_0),.clk(gclk));
	jdff dff_A_FlTTx5ZE9_0(.dout(w_dff_A_xVKWZllH7_0),.din(w_dff_A_FlTTx5ZE9_0),.clk(gclk));
	jdff dff_B_owlxZTpc5_3(.din(n158),.dout(w_dff_B_owlxZTpc5_3),.clk(gclk));
	jdff dff_A_zc2exPZ20_0(.dout(w_n92_1[0]),.din(w_dff_A_zc2exPZ20_0),.clk(gclk));
	jdff dff_A_mNchYbv10_0(.dout(w_dff_A_zc2exPZ20_0),.din(w_dff_A_mNchYbv10_0),.clk(gclk));
	jdff dff_A_OFRntSuX5_2(.dout(w_n92_1[2]),.din(w_dff_A_OFRntSuX5_2),.clk(gclk));
	jdff dff_A_uma05frZ8_2(.dout(w_dff_A_OFRntSuX5_2),.din(w_dff_A_uma05frZ8_2),.clk(gclk));
	jdff dff_B_rjIpW8xh5_2(.din(n286),.dout(w_dff_B_rjIpW8xh5_2),.clk(gclk));
	jdff dff_A_rmQXyUD25_1(.dout(w_n163_0[1]),.din(w_dff_A_rmQXyUD25_1),.clk(gclk));
	jdff dff_A_LI1M4O6h8_1(.dout(w_dff_A_rmQXyUD25_1),.din(w_dff_A_LI1M4O6h8_1),.clk(gclk));
	jdff dff_A_qBFBJK5w9_2(.dout(w_n163_0[2]),.din(w_dff_A_qBFBJK5w9_2),.clk(gclk));
	jdff dff_A_RUEtXAqY8_2(.dout(w_dff_A_qBFBJK5w9_2),.din(w_dff_A_RUEtXAqY8_2),.clk(gclk));
	jdff dff_B_Qp1ZNaVn8_1(.din(n123),.dout(w_dff_B_Qp1ZNaVn8_1),.clk(gclk));
	jdff dff_B_LM6CR5XI4_1(.din(w_dff_B_Qp1ZNaVn8_1),.dout(w_dff_B_LM6CR5XI4_1),.clk(gclk));
	jdff dff_B_HvLhY8AC0_1(.din(w_dff_B_LM6CR5XI4_1),.dout(w_dff_B_HvLhY8AC0_1),.clk(gclk));
	jdff dff_B_5Joslp8J0_1(.din(w_dff_B_HvLhY8AC0_1),.dout(w_dff_B_5Joslp8J0_1),.clk(gclk));
	jdff dff_B_c9ZLC9CU5_1(.din(w_dff_B_5Joslp8J0_1),.dout(w_dff_B_c9ZLC9CU5_1),.clk(gclk));
	jdff dff_A_7J0PynwU1_0(.dout(w_n68_0[0]),.din(w_dff_A_7J0PynwU1_0),.clk(gclk));
	jdff dff_A_mAI8a6530_0(.dout(w_dff_A_7J0PynwU1_0),.din(w_dff_A_mAI8a6530_0),.clk(gclk));
	jdff dff_A_VYcFzFhk6_0(.dout(w_dff_A_mAI8a6530_0),.din(w_dff_A_VYcFzFhk6_0),.clk(gclk));
	jdff dff_A_XWYVQCkV9_0(.dout(w_dff_A_VYcFzFhk6_0),.din(w_dff_A_XWYVQCkV9_0),.clk(gclk));
	jdff dff_A_pF8YWz8c8_0(.dout(w_dff_A_XWYVQCkV9_0),.din(w_dff_A_pF8YWz8c8_0),.clk(gclk));
	jdff dff_A_Exlr2Eoo1_0(.dout(w_dff_A_pF8YWz8c8_0),.din(w_dff_A_Exlr2Eoo1_0),.clk(gclk));
	jdff dff_A_BYVIeeHr4_0(.dout(w_dff_A_Exlr2Eoo1_0),.din(w_dff_A_BYVIeeHr4_0),.clk(gclk));
	jdff dff_A_vjDNgY8s5_0(.dout(w_dff_A_BYVIeeHr4_0),.din(w_dff_A_vjDNgY8s5_0),.clk(gclk));
	jdff dff_A_YlonpCgY7_0(.dout(w_dff_A_vjDNgY8s5_0),.din(w_dff_A_YlonpCgY7_0),.clk(gclk));
	jdff dff_A_TCZ09ifv2_0(.dout(w_dff_A_YlonpCgY7_0),.din(w_dff_A_TCZ09ifv2_0),.clk(gclk));
	jdff dff_A_IrqCsY0U8_0(.dout(w_n281_0[0]),.din(w_dff_A_IrqCsY0U8_0),.clk(gclk));
	jdff dff_A_juWZbGN95_1(.dout(w_n281_0[1]),.din(w_dff_A_juWZbGN95_1),.clk(gclk));
	jdff dff_B_bEywQSYi2_3(.din(n281),.dout(w_dff_B_bEywQSYi2_3),.clk(gclk));
	jdff dff_B_bdT2QtA68_2(.din(n278),.dout(w_dff_B_bdT2QtA68_2),.clk(gclk));
	jdff dff_A_Tz13o3B98_1(.dout(w_n168_0[1]),.din(w_dff_A_Tz13o3B98_1),.clk(gclk));
	jdff dff_A_GoMmkFZB3_1(.dout(w_dff_A_Tz13o3B98_1),.din(w_dff_A_GoMmkFZB3_1),.clk(gclk));
	jdff dff_A_LD3Dv2xE4_2(.dout(w_n168_0[2]),.din(w_dff_A_LD3Dv2xE4_2),.clk(gclk));
	jdff dff_A_5TdxSzju1_2(.dout(w_dff_A_LD3Dv2xE4_2),.din(w_dff_A_5TdxSzju1_2),.clk(gclk));
	jdff dff_B_5bAE8v1W6_1(.din(n133),.dout(w_dff_B_5bAE8v1W6_1),.clk(gclk));
	jdff dff_B_yBRMCjK85_1(.din(w_dff_B_5bAE8v1W6_1),.dout(w_dff_B_yBRMCjK85_1),.clk(gclk));
	jdff dff_B_8L2iblMT8_1(.din(w_dff_B_yBRMCjK85_1),.dout(w_dff_B_8L2iblMT8_1),.clk(gclk));
	jdff dff_B_zqYjqX8i2_1(.din(w_dff_B_8L2iblMT8_1),.dout(w_dff_B_zqYjqX8i2_1),.clk(gclk));
	jdff dff_B_0iPv6gzG1_1(.din(w_dff_B_zqYjqX8i2_1),.dout(w_dff_B_0iPv6gzG1_1),.clk(gclk));
	jdff dff_A_rEBYjwos2_0(.dout(w_n141_0[0]),.din(w_dff_A_rEBYjwos2_0),.clk(gclk));
	jdff dff_A_7e25JeQW8_0(.dout(w_dff_A_rEBYjwos2_0),.din(w_dff_A_7e25JeQW8_0),.clk(gclk));
	jdff dff_A_Bbeih4ml6_0(.dout(w_dff_A_7e25JeQW8_0),.din(w_dff_A_Bbeih4ml6_0),.clk(gclk));
	jdff dff_A_05gUz8eC3_0(.dout(w_dff_A_Bbeih4ml6_0),.din(w_dff_A_05gUz8eC3_0),.clk(gclk));
	jdff dff_A_bH7EHXLC5_0(.dout(w_dff_A_05gUz8eC3_0),.din(w_dff_A_bH7EHXLC5_0),.clk(gclk));
	jdff dff_A_X13iLN897_0(.dout(w_dff_A_bH7EHXLC5_0),.din(w_dff_A_X13iLN897_0),.clk(gclk));
	jdff dff_A_uiojGWRL6_0(.dout(w_dff_A_X13iLN897_0),.din(w_dff_A_uiojGWRL6_0),.clk(gclk));
	jdff dff_A_JjRXqtp87_0(.dout(w_dff_A_uiojGWRL6_0),.din(w_dff_A_JjRXqtp87_0),.clk(gclk));
	jdff dff_A_7x6m75oJ1_0(.dout(w_dff_A_JjRXqtp87_0),.din(w_dff_A_7x6m75oJ1_0),.clk(gclk));
	jdff dff_A_DExDTuAx1_0(.dout(w_dff_A_7x6m75oJ1_0),.din(w_dff_A_DExDTuAx1_0),.clk(gclk));
	jdff dff_A_mk4gPCmd3_0(.dout(w_dff_A_DExDTuAx1_0),.din(w_dff_A_mk4gPCmd3_0),.clk(gclk));
	jdff dff_A_rGr1XINl7_0(.dout(w_dff_A_mk4gPCmd3_0),.din(w_dff_A_rGr1XINl7_0),.clk(gclk));
	jdff dff_B_jnzZwyXB6_1(.din(n134),.dout(w_dff_B_jnzZwyXB6_1),.clk(gclk));
	jdff dff_B_L8QKAwC11_1(.din(w_dff_B_jnzZwyXB6_1),.dout(w_dff_B_L8QKAwC11_1),.clk(gclk));
	jdff dff_A_53JJPNRr4_1(.dout(w_G475_0[1]),.din(w_dff_A_53JJPNRr4_1),.clk(gclk));
	jdff dff_A_o3uS6aLv0_1(.dout(w_dff_A_53JJPNRr4_1),.din(w_dff_A_o3uS6aLv0_1),.clk(gclk));
	jdff dff_A_DM8gqVOJ3_1(.dout(w_dff_A_o3uS6aLv0_1),.din(w_dff_A_DM8gqVOJ3_1),.clk(gclk));
	jdff dff_A_l6FC1KZH0_1(.dout(w_dff_A_DM8gqVOJ3_1),.din(w_dff_A_l6FC1KZH0_1),.clk(gclk));
	jdff dff_A_I28831662_1(.dout(w_dff_A_l6FC1KZH0_1),.din(w_dff_A_I28831662_1),.clk(gclk));
	jdff dff_A_OxoHZ5Ps2_1(.dout(w_dff_A_I28831662_1),.din(w_dff_A_OxoHZ5Ps2_1),.clk(gclk));
	jdff dff_A_LQhley7s3_0(.dout(w_n130_0[0]),.din(w_dff_A_LQhley7s3_0),.clk(gclk));
	jdff dff_A_nnlDv0iF6_0(.dout(w_dff_A_LQhley7s3_0),.din(w_dff_A_nnlDv0iF6_0),.clk(gclk));
	jdff dff_A_UYoiRhCm8_0(.dout(w_dff_A_nnlDv0iF6_0),.din(w_dff_A_UYoiRhCm8_0),.clk(gclk));
	jdff dff_A_GN3tzEEp0_0(.dout(w_dff_A_UYoiRhCm8_0),.din(w_dff_A_GN3tzEEp0_0),.clk(gclk));
	jdff dff_A_DMDHVcJa9_0(.dout(w_dff_A_GN3tzEEp0_0),.din(w_dff_A_DMDHVcJa9_0),.clk(gclk));
	jdff dff_A_Uk705U1L4_0(.dout(w_dff_A_DMDHVcJa9_0),.din(w_dff_A_Uk705U1L4_0),.clk(gclk));
	jdff dff_A_hTrlKjcn8_0(.dout(w_dff_A_Uk705U1L4_0),.din(w_dff_A_hTrlKjcn8_0),.clk(gclk));
	jdff dff_A_ibCtApuJ3_0(.dout(w_dff_A_hTrlKjcn8_0),.din(w_dff_A_ibCtApuJ3_0),.clk(gclk));
	jdff dff_A_32W4jJMI8_0(.dout(w_dff_A_ibCtApuJ3_0),.din(w_dff_A_32W4jJMI8_0),.clk(gclk));
	jdff dff_A_x0jYfg461_0(.dout(w_dff_A_32W4jJMI8_0),.din(w_dff_A_x0jYfg461_0),.clk(gclk));
	jdff dff_A_25ba2pdN7_0(.dout(w_dff_A_x0jYfg461_0),.din(w_dff_A_25ba2pdN7_0),.clk(gclk));
	jdff dff_A_VM9zdHHW2_0(.dout(w_dff_A_25ba2pdN7_0),.din(w_dff_A_VM9zdHHW2_0),.clk(gclk));
	jdff dff_B_bdvoMKgx8_1(.din(n124),.dout(w_dff_B_bdvoMKgx8_1),.clk(gclk));
	jdff dff_B_t0UNrw4Z3_1(.din(w_dff_B_bdvoMKgx8_1),.dout(w_dff_B_t0UNrw4Z3_1),.clk(gclk));
	jdff dff_B_IEDcSjra0_1(.din(w_dff_B_t0UNrw4Z3_1),.dout(w_dff_B_IEDcSjra0_1),.clk(gclk));
	jdff dff_B_fzf9OgLb8_0(.din(n128),.dout(w_dff_B_fzf9OgLb8_0),.clk(gclk));
	jdff dff_A_CtGg71EJ0_1(.dout(w_G478_0[1]),.din(w_dff_A_CtGg71EJ0_1),.clk(gclk));
	jdff dff_A_wXDaLGka3_1(.dout(w_dff_A_CtGg71EJ0_1),.din(w_dff_A_wXDaLGka3_1),.clk(gclk));
	jdff dff_A_p6SYAq3i8_1(.dout(w_dff_A_wXDaLGka3_1),.din(w_dff_A_p6SYAq3i8_1),.clk(gclk));
	jdff dff_A_EeA4weBH6_1(.dout(w_dff_A_p6SYAq3i8_1),.din(w_dff_A_EeA4weBH6_1),.clk(gclk));
	jdff dff_A_A1OTIQDY1_1(.dout(w_dff_A_EeA4weBH6_1),.din(w_dff_A_A1OTIQDY1_1),.clk(gclk));
	jdff dff_A_HidJcISd9_1(.dout(w_dff_A_A1OTIQDY1_1),.din(w_dff_A_HidJcISd9_1),.clk(gclk));
	jdff dff_B_cI1V1wQt5_3(.din(n154),.dout(w_dff_B_cI1V1wQt5_3),.clk(gclk));
	jdff dff_B_TII2KWyq0_3(.din(w_dff_B_cI1V1wQt5_3),.dout(w_dff_B_TII2KWyq0_3),.clk(gclk));
	jdff dff_A_VM14KFsj4_0(.dout(w_n153_0[0]),.din(w_dff_A_VM14KFsj4_0),.clk(gclk));
	jdff dff_A_pt6Y1sLI2_0(.dout(w_dff_A_VM14KFsj4_0),.din(w_dff_A_pt6Y1sLI2_0),.clk(gclk));
	jdff dff_A_7y0MB23R2_0(.dout(w_dff_A_pt6Y1sLI2_0),.din(w_dff_A_7y0MB23R2_0),.clk(gclk));
	jdff dff_A_Da3mUR3W3_1(.dout(w_n153_0[1]),.din(w_dff_A_Da3mUR3W3_1),.clk(gclk));
	jdff dff_A_GVKFDLUy0_1(.dout(w_dff_A_Da3mUR3W3_1),.din(w_dff_A_GVKFDLUy0_1),.clk(gclk));
	jdff dff_A_rICxkPtJ8_1(.dout(w_dff_A_GVKFDLUy0_1),.din(w_dff_A_rICxkPtJ8_1),.clk(gclk));
	jdff dff_B_1zEFzQYj5_1(.din(n148),.dout(w_dff_B_1zEFzQYj5_1),.clk(gclk));
	jdff dff_A_hupSypvR0_0(.dout(w_n151_0[0]),.din(w_dff_A_hupSypvR0_0),.clk(gclk));
	jdff dff_A_9hQcCyMw8_1(.dout(w_n151_0[1]),.din(w_dff_A_9hQcCyMw8_1),.clk(gclk));
	jdff dff_A_Yp6jucyo8_1(.dout(w_dff_A_9hQcCyMw8_1),.din(w_dff_A_Yp6jucyo8_1),.clk(gclk));
	jdff dff_A_VX7vXtxt6_1(.dout(w_dff_A_Yp6jucyo8_1),.din(w_dff_A_VX7vXtxt6_1),.clk(gclk));
	jdff dff_A_6DZDx5TQ8_1(.dout(w_dff_A_VX7vXtxt6_1),.din(w_dff_A_6DZDx5TQ8_1),.clk(gclk));
	jdff dff_A_NrfbGgaG0_1(.dout(w_dff_A_6DZDx5TQ8_1),.din(w_dff_A_NrfbGgaG0_1),.clk(gclk));
	jdff dff_A_XrWe4vcE5_1(.dout(w_dff_A_NrfbGgaG0_1),.din(w_dff_A_XrWe4vcE5_1),.clk(gclk));
	jdff dff_A_8voFaRrL2_1(.dout(w_dff_A_XrWe4vcE5_1),.din(w_dff_A_8voFaRrL2_1),.clk(gclk));
	jdff dff_A_YuDYZB8u6_1(.dout(w_dff_A_8voFaRrL2_1),.din(w_dff_A_YuDYZB8u6_1),.clk(gclk));
	jdff dff_A_11mm1uNl8_1(.dout(w_dff_A_YuDYZB8u6_1),.din(w_dff_A_11mm1uNl8_1),.clk(gclk));
	jdff dff_A_AtNUKxE55_1(.dout(w_dff_A_11mm1uNl8_1),.din(w_dff_A_AtNUKxE55_1),.clk(gclk));
	jdff dff_A_IbXovPq23_1(.dout(w_dff_A_AtNUKxE55_1),.din(w_dff_A_IbXovPq23_1),.clk(gclk));
	jdff dff_A_Tfcn9HTa0_1(.dout(w_G952_0[1]),.din(w_dff_A_Tfcn9HTa0_1),.clk(gclk));
	jdff dff_A_ZMW53MW68_1(.dout(w_dff_A_Tfcn9HTa0_1),.din(w_dff_A_ZMW53MW68_1),.clk(gclk));
	jdff dff_A_Vjc72R8L5_1(.dout(w_dff_A_ZMW53MW68_1),.din(w_dff_A_Vjc72R8L5_1),.clk(gclk));
	jdff dff_A_1vw4cqIS8_1(.dout(w_dff_A_Vjc72R8L5_1),.din(w_dff_A_1vw4cqIS8_1),.clk(gclk));
	jdff dff_A_SUlDxw8x9_1(.dout(w_dff_A_1vw4cqIS8_1),.din(w_dff_A_SUlDxw8x9_1),.clk(gclk));
	jdff dff_A_r5d4qCrU5_1(.dout(w_dff_A_SUlDxw8x9_1),.din(w_dff_A_r5d4qCrU5_1),.clk(gclk));
	jdff dff_A_fWz20p4R0_1(.dout(w_dff_A_r5d4qCrU5_1),.din(w_dff_A_fWz20p4R0_1),.clk(gclk));
	jdff dff_A_7Us8wD3e1_1(.dout(w_dff_A_fWz20p4R0_1),.din(w_dff_A_7Us8wD3e1_1),.clk(gclk));
	jdff dff_A_U131JysR2_1(.dout(w_dff_A_7Us8wD3e1_1),.din(w_dff_A_U131JysR2_1),.clk(gclk));
	jdff dff_A_saO30qQ77_1(.dout(w_dff_A_U131JysR2_1),.din(w_dff_A_saO30qQ77_1),.clk(gclk));
	jdff dff_A_DmHOwzrL9_1(.dout(w_dff_A_saO30qQ77_1),.din(w_dff_A_DmHOwzrL9_1),.clk(gclk));
	jdff dff_A_IoiwkHxL6_1(.dout(w_dff_A_DmHOwzrL9_1),.din(w_dff_A_IoiwkHxL6_1),.clk(gclk));
	jdff dff_A_pNwj3ERr8_1(.dout(w_dff_A_IoiwkHxL6_1),.din(w_dff_A_pNwj3ERr8_1),.clk(gclk));
	jdff dff_A_pv0B8K8e8_1(.dout(w_dff_A_pNwj3ERr8_1),.din(w_dff_A_pv0B8K8e8_1),.clk(gclk));
	jdff dff_A_wWPGREJB6_1(.dout(w_dff_A_pv0B8K8e8_1),.din(w_dff_A_wWPGREJB6_1),.clk(gclk));
	jdff dff_A_tcPEUmQq8_1(.dout(w_dff_A_wWPGREJB6_1),.din(w_dff_A_tcPEUmQq8_1),.clk(gclk));
	jdff dff_B_23RAqRpQ9_3(.din(G952),.dout(w_dff_B_23RAqRpQ9_3),.clk(gclk));
	jdff dff_B_7Y2DWtMV5_1(.din(G898),.dout(w_dff_B_7Y2DWtMV5_1),.clk(gclk));
	jdff dff_A_9iLFHuQA5_2(.dout(w_n253_0[2]),.din(w_dff_A_9iLFHuQA5_2),.clk(gclk));
	jdff dff_A_IAxImSs79_1(.dout(w_n92_0[1]),.din(w_dff_A_IAxImSs79_1),.clk(gclk));
	jdff dff_A_6LwPzpr78_1(.dout(w_dff_A_IAxImSs79_1),.din(w_dff_A_6LwPzpr78_1),.clk(gclk));
	jdff dff_A_QeIaXzPy7_2(.dout(w_n92_0[2]),.din(w_dff_A_QeIaXzPy7_2),.clk(gclk));
	jdff dff_A_j7Zy7O2B8_2(.dout(w_dff_A_QeIaXzPy7_2),.din(w_dff_A_j7Zy7O2B8_2),.clk(gclk));
	jdff dff_A_CvDs9rKb2_1(.dout(w_G472_0[1]),.din(w_dff_A_CvDs9rKb2_1),.clk(gclk));
	jdff dff_A_0p0bzACN2_1(.dout(w_dff_A_CvDs9rKb2_1),.din(w_dff_A_0p0bzACN2_1),.clk(gclk));
	jdff dff_A_cMFhgO2J9_1(.dout(w_dff_A_0p0bzACN2_1),.din(w_dff_A_cMFhgO2J9_1),.clk(gclk));
	jdff dff_A_NTcFWbYE3_1(.dout(w_dff_A_cMFhgO2J9_1),.din(w_dff_A_NTcFWbYE3_1),.clk(gclk));
	jdff dff_A_HvS80Czb7_1(.dout(w_dff_A_NTcFWbYE3_1),.din(w_dff_A_HvS80Czb7_1),.clk(gclk));
	jdff dff_A_j5LbCEsr0_1(.dout(w_dff_A_HvS80Czb7_1),.din(w_dff_A_j5LbCEsr0_1),.clk(gclk));
	jdff dff_B_3HrIOuAs7_2(.din(n73),.dout(w_dff_B_3HrIOuAs7_2),.clk(gclk));
	jdff dff_B_gSd8pB4c1_2(.din(w_dff_B_3HrIOuAs7_2),.dout(w_dff_B_gSd8pB4c1_2),.clk(gclk));
	jdff dff_B_n1oB1xGr7_2(.din(w_dff_B_gSd8pB4c1_2),.dout(w_dff_B_n1oB1xGr7_2),.clk(gclk));
	jdff dff_B_AJ4NIPbd6_2(.din(w_dff_B_n1oB1xGr7_2),.dout(w_dff_B_AJ4NIPbd6_2),.clk(gclk));
	jdff dff_A_B7k92NuB0_1(.dout(w_G217_0[1]),.din(w_dff_A_B7k92NuB0_1),.clk(gclk));
	jdff dff_A_zl8609TL1_1(.dout(w_dff_A_B7k92NuB0_1),.din(w_dff_A_zl8609TL1_1),.clk(gclk));
	jdff dff_A_gAP7lnGJ9_2(.dout(w_G217_0[2]),.din(w_dff_A_gAP7lnGJ9_2),.clk(gclk));
	jdff dff_A_QFYNjmhw9_2(.dout(w_dff_A_gAP7lnGJ9_2),.din(w_dff_A_QFYNjmhw9_2),.clk(gclk));
	jdff dff_A_0FYkV1dJ2_2(.dout(w_dff_A_QFYNjmhw9_2),.din(w_dff_A_0FYkV1dJ2_2),.clk(gclk));
	jdff dff_A_L5vz5Btl7_0(.dout(w_n172_0[0]),.din(w_dff_A_L5vz5Btl7_0),.clk(gclk));
	jdff dff_A_01SBQoWa6_0(.dout(w_dff_A_L5vz5Btl7_0),.din(w_dff_A_01SBQoWa6_0),.clk(gclk));
	jdff dff_A_gE7Nowti9_0(.dout(w_dff_A_01SBQoWa6_0),.din(w_dff_A_gE7Nowti9_0),.clk(gclk));
	jdff dff_A_zBOTKbEV6_0(.dout(w_dff_A_gE7Nowti9_0),.din(w_dff_A_zBOTKbEV6_0),.clk(gclk));
	jdff dff_A_iHmhUX007_0(.dout(w_dff_A_zBOTKbEV6_0),.din(w_dff_A_iHmhUX007_0),.clk(gclk));
	jdff dff_A_6HqoROxp0_0(.dout(w_dff_A_iHmhUX007_0),.din(w_dff_A_6HqoROxp0_0),.clk(gclk));
	jdff dff_A_klwCKbVv7_0(.dout(w_dff_A_6HqoROxp0_0),.din(w_dff_A_klwCKbVv7_0),.clk(gclk));
	jdff dff_A_Cnsov7UN0_0(.dout(w_dff_A_klwCKbVv7_0),.din(w_dff_A_Cnsov7UN0_0),.clk(gclk));
	jdff dff_A_KoiLVggi2_0(.dout(w_dff_A_Cnsov7UN0_0),.din(w_dff_A_KoiLVggi2_0),.clk(gclk));
	jdff dff_A_i59WwYfY7_0(.dout(w_dff_A_KoiLVggi2_0),.din(w_dff_A_i59WwYfY7_0),.clk(gclk));
	jdff dff_B_vGQlEkZ78_1(.din(n171),.dout(w_dff_B_vGQlEkZ78_1),.clk(gclk));
	jdff dff_B_Bw6YcVAi9_1(.din(w_dff_B_vGQlEkZ78_1),.dout(w_dff_B_Bw6YcVAi9_1),.clk(gclk));
	jdff dff_B_MBQeGfwG0_1(.din(w_dff_B_Bw6YcVAi9_1),.dout(w_dff_B_MBQeGfwG0_1),.clk(gclk));
	jdff dff_B_iV8nUqg47_0(.din(n65),.dout(w_dff_B_iV8nUqg47_0),.clk(gclk));
	jdff dff_B_NNq6FVvX2_0(.din(w_dff_B_iV8nUqg47_0),.dout(w_dff_B_NNq6FVvX2_0),.clk(gclk));
	jdff dff_B_BelyrYIz1_0(.din(w_dff_B_NNq6FVvX2_0),.dout(w_dff_B_BelyrYIz1_0),.clk(gclk));
	jdff dff_A_fFZrmiXs5_2(.dout(w_n60_0[2]),.din(w_dff_A_fFZrmiXs5_2),.clk(gclk));
	jdff dff_A_AmL7gSWu2_2(.dout(w_dff_A_fFZrmiXs5_2),.din(w_dff_A_AmL7gSWu2_2),.clk(gclk));
	jdff dff_A_rUkWVoqt7_2(.dout(w_dff_A_AmL7gSWu2_2),.din(w_dff_A_rUkWVoqt7_2),.clk(gclk));
	jdff dff_A_honyHz3o2_2(.dout(w_dff_A_rUkWVoqt7_2),.din(w_dff_A_honyHz3o2_2),.clk(gclk));
	jdff dff_A_rQXRt57y5_0(.dout(w_n59_0[0]),.din(w_dff_A_rQXRt57y5_0),.clk(gclk));
	jdff dff_A_UIGrPf6h3_0(.dout(w_dff_A_rQXRt57y5_0),.din(w_dff_A_UIGrPf6h3_0),.clk(gclk));
	jdff dff_A_NRjXV6Yh0_0(.dout(w_dff_A_UIGrPf6h3_0),.din(w_dff_A_NRjXV6Yh0_0),.clk(gclk));
	jdff dff_A_814i3DzR1_0(.dout(w_n70_1[0]),.din(w_dff_A_814i3DzR1_0),.clk(gclk));
	jdff dff_A_qM7cLgsS9_0(.dout(w_dff_A_814i3DzR1_0),.din(w_dff_A_qM7cLgsS9_0),.clk(gclk));
	jdff dff_A_IQMPX2U20_0(.dout(w_dff_A_qM7cLgsS9_0),.din(w_dff_A_IQMPX2U20_0),.clk(gclk));
	jdff dff_A_YeUhj9EY4_0(.dout(w_dff_A_IQMPX2U20_0),.din(w_dff_A_YeUhj9EY4_0),.clk(gclk));
	jdff dff_A_tjj0vqVn2_0(.dout(w_dff_A_YeUhj9EY4_0),.din(w_dff_A_tjj0vqVn2_0),.clk(gclk));
	jdff dff_A_PyS38Hry9_0(.dout(w_dff_A_tjj0vqVn2_0),.din(w_dff_A_PyS38Hry9_0),.clk(gclk));
	jdff dff_A_W8ddvjR15_2(.dout(w_n70_1[2]),.din(w_dff_A_W8ddvjR15_2),.clk(gclk));
	jdff dff_A_iRp9Pgqu7_2(.dout(w_dff_A_W8ddvjR15_2),.din(w_dff_A_iRp9Pgqu7_2),.clk(gclk));
	jdff dff_A_6Stgew7U1_2(.dout(w_dff_A_iRp9Pgqu7_2),.din(w_dff_A_6Stgew7U1_2),.clk(gclk));
	jdff dff_A_zWlwC2Ou2_2(.dout(w_dff_A_6Stgew7U1_2),.din(w_dff_A_zWlwC2Ou2_2),.clk(gclk));
	jdff dff_A_aK5RmE8l4_0(.dout(w_n276_1[0]),.din(w_dff_A_aK5RmE8l4_0),.clk(gclk));
	jdff dff_B_Noibk2AT2_3(.din(n276),.dout(w_dff_B_Noibk2AT2_3),.clk(gclk));
	jdff dff_B_wO5IPQdQ4_1(.din(n195),.dout(w_dff_B_wO5IPQdQ4_1),.clk(gclk));
	jdff dff_B_DoqiWlGc8_1(.din(w_dff_B_wO5IPQdQ4_1),.dout(w_dff_B_DoqiWlGc8_1),.clk(gclk));
	jdff dff_B_054wAfNi9_1(.din(w_dff_B_DoqiWlGc8_1),.dout(w_dff_B_054wAfNi9_1),.clk(gclk));
	jdff dff_B_YiO9UU9a3_1(.din(w_dff_B_054wAfNi9_1),.dout(w_dff_B_YiO9UU9a3_1),.clk(gclk));
	jdff dff_B_IDrOGnTz9_1(.din(w_dff_B_YiO9UU9a3_1),.dout(w_dff_B_IDrOGnTz9_1),.clk(gclk));
	jdff dff_A_g1zixX7E3_0(.dout(w_n117_0[0]),.din(w_dff_A_g1zixX7E3_0),.clk(gclk));
	jdff dff_A_tpkSHp4F4_0(.dout(w_dff_A_g1zixX7E3_0),.din(w_dff_A_tpkSHp4F4_0),.clk(gclk));
	jdff dff_A_vXyxFrkh0_0(.dout(w_dff_A_tpkSHp4F4_0),.din(w_dff_A_vXyxFrkh0_0),.clk(gclk));
	jdff dff_A_EHajfGsu6_0(.dout(w_dff_A_vXyxFrkh0_0),.din(w_dff_A_EHajfGsu6_0),.clk(gclk));
	jdff dff_A_AUESdjAj7_0(.dout(w_dff_A_EHajfGsu6_0),.din(w_dff_A_AUESdjAj7_0),.clk(gclk));
	jdff dff_A_ehIEWmHZ3_0(.dout(w_dff_A_AUESdjAj7_0),.din(w_dff_A_ehIEWmHZ3_0),.clk(gclk));
	jdff dff_A_2g9Q7j5z3_0(.dout(w_dff_A_ehIEWmHZ3_0),.din(w_dff_A_2g9Q7j5z3_0),.clk(gclk));
	jdff dff_A_B7KGnKDP7_0(.dout(w_dff_A_2g9Q7j5z3_0),.din(w_dff_A_B7KGnKDP7_0),.clk(gclk));
	jdff dff_A_smkwssbt8_0(.dout(w_dff_A_B7KGnKDP7_0),.din(w_dff_A_smkwssbt8_0),.clk(gclk));
	jdff dff_A_mfNqk30O9_0(.dout(w_dff_A_smkwssbt8_0),.din(w_dff_A_mfNqk30O9_0),.clk(gclk));
	jdff dff_A_j87yRcQF3_0(.dout(w_dff_A_mfNqk30O9_0),.din(w_dff_A_j87yRcQF3_0),.clk(gclk));
	jdff dff_A_VzVx22lW7_0(.dout(w_dff_A_j87yRcQF3_0),.din(w_dff_A_VzVx22lW7_0),.clk(gclk));
	jdff dff_B_eKKvfRZ89_1(.din(n113),.dout(w_dff_B_eKKvfRZ89_1),.clk(gclk));
	jdff dff_B_eXj6DoYl4_1(.din(w_dff_B_eKKvfRZ89_1),.dout(w_dff_B_eXj6DoYl4_1),.clk(gclk));
	jdff dff_B_cFSZjj0a2_2(.din(G227),.dout(w_dff_B_cFSZjj0a2_2),.clk(gclk));
	jdff dff_A_leZGNIq02_0(.dout(w_G140_0[0]),.din(w_dff_A_leZGNIq02_0),.clk(gclk));
	jdff dff_A_1PN84TZ54_0(.dout(w_dff_A_leZGNIq02_0),.din(w_dff_A_1PN84TZ54_0),.clk(gclk));
	jdff dff_A_FzLgC7cX9_0(.dout(w_dff_A_1PN84TZ54_0),.din(w_dff_A_FzLgC7cX9_0),.clk(gclk));
	jdff dff_A_4gt6HTaA9_0(.dout(w_dff_A_FzLgC7cX9_0),.din(w_dff_A_4gt6HTaA9_0),.clk(gclk));
	jdff dff_A_AnPH0Xfn5_0(.dout(w_dff_A_4gt6HTaA9_0),.din(w_dff_A_AnPH0Xfn5_0),.clk(gclk));
	jdff dff_A_aVzZ3h7f1_0(.dout(w_dff_A_AnPH0Xfn5_0),.din(w_dff_A_aVzZ3h7f1_0),.clk(gclk));
	jdff dff_A_CFJD27Pf8_0(.dout(w_dff_A_aVzZ3h7f1_0),.din(w_dff_A_CFJD27Pf8_0),.clk(gclk));
	jdff dff_A_0CqJW5CV4_0(.dout(w_dff_A_CFJD27Pf8_0),.din(w_dff_A_0CqJW5CV4_0),.clk(gclk));
	jdff dff_A_VrUYHfgX8_0(.dout(w_dff_A_0CqJW5CV4_0),.din(w_dff_A_VrUYHfgX8_0),.clk(gclk));
	jdff dff_A_w2N3Q8iA4_0(.dout(w_dff_A_VrUYHfgX8_0),.din(w_dff_A_w2N3Q8iA4_0),.clk(gclk));
	jdff dff_A_CmjkHV433_0(.dout(w_dff_A_w2N3Q8iA4_0),.din(w_dff_A_CmjkHV433_0),.clk(gclk));
	jdff dff_A_YVDvWf2Z5_0(.dout(w_dff_A_CmjkHV433_0),.din(w_dff_A_YVDvWf2Z5_0),.clk(gclk));
	jdff dff_A_kYbTGiMo9_2(.dout(w_G469_0[2]),.din(w_dff_A_kYbTGiMo9_2),.clk(gclk));
	jdff dff_A_oZdnrC5n2_2(.dout(w_dff_A_kYbTGiMo9_2),.din(w_dff_A_oZdnrC5n2_2),.clk(gclk));
	jdff dff_A_Ih4YruBg6_2(.dout(w_dff_A_oZdnrC5n2_2),.din(w_dff_A_Ih4YruBg6_2),.clk(gclk));
	jdff dff_A_QMRJReU24_2(.dout(w_dff_A_Ih4YruBg6_2),.din(w_dff_A_QMRJReU24_2),.clk(gclk));
	jdff dff_A_J7KElagk8_2(.dout(w_dff_A_QMRJReU24_2),.din(w_dff_A_J7KElagk8_2),.clk(gclk));
	jdff dff_A_kUKg9n2E9_2(.dout(w_dff_A_J7KElagk8_2),.din(w_dff_A_kUKg9n2E9_2),.clk(gclk));
	jdff dff_B_DmgtZOLf4_2(.din(n274),.dout(w_dff_B_DmgtZOLf4_2),.clk(gclk));
	jdff dff_B_7kQIQ15r4_2(.din(w_dff_B_DmgtZOLf4_2),.dout(w_dff_B_7kQIQ15r4_2),.clk(gclk));
	jdff dff_B_IxfoKFtQ6_2(.din(w_dff_B_7kQIQ15r4_2),.dout(w_dff_B_IxfoKFtQ6_2),.clk(gclk));
	jdff dff_A_EdUnV6IY8_0(.dout(w_n112_0[0]),.din(w_dff_A_EdUnV6IY8_0),.clk(gclk));
	jdff dff_A_u3i1uTpQ7_0(.dout(w_dff_A_EdUnV6IY8_0),.din(w_dff_A_u3i1uTpQ7_0),.clk(gclk));
	jdff dff_A_dcsRzTbO3_0(.dout(w_dff_A_u3i1uTpQ7_0),.din(w_dff_A_dcsRzTbO3_0),.clk(gclk));
	jdff dff_A_QhbAil4O7_0(.dout(w_dff_A_dcsRzTbO3_0),.din(w_dff_A_QhbAil4O7_0),.clk(gclk));
	jdff dff_B_rah6lkTt0_1(.din(n111),.dout(w_dff_B_rah6lkTt0_1),.clk(gclk));
	jdff dff_A_3Rl7pbnY6_0(.dout(w_n70_3[0]),.din(w_dff_A_3Rl7pbnY6_0),.clk(gclk));
	jdff dff_A_redLIpgw6_0(.dout(w_dff_A_3Rl7pbnY6_0),.din(w_dff_A_redLIpgw6_0),.clk(gclk));
	jdff dff_A_WkPdH8WO6_0(.dout(w_dff_A_redLIpgw6_0),.din(w_dff_A_WkPdH8WO6_0),.clk(gclk));
	jdff dff_A_60j5QT485_0(.dout(w_dff_A_WkPdH8WO6_0),.din(w_dff_A_60j5QT485_0),.clk(gclk));
	jdff dff_A_ggVshsIh6_1(.dout(w_G234_0[1]),.din(w_dff_A_ggVshsIh6_1),.clk(gclk));
	jdff dff_A_89kZRE0r3_2(.dout(w_G234_0[2]),.din(w_dff_A_89kZRE0r3_2),.clk(gclk));
	jdff dff_A_2roPytqy0_1(.dout(w_G221_0[1]),.din(w_dff_A_2roPytqy0_1),.clk(gclk));
	jdff dff_A_yCpBk0Y09_1(.dout(w_dff_A_2roPytqy0_1),.din(w_dff_A_yCpBk0Y09_1),.clk(gclk));
	jdff dff_A_sv65aGNS4_1(.dout(w_n216_0[1]),.din(w_dff_A_sv65aGNS4_1),.clk(gclk));
	jdff dff_B_UGeduBdz0_1(.din(n215),.dout(w_dff_B_UGeduBdz0_1),.clk(gclk));
	jdff dff_B_CkLetjez8_1(.din(w_dff_B_UGeduBdz0_1),.dout(w_dff_B_CkLetjez8_1),.clk(gclk));
	jdff dff_B_kUSsOW6B4_1(.din(w_dff_B_CkLetjez8_1),.dout(w_dff_B_kUSsOW6B4_1),.clk(gclk));
	jdff dff_A_ZHkqUpbp4_0(.dout(w_n107_0[0]),.din(w_dff_A_ZHkqUpbp4_0),.clk(gclk));
	jdff dff_A_4k2uxTUi5_0(.dout(w_dff_A_ZHkqUpbp4_0),.din(w_dff_A_4k2uxTUi5_0),.clk(gclk));
	jdff dff_A_Hc370YHl1_0(.dout(w_dff_A_4k2uxTUi5_0),.din(w_dff_A_Hc370YHl1_0),.clk(gclk));
	jdff dff_A_KgxHdDWL2_0(.dout(w_dff_A_Hc370YHl1_0),.din(w_dff_A_KgxHdDWL2_0),.clk(gclk));
	jdff dff_A_JZJ5cXPt2_0(.dout(w_dff_A_KgxHdDWL2_0),.din(w_dff_A_JZJ5cXPt2_0),.clk(gclk));
	jdff dff_A_dTumLa988_0(.dout(w_dff_A_JZJ5cXPt2_0),.din(w_dff_A_dTumLa988_0),.clk(gclk));
	jdff dff_A_EvNMH0Mw6_0(.dout(w_dff_A_dTumLa988_0),.din(w_dff_A_EvNMH0Mw6_0),.clk(gclk));
	jdff dff_A_b34TpyAV9_0(.dout(w_dff_A_EvNMH0Mw6_0),.din(w_dff_A_b34TpyAV9_0),.clk(gclk));
	jdff dff_A_E3sWM7kP7_0(.dout(w_dff_A_b34TpyAV9_0),.din(w_dff_A_E3sWM7kP7_0),.clk(gclk));
	jdff dff_A_f7xTYwhE4_0(.dout(w_dff_A_E3sWM7kP7_0),.din(w_dff_A_f7xTYwhE4_0),.clk(gclk));
	jdff dff_A_hdnF33qb9_0(.dout(w_dff_A_f7xTYwhE4_0),.din(w_dff_A_hdnF33qb9_0),.clk(gclk));
	jdff dff_A_g1ORjDxT3_0(.dout(w_dff_A_hdnF33qb9_0),.din(w_dff_A_g1ORjDxT3_0),.clk(gclk));
	jdff dff_B_FO9vK7AP2_1(.din(n104),.dout(w_dff_B_FO9vK7AP2_1),.clk(gclk));
	jdff dff_A_PnlwhtQw8_0(.dout(w_G125_0[0]),.din(w_dff_A_PnlwhtQw8_0),.clk(gclk));
	jdff dff_A_JZ5m6VnO8_0(.dout(w_dff_A_PnlwhtQw8_0),.din(w_dff_A_JZ5m6VnO8_0),.clk(gclk));
	jdff dff_A_WGfH91Yx6_0(.dout(w_dff_A_JZ5m6VnO8_0),.din(w_dff_A_WGfH91Yx6_0),.clk(gclk));
	jdff dff_A_xGpjIgIh5_0(.dout(w_dff_A_WGfH91Yx6_0),.din(w_dff_A_xGpjIgIh5_0),.clk(gclk));
	jdff dff_A_zKsRrzPj3_0(.dout(w_dff_A_xGpjIgIh5_0),.din(w_dff_A_zKsRrzPj3_0),.clk(gclk));
	jdff dff_A_WDVkUHBz1_0(.dout(w_dff_A_zKsRrzPj3_0),.din(w_dff_A_WDVkUHBz1_0),.clk(gclk));
	jdff dff_A_pi9Y8krL5_0(.dout(w_dff_A_WDVkUHBz1_0),.din(w_dff_A_pi9Y8krL5_0),.clk(gclk));
	jdff dff_A_486T9eco4_0(.dout(w_dff_A_pi9Y8krL5_0),.din(w_dff_A_486T9eco4_0),.clk(gclk));
	jdff dff_A_aqGOVTYM0_0(.dout(w_dff_A_486T9eco4_0),.din(w_dff_A_aqGOVTYM0_0),.clk(gclk));
	jdff dff_A_P29qcHQQ6_0(.dout(w_dff_A_aqGOVTYM0_0),.din(w_dff_A_P29qcHQQ6_0),.clk(gclk));
	jdff dff_A_ArXJfFfX1_0(.dout(w_dff_A_P29qcHQQ6_0),.din(w_dff_A_ArXJfFfX1_0),.clk(gclk));
	jdff dff_A_ZQxUeYFV5_0(.dout(w_dff_A_ArXJfFfX1_0),.din(w_dff_A_ZQxUeYFV5_0),.clk(gclk));
	jdff dff_A_Yo8kznD37_1(.dout(w_G125_0[1]),.din(w_dff_A_Yo8kznD37_1),.clk(gclk));
	jdff dff_A_nAprNfw33_1(.dout(w_dff_A_Yo8kznD37_1),.din(w_dff_A_nAprNfw33_1),.clk(gclk));
	jdff dff_B_Cs8bBDdu8_2(.din(G224),.dout(w_dff_B_Cs8bBDdu8_2),.clk(gclk));
	jdff dff_A_ISIF9isV8_0(.dout(w_n103_0[0]),.din(w_dff_A_ISIF9isV8_0),.clk(gclk));
	jdff dff_A_aIhkJofu7_0(.dout(w_dff_A_ISIF9isV8_0),.din(w_dff_A_aIhkJofu7_0),.clk(gclk));
	jdff dff_A_lNHD9F7Q7_0(.dout(w_dff_A_aIhkJofu7_0),.din(w_dff_A_lNHD9F7Q7_0),.clk(gclk));
	jdff dff_A_SECMuhex4_0(.dout(w_dff_A_lNHD9F7Q7_0),.din(w_dff_A_SECMuhex4_0),.clk(gclk));
	jdff dff_A_hNNPIpT05_0(.dout(w_dff_A_SECMuhex4_0),.din(w_dff_A_hNNPIpT05_0),.clk(gclk));
	jdff dff_A_A4c9U7eH1_0(.dout(w_dff_A_hNNPIpT05_0),.din(w_dff_A_A4c9U7eH1_0),.clk(gclk));
	jdff dff_A_C4HrPy779_0(.dout(w_dff_A_A4c9U7eH1_0),.din(w_dff_A_C4HrPy779_0),.clk(gclk));
	jdff dff_A_EngtZWI63_0(.dout(w_dff_A_C4HrPy779_0),.din(w_dff_A_EngtZWI63_0),.clk(gclk));
	jdff dff_A_guHP7NST5_0(.dout(w_dff_A_EngtZWI63_0),.din(w_dff_A_guHP7NST5_0),.clk(gclk));
	jdff dff_A_jh3iVW3D0_0(.dout(w_dff_A_guHP7NST5_0),.din(w_dff_A_jh3iVW3D0_0),.clk(gclk));
	jdff dff_A_ATqskvdz9_0(.dout(w_dff_A_jh3iVW3D0_0),.din(w_dff_A_ATqskvdz9_0),.clk(gclk));
	jdff dff_A_hCN9fHM94_0(.dout(w_dff_A_ATqskvdz9_0),.din(w_dff_A_hCN9fHM94_0),.clk(gclk));
	jdff dff_A_wN0Zf4xK3_0(.dout(w_dff_A_hCN9fHM94_0),.din(w_dff_A_wN0Zf4xK3_0),.clk(gclk));
	jdff dff_B_dnr6vzjO6_1(.din(n99),.dout(w_dff_B_dnr6vzjO6_1),.clk(gclk));
	jdff dff_A_MDB8iETe1_0(.dout(w_G107_0[0]),.din(w_dff_A_MDB8iETe1_0),.clk(gclk));
	jdff dff_A_ksRPY3xq2_0(.dout(w_dff_A_MDB8iETe1_0),.din(w_dff_A_ksRPY3xq2_0),.clk(gclk));
	jdff dff_A_hWjPEOkq3_0(.dout(w_dff_A_ksRPY3xq2_0),.din(w_dff_A_hWjPEOkq3_0),.clk(gclk));
	jdff dff_A_xpQzUwJK8_0(.dout(w_dff_A_hWjPEOkq3_0),.din(w_dff_A_xpQzUwJK8_0),.clk(gclk));
	jdff dff_A_h3pQ6Ceu2_0(.dout(w_dff_A_xpQzUwJK8_0),.din(w_dff_A_h3pQ6Ceu2_0),.clk(gclk));
	jdff dff_A_APAWADrK7_0(.dout(w_dff_A_h3pQ6Ceu2_0),.din(w_dff_A_APAWADrK7_0),.clk(gclk));
	jdff dff_A_y1czvHnx1_0(.dout(w_dff_A_APAWADrK7_0),.din(w_dff_A_y1czvHnx1_0),.clk(gclk));
	jdff dff_A_NO4oX8BS0_0(.dout(w_dff_A_y1czvHnx1_0),.din(w_dff_A_NO4oX8BS0_0),.clk(gclk));
	jdff dff_A_lahtR6aK2_0(.dout(w_dff_A_NO4oX8BS0_0),.din(w_dff_A_lahtR6aK2_0),.clk(gclk));
	jdff dff_A_OjVz81K20_0(.dout(w_dff_A_lahtR6aK2_0),.din(w_dff_A_OjVz81K20_0),.clk(gclk));
	jdff dff_A_ix3vRjwt2_0(.dout(w_dff_A_OjVz81K20_0),.din(w_dff_A_ix3vRjwt2_0),.clk(gclk));
	jdff dff_A_II0a2sMc3_0(.dout(w_dff_A_ix3vRjwt2_0),.din(w_dff_A_II0a2sMc3_0),.clk(gclk));
	jdff dff_A_o5GIHIjc2_0(.dout(w_G104_0[0]),.din(w_dff_A_o5GIHIjc2_0),.clk(gclk));
	jdff dff_A_yMyujAxK1_0(.dout(w_dff_A_o5GIHIjc2_0),.din(w_dff_A_yMyujAxK1_0),.clk(gclk));
	jdff dff_A_eouqoC498_0(.dout(w_dff_A_yMyujAxK1_0),.din(w_dff_A_eouqoC498_0),.clk(gclk));
	jdff dff_A_DyTSIePs4_0(.dout(w_dff_A_eouqoC498_0),.din(w_dff_A_DyTSIePs4_0),.clk(gclk));
	jdff dff_A_gZPj3fv32_0(.dout(w_dff_A_DyTSIePs4_0),.din(w_dff_A_gZPj3fv32_0),.clk(gclk));
	jdff dff_A_dxVpsDi56_0(.dout(w_dff_A_gZPj3fv32_0),.din(w_dff_A_dxVpsDi56_0),.clk(gclk));
	jdff dff_A_fi8J9VmA6_0(.dout(w_dff_A_dxVpsDi56_0),.din(w_dff_A_fi8J9VmA6_0),.clk(gclk));
	jdff dff_A_o7Kn8B2X4_0(.dout(w_dff_A_fi8J9VmA6_0),.din(w_dff_A_o7Kn8B2X4_0),.clk(gclk));
	jdff dff_A_z5woJNMy4_0(.dout(w_dff_A_o7Kn8B2X4_0),.din(w_dff_A_z5woJNMy4_0),.clk(gclk));
	jdff dff_A_TWFjMZ5A5_0(.dout(w_dff_A_z5woJNMy4_0),.din(w_dff_A_TWFjMZ5A5_0),.clk(gclk));
	jdff dff_A_7wFpHwdV9_0(.dout(w_dff_A_TWFjMZ5A5_0),.din(w_dff_A_7wFpHwdV9_0),.clk(gclk));
	jdff dff_A_JUN6cAtx4_0(.dout(w_dff_A_7wFpHwdV9_0),.din(w_dff_A_JUN6cAtx4_0),.clk(gclk));
	jdff dff_A_p2qQeJRt6_1(.dout(w_G104_0[1]),.din(w_dff_A_p2qQeJRt6_1),.clk(gclk));
	jdff dff_A_L3g0NJor4_1(.dout(w_dff_A_p2qQeJRt6_1),.din(w_dff_A_L3g0NJor4_1),.clk(gclk));
	jdff dff_A_Ddh5DIGQ4_1(.dout(w_G122_1[1]),.din(w_dff_A_Ddh5DIGQ4_1),.clk(gclk));
	jdff dff_A_k3DB6E8w3_1(.dout(w_G122_0[1]),.din(w_dff_A_k3DB6E8w3_1),.clk(gclk));
	jdff dff_A_v1JzMh499_1(.dout(w_dff_A_k3DB6E8w3_1),.din(w_dff_A_v1JzMh499_1),.clk(gclk));
	jdff dff_A_r1xBo5yf9_1(.dout(w_dff_A_v1JzMh499_1),.din(w_dff_A_r1xBo5yf9_1),.clk(gclk));
	jdff dff_A_X5HSDzXy6_1(.dout(w_dff_A_r1xBo5yf9_1),.din(w_dff_A_X5HSDzXy6_1),.clk(gclk));
	jdff dff_A_AMZjBZ5Q2_1(.dout(w_dff_A_X5HSDzXy6_1),.din(w_dff_A_AMZjBZ5Q2_1),.clk(gclk));
	jdff dff_A_kKuEV2AB0_1(.dout(w_dff_A_AMZjBZ5Q2_1),.din(w_dff_A_kKuEV2AB0_1),.clk(gclk));
	jdff dff_A_BVnIvebr8_1(.dout(w_dff_A_kKuEV2AB0_1),.din(w_dff_A_BVnIvebr8_1),.clk(gclk));
	jdff dff_A_YVVRTht70_1(.dout(w_dff_A_BVnIvebr8_1),.din(w_dff_A_YVVRTht70_1),.clk(gclk));
	jdff dff_A_wobpuE6y1_1(.dout(w_dff_A_YVVRTht70_1),.din(w_dff_A_wobpuE6y1_1),.clk(gclk));
	jdff dff_A_2Z629HSC4_1(.dout(w_dff_A_wobpuE6y1_1),.din(w_dff_A_2Z629HSC4_1),.clk(gclk));
	jdff dff_A_SIogjVJG3_1(.dout(w_dff_A_2Z629HSC4_1),.din(w_dff_A_SIogjVJG3_1),.clk(gclk));
	jdff dff_A_w6arXA8v7_1(.dout(w_dff_A_SIogjVJG3_1),.din(w_dff_A_w6arXA8v7_1),.clk(gclk));
	jdff dff_A_Ec8Ld3O35_2(.dout(w_G122_0[2]),.din(w_dff_A_Ec8Ld3O35_2),.clk(gclk));
	jdff dff_A_y6kskGDT1_1(.dout(w_G110_1[1]),.din(w_dff_A_y6kskGDT1_1),.clk(gclk));
	jdff dff_A_YUUqTcvI8_1(.dout(w_dff_A_y6kskGDT1_1),.din(w_dff_A_YUUqTcvI8_1),.clk(gclk));
	jdff dff_A_eKSMDSod0_1(.dout(w_dff_A_YUUqTcvI8_1),.din(w_dff_A_eKSMDSod0_1),.clk(gclk));
	jdff dff_A_MJweIFhr8_1(.dout(w_dff_A_eKSMDSod0_1),.din(w_dff_A_MJweIFhr8_1),.clk(gclk));
	jdff dff_A_aclXEIyw0_1(.dout(w_dff_A_MJweIFhr8_1),.din(w_dff_A_aclXEIyw0_1),.clk(gclk));
	jdff dff_A_BRAQ6cGg2_1(.dout(w_G110_0[1]),.din(w_dff_A_BRAQ6cGg2_1),.clk(gclk));
	jdff dff_A_THMf1PB55_1(.dout(w_dff_A_BRAQ6cGg2_1),.din(w_dff_A_THMf1PB55_1),.clk(gclk));
	jdff dff_A_ZWW6Y2wf2_1(.dout(w_dff_A_THMf1PB55_1),.din(w_dff_A_ZWW6Y2wf2_1),.clk(gclk));
	jdff dff_A_lVBgeQoh8_1(.dout(w_dff_A_ZWW6Y2wf2_1),.din(w_dff_A_lVBgeQoh8_1),.clk(gclk));
	jdff dff_A_9rMQASy27_1(.dout(w_dff_A_lVBgeQoh8_1),.din(w_dff_A_9rMQASy27_1),.clk(gclk));
	jdff dff_A_x4qXe0lD9_1(.dout(w_dff_A_9rMQASy27_1),.din(w_dff_A_x4qXe0lD9_1),.clk(gclk));
	jdff dff_A_j1Zh2E308_1(.dout(w_dff_A_x4qXe0lD9_1),.din(w_dff_A_j1Zh2E308_1),.clk(gclk));
	jdff dff_A_mh9vj8Iq4_1(.dout(w_dff_A_j1Zh2E308_1),.din(w_dff_A_mh9vj8Iq4_1),.clk(gclk));
	jdff dff_A_xdJPCwPR5_1(.dout(w_dff_A_mh9vj8Iq4_1),.din(w_dff_A_xdJPCwPR5_1),.clk(gclk));
	jdff dff_A_nyPTpRkc4_1(.dout(w_dff_A_xdJPCwPR5_1),.din(w_dff_A_nyPTpRkc4_1),.clk(gclk));
	jdff dff_A_QmhLiQbM1_1(.dout(w_dff_A_nyPTpRkc4_1),.din(w_dff_A_QmhLiQbM1_1),.clk(gclk));
	jdff dff_A_DssgHyMX5_1(.dout(w_dff_A_QmhLiQbM1_1),.din(w_dff_A_DssgHyMX5_1),.clk(gclk));
	jdff dff_A_XuI57YRK1_1(.dout(w_n70_0[1]),.din(w_dff_A_XuI57YRK1_1),.clk(gclk));
	jdff dff_A_FWBCGhG24_1(.dout(w_dff_A_XuI57YRK1_1),.din(w_dff_A_FWBCGhG24_1),.clk(gclk));
	jdff dff_A_KmRdp1rA2_1(.dout(w_dff_A_FWBCGhG24_1),.din(w_dff_A_KmRdp1rA2_1),.clk(gclk));
	jdff dff_A_t4wq9cUJ4_1(.dout(w_dff_A_KmRdp1rA2_1),.din(w_dff_A_t4wq9cUJ4_1),.clk(gclk));
	jdff dff_A_iqaD8r9z4_1(.dout(w_n97_0[1]),.din(w_dff_A_iqaD8r9z4_1),.clk(gclk));
	jdff dff_A_lgzrQ1LR2_1(.dout(w_dff_A_iqaD8r9z4_1),.din(w_dff_A_lgzrQ1LR2_1),.clk(gclk));
	jdff dff_A_9tvp1E123_1(.dout(w_dff_A_lgzrQ1LR2_1),.din(w_dff_A_9tvp1E123_1),.clk(gclk));
	jdff dff_A_VhmM6P478_1(.dout(w_dff_A_9tvp1E123_1),.din(w_dff_A_VhmM6P478_1),.clk(gclk));
	jdff dff_A_snbUpo1Z0_0(.dout(w_n95_0[0]),.din(w_dff_A_snbUpo1Z0_0),.clk(gclk));
	jdff dff_A_D50ukLQQ6_0(.dout(w_dff_A_snbUpo1Z0_0),.din(w_dff_A_D50ukLQQ6_0),.clk(gclk));
	jdff dff_A_g6rrSMku3_0(.dout(w_dff_A_D50ukLQQ6_0),.din(w_dff_A_g6rrSMku3_0),.clk(gclk));
	jdff dff_A_Hj9aZnJU9_0(.dout(w_dff_A_g6rrSMku3_0),.din(w_dff_A_Hj9aZnJU9_0),.clk(gclk));
	jdff dff_A_pp7OSwDu3_0(.dout(w_dff_A_Hj9aZnJU9_0),.din(w_dff_A_pp7OSwDu3_0),.clk(gclk));
	jdff dff_A_LIv5uAeB7_1(.dout(w_n95_0[1]),.din(w_dff_A_LIv5uAeB7_1),.clk(gclk));
	jdff dff_A_Tg4ZrqNW5_1(.dout(w_dff_A_LIv5uAeB7_1),.din(w_dff_A_Tg4ZrqNW5_1),.clk(gclk));
	jdff dff_A_nCCG4xHc5_1(.dout(w_dff_A_Tg4ZrqNW5_1),.din(w_dff_A_nCCG4xHc5_1),.clk(gclk));
	jdff dff_A_oqHOa6lF5_1(.dout(w_dff_A_nCCG4xHc5_1),.din(w_dff_A_oqHOa6lF5_1),.clk(gclk));
	jdff dff_A_5I2AiDSb2_1(.dout(w_dff_A_oqHOa6lF5_1),.din(w_dff_A_5I2AiDSb2_1),.clk(gclk));
	jdff dff_A_UFa8GZ8p3_2(.dout(w_G902_3[2]),.din(w_dff_A_UFa8GZ8p3_2),.clk(gclk));
	jdff dff_A_xiag4azV4_2(.dout(w_dff_A_UFa8GZ8p3_2),.din(w_dff_A_xiag4azV4_2),.clk(gclk));
	jdff dff_A_qjYLtkfG3_2(.dout(w_dff_A_xiag4azV4_2),.din(w_dff_A_qjYLtkfG3_2),.clk(gclk));
	jdff dff_A_nDJp6hBW3_2(.dout(w_dff_A_qjYLtkfG3_2),.din(w_dff_A_nDJp6hBW3_2),.clk(gclk));
	jdff dff_A_paufcRPd3_2(.dout(w_dff_A_nDJp6hBW3_2),.din(w_dff_A_paufcRPd3_2),.clk(gclk));
	jdff dff_A_4i9eyJnQ9_2(.dout(w_dff_A_paufcRPd3_2),.din(w_dff_A_4i9eyJnQ9_2),.clk(gclk));
	jdff dff_A_QRdg40aF4_2(.dout(w_dff_A_4i9eyJnQ9_2),.din(w_dff_A_QRdg40aF4_2),.clk(gclk));
	jdff dff_A_WHE8BckL9_1(.dout(w_G214_0[1]),.din(w_dff_A_WHE8BckL9_1),.clk(gclk));
	jdff dff_A_CWymT7yq3_0(.dout(w_n90_0[0]),.din(w_dff_A_CWymT7yq3_0),.clk(gclk));
	jdff dff_A_bO0UbUXO9_0(.dout(w_dff_A_CWymT7yq3_0),.din(w_dff_A_bO0UbUXO9_0),.clk(gclk));
	jdff dff_A_RaerdxAK0_0(.dout(w_dff_A_bO0UbUXO9_0),.din(w_dff_A_RaerdxAK0_0),.clk(gclk));
	jdff dff_A_rjQlVEfz9_0(.dout(w_dff_A_RaerdxAK0_0),.din(w_dff_A_rjQlVEfz9_0),.clk(gclk));
	jdff dff_A_90p0szhD7_0(.dout(w_dff_A_rjQlVEfz9_0),.din(w_dff_A_90p0szhD7_0),.clk(gclk));
	jdff dff_A_HNI1iM831_0(.dout(w_dff_A_90p0szhD7_0),.din(w_dff_A_HNI1iM831_0),.clk(gclk));
	jdff dff_A_Hh7OsBkk2_0(.dout(w_dff_A_HNI1iM831_0),.din(w_dff_A_Hh7OsBkk2_0),.clk(gclk));
	jdff dff_A_9F4TfS4E5_0(.dout(w_dff_A_Hh7OsBkk2_0),.din(w_dff_A_9F4TfS4E5_0),.clk(gclk));
	jdff dff_A_OoH6eD4R6_0(.dout(w_dff_A_9F4TfS4E5_0),.din(w_dff_A_OoH6eD4R6_0),.clk(gclk));
	jdff dff_A_bZCrDLAh8_0(.dout(w_dff_A_OoH6eD4R6_0),.din(w_dff_A_bZCrDLAh8_0),.clk(gclk));
	jdff dff_A_O49NUb3s5_0(.dout(w_dff_A_bZCrDLAh8_0),.din(w_dff_A_O49NUb3s5_0),.clk(gclk));
	jdff dff_A_MCYmCCnC0_0(.dout(w_dff_A_O49NUb3s5_0),.din(w_dff_A_MCYmCCnC0_0),.clk(gclk));
	jdff dff_A_h0Dffoh04_0(.dout(w_G953_1[0]),.din(w_dff_A_h0Dffoh04_0),.clk(gclk));
	jdff dff_A_8nKWwOI41_0(.dout(w_dff_A_h0Dffoh04_0),.din(w_dff_A_8nKWwOI41_0),.clk(gclk));
	jdff dff_A_NSKguIuh7_0(.dout(w_dff_A_8nKWwOI41_0),.din(w_dff_A_NSKguIuh7_0),.clk(gclk));
	jdff dff_A_4naNH1m66_0(.dout(w_dff_A_NSKguIuh7_0),.din(w_dff_A_4naNH1m66_0),.clk(gclk));
	jdff dff_A_4vTOr4r51_0(.dout(w_dff_A_4naNH1m66_0),.din(w_dff_A_4vTOr4r51_0),.clk(gclk));
	jdff dff_A_aeqoslnv0_0(.dout(w_dff_A_4vTOr4r51_0),.din(w_dff_A_aeqoslnv0_0),.clk(gclk));
	jdff dff_A_qhB5ACh29_0(.dout(w_dff_A_aeqoslnv0_0),.din(w_dff_A_qhB5ACh29_0),.clk(gclk));
	jdff dff_A_rIfMH1le8_0(.dout(w_dff_A_qhB5ACh29_0),.din(w_dff_A_rIfMH1le8_0),.clk(gclk));
	jdff dff_A_QTILc4YB6_0(.dout(w_dff_A_rIfMH1le8_0),.din(w_dff_A_QTILc4YB6_0),.clk(gclk));
	jdff dff_A_brTqkjB06_0(.dout(w_dff_A_QTILc4YB6_0),.din(w_dff_A_brTqkjB06_0),.clk(gclk));
	jdff dff_A_w6mxQNlP6_0(.dout(w_dff_A_brTqkjB06_0),.din(w_dff_A_w6mxQNlP6_0),.clk(gclk));
	jdff dff_A_N8483xR91_0(.dout(w_dff_A_w6mxQNlP6_0),.din(w_dff_A_N8483xR91_0),.clk(gclk));
	jdff dff_A_cB1mUdX04_1(.dout(w_G953_0[1]),.din(w_dff_A_cB1mUdX04_1),.clk(gclk));
	jdff dff_A_SEF5qUbG5_1(.dout(w_dff_A_cB1mUdX04_1),.din(w_dff_A_SEF5qUbG5_1),.clk(gclk));
	jdff dff_A_mwoS1c6A6_1(.dout(w_dff_A_SEF5qUbG5_1),.din(w_dff_A_mwoS1c6A6_1),.clk(gclk));
	jdff dff_A_rGZpNTE14_1(.dout(w_dff_A_mwoS1c6A6_1),.din(w_dff_A_rGZpNTE14_1),.clk(gclk));
	jdff dff_A_lY0cgKZ79_1(.dout(w_dff_A_rGZpNTE14_1),.din(w_dff_A_lY0cgKZ79_1),.clk(gclk));
	jdff dff_A_sTKLxUYb7_1(.dout(w_dff_A_lY0cgKZ79_1),.din(w_dff_A_sTKLxUYb7_1),.clk(gclk));
	jdff dff_A_rmas8ajd6_1(.dout(w_dff_A_sTKLxUYb7_1),.din(w_dff_A_rmas8ajd6_1),.clk(gclk));
	jdff dff_A_qVDZP92s6_1(.dout(w_dff_A_rmas8ajd6_1),.din(w_dff_A_qVDZP92s6_1),.clk(gclk));
	jdff dff_A_TJTqvTeT9_1(.dout(w_dff_A_qVDZP92s6_1),.din(w_dff_A_TJTqvTeT9_1),.clk(gclk));
	jdff dff_A_dNVObq0U6_1(.dout(w_dff_A_TJTqvTeT9_1),.din(w_dff_A_dNVObq0U6_1),.clk(gclk));
	jdff dff_A_3dbCYNXb1_1(.dout(w_dff_A_dNVObq0U6_1),.din(w_dff_A_3dbCYNXb1_1),.clk(gclk));
	jdff dff_A_1alljOBI3_1(.dout(w_dff_A_3dbCYNXb1_1),.din(w_dff_A_1alljOBI3_1),.clk(gclk));
	jdff dff_A_8nD2dtlC4_1(.dout(w_dff_A_1alljOBI3_1),.din(w_dff_A_8nD2dtlC4_1),.clk(gclk));
	jdff dff_A_CUgDdtaZ2_1(.dout(w_dff_A_8nD2dtlC4_1),.din(w_dff_A_CUgDdtaZ2_1),.clk(gclk));
	jdff dff_A_v8bqlD7a2_1(.dout(w_dff_A_CUgDdtaZ2_1),.din(w_dff_A_v8bqlD7a2_1),.clk(gclk));
	jdff dff_A_3a2JHqZY5_2(.dout(w_G953_0[2]),.din(w_dff_A_3a2JHqZY5_2),.clk(gclk));
	jdff dff_A_VhO82LPz1_2(.dout(w_dff_A_3a2JHqZY5_2),.din(w_dff_A_VhO82LPz1_2),.clk(gclk));
	jdff dff_A_0YJ11Z8j2_2(.dout(w_dff_A_VhO82LPz1_2),.din(w_dff_A_0YJ11Z8j2_2),.clk(gclk));
	jdff dff_A_bZeC2siw3_2(.dout(w_dff_A_0YJ11Z8j2_2),.din(w_dff_A_bZeC2siw3_2),.clk(gclk));
	jdff dff_A_XlG72CDe4_2(.dout(w_dff_A_bZeC2siw3_2),.din(w_dff_A_XlG72CDe4_2),.clk(gclk));
	jdff dff_A_7mUSggM42_2(.dout(w_dff_A_XlG72CDe4_2),.din(w_dff_A_7mUSggM42_2),.clk(gclk));
	jdff dff_A_2AgwEJ7B3_2(.dout(w_dff_A_7mUSggM42_2),.din(w_dff_A_2AgwEJ7B3_2),.clk(gclk));
	jdff dff_A_VgXDAfB17_2(.dout(w_dff_A_2AgwEJ7B3_2),.din(w_dff_A_VgXDAfB17_2),.clk(gclk));
	jdff dff_A_CIoGP6cw2_2(.dout(w_dff_A_VgXDAfB17_2),.din(w_dff_A_CIoGP6cw2_2),.clk(gclk));
	jdff dff_A_NXFnoskI5_2(.dout(w_dff_A_CIoGP6cw2_2),.din(w_dff_A_NXFnoskI5_2),.clk(gclk));
	jdff dff_A_moeBF56a3_2(.dout(w_dff_A_NXFnoskI5_2),.din(w_dff_A_moeBF56a3_2),.clk(gclk));
	jdff dff_A_oEcTbdz11_2(.dout(w_dff_A_moeBF56a3_2),.din(w_dff_A_oEcTbdz11_2),.clk(gclk));
	jdff dff_A_JhRr7uuN4_2(.dout(w_dff_A_oEcTbdz11_2),.din(w_dff_A_JhRr7uuN4_2),.clk(gclk));
	jdff dff_A_GcbRdbm23_2(.dout(w_dff_A_JhRr7uuN4_2),.din(w_dff_A_GcbRdbm23_2),.clk(gclk));
	jdff dff_A_5XAaL6JI8_2(.dout(w_dff_A_GcbRdbm23_2),.din(w_dff_A_5XAaL6JI8_2),.clk(gclk));
	jdff dff_A_o71ohj0b8_1(.dout(w_G210_0[1]),.din(w_dff_A_o71ohj0b8_1),.clk(gclk));
	jdff dff_A_ZTUYCujP4_0(.dout(w_G101_0[0]),.din(w_dff_A_ZTUYCujP4_0),.clk(gclk));
	jdff dff_A_iCXY3wNZ1_0(.dout(w_dff_A_ZTUYCujP4_0),.din(w_dff_A_iCXY3wNZ1_0),.clk(gclk));
	jdff dff_A_wPhlVCtG5_0(.dout(w_dff_A_iCXY3wNZ1_0),.din(w_dff_A_wPhlVCtG5_0),.clk(gclk));
	jdff dff_A_jig1QCiK7_0(.dout(w_dff_A_wPhlVCtG5_0),.din(w_dff_A_jig1QCiK7_0),.clk(gclk));
	jdff dff_A_gL8JFqHC1_0(.dout(w_dff_A_jig1QCiK7_0),.din(w_dff_A_gL8JFqHC1_0),.clk(gclk));
	jdff dff_A_mn71MHuM9_0(.dout(w_dff_A_gL8JFqHC1_0),.din(w_dff_A_mn71MHuM9_0),.clk(gclk));
	jdff dff_A_F5iUrl6o0_0(.dout(w_dff_A_mn71MHuM9_0),.din(w_dff_A_F5iUrl6o0_0),.clk(gclk));
	jdff dff_A_EkrmMm8i8_0(.dout(w_dff_A_F5iUrl6o0_0),.din(w_dff_A_EkrmMm8i8_0),.clk(gclk));
	jdff dff_A_vMimOC1k9_0(.dout(w_dff_A_EkrmMm8i8_0),.din(w_dff_A_vMimOC1k9_0),.clk(gclk));
	jdff dff_A_KL0o4pkr0_0(.dout(w_dff_A_vMimOC1k9_0),.din(w_dff_A_KL0o4pkr0_0),.clk(gclk));
	jdff dff_A_BD31Yy7l0_0(.dout(w_dff_A_KL0o4pkr0_0),.din(w_dff_A_BD31Yy7l0_0),.clk(gclk));
	jdff dff_A_qpCYztlw5_2(.dout(w_G101_0[2]),.din(w_dff_A_qpCYztlw5_2),.clk(gclk));
	jdff dff_B_Kjj8zeKW6_3(.din(G101),.dout(w_dff_B_Kjj8zeKW6_3),.clk(gclk));
	jdff dff_A_03eJseTV7_1(.dout(w_n84_0[1]),.din(w_dff_A_03eJseTV7_1),.clk(gclk));
	jdff dff_A_RFfJsU3L2_0(.dout(w_G119_0[0]),.din(w_dff_A_RFfJsU3L2_0),.clk(gclk));
	jdff dff_A_NmQBxOPY0_0(.dout(w_dff_A_RFfJsU3L2_0),.din(w_dff_A_NmQBxOPY0_0),.clk(gclk));
	jdff dff_A_DvTUDHWg5_0(.dout(w_dff_A_NmQBxOPY0_0),.din(w_dff_A_DvTUDHWg5_0),.clk(gclk));
	jdff dff_A_DZ3kNWmy3_0(.dout(w_dff_A_DvTUDHWg5_0),.din(w_dff_A_DZ3kNWmy3_0),.clk(gclk));
	jdff dff_A_bBe5pjPZ5_0(.dout(w_dff_A_DZ3kNWmy3_0),.din(w_dff_A_bBe5pjPZ5_0),.clk(gclk));
	jdff dff_A_0HeKcJ4V4_0(.dout(w_dff_A_bBe5pjPZ5_0),.din(w_dff_A_0HeKcJ4V4_0),.clk(gclk));
	jdff dff_A_aPPxyjUa3_0(.dout(w_dff_A_0HeKcJ4V4_0),.din(w_dff_A_aPPxyjUa3_0),.clk(gclk));
	jdff dff_A_RaAq9WJD3_0(.dout(w_dff_A_aPPxyjUa3_0),.din(w_dff_A_RaAq9WJD3_0),.clk(gclk));
	jdff dff_A_JThiMuv48_0(.dout(w_dff_A_RaAq9WJD3_0),.din(w_dff_A_JThiMuv48_0),.clk(gclk));
	jdff dff_A_hp8YCXT01_0(.dout(w_dff_A_JThiMuv48_0),.din(w_dff_A_hp8YCXT01_0),.clk(gclk));
	jdff dff_A_o068Pd0r7_0(.dout(w_dff_A_hp8YCXT01_0),.din(w_dff_A_o068Pd0r7_0),.clk(gclk));
	jdff dff_A_dwW8yMJR4_0(.dout(w_dff_A_o068Pd0r7_0),.din(w_dff_A_dwW8yMJR4_0),.clk(gclk));
	jdff dff_A_fBT6QHjD8_0(.dout(w_G116_0[0]),.din(w_dff_A_fBT6QHjD8_0),.clk(gclk));
	jdff dff_A_r6ZIXBe10_0(.dout(w_dff_A_fBT6QHjD8_0),.din(w_dff_A_r6ZIXBe10_0),.clk(gclk));
	jdff dff_A_RQkaPbBk4_0(.dout(w_dff_A_r6ZIXBe10_0),.din(w_dff_A_RQkaPbBk4_0),.clk(gclk));
	jdff dff_A_ZoSmQTxH3_0(.dout(w_dff_A_RQkaPbBk4_0),.din(w_dff_A_ZoSmQTxH3_0),.clk(gclk));
	jdff dff_A_VCVnypZW6_0(.dout(w_dff_A_ZoSmQTxH3_0),.din(w_dff_A_VCVnypZW6_0),.clk(gclk));
	jdff dff_A_8Bo9Hc4X8_0(.dout(w_dff_A_VCVnypZW6_0),.din(w_dff_A_8Bo9Hc4X8_0),.clk(gclk));
	jdff dff_A_uUoghMSM2_0(.dout(w_dff_A_8Bo9Hc4X8_0),.din(w_dff_A_uUoghMSM2_0),.clk(gclk));
	jdff dff_A_qjS0guJK4_0(.dout(w_dff_A_uUoghMSM2_0),.din(w_dff_A_qjS0guJK4_0),.clk(gclk));
	jdff dff_A_Z6StphLR2_0(.dout(w_dff_A_qjS0guJK4_0),.din(w_dff_A_Z6StphLR2_0),.clk(gclk));
	jdff dff_A_FUBdNWPA0_0(.dout(w_dff_A_Z6StphLR2_0),.din(w_dff_A_FUBdNWPA0_0),.clk(gclk));
	jdff dff_A_kJRBKz5K4_0(.dout(w_dff_A_FUBdNWPA0_0),.din(w_dff_A_kJRBKz5K4_0),.clk(gclk));
	jdff dff_A_ZkCocvNM8_0(.dout(w_dff_A_kJRBKz5K4_0),.din(w_dff_A_ZkCocvNM8_0),.clk(gclk));
	jdff dff_A_JB0yltDU4_0(.dout(w_G113_0[0]),.din(w_dff_A_JB0yltDU4_0),.clk(gclk));
	jdff dff_A_Hih7WZBh5_0(.dout(w_dff_A_JB0yltDU4_0),.din(w_dff_A_Hih7WZBh5_0),.clk(gclk));
	jdff dff_A_z6WDJsky7_0(.dout(w_dff_A_Hih7WZBh5_0),.din(w_dff_A_z6WDJsky7_0),.clk(gclk));
	jdff dff_A_r0EMzGvt8_0(.dout(w_dff_A_z6WDJsky7_0),.din(w_dff_A_r0EMzGvt8_0),.clk(gclk));
	jdff dff_A_oHVSIxFd0_0(.dout(w_dff_A_r0EMzGvt8_0),.din(w_dff_A_oHVSIxFd0_0),.clk(gclk));
	jdff dff_A_vMm4ViDN6_0(.dout(w_dff_A_oHVSIxFd0_0),.din(w_dff_A_vMm4ViDN6_0),.clk(gclk));
	jdff dff_A_vHkAoap27_0(.dout(w_dff_A_vMm4ViDN6_0),.din(w_dff_A_vHkAoap27_0),.clk(gclk));
	jdff dff_A_yqD3fYIL6_0(.dout(w_dff_A_vHkAoap27_0),.din(w_dff_A_yqD3fYIL6_0),.clk(gclk));
	jdff dff_A_LlRkeM6N6_0(.dout(w_dff_A_yqD3fYIL6_0),.din(w_dff_A_LlRkeM6N6_0),.clk(gclk));
	jdff dff_A_AiDsZfnE9_0(.dout(w_dff_A_LlRkeM6N6_0),.din(w_dff_A_AiDsZfnE9_0),.clk(gclk));
	jdff dff_A_4cC0n8LY6_0(.dout(w_dff_A_AiDsZfnE9_0),.din(w_dff_A_4cC0n8LY6_0),.clk(gclk));
	jdff dff_A_J8lUbPxx5_0(.dout(w_dff_A_4cC0n8LY6_0),.din(w_dff_A_J8lUbPxx5_0),.clk(gclk));
	jdff dff_B_6gfZuDbi7_1(.din(n76),.dout(w_dff_B_6gfZuDbi7_1),.clk(gclk));
	jdff dff_A_9eFwGtyh4_0(.dout(w_G146_0[0]),.din(w_dff_A_9eFwGtyh4_0),.clk(gclk));
	jdff dff_A_hdwgpgnO3_0(.dout(w_dff_A_9eFwGtyh4_0),.din(w_dff_A_hdwgpgnO3_0),.clk(gclk));
	jdff dff_A_596yo6Vi2_0(.dout(w_dff_A_hdwgpgnO3_0),.din(w_dff_A_596yo6Vi2_0),.clk(gclk));
	jdff dff_A_j4x7Z8LB3_0(.dout(w_dff_A_596yo6Vi2_0),.din(w_dff_A_j4x7Z8LB3_0),.clk(gclk));
	jdff dff_A_VQFfDJ7K8_0(.dout(w_dff_A_j4x7Z8LB3_0),.din(w_dff_A_VQFfDJ7K8_0),.clk(gclk));
	jdff dff_A_mAbMNXvs3_0(.dout(w_dff_A_VQFfDJ7K8_0),.din(w_dff_A_mAbMNXvs3_0),.clk(gclk));
	jdff dff_A_TmJVRVwT5_0(.dout(w_dff_A_mAbMNXvs3_0),.din(w_dff_A_TmJVRVwT5_0),.clk(gclk));
	jdff dff_A_Ja1R6rpZ0_0(.dout(w_dff_A_TmJVRVwT5_0),.din(w_dff_A_Ja1R6rpZ0_0),.clk(gclk));
	jdff dff_A_nszDdtmS8_0(.dout(w_dff_A_Ja1R6rpZ0_0),.din(w_dff_A_nszDdtmS8_0),.clk(gclk));
	jdff dff_A_XL1cAoy86_0(.dout(w_dff_A_nszDdtmS8_0),.din(w_dff_A_XL1cAoy86_0),.clk(gclk));
	jdff dff_A_PivG70kI5_0(.dout(w_dff_A_XL1cAoy86_0),.din(w_dff_A_PivG70kI5_0),.clk(gclk));
	jdff dff_A_jSIN758f0_0(.dout(w_dff_A_PivG70kI5_0),.din(w_dff_A_jSIN758f0_0),.clk(gclk));
	jdff dff_A_PLIYJFqk0_1(.dout(w_G143_0[1]),.din(w_dff_A_PLIYJFqk0_1),.clk(gclk));
	jdff dff_A_48NzCRVX1_1(.dout(w_dff_A_PLIYJFqk0_1),.din(w_dff_A_48NzCRVX1_1),.clk(gclk));
	jdff dff_A_4eB1vzSh6_1(.dout(w_dff_A_48NzCRVX1_1),.din(w_dff_A_4eB1vzSh6_1),.clk(gclk));
	jdff dff_A_lJ9so47W8_1(.dout(w_dff_A_4eB1vzSh6_1),.din(w_dff_A_lJ9so47W8_1),.clk(gclk));
	jdff dff_A_2Ij2tSQU3_1(.dout(w_dff_A_lJ9so47W8_1),.din(w_dff_A_2Ij2tSQU3_1),.clk(gclk));
	jdff dff_A_dnWcQex08_1(.dout(w_dff_A_2Ij2tSQU3_1),.din(w_dff_A_dnWcQex08_1),.clk(gclk));
	jdff dff_A_Iux8xokn0_1(.dout(w_dff_A_dnWcQex08_1),.din(w_dff_A_Iux8xokn0_1),.clk(gclk));
	jdff dff_A_Xa1wW3WC9_1(.dout(w_dff_A_Iux8xokn0_1),.din(w_dff_A_Xa1wW3WC9_1),.clk(gclk));
	jdff dff_A_Ma8atjKv5_1(.dout(w_dff_A_Xa1wW3WC9_1),.din(w_dff_A_Ma8atjKv5_1),.clk(gclk));
	jdff dff_A_oVoRhqSM1_1(.dout(w_dff_A_Ma8atjKv5_1),.din(w_dff_A_oVoRhqSM1_1),.clk(gclk));
	jdff dff_A_SsHMTVMO1_1(.dout(w_dff_A_oVoRhqSM1_1),.din(w_dff_A_SsHMTVMO1_1),.clk(gclk));
	jdff dff_A_OabsjFqx3_1(.dout(w_dff_A_SsHMTVMO1_1),.din(w_dff_A_OabsjFqx3_1),.clk(gclk));
	jdff dff_A_ew04d99e6_2(.dout(w_G143_0[2]),.din(w_dff_A_ew04d99e6_2),.clk(gclk));
	jdff dff_A_LRvXUAPF7_0(.dout(w_G128_1[0]),.din(w_dff_A_LRvXUAPF7_0),.clk(gclk));
	jdff dff_A_P4TUrj3J0_1(.dout(w_G128_0[1]),.din(w_dff_A_P4TUrj3J0_1),.clk(gclk));
	jdff dff_A_VFoEQOwg3_1(.dout(w_dff_A_P4TUrj3J0_1),.din(w_dff_A_VFoEQOwg3_1),.clk(gclk));
	jdff dff_A_zb5LOJgW4_1(.dout(w_dff_A_VFoEQOwg3_1),.din(w_dff_A_zb5LOJgW4_1),.clk(gclk));
	jdff dff_A_7wRUYp1D7_1(.dout(w_dff_A_zb5LOJgW4_1),.din(w_dff_A_7wRUYp1D7_1),.clk(gclk));
	jdff dff_A_FpzwSYq85_1(.dout(w_dff_A_7wRUYp1D7_1),.din(w_dff_A_FpzwSYq85_1),.clk(gclk));
	jdff dff_A_2ozmdymg6_1(.dout(w_dff_A_FpzwSYq85_1),.din(w_dff_A_2ozmdymg6_1),.clk(gclk));
	jdff dff_A_bunV11Jf6_1(.dout(w_dff_A_2ozmdymg6_1),.din(w_dff_A_bunV11Jf6_1),.clk(gclk));
	jdff dff_A_vMUNhKiV5_1(.dout(w_dff_A_bunV11Jf6_1),.din(w_dff_A_vMUNhKiV5_1),.clk(gclk));
	jdff dff_A_GjTl6uMF1_1(.dout(w_dff_A_vMUNhKiV5_1),.din(w_dff_A_GjTl6uMF1_1),.clk(gclk));
	jdff dff_A_WV88DE9N7_1(.dout(w_dff_A_GjTl6uMF1_1),.din(w_dff_A_WV88DE9N7_1),.clk(gclk));
	jdff dff_A_VLLucF106_1(.dout(w_dff_A_WV88DE9N7_1),.din(w_dff_A_VLLucF106_1),.clk(gclk));
	jdff dff_A_kQaYuDZR3_1(.dout(w_dff_A_VLLucF106_1),.din(w_dff_A_kQaYuDZR3_1),.clk(gclk));
	jdff dff_A_KXZGKMQm0_1(.dout(w_n77_0[1]),.din(w_dff_A_KXZGKMQm0_1),.clk(gclk));
	jdff dff_A_HWVpkStF9_0(.dout(w_G131_0[0]),.din(w_dff_A_HWVpkStF9_0),.clk(gclk));
	jdff dff_A_lEJQRov87_0(.dout(w_dff_A_HWVpkStF9_0),.din(w_dff_A_lEJQRov87_0),.clk(gclk));
	jdff dff_A_GpyikO766_0(.dout(w_dff_A_lEJQRov87_0),.din(w_dff_A_GpyikO766_0),.clk(gclk));
	jdff dff_A_r1sFdeFC2_0(.dout(w_dff_A_GpyikO766_0),.din(w_dff_A_r1sFdeFC2_0),.clk(gclk));
	jdff dff_A_8GxpfENN9_0(.dout(w_dff_A_r1sFdeFC2_0),.din(w_dff_A_8GxpfENN9_0),.clk(gclk));
	jdff dff_A_NMVIQQEQ4_0(.dout(w_dff_A_8GxpfENN9_0),.din(w_dff_A_NMVIQQEQ4_0),.clk(gclk));
	jdff dff_A_81lGVsSg0_0(.dout(w_dff_A_NMVIQQEQ4_0),.din(w_dff_A_81lGVsSg0_0),.clk(gclk));
	jdff dff_A_zV6syvDI7_0(.dout(w_dff_A_81lGVsSg0_0),.din(w_dff_A_zV6syvDI7_0),.clk(gclk));
	jdff dff_A_b4A1Gu0B7_0(.dout(w_dff_A_zV6syvDI7_0),.din(w_dff_A_b4A1Gu0B7_0),.clk(gclk));
	jdff dff_A_RIbDXy913_0(.dout(w_dff_A_b4A1Gu0B7_0),.din(w_dff_A_RIbDXy913_0),.clk(gclk));
	jdff dff_A_4w2dD41U6_0(.dout(w_dff_A_RIbDXy913_0),.din(w_dff_A_4w2dD41U6_0),.clk(gclk));
	jdff dff_A_UxdBwvIm7_0(.dout(w_dff_A_4w2dD41U6_0),.din(w_dff_A_UxdBwvIm7_0),.clk(gclk));
	jdff dff_A_e4gkRgac2_0(.dout(w_G137_0[0]),.din(w_dff_A_e4gkRgac2_0),.clk(gclk));
	jdff dff_A_0kABJPeN4_0(.dout(w_dff_A_e4gkRgac2_0),.din(w_dff_A_0kABJPeN4_0),.clk(gclk));
	jdff dff_A_fPyMpqqX8_0(.dout(w_dff_A_0kABJPeN4_0),.din(w_dff_A_fPyMpqqX8_0),.clk(gclk));
	jdff dff_A_xssdjAiS9_0(.dout(w_dff_A_fPyMpqqX8_0),.din(w_dff_A_xssdjAiS9_0),.clk(gclk));
	jdff dff_A_r7vOCYgc2_0(.dout(w_dff_A_xssdjAiS9_0),.din(w_dff_A_r7vOCYgc2_0),.clk(gclk));
	jdff dff_A_lH6Tg2A75_0(.dout(w_dff_A_r7vOCYgc2_0),.din(w_dff_A_lH6Tg2A75_0),.clk(gclk));
	jdff dff_A_IE0wfjbX8_0(.dout(w_dff_A_lH6Tg2A75_0),.din(w_dff_A_IE0wfjbX8_0),.clk(gclk));
	jdff dff_A_AFQ64MTR9_0(.dout(w_dff_A_IE0wfjbX8_0),.din(w_dff_A_AFQ64MTR9_0),.clk(gclk));
	jdff dff_A_gyiGt1BC9_0(.dout(w_dff_A_AFQ64MTR9_0),.din(w_dff_A_gyiGt1BC9_0),.clk(gclk));
	jdff dff_A_VALhBbBd9_0(.dout(w_dff_A_gyiGt1BC9_0),.din(w_dff_A_VALhBbBd9_0),.clk(gclk));
	jdff dff_A_YExgF0Dl7_0(.dout(w_dff_A_VALhBbBd9_0),.din(w_dff_A_YExgF0Dl7_0),.clk(gclk));
	jdff dff_A_dxOoY1ou1_2(.dout(w_G137_0[2]),.din(w_dff_A_dxOoY1ou1_2),.clk(gclk));
	jdff dff_A_Sb2aoAom9_2(.dout(w_dff_A_dxOoY1ou1_2),.din(w_dff_A_Sb2aoAom9_2),.clk(gclk));
	jdff dff_B_CjQz1sfH8_3(.din(G137),.dout(w_dff_B_CjQz1sfH8_3),.clk(gclk));
	jdff dff_A_t8lApJZ77_0(.dout(w_G134_0[0]),.din(w_dff_A_t8lApJZ77_0),.clk(gclk));
	jdff dff_A_xWUoS5Qy4_0(.dout(w_dff_A_t8lApJZ77_0),.din(w_dff_A_xWUoS5Qy4_0),.clk(gclk));
	jdff dff_A_GO0x0GVu1_0(.dout(w_dff_A_xWUoS5Qy4_0),.din(w_dff_A_GO0x0GVu1_0),.clk(gclk));
	jdff dff_A_MlhHHKkS4_0(.dout(w_dff_A_GO0x0GVu1_0),.din(w_dff_A_MlhHHKkS4_0),.clk(gclk));
	jdff dff_A_et69PjZh9_0(.dout(w_dff_A_MlhHHKkS4_0),.din(w_dff_A_et69PjZh9_0),.clk(gclk));
	jdff dff_A_LEhKMlEW4_0(.dout(w_dff_A_et69PjZh9_0),.din(w_dff_A_LEhKMlEW4_0),.clk(gclk));
	jdff dff_A_yfkd2Jae4_0(.dout(w_dff_A_LEhKMlEW4_0),.din(w_dff_A_yfkd2Jae4_0),.clk(gclk));
	jdff dff_A_GHHk1Mfc7_0(.dout(w_dff_A_yfkd2Jae4_0),.din(w_dff_A_GHHk1Mfc7_0),.clk(gclk));
	jdff dff_A_hGHzXt5B3_0(.dout(w_dff_A_GHHk1Mfc7_0),.din(w_dff_A_hGHzXt5B3_0),.clk(gclk));
	jdff dff_A_ZNmJ56nX8_0(.dout(w_dff_A_hGHzXt5B3_0),.din(w_dff_A_ZNmJ56nX8_0),.clk(gclk));
	jdff dff_A_WTVSMNBA4_0(.dout(w_dff_A_ZNmJ56nX8_0),.din(w_dff_A_WTVSMNBA4_0),.clk(gclk));
	jdff dff_A_3yL4B5kd1_0(.dout(w_dff_A_WTVSMNBA4_0),.din(w_dff_A_3yL4B5kd1_0),.clk(gclk));
	jdff dff_A_ORIxZwkf0_2(.dout(w_dff_A_ycqjFhlk7_0),.din(w_dff_A_ORIxZwkf0_2),.clk(gclk));
	jdff dff_A_ycqjFhlk7_0(.dout(w_dff_A_MpiUFeaL3_0),.din(w_dff_A_ycqjFhlk7_0),.clk(gclk));
	jdff dff_A_MpiUFeaL3_0(.dout(w_dff_A_pOjbguua1_0),.din(w_dff_A_MpiUFeaL3_0),.clk(gclk));
	jdff dff_A_pOjbguua1_0(.dout(w_dff_A_tXrCSyVW4_0),.din(w_dff_A_pOjbguua1_0),.clk(gclk));
	jdff dff_A_tXrCSyVW4_0(.dout(w_dff_A_dHWsy6DF0_0),.din(w_dff_A_tXrCSyVW4_0),.clk(gclk));
	jdff dff_A_dHWsy6DF0_0(.dout(w_dff_A_VI5jphLn7_0),.din(w_dff_A_dHWsy6DF0_0),.clk(gclk));
	jdff dff_A_VI5jphLn7_0(.dout(G3),.din(w_dff_A_VI5jphLn7_0),.clk(gclk));
	jdff dff_A_bKM2r4hu9_2(.dout(w_dff_A_WV8ToBqA8_0),.din(w_dff_A_bKM2r4hu9_2),.clk(gclk));
	jdff dff_A_WV8ToBqA8_0(.dout(w_dff_A_fmigtWPK1_0),.din(w_dff_A_WV8ToBqA8_0),.clk(gclk));
	jdff dff_A_fmigtWPK1_0(.dout(w_dff_A_SSNbB8xX0_0),.din(w_dff_A_fmigtWPK1_0),.clk(gclk));
	jdff dff_A_SSNbB8xX0_0(.dout(w_dff_A_MgTCBivD9_0),.din(w_dff_A_SSNbB8xX0_0),.clk(gclk));
	jdff dff_A_MgTCBivD9_0(.dout(w_dff_A_DqRhxA1J7_0),.din(w_dff_A_MgTCBivD9_0),.clk(gclk));
	jdff dff_A_DqRhxA1J7_0(.dout(w_dff_A_jKIa7hMH7_0),.din(w_dff_A_DqRhxA1J7_0),.clk(gclk));
	jdff dff_A_jKIa7hMH7_0(.dout(G6),.din(w_dff_A_jKIa7hMH7_0),.clk(gclk));
	jdff dff_A_V5YicqZf1_2(.dout(w_dff_A_eRsXNH8k3_0),.din(w_dff_A_V5YicqZf1_2),.clk(gclk));
	jdff dff_A_eRsXNH8k3_0(.dout(w_dff_A_QagbEwuI0_0),.din(w_dff_A_eRsXNH8k3_0),.clk(gclk));
	jdff dff_A_QagbEwuI0_0(.dout(w_dff_A_nUuyKVi23_0),.din(w_dff_A_QagbEwuI0_0),.clk(gclk));
	jdff dff_A_nUuyKVi23_0(.dout(w_dff_A_Pq1YFTcR4_0),.din(w_dff_A_nUuyKVi23_0),.clk(gclk));
	jdff dff_A_Pq1YFTcR4_0(.dout(w_dff_A_WfsOKEuB5_0),.din(w_dff_A_Pq1YFTcR4_0),.clk(gclk));
	jdff dff_A_WfsOKEuB5_0(.dout(w_dff_A_mzd5uUs53_0),.din(w_dff_A_WfsOKEuB5_0),.clk(gclk));
	jdff dff_A_mzd5uUs53_0(.dout(G9),.din(w_dff_A_mzd5uUs53_0),.clk(gclk));
	jdff dff_A_Z87hynQv1_2(.dout(w_dff_A_LPJYAfXf5_0),.din(w_dff_A_Z87hynQv1_2),.clk(gclk));
	jdff dff_A_LPJYAfXf5_0(.dout(w_dff_A_3AWSMHqz1_0),.din(w_dff_A_LPJYAfXf5_0),.clk(gclk));
	jdff dff_A_3AWSMHqz1_0(.dout(w_dff_A_OSD9DhOH8_0),.din(w_dff_A_3AWSMHqz1_0),.clk(gclk));
	jdff dff_A_OSD9DhOH8_0(.dout(w_dff_A_dDXVwRUp2_0),.din(w_dff_A_OSD9DhOH8_0),.clk(gclk));
	jdff dff_A_dDXVwRUp2_0(.dout(w_dff_A_XUJijzqz7_0),.din(w_dff_A_dDXVwRUp2_0),.clk(gclk));
	jdff dff_A_XUJijzqz7_0(.dout(w_dff_A_u5TTwT6p4_0),.din(w_dff_A_XUJijzqz7_0),.clk(gclk));
	jdff dff_A_u5TTwT6p4_0(.dout(G12),.din(w_dff_A_u5TTwT6p4_0),.clk(gclk));
	jdff dff_A_FSygimdF5_2(.dout(w_dff_A_QDNmg8Tt6_0),.din(w_dff_A_FSygimdF5_2),.clk(gclk));
	jdff dff_A_QDNmg8Tt6_0(.dout(w_dff_A_A6W6S7Mx7_0),.din(w_dff_A_QDNmg8Tt6_0),.clk(gclk));
	jdff dff_A_A6W6S7Mx7_0(.dout(w_dff_A_PMweFv0y1_0),.din(w_dff_A_A6W6S7Mx7_0),.clk(gclk));
	jdff dff_A_PMweFv0y1_0(.dout(w_dff_A_HhOoxF5I6_0),.din(w_dff_A_PMweFv0y1_0),.clk(gclk));
	jdff dff_A_HhOoxF5I6_0(.dout(w_dff_A_Spf1me6F2_0),.din(w_dff_A_HhOoxF5I6_0),.clk(gclk));
	jdff dff_A_Spf1me6F2_0(.dout(w_dff_A_BW4y78P94_0),.din(w_dff_A_Spf1me6F2_0),.clk(gclk));
	jdff dff_A_BW4y78P94_0(.dout(G30),.din(w_dff_A_BW4y78P94_0),.clk(gclk));
	jdff dff_A_RZoms0eR5_2(.dout(w_dff_A_YZJptP9c8_0),.din(w_dff_A_RZoms0eR5_2),.clk(gclk));
	jdff dff_A_YZJptP9c8_0(.dout(w_dff_A_lVVxvWyr1_0),.din(w_dff_A_YZJptP9c8_0),.clk(gclk));
	jdff dff_A_lVVxvWyr1_0(.dout(w_dff_A_7sneRSUN9_0),.din(w_dff_A_lVVxvWyr1_0),.clk(gclk));
	jdff dff_A_7sneRSUN9_0(.dout(w_dff_A_vVhtA5lP9_0),.din(w_dff_A_7sneRSUN9_0),.clk(gclk));
	jdff dff_A_vVhtA5lP9_0(.dout(w_dff_A_T9bLOFgY9_0),.din(w_dff_A_vVhtA5lP9_0),.clk(gclk));
	jdff dff_A_T9bLOFgY9_0(.dout(w_dff_A_CcrjtClQ3_0),.din(w_dff_A_T9bLOFgY9_0),.clk(gclk));
	jdff dff_A_CcrjtClQ3_0(.dout(G45),.din(w_dff_A_CcrjtClQ3_0),.clk(gclk));
	jdff dff_A_NQySwvJu6_2(.dout(w_dff_A_p55143YZ7_0),.din(w_dff_A_NQySwvJu6_2),.clk(gclk));
	jdff dff_A_p55143YZ7_0(.dout(w_dff_A_IDYeaL2B4_0),.din(w_dff_A_p55143YZ7_0),.clk(gclk));
	jdff dff_A_IDYeaL2B4_0(.dout(w_dff_A_7dEOFYhG3_0),.din(w_dff_A_IDYeaL2B4_0),.clk(gclk));
	jdff dff_A_7dEOFYhG3_0(.dout(w_dff_A_H9lozehi6_0),.din(w_dff_A_7dEOFYhG3_0),.clk(gclk));
	jdff dff_A_H9lozehi6_0(.dout(w_dff_A_mQYWtEAA9_0),.din(w_dff_A_H9lozehi6_0),.clk(gclk));
	jdff dff_A_mQYWtEAA9_0(.dout(w_dff_A_bcjyiXsn8_0),.din(w_dff_A_mQYWtEAA9_0),.clk(gclk));
	jdff dff_A_bcjyiXsn8_0(.dout(G48),.din(w_dff_A_bcjyiXsn8_0),.clk(gclk));
	jdff dff_A_TQOLLgwC9_2(.dout(w_dff_A_pmEkwUVb2_0),.din(w_dff_A_TQOLLgwC9_2),.clk(gclk));
	jdff dff_A_pmEkwUVb2_0(.dout(w_dff_A_9aFBBIwN7_0),.din(w_dff_A_pmEkwUVb2_0),.clk(gclk));
	jdff dff_A_9aFBBIwN7_0(.dout(w_dff_A_POutuJXy3_0),.din(w_dff_A_9aFBBIwN7_0),.clk(gclk));
	jdff dff_A_POutuJXy3_0(.dout(w_dff_A_M7NiAXy27_0),.din(w_dff_A_POutuJXy3_0),.clk(gclk));
	jdff dff_A_M7NiAXy27_0(.dout(w_dff_A_9FGCjAMl1_0),.din(w_dff_A_M7NiAXy27_0),.clk(gclk));
	jdff dff_A_9FGCjAMl1_0(.dout(w_dff_A_3iU71VsT9_0),.din(w_dff_A_9FGCjAMl1_0),.clk(gclk));
	jdff dff_A_3iU71VsT9_0(.dout(G15),.din(w_dff_A_3iU71VsT9_0),.clk(gclk));
	jdff dff_A_5Ycg22Kv1_2(.dout(w_dff_A_qIqGPx9B2_0),.din(w_dff_A_5Ycg22Kv1_2),.clk(gclk));
	jdff dff_A_qIqGPx9B2_0(.dout(w_dff_A_AXvst8434_0),.din(w_dff_A_qIqGPx9B2_0),.clk(gclk));
	jdff dff_A_AXvst8434_0(.dout(w_dff_A_ZGdw4PWF5_0),.din(w_dff_A_AXvst8434_0),.clk(gclk));
	jdff dff_A_ZGdw4PWF5_0(.dout(w_dff_A_YI3b27bo9_0),.din(w_dff_A_ZGdw4PWF5_0),.clk(gclk));
	jdff dff_A_YI3b27bo9_0(.dout(w_dff_A_vcZyp59v1_0),.din(w_dff_A_YI3b27bo9_0),.clk(gclk));
	jdff dff_A_vcZyp59v1_0(.dout(w_dff_A_mwCnbsbj3_0),.din(w_dff_A_vcZyp59v1_0),.clk(gclk));
	jdff dff_A_mwCnbsbj3_0(.dout(G18),.din(w_dff_A_mwCnbsbj3_0),.clk(gclk));
	jdff dff_A_lzIT8M3g4_2(.dout(w_dff_A_rfh8kOMA4_0),.din(w_dff_A_lzIT8M3g4_2),.clk(gclk));
	jdff dff_A_rfh8kOMA4_0(.dout(w_dff_A_CYnUaVIB6_0),.din(w_dff_A_rfh8kOMA4_0),.clk(gclk));
	jdff dff_A_CYnUaVIB6_0(.dout(w_dff_A_7Pa96jhw6_0),.din(w_dff_A_CYnUaVIB6_0),.clk(gclk));
	jdff dff_A_7Pa96jhw6_0(.dout(w_dff_A_sEGMMIQM9_0),.din(w_dff_A_7Pa96jhw6_0),.clk(gclk));
	jdff dff_A_sEGMMIQM9_0(.dout(w_dff_A_VHQRqxOg6_0),.din(w_dff_A_sEGMMIQM9_0),.clk(gclk));
	jdff dff_A_VHQRqxOg6_0(.dout(w_dff_A_Sj71KOIq9_0),.din(w_dff_A_VHQRqxOg6_0),.clk(gclk));
	jdff dff_A_Sj71KOIq9_0(.dout(G21),.din(w_dff_A_Sj71KOIq9_0),.clk(gclk));
	jdff dff_A_uvUXLcwz5_2(.dout(w_dff_A_iRljTdW81_0),.din(w_dff_A_uvUXLcwz5_2),.clk(gclk));
	jdff dff_A_iRljTdW81_0(.dout(w_dff_A_JxUgbM0U2_0),.din(w_dff_A_iRljTdW81_0),.clk(gclk));
	jdff dff_A_JxUgbM0U2_0(.dout(w_dff_A_Z5XN34oW7_0),.din(w_dff_A_JxUgbM0U2_0),.clk(gclk));
	jdff dff_A_Z5XN34oW7_0(.dout(w_dff_A_io1Mu50u3_0),.din(w_dff_A_Z5XN34oW7_0),.clk(gclk));
	jdff dff_A_io1Mu50u3_0(.dout(w_dff_A_4YK3SS4q2_0),.din(w_dff_A_io1Mu50u3_0),.clk(gclk));
	jdff dff_A_4YK3SS4q2_0(.dout(w_dff_A_LLu33uYp7_0),.din(w_dff_A_4YK3SS4q2_0),.clk(gclk));
	jdff dff_A_LLu33uYp7_0(.dout(G24),.din(w_dff_A_LLu33uYp7_0),.clk(gclk));
	jdff dff_A_P2cnVXRN3_2(.dout(w_dff_A_XxmygrCQ4_0),.din(w_dff_A_P2cnVXRN3_2),.clk(gclk));
	jdff dff_A_XxmygrCQ4_0(.dout(w_dff_A_q5q0f57m1_0),.din(w_dff_A_XxmygrCQ4_0),.clk(gclk));
	jdff dff_A_q5q0f57m1_0(.dout(w_dff_A_nbWLKJ4h0_0),.din(w_dff_A_q5q0f57m1_0),.clk(gclk));
	jdff dff_A_nbWLKJ4h0_0(.dout(w_dff_A_hbjlsx3U7_0),.din(w_dff_A_nbWLKJ4h0_0),.clk(gclk));
	jdff dff_A_hbjlsx3U7_0(.dout(w_dff_A_BmdcwmAi6_0),.din(w_dff_A_hbjlsx3U7_0),.clk(gclk));
	jdff dff_A_BmdcwmAi6_0(.dout(w_dff_A_9UcKii0l6_0),.din(w_dff_A_BmdcwmAi6_0),.clk(gclk));
	jdff dff_A_9UcKii0l6_0(.dout(G27),.din(w_dff_A_9UcKii0l6_0),.clk(gclk));
	jdff dff_A_AZ2yvGcJ3_2(.dout(w_dff_A_vAuxRXTY8_0),.din(w_dff_A_AZ2yvGcJ3_2),.clk(gclk));
	jdff dff_A_vAuxRXTY8_0(.dout(w_dff_A_FBZA62DK0_0),.din(w_dff_A_vAuxRXTY8_0),.clk(gclk));
	jdff dff_A_FBZA62DK0_0(.dout(w_dff_A_5VW6dXCi3_0),.din(w_dff_A_FBZA62DK0_0),.clk(gclk));
	jdff dff_A_5VW6dXCi3_0(.dout(w_dff_A_lMWWcJgq9_0),.din(w_dff_A_5VW6dXCi3_0),.clk(gclk));
	jdff dff_A_lMWWcJgq9_0(.dout(w_dff_A_KBalGWIV8_0),.din(w_dff_A_lMWWcJgq9_0),.clk(gclk));
	jdff dff_A_KBalGWIV8_0(.dout(w_dff_A_RuziirYU4_0),.din(w_dff_A_KBalGWIV8_0),.clk(gclk));
	jdff dff_A_RuziirYU4_0(.dout(G33),.din(w_dff_A_RuziirYU4_0),.clk(gclk));
	jdff dff_A_h1KbCkLi7_2(.dout(w_dff_A_csfwnwYU8_0),.din(w_dff_A_h1KbCkLi7_2),.clk(gclk));
	jdff dff_A_csfwnwYU8_0(.dout(w_dff_A_IAoeHS3R0_0),.din(w_dff_A_csfwnwYU8_0),.clk(gclk));
	jdff dff_A_IAoeHS3R0_0(.dout(w_dff_A_dyyzbw0S6_0),.din(w_dff_A_IAoeHS3R0_0),.clk(gclk));
	jdff dff_A_dyyzbw0S6_0(.dout(w_dff_A_4lSJi6Dc8_0),.din(w_dff_A_dyyzbw0S6_0),.clk(gclk));
	jdff dff_A_4lSJi6Dc8_0(.dout(w_dff_A_nKg3xQLb8_0),.din(w_dff_A_4lSJi6Dc8_0),.clk(gclk));
	jdff dff_A_nKg3xQLb8_0(.dout(w_dff_A_6Jvh7HyU0_0),.din(w_dff_A_nKg3xQLb8_0),.clk(gclk));
	jdff dff_A_6Jvh7HyU0_0(.dout(G36),.din(w_dff_A_6Jvh7HyU0_0),.clk(gclk));
	jdff dff_A_FiQj09nF1_2(.dout(w_dff_A_jdMXLw3G7_0),.din(w_dff_A_FiQj09nF1_2),.clk(gclk));
	jdff dff_A_jdMXLw3G7_0(.dout(w_dff_A_ig4vAVge4_0),.din(w_dff_A_jdMXLw3G7_0),.clk(gclk));
	jdff dff_A_ig4vAVge4_0(.dout(w_dff_A_yJtbTHFj1_0),.din(w_dff_A_ig4vAVge4_0),.clk(gclk));
	jdff dff_A_yJtbTHFj1_0(.dout(w_dff_A_1zMHCGuL5_0),.din(w_dff_A_yJtbTHFj1_0),.clk(gclk));
	jdff dff_A_1zMHCGuL5_0(.dout(w_dff_A_bORZuoLS6_0),.din(w_dff_A_1zMHCGuL5_0),.clk(gclk));
	jdff dff_A_bORZuoLS6_0(.dout(w_dff_A_6BPlr4yS6_0),.din(w_dff_A_bORZuoLS6_0),.clk(gclk));
	jdff dff_A_6BPlr4yS6_0(.dout(G39),.din(w_dff_A_6BPlr4yS6_0),.clk(gclk));
	jdff dff_A_WA84vgUW7_2(.dout(w_dff_A_jPhWAmZk1_0),.din(w_dff_A_WA84vgUW7_2),.clk(gclk));
	jdff dff_A_jPhWAmZk1_0(.dout(w_dff_A_XPGCH2QZ1_0),.din(w_dff_A_jPhWAmZk1_0),.clk(gclk));
	jdff dff_A_XPGCH2QZ1_0(.dout(w_dff_A_pGX9e0om2_0),.din(w_dff_A_XPGCH2QZ1_0),.clk(gclk));
	jdff dff_A_pGX9e0om2_0(.dout(w_dff_A_Wti0b0ev4_0),.din(w_dff_A_pGX9e0om2_0),.clk(gclk));
	jdff dff_A_Wti0b0ev4_0(.dout(w_dff_A_UMJhHJEx7_0),.din(w_dff_A_Wti0b0ev4_0),.clk(gclk));
	jdff dff_A_UMJhHJEx7_0(.dout(w_dff_A_YNLFgSwq3_0),.din(w_dff_A_UMJhHJEx7_0),.clk(gclk));
	jdff dff_A_YNLFgSwq3_0(.dout(G42),.din(w_dff_A_YNLFgSwq3_0),.clk(gclk));
	jdff dff_A_sQC4fYt42_2(.dout(G75),.din(w_dff_A_sQC4fYt42_2),.clk(gclk));
	jdff dff_A_V1e0H1oc8_2(.dout(G69),.din(w_dff_A_V1e0H1oc8_2),.clk(gclk));
	jdff dff_A_uG0hByNW5_2(.dout(w_dff_A_2ICqsIVK0_0),.din(w_dff_A_uG0hByNW5_2),.clk(gclk));
	jdff dff_A_2ICqsIVK0_0(.dout(G72),.din(w_dff_A_2ICqsIVK0_0),.clk(gclk));
endmodule

