/*

c880:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 1127
	jand: 153
	jor: 119

Summary:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 1127
	jand: 153
	jor: 119
*/

module c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n101;
	wire n102;
	wire n103;
	wire n105;
	wire n106;
	wire n107;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n118;
	wire n119;
	wire n121;
	wire n122;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire[2:0] w_G1gat_0;
	wire[1:0] w_G1gat_1;
	wire[1:0] w_G8gat_0;
	wire[1:0] w_G13gat_0;
	wire[2:0] w_G17gat_0;
	wire[2:0] w_G17gat_1;
	wire[2:0] w_G17gat_2;
	wire[1:0] w_G26gat_0;
	wire[2:0] w_G29gat_0;
	wire[1:0] w_G36gat_0;
	wire[2:0] w_G42gat_0;
	wire[2:0] w_G42gat_1;
	wire[1:0] w_G42gat_2;
	wire[2:0] w_G51gat_0;
	wire[1:0] w_G51gat_1;
	wire[2:0] w_G55gat_0;
	wire[2:0] w_G59gat_0;
	wire[1:0] w_G59gat_1;
	wire[1:0] w_G68gat_0;
	wire[1:0] w_G75gat_0;
	wire[2:0] w_G80gat_0;
	wire[2:0] w_G91gat_0;
	wire[2:0] w_G96gat_0;
	wire[2:0] w_G101gat_0;
	wire[2:0] w_G106gat_0;
	wire[2:0] w_G111gat_0;
	wire[2:0] w_G116gat_0;
	wire[2:0] w_G121gat_0;
	wire[1:0] w_G126gat_0;
	wire[1:0] w_G130gat_0;
	wire[2:0] w_G138gat_0;
	wire[1:0] w_G138gat_1;
	wire[1:0] w_G143gat_0;
	wire[1:0] w_G146gat_0;
	wire[1:0] w_G149gat_0;
	wire[2:0] w_G153gat_0;
	wire[1:0] w_G156gat_0;
	wire[2:0] w_G159gat_0;
	wire[2:0] w_G159gat_1;
	wire[1:0] w_G159gat_2;
	wire[2:0] w_G165gat_0;
	wire[2:0] w_G165gat_1;
	wire[1:0] w_G165gat_2;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[1:0] w_G171gat_2;
	wire[2:0] w_G177gat_0;
	wire[2:0] w_G177gat_1;
	wire[1:0] w_G177gat_2;
	wire[2:0] w_G183gat_0;
	wire[2:0] w_G183gat_1;
	wire[1:0] w_G183gat_2;
	wire[2:0] w_G189gat_0;
	wire[2:0] w_G189gat_1;
	wire[1:0] w_G189gat_2;
	wire[2:0] w_G195gat_0;
	wire[2:0] w_G195gat_1;
	wire[1:0] w_G195gat_2;
	wire[2:0] w_G201gat_0;
	wire[2:0] w_G201gat_1;
	wire[2:0] w_G201gat_2;
	wire[2:0] w_G210gat_0;
	wire[2:0] w_G210gat_1;
	wire[2:0] w_G210gat_2;
	wire[1:0] w_G210gat_3;
	wire[2:0] w_G219gat_0;
	wire[2:0] w_G219gat_1;
	wire[2:0] w_G219gat_2;
	wire[1:0] w_G219gat_3;
	wire[2:0] w_G228gat_0;
	wire[2:0] w_G228gat_1;
	wire[2:0] w_G228gat_2;
	wire[1:0] w_G228gat_3;
	wire[2:0] w_G237gat_0;
	wire[2:0] w_G237gat_1;
	wire[2:0] w_G237gat_2;
	wire[1:0] w_G237gat_3;
	wire[2:0] w_G246gat_0;
	wire[2:0] w_G246gat_1;
	wire[2:0] w_G246gat_2;
	wire[1:0] w_G246gat_3;
	wire[2:0] w_G255gat_0;
	wire[2:0] w_G261gat_0;
	wire[1:0] w_G268gat_0;
	wire[1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire[2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire[1:0] w_n86_0;
	wire[1:0] w_n88_0;
	wire[2:0] w_n92_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n96_0;
	wire[1:0] w_n98_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n101_0;
	wire[1:0] w_n102_0;
	wire[1:0] w_n106_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n111_0;
	wire[2:0] w_n118_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n143_0;
	wire[1:0] w_n149_0;
	wire[2:0] w_n153_0;
	wire[2:0] w_n153_1;
	wire[2:0] w_n153_2;
	wire[1:0] w_n153_3;
	wire[1:0] w_n154_0;
	wire[1:0] w_n157_0;
	wire[2:0] w_n159_0;
	wire[1:0] w_n159_1;
	wire[1:0] w_n162_0;
	wire[1:0] w_n163_0;
	wire[2:0] w_n165_0;
	wire[2:0] w_n165_1;
	wire[2:0] w_n167_0;
	wire[1:0] w_n167_1;
	wire[2:0] w_n168_0;
	wire[2:0] w_n181_0;
	wire[2:0] w_n181_1;
	wire[2:0] w_n181_2;
	wire[1:0] w_n181_3;
	wire[2:0] w_n193_0;
	wire[1:0] w_n193_1;
	wire[2:0] w_n194_0;
	wire[1:0] w_n196_0;
	wire[1:0] w_n213_0;
	wire[2:0] w_n217_0;
	wire[1:0] w_n217_1;
	wire[1:0] w_n218_0;
	wire[2:0] w_n222_0;
	wire[1:0] w_n222_1;
	wire[1:0] w_n223_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n228_0;
	wire[1:0] w_n230_0;
	wire[1:0] w_n232_0;
	wire[2:0] w_n236_0;
	wire[1:0] w_n238_0;
	wire[2:0] w_n252_0;
	wire[1:0] w_n255_0;
	wire[2:0] w_n273_0;
	wire[2:0] w_n292_0;
	wire[1:0] w_n292_1;
	wire[2:0] w_n296_0;
	wire[1:0] w_n296_1;
	wire[2:0] w_n299_0;
	wire[1:0] w_n299_1;
	wire[1:0] w_n302_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n305_0;
	wire[1:0] w_n305_1;
	wire[2:0] w_n312_0;
	wire[1:0] w_n312_1;
	wire[1:0] w_n315_0;
	wire[2:0] w_n321_0;
	wire[1:0] w_n321_1;
	wire[1:0] w_n322_0;
	wire[2:0] w_n328_0;
	wire[1:0] w_n328_1;
	wire[2:0] w_n329_0;
	wire[2:0] w_n330_0;
	wire[1:0] w_n331_0;
	wire[2:0] w_n335_0;
	wire[2:0] w_n337_0;
	wire[1:0] w_n339_0;
	wire[1:0] w_n340_0;
	wire[2:0] w_n346_0;
	wire[1:0] w_n346_1;
	wire[2:0] w_n347_0;
	wire[2:0] w_n367_0;
	wire[2:0] w_n383_0;
	wire[2:0] w_n405_0;
	wire w_dff_B_CyKwyphr1_2;
	wire w_dff_B_iugJthxE1_1;
	wire w_dff_B_tDtNnlHu9_1;
	wire w_dff_A_jjSD3FkA1_1;
	wire w_dff_B_2w2NwKet5_0;
	wire w_dff_B_GdgUF8cQ0_1;
	wire w_dff_B_WLWUl7eF7_1;
	wire w_dff_B_xwH9UetB0_0;
	wire w_dff_B_bU6U96DH3_1;
	wire w_dff_B_ESnsRQaR5_0;
	wire w_dff_B_8vDVZbqX9_0;
	wire w_dff_B_4fXyhJE60_1;
	wire w_dff_B_PNiG9O2k8_0;
	wire w_dff_B_cH2q8aK22_2;
	wire w_dff_B_6PGRgfmA5_0;
	wire w_dff_B_Rj7S9AwS4_0;
	wire w_dff_B_5PkVdPCL5_0;
	wire w_dff_B_mzqr1oNS7_0;
	wire w_dff_B_GA4BDbyK5_0;
	wire w_dff_B_UNalbLpO1_0;
	wire w_dff_B_auSpZ2Q82_0;
	wire w_dff_B_G2xuKXNM6_0;
	wire w_dff_B_ircdiJlw5_0;
	wire w_dff_B_DdFX4hTk6_0;
	wire w_dff_B_XUZUtypu5_0;
	wire w_dff_B_hORW2yly9_0;
	wire w_dff_B_LAkMJVPZ7_0;
	wire w_dff_A_DJcKU5pm5_1;
	wire w_dff_A_76OVWLZU0_1;
	wire w_dff_A_drbIm2M96_1;
	wire w_dff_A_Va0bTc9T9_1;
	wire w_dff_A_dM5i8yYs9_1;
	wire w_dff_A_Fqq71yoJ7_1;
	wire w_dff_A_gMwGrmXA5_1;
	wire w_dff_A_8LuQ0HYn9_1;
	wire w_dff_B_n3B4a7lS8_0;
	wire w_dff_B_1LaZuo0X7_0;
	wire w_dff_B_vEOIMitj1_0;
	wire w_dff_B_RFRaNVNs6_0;
	wire w_dff_B_tMPfvelr4_0;
	wire w_dff_B_O3NwFjze2_0;
	wire w_dff_B_nkSNQtUL6_0;
	wire w_dff_B_ZTIf6Wlo2_0;
	wire w_dff_B_2a9wlo0A4_0;
	wire w_dff_B_RPP6nf8I6_0;
	wire w_dff_B_v7bZx6Pu4_0;
	wire w_dff_B_FPQEmp059_0;
	wire w_dff_B_LJog64C59_0;
	wire w_dff_B_AqlrS1L85_0;
	wire w_dff_B_0Q2cIPyv4_0;
	wire w_dff_B_IthI9RXJ2_0;
	wire w_dff_B_4CEbYnw38_0;
	wire w_dff_B_jzXK16sE8_0;
	wire w_dff_A_Ucd6nBB01_0;
	wire w_dff_A_iyftkq4J4_0;
	wire w_dff_A_r3WWknnc7_0;
	wire w_dff_A_hYga5udw7_0;
	wire w_dff_B_YE4IuKer1_1;
	wire w_dff_B_vwZ6j0gl8_1;
	wire w_dff_B_ezsaci3V1_1;
	wire w_dff_B_FmOh0vb39_1;
	wire w_dff_A_Ku7EBwKj6_1;
	wire w_dff_A_74RdxEXT9_1;
	wire w_dff_A_ju7K1gXA5_1;
	wire w_dff_A_9WwPqc2N7_1;
	wire w_dff_A_GOqi5TUC6_0;
	wire w_dff_A_LT5vWtVn3_0;
	wire w_dff_A_U74bqfG07_0;
	wire w_dff_A_yFkepAiF0_0;
	wire w_dff_A_i3TYDPGR4_0;
	wire w_dff_A_64gn8B5s4_0;
	wire w_dff_A_JVbeLkoD2_0;
	wire w_dff_A_XUvNKZBq2_0;
	wire w_dff_B_gXBZupkW3_0;
	wire w_dff_B_hKoZQoUf9_0;
	wire w_dff_B_Z32LhIcC5_0;
	wire w_dff_B_N27f2amn7_0;
	wire w_dff_B_sot1kt8j9_0;
	wire w_dff_B_gRK9DI3U2_0;
	wire w_dff_B_DIj5wJvP7_0;
	wire w_dff_B_xrA1lCIC7_0;
	wire w_dff_B_sj7NpmzF7_0;
	wire w_dff_B_usRYsrWj5_0;
	wire w_dff_B_gQ6iSmGV4_0;
	wire w_dff_B_qJEnLQRc6_0;
	wire w_dff_B_O6om52v94_0;
	wire w_dff_B_kSfSpbUW3_0;
	wire w_dff_B_wNHw4sdd2_0;
	wire w_dff_B_NXeFrPuv1_0;
	wire w_dff_B_wyNBG4UK4_0;
	wire w_dff_B_pvGs5Tpn8_1;
	wire w_dff_B_0Sr4TRom6_1;
	wire w_dff_B_I9xaJ2Vs3_1;
	wire w_dff_B_7RiwbCrg6_1;
	wire w_dff_A_MBRSfp1H7_1;
	wire w_dff_A_ZNgEiuxT4_1;
	wire w_dff_A_c2K6wtFV0_1;
	wire w_dff_A_wDsjkRMa9_1;
	wire w_dff_B_ilJVTnfp2_0;
	wire w_dff_B_hqe7xUh36_0;
	wire w_dff_B_taZEckL56_0;
	wire w_dff_B_rwO8bQQN1_0;
	wire w_dff_B_jlcST0ad6_0;
	wire w_dff_B_nmyHmH251_0;
	wire w_dff_B_bF6rdf6s2_0;
	wire w_dff_B_Y6OtWTIO5_0;
	wire w_dff_B_EkS5AOkG9_0;
	wire w_dff_B_7KNDYjcd5_0;
	wire w_dff_B_f27Rd26J6_0;
	wire w_dff_B_RSLK5cRb2_0;
	wire w_dff_B_WTCjI5Ai7_0;
	wire w_dff_B_G9BcWP8M4_0;
	wire w_dff_B_VSJf4baY0_0;
	wire w_dff_B_Njkvh2yk1_0;
	wire w_dff_B_5J4qcP2F2_0;
	wire w_dff_A_AneMG0E56_1;
	wire w_dff_A_gIRiRx1j2_1;
	wire w_dff_B_c6VKpkoU6_1;
	wire w_dff_B_vFuiJCzA9_1;
	wire w_dff_B_wI1HhxIi1_1;
	wire w_dff_B_r5HwmhLs8_1;
	wire w_dff_B_pLQsUUeC0_1;
	wire w_dff_B_OtGd4gEO3_1;
	wire w_dff_B_uXvqC6gh2_1;
	wire w_dff_B_joR9MMqD7_1;
	wire w_dff_B_Aa0b0IwG6_1;
	wire w_dff_B_S5Soqeu77_1;
	wire w_dff_B_WAM8w3rF1_1;
	wire w_dff_B_cx6ixeKO8_1;
	wire w_dff_B_EapkadzS9_1;
	wire w_dff_B_7Bv86fkV0_1;
	wire w_dff_B_vQVTNHeQ5_1;
	wire w_dff_B_LvU4dEk43_1;
	wire w_dff_B_SftK35936_1;
	wire w_dff_B_BJUthwO50_1;
	wire w_dff_B_TPc0ucj43_1;
	wire w_dff_A_h16rlwVR8_0;
	wire w_dff_A_XXvf1WCp3_0;
	wire w_dff_A_qolJqMAb1_0;
	wire w_dff_A_WWX9KilH4_0;
	wire w_dff_A_bnoQoq9v7_0;
	wire w_dff_A_5gsQMc7H6_0;
	wire w_dff_A_Zph5uTU19_0;
	wire w_dff_B_IXoUkkfG5_0;
	wire w_dff_B_QdShgpTW3_0;
	wire w_dff_B_TpwtzfxI7_0;
	wire w_dff_B_T0q9xtsL5_0;
	wire w_dff_B_oCAS8xxo5_0;
	wire w_dff_B_PG58jnzw4_0;
	wire w_dff_B_Ys9LyCPv1_0;
	wire w_dff_B_YdjaX97Q5_0;
	wire w_dff_B_aR1sYrKA9_0;
	wire w_dff_B_mT3mTevV1_0;
	wire w_dff_B_aaZdzcYZ6_0;
	wire w_dff_B_dVkW5Q0U2_0;
	wire w_dff_B_BrptghCx9_0;
	wire w_dff_B_bDjocvHb4_0;
	wire w_dff_B_swn9wA5a8_0;
	wire w_dff_B_8luZ1cp45_0;
	wire w_dff_B_Ie2yRgld1_0;
	wire w_dff_B_RTMFee0S6_0;
	wire w_dff_B_nusyD60S3_0;
	wire w_dff_A_8BBT3WcH8_1;
	wire w_dff_A_LGmn9IrG1_2;
	wire w_dff_A_eb2a4rMR8_0;
	wire w_dff_A_CgLMGN279_0;
	wire w_dff_A_hesCPpLD5_0;
	wire w_dff_A_B2yRUTx84_0;
	wire w_dff_A_UVL9DDTW0_2;
	wire w_dff_A_ix8qC5Da8_2;
	wire w_dff_B_v9e0R0VX8_0;
	wire w_dff_B_sSEyuvey6_0;
	wire w_dff_B_qZaEHHNq0_0;
	wire w_dff_B_XZetI1kQ9_0;
	wire w_dff_B_vlfLJufO0_0;
	wire w_dff_B_3Di8qKXO4_0;
	wire w_dff_B_fbJ5YCMu6_0;
	wire w_dff_A_lWudaLyD8_1;
	wire w_dff_A_3sWm1OLd7_1;
	wire w_dff_A_LuSFRLYE3_1;
	wire w_dff_A_8RUE70Lh5_1;
	wire w_dff_A_zs2itGKQ5_1;
	wire w_dff_A_BgCQorEw5_1;
	wire w_dff_A_Bw1e8Sbi0_1;
	wire w_dff_B_KRRdZg4H6_0;
	wire w_dff_B_l9GxMlbw1_0;
	wire w_dff_B_MIs4jiPP3_0;
	wire w_dff_B_Wtgiavdv5_0;
	wire w_dff_B_z0l5yEZX2_0;
	wire w_dff_B_ImFGVWlM8_0;
	wire w_dff_B_3Bbl0ugy4_0;
	wire w_dff_B_RHfbd8kW2_0;
	wire w_dff_B_pD1CfkvY9_0;
	wire w_dff_B_zEyI8zSt7_0;
	wire w_dff_B_P0wL9Awp2_0;
	wire w_dff_B_3nBWanky2_0;
	wire w_dff_B_nq3fvDGS9_0;
	wire w_dff_B_fHAgzPVK0_0;
	wire w_dff_B_sAGoI8hL6_0;
	wire w_dff_B_7a9JN6SX4_0;
	wire w_dff_B_XGKfbu7B3_0;
	wire w_dff_B_kobm6ENd0_0;
	wire w_dff_B_pZXeD6dm7_0;
	wire w_dff_B_hosz5vSi9_0;
	wire w_dff_B_FNrHhMWb6_0;
	wire w_dff_B_p4N9zMSy3_0;
	wire w_dff_B_pi2wFGve7_0;
	wire w_dff_B_IlWIID078_0;
	wire w_dff_B_DQGuZUL71_0;
	wire w_dff_B_4oR1tRUd7_0;
	wire w_dff_B_LBG5OWJQ7_0;
	wire w_dff_B_WdIU6xvz1_0;
	wire w_dff_B_OcyUjgvv4_0;
	wire w_dff_B_NgN9tBnN1_0;
	wire w_dff_A_V6zhMGb76_1;
	wire w_dff_A_K4s2Dg1J8_1;
	wire w_dff_A_WN9MZPBm3_1;
	wire w_dff_A_J06Ca8h29_1;
	wire w_dff_A_prDYwrzb7_1;
	wire w_dff_A_jPujGZjQ0_1;
	wire w_dff_A_BDMPWaHy9_1;
	wire w_dff_A_hj6QrRjR0_1;
	wire w_dff_A_I9eTOsSs8_1;
	wire w_dff_B_6G9LXMK19_1;
	wire w_dff_B_1RVjmJHb9_1;
	wire w_dff_B_oKw6tXG59_1;
	wire w_dff_A_CUi5cSKk9_1;
	wire w_dff_A_Uld0OURf3_1;
	wire w_dff_A_2EdkuGeC3_1;
	wire w_dff_A_hXGbQzsN6_1;
	wire w_dff_A_5wYUwuVt7_1;
	wire w_dff_A_ZUa6FsL69_1;
	wire w_dff_A_9OHafTkt0_1;
	wire w_dff_A_201kpSRp5_2;
	wire w_dff_A_259hgUSJ5_2;
	wire w_dff_A_CCTWhhIh1_2;
	wire w_dff_A_hBuj7yyj4_2;
	wire w_dff_A_ZNSlLW4L0_2;
	wire w_dff_A_kMFyP6AF2_2;
	wire w_dff_A_vqEMsjDs5_2;
	wire w_dff_A_CFrdlXM94_2;
	wire w_dff_A_5lW1YvpY6_2;
	wire w_dff_A_9SqySWtc3_2;
	wire w_dff_A_lL6cgLL13_2;
	wire w_dff_B_XR8PMdAH1_0;
	wire w_dff_B_a33JBwVM7_0;
	wire w_dff_B_k4kf8T8c1_0;
	wire w_dff_B_Oj41tBd14_0;
	wire w_dff_A_1bvlYosF7_1;
	wire w_dff_A_7TCj7ijA7_1;
	wire w_dff_A_RrDniVTh0_1;
	wire w_dff_A_16O2qm1c0_1;
	wire w_dff_B_C4Dvv0t19_1;
	wire w_dff_B_sgQOOH0F8_1;
	wire w_dff_B_jLQujL9a6_1;
	wire w_dff_B_ukEnEh6a8_0;
	wire w_dff_B_f95Zyvt28_0;
	wire w_dff_B_maOir8CZ6_0;
	wire w_dff_B_XoYr91NN9_0;
	wire w_dff_A_i04SvP2Y7_1;
	wire w_dff_A_8dkBumGM4_1;
	wire w_dff_A_Dhx21nBw0_1;
	wire w_dff_A_wH5Gg4sN4_1;
	wire w_dff_B_GPgp6nAp4_1;
	wire w_dff_B_iJn8jKKa6_1;
	wire w_dff_B_20IZbmUG6_1;
	wire w_dff_B_HkS9qsD45_1;
	wire w_dff_B_BUPKsVHh9_1;
	wire w_dff_B_kRLr6eC78_1;
	wire w_dff_B_ZsmjwWGx2_1;
	wire w_dff_B_VgUtxseO0_0;
	wire w_dff_B_NHLTXGZ07_0;
	wire w_dff_B_COiCVePz9_0;
	wire w_dff_B_0fUM2BM80_0;
	wire w_dff_B_DXuKsD0O9_0;
	wire w_dff_B_7AdnsBA27_0;
	wire w_dff_B_KvpcJOkT2_0;
	wire w_dff_B_zCYoDjUN4_0;
	wire w_dff_B_aHLx74Sb4_0;
	wire w_dff_B_ObHH3cAX7_0;
	wire w_dff_B_dKybQjpE7_0;
	wire w_dff_B_0DzC5rDp0_0;
	wire w_dff_B_2t9vMCFu3_0;
	wire w_dff_B_gTN7xQnf8_0;
	wire w_dff_B_pwnW2eiY9_0;
	wire w_dff_B_ImGLq4gj7_0;
	wire w_dff_A_1j4UG0cm6_1;
	wire w_dff_A_4OOSH44w8_1;
	wire w_dff_A_IrK88W3t1_1;
	wire w_dff_A_9qqrJkE60_1;
	wire w_dff_A_X1OJdXbj3_1;
	wire w_dff_B_JiGp95Kg4_0;
	wire w_dff_B_TFm4noDO6_0;
	wire w_dff_B_RTezwXI73_0;
	wire w_dff_B_lNHmu34x3_0;
	wire w_dff_B_jvsOuxFA9_0;
	wire w_dff_B_4rke9fUf9_1;
	wire w_dff_B_sV1MvrWv7_1;
	wire w_dff_B_Gkam16Qx8_1;
	wire w_dff_B_rGM53A5o9_1;
	wire w_dff_B_VZdcpzdW2_1;
	wire w_dff_B_eZK03X1m8_1;
	wire w_dff_B_gK09yN0x5_1;
	wire w_dff_B_qvWiE8fs9_1;
	wire w_dff_B_1pd4Ccwh2_1;
	wire w_dff_B_prFWXAF80_1;
	wire w_dff_B_g8rE8TPU0_1;
	wire w_dff_B_mTeFZ3c33_1;
	wire w_dff_B_gPEb4QjS6_1;
	wire w_dff_B_ozykzldL0_1;
	wire w_dff_B_7R9s9ooO7_1;
	wire w_dff_B_zPTo8wku1_0;
	wire w_dff_B_PBYuE5wH7_0;
	wire w_dff_B_N1VuPPoD6_0;
	wire w_dff_B_vRlCJ29I2_0;
	wire w_dff_B_cs0Dx8UG2_0;
	wire w_dff_B_YUvVzvXC8_0;
	wire w_dff_A_s5rCXlAG6_0;
	wire w_dff_A_6mVfejcr1_0;
	wire w_dff_A_KrcYq9679_0;
	wire w_dff_A_AZb9FAO09_0;
	wire w_dff_A_DYCW0Jmy5_0;
	wire w_dff_A_cIMVAcIE0_0;
	wire w_dff_A_YIhTZkIK0_2;
	wire w_dff_A_mNcjiUTS4_0;
	wire w_dff_A_zPYlU2wa5_0;
	wire w_dff_A_8OGcqSg49_0;
	wire w_dff_A_gw4B2maH7_0;
	wire w_dff_A_2UTuchFl9_0;
	wire w_dff_A_NjUnijN24_0;
	wire w_dff_B_FE3FwbSM1_1;
	wire w_dff_A_5nyxg60e1_0;
	wire w_dff_A_IuWTlpDl7_0;
	wire w_dff_A_z1KooGNv4_0;
	wire w_dff_A_u0cpHpTX4_0;
	wire w_dff_A_mZxIiWQ83_0;
	wire w_dff_A_pW4y1Ak80_0;
	wire w_dff_A_k6DoSIxV4_0;
	wire w_dff_A_zVmWF26z1_1;
	wire w_dff_A_BRUnb4Ww5_1;
	wire w_dff_A_d7y0z4AG3_1;
	wire w_dff_A_OBdixHz37_1;
	wire w_dff_A_xZZX1C1g8_1;
	wire w_dff_A_Yi1MI5Qq2_1;
	wire w_dff_A_cZ3dTSwV8_1;
	wire w_dff_A_QKmOS0196_1;
	wire w_dff_A_hma2NagD0_1;
	wire w_dff_B_spsMgE7k2_0;
	wire w_dff_B_HxHEbcII6_0;
	wire w_dff_B_lCxEUWz72_0;
	wire w_dff_A_CVFts5Eh3_1;
	wire w_dff_A_6rQmRFlr7_1;
	wire w_dff_A_bNm6HBDy8_1;
	wire w_dff_A_SNkIjNkL5_1;
	wire w_dff_A_wgtPdGVE7_1;
	wire w_dff_A_00tgw1860_1;
	wire w_dff_A_4yaqyCEp6_1;
	wire w_dff_A_EWSSpqNB4_2;
	wire w_dff_A_mvQ2J5K39_2;
	wire w_dff_A_FgcSLf711_2;
	wire w_dff_A_6uBggni70_2;
	wire w_dff_A_1wDC8Hp87_2;
	wire w_dff_A_sENeX9xq0_2;
	wire w_dff_A_ZrpWIYCz2_2;
	wire w_dff_A_51SqRrIP5_2;
	wire w_dff_A_Fr8kzAYO2_2;
	wire w_dff_A_pkDTK9Bw3_2;
	wire w_dff_A_jWD1m8Ga0_2;
	wire w_dff_B_LewbkPHH6_0;
	wire w_dff_B_3AECi5ED9_0;
	wire w_dff_B_iE6YmXYw3_0;
	wire w_dff_B_oz6HQKjY0_0;
	wire w_dff_B_jVvkZzmh1_0;
	wire w_dff_B_TDcSGP7N1_0;
	wire w_dff_B_WlDYEft91_0;
	wire w_dff_B_XtXhwEY92_0;
	wire w_dff_B_0hzHmD3M5_0;
	wire w_dff_B_Nigc0Z265_0;
	wire w_dff_B_QbUYHx6i4_0;
	wire w_dff_B_7HwCOTBq1_0;
	wire w_dff_B_QN60WPBm1_0;
	wire w_dff_B_ee4C7dX55_0;
	wire w_dff_B_IJFyViog8_0;
	wire w_dff_B_PMLc6udB4_0;
	wire w_dff_A_oKlz0ELJ7_1;
	wire w_dff_A_F6F0Br6R1_1;
	wire w_dff_A_rkVxnocP7_1;
	wire w_dff_A_p2C2SppA4_1;
	wire w_dff_A_vfPBbFAz9_1;
	wire w_dff_B_v1xyCebV4_1;
	wire w_dff_A_OM48yGBA4_0;
	wire w_dff_A_SA7BZnPm1_0;
	wire w_dff_B_wfkIujoZ8_0;
	wire w_dff_B_ckaEptPj1_0;
	wire w_dff_B_eeW5rn2X8_0;
	wire w_dff_B_O67J6Nxd7_0;
	wire w_dff_B_UyJSPswS6_0;
	wire w_dff_B_whdvNOk09_3;
	wire w_dff_A_Nhdao0Dr4_2;
	wire w_dff_B_jOd7JQF56_3;
	wire w_dff_B_daADxTze6_3;
	wire w_dff_B_FqcmaZdc7_3;
	wire w_dff_B_FZZmvEat2_3;
	wire w_dff_B_nvMgiuIL2_3;
	wire w_dff_B_YuRNS4hx1_3;
	wire w_dff_B_J8ljZcny0_3;
	wire w_dff_B_T91JKijC2_3;
	wire w_dff_A_rVAjY0GK0_0;
	wire w_dff_A_3Oqe3ufH6_0;
	wire w_dff_A_b5e1wHnW1_0;
	wire w_dff_A_yx6M2I7s5_0;
	wire w_dff_A_eVvwObL41_0;
	wire w_dff_A_RYFJvG568_0;
	wire w_dff_A_5dfcbgM47_0;
	wire w_dff_A_t7KS4ed80_0;
	wire w_dff_A_18ZhxSlV5_1;
	wire w_dff_A_lIgj2OvW9_1;
	wire w_dff_B_O9oLpDuU0_3;
	wire w_dff_B_R02UGAWA1_3;
	wire w_dff_B_1MraEhNs2_3;
	wire w_dff_B_x57ofOHd6_3;
	wire w_dff_B_Zgzw6iPU8_3;
	wire w_dff_B_t2zJa4iU9_3;
	wire w_dff_B_UfnRBDC88_3;
	wire w_dff_B_wlsGuj6l3_3;
	wire w_dff_B_uGQMOXZ37_3;
	wire w_dff_B_nzN8IDbZ5_3;
	wire w_dff_B_V3pupD2l2_1;
	wire w_dff_B_kkK3U1ve9_1;
	wire w_dff_B_qV8ONmbE7_1;
	wire w_dff_B_ymLB1aEk1_1;
	wire w_dff_B_OhUSpVA47_1;
	wire w_dff_B_Co37Av8c6_1;
	wire w_dff_B_pF0LVP5R3_1;
	wire w_dff_B_N4REVMAn7_1;
	wire w_dff_B_bRPOcEi75_1;
	wire w_dff_B_H1BwVxyk3_1;
	wire w_dff_B_OV6HhMtM7_1;
	wire w_dff_B_zw978dEx9_1;
	wire w_dff_B_ozOiaOpt3_1;
	wire w_dff_B_soCIg1hW9_1;
	wire w_dff_B_JwetYlcX5_1;
	wire w_dff_B_AY2Mtqzl2_1;
	wire w_dff_B_WfuUDdre2_1;
	wire w_dff_B_qQiaIzkt0_0;
	wire w_dff_B_PPO2YRwi6_0;
	wire w_dff_B_dRZnWDra1_0;
	wire w_dff_B_gacHT41n2_0;
	wire w_dff_B_TFk3Smfx4_0;
	wire w_dff_B_LIcxoJsr7_0;
	wire w_dff_B_zhzCgr9l2_0;
	wire w_dff_A_C5PfbyWd0_0;
	wire w_dff_A_6P6xMBd96_0;
	wire w_dff_A_mDgRez6e5_0;
	wire w_dff_A_S9rtRJqS2_0;
	wire w_dff_A_F09O55e07_0;
	wire w_dff_A_vNIgRCAi0_0;
	wire w_dff_A_sEYTIeD96_0;
	wire w_dff_A_E9Adb3CX6_0;
	wire w_dff_A_Ifgm6QmN8_0;
	wire w_dff_A_I1hxqBkG5_0;
	wire w_dff_A_bS7DxMq41_0;
	wire w_dff_A_OFRLRvej8_0;
	wire w_dff_A_nrjRGeno0_0;
	wire w_dff_A_oj9M9gvy2_0;
	wire w_dff_B_1uOhd1uu6_1;
	wire w_dff_B_o8rM7Yca6_1;
	wire w_dff_B_IyqeUokb7_1;
	wire w_dff_B_hvMQNGkC2_1;
	wire w_dff_B_xNk9LDaO0_1;
	wire w_dff_B_zKiMtKk26_1;
	wire w_dff_B_whaycpAI9_1;
	wire w_dff_B_fILuNpqi9_1;
	wire w_dff_B_GIwfvGCa0_1;
	wire w_dff_B_q2cswN5H8_0;
	wire w_dff_A_rPv8zhsi0_0;
	wire w_dff_B_QlEQ6RiZ3_1;
	wire w_dff_A_WOVoZcG36_0;
	wire w_dff_A_84d0TDkI9_0;
	wire w_dff_A_gvbS2i9b2_0;
	wire w_dff_A_4EQMkSy42_1;
	wire w_dff_A_3L7vHM4g2_1;
	wire w_dff_A_bC5DtVfh7_1;
	wire w_dff_A_JsRBExNr4_1;
	wire w_dff_A_OLHkUQAD4_1;
	wire w_dff_A_ImafkSlk0_1;
	wire w_dff_A_MYpj7YG87_1;
	wire w_dff_A_YXUvDKir7_1;
	wire w_dff_A_Ex86Bgfe7_2;
	wire w_dff_A_47uOJb8k8_2;
	wire w_dff_A_VoIcRHx63_2;
	wire w_dff_A_MOS8ERis5_2;
	wire w_dff_A_AeIcqstQ4_2;
	wire w_dff_A_U9wheQsN1_2;
	wire w_dff_A_kBTG5W2H9_2;
	wire w_dff_A_PvdxKnbG1_2;
	wire w_dff_A_jpLbGSZ38_1;
	wire w_dff_A_HkXStBlK6_1;
	wire w_dff_A_ITAYOnLV4_1;
	wire w_dff_A_cKpffvdx4_1;
	wire w_dff_A_uewzBx6T7_1;
	wire w_dff_A_XbUo13MA8_1;
	wire w_dff_A_YtUhTfeo9_1;
	wire w_dff_A_galFhZhB6_1;
	wire w_dff_A_TJPkR2Tu3_2;
	wire w_dff_A_5U9LdHQq1_2;
	wire w_dff_A_ZUSVhw7t6_2;
	wire w_dff_A_vHo74eu67_2;
	wire w_dff_A_hGdyEgPe1_2;
	wire w_dff_A_XJNc4xWq8_2;
	wire w_dff_A_c8oc95er8_2;
	wire w_dff_A_aq6BOP380_2;
	wire w_dff_B_TEqq0CvK2_0;
	wire w_dff_A_ythxWxRF6_0;
	wire w_dff_A_ugzhzE3Q9_0;
	wire w_dff_A_6UN2C2Xw2_0;
	wire w_dff_B_uESYCf1D5_1;
	wire w_dff_A_Mdeczmo63_0;
	wire w_dff_A_wQEL6ZLk0_0;
	wire w_dff_A_E1MrlAA19_0;
	wire w_dff_A_TfGSNyHS9_0;
	wire w_dff_A_FKKbzkpB8_0;
	wire w_dff_A_TxQbYvda3_0;
	wire w_dff_A_gZx3R28Z2_0;
	wire w_dff_A_LxCX8sQ08_0;
	wire w_dff_A_wP8LvX911_0;
	wire w_dff_A_1drCJS6Y4_0;
	wire w_dff_A_h75rBSBt9_0;
	wire w_dff_A_r67ewH9Y4_0;
	wire w_dff_A_p7ylLqnr5_0;
	wire w_dff_A_9GKFZAmg5_2;
	wire w_dff_A_lU0Cntqy3_2;
	wire w_dff_A_DuzjXoJW8_2;
	wire w_dff_A_rdzFG80g1_2;
	wire w_dff_B_aqjt3HhL1_1;
	wire w_dff_A_PkIF8hws6_1;
	wire w_dff_A_L6Dd8G5R1_1;
	wire w_dff_A_ShOk8JTM8_1;
	wire w_dff_A_VNB054K53_1;
	wire w_dff_A_RO9ze0Q51_1;
	wire w_dff_A_9OjhhdMe0_1;
	wire w_dff_B_cuGwXApU3_2;
	wire w_dff_B_o2S9G4eD4_2;
	wire w_dff_B_1cNUGuJs7_2;
	wire w_dff_B_0BQ6LSLO5_2;
	wire w_dff_A_Y5f2zBtt0_0;
	wire w_dff_A_ikf9a0rw9_0;
	wire w_dff_A_gqB3bEwg7_0;
	wire w_dff_A_n27r3JlS9_0;
	wire w_dff_A_N9bhLb198_0;
	wire w_dff_A_pgeauC2i2_0;
	wire w_dff_A_GIMa11pH2_0;
	wire w_dff_A_M4yjlATT5_0;
	wire w_dff_A_coz4d7269_2;
	wire w_dff_A_pBmMvaYD8_2;
	wire w_dff_A_nXnt9UZ37_2;
	wire w_dff_A_XBC0j54E6_2;
	wire w_dff_B_clXIMNx08_1;
	wire w_dff_B_uNIxL1w15_1;
	wire w_dff_B_NEJpFa1Y4_1;
	wire w_dff_B_dHmHW6Ni5_1;
	wire w_dff_B_6g7n988u1_1;
	wire w_dff_B_acWBpf4X8_1;
	wire w_dff_B_3DsWS1yx8_1;
	wire w_dff_B_aQp2wqku5_1;
	wire w_dff_B_kgLBemVM5_1;
	wire w_dff_B_ZEfKWUgn0_1;
	wire w_dff_B_5tU4TEeO2_0;
	wire w_dff_B_7ZCE6cac4_0;
	wire w_dff_B_bmyX14cA2_1;
	wire w_dff_B_yHh7Pf790_1;
	wire w_dff_B_gRf1Ty346_1;
	wire w_dff_B_BN4xaQeZ1_1;
	wire w_dff_B_vr0TsmQz8_1;
	wire w_dff_B_sgSxXV373_1;
	wire w_dff_B_X9XwSFDQ9_1;
	wire w_dff_B_AYIgoPJz7_1;
	wire w_dff_B_WPPIywU42_1;
	wire w_dff_B_FG5AiP5E0_2;
	wire w_dff_B_JfsPZuPH7_2;
	wire w_dff_B_QMQtV8nj2_2;
	wire w_dff_B_snVtZAwb5_2;
	wire w_dff_B_gCXJgSho5_2;
	wire w_dff_B_h0h555jf1_2;
	wire w_dff_B_ffpzhXNI9_2;
	wire w_dff_B_MyAcuUYg3_2;
	wire w_dff_B_Kewu7pk98_2;
	wire w_dff_A_XZbDj4xZ5_0;
	wire w_dff_A_OMy2n1rb9_0;
	wire w_dff_A_VmgtsNXi3_0;
	wire w_dff_A_l5M72jJp2_0;
	wire w_dff_A_pVfSXInm1_0;
	wire w_dff_A_it8krLq24_0;
	wire w_dff_A_OpWZAwtm4_0;
	wire w_dff_A_HHefhRMK2_0;
	wire w_dff_A_VD6wq4HN3_0;
	wire w_dff_A_QNE8kluf0_1;
	wire w_dff_A_xClHQgzr7_1;
	wire w_dff_A_HeqR0W707_1;
	wire w_dff_A_7kdvXk797_1;
	wire w_dff_A_28rE5bO83_1;
	wire w_dff_A_lsXK59Mm0_1;
	wire w_dff_A_dplABmtu7_1;
	wire w_dff_A_wvSjaXfD5_1;
	wire w_dff_A_iiGZ1f197_1;
	wire w_dff_A_P9E7V1247_0;
	wire w_dff_A_rxtSPeVE2_1;
	wire w_dff_A_50LvCA3d3_0;
	wire w_dff_A_RUMYQ1GU7_0;
	wire w_dff_A_SkUdZt1p7_0;
	wire w_dff_A_mL6SUM955_0;
	wire w_dff_A_SU8vcFnq8_0;
	wire w_dff_A_1septHAP6_1;
	wire w_dff_A_dLeIfbgb5_1;
	wire w_dff_A_7WQ57LK56_1;
	wire w_dff_A_ik8YJjHT4_1;
	wire w_dff_A_acYFoEt74_1;
	wire w_dff_A_hHlQe7d67_1;
	wire w_dff_A_LbhkGPRU4_1;
	wire w_dff_A_RkxdeWDZ7_1;
	wire w_dff_A_HcbnxuwG3_2;
	wire w_dff_A_JLQFQzWD1_2;
	wire w_dff_A_NLHx8rSA3_2;
	wire w_dff_A_yuUaDZct5_2;
	wire w_dff_A_ZrXyeeNW3_2;
	wire w_dff_A_nDANibwo2_2;
	wire w_dff_A_pcTaRTIg6_2;
	wire w_dff_A_jR9fRiDK2_2;
	wire w_dff_A_CaeuMWeM4_2;
	wire w_dff_A_K5QYDIK07_2;
	wire w_dff_A_9ga3GXDX0_2;
	wire w_dff_A_WAjYHuCH9_2;
	wire w_dff_A_5RgSses18_1;
	wire w_dff_A_SKGtrvqT2_1;
	wire w_dff_A_uY4irrfR3_1;
	wire w_dff_A_JO6lxcXS8_1;
	wire w_dff_A_RLcVChcq6_1;
	wire w_dff_A_IRRUgXBZ4_1;
	wire w_dff_A_KNWiplwD2_1;
	wire w_dff_A_llG7awQD0_1;
	wire w_dff_A_GyEHmUoP2_1;
	wire w_dff_B_41bkNbQJ2_1;
	wire w_dff_A_wmwB03id7_1;
	wire w_dff_A_S1hGICed4_1;
	wire w_dff_A_e02uxWhd3_1;
	wire w_dff_A_w79Okj218_1;
	wire w_dff_A_DZe664RI1_1;
	wire w_dff_A_yBSFLR1Y2_1;
	wire w_dff_A_JMRI1rol2_1;
	wire w_dff_A_rwupaW538_2;
	wire w_dff_A_ksVZSOd59_2;
	wire w_dff_A_Ar8F1l249_1;
	wire w_dff_A_KLPTewSx0_1;
	wire w_dff_A_pQu9YZul1_2;
	wire w_dff_A_WXfcxGc05_2;
	wire w_dff_B_YXTVlwAl6_0;
	wire w_dff_A_DSxhz7Xv4_0;
	wire w_dff_A_fd6vNQtk6_0;
	wire w_dff_A_i1fXFduF3_0;
	wire w_dff_A_auBPxiDF9_1;
	wire w_dff_B_URNE08AT0_2;
	wire w_dff_B_hCGwS8mQ1_2;
	wire w_dff_B_gxKLwhGZ4_2;
	wire w_dff_B_FlFqBa146_2;
	wire w_dff_A_KpLc9riO5_0;
	wire w_dff_A_ZDoMkGcH7_0;
	wire w_dff_A_2Ofwe7XL4_0;
	wire w_dff_A_FXonsxuv3_0;
	wire w_dff_A_1X3uMO1W8_0;
	wire w_dff_A_ITZ0XuNp3_0;
	wire w_dff_A_914qiOEl3_0;
	wire w_dff_A_jGGLLWCh5_0;
	wire w_dff_A_46jUHdup2_1;
	wire w_dff_A_2Vjpfe6O8_1;
	wire w_dff_A_O4OTqwSL0_1;
	wire w_dff_A_5HyzhKfF7_1;
	wire w_dff_A_4M1fZEW37_2;
	wire w_dff_A_4hyzWsZI6_2;
	wire w_dff_A_Dt3WrPyW9_2;
	wire w_dff_A_fMtRVZPj4_2;
	wire w_dff_A_RJifzXoI1_2;
	wire w_dff_A_oVk6XzCn2_2;
	wire w_dff_A_wNamG5Jj6_2;
	wire w_dff_A_yNv5bI6Q9_2;
	wire w_dff_A_ZqyevI922_0;
	wire w_dff_A_k2fe3CQF4_0;
	wire w_dff_A_36VZNr936_0;
	wire w_dff_A_TldeYhD49_0;
	wire w_dff_A_37W5QOov8_0;
	wire w_dff_A_34NJyDMq2_0;
	wire w_dff_A_dAWNpyVM0_0;
	wire w_dff_A_rvGRHzXk8_0;
	wire w_dff_B_d0rmJPO08_0;
	wire w_dff_B_lj9VG66f1_0;
	wire w_dff_B_6AOg5QhU1_0;
	wire w_dff_A_E5PkoBVc7_0;
	wire w_dff_A_gXaunhRy7_0;
	wire w_dff_A_XNiufU1F4_0;
	wire w_dff_A_x4rl85sv9_0;
	wire w_dff_A_9ClFW5Z38_2;
	wire w_dff_A_Ya1aMsvR2_2;
	wire w_dff_A_h5TVYHoT7_2;
	wire w_dff_A_gwjujEoB2_2;
	wire w_dff_A_GboRYmrx5_2;
	wire w_dff_A_JTiRaHTM1_0;
	wire w_dff_A_gd0sAq6F5_0;
	wire w_dff_A_guMaubLw1_0;
	wire w_dff_A_xzquZ7UM4_0;
	wire w_dff_A_Vk9D0hN00_0;
	wire w_dff_A_qNPOQFP58_1;
	wire w_dff_A_bjnGDSPe2_1;
	wire w_dff_A_wjyKYs0U3_1;
	wire w_dff_A_C4m0W6bJ3_1;
	wire w_dff_A_Q1AbWXoR0_1;
	wire w_dff_A_zOacub3q2_1;
	wire w_dff_A_jGoQ9h4C1_1;
	wire w_dff_A_hNoLYn6H2_2;
	wire w_dff_A_NX7RPgNm3_2;
	wire w_dff_A_7ZSdWsH67_2;
	wire w_dff_A_dTZzk9vt5_2;
	wire w_dff_A_Dar61H9R8_2;
	wire w_dff_A_0vDvbFg78_2;
	wire w_dff_A_h9WWGJRw2_2;
	wire w_dff_A_lwGGzGvu8_2;
	wire w_dff_A_4ZnhGBAl6_2;
	wire w_dff_A_456Kl9v00_2;
	wire w_dff_A_08epPKth5_2;
	wire w_dff_A_vgQnunVY8_1;
	wire w_dff_A_1vBoSNfe5_1;
	wire w_dff_A_CcRdQOYK7_1;
	wire w_dff_A_HiSFdrFZ0_1;
	wire w_dff_A_xqDhygg53_1;
	wire w_dff_A_btL9Agcb8_1;
	wire w_dff_A_XbtpfE8j7_1;
	wire w_dff_A_iH9anqzM4_1;
	wire w_dff_A_HARwFZmJ1_1;
	wire w_dff_B_mZPw0CLR8_0;
	wire w_dff_B_BTqafFDX7_0;
	wire w_dff_B_2NlrS6577_0;
	wire w_dff_B_XdB8JRhX9_0;
	wire w_dff_A_jk2LrdXk9_0;
	wire w_dff_A_K71u5oYo0_2;
	wire w_dff_A_VJz64C2M0_2;
	wire w_dff_A_Ol41ZdeR4_2;
	wire w_dff_A_pFaqW4Nf0_0;
	wire w_dff_A_QtnwI8EJ5_2;
	wire w_dff_A_spW4h4da2_0;
	wire w_dff_A_gbFP4Yft7_0;
	wire w_dff_A_OxXuaSf93_0;
	wire w_dff_A_JJjKsZ4p2_1;
	wire w_dff_A_m7f1IMZA8_1;
	wire w_dff_B_rUjrGK0s1_2;
	wire w_dff_B_qtDbI3Zt3_2;
	wire w_dff_B_EToVaKBN7_2;
	wire w_dff_B_mmKJ5qqi8_2;
	wire w_dff_B_MeCVlgJM3_0;
	wire w_dff_A_3LGUGYRd9_0;
	wire w_dff_A_EsLHXE3L0_0;
	wire w_dff_B_xe2q5kHB6_0;
	wire w_dff_A_XqHtVFsO4_1;
	wire w_dff_A_W1c1TVdY3_1;
	wire w_dff_A_9YLdQILM7_1;
	wire w_dff_A_3C4k9QRd6_1;
	wire w_dff_A_Dm3H6giZ3_1;
	wire w_dff_A_qsl1bnTk2_1;
	wire w_dff_A_Q65ouTAs2_1;
	wire w_dff_A_SozBqppf7_1;
	wire w_dff_A_lPLd9Pn27_1;
	wire w_dff_A_7k64b6kS6_1;
	wire w_dff_A_dKiqw83U8_1;
	wire w_dff_A_hW804BSL3_1;
	wire w_dff_A_eI78CFqv4_1;
	wire w_dff_A_3QYhKI754_1;
	wire w_dff_A_3QvyCeFi8_1;
	wire w_dff_A_CemPURmK5_1;
	wire w_dff_A_eXwJdX2V7_1;
	wire w_dff_A_mNaXwtfb0_1;
	wire w_dff_A_jfCAJBeO5_1;
	wire w_dff_A_y1U3RlEq9_1;
	wire w_dff_A_tS7ni6pF2_2;
	wire w_dff_A_sHcYbj7c1_2;
	wire w_dff_A_YaR9Amxy9_2;
	wire w_dff_A_oS1obBMh2_2;
	wire w_dff_A_Am7Ml6aC2_2;
	wire w_dff_A_lnV5gdjH3_2;
	wire w_dff_A_OMzKAEPm8_2;
	wire w_dff_A_k6jXxjeM9_2;
	wire w_dff_A_vNKgmZij1_2;
	wire w_dff_A_CLRnVBti7_2;
	wire w_dff_A_W5CMpLB79_2;
	wire w_dff_A_v0x2Em3E2_2;
	wire w_dff_A_xtkQUYuL6_0;
	wire w_dff_A_KdmmqOod6_0;
	wire w_dff_A_lmLj9Lys5_0;
	wire w_dff_A_hDrs1Hc01_0;
	wire w_dff_A_WnumbqER2_0;
	wire w_dff_A_ladQDdBe3_0;
	wire w_dff_A_xG3u0NB46_0;
	wire w_dff_A_DUrS3OY56_0;
	wire w_dff_A_89cFRmeR0_0;
	wire w_dff_A_J3g2x2e91_0;
	wire w_dff_A_DQsXNwKp4_0;
	wire w_dff_A_liEfg0Qt9_0;
	wire w_dff_A_DGHc9F6a3_0;
	wire w_dff_A_SJjSEmZ87_0;
	wire w_dff_A_9t8R4aYe8_0;
	wire w_dff_A_DJVy1Vj43_0;
	wire w_dff_A_P4z0Z6u07_0;
	wire w_dff_A_JFbBJjwL8_0;
	wire w_dff_A_2Vs49HL71_2;
	wire w_dff_A_Zvluu8NA5_0;
	wire w_dff_A_vfa2d84t6_0;
	wire w_dff_A_9n1AUUg50_0;
	wire w_dff_A_xDP9o8427_0;
	wire w_dff_A_mXAxSiCI5_0;
	wire w_dff_A_f0lOnMoU3_0;
	wire w_dff_A_n8OxAATE0_0;
	wire w_dff_A_jCUKFyHl9_0;
	wire w_dff_A_0aUvTdKl0_0;
	wire w_dff_A_rQd0gKmE4_0;
	wire w_dff_A_G6W5veAp4_0;
	wire w_dff_A_MkuOaLul8_0;
	wire w_dff_A_7bMKgShr7_0;
	wire w_dff_A_hPT0rcx76_0;
	wire w_dff_A_aqE72HcN8_0;
	wire w_dff_A_WManN0r55_0;
	wire w_dff_A_4cToR0fG3_0;
	wire w_dff_A_hft1OadK4_0;
	wire w_dff_A_CX6SNnSY4_2;
	wire w_dff_A_E4w2Cg7B7_0;
	wire w_dff_A_sJiKNRuu5_0;
	wire w_dff_A_LYXWeyiV4_0;
	wire w_dff_A_IVzQps155_0;
	wire w_dff_A_XYs2lv1G6_0;
	wire w_dff_A_lsVcQylp4_0;
	wire w_dff_A_nriLEvHh8_0;
	wire w_dff_A_iymqAfR47_0;
	wire w_dff_A_RGoTqBv61_0;
	wire w_dff_A_9wsH7zyo4_0;
	wire w_dff_A_J8nQqiQK1_0;
	wire w_dff_A_AuJeQc7Z9_0;
	wire w_dff_A_9trUj2dj2_0;
	wire w_dff_A_ZYTG7bga4_0;
	wire w_dff_A_VkeoxyuL1_0;
	wire w_dff_A_E1YH34Hz8_0;
	wire w_dff_A_rT324FG03_0;
	wire w_dff_A_iUxU1lmx4_0;
	wire w_dff_A_Xh2ELakS9_2;
	wire w_dff_A_RcxGboRk1_0;
	wire w_dff_A_wYF4a9w83_0;
	wire w_dff_A_JHzzZ78h0_0;
	wire w_dff_A_uSIQMkia0_0;
	wire w_dff_A_PrbXm2LQ2_0;
	wire w_dff_A_ivyqjlCB7_0;
	wire w_dff_A_U2ptytqh7_0;
	wire w_dff_A_xEV7E2Dx5_0;
	wire w_dff_A_pECFW0EF4_0;
	wire w_dff_A_nMDLpxkd2_0;
	wire w_dff_A_HTPJ8ZFe9_0;
	wire w_dff_A_hJzaNZo99_0;
	wire w_dff_A_XA9uKdIl9_0;
	wire w_dff_A_WCkSSlC85_0;
	wire w_dff_A_WbkkA9fY0_0;
	wire w_dff_A_u7QlEQN13_0;
	wire w_dff_A_WReXI3mr5_0;
	wire w_dff_A_GBtaoWwc3_0;
	wire w_dff_A_itv1kqrl8_0;
	wire w_dff_A_FDWFIrl16_2;
	wire w_dff_A_D5WWLe269_0;
	wire w_dff_A_D1ILTAvo4_0;
	wire w_dff_A_3K0vDBkf2_0;
	wire w_dff_A_5kUjCC0O9_0;
	wire w_dff_A_ows4u9JO5_0;
	wire w_dff_A_uVPYN4iP4_0;
	wire w_dff_A_kzKSYTzO7_0;
	wire w_dff_A_WSNnWOHh0_0;
	wire w_dff_A_KyyocGZe6_0;
	wire w_dff_A_THNrH40Q5_0;
	wire w_dff_A_qXSwfnKp8_0;
	wire w_dff_A_5XdKHzDI6_0;
	wire w_dff_A_bt9xHAmH3_0;
	wire w_dff_A_0SO10ped5_0;
	wire w_dff_A_0Cl95lyv3_0;
	wire w_dff_A_tinlgHgA4_0;
	wire w_dff_A_imctwPHn3_0;
	wire w_dff_A_QRMKaVJk5_0;
	wire w_dff_A_tqHLL7uK6_2;
	wire w_dff_A_KACSFeVn6_0;
	wire w_dff_A_IJbXFV4b9_0;
	wire w_dff_A_AiP1ikyE7_0;
	wire w_dff_A_tH3EmEVv1_0;
	wire w_dff_A_jTuRkaIz4_0;
	wire w_dff_A_n3cnsbSD6_0;
	wire w_dff_A_CJlwXQdA8_0;
	wire w_dff_A_3AKbhcvO5_0;
	wire w_dff_A_mJodgsau7_0;
	wire w_dff_A_HfTbvByc6_0;
	wire w_dff_A_anntVTbu3_0;
	wire w_dff_A_MMJYSJ0X6_0;
	wire w_dff_A_F5vSktkQ3_0;
	wire w_dff_A_asiu61cE3_0;
	wire w_dff_A_TiJ0vDt26_0;
	wire w_dff_A_Q9Mm0WCy1_0;
	wire w_dff_A_3Vj6ap9D4_2;
	wire w_dff_A_wNpyU6gF4_0;
	wire w_dff_A_wxn9bf7a8_0;
	wire w_dff_A_T9CsQu4l1_0;
	wire w_dff_A_d5QdZfZp7_0;
	wire w_dff_A_y8Yu9Aez5_0;
	wire w_dff_A_2EvaerIa6_0;
	wire w_dff_A_CjJUkOXJ7_0;
	wire w_dff_A_FOww7t603_0;
	wire w_dff_A_X2QbrQik8_0;
	wire w_dff_A_25avs1oa0_0;
	wire w_dff_A_tecoaT1k6_0;
	wire w_dff_A_4UgBqPiN4_0;
	wire w_dff_A_kfZWxZa49_0;
	wire w_dff_A_a5YZHejn2_0;
	wire w_dff_A_eyzhNh3I2_0;
	wire w_dff_A_IaD2PxtD0_0;
	wire w_dff_A_kZ9MkF7H9_0;
	wire w_dff_A_XFUZnNOl3_2;
	wire w_dff_A_rPTjTisk5_0;
	wire w_dff_A_p5xzbR8Z7_0;
	wire w_dff_A_XNugZ0bg6_0;
	wire w_dff_A_3q1Aja3K1_0;
	wire w_dff_A_UrIQz1AP4_0;
	wire w_dff_A_du7xO8RR3_0;
	wire w_dff_A_kjdfwjxG3_0;
	wire w_dff_A_9AXVyoWV3_0;
	wire w_dff_A_X0u2I49y7_0;
	wire w_dff_A_6tq8lMEF6_0;
	wire w_dff_A_6SniNiZx7_0;
	wire w_dff_A_lxLJ1r8X9_0;
	wire w_dff_A_PpOKEoAJ1_0;
	wire w_dff_A_P1ybqFjO2_0;
	wire w_dff_A_4zWGkNDC0_0;
	wire w_dff_A_fvTmgAWN7_0;
	wire w_dff_A_ODiXCupA7_0;
	wire w_dff_A_g6bXiTJg5_2;
	wire w_dff_A_mcPsRd1K9_0;
	wire w_dff_A_hN4nzfMg3_0;
	wire w_dff_A_wfoY278h7_0;
	wire w_dff_A_axWIUTCu1_0;
	wire w_dff_A_xZA8gvVV4_0;
	wire w_dff_A_0ex4AtiZ6_0;
	wire w_dff_A_oaK77J3U7_0;
	wire w_dff_A_Ibf4GOqP4_0;
	wire w_dff_A_y82YZVhN4_0;
	wire w_dff_A_sCzAckFO8_0;
	wire w_dff_A_c82g1weT7_0;
	wire w_dff_A_Ucp7WZ6P4_0;
	wire w_dff_A_kw1IApWj5_0;
	wire w_dff_A_RLRdFeb08_0;
	wire w_dff_A_aQ99LbxA2_0;
	wire w_dff_A_eM4weOKO9_0;
	wire w_dff_A_2Z61ps791_0;
	wire w_dff_A_2F8BBGCp1_2;
	wire w_dff_A_8ab2RlK79_0;
	wire w_dff_A_hE6bpMsx8_0;
	wire w_dff_A_h5cCdXKr6_0;
	wire w_dff_A_nWQERbPz9_0;
	wire w_dff_A_IpZ0lVAO4_0;
	wire w_dff_A_tW4eTduQ6_0;
	wire w_dff_A_AVG8HZr79_0;
	wire w_dff_A_D65CF86p1_0;
	wire w_dff_A_oJTu87Dn6_0;
	wire w_dff_A_8Xr1gNFM8_0;
	wire w_dff_A_tHBMkvBX5_0;
	wire w_dff_A_ALvt2Tr15_0;
	wire w_dff_A_4bYeS8tP7_0;
	wire w_dff_A_AZUh64Lp7_0;
	wire w_dff_A_WFk6BzR51_0;
	wire w_dff_A_ZRHcwRTJ9_0;
	wire w_dff_A_YZvl8Xfh8_0;
	wire w_dff_A_Jy0JyhUZ8_0;
	wire w_dff_A_NowZgrpN0_2;
	wire w_dff_A_ez5JPiF32_0;
	wire w_dff_A_aJhmc3KS9_0;
	wire w_dff_A_Mqbvvkrg6_0;
	wire w_dff_A_ua8wzgOT2_0;
	wire w_dff_A_y8GMdNal9_0;
	wire w_dff_A_7abAmPvm7_0;
	wire w_dff_A_vRKz4I905_0;
	wire w_dff_A_hJ98fB685_0;
	wire w_dff_A_ps25jzSs5_0;
	wire w_dff_A_Xe6d9Sok1_0;
	wire w_dff_A_mQzREqH25_0;
	wire w_dff_A_V9ltStEh0_0;
	wire w_dff_A_hMqEYEQA0_0;
	wire w_dff_A_zhbMisoT8_0;
	wire w_dff_A_BMLBQxe45_0;
	wire w_dff_A_0R5U5ofJ9_0;
	wire w_dff_A_wbw40VA04_1;
	wire w_dff_A_RWWMBmUX0_0;
	wire w_dff_A_Y9HYAg1j0_0;
	wire w_dff_A_pFwygKjG0_0;
	wire w_dff_A_XQlQGsfQ8_0;
	wire w_dff_A_NtPzn7Qf6_0;
	wire w_dff_A_JseRuWVB6_0;
	wire w_dff_A_LNObQEut7_0;
	wire w_dff_A_ncz4YBQL5_0;
	wire w_dff_A_VYVtXc3e4_0;
	wire w_dff_A_X8vKrcpy5_0;
	wire w_dff_A_V4wPDe5y5_0;
	wire w_dff_A_c0InGZ4f6_0;
	wire w_dff_A_ZJF1DjtW6_0;
	wire w_dff_A_tKPTQEpc5_0;
	wire w_dff_A_FtQx97CX7_0;
	wire w_dff_A_4TUbB0vq3_0;
	wire w_dff_A_orJTJbDA6_0;
	wire w_dff_A_J8xnWMmK8_0;
	wire w_dff_A_vEUawqo43_2;
	wire w_dff_A_U977mjRo7_0;
	wire w_dff_A_lCKS3kqa6_0;
	wire w_dff_A_OMh5MYx10_0;
	wire w_dff_A_wPmuxMqR3_0;
	wire w_dff_A_7BDasKBt7_0;
	wire w_dff_A_V8PNeLYQ6_0;
	wire w_dff_A_jx1ARsVy3_0;
	wire w_dff_A_EtJyfVQ54_0;
	wire w_dff_A_Mtk3Onhd8_0;
	wire w_dff_A_DiFH2RKg5_0;
	wire w_dff_A_7rYLz2Pt3_0;
	wire w_dff_A_7hPpqPks9_0;
	wire w_dff_A_oz5oGohB1_0;
	wire w_dff_A_4z4pNh510_0;
	wire w_dff_A_hqi8BIDZ9_0;
	wire w_dff_A_Im0opok21_0;
	wire w_dff_A_O1IwgoSl3_0;
	wire w_dff_A_pKviZhew7_2;
	wire w_dff_A_WUwHDdlA5_0;
	wire w_dff_A_MLBTSbsZ3_0;
	wire w_dff_A_rpJgTuYi0_0;
	wire w_dff_A_wK7XOcnt3_0;
	wire w_dff_A_lev5a7F41_0;
	wire w_dff_A_UJJdBNSA1_0;
	wire w_dff_A_1t61mpq78_0;
	wire w_dff_A_Uta5chsW1_0;
	wire w_dff_A_83cjwK6v0_0;
	wire w_dff_A_FH7ENENa4_0;
	wire w_dff_A_CaQfbgwv1_0;
	wire w_dff_A_9aTiXfNm9_0;
	wire w_dff_A_fGAdYluU9_0;
	wire w_dff_A_KFEV1lyz5_0;
	wire w_dff_A_Of2s9mnT3_0;
	wire w_dff_A_vTgbgUFr0_0;
	wire w_dff_A_MsihI2xx3_0;
	wire w_dff_A_DXYPJYMd4_2;
	wire w_dff_A_N7fzxBil4_0;
	wire w_dff_A_LZTHB2zd1_0;
	wire w_dff_A_aVmaBTBD5_0;
	wire w_dff_A_0RK32nxr3_0;
	wire w_dff_A_XoEkWgyZ5_0;
	wire w_dff_A_RTHDuTM76_0;
	wire w_dff_A_eaZyWBaK5_0;
	wire w_dff_A_4FoVSiQL7_0;
	wire w_dff_A_Loi7ElGu3_0;
	wire w_dff_A_5Xz8bkrc5_0;
	wire w_dff_A_0ksjWoiW1_0;
	wire w_dff_A_yS1bS6Kz8_0;
	wire w_dff_A_tIx92P8k7_0;
	wire w_dff_A_5dtrpx958_0;
	wire w_dff_A_d34oFi6j6_0;
	wire w_dff_A_NUPHI5O48_0;
	wire w_dff_A_z2k2FgAq9_0;
	wire w_dff_A_qE32jqNx9_0;
	wire w_dff_A_OLTbHvvH0_2;
	wire w_dff_A_7LwcjK0y0_0;
	wire w_dff_A_XYr7xw2H7_0;
	wire w_dff_A_QJtNXSHq5_0;
	wire w_dff_A_OOk4ScND3_0;
	wire w_dff_A_8Fg2Lyhj1_0;
	wire w_dff_A_XMianCNc7_0;
	wire w_dff_A_fNWX4ibp4_0;
	wire w_dff_A_oWhyp7Er3_0;
	wire w_dff_A_RF5GxOWV6_0;
	wire w_dff_A_zNJCibHF9_0;
	wire w_dff_A_6Bnlvj034_0;
	wire w_dff_A_tt1CmXvZ1_0;
	wire w_dff_A_7BoktcCx1_0;
	wire w_dff_A_NRtespHK1_0;
	wire w_dff_A_FScb5QMa7_0;
	wire w_dff_A_xRMhYuOI2_0;
	wire w_dff_A_eFK7LroM1_2;
	wire w_dff_A_sZxFQNy83_0;
	wire w_dff_A_X6bNZAtW3_0;
	wire w_dff_A_Oyh92nqn6_0;
	wire w_dff_A_WKw2PRZy7_0;
	wire w_dff_A_HKqw4KX41_0;
	wire w_dff_A_v4nydyvP1_0;
	wire w_dff_A_VUMnKgYs3_0;
	wire w_dff_A_wlkJxLG59_0;
	wire w_dff_A_SLq7dLTq7_0;
	wire w_dff_A_rK3mPQif7_0;
	wire w_dff_A_vztwDrbc9_0;
	wire w_dff_A_cDf4RW9v0_0;
	wire w_dff_A_dmMIlVwQ1_0;
	wire w_dff_A_T894taxk0_0;
	wire w_dff_A_zSOToXXM2_0;
	wire w_dff_A_s3u7Ckjo0_0;
	wire w_dff_A_pS0wowaN6_2;
	wire w_dff_A_ks4a92Wh9_0;
	wire w_dff_A_0vVOKW4o9_0;
	wire w_dff_A_mvXaCdjZ6_0;
	wire w_dff_A_b5KCODrM2_0;
	wire w_dff_A_wL26Jx331_0;
	wire w_dff_A_hp7UmHj04_0;
	wire w_dff_A_jfC4LkO81_0;
	wire w_dff_A_uKd4HO2L8_2;
	wire w_dff_A_HgCi46kM4_0;
	wire w_dff_A_YpNUobZl3_0;
	wire w_dff_A_rAiVBEsX2_0;
	wire w_dff_A_osBm35gL3_2;
	wire w_dff_A_SF9iIUlC6_0;
	wire w_dff_A_5JSJaS396_0;
	wire w_dff_A_aatVJbvH0_0;
	wire w_dff_A_TGjlIEZu5_2;
	wire w_dff_A_OZvexL6z0_0;
	wire w_dff_A_2fore71h0_0;
	wire w_dff_A_hncFd4F85_0;
	wire w_dff_A_ZHe4fB7d1_0;
	wire w_dff_A_Hj0sHmmF5_0;
	wire w_dff_A_pjkRVhk99_2;
	wire w_dff_A_Ve8CQfh89_0;
	wire w_dff_A_cQvl11VV9_2;
	wire w_dff_A_X7xuBf9F5_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_v0x2Em3E2_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_2Vs49HL71_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_Xh2ELakS9_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_G17gat_2[2]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_n92_0[2]),.dout(w_dff_A_FDWFIrl16_2),.clk(gclk));
	jnot g009(.din(w_n93_0[0]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G1gat_1[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G26gat_0[1]),.dout(n97),.clk(gclk));
	jor g012(.dina(n97),.dinb(w_n96_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(w_n98_0[1]),.dinb(n95),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_tqHLL7uK6_2),.clk(gclk));
	jnot g015(.din(w_G80gat_0[1]),.dout(n101),.clk(gclk));
	jand g016(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n102),.clk(gclk));
	jnot g017(.din(w_n102_0[1]),.dout(n103),.clk(gclk));
	jor g018(.dina(n103),.dinb(w_n101_0[1]),.dout(w_dff_A_3Vj6ap9D4_2),.clk(gclk));
	jnot g019(.din(w_G36gat_0[0]),.dout(n105),.clk(gclk));
	jnot g020(.din(w_G59gat_1[0]),.dout(n106),.clk(gclk));
	jor g021(.dina(w_n106_0[1]),.dinb(n105),.dout(n107),.clk(gclk));
	jor g022(.dina(w_n107_0[1]),.dinb(w_n101_0[0]),.dout(w_dff_A_XFUZnNOl3_2),.clk(gclk));
	jnot g023(.din(w_G42gat_1[2]),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n107_0[0]),.dinb(w_dff_B_iugJthxE1_1),.dout(w_dff_A_g6bXiTJg5_2),.clk(gclk));
	jor g025(.dina(G88gat),.dinb(G87gat),.dout(n111),.clk(gclk));
	jand g026(.dina(w_n111_0[1]),.dinb(w_dff_B_tDtNnlHu9_1),.dout(w_dff_A_2F8BBGCp1_2),.clk(gclk));
	jnot g027(.din(w_G390gat_0[0]),.dout(n113),.clk(gclk));
	jor g028(.dina(w_n99_0[0]),.dinb(n113),.dout(w_dff_A_NowZgrpN0_2),.clk(gclk));
	jand g029(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n115),.clk(gclk));
	jand g030(.dina(n115),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g031(.dina(w_G55gat_0[2]),.dinb(w_G13gat_0[0]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_n92_0[1]),.dout(n118),.clk(gclk));
	jand g033(.dina(w_G68gat_0[1]),.dinb(w_G29gat_0[0]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_dff_B_2w2NwKet5_0),.dinb(w_n118_0[2]),.dout(w_dff_A_vEUawqo43_2),.clk(gclk));
	jand g035(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n121),.clk(gclk));
	jand g036(.dina(w_n121_0[1]),.dinb(w_dff_B_GdgUF8cQ0_1),.dout(n122),.clk(gclk));
	jand g037(.dina(n122),.dinb(w_n118_0[1]),.dout(w_dff_A_pKviZhew7_2),.clk(gclk));
	jand g038(.dina(w_n111_0[0]),.dinb(w_dff_B_WLWUl7eF7_1),.dout(w_dff_A_DXYPJYMd4_2),.clk(gclk));
	jxor g039(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n125),.clk(gclk));
	jxor g040(.dina(n125),.dinb(w_G130gat_0[1]),.dout(n126),.clk(gclk));
	jxor g041(.dina(w_G126gat_0[1]),.dinb(w_G121gat_0[2]),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_dff_B_ESnsRQaR5_0),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g043(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n129),.clk(gclk));
	jxor g044(.dina(n129),.dinb(w_dff_B_bU6U96DH3_1),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(w_dff_B_xwH9UetB0_0),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n128),.dout(w_dff_A_OLTbHvvH0_2),.clk(gclk));
	jxor g048(.dina(w_G165gat_2[1]),.dinb(w_G159gat_2[1]),.dout(n134),.clk(gclk));
	jxor g049(.dina(n134),.dinb(w_G130gat_0[0]),.dout(n135),.clk(gclk));
	jxor g050(.dina(w_G201gat_2[2]),.dinb(w_G195gat_2[1]),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_dff_B_PNiG9O2k8_0),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g052(.dina(w_G189gat_2[1]),.dinb(w_G183gat_2[1]),.dout(n138),.clk(gclk));
	jxor g053(.dina(n138),.dinb(w_dff_B_4fXyhJE60_1),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G177gat_2[1]),.dinb(w_G171gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(w_dff_B_8vDVZbqX9_0),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n137),.dout(w_dff_A_eFK7LroM1_2),.clk(gclk));
	jnot g057(.din(w_G261gat_0[2]),.dout(n143),.clk(gclk));
	jand g058(.dina(w_n102_0[0]),.dinb(w_G42gat_1[1]),.dout(n144),.clk(gclk));
	jnot g059(.din(n144),.dout(n145),.clk(gclk));
	jand g060(.dina(w_G51gat_1[0]),.dinb(w_G17gat_2[1]),.dout(n146),.clk(gclk));
	jand g061(.dina(n146),.dinb(w_n92_0[0]),.dout(n147),.clk(gclk));
	jand g062(.dina(w_dff_B_xe2q5kHB6_0),.dinb(n145),.dout(n148),.clk(gclk));
	jand g063(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n149),.clk(gclk));
	jxor g064(.dina(w_G42gat_1[0]),.dinb(w_G17gat_2[0]),.dout(n150),.clk(gclk));
	jand g065(.dina(n150),.dinb(w_n149_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(n151),.dinb(w_G447gat_1),.dout(n152),.clk(gclk));
	jor g067(.dina(w_dff_B_MeCVlgJM3_0),.dinb(n148),.dout(n153),.clk(gclk));
	jand g068(.dina(w_n153_3[1]),.dinb(w_G126gat_0[0]),.dout(n154),.clk(gclk));
	jnot g069(.din(w_G156gat_0[0]),.dout(n155),.clk(gclk));
	jor g070(.dina(n155),.dinb(w_n106_0[0]),.dout(n156),.clk(gclk));
	jand g071(.dina(n156),.dinb(w_G447gat_0[2]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n157_0[1]),.dinb(w_G17gat_1[2]),.dout(n158),.clk(gclk));
	jor g073(.dina(n158),.dinb(w_n96_0[0]),.dout(n159),.clk(gclk));
	jand g074(.dina(w_n159_1[1]),.dinb(w_G153gat_0[2]),.dout(n160),.clk(gclk));
	jand g075(.dina(w_n86_0[0]),.dinb(w_G80gat_0[0]),.dout(n161),.clk(gclk));
	jand g076(.dina(n161),.dinb(w_G447gat_0[1]),.dout(n162),.clk(gclk));
	jnot g077(.din(w_G268gat_0[1]),.dout(n163),.clk(gclk));
	jand g078(.dina(w_n163_0[1]),.dinb(w_G55gat_0[1]),.dout(n164),.clk(gclk));
	jand g079(.dina(w_dff_B_YXTVlwAl6_0),.dinb(w_n162_0[1]),.dout(n165),.clk(gclk));
	jor g080(.dina(w_n165_1[2]),.dinb(n160),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n154_0[1]),.dout(n167),.clk(gclk));
	jxor g082(.dina(w_n167_1[1]),.dinb(w_G201gat_2[1]),.dout(n168),.clk(gclk));
	jnot g083(.din(w_n168_0[2]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n143_0[1]),.dout(n170),.clk(gclk));
	jor g085(.dina(w_n168_0[1]),.dinb(w_G261gat_0[1]),.dout(n171),.clk(gclk));
	jand g086(.dina(n171),.dinb(w_G219gat_3[1]),.dout(n172),.clk(gclk));
	jand g087(.dina(n172),.dinb(n170),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n168_0[0]),.dinb(w_G228gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_G237gat_3[1]),.dinb(w_G201gat_2[0]),.dout(n175),.clk(gclk));
	jor g090(.dina(n175),.dinb(w_G246gat_3[1]),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_LAkMJVPZ7_0),.dinb(w_n167_1[0]),.dout(n177),.clk(gclk));
	jand g092(.dina(G72gat),.dinb(w_G42gat_0[2]),.dout(n178),.clk(gclk));
	jand g093(.dina(n178),.dinb(w_dff_B_v1xyCebV4_1),.dout(n179),.clk(gclk));
	jand g094(.dina(n179),.dinb(w_n121_0[0]),.dout(n180),.clk(gclk));
	jand g095(.dina(n180),.dinb(w_n118_0[0]),.dout(n181),.clk(gclk));
	jand g096(.dina(w_n181_3[1]),.dinb(w_G201gat_1[2]),.dout(n182),.clk(gclk));
	jand g097(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n183),.clk(gclk));
	jand g098(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(n184),.dinb(n183),.dout(n185),.clk(gclk));
	jor g100(.dina(w_dff_B_auSpZ2Q82_0),.dinb(n182),.dout(n186),.clk(gclk));
	jor g101(.dina(w_dff_B_mzqr1oNS7_0),.dinb(n177),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(n174),.dout(n188),.clk(gclk));
	jor g103(.dina(w_dff_B_6PGRgfmA5_0),.dinb(n173),.dout(w_dff_A_pS0wowaN6_2),.clk(gclk));
	jand g104(.dina(w_n159_1[0]),.dinb(w_G143gat_0[1]),.dout(n190),.clk(gclk));
	jand g105(.dina(w_n153_3[0]),.dinb(w_G111gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(n191),.dinb(w_n165_1[1]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_dff_B_41bkNbQJ2_1),.dout(n193),.clk(gclk));
	jxor g108(.dina(w_n193_1[1]),.dinb(w_G183gat_2[0]),.dout(n194),.clk(gclk));
	jnot g109(.din(w_n194_0[2]),.dout(n195),.clk(gclk));
	jand g110(.dina(w_n167_0[2]),.dinb(w_G201gat_1[1]),.dout(n196),.clk(gclk));
	jnot g111(.din(w_n196_0[1]),.dout(n197),.clk(gclk));
	jnot g112(.din(w_G201gat_1[0]),.dout(n198),.clk(gclk));
	jnot g113(.din(w_n154_0[0]),.dout(n199),.clk(gclk));
	jnot g114(.din(w_G153gat_0[1]),.dout(n200),.clk(gclk));
	jnot g115(.din(w_G17gat_1[1]),.dout(n201),.clk(gclk));
	jnot g116(.din(w_G51gat_0[2]),.dout(n202),.clk(gclk));
	jor g117(.dina(w_n98_0[0]),.dinb(w_dff_B_WPPIywU42_1),.dout(n203),.clk(gclk));
	jor g118(.dina(w_n149_0[0]),.dinb(n203),.dout(n204),.clk(gclk));
	jor g119(.dina(n204),.dinb(w_dff_B_AYIgoPJz7_1),.dout(n205),.clk(gclk));
	jand g120(.dina(n205),.dinb(w_G1gat_0[1]),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(w_dff_B_vr0TsmQz8_1),.dout(n207),.clk(gclk));
	jnot g122(.din(w_n165_1[0]),.dout(n208),.clk(gclk));
	jand g123(.dina(w_dff_B_7ZCE6cac4_0),.dinb(n207),.dout(n209),.clk(gclk));
	jand g124(.dina(n209),.dinb(w_dff_B_ZEfKWUgn0_1),.dout(n210),.clk(gclk));
	jand g125(.dina(n210),.dinb(w_dff_B_kgLBemVM5_1),.dout(n211),.clk(gclk));
	jor g126(.dina(n211),.dinb(w_n143_0[0]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_clXIMNx08_1),.dout(n213),.clk(gclk));
	jand g128(.dina(w_n159_0[2]),.dinb(w_G146gat_0[1]),.dout(n214),.clk(gclk));
	jand g129(.dina(w_n153_2[2]),.dinb(w_G116gat_0[1]),.dout(n215),.clk(gclk));
	jor g130(.dina(n215),.dinb(w_n165_0[2]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_dff_B_aqjt3HhL1_1),.dout(n217),.clk(gclk));
	jor g132(.dina(w_n217_1[1]),.dinb(w_G189gat_2[0]),.dout(n218),.clk(gclk));
	jand g133(.dina(w_n159_0[1]),.dinb(w_G149gat_0[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n153_2[1]),.dinb(w_G121gat_0[0]),.dout(n220),.clk(gclk));
	jor g135(.dina(n220),.dinb(w_n165_0[1]),.dout(n221),.clk(gclk));
	jor g136(.dina(n221),.dinb(w_dff_B_uESYCf1D5_1),.dout(n222),.clk(gclk));
	jor g137(.dina(w_n222_1[1]),.dinb(w_G195gat_2[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n223_0[1]),.dinb(w_n218_0[1]),.dout(n224),.clk(gclk));
	jnot g139(.din(w_n224_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_TEqq0CvK2_0),.dinb(w_n213_0[1]),.dout(n226),.clk(gclk));
	jand g141(.dina(w_n217_1[0]),.dinb(w_G189gat_1[2]),.dout(n227),.clk(gclk));
	jand g142(.dina(w_n222_1[0]),.dinb(w_G195gat_1[2]),.dout(n228),.clk(gclk));
	jand g143(.dina(w_n228_0[1]),.dinb(w_n218_0[0]),.dout(n229),.clk(gclk));
	jor g144(.dina(n229),.dinb(w_dff_B_QlEQ6RiZ3_1),.dout(n230),.clk(gclk));
	jnot g145(.din(w_n230_0[1]),.dout(n231),.clk(gclk));
	jand g146(.dina(w_dff_B_q2cswN5H8_0),.dinb(n226),.dout(n232),.clk(gclk));
	jor g147(.dina(w_n232_0[1]),.dinb(w_dff_B_FmOh0vb39_1),.dout(n233),.clk(gclk));
	jor g148(.dina(w_n167_0[1]),.dinb(w_G201gat_0[2]),.dout(n234),.clk(gclk));
	jand g149(.dina(n234),.dinb(w_G261gat_0[0]),.dout(n235),.clk(gclk));
	jor g150(.dina(n235),.dinb(w_n196_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n224_0[0]),.dinb(w_n236_0[2]),.dout(n237),.clk(gclk));
	jor g152(.dina(w_n230_0[0]),.dinb(n237),.dout(n238),.clk(gclk));
	jor g153(.dina(w_n238_0[1]),.dinb(w_n194_0[1]),.dout(n239),.clk(gclk));
	jand g154(.dina(n239),.dinb(w_G219gat_3[0]),.dout(n240),.clk(gclk));
	jand g155(.dina(n240),.dinb(n233),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n194_0[0]),.dinb(w_G228gat_3[0]),.dout(n242),.clk(gclk));
	jand g157(.dina(w_G237gat_3[0]),.dinb(w_G183gat_1[2]),.dout(n243),.clk(gclk));
	jor g158(.dina(n243),.dinb(w_G246gat_3[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(w_dff_B_jzXK16sE8_0),.dinb(w_n193_1[0]),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n181_3[0]),.dinb(w_G183gat_1[1]),.dout(n246),.clk(gclk));
	jand g161(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n247),.clk(gclk));
	jor g162(.dina(w_dff_B_FPQEmp059_0),.dinb(n246),.dout(n248),.clk(gclk));
	jor g163(.dina(w_dff_B_ZTIf6Wlo2_0),.dinb(n245),.dout(n249),.clk(gclk));
	jor g164(.dina(n249),.dinb(n242),.dout(n250),.clk(gclk));
	jor g165(.dina(w_dff_B_tMPfvelr4_0),.dinb(n241),.dout(w_dff_A_uKd4HO2L8_2),.clk(gclk));
	jxor g166(.dina(w_n217_0[2]),.dinb(w_G189gat_1[1]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n252_0[2]),.dout(n253),.clk(gclk));
	jand g168(.dina(w_n223_0[0]),.dinb(w_n236_0[1]),.dout(n254),.clk(gclk));
	jor g169(.dina(n254),.dinb(w_n228_0[0]),.dout(n255),.clk(gclk));
	jnot g170(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jor g171(.dina(n256),.dinb(w_dff_B_7RiwbCrg6_1),.dout(n257),.clk(gclk));
	jor g172(.dina(w_n255_0[0]),.dinb(w_n252_0[1]),.dout(n258),.clk(gclk));
	jand g173(.dina(n258),.dinb(w_G219gat_2[2]),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(n257),.dout(n260),.clk(gclk));
	jand g175(.dina(w_n252_0[0]),.dinb(w_G228gat_2[2]),.dout(n261),.clk(gclk));
	jand g176(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n262),.clk(gclk));
	jor g177(.dina(n262),.dinb(w_G246gat_2[2]),.dout(n263),.clk(gclk));
	jand g178(.dina(w_dff_B_wyNBG4UK4_0),.dinb(w_n217_0[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(w_n181_2[2]),.dinb(w_G189gat_0[2]),.dout(n265),.clk(gclk));
	jand g180(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n266),.clk(gclk));
	jand g181(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n267),.clk(gclk));
	jor g182(.dina(n267),.dinb(n266),.dout(n268),.clk(gclk));
	jor g183(.dina(w_dff_B_gQ6iSmGV4_0),.dinb(n265),.dout(n269),.clk(gclk));
	jor g184(.dina(w_dff_B_xrA1lCIC7_0),.dinb(n264),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(n261),.dout(n271),.clk(gclk));
	jor g186(.dina(w_dff_B_sot1kt8j9_0),.dinb(n260),.dout(w_dff_A_osBm35gL3_2),.clk(gclk));
	jxor g187(.dina(w_n222_0[2]),.dinb(w_G195gat_1[1]),.dout(n273),.clk(gclk));
	jnot g188(.din(w_n273_0[2]),.dout(n274),.clk(gclk));
	jor g189(.dina(w_dff_B_5J4qcP2F2_0),.dinb(w_n213_0[0]),.dout(n275),.clk(gclk));
	jor g190(.dina(w_n273_0[1]),.dinb(w_n236_0[0]),.dout(n276),.clk(gclk));
	jand g191(.dina(n276),.dinb(w_G219gat_2[1]),.dout(n277),.clk(gclk));
	jand g192(.dina(n277),.dinb(n275),.dout(n278),.clk(gclk));
	jand g193(.dina(w_n273_0[0]),.dinb(w_G228gat_2[1]),.dout(n279),.clk(gclk));
	jand g194(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(n280),.dinb(w_G246gat_2[1]),.dout(n281),.clk(gclk));
	jand g196(.dina(w_dff_B_VSJf4baY0_0),.dinb(w_n222_0[1]),.dout(n282),.clk(gclk));
	jand g197(.dina(w_n181_2[1]),.dinb(w_G195gat_0[2]),.dout(n283),.clk(gclk));
	jand g198(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n284),.clk(gclk));
	jand g199(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n285),.clk(gclk));
	jor g200(.dina(n285),.dinb(n284),.dout(n286),.clk(gclk));
	jor g201(.dina(w_dff_B_EkS5AOkG9_0),.dinb(n283),.dout(n287),.clk(gclk));
	jor g202(.dina(w_dff_B_nmyHmH251_0),.dinb(n282),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(n279),.dout(n289),.clk(gclk));
	jor g204(.dina(w_dff_B_taZEckL56_0),.dinb(n278),.dout(w_dff_A_TGjlIEZu5_2),.clk(gclk));
	jand g205(.dina(w_n153_2[0]),.dinb(w_G91gat_0[1]),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n157_0[0]),.dinb(w_G55gat_0[0]),.dout(n292),.clk(gclk));
	jand g207(.dina(w_n292_1[1]),.dinb(w_G143gat_0[0]),.dout(n293),.clk(gclk));
	jand g208(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n294),.clk(gclk));
	jand g209(.dina(w_n163_0[0]),.dinb(w_G17gat_1[0]),.dout(n295),.clk(gclk));
	jand g210(.dina(w_dff_B_XdB8JRhX9_0),.dinb(w_n162_0[0]),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n296_1[1]),.dinb(w_dff_B_oKw6tXG59_1),.dout(n297),.clk(gclk));
	jor g212(.dina(n297),.dinb(n293),.dout(n298),.clk(gclk));
	jor g213(.dina(n298),.dinb(n291),.dout(n299),.clk(gclk));
	jand g214(.dina(w_n299_1[1]),.dinb(w_G159gat_2[0]),.dout(n300),.clk(gclk));
	jor g215(.dina(w_n299_1[0]),.dinb(w_G159gat_1[2]),.dout(n301),.clk(gclk));
	jand g216(.dina(w_n193_0[2]),.dinb(w_G183gat_1[0]),.dout(n302),.clk(gclk));
	jor g217(.dina(w_n193_0[1]),.dinb(w_G183gat_0[2]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n238_0[0]),.dinb(w_n303_0[1]),.dout(n304),.clk(gclk));
	jor g219(.dina(n304),.dinb(w_n302_0[1]),.dout(n305),.clk(gclk));
	jnot g220(.din(w_G165gat_2[0]),.dout(n306),.clk(gclk));
	jand g221(.dina(w_n153_1[2]),.dinb(w_G96gat_0[1]),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n292_1[0]),.dinb(w_G146gat_0[0]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_lCxEUWz72_0),.dinb(w_n296_1[0]),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(n308),.dout(n311),.clk(gclk));
	jor g226(.dina(n311),.dinb(n307),.dout(n312),.clk(gclk));
	jnot g227(.din(w_n312_1[1]),.dout(n313),.clk(gclk));
	jand g228(.dina(n313),.dinb(w_dff_B_ZsmjwWGx2_1),.dout(n314),.clk(gclk));
	jnot g229(.din(n314),.dout(n315),.clk(gclk));
	jand g230(.dina(w_n153_1[1]),.dinb(w_G101gat_0[1]),.dout(n316),.clk(gclk));
	jand g231(.dina(w_n292_0[2]),.dinb(w_G149gat_0[0]),.dout(n317),.clk(gclk));
	jand g232(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n318),.clk(gclk));
	jor g233(.dina(w_dff_B_2NlrS6577_0),.dinb(w_n296_0[2]),.dout(n319),.clk(gclk));
	jor g234(.dina(n319),.dinb(n317),.dout(n320),.clk(gclk));
	jor g235(.dina(n320),.dinb(n316),.dout(n321),.clk(gclk));
	jor g236(.dina(w_n321_1[1]),.dinb(w_G171gat_2[0]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n153_1[0]),.dinb(w_G106gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_n292_0[1]),.dinb(w_G153gat_0[0]),.dout(n324),.clk(gclk));
	jand g239(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_6AOg5QhU1_0),.dinb(w_n296_0[1]),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g242(.dina(n327),.dinb(n323),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n328_1[1]),.dinb(w_G177gat_2[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n329_0[2]),.dinb(w_n322_0[1]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n330_0[2]),.dinb(w_n315_0[1]),.dout(n331),.clk(gclk));
	jand g246(.dina(w_n331_0[1]),.dinb(w_n305_1[1]),.dout(n332),.clk(gclk));
	jand g247(.dina(w_n312_1[0]),.dinb(w_G165gat_1[2]),.dout(n333),.clk(gclk));
	jand g248(.dina(w_n321_1[0]),.dinb(w_G171gat_1[2]),.dout(n334),.clk(gclk));
	jand g249(.dina(w_n328_1[0]),.dinb(w_G177gat_1[2]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_0[2]),.dinb(w_n322_0[0]),.dout(n336),.clk(gclk));
	jor g251(.dina(n336),.dinb(w_dff_B_FE3FwbSM1_1),.dout(n337),.clk(gclk));
	jand g252(.dina(w_n337_0[2]),.dinb(w_n315_0[0]),.dout(n338),.clk(gclk));
	jor g253(.dina(n338),.dinb(w_dff_B_jLQujL9a6_1),.dout(n339),.clk(gclk));
	jor g254(.dina(w_n339_0[1]),.dinb(n332),.dout(n340),.clk(gclk));
	jand g255(.dina(w_n340_0[1]),.dinb(w_dff_B_TPc0ucj43_1),.dout(n341),.clk(gclk));
	jor g256(.dina(n341),.dinb(w_dff_B_S5Soqeu77_1),.dout(w_dff_A_pjkRVhk99_2),.clk(gclk));
	jnot g257(.din(w_n302_0[0]),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n303_0[0]),.dout(n344),.clk(gclk));
	jor g259(.dina(w_n232_0[0]),.dinb(w_dff_B_GIwfvGCa0_1),.dout(n345),.clk(gclk));
	jand g260(.dina(n345),.dinb(w_dff_B_xNk9LDaO0_1),.dout(n346),.clk(gclk));
	jxor g261(.dina(w_n328_0[2]),.dinb(w_G177gat_1[1]),.dout(n347),.clk(gclk));
	jnot g262(.din(w_n347_0[2]),.dout(n348),.clk(gclk));
	jor g263(.dina(w_dff_B_fbJ5YCMu6_0),.dinb(w_n346_1[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(w_n347_0[1]),.dinb(w_n305_1[0]),.dout(n350),.clk(gclk));
	jand g265(.dina(n350),.dinb(w_G219gat_2[0]),.dout(n351),.clk(gclk));
	jand g266(.dina(n351),.dinb(n349),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n347_0[0]),.dinb(w_G228gat_2[0]),.dout(n353),.clk(gclk));
	jand g268(.dina(w_G237gat_2[0]),.dinb(w_G177gat_1[0]),.dout(n354),.clk(gclk));
	jor g269(.dina(n354),.dinb(w_G246gat_2[0]),.dout(n355),.clk(gclk));
	jand g270(.dina(w_dff_B_nusyD60S3_0),.dinb(w_n328_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n181_2[0]),.dinb(w_G177gat_0[2]),.dout(n357),.clk(gclk));
	jand g272(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n358),.clk(gclk));
	jor g273(.dina(w_dff_B_bDjocvHb4_0),.dinb(n357),.dout(n359),.clk(gclk));
	jor g274(.dina(w_dff_B_mT3mTevV1_0),.dinb(n356),.dout(n360),.clk(gclk));
	jor g275(.dina(n360),.dinb(n353),.dout(n361),.clk(gclk));
	jor g276(.dina(w_dff_B_YdjaX97Q5_0),.dinb(n352),.dout(w_dff_A_cQvl11VV9_2),.clk(gclk));
	jnot g277(.din(w_n331_0[0]),.dout(n363),.clk(gclk));
	jor g278(.dina(w_dff_B_XoYr91NN9_0),.dinb(w_n346_1[0]),.dout(n364),.clk(gclk));
	jnot g279(.din(w_n339_0[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_dff_B_Oj41tBd14_0),.dinb(n364),.dout(n366),.clk(gclk));
	jxor g281(.dina(w_n299_0[2]),.dinb(w_G159gat_1[1]),.dout(n367),.clk(gclk));
	jnot g282(.din(w_n367_0[2]),.dout(n368),.clk(gclk));
	jor g283(.dina(w_dff_B_NgN9tBnN1_0),.dinb(n366),.dout(n369),.clk(gclk));
	jor g284(.dina(w_n367_0[1]),.dinb(w_n340_0[0]),.dout(n370),.clk(gclk));
	jand g285(.dina(n370),.dinb(w_G219gat_1[2]),.dout(n371),.clk(gclk));
	jand g286(.dina(n371),.dinb(n369),.dout(n372),.clk(gclk));
	jand g287(.dina(w_n367_0[0]),.dinb(w_G228gat_1[2]),.dout(n373),.clk(gclk));
	jand g288(.dina(w_G237gat_1[2]),.dinb(w_G159gat_1[0]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_G246gat_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(w_dff_B_FNrHhMWb6_0),.dinb(w_n299_0[1]),.dout(n376),.clk(gclk));
	jand g291(.dina(w_n181_1[2]),.dinb(w_G159gat_0[2]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n378),.clk(gclk));
	jor g293(.dina(w_dff_B_7a9JN6SX4_0),.dinb(n377),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_3nBWanky2_0),.dinb(n376),.dout(n380),.clk(gclk));
	jor g295(.dina(n380),.dinb(n373),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_zEyI8zSt7_0),.dinb(n372),.dout(G878gat),.clk(gclk));
	jxor g297(.dina(w_n312_0[2]),.dinb(w_G165gat_1[1]),.dout(n383),.clk(gclk));
	jnot g298(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n337_0[1]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n330_0[1]),.dout(n386),.clk(gclk));
	jor g301(.dina(w_dff_B_YUvVzvXC8_0),.dinb(w_n346_0[2]),.dout(n387),.clk(gclk));
	jand g302(.dina(n387),.dinb(w_dff_B_7R9s9ooO7_1),.dout(n388),.clk(gclk));
	jor g303(.dina(n388),.dinb(w_dff_B_1pd4Ccwh2_1),.dout(n389),.clk(gclk));
	jand g304(.dina(w_n330_0[0]),.dinb(w_n305_0[2]),.dout(n390),.clk(gclk));
	jor g305(.dina(n390),.dinb(w_n337_0[0]),.dout(n391),.clk(gclk));
	jor g306(.dina(n391),.dinb(w_n383_0[1]),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_G219gat_1[1]),.dout(n393),.clk(gclk));
	jand g308(.dina(n393),.dinb(n389),.dout(n394),.clk(gclk));
	jand g309(.dina(w_n383_0[0]),.dinb(w_G228gat_1[1]),.dout(n395),.clk(gclk));
	jand g310(.dina(w_G237gat_1[1]),.dinb(w_G165gat_1[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(n396),.dinb(w_G246gat_1[1]),.dout(n397),.clk(gclk));
	jand g312(.dina(w_dff_B_jvsOuxFA9_0),.dinb(w_n312_0[1]),.dout(n398),.clk(gclk));
	jand g313(.dina(w_n181_1[1]),.dinb(w_G165gat_0[2]),.dout(n399),.clk(gclk));
	jand g314(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n400),.clk(gclk));
	jor g315(.dina(w_dff_B_ImGLq4gj7_0),.dinb(n399),.dout(n401),.clk(gclk));
	jor g316(.dina(w_dff_B_0DzC5rDp0_0),.dinb(n398),.dout(n402),.clk(gclk));
	jor g317(.dina(n402),.dinb(n395),.dout(n403),.clk(gclk));
	jor g318(.dina(w_dff_B_ObHH3cAX7_0),.dinb(n394),.dout(G879gat),.clk(gclk));
	jxor g319(.dina(w_n321_0[2]),.dinb(w_G171gat_1[1]),.dout(n405),.clk(gclk));
	jnot g320(.din(w_n405_0[2]),.dout(n406),.clk(gclk));
	jnot g321(.din(w_n335_0[1]),.dout(n407),.clk(gclk));
	jnot g322(.din(w_n329_0[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_zhzCgr9l2_0),.dinb(w_n346_0[1]),.dout(n409),.clk(gclk));
	jand g324(.dina(n409),.dinb(w_dff_B_WfuUDdre2_1),.dout(n410),.clk(gclk));
	jor g325(.dina(n410),.dinb(w_dff_B_bRPOcEi75_1),.dout(n411),.clk(gclk));
	jand g326(.dina(w_n329_0[0]),.dinb(w_n305_0[1]),.dout(n412),.clk(gclk));
	jor g327(.dina(n412),.dinb(w_n335_0[0]),.dout(n413),.clk(gclk));
	jor g328(.dina(n413),.dinb(w_n405_0[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_G219gat_1[0]),.dout(n415),.clk(gclk));
	jand g330(.dina(n415),.dinb(n411),.dout(n416),.clk(gclk));
	jand g331(.dina(w_n405_0[0]),.dinb(w_G228gat_1[0]),.dout(n417),.clk(gclk));
	jand g332(.dina(w_G237gat_1[0]),.dinb(w_G171gat_1[0]),.dout(n418),.clk(gclk));
	jor g333(.dina(n418),.dinb(w_G246gat_1[0]),.dout(n419),.clk(gclk));
	jand g334(.dina(w_dff_B_UyJSPswS6_0),.dinb(w_n321_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n181_1[0]),.dinb(w_G171gat_0[2]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(w_dff_B_PMLc6udB4_0),.dinb(n421),.dout(n423),.clk(gclk));
	jor g338(.dina(w_dff_B_7HwCOTBq1_0),.dinb(n420),.dout(n424),.clk(gclk));
	jor g339(.dina(n424),.dinb(n417),.dout(n425),.clk(gclk));
	jor g340(.dina(w_dff_B_Nigc0Z265_0),.dinb(n416),.dout(G880gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_qsl1bnTk2_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_G13gat_0[1]),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_jk2LrdXk9_0),.doutb(w_G17gat_1[1]),.doutc(w_dff_A_Ol41ZdeR4_2),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_G17gat_2[2]),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_G29gat_0[0]),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_SozBqppf7_1),.doutc(w_G42gat_0[2]),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_G42gat_1[0]),.doutb(w_dff_A_Q65ouTAs2_1),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_XqHtVFsO4_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_OxXuaSf93_0),.doutb(w_dff_A_JJjKsZ4p2_1),.doutc(w_G55gat_0[2]),.din(G55gat));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_G68gat_0[1]),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_pFaqW4Nf0_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_QtnwI8EJ5_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_X1OJdXbj3_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_vfPBbFAz9_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_eI78CFqv4_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_Vk9D0hN00_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_DZe664RI1_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_RO9ze0Q51_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_FKKbzkpB8_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl jspl_w_G126gat_0(.douta(w_dff_A_SU8vcFnq8_0),.doutb(w_G126gat_0[1]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_G130gat_0[1]),.din(w_dff_B_cH2q8aK22_2));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_auBPxiDF9_1),.din(w_dff_B_FlFqBa146_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_9OjhhdMe0_1),.din(w_dff_B_0BQ6LSLO5_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_m7f1IMZA8_1),.din(w_dff_B_mmKJ5qqi8_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_x4rl85sv9_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_GboRYmrx5_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_G159gat_0[1]),.doutc(w_dff_A_lL6cgLL13_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_G159gat_1[0]),.doutb(w_dff_A_9OHafTkt0_1),.doutc(w_dff_A_vqEMsjDs5_2),.din(w_G159gat_0[0]));
	jspl jspl_w_G159gat_2(.douta(w_dff_A_Zph5uTU19_0),.doutb(w_G159gat_2[1]),.din(w_G159gat_0[1]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_G165gat_0[1]),.doutc(w_dff_A_jWD1m8Ga0_2),.din(G165gat));
	jspl3 jspl3_w_G165gat_1(.douta(w_G165gat_1[0]),.doutb(w_dff_A_4yaqyCEp6_1),.doutc(w_dff_A_ZrpWIYCz2_2),.din(w_G165gat_0[0]));
	jspl jspl_w_G165gat_2(.douta(w_G165gat_2[0]),.doutb(w_G165gat_2[1]),.din(w_G165gat_0[1]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_dff_A_W5CMpLB79_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_dff_A_y1U3RlEq9_1),.doutc(w_dff_A_OMzKAEPm8_2),.din(w_G171gat_0[0]));
	jspl jspl_w_G171gat_2(.douta(w_dff_A_k6DoSIxV4_0),.doutb(w_G171gat_2[1]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_G177gat_0[1]),.doutc(w_dff_A_08epPKth5_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_jGoQ9h4C1_1),.doutc(w_dff_A_h9WWGJRw2_2),.din(w_G177gat_0[0]));
	jspl jspl_w_G177gat_2(.douta(w_dff_A_oj9M9gvy2_0),.doutb(w_G177gat_2[1]),.din(w_G177gat_0[1]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_yNv5bI6Q9_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_jGGLLWCh5_0),.doutb(w_dff_A_5HyzhKfF7_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl jspl_w_G183gat_2(.douta(w_dff_A_XUvNKZBq2_0),.doutb(w_G183gat_2[1]),.din(w_G183gat_0[1]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_XBC0j54E6_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_galFhZhB6_1),.doutc(w_dff_A_aq6BOP380_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_M4yjlATT5_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_rdzFG80g1_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_YXUvDKir7_1),.doutc(w_dff_A_PvdxKnbG1_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_p7ylLqnr5_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_G201gat_0[1]),.doutc(w_dff_A_WAjYHuCH9_2),.din(G201gat));
	jspl3 jspl3_w_G201gat_1(.douta(w_G201gat_1[0]),.doutb(w_dff_A_RkxdeWDZ7_1),.doutc(w_dff_A_yuUaDZct5_2),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G201gat_2(.douta(w_G201gat_2[0]),.doutb(w_dff_A_8LuQ0HYn9_1),.doutc(w_G201gat_2[2]),.din(w_G201gat_0[1]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_t7KS4ed80_0),.doutb(w_dff_A_lIgj2OvW9_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_nzN8IDbZ5_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_G219gat_1[1]),.doutc(w_G219gat_1[2]),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_B2yRUTx84_0),.doutb(w_G219gat_2[1]),.doutc(w_dff_A_ix8qC5Da8_2),.din(w_G219gat_0[1]));
	jspl jspl_w_G219gat_3(.douta(w_dff_A_hYga5udw7_0),.doutb(w_G219gat_3[1]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_G228gat_0[0]),.doutb(w_G228gat_0[1]),.doutc(w_dff_A_Nhdao0Dr4_2),.din(w_dff_B_T91JKijC2_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_G228gat_2[0]),.doutb(w_dff_A_8BBT3WcH8_1),.doutc(w_dff_A_LGmn9IrG1_2),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_G228gat_3[1]),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_G237gat_0[0]),.doutb(w_G237gat_0[1]),.doutc(w_G237gat_0[2]),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_G237gat_2[0]),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_G237gat_3[1]),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_G246gat_0[0]),.doutb(w_G246gat_0[1]),.doutc(w_G246gat_0[2]),.din(w_dff_B_whdvNOk09_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_G246gat_2[0]),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_G246gat_3[1]),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_VD6wq4HN3_0),.doutb(w_dff_A_iiGZ1f197_1),.doutc(w_G261gat_0[2]),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_jjSD3FkA1_1),.doutc(w_dff_A_CX6SNnSY4_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_G447gat_0[2]),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_wbw40VA04_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n96_0(.douta(w_dff_A_i1fXFduF3_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(w_dff_B_CyKwyphr1_2));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n118_0(.douta(w_dff_A_SA7BZnPm1_0),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n121_0(.douta(w_dff_A_OM48yGBA4_0),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(w_dff_B_Kewu7pk98_2));
	jspl jspl_w_n149_0(.douta(w_dff_A_EsLHXE3L0_0),.doutb(w_n149_0[1]),.din(n149));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_n153_2[2]),.din(w_n153_0[1]));
	jspl jspl_w_n153_3(.douta(w_n153_3[0]),.doutb(w_n153_3[1]),.din(w_n153_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_dff_A_rxtSPeVE2_1),.din(n154));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_KLPTewSx0_1),.doutc(w_dff_A_WXfcxGc05_2),.din(n165));
	jspl3 jspl3_w_n165_1(.douta(w_n165_1[0]),.doutb(w_dff_A_JMRI1rol2_1),.doutc(w_dff_A_ksVZSOd59_2),.din(w_n165_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n181_3(.douta(w_n181_3[0]),.doutb(w_n181_3[1]),.din(w_n181_0[2]));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.doutc(w_n193_0[2]),.din(n193));
	jspl jspl_w_n193_1(.douta(w_n193_1[0]),.doutb(w_n193_1[1]),.din(w_n193_0[0]));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_dff_A_9WwPqc2N7_1),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_dff_A_P9E7V1247_0),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl jspl_w_n217_1(.douta(w_n217_1[0]),.doutb(w_n217_1[1]),.din(w_n217_0[0]));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.doutc(w_n222_0[2]),.din(n222));
	jspl jspl_w_n222_1(.douta(w_n222_1[0]),.doutb(w_n222_1[1]),.din(w_n222_0[0]));
	jspl jspl_w_n223_0(.douta(w_dff_A_6UN2C2Xw2_0),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n224_0(.douta(w_dff_A_ythxWxRF6_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n228_0(.douta(w_dff_A_gvbS2i9b2_0),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_dff_A_rPv8zhsi0_0),.doutb(w_n230_0[1]),.din(n230));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_n238_0[1]),.din(n238));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_wDsjkRMa9_1),.doutc(w_n252_0[2]),.din(n252));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_dff_A_gIRiRx1j2_1),.doutc(w_n273_0[2]),.din(n273));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.doutc(w_n296_0[2]),.din(n296));
	jspl jspl_w_n296_1(.douta(w_n296_1[0]),.doutb(w_n296_1[1]),.din(w_n296_0[0]));
	jspl3 jspl3_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.doutc(w_n299_0[2]),.din(n299));
	jspl jspl_w_n299_1(.douta(w_n299_1[0]),.doutb(w_n299_1[1]),.din(w_n299_0[0]));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_dff_A_GyEHmUoP2_1),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_JO6lxcXS8_1),.din(n303));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl jspl_w_n305_1(.douta(w_n305_1[0]),.doutb(w_n305_1[1]),.din(w_n305_0[0]));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl3 jspl3_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.doutc(w_n321_0[2]),.din(n321));
	jspl jspl_w_n321_1(.douta(w_n321_1[0]),.doutb(w_n321_1[1]),.din(w_n321_0[0]));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n328_1(.douta(w_n328_1[0]),.doutb(w_n328_1[1]),.din(w_n328_0[0]));
	jspl3 jspl3_w_n329_0(.douta(w_dff_A_sEYTIeD96_0),.doutb(w_n329_0[1]),.doutc(w_n329_0[2]),.din(n329));
	jspl3 jspl3_w_n330_0(.douta(w_dff_A_cIMVAcIE0_0),.doutb(w_n330_0[1]),.doutc(w_dff_A_YIhTZkIK0_2),.din(n330));
	jspl jspl_w_n331_0(.douta(w_n331_0[0]),.doutb(w_dff_A_wH5Gg4sN4_1),.din(n331));
	jspl3 jspl3_w_n335_0(.douta(w_dff_A_rvGRHzXk8_0),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n337_0(.douta(w_dff_A_NjUnijN24_0),.doutb(w_n337_0[1]),.doutc(w_n337_0[2]),.din(n337));
	jspl jspl_w_n339_0(.douta(w_n339_0[0]),.doutb(w_dff_A_16O2qm1c0_1),.din(n339));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n347_0(.douta(w_n347_0[0]),.doutb(w_dff_A_Bw1e8Sbi0_1),.doutc(w_n347_0[2]),.din(n347));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_dff_A_I9eTOsSs8_1),.doutc(w_n367_0[2]),.din(n367));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_hma2NagD0_1),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_dff_A_HARwFZmJ1_1),.doutc(w_n405_0[2]),.din(n405));
	jdff dff_B_CyKwyphr1_2(.din(n101),.dout(w_dff_B_CyKwyphr1_2),.clk(gclk));
	jdff dff_B_iugJthxE1_1(.din(n109),.dout(w_dff_B_iugJthxE1_1),.clk(gclk));
	jdff dff_B_tDtNnlHu9_1(.din(G90gat),.dout(w_dff_B_tDtNnlHu9_1),.clk(gclk));
	jdff dff_A_jjSD3FkA1_1(.dout(w_G390gat_0[1]),.din(w_dff_A_jjSD3FkA1_1),.clk(gclk));
	jdff dff_B_2w2NwKet5_0(.din(n119),.dout(w_dff_B_2w2NwKet5_0),.clk(gclk));
	jdff dff_B_GdgUF8cQ0_1(.din(G74gat),.dout(w_dff_B_GdgUF8cQ0_1),.clk(gclk));
	jdff dff_B_WLWUl7eF7_1(.din(G89gat),.dout(w_dff_B_WLWUl7eF7_1),.clk(gclk));
	jdff dff_B_xwH9UetB0_0(.din(n131),.dout(w_dff_B_xwH9UetB0_0),.clk(gclk));
	jdff dff_B_bU6U96DH3_1(.din(G135gat),.dout(w_dff_B_bU6U96DH3_1),.clk(gclk));
	jdff dff_B_ESnsRQaR5_0(.din(n127),.dout(w_dff_B_ESnsRQaR5_0),.clk(gclk));
	jdff dff_B_8vDVZbqX9_0(.din(n140),.dout(w_dff_B_8vDVZbqX9_0),.clk(gclk));
	jdff dff_B_4fXyhJE60_1(.din(G207gat),.dout(w_dff_B_4fXyhJE60_1),.clk(gclk));
	jdff dff_B_PNiG9O2k8_0(.din(n136),.dout(w_dff_B_PNiG9O2k8_0),.clk(gclk));
	jdff dff_B_cH2q8aK22_2(.din(G130gat),.dout(w_dff_B_cH2q8aK22_2),.clk(gclk));
	jdff dff_B_6PGRgfmA5_0(.din(n188),.dout(w_dff_B_6PGRgfmA5_0),.clk(gclk));
	jdff dff_B_Rj7S9AwS4_0(.din(n186),.dout(w_dff_B_Rj7S9AwS4_0),.clk(gclk));
	jdff dff_B_5PkVdPCL5_0(.din(w_dff_B_Rj7S9AwS4_0),.dout(w_dff_B_5PkVdPCL5_0),.clk(gclk));
	jdff dff_B_mzqr1oNS7_0(.din(w_dff_B_5PkVdPCL5_0),.dout(w_dff_B_mzqr1oNS7_0),.clk(gclk));
	jdff dff_B_GA4BDbyK5_0(.din(n185),.dout(w_dff_B_GA4BDbyK5_0),.clk(gclk));
	jdff dff_B_UNalbLpO1_0(.din(w_dff_B_GA4BDbyK5_0),.dout(w_dff_B_UNalbLpO1_0),.clk(gclk));
	jdff dff_B_auSpZ2Q82_0(.din(w_dff_B_UNalbLpO1_0),.dout(w_dff_B_auSpZ2Q82_0),.clk(gclk));
	jdff dff_B_G2xuKXNM6_0(.din(n176),.dout(w_dff_B_G2xuKXNM6_0),.clk(gclk));
	jdff dff_B_ircdiJlw5_0(.din(w_dff_B_G2xuKXNM6_0),.dout(w_dff_B_ircdiJlw5_0),.clk(gclk));
	jdff dff_B_DdFX4hTk6_0(.din(w_dff_B_ircdiJlw5_0),.dout(w_dff_B_DdFX4hTk6_0),.clk(gclk));
	jdff dff_B_XUZUtypu5_0(.din(w_dff_B_DdFX4hTk6_0),.dout(w_dff_B_XUZUtypu5_0),.clk(gclk));
	jdff dff_B_hORW2yly9_0(.din(w_dff_B_XUZUtypu5_0),.dout(w_dff_B_hORW2yly9_0),.clk(gclk));
	jdff dff_B_LAkMJVPZ7_0(.din(w_dff_B_hORW2yly9_0),.dout(w_dff_B_LAkMJVPZ7_0),.clk(gclk));
	jdff dff_A_DJcKU5pm5_1(.dout(w_G201gat_2[1]),.din(w_dff_A_DJcKU5pm5_1),.clk(gclk));
	jdff dff_A_76OVWLZU0_1(.dout(w_dff_A_DJcKU5pm5_1),.din(w_dff_A_76OVWLZU0_1),.clk(gclk));
	jdff dff_A_drbIm2M96_1(.dout(w_dff_A_76OVWLZU0_1),.din(w_dff_A_drbIm2M96_1),.clk(gclk));
	jdff dff_A_Va0bTc9T9_1(.dout(w_dff_A_drbIm2M96_1),.din(w_dff_A_Va0bTc9T9_1),.clk(gclk));
	jdff dff_A_dM5i8yYs9_1(.dout(w_dff_A_Va0bTc9T9_1),.din(w_dff_A_dM5i8yYs9_1),.clk(gclk));
	jdff dff_A_Fqq71yoJ7_1(.dout(w_dff_A_dM5i8yYs9_1),.din(w_dff_A_Fqq71yoJ7_1),.clk(gclk));
	jdff dff_A_gMwGrmXA5_1(.dout(w_dff_A_Fqq71yoJ7_1),.din(w_dff_A_gMwGrmXA5_1),.clk(gclk));
	jdff dff_A_8LuQ0HYn9_1(.dout(w_dff_A_gMwGrmXA5_1),.din(w_dff_A_8LuQ0HYn9_1),.clk(gclk));
	jdff dff_B_n3B4a7lS8_0(.din(n250),.dout(w_dff_B_n3B4a7lS8_0),.clk(gclk));
	jdff dff_B_1LaZuo0X7_0(.din(w_dff_B_n3B4a7lS8_0),.dout(w_dff_B_1LaZuo0X7_0),.clk(gclk));
	jdff dff_B_vEOIMitj1_0(.din(w_dff_B_1LaZuo0X7_0),.dout(w_dff_B_vEOIMitj1_0),.clk(gclk));
	jdff dff_B_RFRaNVNs6_0(.din(w_dff_B_vEOIMitj1_0),.dout(w_dff_B_RFRaNVNs6_0),.clk(gclk));
	jdff dff_B_tMPfvelr4_0(.din(w_dff_B_RFRaNVNs6_0),.dout(w_dff_B_tMPfvelr4_0),.clk(gclk));
	jdff dff_B_O3NwFjze2_0(.din(n248),.dout(w_dff_B_O3NwFjze2_0),.clk(gclk));
	jdff dff_B_nkSNQtUL6_0(.din(w_dff_B_O3NwFjze2_0),.dout(w_dff_B_nkSNQtUL6_0),.clk(gclk));
	jdff dff_B_ZTIf6Wlo2_0(.din(w_dff_B_nkSNQtUL6_0),.dout(w_dff_B_ZTIf6Wlo2_0),.clk(gclk));
	jdff dff_B_2a9wlo0A4_0(.din(n247),.dout(w_dff_B_2a9wlo0A4_0),.clk(gclk));
	jdff dff_B_RPP6nf8I6_0(.din(w_dff_B_2a9wlo0A4_0),.dout(w_dff_B_RPP6nf8I6_0),.clk(gclk));
	jdff dff_B_v7bZx6Pu4_0(.din(w_dff_B_RPP6nf8I6_0),.dout(w_dff_B_v7bZx6Pu4_0),.clk(gclk));
	jdff dff_B_FPQEmp059_0(.din(w_dff_B_v7bZx6Pu4_0),.dout(w_dff_B_FPQEmp059_0),.clk(gclk));
	jdff dff_B_LJog64C59_0(.din(n244),.dout(w_dff_B_LJog64C59_0),.clk(gclk));
	jdff dff_B_AqlrS1L85_0(.din(w_dff_B_LJog64C59_0),.dout(w_dff_B_AqlrS1L85_0),.clk(gclk));
	jdff dff_B_0Q2cIPyv4_0(.din(w_dff_B_AqlrS1L85_0),.dout(w_dff_B_0Q2cIPyv4_0),.clk(gclk));
	jdff dff_B_IthI9RXJ2_0(.din(w_dff_B_0Q2cIPyv4_0),.dout(w_dff_B_IthI9RXJ2_0),.clk(gclk));
	jdff dff_B_4CEbYnw38_0(.din(w_dff_B_IthI9RXJ2_0),.dout(w_dff_B_4CEbYnw38_0),.clk(gclk));
	jdff dff_B_jzXK16sE8_0(.din(w_dff_B_4CEbYnw38_0),.dout(w_dff_B_jzXK16sE8_0),.clk(gclk));
	jdff dff_A_Ucd6nBB01_0(.dout(w_G219gat_3[0]),.din(w_dff_A_Ucd6nBB01_0),.clk(gclk));
	jdff dff_A_iyftkq4J4_0(.dout(w_dff_A_Ucd6nBB01_0),.din(w_dff_A_iyftkq4J4_0),.clk(gclk));
	jdff dff_A_r3WWknnc7_0(.dout(w_dff_A_iyftkq4J4_0),.din(w_dff_A_r3WWknnc7_0),.clk(gclk));
	jdff dff_A_hYga5udw7_0(.dout(w_dff_A_r3WWknnc7_0),.din(w_dff_A_hYga5udw7_0),.clk(gclk));
	jdff dff_B_YE4IuKer1_1(.din(n195),.dout(w_dff_B_YE4IuKer1_1),.clk(gclk));
	jdff dff_B_vwZ6j0gl8_1(.din(w_dff_B_YE4IuKer1_1),.dout(w_dff_B_vwZ6j0gl8_1),.clk(gclk));
	jdff dff_B_ezsaci3V1_1(.din(w_dff_B_vwZ6j0gl8_1),.dout(w_dff_B_ezsaci3V1_1),.clk(gclk));
	jdff dff_B_FmOh0vb39_1(.din(w_dff_B_ezsaci3V1_1),.dout(w_dff_B_FmOh0vb39_1),.clk(gclk));
	jdff dff_A_Ku7EBwKj6_1(.dout(w_n194_0[1]),.din(w_dff_A_Ku7EBwKj6_1),.clk(gclk));
	jdff dff_A_74RdxEXT9_1(.dout(w_dff_A_Ku7EBwKj6_1),.din(w_dff_A_74RdxEXT9_1),.clk(gclk));
	jdff dff_A_ju7K1gXA5_1(.dout(w_dff_A_74RdxEXT9_1),.din(w_dff_A_ju7K1gXA5_1),.clk(gclk));
	jdff dff_A_9WwPqc2N7_1(.dout(w_dff_A_ju7K1gXA5_1),.din(w_dff_A_9WwPqc2N7_1),.clk(gclk));
	jdff dff_A_GOqi5TUC6_0(.dout(w_G183gat_2[0]),.din(w_dff_A_GOqi5TUC6_0),.clk(gclk));
	jdff dff_A_LT5vWtVn3_0(.dout(w_dff_A_GOqi5TUC6_0),.din(w_dff_A_LT5vWtVn3_0),.clk(gclk));
	jdff dff_A_U74bqfG07_0(.dout(w_dff_A_LT5vWtVn3_0),.din(w_dff_A_U74bqfG07_0),.clk(gclk));
	jdff dff_A_yFkepAiF0_0(.dout(w_dff_A_U74bqfG07_0),.din(w_dff_A_yFkepAiF0_0),.clk(gclk));
	jdff dff_A_i3TYDPGR4_0(.dout(w_dff_A_yFkepAiF0_0),.din(w_dff_A_i3TYDPGR4_0),.clk(gclk));
	jdff dff_A_64gn8B5s4_0(.dout(w_dff_A_i3TYDPGR4_0),.din(w_dff_A_64gn8B5s4_0),.clk(gclk));
	jdff dff_A_JVbeLkoD2_0(.dout(w_dff_A_64gn8B5s4_0),.din(w_dff_A_JVbeLkoD2_0),.clk(gclk));
	jdff dff_A_XUvNKZBq2_0(.dout(w_dff_A_JVbeLkoD2_0),.din(w_dff_A_XUvNKZBq2_0),.clk(gclk));
	jdff dff_B_gXBZupkW3_0(.din(n271),.dout(w_dff_B_gXBZupkW3_0),.clk(gclk));
	jdff dff_B_hKoZQoUf9_0(.din(w_dff_B_gXBZupkW3_0),.dout(w_dff_B_hKoZQoUf9_0),.clk(gclk));
	jdff dff_B_Z32LhIcC5_0(.din(w_dff_B_hKoZQoUf9_0),.dout(w_dff_B_Z32LhIcC5_0),.clk(gclk));
	jdff dff_B_N27f2amn7_0(.din(w_dff_B_Z32LhIcC5_0),.dout(w_dff_B_N27f2amn7_0),.clk(gclk));
	jdff dff_B_sot1kt8j9_0(.din(w_dff_B_N27f2amn7_0),.dout(w_dff_B_sot1kt8j9_0),.clk(gclk));
	jdff dff_B_gRK9DI3U2_0(.din(n269),.dout(w_dff_B_gRK9DI3U2_0),.clk(gclk));
	jdff dff_B_DIj5wJvP7_0(.din(w_dff_B_gRK9DI3U2_0),.dout(w_dff_B_DIj5wJvP7_0),.clk(gclk));
	jdff dff_B_xrA1lCIC7_0(.din(w_dff_B_DIj5wJvP7_0),.dout(w_dff_B_xrA1lCIC7_0),.clk(gclk));
	jdff dff_B_sj7NpmzF7_0(.din(n268),.dout(w_dff_B_sj7NpmzF7_0),.clk(gclk));
	jdff dff_B_usRYsrWj5_0(.din(w_dff_B_sj7NpmzF7_0),.dout(w_dff_B_usRYsrWj5_0),.clk(gclk));
	jdff dff_B_gQ6iSmGV4_0(.din(w_dff_B_usRYsrWj5_0),.dout(w_dff_B_gQ6iSmGV4_0),.clk(gclk));
	jdff dff_B_qJEnLQRc6_0(.din(n263),.dout(w_dff_B_qJEnLQRc6_0),.clk(gclk));
	jdff dff_B_O6om52v94_0(.din(w_dff_B_qJEnLQRc6_0),.dout(w_dff_B_O6om52v94_0),.clk(gclk));
	jdff dff_B_kSfSpbUW3_0(.din(w_dff_B_O6om52v94_0),.dout(w_dff_B_kSfSpbUW3_0),.clk(gclk));
	jdff dff_B_wNHw4sdd2_0(.din(w_dff_B_kSfSpbUW3_0),.dout(w_dff_B_wNHw4sdd2_0),.clk(gclk));
	jdff dff_B_NXeFrPuv1_0(.din(w_dff_B_wNHw4sdd2_0),.dout(w_dff_B_NXeFrPuv1_0),.clk(gclk));
	jdff dff_B_wyNBG4UK4_0(.din(w_dff_B_NXeFrPuv1_0),.dout(w_dff_B_wyNBG4UK4_0),.clk(gclk));
	jdff dff_B_pvGs5Tpn8_1(.din(n253),.dout(w_dff_B_pvGs5Tpn8_1),.clk(gclk));
	jdff dff_B_0Sr4TRom6_1(.din(w_dff_B_pvGs5Tpn8_1),.dout(w_dff_B_0Sr4TRom6_1),.clk(gclk));
	jdff dff_B_I9xaJ2Vs3_1(.din(w_dff_B_0Sr4TRom6_1),.dout(w_dff_B_I9xaJ2Vs3_1),.clk(gclk));
	jdff dff_B_7RiwbCrg6_1(.din(w_dff_B_I9xaJ2Vs3_1),.dout(w_dff_B_7RiwbCrg6_1),.clk(gclk));
	jdff dff_A_MBRSfp1H7_1(.dout(w_n252_0[1]),.din(w_dff_A_MBRSfp1H7_1),.clk(gclk));
	jdff dff_A_ZNgEiuxT4_1(.dout(w_dff_A_MBRSfp1H7_1),.din(w_dff_A_ZNgEiuxT4_1),.clk(gclk));
	jdff dff_A_c2K6wtFV0_1(.dout(w_dff_A_ZNgEiuxT4_1),.din(w_dff_A_c2K6wtFV0_1),.clk(gclk));
	jdff dff_A_wDsjkRMa9_1(.dout(w_dff_A_c2K6wtFV0_1),.din(w_dff_A_wDsjkRMa9_1),.clk(gclk));
	jdff dff_B_ilJVTnfp2_0(.din(n289),.dout(w_dff_B_ilJVTnfp2_0),.clk(gclk));
	jdff dff_B_hqe7xUh36_0(.din(w_dff_B_ilJVTnfp2_0),.dout(w_dff_B_hqe7xUh36_0),.clk(gclk));
	jdff dff_B_taZEckL56_0(.din(w_dff_B_hqe7xUh36_0),.dout(w_dff_B_taZEckL56_0),.clk(gclk));
	jdff dff_B_rwO8bQQN1_0(.din(n287),.dout(w_dff_B_rwO8bQQN1_0),.clk(gclk));
	jdff dff_B_jlcST0ad6_0(.din(w_dff_B_rwO8bQQN1_0),.dout(w_dff_B_jlcST0ad6_0),.clk(gclk));
	jdff dff_B_nmyHmH251_0(.din(w_dff_B_jlcST0ad6_0),.dout(w_dff_B_nmyHmH251_0),.clk(gclk));
	jdff dff_B_bF6rdf6s2_0(.din(n286),.dout(w_dff_B_bF6rdf6s2_0),.clk(gclk));
	jdff dff_B_Y6OtWTIO5_0(.din(w_dff_B_bF6rdf6s2_0),.dout(w_dff_B_Y6OtWTIO5_0),.clk(gclk));
	jdff dff_B_EkS5AOkG9_0(.din(w_dff_B_Y6OtWTIO5_0),.dout(w_dff_B_EkS5AOkG9_0),.clk(gclk));
	jdff dff_B_7KNDYjcd5_0(.din(n281),.dout(w_dff_B_7KNDYjcd5_0),.clk(gclk));
	jdff dff_B_f27Rd26J6_0(.din(w_dff_B_7KNDYjcd5_0),.dout(w_dff_B_f27Rd26J6_0),.clk(gclk));
	jdff dff_B_RSLK5cRb2_0(.din(w_dff_B_f27Rd26J6_0),.dout(w_dff_B_RSLK5cRb2_0),.clk(gclk));
	jdff dff_B_WTCjI5Ai7_0(.din(w_dff_B_RSLK5cRb2_0),.dout(w_dff_B_WTCjI5Ai7_0),.clk(gclk));
	jdff dff_B_G9BcWP8M4_0(.din(w_dff_B_WTCjI5Ai7_0),.dout(w_dff_B_G9BcWP8M4_0),.clk(gclk));
	jdff dff_B_VSJf4baY0_0(.din(w_dff_B_G9BcWP8M4_0),.dout(w_dff_B_VSJf4baY0_0),.clk(gclk));
	jdff dff_B_Njkvh2yk1_0(.din(n274),.dout(w_dff_B_Njkvh2yk1_0),.clk(gclk));
	jdff dff_B_5J4qcP2F2_0(.din(w_dff_B_Njkvh2yk1_0),.dout(w_dff_B_5J4qcP2F2_0),.clk(gclk));
	jdff dff_A_AneMG0E56_1(.dout(w_n273_0[1]),.din(w_dff_A_AneMG0E56_1),.clk(gclk));
	jdff dff_A_gIRiRx1j2_1(.dout(w_dff_A_AneMG0E56_1),.din(w_dff_A_gIRiRx1j2_1),.clk(gclk));
	jdff dff_B_c6VKpkoU6_1(.din(n300),.dout(w_dff_B_c6VKpkoU6_1),.clk(gclk));
	jdff dff_B_vFuiJCzA9_1(.din(w_dff_B_c6VKpkoU6_1),.dout(w_dff_B_vFuiJCzA9_1),.clk(gclk));
	jdff dff_B_wI1HhxIi1_1(.din(w_dff_B_vFuiJCzA9_1),.dout(w_dff_B_wI1HhxIi1_1),.clk(gclk));
	jdff dff_B_r5HwmhLs8_1(.din(w_dff_B_wI1HhxIi1_1),.dout(w_dff_B_r5HwmhLs8_1),.clk(gclk));
	jdff dff_B_pLQsUUeC0_1(.din(w_dff_B_r5HwmhLs8_1),.dout(w_dff_B_pLQsUUeC0_1),.clk(gclk));
	jdff dff_B_OtGd4gEO3_1(.din(w_dff_B_pLQsUUeC0_1),.dout(w_dff_B_OtGd4gEO3_1),.clk(gclk));
	jdff dff_B_uXvqC6gh2_1(.din(w_dff_B_OtGd4gEO3_1),.dout(w_dff_B_uXvqC6gh2_1),.clk(gclk));
	jdff dff_B_joR9MMqD7_1(.din(w_dff_B_uXvqC6gh2_1),.dout(w_dff_B_joR9MMqD7_1),.clk(gclk));
	jdff dff_B_Aa0b0IwG6_1(.din(w_dff_B_joR9MMqD7_1),.dout(w_dff_B_Aa0b0IwG6_1),.clk(gclk));
	jdff dff_B_S5Soqeu77_1(.din(w_dff_B_Aa0b0IwG6_1),.dout(w_dff_B_S5Soqeu77_1),.clk(gclk));
	jdff dff_B_WAM8w3rF1_1(.din(n301),.dout(w_dff_B_WAM8w3rF1_1),.clk(gclk));
	jdff dff_B_cx6ixeKO8_1(.din(w_dff_B_WAM8w3rF1_1),.dout(w_dff_B_cx6ixeKO8_1),.clk(gclk));
	jdff dff_B_EapkadzS9_1(.din(w_dff_B_cx6ixeKO8_1),.dout(w_dff_B_EapkadzS9_1),.clk(gclk));
	jdff dff_B_7Bv86fkV0_1(.din(w_dff_B_EapkadzS9_1),.dout(w_dff_B_7Bv86fkV0_1),.clk(gclk));
	jdff dff_B_vQVTNHeQ5_1(.din(w_dff_B_7Bv86fkV0_1),.dout(w_dff_B_vQVTNHeQ5_1),.clk(gclk));
	jdff dff_B_LvU4dEk43_1(.din(w_dff_B_vQVTNHeQ5_1),.dout(w_dff_B_LvU4dEk43_1),.clk(gclk));
	jdff dff_B_SftK35936_1(.din(w_dff_B_LvU4dEk43_1),.dout(w_dff_B_SftK35936_1),.clk(gclk));
	jdff dff_B_BJUthwO50_1(.din(w_dff_B_SftK35936_1),.dout(w_dff_B_BJUthwO50_1),.clk(gclk));
	jdff dff_B_TPc0ucj43_1(.din(w_dff_B_BJUthwO50_1),.dout(w_dff_B_TPc0ucj43_1),.clk(gclk));
	jdff dff_A_h16rlwVR8_0(.dout(w_G159gat_2[0]),.din(w_dff_A_h16rlwVR8_0),.clk(gclk));
	jdff dff_A_XXvf1WCp3_0(.dout(w_dff_A_h16rlwVR8_0),.din(w_dff_A_XXvf1WCp3_0),.clk(gclk));
	jdff dff_A_qolJqMAb1_0(.dout(w_dff_A_XXvf1WCp3_0),.din(w_dff_A_qolJqMAb1_0),.clk(gclk));
	jdff dff_A_WWX9KilH4_0(.dout(w_dff_A_qolJqMAb1_0),.din(w_dff_A_WWX9KilH4_0),.clk(gclk));
	jdff dff_A_bnoQoq9v7_0(.dout(w_dff_A_WWX9KilH4_0),.din(w_dff_A_bnoQoq9v7_0),.clk(gclk));
	jdff dff_A_5gsQMc7H6_0(.dout(w_dff_A_bnoQoq9v7_0),.din(w_dff_A_5gsQMc7H6_0),.clk(gclk));
	jdff dff_A_Zph5uTU19_0(.dout(w_dff_A_5gsQMc7H6_0),.din(w_dff_A_Zph5uTU19_0),.clk(gclk));
	jdff dff_B_IXoUkkfG5_0(.din(n361),.dout(w_dff_B_IXoUkkfG5_0),.clk(gclk));
	jdff dff_B_QdShgpTW3_0(.din(w_dff_B_IXoUkkfG5_0),.dout(w_dff_B_QdShgpTW3_0),.clk(gclk));
	jdff dff_B_TpwtzfxI7_0(.din(w_dff_B_QdShgpTW3_0),.dout(w_dff_B_TpwtzfxI7_0),.clk(gclk));
	jdff dff_B_T0q9xtsL5_0(.din(w_dff_B_TpwtzfxI7_0),.dout(w_dff_B_T0q9xtsL5_0),.clk(gclk));
	jdff dff_B_oCAS8xxo5_0(.din(w_dff_B_T0q9xtsL5_0),.dout(w_dff_B_oCAS8xxo5_0),.clk(gclk));
	jdff dff_B_PG58jnzw4_0(.din(w_dff_B_oCAS8xxo5_0),.dout(w_dff_B_PG58jnzw4_0),.clk(gclk));
	jdff dff_B_Ys9LyCPv1_0(.din(w_dff_B_PG58jnzw4_0),.dout(w_dff_B_Ys9LyCPv1_0),.clk(gclk));
	jdff dff_B_YdjaX97Q5_0(.din(w_dff_B_Ys9LyCPv1_0),.dout(w_dff_B_YdjaX97Q5_0),.clk(gclk));
	jdff dff_B_aR1sYrKA9_0(.din(n359),.dout(w_dff_B_aR1sYrKA9_0),.clk(gclk));
	jdff dff_B_mT3mTevV1_0(.din(w_dff_B_aR1sYrKA9_0),.dout(w_dff_B_mT3mTevV1_0),.clk(gclk));
	jdff dff_B_aaZdzcYZ6_0(.din(n358),.dout(w_dff_B_aaZdzcYZ6_0),.clk(gclk));
	jdff dff_B_dVkW5Q0U2_0(.din(w_dff_B_aaZdzcYZ6_0),.dout(w_dff_B_dVkW5Q0U2_0),.clk(gclk));
	jdff dff_B_BrptghCx9_0(.din(w_dff_B_dVkW5Q0U2_0),.dout(w_dff_B_BrptghCx9_0),.clk(gclk));
	jdff dff_B_bDjocvHb4_0(.din(w_dff_B_BrptghCx9_0),.dout(w_dff_B_bDjocvHb4_0),.clk(gclk));
	jdff dff_B_swn9wA5a8_0(.din(n355),.dout(w_dff_B_swn9wA5a8_0),.clk(gclk));
	jdff dff_B_8luZ1cp45_0(.din(w_dff_B_swn9wA5a8_0),.dout(w_dff_B_8luZ1cp45_0),.clk(gclk));
	jdff dff_B_Ie2yRgld1_0(.din(w_dff_B_8luZ1cp45_0),.dout(w_dff_B_Ie2yRgld1_0),.clk(gclk));
	jdff dff_B_RTMFee0S6_0(.din(w_dff_B_Ie2yRgld1_0),.dout(w_dff_B_RTMFee0S6_0),.clk(gclk));
	jdff dff_B_nusyD60S3_0(.din(w_dff_B_RTMFee0S6_0),.dout(w_dff_B_nusyD60S3_0),.clk(gclk));
	jdff dff_A_8BBT3WcH8_1(.dout(w_G228gat_2[1]),.din(w_dff_A_8BBT3WcH8_1),.clk(gclk));
	jdff dff_A_LGmn9IrG1_2(.dout(w_G228gat_2[2]),.din(w_dff_A_LGmn9IrG1_2),.clk(gclk));
	jdff dff_A_eb2a4rMR8_0(.dout(w_G219gat_2[0]),.din(w_dff_A_eb2a4rMR8_0),.clk(gclk));
	jdff dff_A_CgLMGN279_0(.dout(w_dff_A_eb2a4rMR8_0),.din(w_dff_A_CgLMGN279_0),.clk(gclk));
	jdff dff_A_hesCPpLD5_0(.dout(w_dff_A_CgLMGN279_0),.din(w_dff_A_hesCPpLD5_0),.clk(gclk));
	jdff dff_A_B2yRUTx84_0(.dout(w_dff_A_hesCPpLD5_0),.din(w_dff_A_B2yRUTx84_0),.clk(gclk));
	jdff dff_A_UVL9DDTW0_2(.dout(w_G219gat_2[2]),.din(w_dff_A_UVL9DDTW0_2),.clk(gclk));
	jdff dff_A_ix8qC5Da8_2(.dout(w_dff_A_UVL9DDTW0_2),.din(w_dff_A_ix8qC5Da8_2),.clk(gclk));
	jdff dff_B_v9e0R0VX8_0(.din(n348),.dout(w_dff_B_v9e0R0VX8_0),.clk(gclk));
	jdff dff_B_sSEyuvey6_0(.din(w_dff_B_v9e0R0VX8_0),.dout(w_dff_B_sSEyuvey6_0),.clk(gclk));
	jdff dff_B_qZaEHHNq0_0(.din(w_dff_B_sSEyuvey6_0),.dout(w_dff_B_qZaEHHNq0_0),.clk(gclk));
	jdff dff_B_XZetI1kQ9_0(.din(w_dff_B_qZaEHHNq0_0),.dout(w_dff_B_XZetI1kQ9_0),.clk(gclk));
	jdff dff_B_vlfLJufO0_0(.din(w_dff_B_XZetI1kQ9_0),.dout(w_dff_B_vlfLJufO0_0),.clk(gclk));
	jdff dff_B_3Di8qKXO4_0(.din(w_dff_B_vlfLJufO0_0),.dout(w_dff_B_3Di8qKXO4_0),.clk(gclk));
	jdff dff_B_fbJ5YCMu6_0(.din(w_dff_B_3Di8qKXO4_0),.dout(w_dff_B_fbJ5YCMu6_0),.clk(gclk));
	jdff dff_A_lWudaLyD8_1(.dout(w_n347_0[1]),.din(w_dff_A_lWudaLyD8_1),.clk(gclk));
	jdff dff_A_3sWm1OLd7_1(.dout(w_dff_A_lWudaLyD8_1),.din(w_dff_A_3sWm1OLd7_1),.clk(gclk));
	jdff dff_A_LuSFRLYE3_1(.dout(w_dff_A_3sWm1OLd7_1),.din(w_dff_A_LuSFRLYE3_1),.clk(gclk));
	jdff dff_A_8RUE70Lh5_1(.dout(w_dff_A_LuSFRLYE3_1),.din(w_dff_A_8RUE70Lh5_1),.clk(gclk));
	jdff dff_A_zs2itGKQ5_1(.dout(w_dff_A_8RUE70Lh5_1),.din(w_dff_A_zs2itGKQ5_1),.clk(gclk));
	jdff dff_A_BgCQorEw5_1(.dout(w_dff_A_zs2itGKQ5_1),.din(w_dff_A_BgCQorEw5_1),.clk(gclk));
	jdff dff_A_Bw1e8Sbi0_1(.dout(w_dff_A_BgCQorEw5_1),.din(w_dff_A_Bw1e8Sbi0_1),.clk(gclk));
	jdff dff_B_KRRdZg4H6_0(.din(n381),.dout(w_dff_B_KRRdZg4H6_0),.clk(gclk));
	jdff dff_B_l9GxMlbw1_0(.din(w_dff_B_KRRdZg4H6_0),.dout(w_dff_B_l9GxMlbw1_0),.clk(gclk));
	jdff dff_B_MIs4jiPP3_0(.din(w_dff_B_l9GxMlbw1_0),.dout(w_dff_B_MIs4jiPP3_0),.clk(gclk));
	jdff dff_B_Wtgiavdv5_0(.din(w_dff_B_MIs4jiPP3_0),.dout(w_dff_B_Wtgiavdv5_0),.clk(gclk));
	jdff dff_B_z0l5yEZX2_0(.din(w_dff_B_Wtgiavdv5_0),.dout(w_dff_B_z0l5yEZX2_0),.clk(gclk));
	jdff dff_B_ImFGVWlM8_0(.din(w_dff_B_z0l5yEZX2_0),.dout(w_dff_B_ImFGVWlM8_0),.clk(gclk));
	jdff dff_B_3Bbl0ugy4_0(.din(w_dff_B_ImFGVWlM8_0),.dout(w_dff_B_3Bbl0ugy4_0),.clk(gclk));
	jdff dff_B_RHfbd8kW2_0(.din(w_dff_B_3Bbl0ugy4_0),.dout(w_dff_B_RHfbd8kW2_0),.clk(gclk));
	jdff dff_B_pD1CfkvY9_0(.din(w_dff_B_RHfbd8kW2_0),.dout(w_dff_B_pD1CfkvY9_0),.clk(gclk));
	jdff dff_B_zEyI8zSt7_0(.din(w_dff_B_pD1CfkvY9_0),.dout(w_dff_B_zEyI8zSt7_0),.clk(gclk));
	jdff dff_B_P0wL9Awp2_0(.din(n379),.dout(w_dff_B_P0wL9Awp2_0),.clk(gclk));
	jdff dff_B_3nBWanky2_0(.din(w_dff_B_P0wL9Awp2_0),.dout(w_dff_B_3nBWanky2_0),.clk(gclk));
	jdff dff_B_nq3fvDGS9_0(.din(n378),.dout(w_dff_B_nq3fvDGS9_0),.clk(gclk));
	jdff dff_B_fHAgzPVK0_0(.din(w_dff_B_nq3fvDGS9_0),.dout(w_dff_B_fHAgzPVK0_0),.clk(gclk));
	jdff dff_B_sAGoI8hL6_0(.din(w_dff_B_fHAgzPVK0_0),.dout(w_dff_B_sAGoI8hL6_0),.clk(gclk));
	jdff dff_B_7a9JN6SX4_0(.din(w_dff_B_sAGoI8hL6_0),.dout(w_dff_B_7a9JN6SX4_0),.clk(gclk));
	jdff dff_B_XGKfbu7B3_0(.din(n375),.dout(w_dff_B_XGKfbu7B3_0),.clk(gclk));
	jdff dff_B_kobm6ENd0_0(.din(w_dff_B_XGKfbu7B3_0),.dout(w_dff_B_kobm6ENd0_0),.clk(gclk));
	jdff dff_B_pZXeD6dm7_0(.din(w_dff_B_kobm6ENd0_0),.dout(w_dff_B_pZXeD6dm7_0),.clk(gclk));
	jdff dff_B_hosz5vSi9_0(.din(w_dff_B_pZXeD6dm7_0),.dout(w_dff_B_hosz5vSi9_0),.clk(gclk));
	jdff dff_B_FNrHhMWb6_0(.din(w_dff_B_hosz5vSi9_0),.dout(w_dff_B_FNrHhMWb6_0),.clk(gclk));
	jdff dff_B_p4N9zMSy3_0(.din(n368),.dout(w_dff_B_p4N9zMSy3_0),.clk(gclk));
	jdff dff_B_pi2wFGve7_0(.din(w_dff_B_p4N9zMSy3_0),.dout(w_dff_B_pi2wFGve7_0),.clk(gclk));
	jdff dff_B_IlWIID078_0(.din(w_dff_B_pi2wFGve7_0),.dout(w_dff_B_IlWIID078_0),.clk(gclk));
	jdff dff_B_DQGuZUL71_0(.din(w_dff_B_IlWIID078_0),.dout(w_dff_B_DQGuZUL71_0),.clk(gclk));
	jdff dff_B_4oR1tRUd7_0(.din(w_dff_B_DQGuZUL71_0),.dout(w_dff_B_4oR1tRUd7_0),.clk(gclk));
	jdff dff_B_LBG5OWJQ7_0(.din(w_dff_B_4oR1tRUd7_0),.dout(w_dff_B_LBG5OWJQ7_0),.clk(gclk));
	jdff dff_B_WdIU6xvz1_0(.din(w_dff_B_LBG5OWJQ7_0),.dout(w_dff_B_WdIU6xvz1_0),.clk(gclk));
	jdff dff_B_OcyUjgvv4_0(.din(w_dff_B_WdIU6xvz1_0),.dout(w_dff_B_OcyUjgvv4_0),.clk(gclk));
	jdff dff_B_NgN9tBnN1_0(.din(w_dff_B_OcyUjgvv4_0),.dout(w_dff_B_NgN9tBnN1_0),.clk(gclk));
	jdff dff_A_V6zhMGb76_1(.dout(w_n367_0[1]),.din(w_dff_A_V6zhMGb76_1),.clk(gclk));
	jdff dff_A_K4s2Dg1J8_1(.dout(w_dff_A_V6zhMGb76_1),.din(w_dff_A_K4s2Dg1J8_1),.clk(gclk));
	jdff dff_A_WN9MZPBm3_1(.dout(w_dff_A_K4s2Dg1J8_1),.din(w_dff_A_WN9MZPBm3_1),.clk(gclk));
	jdff dff_A_J06Ca8h29_1(.dout(w_dff_A_WN9MZPBm3_1),.din(w_dff_A_J06Ca8h29_1),.clk(gclk));
	jdff dff_A_prDYwrzb7_1(.dout(w_dff_A_J06Ca8h29_1),.din(w_dff_A_prDYwrzb7_1),.clk(gclk));
	jdff dff_A_jPujGZjQ0_1(.dout(w_dff_A_prDYwrzb7_1),.din(w_dff_A_jPujGZjQ0_1),.clk(gclk));
	jdff dff_A_BDMPWaHy9_1(.dout(w_dff_A_jPujGZjQ0_1),.din(w_dff_A_BDMPWaHy9_1),.clk(gclk));
	jdff dff_A_hj6QrRjR0_1(.dout(w_dff_A_BDMPWaHy9_1),.din(w_dff_A_hj6QrRjR0_1),.clk(gclk));
	jdff dff_A_I9eTOsSs8_1(.dout(w_dff_A_hj6QrRjR0_1),.din(w_dff_A_I9eTOsSs8_1),.clk(gclk));
	jdff dff_B_6G9LXMK19_1(.din(n294),.dout(w_dff_B_6G9LXMK19_1),.clk(gclk));
	jdff dff_B_1RVjmJHb9_1(.din(w_dff_B_6G9LXMK19_1),.dout(w_dff_B_1RVjmJHb9_1),.clk(gclk));
	jdff dff_B_oKw6tXG59_1(.din(w_dff_B_1RVjmJHb9_1),.dout(w_dff_B_oKw6tXG59_1),.clk(gclk));
	jdff dff_A_CUi5cSKk9_1(.dout(w_G159gat_1[1]),.din(w_dff_A_CUi5cSKk9_1),.clk(gclk));
	jdff dff_A_Uld0OURf3_1(.dout(w_dff_A_CUi5cSKk9_1),.din(w_dff_A_Uld0OURf3_1),.clk(gclk));
	jdff dff_A_2EdkuGeC3_1(.dout(w_dff_A_Uld0OURf3_1),.din(w_dff_A_2EdkuGeC3_1),.clk(gclk));
	jdff dff_A_hXGbQzsN6_1(.dout(w_dff_A_2EdkuGeC3_1),.din(w_dff_A_hXGbQzsN6_1),.clk(gclk));
	jdff dff_A_5wYUwuVt7_1(.dout(w_dff_A_hXGbQzsN6_1),.din(w_dff_A_5wYUwuVt7_1),.clk(gclk));
	jdff dff_A_ZUa6FsL69_1(.dout(w_dff_A_5wYUwuVt7_1),.din(w_dff_A_ZUa6FsL69_1),.clk(gclk));
	jdff dff_A_9OHafTkt0_1(.dout(w_dff_A_ZUa6FsL69_1),.din(w_dff_A_9OHafTkt0_1),.clk(gclk));
	jdff dff_A_201kpSRp5_2(.dout(w_G159gat_1[2]),.din(w_dff_A_201kpSRp5_2),.clk(gclk));
	jdff dff_A_259hgUSJ5_2(.dout(w_dff_A_201kpSRp5_2),.din(w_dff_A_259hgUSJ5_2),.clk(gclk));
	jdff dff_A_CCTWhhIh1_2(.dout(w_dff_A_259hgUSJ5_2),.din(w_dff_A_CCTWhhIh1_2),.clk(gclk));
	jdff dff_A_hBuj7yyj4_2(.dout(w_dff_A_CCTWhhIh1_2),.din(w_dff_A_hBuj7yyj4_2),.clk(gclk));
	jdff dff_A_ZNSlLW4L0_2(.dout(w_dff_A_hBuj7yyj4_2),.din(w_dff_A_ZNSlLW4L0_2),.clk(gclk));
	jdff dff_A_kMFyP6AF2_2(.dout(w_dff_A_ZNSlLW4L0_2),.din(w_dff_A_kMFyP6AF2_2),.clk(gclk));
	jdff dff_A_vqEMsjDs5_2(.dout(w_dff_A_kMFyP6AF2_2),.din(w_dff_A_vqEMsjDs5_2),.clk(gclk));
	jdff dff_A_CFrdlXM94_2(.dout(w_G159gat_0[2]),.din(w_dff_A_CFrdlXM94_2),.clk(gclk));
	jdff dff_A_5lW1YvpY6_2(.dout(w_dff_A_CFrdlXM94_2),.din(w_dff_A_5lW1YvpY6_2),.clk(gclk));
	jdff dff_A_9SqySWtc3_2(.dout(w_dff_A_5lW1YvpY6_2),.din(w_dff_A_9SqySWtc3_2),.clk(gclk));
	jdff dff_A_lL6cgLL13_2(.dout(w_dff_A_9SqySWtc3_2),.din(w_dff_A_lL6cgLL13_2),.clk(gclk));
	jdff dff_B_XR8PMdAH1_0(.din(n365),.dout(w_dff_B_XR8PMdAH1_0),.clk(gclk));
	jdff dff_B_a33JBwVM7_0(.din(w_dff_B_XR8PMdAH1_0),.dout(w_dff_B_a33JBwVM7_0),.clk(gclk));
	jdff dff_B_k4kf8T8c1_0(.din(w_dff_B_a33JBwVM7_0),.dout(w_dff_B_k4kf8T8c1_0),.clk(gclk));
	jdff dff_B_Oj41tBd14_0(.din(w_dff_B_k4kf8T8c1_0),.dout(w_dff_B_Oj41tBd14_0),.clk(gclk));
	jdff dff_A_1bvlYosF7_1(.dout(w_n339_0[1]),.din(w_dff_A_1bvlYosF7_1),.clk(gclk));
	jdff dff_A_7TCj7ijA7_1(.dout(w_dff_A_1bvlYosF7_1),.din(w_dff_A_7TCj7ijA7_1),.clk(gclk));
	jdff dff_A_RrDniVTh0_1(.dout(w_dff_A_7TCj7ijA7_1),.din(w_dff_A_RrDniVTh0_1),.clk(gclk));
	jdff dff_A_16O2qm1c0_1(.dout(w_dff_A_RrDniVTh0_1),.din(w_dff_A_16O2qm1c0_1),.clk(gclk));
	jdff dff_B_C4Dvv0t19_1(.din(n333),.dout(w_dff_B_C4Dvv0t19_1),.clk(gclk));
	jdff dff_B_sgQOOH0F8_1(.din(w_dff_B_C4Dvv0t19_1),.dout(w_dff_B_sgQOOH0F8_1),.clk(gclk));
	jdff dff_B_jLQujL9a6_1(.din(w_dff_B_sgQOOH0F8_1),.dout(w_dff_B_jLQujL9a6_1),.clk(gclk));
	jdff dff_B_ukEnEh6a8_0(.din(n363),.dout(w_dff_B_ukEnEh6a8_0),.clk(gclk));
	jdff dff_B_f95Zyvt28_0(.din(w_dff_B_ukEnEh6a8_0),.dout(w_dff_B_f95Zyvt28_0),.clk(gclk));
	jdff dff_B_maOir8CZ6_0(.din(w_dff_B_f95Zyvt28_0),.dout(w_dff_B_maOir8CZ6_0),.clk(gclk));
	jdff dff_B_XoYr91NN9_0(.din(w_dff_B_maOir8CZ6_0),.dout(w_dff_B_XoYr91NN9_0),.clk(gclk));
	jdff dff_A_i04SvP2Y7_1(.dout(w_n331_0[1]),.din(w_dff_A_i04SvP2Y7_1),.clk(gclk));
	jdff dff_A_8dkBumGM4_1(.dout(w_dff_A_i04SvP2Y7_1),.din(w_dff_A_8dkBumGM4_1),.clk(gclk));
	jdff dff_A_Dhx21nBw0_1(.dout(w_dff_A_8dkBumGM4_1),.din(w_dff_A_Dhx21nBw0_1),.clk(gclk));
	jdff dff_A_wH5Gg4sN4_1(.dout(w_dff_A_Dhx21nBw0_1),.din(w_dff_A_wH5Gg4sN4_1),.clk(gclk));
	jdff dff_B_GPgp6nAp4_1(.din(n306),.dout(w_dff_B_GPgp6nAp4_1),.clk(gclk));
	jdff dff_B_iJn8jKKa6_1(.din(w_dff_B_GPgp6nAp4_1),.dout(w_dff_B_iJn8jKKa6_1),.clk(gclk));
	jdff dff_B_20IZbmUG6_1(.din(w_dff_B_iJn8jKKa6_1),.dout(w_dff_B_20IZbmUG6_1),.clk(gclk));
	jdff dff_B_HkS9qsD45_1(.din(w_dff_B_20IZbmUG6_1),.dout(w_dff_B_HkS9qsD45_1),.clk(gclk));
	jdff dff_B_BUPKsVHh9_1(.din(w_dff_B_HkS9qsD45_1),.dout(w_dff_B_BUPKsVHh9_1),.clk(gclk));
	jdff dff_B_kRLr6eC78_1(.din(w_dff_B_BUPKsVHh9_1),.dout(w_dff_B_kRLr6eC78_1),.clk(gclk));
	jdff dff_B_ZsmjwWGx2_1(.din(w_dff_B_kRLr6eC78_1),.dout(w_dff_B_ZsmjwWGx2_1),.clk(gclk));
	jdff dff_B_VgUtxseO0_0(.din(n403),.dout(w_dff_B_VgUtxseO0_0),.clk(gclk));
	jdff dff_B_NHLTXGZ07_0(.din(w_dff_B_VgUtxseO0_0),.dout(w_dff_B_NHLTXGZ07_0),.clk(gclk));
	jdff dff_B_COiCVePz9_0(.din(w_dff_B_NHLTXGZ07_0),.dout(w_dff_B_COiCVePz9_0),.clk(gclk));
	jdff dff_B_0fUM2BM80_0(.din(w_dff_B_COiCVePz9_0),.dout(w_dff_B_0fUM2BM80_0),.clk(gclk));
	jdff dff_B_DXuKsD0O9_0(.din(w_dff_B_0fUM2BM80_0),.dout(w_dff_B_DXuKsD0O9_0),.clk(gclk));
	jdff dff_B_7AdnsBA27_0(.din(w_dff_B_DXuKsD0O9_0),.dout(w_dff_B_7AdnsBA27_0),.clk(gclk));
	jdff dff_B_KvpcJOkT2_0(.din(w_dff_B_7AdnsBA27_0),.dout(w_dff_B_KvpcJOkT2_0),.clk(gclk));
	jdff dff_B_zCYoDjUN4_0(.din(w_dff_B_KvpcJOkT2_0),.dout(w_dff_B_zCYoDjUN4_0),.clk(gclk));
	jdff dff_B_aHLx74Sb4_0(.din(w_dff_B_zCYoDjUN4_0),.dout(w_dff_B_aHLx74Sb4_0),.clk(gclk));
	jdff dff_B_ObHH3cAX7_0(.din(w_dff_B_aHLx74Sb4_0),.dout(w_dff_B_ObHH3cAX7_0),.clk(gclk));
	jdff dff_B_dKybQjpE7_0(.din(n401),.dout(w_dff_B_dKybQjpE7_0),.clk(gclk));
	jdff dff_B_0DzC5rDp0_0(.din(w_dff_B_dKybQjpE7_0),.dout(w_dff_B_0DzC5rDp0_0),.clk(gclk));
	jdff dff_B_2t9vMCFu3_0(.din(n400),.dout(w_dff_B_2t9vMCFu3_0),.clk(gclk));
	jdff dff_B_gTN7xQnf8_0(.din(w_dff_B_2t9vMCFu3_0),.dout(w_dff_B_gTN7xQnf8_0),.clk(gclk));
	jdff dff_B_pwnW2eiY9_0(.din(w_dff_B_gTN7xQnf8_0),.dout(w_dff_B_pwnW2eiY9_0),.clk(gclk));
	jdff dff_B_ImGLq4gj7_0(.din(w_dff_B_pwnW2eiY9_0),.dout(w_dff_B_ImGLq4gj7_0),.clk(gclk));
	jdff dff_A_1j4UG0cm6_1(.dout(w_G91gat_0[1]),.din(w_dff_A_1j4UG0cm6_1),.clk(gclk));
	jdff dff_A_4OOSH44w8_1(.dout(w_dff_A_1j4UG0cm6_1),.din(w_dff_A_4OOSH44w8_1),.clk(gclk));
	jdff dff_A_IrK88W3t1_1(.dout(w_dff_A_4OOSH44w8_1),.din(w_dff_A_IrK88W3t1_1),.clk(gclk));
	jdff dff_A_9qqrJkE60_1(.dout(w_dff_A_IrK88W3t1_1),.din(w_dff_A_9qqrJkE60_1),.clk(gclk));
	jdff dff_A_X1OJdXbj3_1(.dout(w_dff_A_9qqrJkE60_1),.din(w_dff_A_X1OJdXbj3_1),.clk(gclk));
	jdff dff_B_JiGp95Kg4_0(.din(n397),.dout(w_dff_B_JiGp95Kg4_0),.clk(gclk));
	jdff dff_B_TFm4noDO6_0(.din(w_dff_B_JiGp95Kg4_0),.dout(w_dff_B_TFm4noDO6_0),.clk(gclk));
	jdff dff_B_RTezwXI73_0(.din(w_dff_B_TFm4noDO6_0),.dout(w_dff_B_RTezwXI73_0),.clk(gclk));
	jdff dff_B_lNHmu34x3_0(.din(w_dff_B_RTezwXI73_0),.dout(w_dff_B_lNHmu34x3_0),.clk(gclk));
	jdff dff_B_jvsOuxFA9_0(.din(w_dff_B_lNHmu34x3_0),.dout(w_dff_B_jvsOuxFA9_0),.clk(gclk));
	jdff dff_B_4rke9fUf9_1(.din(n384),.dout(w_dff_B_4rke9fUf9_1),.clk(gclk));
	jdff dff_B_sV1MvrWv7_1(.din(w_dff_B_4rke9fUf9_1),.dout(w_dff_B_sV1MvrWv7_1),.clk(gclk));
	jdff dff_B_Gkam16Qx8_1(.din(w_dff_B_sV1MvrWv7_1),.dout(w_dff_B_Gkam16Qx8_1),.clk(gclk));
	jdff dff_B_rGM53A5o9_1(.din(w_dff_B_Gkam16Qx8_1),.dout(w_dff_B_rGM53A5o9_1),.clk(gclk));
	jdff dff_B_VZdcpzdW2_1(.din(w_dff_B_rGM53A5o9_1),.dout(w_dff_B_VZdcpzdW2_1),.clk(gclk));
	jdff dff_B_eZK03X1m8_1(.din(w_dff_B_VZdcpzdW2_1),.dout(w_dff_B_eZK03X1m8_1),.clk(gclk));
	jdff dff_B_gK09yN0x5_1(.din(w_dff_B_eZK03X1m8_1),.dout(w_dff_B_gK09yN0x5_1),.clk(gclk));
	jdff dff_B_qvWiE8fs9_1(.din(w_dff_B_gK09yN0x5_1),.dout(w_dff_B_qvWiE8fs9_1),.clk(gclk));
	jdff dff_B_1pd4Ccwh2_1(.din(w_dff_B_qvWiE8fs9_1),.dout(w_dff_B_1pd4Ccwh2_1),.clk(gclk));
	jdff dff_B_prFWXAF80_1(.din(n385),.dout(w_dff_B_prFWXAF80_1),.clk(gclk));
	jdff dff_B_g8rE8TPU0_1(.din(w_dff_B_prFWXAF80_1),.dout(w_dff_B_g8rE8TPU0_1),.clk(gclk));
	jdff dff_B_mTeFZ3c33_1(.din(w_dff_B_g8rE8TPU0_1),.dout(w_dff_B_mTeFZ3c33_1),.clk(gclk));
	jdff dff_B_gPEb4QjS6_1(.din(w_dff_B_mTeFZ3c33_1),.dout(w_dff_B_gPEb4QjS6_1),.clk(gclk));
	jdff dff_B_ozykzldL0_1(.din(w_dff_B_gPEb4QjS6_1),.dout(w_dff_B_ozykzldL0_1),.clk(gclk));
	jdff dff_B_7R9s9ooO7_1(.din(w_dff_B_ozykzldL0_1),.dout(w_dff_B_7R9s9ooO7_1),.clk(gclk));
	jdff dff_B_zPTo8wku1_0(.din(n386),.dout(w_dff_B_zPTo8wku1_0),.clk(gclk));
	jdff dff_B_PBYuE5wH7_0(.din(w_dff_B_zPTo8wku1_0),.dout(w_dff_B_PBYuE5wH7_0),.clk(gclk));
	jdff dff_B_N1VuPPoD6_0(.din(w_dff_B_PBYuE5wH7_0),.dout(w_dff_B_N1VuPPoD6_0),.clk(gclk));
	jdff dff_B_vRlCJ29I2_0(.din(w_dff_B_N1VuPPoD6_0),.dout(w_dff_B_vRlCJ29I2_0),.clk(gclk));
	jdff dff_B_cs0Dx8UG2_0(.din(w_dff_B_vRlCJ29I2_0),.dout(w_dff_B_cs0Dx8UG2_0),.clk(gclk));
	jdff dff_B_YUvVzvXC8_0(.din(w_dff_B_cs0Dx8UG2_0),.dout(w_dff_B_YUvVzvXC8_0),.clk(gclk));
	jdff dff_A_s5rCXlAG6_0(.dout(w_n330_0[0]),.din(w_dff_A_s5rCXlAG6_0),.clk(gclk));
	jdff dff_A_6mVfejcr1_0(.dout(w_dff_A_s5rCXlAG6_0),.din(w_dff_A_6mVfejcr1_0),.clk(gclk));
	jdff dff_A_KrcYq9679_0(.dout(w_dff_A_6mVfejcr1_0),.din(w_dff_A_KrcYq9679_0),.clk(gclk));
	jdff dff_A_AZb9FAO09_0(.dout(w_dff_A_KrcYq9679_0),.din(w_dff_A_AZb9FAO09_0),.clk(gclk));
	jdff dff_A_DYCW0Jmy5_0(.dout(w_dff_A_AZb9FAO09_0),.din(w_dff_A_DYCW0Jmy5_0),.clk(gclk));
	jdff dff_A_cIMVAcIE0_0(.dout(w_dff_A_DYCW0Jmy5_0),.din(w_dff_A_cIMVAcIE0_0),.clk(gclk));
	jdff dff_A_YIhTZkIK0_2(.dout(w_n330_0[2]),.din(w_dff_A_YIhTZkIK0_2),.clk(gclk));
	jdff dff_A_mNcjiUTS4_0(.dout(w_n337_0[0]),.din(w_dff_A_mNcjiUTS4_0),.clk(gclk));
	jdff dff_A_zPYlU2wa5_0(.dout(w_dff_A_mNcjiUTS4_0),.din(w_dff_A_zPYlU2wa5_0),.clk(gclk));
	jdff dff_A_8OGcqSg49_0(.dout(w_dff_A_zPYlU2wa5_0),.din(w_dff_A_8OGcqSg49_0),.clk(gclk));
	jdff dff_A_gw4B2maH7_0(.dout(w_dff_A_8OGcqSg49_0),.din(w_dff_A_gw4B2maH7_0),.clk(gclk));
	jdff dff_A_2UTuchFl9_0(.dout(w_dff_A_gw4B2maH7_0),.din(w_dff_A_2UTuchFl9_0),.clk(gclk));
	jdff dff_A_NjUnijN24_0(.dout(w_dff_A_2UTuchFl9_0),.din(w_dff_A_NjUnijN24_0),.clk(gclk));
	jdff dff_B_FE3FwbSM1_1(.din(n334),.dout(w_dff_B_FE3FwbSM1_1),.clk(gclk));
	jdff dff_A_5nyxg60e1_0(.dout(w_G171gat_2[0]),.din(w_dff_A_5nyxg60e1_0),.clk(gclk));
	jdff dff_A_IuWTlpDl7_0(.dout(w_dff_A_5nyxg60e1_0),.din(w_dff_A_IuWTlpDl7_0),.clk(gclk));
	jdff dff_A_z1KooGNv4_0(.dout(w_dff_A_IuWTlpDl7_0),.din(w_dff_A_z1KooGNv4_0),.clk(gclk));
	jdff dff_A_u0cpHpTX4_0(.dout(w_dff_A_z1KooGNv4_0),.din(w_dff_A_u0cpHpTX4_0),.clk(gclk));
	jdff dff_A_mZxIiWQ83_0(.dout(w_dff_A_u0cpHpTX4_0),.din(w_dff_A_mZxIiWQ83_0),.clk(gclk));
	jdff dff_A_pW4y1Ak80_0(.dout(w_dff_A_mZxIiWQ83_0),.din(w_dff_A_pW4y1Ak80_0),.clk(gclk));
	jdff dff_A_k6DoSIxV4_0(.dout(w_dff_A_pW4y1Ak80_0),.din(w_dff_A_k6DoSIxV4_0),.clk(gclk));
	jdff dff_A_zVmWF26z1_1(.dout(w_n383_0[1]),.din(w_dff_A_zVmWF26z1_1),.clk(gclk));
	jdff dff_A_BRUnb4Ww5_1(.dout(w_dff_A_zVmWF26z1_1),.din(w_dff_A_BRUnb4Ww5_1),.clk(gclk));
	jdff dff_A_d7y0z4AG3_1(.dout(w_dff_A_BRUnb4Ww5_1),.din(w_dff_A_d7y0z4AG3_1),.clk(gclk));
	jdff dff_A_OBdixHz37_1(.dout(w_dff_A_d7y0z4AG3_1),.din(w_dff_A_OBdixHz37_1),.clk(gclk));
	jdff dff_A_xZZX1C1g8_1(.dout(w_dff_A_OBdixHz37_1),.din(w_dff_A_xZZX1C1g8_1),.clk(gclk));
	jdff dff_A_Yi1MI5Qq2_1(.dout(w_dff_A_xZZX1C1g8_1),.din(w_dff_A_Yi1MI5Qq2_1),.clk(gclk));
	jdff dff_A_cZ3dTSwV8_1(.dout(w_dff_A_Yi1MI5Qq2_1),.din(w_dff_A_cZ3dTSwV8_1),.clk(gclk));
	jdff dff_A_QKmOS0196_1(.dout(w_dff_A_cZ3dTSwV8_1),.din(w_dff_A_QKmOS0196_1),.clk(gclk));
	jdff dff_A_hma2NagD0_1(.dout(w_dff_A_QKmOS0196_1),.din(w_dff_A_hma2NagD0_1),.clk(gclk));
	jdff dff_B_spsMgE7k2_0(.din(n309),.dout(w_dff_B_spsMgE7k2_0),.clk(gclk));
	jdff dff_B_HxHEbcII6_0(.din(w_dff_B_spsMgE7k2_0),.dout(w_dff_B_HxHEbcII6_0),.clk(gclk));
	jdff dff_B_lCxEUWz72_0(.din(w_dff_B_HxHEbcII6_0),.dout(w_dff_B_lCxEUWz72_0),.clk(gclk));
	jdff dff_A_CVFts5Eh3_1(.dout(w_G165gat_1[1]),.din(w_dff_A_CVFts5Eh3_1),.clk(gclk));
	jdff dff_A_6rQmRFlr7_1(.dout(w_dff_A_CVFts5Eh3_1),.din(w_dff_A_6rQmRFlr7_1),.clk(gclk));
	jdff dff_A_bNm6HBDy8_1(.dout(w_dff_A_6rQmRFlr7_1),.din(w_dff_A_bNm6HBDy8_1),.clk(gclk));
	jdff dff_A_SNkIjNkL5_1(.dout(w_dff_A_bNm6HBDy8_1),.din(w_dff_A_SNkIjNkL5_1),.clk(gclk));
	jdff dff_A_wgtPdGVE7_1(.dout(w_dff_A_SNkIjNkL5_1),.din(w_dff_A_wgtPdGVE7_1),.clk(gclk));
	jdff dff_A_00tgw1860_1(.dout(w_dff_A_wgtPdGVE7_1),.din(w_dff_A_00tgw1860_1),.clk(gclk));
	jdff dff_A_4yaqyCEp6_1(.dout(w_dff_A_00tgw1860_1),.din(w_dff_A_4yaqyCEp6_1),.clk(gclk));
	jdff dff_A_EWSSpqNB4_2(.dout(w_G165gat_1[2]),.din(w_dff_A_EWSSpqNB4_2),.clk(gclk));
	jdff dff_A_mvQ2J5K39_2(.dout(w_dff_A_EWSSpqNB4_2),.din(w_dff_A_mvQ2J5K39_2),.clk(gclk));
	jdff dff_A_FgcSLf711_2(.dout(w_dff_A_mvQ2J5K39_2),.din(w_dff_A_FgcSLf711_2),.clk(gclk));
	jdff dff_A_6uBggni70_2(.dout(w_dff_A_FgcSLf711_2),.din(w_dff_A_6uBggni70_2),.clk(gclk));
	jdff dff_A_1wDC8Hp87_2(.dout(w_dff_A_6uBggni70_2),.din(w_dff_A_1wDC8Hp87_2),.clk(gclk));
	jdff dff_A_sENeX9xq0_2(.dout(w_dff_A_1wDC8Hp87_2),.din(w_dff_A_sENeX9xq0_2),.clk(gclk));
	jdff dff_A_ZrpWIYCz2_2(.dout(w_dff_A_sENeX9xq0_2),.din(w_dff_A_ZrpWIYCz2_2),.clk(gclk));
	jdff dff_A_51SqRrIP5_2(.dout(w_G165gat_0[2]),.din(w_dff_A_51SqRrIP5_2),.clk(gclk));
	jdff dff_A_Fr8kzAYO2_2(.dout(w_dff_A_51SqRrIP5_2),.din(w_dff_A_Fr8kzAYO2_2),.clk(gclk));
	jdff dff_A_pkDTK9Bw3_2(.dout(w_dff_A_Fr8kzAYO2_2),.din(w_dff_A_pkDTK9Bw3_2),.clk(gclk));
	jdff dff_A_jWD1m8Ga0_2(.dout(w_dff_A_pkDTK9Bw3_2),.din(w_dff_A_jWD1m8Ga0_2),.clk(gclk));
	jdff dff_B_LewbkPHH6_0(.din(n425),.dout(w_dff_B_LewbkPHH6_0),.clk(gclk));
	jdff dff_B_3AECi5ED9_0(.din(w_dff_B_LewbkPHH6_0),.dout(w_dff_B_3AECi5ED9_0),.clk(gclk));
	jdff dff_B_iE6YmXYw3_0(.din(w_dff_B_3AECi5ED9_0),.dout(w_dff_B_iE6YmXYw3_0),.clk(gclk));
	jdff dff_B_oz6HQKjY0_0(.din(w_dff_B_iE6YmXYw3_0),.dout(w_dff_B_oz6HQKjY0_0),.clk(gclk));
	jdff dff_B_jVvkZzmh1_0(.din(w_dff_B_oz6HQKjY0_0),.dout(w_dff_B_jVvkZzmh1_0),.clk(gclk));
	jdff dff_B_TDcSGP7N1_0(.din(w_dff_B_jVvkZzmh1_0),.dout(w_dff_B_TDcSGP7N1_0),.clk(gclk));
	jdff dff_B_WlDYEft91_0(.din(w_dff_B_TDcSGP7N1_0),.dout(w_dff_B_WlDYEft91_0),.clk(gclk));
	jdff dff_B_XtXhwEY92_0(.din(w_dff_B_WlDYEft91_0),.dout(w_dff_B_XtXhwEY92_0),.clk(gclk));
	jdff dff_B_0hzHmD3M5_0(.din(w_dff_B_XtXhwEY92_0),.dout(w_dff_B_0hzHmD3M5_0),.clk(gclk));
	jdff dff_B_Nigc0Z265_0(.din(w_dff_B_0hzHmD3M5_0),.dout(w_dff_B_Nigc0Z265_0),.clk(gclk));
	jdff dff_B_QbUYHx6i4_0(.din(n423),.dout(w_dff_B_QbUYHx6i4_0),.clk(gclk));
	jdff dff_B_7HwCOTBq1_0(.din(w_dff_B_QbUYHx6i4_0),.dout(w_dff_B_7HwCOTBq1_0),.clk(gclk));
	jdff dff_B_QN60WPBm1_0(.din(n422),.dout(w_dff_B_QN60WPBm1_0),.clk(gclk));
	jdff dff_B_ee4C7dX55_0(.din(w_dff_B_QN60WPBm1_0),.dout(w_dff_B_ee4C7dX55_0),.clk(gclk));
	jdff dff_B_IJFyViog8_0(.din(w_dff_B_ee4C7dX55_0),.dout(w_dff_B_IJFyViog8_0),.clk(gclk));
	jdff dff_B_PMLc6udB4_0(.din(w_dff_B_IJFyViog8_0),.dout(w_dff_B_PMLc6udB4_0),.clk(gclk));
	jdff dff_A_oKlz0ELJ7_1(.dout(w_G96gat_0[1]),.din(w_dff_A_oKlz0ELJ7_1),.clk(gclk));
	jdff dff_A_F6F0Br6R1_1(.dout(w_dff_A_oKlz0ELJ7_1),.din(w_dff_A_F6F0Br6R1_1),.clk(gclk));
	jdff dff_A_rkVxnocP7_1(.dout(w_dff_A_F6F0Br6R1_1),.din(w_dff_A_rkVxnocP7_1),.clk(gclk));
	jdff dff_A_p2C2SppA4_1(.dout(w_dff_A_rkVxnocP7_1),.din(w_dff_A_p2C2SppA4_1),.clk(gclk));
	jdff dff_A_vfPBbFAz9_1(.dout(w_dff_A_p2C2SppA4_1),.din(w_dff_A_vfPBbFAz9_1),.clk(gclk));
	jdff dff_B_v1xyCebV4_1(.din(G73gat),.dout(w_dff_B_v1xyCebV4_1),.clk(gclk));
	jdff dff_A_OM48yGBA4_0(.dout(w_n121_0[0]),.din(w_dff_A_OM48yGBA4_0),.clk(gclk));
	jdff dff_A_SA7BZnPm1_0(.dout(w_n118_0[0]),.din(w_dff_A_SA7BZnPm1_0),.clk(gclk));
	jdff dff_B_wfkIujoZ8_0(.din(n419),.dout(w_dff_B_wfkIujoZ8_0),.clk(gclk));
	jdff dff_B_ckaEptPj1_0(.din(w_dff_B_wfkIujoZ8_0),.dout(w_dff_B_ckaEptPj1_0),.clk(gclk));
	jdff dff_B_eeW5rn2X8_0(.din(w_dff_B_ckaEptPj1_0),.dout(w_dff_B_eeW5rn2X8_0),.clk(gclk));
	jdff dff_B_O67J6Nxd7_0(.din(w_dff_B_eeW5rn2X8_0),.dout(w_dff_B_O67J6Nxd7_0),.clk(gclk));
	jdff dff_B_UyJSPswS6_0(.din(w_dff_B_O67J6Nxd7_0),.dout(w_dff_B_UyJSPswS6_0),.clk(gclk));
	jdff dff_B_whdvNOk09_3(.din(G246gat),.dout(w_dff_B_whdvNOk09_3),.clk(gclk));
	jdff dff_A_Nhdao0Dr4_2(.dout(w_G228gat_0[2]),.din(w_dff_A_Nhdao0Dr4_2),.clk(gclk));
	jdff dff_B_jOd7JQF56_3(.din(G228gat),.dout(w_dff_B_jOd7JQF56_3),.clk(gclk));
	jdff dff_B_daADxTze6_3(.din(w_dff_B_jOd7JQF56_3),.dout(w_dff_B_daADxTze6_3),.clk(gclk));
	jdff dff_B_FqcmaZdc7_3(.din(w_dff_B_daADxTze6_3),.dout(w_dff_B_FqcmaZdc7_3),.clk(gclk));
	jdff dff_B_FZZmvEat2_3(.din(w_dff_B_FqcmaZdc7_3),.dout(w_dff_B_FZZmvEat2_3),.clk(gclk));
	jdff dff_B_nvMgiuIL2_3(.din(w_dff_B_FZZmvEat2_3),.dout(w_dff_B_nvMgiuIL2_3),.clk(gclk));
	jdff dff_B_YuRNS4hx1_3(.din(w_dff_B_nvMgiuIL2_3),.dout(w_dff_B_YuRNS4hx1_3),.clk(gclk));
	jdff dff_B_J8ljZcny0_3(.din(w_dff_B_YuRNS4hx1_3),.dout(w_dff_B_J8ljZcny0_3),.clk(gclk));
	jdff dff_B_T91JKijC2_3(.din(w_dff_B_J8ljZcny0_3),.dout(w_dff_B_T91JKijC2_3),.clk(gclk));
	jdff dff_A_rVAjY0GK0_0(.dout(w_G219gat_0[0]),.din(w_dff_A_rVAjY0GK0_0),.clk(gclk));
	jdff dff_A_3Oqe3ufH6_0(.dout(w_dff_A_rVAjY0GK0_0),.din(w_dff_A_3Oqe3ufH6_0),.clk(gclk));
	jdff dff_A_b5e1wHnW1_0(.dout(w_dff_A_3Oqe3ufH6_0),.din(w_dff_A_b5e1wHnW1_0),.clk(gclk));
	jdff dff_A_yx6M2I7s5_0(.dout(w_dff_A_b5e1wHnW1_0),.din(w_dff_A_yx6M2I7s5_0),.clk(gclk));
	jdff dff_A_eVvwObL41_0(.dout(w_dff_A_yx6M2I7s5_0),.din(w_dff_A_eVvwObL41_0),.clk(gclk));
	jdff dff_A_RYFJvG568_0(.dout(w_dff_A_eVvwObL41_0),.din(w_dff_A_RYFJvG568_0),.clk(gclk));
	jdff dff_A_5dfcbgM47_0(.dout(w_dff_A_RYFJvG568_0),.din(w_dff_A_5dfcbgM47_0),.clk(gclk));
	jdff dff_A_t7KS4ed80_0(.dout(w_dff_A_5dfcbgM47_0),.din(w_dff_A_t7KS4ed80_0),.clk(gclk));
	jdff dff_A_18ZhxSlV5_1(.dout(w_G219gat_0[1]),.din(w_dff_A_18ZhxSlV5_1),.clk(gclk));
	jdff dff_A_lIgj2OvW9_1(.dout(w_dff_A_18ZhxSlV5_1),.din(w_dff_A_lIgj2OvW9_1),.clk(gclk));
	jdff dff_B_O9oLpDuU0_3(.din(G219gat),.dout(w_dff_B_O9oLpDuU0_3),.clk(gclk));
	jdff dff_B_R02UGAWA1_3(.din(w_dff_B_O9oLpDuU0_3),.dout(w_dff_B_R02UGAWA1_3),.clk(gclk));
	jdff dff_B_1MraEhNs2_3(.din(w_dff_B_R02UGAWA1_3),.dout(w_dff_B_1MraEhNs2_3),.clk(gclk));
	jdff dff_B_x57ofOHd6_3(.din(w_dff_B_1MraEhNs2_3),.dout(w_dff_B_x57ofOHd6_3),.clk(gclk));
	jdff dff_B_Zgzw6iPU8_3(.din(w_dff_B_x57ofOHd6_3),.dout(w_dff_B_Zgzw6iPU8_3),.clk(gclk));
	jdff dff_B_t2zJa4iU9_3(.din(w_dff_B_Zgzw6iPU8_3),.dout(w_dff_B_t2zJa4iU9_3),.clk(gclk));
	jdff dff_B_UfnRBDC88_3(.din(w_dff_B_t2zJa4iU9_3),.dout(w_dff_B_UfnRBDC88_3),.clk(gclk));
	jdff dff_B_wlsGuj6l3_3(.din(w_dff_B_UfnRBDC88_3),.dout(w_dff_B_wlsGuj6l3_3),.clk(gclk));
	jdff dff_B_uGQMOXZ37_3(.din(w_dff_B_wlsGuj6l3_3),.dout(w_dff_B_uGQMOXZ37_3),.clk(gclk));
	jdff dff_B_nzN8IDbZ5_3(.din(w_dff_B_uGQMOXZ37_3),.dout(w_dff_B_nzN8IDbZ5_3),.clk(gclk));
	jdff dff_B_V3pupD2l2_1(.din(n406),.dout(w_dff_B_V3pupD2l2_1),.clk(gclk));
	jdff dff_B_kkK3U1ve9_1(.din(w_dff_B_V3pupD2l2_1),.dout(w_dff_B_kkK3U1ve9_1),.clk(gclk));
	jdff dff_B_qV8ONmbE7_1(.din(w_dff_B_kkK3U1ve9_1),.dout(w_dff_B_qV8ONmbE7_1),.clk(gclk));
	jdff dff_B_ymLB1aEk1_1(.din(w_dff_B_qV8ONmbE7_1),.dout(w_dff_B_ymLB1aEk1_1),.clk(gclk));
	jdff dff_B_OhUSpVA47_1(.din(w_dff_B_ymLB1aEk1_1),.dout(w_dff_B_OhUSpVA47_1),.clk(gclk));
	jdff dff_B_Co37Av8c6_1(.din(w_dff_B_OhUSpVA47_1),.dout(w_dff_B_Co37Av8c6_1),.clk(gclk));
	jdff dff_B_pF0LVP5R3_1(.din(w_dff_B_Co37Av8c6_1),.dout(w_dff_B_pF0LVP5R3_1),.clk(gclk));
	jdff dff_B_N4REVMAn7_1(.din(w_dff_B_pF0LVP5R3_1),.dout(w_dff_B_N4REVMAn7_1),.clk(gclk));
	jdff dff_B_bRPOcEi75_1(.din(w_dff_B_N4REVMAn7_1),.dout(w_dff_B_bRPOcEi75_1),.clk(gclk));
	jdff dff_B_H1BwVxyk3_1(.din(n407),.dout(w_dff_B_H1BwVxyk3_1),.clk(gclk));
	jdff dff_B_OV6HhMtM7_1(.din(w_dff_B_H1BwVxyk3_1),.dout(w_dff_B_OV6HhMtM7_1),.clk(gclk));
	jdff dff_B_zw978dEx9_1(.din(w_dff_B_OV6HhMtM7_1),.dout(w_dff_B_zw978dEx9_1),.clk(gclk));
	jdff dff_B_ozOiaOpt3_1(.din(w_dff_B_zw978dEx9_1),.dout(w_dff_B_ozOiaOpt3_1),.clk(gclk));
	jdff dff_B_soCIg1hW9_1(.din(w_dff_B_ozOiaOpt3_1),.dout(w_dff_B_soCIg1hW9_1),.clk(gclk));
	jdff dff_B_JwetYlcX5_1(.din(w_dff_B_soCIg1hW9_1),.dout(w_dff_B_JwetYlcX5_1),.clk(gclk));
	jdff dff_B_AY2Mtqzl2_1(.din(w_dff_B_JwetYlcX5_1),.dout(w_dff_B_AY2Mtqzl2_1),.clk(gclk));
	jdff dff_B_WfuUDdre2_1(.din(w_dff_B_AY2Mtqzl2_1),.dout(w_dff_B_WfuUDdre2_1),.clk(gclk));
	jdff dff_B_qQiaIzkt0_0(.din(n408),.dout(w_dff_B_qQiaIzkt0_0),.clk(gclk));
	jdff dff_B_PPO2YRwi6_0(.din(w_dff_B_qQiaIzkt0_0),.dout(w_dff_B_PPO2YRwi6_0),.clk(gclk));
	jdff dff_B_dRZnWDra1_0(.din(w_dff_B_PPO2YRwi6_0),.dout(w_dff_B_dRZnWDra1_0),.clk(gclk));
	jdff dff_B_gacHT41n2_0(.din(w_dff_B_dRZnWDra1_0),.dout(w_dff_B_gacHT41n2_0),.clk(gclk));
	jdff dff_B_TFk3Smfx4_0(.din(w_dff_B_gacHT41n2_0),.dout(w_dff_B_TFk3Smfx4_0),.clk(gclk));
	jdff dff_B_LIcxoJsr7_0(.din(w_dff_B_TFk3Smfx4_0),.dout(w_dff_B_LIcxoJsr7_0),.clk(gclk));
	jdff dff_B_zhzCgr9l2_0(.din(w_dff_B_LIcxoJsr7_0),.dout(w_dff_B_zhzCgr9l2_0),.clk(gclk));
	jdff dff_A_C5PfbyWd0_0(.dout(w_n329_0[0]),.din(w_dff_A_C5PfbyWd0_0),.clk(gclk));
	jdff dff_A_6P6xMBd96_0(.dout(w_dff_A_C5PfbyWd0_0),.din(w_dff_A_6P6xMBd96_0),.clk(gclk));
	jdff dff_A_mDgRez6e5_0(.dout(w_dff_A_6P6xMBd96_0),.din(w_dff_A_mDgRez6e5_0),.clk(gclk));
	jdff dff_A_S9rtRJqS2_0(.dout(w_dff_A_mDgRez6e5_0),.din(w_dff_A_S9rtRJqS2_0),.clk(gclk));
	jdff dff_A_F09O55e07_0(.dout(w_dff_A_S9rtRJqS2_0),.din(w_dff_A_F09O55e07_0),.clk(gclk));
	jdff dff_A_vNIgRCAi0_0(.dout(w_dff_A_F09O55e07_0),.din(w_dff_A_vNIgRCAi0_0),.clk(gclk));
	jdff dff_A_sEYTIeD96_0(.dout(w_dff_A_vNIgRCAi0_0),.din(w_dff_A_sEYTIeD96_0),.clk(gclk));
	jdff dff_A_E9Adb3CX6_0(.dout(w_G177gat_2[0]),.din(w_dff_A_E9Adb3CX6_0),.clk(gclk));
	jdff dff_A_Ifgm6QmN8_0(.dout(w_dff_A_E9Adb3CX6_0),.din(w_dff_A_Ifgm6QmN8_0),.clk(gclk));
	jdff dff_A_I1hxqBkG5_0(.dout(w_dff_A_Ifgm6QmN8_0),.din(w_dff_A_I1hxqBkG5_0),.clk(gclk));
	jdff dff_A_bS7DxMq41_0(.dout(w_dff_A_I1hxqBkG5_0),.din(w_dff_A_bS7DxMq41_0),.clk(gclk));
	jdff dff_A_OFRLRvej8_0(.dout(w_dff_A_bS7DxMq41_0),.din(w_dff_A_OFRLRvej8_0),.clk(gclk));
	jdff dff_A_nrjRGeno0_0(.dout(w_dff_A_OFRLRvej8_0),.din(w_dff_A_nrjRGeno0_0),.clk(gclk));
	jdff dff_A_oj9M9gvy2_0(.dout(w_dff_A_nrjRGeno0_0),.din(w_dff_A_oj9M9gvy2_0),.clk(gclk));
	jdff dff_B_1uOhd1uu6_1(.din(n343),.dout(w_dff_B_1uOhd1uu6_1),.clk(gclk));
	jdff dff_B_o8rM7Yca6_1(.din(w_dff_B_1uOhd1uu6_1),.dout(w_dff_B_o8rM7Yca6_1),.clk(gclk));
	jdff dff_B_IyqeUokb7_1(.din(w_dff_B_o8rM7Yca6_1),.dout(w_dff_B_IyqeUokb7_1),.clk(gclk));
	jdff dff_B_hvMQNGkC2_1(.din(w_dff_B_IyqeUokb7_1),.dout(w_dff_B_hvMQNGkC2_1),.clk(gclk));
	jdff dff_B_xNk9LDaO0_1(.din(w_dff_B_hvMQNGkC2_1),.dout(w_dff_B_xNk9LDaO0_1),.clk(gclk));
	jdff dff_B_zKiMtKk26_1(.din(n344),.dout(w_dff_B_zKiMtKk26_1),.clk(gclk));
	jdff dff_B_whaycpAI9_1(.din(w_dff_B_zKiMtKk26_1),.dout(w_dff_B_whaycpAI9_1),.clk(gclk));
	jdff dff_B_fILuNpqi9_1(.din(w_dff_B_whaycpAI9_1),.dout(w_dff_B_fILuNpqi9_1),.clk(gclk));
	jdff dff_B_GIwfvGCa0_1(.din(w_dff_B_fILuNpqi9_1),.dout(w_dff_B_GIwfvGCa0_1),.clk(gclk));
	jdff dff_B_q2cswN5H8_0(.din(n231),.dout(w_dff_B_q2cswN5H8_0),.clk(gclk));
	jdff dff_A_rPv8zhsi0_0(.dout(w_n230_0[0]),.din(w_dff_A_rPv8zhsi0_0),.clk(gclk));
	jdff dff_B_QlEQ6RiZ3_1(.din(n227),.dout(w_dff_B_QlEQ6RiZ3_1),.clk(gclk));
	jdff dff_A_WOVoZcG36_0(.dout(w_n228_0[0]),.din(w_dff_A_WOVoZcG36_0),.clk(gclk));
	jdff dff_A_84d0TDkI9_0(.dout(w_dff_A_WOVoZcG36_0),.din(w_dff_A_84d0TDkI9_0),.clk(gclk));
	jdff dff_A_gvbS2i9b2_0(.dout(w_dff_A_84d0TDkI9_0),.din(w_dff_A_gvbS2i9b2_0),.clk(gclk));
	jdff dff_A_4EQMkSy42_1(.dout(w_G195gat_1[1]),.din(w_dff_A_4EQMkSy42_1),.clk(gclk));
	jdff dff_A_3L7vHM4g2_1(.dout(w_dff_A_4EQMkSy42_1),.din(w_dff_A_3L7vHM4g2_1),.clk(gclk));
	jdff dff_A_bC5DtVfh7_1(.dout(w_dff_A_3L7vHM4g2_1),.din(w_dff_A_bC5DtVfh7_1),.clk(gclk));
	jdff dff_A_JsRBExNr4_1(.dout(w_dff_A_bC5DtVfh7_1),.din(w_dff_A_JsRBExNr4_1),.clk(gclk));
	jdff dff_A_OLHkUQAD4_1(.dout(w_dff_A_JsRBExNr4_1),.din(w_dff_A_OLHkUQAD4_1),.clk(gclk));
	jdff dff_A_ImafkSlk0_1(.dout(w_dff_A_OLHkUQAD4_1),.din(w_dff_A_ImafkSlk0_1),.clk(gclk));
	jdff dff_A_MYpj7YG87_1(.dout(w_dff_A_ImafkSlk0_1),.din(w_dff_A_MYpj7YG87_1),.clk(gclk));
	jdff dff_A_YXUvDKir7_1(.dout(w_dff_A_MYpj7YG87_1),.din(w_dff_A_YXUvDKir7_1),.clk(gclk));
	jdff dff_A_Ex86Bgfe7_2(.dout(w_G195gat_1[2]),.din(w_dff_A_Ex86Bgfe7_2),.clk(gclk));
	jdff dff_A_47uOJb8k8_2(.dout(w_dff_A_Ex86Bgfe7_2),.din(w_dff_A_47uOJb8k8_2),.clk(gclk));
	jdff dff_A_VoIcRHx63_2(.dout(w_dff_A_47uOJb8k8_2),.din(w_dff_A_VoIcRHx63_2),.clk(gclk));
	jdff dff_A_MOS8ERis5_2(.dout(w_dff_A_VoIcRHx63_2),.din(w_dff_A_MOS8ERis5_2),.clk(gclk));
	jdff dff_A_AeIcqstQ4_2(.dout(w_dff_A_MOS8ERis5_2),.din(w_dff_A_AeIcqstQ4_2),.clk(gclk));
	jdff dff_A_U9wheQsN1_2(.dout(w_dff_A_AeIcqstQ4_2),.din(w_dff_A_U9wheQsN1_2),.clk(gclk));
	jdff dff_A_kBTG5W2H9_2(.dout(w_dff_A_U9wheQsN1_2),.din(w_dff_A_kBTG5W2H9_2),.clk(gclk));
	jdff dff_A_PvdxKnbG1_2(.dout(w_dff_A_kBTG5W2H9_2),.din(w_dff_A_PvdxKnbG1_2),.clk(gclk));
	jdff dff_A_jpLbGSZ38_1(.dout(w_G189gat_1[1]),.din(w_dff_A_jpLbGSZ38_1),.clk(gclk));
	jdff dff_A_HkXStBlK6_1(.dout(w_dff_A_jpLbGSZ38_1),.din(w_dff_A_HkXStBlK6_1),.clk(gclk));
	jdff dff_A_ITAYOnLV4_1(.dout(w_dff_A_HkXStBlK6_1),.din(w_dff_A_ITAYOnLV4_1),.clk(gclk));
	jdff dff_A_cKpffvdx4_1(.dout(w_dff_A_ITAYOnLV4_1),.din(w_dff_A_cKpffvdx4_1),.clk(gclk));
	jdff dff_A_uewzBx6T7_1(.dout(w_dff_A_cKpffvdx4_1),.din(w_dff_A_uewzBx6T7_1),.clk(gclk));
	jdff dff_A_XbUo13MA8_1(.dout(w_dff_A_uewzBx6T7_1),.din(w_dff_A_XbUo13MA8_1),.clk(gclk));
	jdff dff_A_YtUhTfeo9_1(.dout(w_dff_A_XbUo13MA8_1),.din(w_dff_A_YtUhTfeo9_1),.clk(gclk));
	jdff dff_A_galFhZhB6_1(.dout(w_dff_A_YtUhTfeo9_1),.din(w_dff_A_galFhZhB6_1),.clk(gclk));
	jdff dff_A_TJPkR2Tu3_2(.dout(w_G189gat_1[2]),.din(w_dff_A_TJPkR2Tu3_2),.clk(gclk));
	jdff dff_A_5U9LdHQq1_2(.dout(w_dff_A_TJPkR2Tu3_2),.din(w_dff_A_5U9LdHQq1_2),.clk(gclk));
	jdff dff_A_ZUSVhw7t6_2(.dout(w_dff_A_5U9LdHQq1_2),.din(w_dff_A_ZUSVhw7t6_2),.clk(gclk));
	jdff dff_A_vHo74eu67_2(.dout(w_dff_A_ZUSVhw7t6_2),.din(w_dff_A_vHo74eu67_2),.clk(gclk));
	jdff dff_A_hGdyEgPe1_2(.dout(w_dff_A_vHo74eu67_2),.din(w_dff_A_hGdyEgPe1_2),.clk(gclk));
	jdff dff_A_XJNc4xWq8_2(.dout(w_dff_A_hGdyEgPe1_2),.din(w_dff_A_XJNc4xWq8_2),.clk(gclk));
	jdff dff_A_c8oc95er8_2(.dout(w_dff_A_XJNc4xWq8_2),.din(w_dff_A_c8oc95er8_2),.clk(gclk));
	jdff dff_A_aq6BOP380_2(.dout(w_dff_A_c8oc95er8_2),.din(w_dff_A_aq6BOP380_2),.clk(gclk));
	jdff dff_B_TEqq0CvK2_0(.din(n225),.dout(w_dff_B_TEqq0CvK2_0),.clk(gclk));
	jdff dff_A_ythxWxRF6_0(.dout(w_n224_0[0]),.din(w_dff_A_ythxWxRF6_0),.clk(gclk));
	jdff dff_A_ugzhzE3Q9_0(.dout(w_n223_0[0]),.din(w_dff_A_ugzhzE3Q9_0),.clk(gclk));
	jdff dff_A_6UN2C2Xw2_0(.dout(w_dff_A_ugzhzE3Q9_0),.din(w_dff_A_6UN2C2Xw2_0),.clk(gclk));
	jdff dff_B_uESYCf1D5_1(.din(n219),.dout(w_dff_B_uESYCf1D5_1),.clk(gclk));
	jdff dff_A_Mdeczmo63_0(.dout(w_G121gat_0[0]),.din(w_dff_A_Mdeczmo63_0),.clk(gclk));
	jdff dff_A_wQEL6ZLk0_0(.dout(w_dff_A_Mdeczmo63_0),.din(w_dff_A_wQEL6ZLk0_0),.clk(gclk));
	jdff dff_A_E1MrlAA19_0(.dout(w_dff_A_wQEL6ZLk0_0),.din(w_dff_A_E1MrlAA19_0),.clk(gclk));
	jdff dff_A_TfGSNyHS9_0(.dout(w_dff_A_E1MrlAA19_0),.din(w_dff_A_TfGSNyHS9_0),.clk(gclk));
	jdff dff_A_FKKbzkpB8_0(.dout(w_dff_A_TfGSNyHS9_0),.din(w_dff_A_FKKbzkpB8_0),.clk(gclk));
	jdff dff_A_TxQbYvda3_0(.dout(w_G195gat_2[0]),.din(w_dff_A_TxQbYvda3_0),.clk(gclk));
	jdff dff_A_gZx3R28Z2_0(.dout(w_dff_A_TxQbYvda3_0),.din(w_dff_A_gZx3R28Z2_0),.clk(gclk));
	jdff dff_A_LxCX8sQ08_0(.dout(w_dff_A_gZx3R28Z2_0),.din(w_dff_A_LxCX8sQ08_0),.clk(gclk));
	jdff dff_A_wP8LvX911_0(.dout(w_dff_A_LxCX8sQ08_0),.din(w_dff_A_wP8LvX911_0),.clk(gclk));
	jdff dff_A_1drCJS6Y4_0(.dout(w_dff_A_wP8LvX911_0),.din(w_dff_A_1drCJS6Y4_0),.clk(gclk));
	jdff dff_A_h75rBSBt9_0(.dout(w_dff_A_1drCJS6Y4_0),.din(w_dff_A_h75rBSBt9_0),.clk(gclk));
	jdff dff_A_r67ewH9Y4_0(.dout(w_dff_A_h75rBSBt9_0),.din(w_dff_A_r67ewH9Y4_0),.clk(gclk));
	jdff dff_A_p7ylLqnr5_0(.dout(w_dff_A_r67ewH9Y4_0),.din(w_dff_A_p7ylLqnr5_0),.clk(gclk));
	jdff dff_A_9GKFZAmg5_2(.dout(w_G195gat_0[2]),.din(w_dff_A_9GKFZAmg5_2),.clk(gclk));
	jdff dff_A_lU0Cntqy3_2(.dout(w_dff_A_9GKFZAmg5_2),.din(w_dff_A_lU0Cntqy3_2),.clk(gclk));
	jdff dff_A_DuzjXoJW8_2(.dout(w_dff_A_lU0Cntqy3_2),.din(w_dff_A_DuzjXoJW8_2),.clk(gclk));
	jdff dff_A_rdzFG80g1_2(.dout(w_dff_A_DuzjXoJW8_2),.din(w_dff_A_rdzFG80g1_2),.clk(gclk));
	jdff dff_B_aqjt3HhL1_1(.din(n214),.dout(w_dff_B_aqjt3HhL1_1),.clk(gclk));
	jdff dff_A_PkIF8hws6_1(.dout(w_G116gat_0[1]),.din(w_dff_A_PkIF8hws6_1),.clk(gclk));
	jdff dff_A_L6Dd8G5R1_1(.dout(w_dff_A_PkIF8hws6_1),.din(w_dff_A_L6Dd8G5R1_1),.clk(gclk));
	jdff dff_A_ShOk8JTM8_1(.dout(w_dff_A_L6Dd8G5R1_1),.din(w_dff_A_ShOk8JTM8_1),.clk(gclk));
	jdff dff_A_VNB054K53_1(.dout(w_dff_A_ShOk8JTM8_1),.din(w_dff_A_VNB054K53_1),.clk(gclk));
	jdff dff_A_RO9ze0Q51_1(.dout(w_dff_A_VNB054K53_1),.din(w_dff_A_RO9ze0Q51_1),.clk(gclk));
	jdff dff_A_9OjhhdMe0_1(.dout(w_G146gat_0[1]),.din(w_dff_A_9OjhhdMe0_1),.clk(gclk));
	jdff dff_B_cuGwXApU3_2(.din(G146gat),.dout(w_dff_B_cuGwXApU3_2),.clk(gclk));
	jdff dff_B_o2S9G4eD4_2(.din(w_dff_B_cuGwXApU3_2),.dout(w_dff_B_o2S9G4eD4_2),.clk(gclk));
	jdff dff_B_1cNUGuJs7_2(.din(w_dff_B_o2S9G4eD4_2),.dout(w_dff_B_1cNUGuJs7_2),.clk(gclk));
	jdff dff_B_0BQ6LSLO5_2(.din(w_dff_B_1cNUGuJs7_2),.dout(w_dff_B_0BQ6LSLO5_2),.clk(gclk));
	jdff dff_A_Y5f2zBtt0_0(.dout(w_G189gat_2[0]),.din(w_dff_A_Y5f2zBtt0_0),.clk(gclk));
	jdff dff_A_ikf9a0rw9_0(.dout(w_dff_A_Y5f2zBtt0_0),.din(w_dff_A_ikf9a0rw9_0),.clk(gclk));
	jdff dff_A_gqB3bEwg7_0(.dout(w_dff_A_ikf9a0rw9_0),.din(w_dff_A_gqB3bEwg7_0),.clk(gclk));
	jdff dff_A_n27r3JlS9_0(.dout(w_dff_A_gqB3bEwg7_0),.din(w_dff_A_n27r3JlS9_0),.clk(gclk));
	jdff dff_A_N9bhLb198_0(.dout(w_dff_A_n27r3JlS9_0),.din(w_dff_A_N9bhLb198_0),.clk(gclk));
	jdff dff_A_pgeauC2i2_0(.dout(w_dff_A_N9bhLb198_0),.din(w_dff_A_pgeauC2i2_0),.clk(gclk));
	jdff dff_A_GIMa11pH2_0(.dout(w_dff_A_pgeauC2i2_0),.din(w_dff_A_GIMa11pH2_0),.clk(gclk));
	jdff dff_A_M4yjlATT5_0(.dout(w_dff_A_GIMa11pH2_0),.din(w_dff_A_M4yjlATT5_0),.clk(gclk));
	jdff dff_A_coz4d7269_2(.dout(w_G189gat_0[2]),.din(w_dff_A_coz4d7269_2),.clk(gclk));
	jdff dff_A_pBmMvaYD8_2(.dout(w_dff_A_coz4d7269_2),.din(w_dff_A_pBmMvaYD8_2),.clk(gclk));
	jdff dff_A_nXnt9UZ37_2(.dout(w_dff_A_pBmMvaYD8_2),.din(w_dff_A_nXnt9UZ37_2),.clk(gclk));
	jdff dff_A_XBC0j54E6_2(.dout(w_dff_A_nXnt9UZ37_2),.din(w_dff_A_XBC0j54E6_2),.clk(gclk));
	jdff dff_B_clXIMNx08_1(.din(n197),.dout(w_dff_B_clXIMNx08_1),.clk(gclk));
	jdff dff_B_uNIxL1w15_1(.din(n198),.dout(w_dff_B_uNIxL1w15_1),.clk(gclk));
	jdff dff_B_NEJpFa1Y4_1(.din(w_dff_B_uNIxL1w15_1),.dout(w_dff_B_NEJpFa1Y4_1),.clk(gclk));
	jdff dff_B_dHmHW6Ni5_1(.din(w_dff_B_NEJpFa1Y4_1),.dout(w_dff_B_dHmHW6Ni5_1),.clk(gclk));
	jdff dff_B_6g7n988u1_1(.din(w_dff_B_dHmHW6Ni5_1),.dout(w_dff_B_6g7n988u1_1),.clk(gclk));
	jdff dff_B_acWBpf4X8_1(.din(w_dff_B_6g7n988u1_1),.dout(w_dff_B_acWBpf4X8_1),.clk(gclk));
	jdff dff_B_3DsWS1yx8_1(.din(w_dff_B_acWBpf4X8_1),.dout(w_dff_B_3DsWS1yx8_1),.clk(gclk));
	jdff dff_B_aQp2wqku5_1(.din(w_dff_B_3DsWS1yx8_1),.dout(w_dff_B_aQp2wqku5_1),.clk(gclk));
	jdff dff_B_kgLBemVM5_1(.din(w_dff_B_aQp2wqku5_1),.dout(w_dff_B_kgLBemVM5_1),.clk(gclk));
	jdff dff_B_ZEfKWUgn0_1(.din(n199),.dout(w_dff_B_ZEfKWUgn0_1),.clk(gclk));
	jdff dff_B_5tU4TEeO2_0(.din(n208),.dout(w_dff_B_5tU4TEeO2_0),.clk(gclk));
	jdff dff_B_7ZCE6cac4_0(.din(w_dff_B_5tU4TEeO2_0),.dout(w_dff_B_7ZCE6cac4_0),.clk(gclk));
	jdff dff_B_bmyX14cA2_1(.din(n200),.dout(w_dff_B_bmyX14cA2_1),.clk(gclk));
	jdff dff_B_yHh7Pf790_1(.din(w_dff_B_bmyX14cA2_1),.dout(w_dff_B_yHh7Pf790_1),.clk(gclk));
	jdff dff_B_gRf1Ty346_1(.din(w_dff_B_yHh7Pf790_1),.dout(w_dff_B_gRf1Ty346_1),.clk(gclk));
	jdff dff_B_BN4xaQeZ1_1(.din(w_dff_B_gRf1Ty346_1),.dout(w_dff_B_BN4xaQeZ1_1),.clk(gclk));
	jdff dff_B_vr0TsmQz8_1(.din(w_dff_B_BN4xaQeZ1_1),.dout(w_dff_B_vr0TsmQz8_1),.clk(gclk));
	jdff dff_B_sgSxXV373_1(.din(n201),.dout(w_dff_B_sgSxXV373_1),.clk(gclk));
	jdff dff_B_X9XwSFDQ9_1(.din(w_dff_B_sgSxXV373_1),.dout(w_dff_B_X9XwSFDQ9_1),.clk(gclk));
	jdff dff_B_AYIgoPJz7_1(.din(w_dff_B_X9XwSFDQ9_1),.dout(w_dff_B_AYIgoPJz7_1),.clk(gclk));
	jdff dff_B_WPPIywU42_1(.din(n202),.dout(w_dff_B_WPPIywU42_1),.clk(gclk));
	jdff dff_B_FG5AiP5E0_2(.din(n143),.dout(w_dff_B_FG5AiP5E0_2),.clk(gclk));
	jdff dff_B_JfsPZuPH7_2(.din(w_dff_B_FG5AiP5E0_2),.dout(w_dff_B_JfsPZuPH7_2),.clk(gclk));
	jdff dff_B_QMQtV8nj2_2(.din(w_dff_B_JfsPZuPH7_2),.dout(w_dff_B_QMQtV8nj2_2),.clk(gclk));
	jdff dff_B_snVtZAwb5_2(.din(w_dff_B_QMQtV8nj2_2),.dout(w_dff_B_snVtZAwb5_2),.clk(gclk));
	jdff dff_B_gCXJgSho5_2(.din(w_dff_B_snVtZAwb5_2),.dout(w_dff_B_gCXJgSho5_2),.clk(gclk));
	jdff dff_B_h0h555jf1_2(.din(w_dff_B_gCXJgSho5_2),.dout(w_dff_B_h0h555jf1_2),.clk(gclk));
	jdff dff_B_ffpzhXNI9_2(.din(w_dff_B_h0h555jf1_2),.dout(w_dff_B_ffpzhXNI9_2),.clk(gclk));
	jdff dff_B_MyAcuUYg3_2(.din(w_dff_B_ffpzhXNI9_2),.dout(w_dff_B_MyAcuUYg3_2),.clk(gclk));
	jdff dff_B_Kewu7pk98_2(.din(w_dff_B_MyAcuUYg3_2),.dout(w_dff_B_Kewu7pk98_2),.clk(gclk));
	jdff dff_A_XZbDj4xZ5_0(.dout(w_G261gat_0[0]),.din(w_dff_A_XZbDj4xZ5_0),.clk(gclk));
	jdff dff_A_OMy2n1rb9_0(.dout(w_dff_A_XZbDj4xZ5_0),.din(w_dff_A_OMy2n1rb9_0),.clk(gclk));
	jdff dff_A_VmgtsNXi3_0(.dout(w_dff_A_OMy2n1rb9_0),.din(w_dff_A_VmgtsNXi3_0),.clk(gclk));
	jdff dff_A_l5M72jJp2_0(.dout(w_dff_A_VmgtsNXi3_0),.din(w_dff_A_l5M72jJp2_0),.clk(gclk));
	jdff dff_A_pVfSXInm1_0(.dout(w_dff_A_l5M72jJp2_0),.din(w_dff_A_pVfSXInm1_0),.clk(gclk));
	jdff dff_A_it8krLq24_0(.dout(w_dff_A_pVfSXInm1_0),.din(w_dff_A_it8krLq24_0),.clk(gclk));
	jdff dff_A_OpWZAwtm4_0(.dout(w_dff_A_it8krLq24_0),.din(w_dff_A_OpWZAwtm4_0),.clk(gclk));
	jdff dff_A_HHefhRMK2_0(.dout(w_dff_A_OpWZAwtm4_0),.din(w_dff_A_HHefhRMK2_0),.clk(gclk));
	jdff dff_A_VD6wq4HN3_0(.dout(w_dff_A_HHefhRMK2_0),.din(w_dff_A_VD6wq4HN3_0),.clk(gclk));
	jdff dff_A_QNE8kluf0_1(.dout(w_G261gat_0[1]),.din(w_dff_A_QNE8kluf0_1),.clk(gclk));
	jdff dff_A_xClHQgzr7_1(.dout(w_dff_A_QNE8kluf0_1),.din(w_dff_A_xClHQgzr7_1),.clk(gclk));
	jdff dff_A_HeqR0W707_1(.dout(w_dff_A_xClHQgzr7_1),.din(w_dff_A_HeqR0W707_1),.clk(gclk));
	jdff dff_A_7kdvXk797_1(.dout(w_dff_A_HeqR0W707_1),.din(w_dff_A_7kdvXk797_1),.clk(gclk));
	jdff dff_A_28rE5bO83_1(.dout(w_dff_A_7kdvXk797_1),.din(w_dff_A_28rE5bO83_1),.clk(gclk));
	jdff dff_A_lsXK59Mm0_1(.dout(w_dff_A_28rE5bO83_1),.din(w_dff_A_lsXK59Mm0_1),.clk(gclk));
	jdff dff_A_dplABmtu7_1(.dout(w_dff_A_lsXK59Mm0_1),.din(w_dff_A_dplABmtu7_1),.clk(gclk));
	jdff dff_A_wvSjaXfD5_1(.dout(w_dff_A_dplABmtu7_1),.din(w_dff_A_wvSjaXfD5_1),.clk(gclk));
	jdff dff_A_iiGZ1f197_1(.dout(w_dff_A_wvSjaXfD5_1),.din(w_dff_A_iiGZ1f197_1),.clk(gclk));
	jdff dff_A_P9E7V1247_0(.dout(w_n196_0[0]),.din(w_dff_A_P9E7V1247_0),.clk(gclk));
	jdff dff_A_rxtSPeVE2_1(.dout(w_n154_0[1]),.din(w_dff_A_rxtSPeVE2_1),.clk(gclk));
	jdff dff_A_50LvCA3d3_0(.dout(w_G126gat_0[0]),.din(w_dff_A_50LvCA3d3_0),.clk(gclk));
	jdff dff_A_RUMYQ1GU7_0(.dout(w_dff_A_50LvCA3d3_0),.din(w_dff_A_RUMYQ1GU7_0),.clk(gclk));
	jdff dff_A_SkUdZt1p7_0(.dout(w_dff_A_RUMYQ1GU7_0),.din(w_dff_A_SkUdZt1p7_0),.clk(gclk));
	jdff dff_A_mL6SUM955_0(.dout(w_dff_A_SkUdZt1p7_0),.din(w_dff_A_mL6SUM955_0),.clk(gclk));
	jdff dff_A_SU8vcFnq8_0(.dout(w_dff_A_mL6SUM955_0),.din(w_dff_A_SU8vcFnq8_0),.clk(gclk));
	jdff dff_A_1septHAP6_1(.dout(w_G201gat_1[1]),.din(w_dff_A_1septHAP6_1),.clk(gclk));
	jdff dff_A_dLeIfbgb5_1(.dout(w_dff_A_1septHAP6_1),.din(w_dff_A_dLeIfbgb5_1),.clk(gclk));
	jdff dff_A_7WQ57LK56_1(.dout(w_dff_A_dLeIfbgb5_1),.din(w_dff_A_7WQ57LK56_1),.clk(gclk));
	jdff dff_A_ik8YJjHT4_1(.dout(w_dff_A_7WQ57LK56_1),.din(w_dff_A_ik8YJjHT4_1),.clk(gclk));
	jdff dff_A_acYFoEt74_1(.dout(w_dff_A_ik8YJjHT4_1),.din(w_dff_A_acYFoEt74_1),.clk(gclk));
	jdff dff_A_hHlQe7d67_1(.dout(w_dff_A_acYFoEt74_1),.din(w_dff_A_hHlQe7d67_1),.clk(gclk));
	jdff dff_A_LbhkGPRU4_1(.dout(w_dff_A_hHlQe7d67_1),.din(w_dff_A_LbhkGPRU4_1),.clk(gclk));
	jdff dff_A_RkxdeWDZ7_1(.dout(w_dff_A_LbhkGPRU4_1),.din(w_dff_A_RkxdeWDZ7_1),.clk(gclk));
	jdff dff_A_HcbnxuwG3_2(.dout(w_G201gat_1[2]),.din(w_dff_A_HcbnxuwG3_2),.clk(gclk));
	jdff dff_A_JLQFQzWD1_2(.dout(w_dff_A_HcbnxuwG3_2),.din(w_dff_A_JLQFQzWD1_2),.clk(gclk));
	jdff dff_A_NLHx8rSA3_2(.dout(w_dff_A_JLQFQzWD1_2),.din(w_dff_A_NLHx8rSA3_2),.clk(gclk));
	jdff dff_A_yuUaDZct5_2(.dout(w_dff_A_NLHx8rSA3_2),.din(w_dff_A_yuUaDZct5_2),.clk(gclk));
	jdff dff_A_ZrXyeeNW3_2(.dout(w_G201gat_0[2]),.din(w_dff_A_ZrXyeeNW3_2),.clk(gclk));
	jdff dff_A_nDANibwo2_2(.dout(w_dff_A_ZrXyeeNW3_2),.din(w_dff_A_nDANibwo2_2),.clk(gclk));
	jdff dff_A_pcTaRTIg6_2(.dout(w_dff_A_nDANibwo2_2),.din(w_dff_A_pcTaRTIg6_2),.clk(gclk));
	jdff dff_A_jR9fRiDK2_2(.dout(w_dff_A_pcTaRTIg6_2),.din(w_dff_A_jR9fRiDK2_2),.clk(gclk));
	jdff dff_A_CaeuMWeM4_2(.dout(w_dff_A_jR9fRiDK2_2),.din(w_dff_A_CaeuMWeM4_2),.clk(gclk));
	jdff dff_A_K5QYDIK07_2(.dout(w_dff_A_CaeuMWeM4_2),.din(w_dff_A_K5QYDIK07_2),.clk(gclk));
	jdff dff_A_9ga3GXDX0_2(.dout(w_dff_A_K5QYDIK07_2),.din(w_dff_A_9ga3GXDX0_2),.clk(gclk));
	jdff dff_A_WAjYHuCH9_2(.dout(w_dff_A_9ga3GXDX0_2),.din(w_dff_A_WAjYHuCH9_2),.clk(gclk));
	jdff dff_A_5RgSses18_1(.dout(w_n303_0[1]),.din(w_dff_A_5RgSses18_1),.clk(gclk));
	jdff dff_A_SKGtrvqT2_1(.dout(w_dff_A_5RgSses18_1),.din(w_dff_A_SKGtrvqT2_1),.clk(gclk));
	jdff dff_A_uY4irrfR3_1(.dout(w_dff_A_SKGtrvqT2_1),.din(w_dff_A_uY4irrfR3_1),.clk(gclk));
	jdff dff_A_JO6lxcXS8_1(.dout(w_dff_A_uY4irrfR3_1),.din(w_dff_A_JO6lxcXS8_1),.clk(gclk));
	jdff dff_A_RLcVChcq6_1(.dout(w_n302_0[1]),.din(w_dff_A_RLcVChcq6_1),.clk(gclk));
	jdff dff_A_IRRUgXBZ4_1(.dout(w_dff_A_RLcVChcq6_1),.din(w_dff_A_IRRUgXBZ4_1),.clk(gclk));
	jdff dff_A_KNWiplwD2_1(.dout(w_dff_A_IRRUgXBZ4_1),.din(w_dff_A_KNWiplwD2_1),.clk(gclk));
	jdff dff_A_llG7awQD0_1(.dout(w_dff_A_KNWiplwD2_1),.din(w_dff_A_llG7awQD0_1),.clk(gclk));
	jdff dff_A_GyEHmUoP2_1(.dout(w_dff_A_llG7awQD0_1),.din(w_dff_A_GyEHmUoP2_1),.clk(gclk));
	jdff dff_B_41bkNbQJ2_1(.din(n190),.dout(w_dff_B_41bkNbQJ2_1),.clk(gclk));
	jdff dff_A_wmwB03id7_1(.dout(w_G111gat_0[1]),.din(w_dff_A_wmwB03id7_1),.clk(gclk));
	jdff dff_A_S1hGICed4_1(.dout(w_dff_A_wmwB03id7_1),.din(w_dff_A_S1hGICed4_1),.clk(gclk));
	jdff dff_A_e02uxWhd3_1(.dout(w_dff_A_S1hGICed4_1),.din(w_dff_A_e02uxWhd3_1),.clk(gclk));
	jdff dff_A_w79Okj218_1(.dout(w_dff_A_e02uxWhd3_1),.din(w_dff_A_w79Okj218_1),.clk(gclk));
	jdff dff_A_DZe664RI1_1(.dout(w_dff_A_w79Okj218_1),.din(w_dff_A_DZe664RI1_1),.clk(gclk));
	jdff dff_A_yBSFLR1Y2_1(.dout(w_n165_1[1]),.din(w_dff_A_yBSFLR1Y2_1),.clk(gclk));
	jdff dff_A_JMRI1rol2_1(.dout(w_dff_A_yBSFLR1Y2_1),.din(w_dff_A_JMRI1rol2_1),.clk(gclk));
	jdff dff_A_rwupaW538_2(.dout(w_n165_1[2]),.din(w_dff_A_rwupaW538_2),.clk(gclk));
	jdff dff_A_ksVZSOd59_2(.dout(w_dff_A_rwupaW538_2),.din(w_dff_A_ksVZSOd59_2),.clk(gclk));
	jdff dff_A_Ar8F1l249_1(.dout(w_n165_0[1]),.din(w_dff_A_Ar8F1l249_1),.clk(gclk));
	jdff dff_A_KLPTewSx0_1(.dout(w_dff_A_Ar8F1l249_1),.din(w_dff_A_KLPTewSx0_1),.clk(gclk));
	jdff dff_A_pQu9YZul1_2(.dout(w_n165_0[2]),.din(w_dff_A_pQu9YZul1_2),.clk(gclk));
	jdff dff_A_WXfcxGc05_2(.dout(w_dff_A_pQu9YZul1_2),.din(w_dff_A_WXfcxGc05_2),.clk(gclk));
	jdff dff_B_YXTVlwAl6_0(.din(n164),.dout(w_dff_B_YXTVlwAl6_0),.clk(gclk));
	jdff dff_A_DSxhz7Xv4_0(.dout(w_n96_0[0]),.din(w_dff_A_DSxhz7Xv4_0),.clk(gclk));
	jdff dff_A_fd6vNQtk6_0(.dout(w_dff_A_DSxhz7Xv4_0),.din(w_dff_A_fd6vNQtk6_0),.clk(gclk));
	jdff dff_A_i1fXFduF3_0(.dout(w_dff_A_fd6vNQtk6_0),.din(w_dff_A_i1fXFduF3_0),.clk(gclk));
	jdff dff_A_auBPxiDF9_1(.dout(w_G143gat_0[1]),.din(w_dff_A_auBPxiDF9_1),.clk(gclk));
	jdff dff_B_URNE08AT0_2(.din(G143gat),.dout(w_dff_B_URNE08AT0_2),.clk(gclk));
	jdff dff_B_hCGwS8mQ1_2(.din(w_dff_B_URNE08AT0_2),.dout(w_dff_B_hCGwS8mQ1_2),.clk(gclk));
	jdff dff_B_gxKLwhGZ4_2(.din(w_dff_B_hCGwS8mQ1_2),.dout(w_dff_B_gxKLwhGZ4_2),.clk(gclk));
	jdff dff_B_FlFqBa146_2(.din(w_dff_B_gxKLwhGZ4_2),.dout(w_dff_B_FlFqBa146_2),.clk(gclk));
	jdff dff_A_KpLc9riO5_0(.dout(w_G183gat_1[0]),.din(w_dff_A_KpLc9riO5_0),.clk(gclk));
	jdff dff_A_ZDoMkGcH7_0(.dout(w_dff_A_KpLc9riO5_0),.din(w_dff_A_ZDoMkGcH7_0),.clk(gclk));
	jdff dff_A_2Ofwe7XL4_0(.dout(w_dff_A_ZDoMkGcH7_0),.din(w_dff_A_2Ofwe7XL4_0),.clk(gclk));
	jdff dff_A_FXonsxuv3_0(.dout(w_dff_A_2Ofwe7XL4_0),.din(w_dff_A_FXonsxuv3_0),.clk(gclk));
	jdff dff_A_1X3uMO1W8_0(.dout(w_dff_A_FXonsxuv3_0),.din(w_dff_A_1X3uMO1W8_0),.clk(gclk));
	jdff dff_A_ITZ0XuNp3_0(.dout(w_dff_A_1X3uMO1W8_0),.din(w_dff_A_ITZ0XuNp3_0),.clk(gclk));
	jdff dff_A_914qiOEl3_0(.dout(w_dff_A_ITZ0XuNp3_0),.din(w_dff_A_914qiOEl3_0),.clk(gclk));
	jdff dff_A_jGGLLWCh5_0(.dout(w_dff_A_914qiOEl3_0),.din(w_dff_A_jGGLLWCh5_0),.clk(gclk));
	jdff dff_A_46jUHdup2_1(.dout(w_G183gat_1[1]),.din(w_dff_A_46jUHdup2_1),.clk(gclk));
	jdff dff_A_2Vjpfe6O8_1(.dout(w_dff_A_46jUHdup2_1),.din(w_dff_A_2Vjpfe6O8_1),.clk(gclk));
	jdff dff_A_O4OTqwSL0_1(.dout(w_dff_A_2Vjpfe6O8_1),.din(w_dff_A_O4OTqwSL0_1),.clk(gclk));
	jdff dff_A_5HyzhKfF7_1(.dout(w_dff_A_O4OTqwSL0_1),.din(w_dff_A_5HyzhKfF7_1),.clk(gclk));
	jdff dff_A_4M1fZEW37_2(.dout(w_G183gat_0[2]),.din(w_dff_A_4M1fZEW37_2),.clk(gclk));
	jdff dff_A_4hyzWsZI6_2(.dout(w_dff_A_4M1fZEW37_2),.din(w_dff_A_4hyzWsZI6_2),.clk(gclk));
	jdff dff_A_Dt3WrPyW9_2(.dout(w_dff_A_4hyzWsZI6_2),.din(w_dff_A_Dt3WrPyW9_2),.clk(gclk));
	jdff dff_A_fMtRVZPj4_2(.dout(w_dff_A_Dt3WrPyW9_2),.din(w_dff_A_fMtRVZPj4_2),.clk(gclk));
	jdff dff_A_RJifzXoI1_2(.dout(w_dff_A_fMtRVZPj4_2),.din(w_dff_A_RJifzXoI1_2),.clk(gclk));
	jdff dff_A_oVk6XzCn2_2(.dout(w_dff_A_RJifzXoI1_2),.din(w_dff_A_oVk6XzCn2_2),.clk(gclk));
	jdff dff_A_wNamG5Jj6_2(.dout(w_dff_A_oVk6XzCn2_2),.din(w_dff_A_wNamG5Jj6_2),.clk(gclk));
	jdff dff_A_yNv5bI6Q9_2(.dout(w_dff_A_wNamG5Jj6_2),.din(w_dff_A_yNv5bI6Q9_2),.clk(gclk));
	jdff dff_A_ZqyevI922_0(.dout(w_n335_0[0]),.din(w_dff_A_ZqyevI922_0),.clk(gclk));
	jdff dff_A_k2fe3CQF4_0(.dout(w_dff_A_ZqyevI922_0),.din(w_dff_A_k2fe3CQF4_0),.clk(gclk));
	jdff dff_A_36VZNr936_0(.dout(w_dff_A_k2fe3CQF4_0),.din(w_dff_A_36VZNr936_0),.clk(gclk));
	jdff dff_A_TldeYhD49_0(.dout(w_dff_A_36VZNr936_0),.din(w_dff_A_TldeYhD49_0),.clk(gclk));
	jdff dff_A_37W5QOov8_0(.dout(w_dff_A_TldeYhD49_0),.din(w_dff_A_37W5QOov8_0),.clk(gclk));
	jdff dff_A_34NJyDMq2_0(.dout(w_dff_A_37W5QOov8_0),.din(w_dff_A_34NJyDMq2_0),.clk(gclk));
	jdff dff_A_dAWNpyVM0_0(.dout(w_dff_A_34NJyDMq2_0),.din(w_dff_A_dAWNpyVM0_0),.clk(gclk));
	jdff dff_A_rvGRHzXk8_0(.dout(w_dff_A_dAWNpyVM0_0),.din(w_dff_A_rvGRHzXk8_0),.clk(gclk));
	jdff dff_B_d0rmJPO08_0(.din(n325),.dout(w_dff_B_d0rmJPO08_0),.clk(gclk));
	jdff dff_B_lj9VG66f1_0(.din(w_dff_B_d0rmJPO08_0),.dout(w_dff_B_lj9VG66f1_0),.clk(gclk));
	jdff dff_B_6AOg5QhU1_0(.din(w_dff_B_lj9VG66f1_0),.dout(w_dff_B_6AOg5QhU1_0),.clk(gclk));
	jdff dff_A_E5PkoBVc7_0(.dout(w_G153gat_0[0]),.din(w_dff_A_E5PkoBVc7_0),.clk(gclk));
	jdff dff_A_gXaunhRy7_0(.dout(w_dff_A_E5PkoBVc7_0),.din(w_dff_A_gXaunhRy7_0),.clk(gclk));
	jdff dff_A_XNiufU1F4_0(.dout(w_dff_A_gXaunhRy7_0),.din(w_dff_A_XNiufU1F4_0),.clk(gclk));
	jdff dff_A_x4rl85sv9_0(.dout(w_dff_A_XNiufU1F4_0),.din(w_dff_A_x4rl85sv9_0),.clk(gclk));
	jdff dff_A_9ClFW5Z38_2(.dout(w_G153gat_0[2]),.din(w_dff_A_9ClFW5Z38_2),.clk(gclk));
	jdff dff_A_Ya1aMsvR2_2(.dout(w_dff_A_9ClFW5Z38_2),.din(w_dff_A_Ya1aMsvR2_2),.clk(gclk));
	jdff dff_A_h5TVYHoT7_2(.dout(w_dff_A_Ya1aMsvR2_2),.din(w_dff_A_h5TVYHoT7_2),.clk(gclk));
	jdff dff_A_gwjujEoB2_2(.dout(w_dff_A_h5TVYHoT7_2),.din(w_dff_A_gwjujEoB2_2),.clk(gclk));
	jdff dff_A_GboRYmrx5_2(.dout(w_dff_A_gwjujEoB2_2),.din(w_dff_A_GboRYmrx5_2),.clk(gclk));
	jdff dff_A_JTiRaHTM1_0(.dout(w_G106gat_0[0]),.din(w_dff_A_JTiRaHTM1_0),.clk(gclk));
	jdff dff_A_gd0sAq6F5_0(.dout(w_dff_A_JTiRaHTM1_0),.din(w_dff_A_gd0sAq6F5_0),.clk(gclk));
	jdff dff_A_guMaubLw1_0(.dout(w_dff_A_gd0sAq6F5_0),.din(w_dff_A_guMaubLw1_0),.clk(gclk));
	jdff dff_A_xzquZ7UM4_0(.dout(w_dff_A_guMaubLw1_0),.din(w_dff_A_xzquZ7UM4_0),.clk(gclk));
	jdff dff_A_Vk9D0hN00_0(.dout(w_dff_A_xzquZ7UM4_0),.din(w_dff_A_Vk9D0hN00_0),.clk(gclk));
	jdff dff_A_qNPOQFP58_1(.dout(w_G177gat_1[1]),.din(w_dff_A_qNPOQFP58_1),.clk(gclk));
	jdff dff_A_bjnGDSPe2_1(.dout(w_dff_A_qNPOQFP58_1),.din(w_dff_A_bjnGDSPe2_1),.clk(gclk));
	jdff dff_A_wjyKYs0U3_1(.dout(w_dff_A_bjnGDSPe2_1),.din(w_dff_A_wjyKYs0U3_1),.clk(gclk));
	jdff dff_A_C4m0W6bJ3_1(.dout(w_dff_A_wjyKYs0U3_1),.din(w_dff_A_C4m0W6bJ3_1),.clk(gclk));
	jdff dff_A_Q1AbWXoR0_1(.dout(w_dff_A_C4m0W6bJ3_1),.din(w_dff_A_Q1AbWXoR0_1),.clk(gclk));
	jdff dff_A_zOacub3q2_1(.dout(w_dff_A_Q1AbWXoR0_1),.din(w_dff_A_zOacub3q2_1),.clk(gclk));
	jdff dff_A_jGoQ9h4C1_1(.dout(w_dff_A_zOacub3q2_1),.din(w_dff_A_jGoQ9h4C1_1),.clk(gclk));
	jdff dff_A_hNoLYn6H2_2(.dout(w_G177gat_1[2]),.din(w_dff_A_hNoLYn6H2_2),.clk(gclk));
	jdff dff_A_NX7RPgNm3_2(.dout(w_dff_A_hNoLYn6H2_2),.din(w_dff_A_NX7RPgNm3_2),.clk(gclk));
	jdff dff_A_7ZSdWsH67_2(.dout(w_dff_A_NX7RPgNm3_2),.din(w_dff_A_7ZSdWsH67_2),.clk(gclk));
	jdff dff_A_dTZzk9vt5_2(.dout(w_dff_A_7ZSdWsH67_2),.din(w_dff_A_dTZzk9vt5_2),.clk(gclk));
	jdff dff_A_Dar61H9R8_2(.dout(w_dff_A_dTZzk9vt5_2),.din(w_dff_A_Dar61H9R8_2),.clk(gclk));
	jdff dff_A_0vDvbFg78_2(.dout(w_dff_A_Dar61H9R8_2),.din(w_dff_A_0vDvbFg78_2),.clk(gclk));
	jdff dff_A_h9WWGJRw2_2(.dout(w_dff_A_0vDvbFg78_2),.din(w_dff_A_h9WWGJRw2_2),.clk(gclk));
	jdff dff_A_lwGGzGvu8_2(.dout(w_G177gat_0[2]),.din(w_dff_A_lwGGzGvu8_2),.clk(gclk));
	jdff dff_A_4ZnhGBAl6_2(.dout(w_dff_A_lwGGzGvu8_2),.din(w_dff_A_4ZnhGBAl6_2),.clk(gclk));
	jdff dff_A_456Kl9v00_2(.dout(w_dff_A_4ZnhGBAl6_2),.din(w_dff_A_456Kl9v00_2),.clk(gclk));
	jdff dff_A_08epPKth5_2(.dout(w_dff_A_456Kl9v00_2),.din(w_dff_A_08epPKth5_2),.clk(gclk));
	jdff dff_A_vgQnunVY8_1(.dout(w_n405_0[1]),.din(w_dff_A_vgQnunVY8_1),.clk(gclk));
	jdff dff_A_1vBoSNfe5_1(.dout(w_dff_A_vgQnunVY8_1),.din(w_dff_A_1vBoSNfe5_1),.clk(gclk));
	jdff dff_A_CcRdQOYK7_1(.dout(w_dff_A_1vBoSNfe5_1),.din(w_dff_A_CcRdQOYK7_1),.clk(gclk));
	jdff dff_A_HiSFdrFZ0_1(.dout(w_dff_A_CcRdQOYK7_1),.din(w_dff_A_HiSFdrFZ0_1),.clk(gclk));
	jdff dff_A_xqDhygg53_1(.dout(w_dff_A_HiSFdrFZ0_1),.din(w_dff_A_xqDhygg53_1),.clk(gclk));
	jdff dff_A_btL9Agcb8_1(.dout(w_dff_A_xqDhygg53_1),.din(w_dff_A_btL9Agcb8_1),.clk(gclk));
	jdff dff_A_XbtpfE8j7_1(.dout(w_dff_A_btL9Agcb8_1),.din(w_dff_A_XbtpfE8j7_1),.clk(gclk));
	jdff dff_A_iH9anqzM4_1(.dout(w_dff_A_XbtpfE8j7_1),.din(w_dff_A_iH9anqzM4_1),.clk(gclk));
	jdff dff_A_HARwFZmJ1_1(.dout(w_dff_A_iH9anqzM4_1),.din(w_dff_A_HARwFZmJ1_1),.clk(gclk));
	jdff dff_B_mZPw0CLR8_0(.din(n318),.dout(w_dff_B_mZPw0CLR8_0),.clk(gclk));
	jdff dff_B_BTqafFDX7_0(.din(w_dff_B_mZPw0CLR8_0),.dout(w_dff_B_BTqafFDX7_0),.clk(gclk));
	jdff dff_B_2NlrS6577_0(.din(w_dff_B_BTqafFDX7_0),.dout(w_dff_B_2NlrS6577_0),.clk(gclk));
	jdff dff_B_XdB8JRhX9_0(.din(n295),.dout(w_dff_B_XdB8JRhX9_0),.clk(gclk));
	jdff dff_A_jk2LrdXk9_0(.dout(w_G17gat_1[0]),.din(w_dff_A_jk2LrdXk9_0),.clk(gclk));
	jdff dff_A_K71u5oYo0_2(.dout(w_G17gat_1[2]),.din(w_dff_A_K71u5oYo0_2),.clk(gclk));
	jdff dff_A_VJz64C2M0_2(.dout(w_dff_A_K71u5oYo0_2),.din(w_dff_A_VJz64C2M0_2),.clk(gclk));
	jdff dff_A_Ol41ZdeR4_2(.dout(w_dff_A_VJz64C2M0_2),.din(w_dff_A_Ol41ZdeR4_2),.clk(gclk));
	jdff dff_A_pFaqW4Nf0_0(.dout(w_G80gat_0[0]),.din(w_dff_A_pFaqW4Nf0_0),.clk(gclk));
	jdff dff_A_QtnwI8EJ5_2(.dout(w_G80gat_0[2]),.din(w_dff_A_QtnwI8EJ5_2),.clk(gclk));
	jdff dff_A_spW4h4da2_0(.dout(w_G55gat_0[0]),.din(w_dff_A_spW4h4da2_0),.clk(gclk));
	jdff dff_A_gbFP4Yft7_0(.dout(w_dff_A_spW4h4da2_0),.din(w_dff_A_gbFP4Yft7_0),.clk(gclk));
	jdff dff_A_OxXuaSf93_0(.dout(w_dff_A_gbFP4Yft7_0),.din(w_dff_A_OxXuaSf93_0),.clk(gclk));
	jdff dff_A_JJjKsZ4p2_1(.dout(w_G55gat_0[1]),.din(w_dff_A_JJjKsZ4p2_1),.clk(gclk));
	jdff dff_A_m7f1IMZA8_1(.dout(w_G149gat_0[1]),.din(w_dff_A_m7f1IMZA8_1),.clk(gclk));
	jdff dff_B_rUjrGK0s1_2(.din(G149gat),.dout(w_dff_B_rUjrGK0s1_2),.clk(gclk));
	jdff dff_B_qtDbI3Zt3_2(.din(w_dff_B_rUjrGK0s1_2),.dout(w_dff_B_qtDbI3Zt3_2),.clk(gclk));
	jdff dff_B_EToVaKBN7_2(.din(w_dff_B_qtDbI3Zt3_2),.dout(w_dff_B_EToVaKBN7_2),.clk(gclk));
	jdff dff_B_mmKJ5qqi8_2(.din(w_dff_B_EToVaKBN7_2),.dout(w_dff_B_mmKJ5qqi8_2),.clk(gclk));
	jdff dff_B_MeCVlgJM3_0(.din(n152),.dout(w_dff_B_MeCVlgJM3_0),.clk(gclk));
	jdff dff_A_3LGUGYRd9_0(.dout(w_n149_0[0]),.din(w_dff_A_3LGUGYRd9_0),.clk(gclk));
	jdff dff_A_EsLHXE3L0_0(.dout(w_dff_A_3LGUGYRd9_0),.din(w_dff_A_EsLHXE3L0_0),.clk(gclk));
	jdff dff_B_xe2q5kHB6_0(.din(n147),.dout(w_dff_B_xe2q5kHB6_0),.clk(gclk));
	jdff dff_A_XqHtVFsO4_1(.dout(w_G51gat_1[1]),.din(w_dff_A_XqHtVFsO4_1),.clk(gclk));
	jdff dff_A_W1c1TVdY3_1(.dout(w_G1gat_0[1]),.din(w_dff_A_W1c1TVdY3_1),.clk(gclk));
	jdff dff_A_9YLdQILM7_1(.dout(w_dff_A_W1c1TVdY3_1),.din(w_dff_A_9YLdQILM7_1),.clk(gclk));
	jdff dff_A_3C4k9QRd6_1(.dout(w_dff_A_9YLdQILM7_1),.din(w_dff_A_3C4k9QRd6_1),.clk(gclk));
	jdff dff_A_Dm3H6giZ3_1(.dout(w_dff_A_3C4k9QRd6_1),.din(w_dff_A_Dm3H6giZ3_1),.clk(gclk));
	jdff dff_A_qsl1bnTk2_1(.dout(w_dff_A_Dm3H6giZ3_1),.din(w_dff_A_qsl1bnTk2_1),.clk(gclk));
	jdff dff_A_Q65ouTAs2_1(.dout(w_G42gat_1[1]),.din(w_dff_A_Q65ouTAs2_1),.clk(gclk));
	jdff dff_A_SozBqppf7_1(.dout(w_G42gat_0[1]),.din(w_dff_A_SozBqppf7_1),.clk(gclk));
	jdff dff_A_lPLd9Pn27_1(.dout(w_G101gat_0[1]),.din(w_dff_A_lPLd9Pn27_1),.clk(gclk));
	jdff dff_A_7k64b6kS6_1(.dout(w_dff_A_lPLd9Pn27_1),.din(w_dff_A_7k64b6kS6_1),.clk(gclk));
	jdff dff_A_dKiqw83U8_1(.dout(w_dff_A_7k64b6kS6_1),.din(w_dff_A_dKiqw83U8_1),.clk(gclk));
	jdff dff_A_hW804BSL3_1(.dout(w_dff_A_dKiqw83U8_1),.din(w_dff_A_hW804BSL3_1),.clk(gclk));
	jdff dff_A_eI78CFqv4_1(.dout(w_dff_A_hW804BSL3_1),.din(w_dff_A_eI78CFqv4_1),.clk(gclk));
	jdff dff_A_3QYhKI754_1(.dout(w_G171gat_1[1]),.din(w_dff_A_3QYhKI754_1),.clk(gclk));
	jdff dff_A_3QvyCeFi8_1(.dout(w_dff_A_3QYhKI754_1),.din(w_dff_A_3QvyCeFi8_1),.clk(gclk));
	jdff dff_A_CemPURmK5_1(.dout(w_dff_A_3QvyCeFi8_1),.din(w_dff_A_CemPURmK5_1),.clk(gclk));
	jdff dff_A_eXwJdX2V7_1(.dout(w_dff_A_CemPURmK5_1),.din(w_dff_A_eXwJdX2V7_1),.clk(gclk));
	jdff dff_A_mNaXwtfb0_1(.dout(w_dff_A_eXwJdX2V7_1),.din(w_dff_A_mNaXwtfb0_1),.clk(gclk));
	jdff dff_A_jfCAJBeO5_1(.dout(w_dff_A_mNaXwtfb0_1),.din(w_dff_A_jfCAJBeO5_1),.clk(gclk));
	jdff dff_A_y1U3RlEq9_1(.dout(w_dff_A_jfCAJBeO5_1),.din(w_dff_A_y1U3RlEq9_1),.clk(gclk));
	jdff dff_A_tS7ni6pF2_2(.dout(w_G171gat_1[2]),.din(w_dff_A_tS7ni6pF2_2),.clk(gclk));
	jdff dff_A_sHcYbj7c1_2(.dout(w_dff_A_tS7ni6pF2_2),.din(w_dff_A_sHcYbj7c1_2),.clk(gclk));
	jdff dff_A_YaR9Amxy9_2(.dout(w_dff_A_sHcYbj7c1_2),.din(w_dff_A_YaR9Amxy9_2),.clk(gclk));
	jdff dff_A_oS1obBMh2_2(.dout(w_dff_A_YaR9Amxy9_2),.din(w_dff_A_oS1obBMh2_2),.clk(gclk));
	jdff dff_A_Am7Ml6aC2_2(.dout(w_dff_A_oS1obBMh2_2),.din(w_dff_A_Am7Ml6aC2_2),.clk(gclk));
	jdff dff_A_lnV5gdjH3_2(.dout(w_dff_A_Am7Ml6aC2_2),.din(w_dff_A_lnV5gdjH3_2),.clk(gclk));
	jdff dff_A_OMzKAEPm8_2(.dout(w_dff_A_lnV5gdjH3_2),.din(w_dff_A_OMzKAEPm8_2),.clk(gclk));
	jdff dff_A_k6jXxjeM9_2(.dout(w_G171gat_0[2]),.din(w_dff_A_k6jXxjeM9_2),.clk(gclk));
	jdff dff_A_vNKgmZij1_2(.dout(w_dff_A_k6jXxjeM9_2),.din(w_dff_A_vNKgmZij1_2),.clk(gclk));
	jdff dff_A_CLRnVBti7_2(.dout(w_dff_A_vNKgmZij1_2),.din(w_dff_A_CLRnVBti7_2),.clk(gclk));
	jdff dff_A_W5CMpLB79_2(.dout(w_dff_A_CLRnVBti7_2),.din(w_dff_A_W5CMpLB79_2),.clk(gclk));
	jdff dff_A_v0x2Em3E2_2(.dout(w_dff_A_xtkQUYuL6_0),.din(w_dff_A_v0x2Em3E2_2),.clk(gclk));
	jdff dff_A_xtkQUYuL6_0(.dout(w_dff_A_KdmmqOod6_0),.din(w_dff_A_xtkQUYuL6_0),.clk(gclk));
	jdff dff_A_KdmmqOod6_0(.dout(w_dff_A_lmLj9Lys5_0),.din(w_dff_A_KdmmqOod6_0),.clk(gclk));
	jdff dff_A_lmLj9Lys5_0(.dout(w_dff_A_hDrs1Hc01_0),.din(w_dff_A_lmLj9Lys5_0),.clk(gclk));
	jdff dff_A_hDrs1Hc01_0(.dout(w_dff_A_WnumbqER2_0),.din(w_dff_A_hDrs1Hc01_0),.clk(gclk));
	jdff dff_A_WnumbqER2_0(.dout(w_dff_A_ladQDdBe3_0),.din(w_dff_A_WnumbqER2_0),.clk(gclk));
	jdff dff_A_ladQDdBe3_0(.dout(w_dff_A_xG3u0NB46_0),.din(w_dff_A_ladQDdBe3_0),.clk(gclk));
	jdff dff_A_xG3u0NB46_0(.dout(w_dff_A_DUrS3OY56_0),.din(w_dff_A_xG3u0NB46_0),.clk(gclk));
	jdff dff_A_DUrS3OY56_0(.dout(w_dff_A_89cFRmeR0_0),.din(w_dff_A_DUrS3OY56_0),.clk(gclk));
	jdff dff_A_89cFRmeR0_0(.dout(w_dff_A_J3g2x2e91_0),.din(w_dff_A_89cFRmeR0_0),.clk(gclk));
	jdff dff_A_J3g2x2e91_0(.dout(w_dff_A_DQsXNwKp4_0),.din(w_dff_A_J3g2x2e91_0),.clk(gclk));
	jdff dff_A_DQsXNwKp4_0(.dout(w_dff_A_liEfg0Qt9_0),.din(w_dff_A_DQsXNwKp4_0),.clk(gclk));
	jdff dff_A_liEfg0Qt9_0(.dout(w_dff_A_DGHc9F6a3_0),.din(w_dff_A_liEfg0Qt9_0),.clk(gclk));
	jdff dff_A_DGHc9F6a3_0(.dout(w_dff_A_SJjSEmZ87_0),.din(w_dff_A_DGHc9F6a3_0),.clk(gclk));
	jdff dff_A_SJjSEmZ87_0(.dout(w_dff_A_9t8R4aYe8_0),.din(w_dff_A_SJjSEmZ87_0),.clk(gclk));
	jdff dff_A_9t8R4aYe8_0(.dout(w_dff_A_DJVy1Vj43_0),.din(w_dff_A_9t8R4aYe8_0),.clk(gclk));
	jdff dff_A_DJVy1Vj43_0(.dout(w_dff_A_P4z0Z6u07_0),.din(w_dff_A_DJVy1Vj43_0),.clk(gclk));
	jdff dff_A_P4z0Z6u07_0(.dout(w_dff_A_JFbBJjwL8_0),.din(w_dff_A_P4z0Z6u07_0),.clk(gclk));
	jdff dff_A_JFbBJjwL8_0(.dout(G388gat),.din(w_dff_A_JFbBJjwL8_0),.clk(gclk));
	jdff dff_A_2Vs49HL71_2(.dout(w_dff_A_Zvluu8NA5_0),.din(w_dff_A_2Vs49HL71_2),.clk(gclk));
	jdff dff_A_Zvluu8NA5_0(.dout(w_dff_A_vfa2d84t6_0),.din(w_dff_A_Zvluu8NA5_0),.clk(gclk));
	jdff dff_A_vfa2d84t6_0(.dout(w_dff_A_9n1AUUg50_0),.din(w_dff_A_vfa2d84t6_0),.clk(gclk));
	jdff dff_A_9n1AUUg50_0(.dout(w_dff_A_xDP9o8427_0),.din(w_dff_A_9n1AUUg50_0),.clk(gclk));
	jdff dff_A_xDP9o8427_0(.dout(w_dff_A_mXAxSiCI5_0),.din(w_dff_A_xDP9o8427_0),.clk(gclk));
	jdff dff_A_mXAxSiCI5_0(.dout(w_dff_A_f0lOnMoU3_0),.din(w_dff_A_mXAxSiCI5_0),.clk(gclk));
	jdff dff_A_f0lOnMoU3_0(.dout(w_dff_A_n8OxAATE0_0),.din(w_dff_A_f0lOnMoU3_0),.clk(gclk));
	jdff dff_A_n8OxAATE0_0(.dout(w_dff_A_jCUKFyHl9_0),.din(w_dff_A_n8OxAATE0_0),.clk(gclk));
	jdff dff_A_jCUKFyHl9_0(.dout(w_dff_A_0aUvTdKl0_0),.din(w_dff_A_jCUKFyHl9_0),.clk(gclk));
	jdff dff_A_0aUvTdKl0_0(.dout(w_dff_A_rQd0gKmE4_0),.din(w_dff_A_0aUvTdKl0_0),.clk(gclk));
	jdff dff_A_rQd0gKmE4_0(.dout(w_dff_A_G6W5veAp4_0),.din(w_dff_A_rQd0gKmE4_0),.clk(gclk));
	jdff dff_A_G6W5veAp4_0(.dout(w_dff_A_MkuOaLul8_0),.din(w_dff_A_G6W5veAp4_0),.clk(gclk));
	jdff dff_A_MkuOaLul8_0(.dout(w_dff_A_7bMKgShr7_0),.din(w_dff_A_MkuOaLul8_0),.clk(gclk));
	jdff dff_A_7bMKgShr7_0(.dout(w_dff_A_hPT0rcx76_0),.din(w_dff_A_7bMKgShr7_0),.clk(gclk));
	jdff dff_A_hPT0rcx76_0(.dout(w_dff_A_aqE72HcN8_0),.din(w_dff_A_hPT0rcx76_0),.clk(gclk));
	jdff dff_A_aqE72HcN8_0(.dout(w_dff_A_WManN0r55_0),.din(w_dff_A_aqE72HcN8_0),.clk(gclk));
	jdff dff_A_WManN0r55_0(.dout(w_dff_A_4cToR0fG3_0),.din(w_dff_A_WManN0r55_0),.clk(gclk));
	jdff dff_A_4cToR0fG3_0(.dout(w_dff_A_hft1OadK4_0),.din(w_dff_A_4cToR0fG3_0),.clk(gclk));
	jdff dff_A_hft1OadK4_0(.dout(G389gat),.din(w_dff_A_hft1OadK4_0),.clk(gclk));
	jdff dff_A_CX6SNnSY4_2(.dout(w_dff_A_E4w2Cg7B7_0),.din(w_dff_A_CX6SNnSY4_2),.clk(gclk));
	jdff dff_A_E4w2Cg7B7_0(.dout(w_dff_A_sJiKNRuu5_0),.din(w_dff_A_E4w2Cg7B7_0),.clk(gclk));
	jdff dff_A_sJiKNRuu5_0(.dout(w_dff_A_LYXWeyiV4_0),.din(w_dff_A_sJiKNRuu5_0),.clk(gclk));
	jdff dff_A_LYXWeyiV4_0(.dout(w_dff_A_IVzQps155_0),.din(w_dff_A_LYXWeyiV4_0),.clk(gclk));
	jdff dff_A_IVzQps155_0(.dout(w_dff_A_XYs2lv1G6_0),.din(w_dff_A_IVzQps155_0),.clk(gclk));
	jdff dff_A_XYs2lv1G6_0(.dout(w_dff_A_lsVcQylp4_0),.din(w_dff_A_XYs2lv1G6_0),.clk(gclk));
	jdff dff_A_lsVcQylp4_0(.dout(w_dff_A_nriLEvHh8_0),.din(w_dff_A_lsVcQylp4_0),.clk(gclk));
	jdff dff_A_nriLEvHh8_0(.dout(w_dff_A_iymqAfR47_0),.din(w_dff_A_nriLEvHh8_0),.clk(gclk));
	jdff dff_A_iymqAfR47_0(.dout(w_dff_A_RGoTqBv61_0),.din(w_dff_A_iymqAfR47_0),.clk(gclk));
	jdff dff_A_RGoTqBv61_0(.dout(w_dff_A_9wsH7zyo4_0),.din(w_dff_A_RGoTqBv61_0),.clk(gclk));
	jdff dff_A_9wsH7zyo4_0(.dout(w_dff_A_J8nQqiQK1_0),.din(w_dff_A_9wsH7zyo4_0),.clk(gclk));
	jdff dff_A_J8nQqiQK1_0(.dout(w_dff_A_AuJeQc7Z9_0),.din(w_dff_A_J8nQqiQK1_0),.clk(gclk));
	jdff dff_A_AuJeQc7Z9_0(.dout(w_dff_A_9trUj2dj2_0),.din(w_dff_A_AuJeQc7Z9_0),.clk(gclk));
	jdff dff_A_9trUj2dj2_0(.dout(w_dff_A_ZYTG7bga4_0),.din(w_dff_A_9trUj2dj2_0),.clk(gclk));
	jdff dff_A_ZYTG7bga4_0(.dout(w_dff_A_VkeoxyuL1_0),.din(w_dff_A_ZYTG7bga4_0),.clk(gclk));
	jdff dff_A_VkeoxyuL1_0(.dout(w_dff_A_E1YH34Hz8_0),.din(w_dff_A_VkeoxyuL1_0),.clk(gclk));
	jdff dff_A_E1YH34Hz8_0(.dout(w_dff_A_rT324FG03_0),.din(w_dff_A_E1YH34Hz8_0),.clk(gclk));
	jdff dff_A_rT324FG03_0(.dout(w_dff_A_iUxU1lmx4_0),.din(w_dff_A_rT324FG03_0),.clk(gclk));
	jdff dff_A_iUxU1lmx4_0(.dout(G390gat),.din(w_dff_A_iUxU1lmx4_0),.clk(gclk));
	jdff dff_A_Xh2ELakS9_2(.dout(w_dff_A_RcxGboRk1_0),.din(w_dff_A_Xh2ELakS9_2),.clk(gclk));
	jdff dff_A_RcxGboRk1_0(.dout(w_dff_A_wYF4a9w83_0),.din(w_dff_A_RcxGboRk1_0),.clk(gclk));
	jdff dff_A_wYF4a9w83_0(.dout(w_dff_A_JHzzZ78h0_0),.din(w_dff_A_wYF4a9w83_0),.clk(gclk));
	jdff dff_A_JHzzZ78h0_0(.dout(w_dff_A_uSIQMkia0_0),.din(w_dff_A_JHzzZ78h0_0),.clk(gclk));
	jdff dff_A_uSIQMkia0_0(.dout(w_dff_A_PrbXm2LQ2_0),.din(w_dff_A_uSIQMkia0_0),.clk(gclk));
	jdff dff_A_PrbXm2LQ2_0(.dout(w_dff_A_ivyqjlCB7_0),.din(w_dff_A_PrbXm2LQ2_0),.clk(gclk));
	jdff dff_A_ivyqjlCB7_0(.dout(w_dff_A_U2ptytqh7_0),.din(w_dff_A_ivyqjlCB7_0),.clk(gclk));
	jdff dff_A_U2ptytqh7_0(.dout(w_dff_A_xEV7E2Dx5_0),.din(w_dff_A_U2ptytqh7_0),.clk(gclk));
	jdff dff_A_xEV7E2Dx5_0(.dout(w_dff_A_pECFW0EF4_0),.din(w_dff_A_xEV7E2Dx5_0),.clk(gclk));
	jdff dff_A_pECFW0EF4_0(.dout(w_dff_A_nMDLpxkd2_0),.din(w_dff_A_pECFW0EF4_0),.clk(gclk));
	jdff dff_A_nMDLpxkd2_0(.dout(w_dff_A_HTPJ8ZFe9_0),.din(w_dff_A_nMDLpxkd2_0),.clk(gclk));
	jdff dff_A_HTPJ8ZFe9_0(.dout(w_dff_A_hJzaNZo99_0),.din(w_dff_A_HTPJ8ZFe9_0),.clk(gclk));
	jdff dff_A_hJzaNZo99_0(.dout(w_dff_A_XA9uKdIl9_0),.din(w_dff_A_hJzaNZo99_0),.clk(gclk));
	jdff dff_A_XA9uKdIl9_0(.dout(w_dff_A_WCkSSlC85_0),.din(w_dff_A_XA9uKdIl9_0),.clk(gclk));
	jdff dff_A_WCkSSlC85_0(.dout(w_dff_A_WbkkA9fY0_0),.din(w_dff_A_WCkSSlC85_0),.clk(gclk));
	jdff dff_A_WbkkA9fY0_0(.dout(w_dff_A_u7QlEQN13_0),.din(w_dff_A_WbkkA9fY0_0),.clk(gclk));
	jdff dff_A_u7QlEQN13_0(.dout(w_dff_A_WReXI3mr5_0),.din(w_dff_A_u7QlEQN13_0),.clk(gclk));
	jdff dff_A_WReXI3mr5_0(.dout(w_dff_A_GBtaoWwc3_0),.din(w_dff_A_WReXI3mr5_0),.clk(gclk));
	jdff dff_A_GBtaoWwc3_0(.dout(w_dff_A_itv1kqrl8_0),.din(w_dff_A_GBtaoWwc3_0),.clk(gclk));
	jdff dff_A_itv1kqrl8_0(.dout(G391gat),.din(w_dff_A_itv1kqrl8_0),.clk(gclk));
	jdff dff_A_FDWFIrl16_2(.dout(w_dff_A_D5WWLe269_0),.din(w_dff_A_FDWFIrl16_2),.clk(gclk));
	jdff dff_A_D5WWLe269_0(.dout(w_dff_A_D1ILTAvo4_0),.din(w_dff_A_D5WWLe269_0),.clk(gclk));
	jdff dff_A_D1ILTAvo4_0(.dout(w_dff_A_3K0vDBkf2_0),.din(w_dff_A_D1ILTAvo4_0),.clk(gclk));
	jdff dff_A_3K0vDBkf2_0(.dout(w_dff_A_5kUjCC0O9_0),.din(w_dff_A_3K0vDBkf2_0),.clk(gclk));
	jdff dff_A_5kUjCC0O9_0(.dout(w_dff_A_ows4u9JO5_0),.din(w_dff_A_5kUjCC0O9_0),.clk(gclk));
	jdff dff_A_ows4u9JO5_0(.dout(w_dff_A_uVPYN4iP4_0),.din(w_dff_A_ows4u9JO5_0),.clk(gclk));
	jdff dff_A_uVPYN4iP4_0(.dout(w_dff_A_kzKSYTzO7_0),.din(w_dff_A_uVPYN4iP4_0),.clk(gclk));
	jdff dff_A_kzKSYTzO7_0(.dout(w_dff_A_WSNnWOHh0_0),.din(w_dff_A_kzKSYTzO7_0),.clk(gclk));
	jdff dff_A_WSNnWOHh0_0(.dout(w_dff_A_KyyocGZe6_0),.din(w_dff_A_WSNnWOHh0_0),.clk(gclk));
	jdff dff_A_KyyocGZe6_0(.dout(w_dff_A_THNrH40Q5_0),.din(w_dff_A_KyyocGZe6_0),.clk(gclk));
	jdff dff_A_THNrH40Q5_0(.dout(w_dff_A_qXSwfnKp8_0),.din(w_dff_A_THNrH40Q5_0),.clk(gclk));
	jdff dff_A_qXSwfnKp8_0(.dout(w_dff_A_5XdKHzDI6_0),.din(w_dff_A_qXSwfnKp8_0),.clk(gclk));
	jdff dff_A_5XdKHzDI6_0(.dout(w_dff_A_bt9xHAmH3_0),.din(w_dff_A_5XdKHzDI6_0),.clk(gclk));
	jdff dff_A_bt9xHAmH3_0(.dout(w_dff_A_0SO10ped5_0),.din(w_dff_A_bt9xHAmH3_0),.clk(gclk));
	jdff dff_A_0SO10ped5_0(.dout(w_dff_A_0Cl95lyv3_0),.din(w_dff_A_0SO10ped5_0),.clk(gclk));
	jdff dff_A_0Cl95lyv3_0(.dout(w_dff_A_tinlgHgA4_0),.din(w_dff_A_0Cl95lyv3_0),.clk(gclk));
	jdff dff_A_tinlgHgA4_0(.dout(w_dff_A_imctwPHn3_0),.din(w_dff_A_tinlgHgA4_0),.clk(gclk));
	jdff dff_A_imctwPHn3_0(.dout(w_dff_A_QRMKaVJk5_0),.din(w_dff_A_imctwPHn3_0),.clk(gclk));
	jdff dff_A_QRMKaVJk5_0(.dout(G418gat),.din(w_dff_A_QRMKaVJk5_0),.clk(gclk));
	jdff dff_A_tqHLL7uK6_2(.dout(w_dff_A_KACSFeVn6_0),.din(w_dff_A_tqHLL7uK6_2),.clk(gclk));
	jdff dff_A_KACSFeVn6_0(.dout(w_dff_A_IJbXFV4b9_0),.din(w_dff_A_KACSFeVn6_0),.clk(gclk));
	jdff dff_A_IJbXFV4b9_0(.dout(w_dff_A_AiP1ikyE7_0),.din(w_dff_A_IJbXFV4b9_0),.clk(gclk));
	jdff dff_A_AiP1ikyE7_0(.dout(w_dff_A_tH3EmEVv1_0),.din(w_dff_A_AiP1ikyE7_0),.clk(gclk));
	jdff dff_A_tH3EmEVv1_0(.dout(w_dff_A_jTuRkaIz4_0),.din(w_dff_A_tH3EmEVv1_0),.clk(gclk));
	jdff dff_A_jTuRkaIz4_0(.dout(w_dff_A_n3cnsbSD6_0),.din(w_dff_A_jTuRkaIz4_0),.clk(gclk));
	jdff dff_A_n3cnsbSD6_0(.dout(w_dff_A_CJlwXQdA8_0),.din(w_dff_A_n3cnsbSD6_0),.clk(gclk));
	jdff dff_A_CJlwXQdA8_0(.dout(w_dff_A_3AKbhcvO5_0),.din(w_dff_A_CJlwXQdA8_0),.clk(gclk));
	jdff dff_A_3AKbhcvO5_0(.dout(w_dff_A_mJodgsau7_0),.din(w_dff_A_3AKbhcvO5_0),.clk(gclk));
	jdff dff_A_mJodgsau7_0(.dout(w_dff_A_HfTbvByc6_0),.din(w_dff_A_mJodgsau7_0),.clk(gclk));
	jdff dff_A_HfTbvByc6_0(.dout(w_dff_A_anntVTbu3_0),.din(w_dff_A_HfTbvByc6_0),.clk(gclk));
	jdff dff_A_anntVTbu3_0(.dout(w_dff_A_MMJYSJ0X6_0),.din(w_dff_A_anntVTbu3_0),.clk(gclk));
	jdff dff_A_MMJYSJ0X6_0(.dout(w_dff_A_F5vSktkQ3_0),.din(w_dff_A_MMJYSJ0X6_0),.clk(gclk));
	jdff dff_A_F5vSktkQ3_0(.dout(w_dff_A_asiu61cE3_0),.din(w_dff_A_F5vSktkQ3_0),.clk(gclk));
	jdff dff_A_asiu61cE3_0(.dout(w_dff_A_TiJ0vDt26_0),.din(w_dff_A_asiu61cE3_0),.clk(gclk));
	jdff dff_A_TiJ0vDt26_0(.dout(w_dff_A_Q9Mm0WCy1_0),.din(w_dff_A_TiJ0vDt26_0),.clk(gclk));
	jdff dff_A_Q9Mm0WCy1_0(.dout(G419gat),.din(w_dff_A_Q9Mm0WCy1_0),.clk(gclk));
	jdff dff_A_3Vj6ap9D4_2(.dout(w_dff_A_wNpyU6gF4_0),.din(w_dff_A_3Vj6ap9D4_2),.clk(gclk));
	jdff dff_A_wNpyU6gF4_0(.dout(w_dff_A_wxn9bf7a8_0),.din(w_dff_A_wNpyU6gF4_0),.clk(gclk));
	jdff dff_A_wxn9bf7a8_0(.dout(w_dff_A_T9CsQu4l1_0),.din(w_dff_A_wxn9bf7a8_0),.clk(gclk));
	jdff dff_A_T9CsQu4l1_0(.dout(w_dff_A_d5QdZfZp7_0),.din(w_dff_A_T9CsQu4l1_0),.clk(gclk));
	jdff dff_A_d5QdZfZp7_0(.dout(w_dff_A_y8Yu9Aez5_0),.din(w_dff_A_d5QdZfZp7_0),.clk(gclk));
	jdff dff_A_y8Yu9Aez5_0(.dout(w_dff_A_2EvaerIa6_0),.din(w_dff_A_y8Yu9Aez5_0),.clk(gclk));
	jdff dff_A_2EvaerIa6_0(.dout(w_dff_A_CjJUkOXJ7_0),.din(w_dff_A_2EvaerIa6_0),.clk(gclk));
	jdff dff_A_CjJUkOXJ7_0(.dout(w_dff_A_FOww7t603_0),.din(w_dff_A_CjJUkOXJ7_0),.clk(gclk));
	jdff dff_A_FOww7t603_0(.dout(w_dff_A_X2QbrQik8_0),.din(w_dff_A_FOww7t603_0),.clk(gclk));
	jdff dff_A_X2QbrQik8_0(.dout(w_dff_A_25avs1oa0_0),.din(w_dff_A_X2QbrQik8_0),.clk(gclk));
	jdff dff_A_25avs1oa0_0(.dout(w_dff_A_tecoaT1k6_0),.din(w_dff_A_25avs1oa0_0),.clk(gclk));
	jdff dff_A_tecoaT1k6_0(.dout(w_dff_A_4UgBqPiN4_0),.din(w_dff_A_tecoaT1k6_0),.clk(gclk));
	jdff dff_A_4UgBqPiN4_0(.dout(w_dff_A_kfZWxZa49_0),.din(w_dff_A_4UgBqPiN4_0),.clk(gclk));
	jdff dff_A_kfZWxZa49_0(.dout(w_dff_A_a5YZHejn2_0),.din(w_dff_A_kfZWxZa49_0),.clk(gclk));
	jdff dff_A_a5YZHejn2_0(.dout(w_dff_A_eyzhNh3I2_0),.din(w_dff_A_a5YZHejn2_0),.clk(gclk));
	jdff dff_A_eyzhNh3I2_0(.dout(w_dff_A_IaD2PxtD0_0),.din(w_dff_A_eyzhNh3I2_0),.clk(gclk));
	jdff dff_A_IaD2PxtD0_0(.dout(w_dff_A_kZ9MkF7H9_0),.din(w_dff_A_IaD2PxtD0_0),.clk(gclk));
	jdff dff_A_kZ9MkF7H9_0(.dout(G420gat),.din(w_dff_A_kZ9MkF7H9_0),.clk(gclk));
	jdff dff_A_XFUZnNOl3_2(.dout(w_dff_A_rPTjTisk5_0),.din(w_dff_A_XFUZnNOl3_2),.clk(gclk));
	jdff dff_A_rPTjTisk5_0(.dout(w_dff_A_p5xzbR8Z7_0),.din(w_dff_A_rPTjTisk5_0),.clk(gclk));
	jdff dff_A_p5xzbR8Z7_0(.dout(w_dff_A_XNugZ0bg6_0),.din(w_dff_A_p5xzbR8Z7_0),.clk(gclk));
	jdff dff_A_XNugZ0bg6_0(.dout(w_dff_A_3q1Aja3K1_0),.din(w_dff_A_XNugZ0bg6_0),.clk(gclk));
	jdff dff_A_3q1Aja3K1_0(.dout(w_dff_A_UrIQz1AP4_0),.din(w_dff_A_3q1Aja3K1_0),.clk(gclk));
	jdff dff_A_UrIQz1AP4_0(.dout(w_dff_A_du7xO8RR3_0),.din(w_dff_A_UrIQz1AP4_0),.clk(gclk));
	jdff dff_A_du7xO8RR3_0(.dout(w_dff_A_kjdfwjxG3_0),.din(w_dff_A_du7xO8RR3_0),.clk(gclk));
	jdff dff_A_kjdfwjxG3_0(.dout(w_dff_A_9AXVyoWV3_0),.din(w_dff_A_kjdfwjxG3_0),.clk(gclk));
	jdff dff_A_9AXVyoWV3_0(.dout(w_dff_A_X0u2I49y7_0),.din(w_dff_A_9AXVyoWV3_0),.clk(gclk));
	jdff dff_A_X0u2I49y7_0(.dout(w_dff_A_6tq8lMEF6_0),.din(w_dff_A_X0u2I49y7_0),.clk(gclk));
	jdff dff_A_6tq8lMEF6_0(.dout(w_dff_A_6SniNiZx7_0),.din(w_dff_A_6tq8lMEF6_0),.clk(gclk));
	jdff dff_A_6SniNiZx7_0(.dout(w_dff_A_lxLJ1r8X9_0),.din(w_dff_A_6SniNiZx7_0),.clk(gclk));
	jdff dff_A_lxLJ1r8X9_0(.dout(w_dff_A_PpOKEoAJ1_0),.din(w_dff_A_lxLJ1r8X9_0),.clk(gclk));
	jdff dff_A_PpOKEoAJ1_0(.dout(w_dff_A_P1ybqFjO2_0),.din(w_dff_A_PpOKEoAJ1_0),.clk(gclk));
	jdff dff_A_P1ybqFjO2_0(.dout(w_dff_A_4zWGkNDC0_0),.din(w_dff_A_P1ybqFjO2_0),.clk(gclk));
	jdff dff_A_4zWGkNDC0_0(.dout(w_dff_A_fvTmgAWN7_0),.din(w_dff_A_4zWGkNDC0_0),.clk(gclk));
	jdff dff_A_fvTmgAWN7_0(.dout(w_dff_A_ODiXCupA7_0),.din(w_dff_A_fvTmgAWN7_0),.clk(gclk));
	jdff dff_A_ODiXCupA7_0(.dout(G421gat),.din(w_dff_A_ODiXCupA7_0),.clk(gclk));
	jdff dff_A_g6bXiTJg5_2(.dout(w_dff_A_mcPsRd1K9_0),.din(w_dff_A_g6bXiTJg5_2),.clk(gclk));
	jdff dff_A_mcPsRd1K9_0(.dout(w_dff_A_hN4nzfMg3_0),.din(w_dff_A_mcPsRd1K9_0),.clk(gclk));
	jdff dff_A_hN4nzfMg3_0(.dout(w_dff_A_wfoY278h7_0),.din(w_dff_A_hN4nzfMg3_0),.clk(gclk));
	jdff dff_A_wfoY278h7_0(.dout(w_dff_A_axWIUTCu1_0),.din(w_dff_A_wfoY278h7_0),.clk(gclk));
	jdff dff_A_axWIUTCu1_0(.dout(w_dff_A_xZA8gvVV4_0),.din(w_dff_A_axWIUTCu1_0),.clk(gclk));
	jdff dff_A_xZA8gvVV4_0(.dout(w_dff_A_0ex4AtiZ6_0),.din(w_dff_A_xZA8gvVV4_0),.clk(gclk));
	jdff dff_A_0ex4AtiZ6_0(.dout(w_dff_A_oaK77J3U7_0),.din(w_dff_A_0ex4AtiZ6_0),.clk(gclk));
	jdff dff_A_oaK77J3U7_0(.dout(w_dff_A_Ibf4GOqP4_0),.din(w_dff_A_oaK77J3U7_0),.clk(gclk));
	jdff dff_A_Ibf4GOqP4_0(.dout(w_dff_A_y82YZVhN4_0),.din(w_dff_A_Ibf4GOqP4_0),.clk(gclk));
	jdff dff_A_y82YZVhN4_0(.dout(w_dff_A_sCzAckFO8_0),.din(w_dff_A_y82YZVhN4_0),.clk(gclk));
	jdff dff_A_sCzAckFO8_0(.dout(w_dff_A_c82g1weT7_0),.din(w_dff_A_sCzAckFO8_0),.clk(gclk));
	jdff dff_A_c82g1weT7_0(.dout(w_dff_A_Ucp7WZ6P4_0),.din(w_dff_A_c82g1weT7_0),.clk(gclk));
	jdff dff_A_Ucp7WZ6P4_0(.dout(w_dff_A_kw1IApWj5_0),.din(w_dff_A_Ucp7WZ6P4_0),.clk(gclk));
	jdff dff_A_kw1IApWj5_0(.dout(w_dff_A_RLRdFeb08_0),.din(w_dff_A_kw1IApWj5_0),.clk(gclk));
	jdff dff_A_RLRdFeb08_0(.dout(w_dff_A_aQ99LbxA2_0),.din(w_dff_A_RLRdFeb08_0),.clk(gclk));
	jdff dff_A_aQ99LbxA2_0(.dout(w_dff_A_eM4weOKO9_0),.din(w_dff_A_aQ99LbxA2_0),.clk(gclk));
	jdff dff_A_eM4weOKO9_0(.dout(w_dff_A_2Z61ps791_0),.din(w_dff_A_eM4weOKO9_0),.clk(gclk));
	jdff dff_A_2Z61ps791_0(.dout(G422gat),.din(w_dff_A_2Z61ps791_0),.clk(gclk));
	jdff dff_A_2F8BBGCp1_2(.dout(w_dff_A_8ab2RlK79_0),.din(w_dff_A_2F8BBGCp1_2),.clk(gclk));
	jdff dff_A_8ab2RlK79_0(.dout(w_dff_A_hE6bpMsx8_0),.din(w_dff_A_8ab2RlK79_0),.clk(gclk));
	jdff dff_A_hE6bpMsx8_0(.dout(w_dff_A_h5cCdXKr6_0),.din(w_dff_A_hE6bpMsx8_0),.clk(gclk));
	jdff dff_A_h5cCdXKr6_0(.dout(w_dff_A_nWQERbPz9_0),.din(w_dff_A_h5cCdXKr6_0),.clk(gclk));
	jdff dff_A_nWQERbPz9_0(.dout(w_dff_A_IpZ0lVAO4_0),.din(w_dff_A_nWQERbPz9_0),.clk(gclk));
	jdff dff_A_IpZ0lVAO4_0(.dout(w_dff_A_tW4eTduQ6_0),.din(w_dff_A_IpZ0lVAO4_0),.clk(gclk));
	jdff dff_A_tW4eTduQ6_0(.dout(w_dff_A_AVG8HZr79_0),.din(w_dff_A_tW4eTduQ6_0),.clk(gclk));
	jdff dff_A_AVG8HZr79_0(.dout(w_dff_A_D65CF86p1_0),.din(w_dff_A_AVG8HZr79_0),.clk(gclk));
	jdff dff_A_D65CF86p1_0(.dout(w_dff_A_oJTu87Dn6_0),.din(w_dff_A_D65CF86p1_0),.clk(gclk));
	jdff dff_A_oJTu87Dn6_0(.dout(w_dff_A_8Xr1gNFM8_0),.din(w_dff_A_oJTu87Dn6_0),.clk(gclk));
	jdff dff_A_8Xr1gNFM8_0(.dout(w_dff_A_tHBMkvBX5_0),.din(w_dff_A_8Xr1gNFM8_0),.clk(gclk));
	jdff dff_A_tHBMkvBX5_0(.dout(w_dff_A_ALvt2Tr15_0),.din(w_dff_A_tHBMkvBX5_0),.clk(gclk));
	jdff dff_A_ALvt2Tr15_0(.dout(w_dff_A_4bYeS8tP7_0),.din(w_dff_A_ALvt2Tr15_0),.clk(gclk));
	jdff dff_A_4bYeS8tP7_0(.dout(w_dff_A_AZUh64Lp7_0),.din(w_dff_A_4bYeS8tP7_0),.clk(gclk));
	jdff dff_A_AZUh64Lp7_0(.dout(w_dff_A_WFk6BzR51_0),.din(w_dff_A_AZUh64Lp7_0),.clk(gclk));
	jdff dff_A_WFk6BzR51_0(.dout(w_dff_A_ZRHcwRTJ9_0),.din(w_dff_A_WFk6BzR51_0),.clk(gclk));
	jdff dff_A_ZRHcwRTJ9_0(.dout(w_dff_A_YZvl8Xfh8_0),.din(w_dff_A_ZRHcwRTJ9_0),.clk(gclk));
	jdff dff_A_YZvl8Xfh8_0(.dout(w_dff_A_Jy0JyhUZ8_0),.din(w_dff_A_YZvl8Xfh8_0),.clk(gclk));
	jdff dff_A_Jy0JyhUZ8_0(.dout(G423gat),.din(w_dff_A_Jy0JyhUZ8_0),.clk(gclk));
	jdff dff_A_NowZgrpN0_2(.dout(w_dff_A_ez5JPiF32_0),.din(w_dff_A_NowZgrpN0_2),.clk(gclk));
	jdff dff_A_ez5JPiF32_0(.dout(w_dff_A_aJhmc3KS9_0),.din(w_dff_A_ez5JPiF32_0),.clk(gclk));
	jdff dff_A_aJhmc3KS9_0(.dout(w_dff_A_Mqbvvkrg6_0),.din(w_dff_A_aJhmc3KS9_0),.clk(gclk));
	jdff dff_A_Mqbvvkrg6_0(.dout(w_dff_A_ua8wzgOT2_0),.din(w_dff_A_Mqbvvkrg6_0),.clk(gclk));
	jdff dff_A_ua8wzgOT2_0(.dout(w_dff_A_y8GMdNal9_0),.din(w_dff_A_ua8wzgOT2_0),.clk(gclk));
	jdff dff_A_y8GMdNal9_0(.dout(w_dff_A_7abAmPvm7_0),.din(w_dff_A_y8GMdNal9_0),.clk(gclk));
	jdff dff_A_7abAmPvm7_0(.dout(w_dff_A_vRKz4I905_0),.din(w_dff_A_7abAmPvm7_0),.clk(gclk));
	jdff dff_A_vRKz4I905_0(.dout(w_dff_A_hJ98fB685_0),.din(w_dff_A_vRKz4I905_0),.clk(gclk));
	jdff dff_A_hJ98fB685_0(.dout(w_dff_A_ps25jzSs5_0),.din(w_dff_A_hJ98fB685_0),.clk(gclk));
	jdff dff_A_ps25jzSs5_0(.dout(w_dff_A_Xe6d9Sok1_0),.din(w_dff_A_ps25jzSs5_0),.clk(gclk));
	jdff dff_A_Xe6d9Sok1_0(.dout(w_dff_A_mQzREqH25_0),.din(w_dff_A_Xe6d9Sok1_0),.clk(gclk));
	jdff dff_A_mQzREqH25_0(.dout(w_dff_A_V9ltStEh0_0),.din(w_dff_A_mQzREqH25_0),.clk(gclk));
	jdff dff_A_V9ltStEh0_0(.dout(w_dff_A_hMqEYEQA0_0),.din(w_dff_A_V9ltStEh0_0),.clk(gclk));
	jdff dff_A_hMqEYEQA0_0(.dout(w_dff_A_zhbMisoT8_0),.din(w_dff_A_hMqEYEQA0_0),.clk(gclk));
	jdff dff_A_zhbMisoT8_0(.dout(w_dff_A_BMLBQxe45_0),.din(w_dff_A_zhbMisoT8_0),.clk(gclk));
	jdff dff_A_BMLBQxe45_0(.dout(w_dff_A_0R5U5ofJ9_0),.din(w_dff_A_BMLBQxe45_0),.clk(gclk));
	jdff dff_A_0R5U5ofJ9_0(.dout(G446gat),.din(w_dff_A_0R5U5ofJ9_0),.clk(gclk));
	jdff dff_A_wbw40VA04_1(.dout(w_dff_A_RWWMBmUX0_0),.din(w_dff_A_wbw40VA04_1),.clk(gclk));
	jdff dff_A_RWWMBmUX0_0(.dout(w_dff_A_Y9HYAg1j0_0),.din(w_dff_A_RWWMBmUX0_0),.clk(gclk));
	jdff dff_A_Y9HYAg1j0_0(.dout(w_dff_A_pFwygKjG0_0),.din(w_dff_A_Y9HYAg1j0_0),.clk(gclk));
	jdff dff_A_pFwygKjG0_0(.dout(w_dff_A_XQlQGsfQ8_0),.din(w_dff_A_pFwygKjG0_0),.clk(gclk));
	jdff dff_A_XQlQGsfQ8_0(.dout(w_dff_A_NtPzn7Qf6_0),.din(w_dff_A_XQlQGsfQ8_0),.clk(gclk));
	jdff dff_A_NtPzn7Qf6_0(.dout(w_dff_A_JseRuWVB6_0),.din(w_dff_A_NtPzn7Qf6_0),.clk(gclk));
	jdff dff_A_JseRuWVB6_0(.dout(w_dff_A_LNObQEut7_0),.din(w_dff_A_JseRuWVB6_0),.clk(gclk));
	jdff dff_A_LNObQEut7_0(.dout(w_dff_A_ncz4YBQL5_0),.din(w_dff_A_LNObQEut7_0),.clk(gclk));
	jdff dff_A_ncz4YBQL5_0(.dout(w_dff_A_VYVtXc3e4_0),.din(w_dff_A_ncz4YBQL5_0),.clk(gclk));
	jdff dff_A_VYVtXc3e4_0(.dout(w_dff_A_X8vKrcpy5_0),.din(w_dff_A_VYVtXc3e4_0),.clk(gclk));
	jdff dff_A_X8vKrcpy5_0(.dout(w_dff_A_V4wPDe5y5_0),.din(w_dff_A_X8vKrcpy5_0),.clk(gclk));
	jdff dff_A_V4wPDe5y5_0(.dout(w_dff_A_c0InGZ4f6_0),.din(w_dff_A_V4wPDe5y5_0),.clk(gclk));
	jdff dff_A_c0InGZ4f6_0(.dout(w_dff_A_ZJF1DjtW6_0),.din(w_dff_A_c0InGZ4f6_0),.clk(gclk));
	jdff dff_A_ZJF1DjtW6_0(.dout(w_dff_A_tKPTQEpc5_0),.din(w_dff_A_ZJF1DjtW6_0),.clk(gclk));
	jdff dff_A_tKPTQEpc5_0(.dout(w_dff_A_FtQx97CX7_0),.din(w_dff_A_tKPTQEpc5_0),.clk(gclk));
	jdff dff_A_FtQx97CX7_0(.dout(w_dff_A_4TUbB0vq3_0),.din(w_dff_A_FtQx97CX7_0),.clk(gclk));
	jdff dff_A_4TUbB0vq3_0(.dout(w_dff_A_orJTJbDA6_0),.din(w_dff_A_4TUbB0vq3_0),.clk(gclk));
	jdff dff_A_orJTJbDA6_0(.dout(w_dff_A_J8xnWMmK8_0),.din(w_dff_A_orJTJbDA6_0),.clk(gclk));
	jdff dff_A_J8xnWMmK8_0(.dout(G447gat),.din(w_dff_A_J8xnWMmK8_0),.clk(gclk));
	jdff dff_A_vEUawqo43_2(.dout(w_dff_A_U977mjRo7_0),.din(w_dff_A_vEUawqo43_2),.clk(gclk));
	jdff dff_A_U977mjRo7_0(.dout(w_dff_A_lCKS3kqa6_0),.din(w_dff_A_U977mjRo7_0),.clk(gclk));
	jdff dff_A_lCKS3kqa6_0(.dout(w_dff_A_OMh5MYx10_0),.din(w_dff_A_lCKS3kqa6_0),.clk(gclk));
	jdff dff_A_OMh5MYx10_0(.dout(w_dff_A_wPmuxMqR3_0),.din(w_dff_A_OMh5MYx10_0),.clk(gclk));
	jdff dff_A_wPmuxMqR3_0(.dout(w_dff_A_7BDasKBt7_0),.din(w_dff_A_wPmuxMqR3_0),.clk(gclk));
	jdff dff_A_7BDasKBt7_0(.dout(w_dff_A_V8PNeLYQ6_0),.din(w_dff_A_7BDasKBt7_0),.clk(gclk));
	jdff dff_A_V8PNeLYQ6_0(.dout(w_dff_A_jx1ARsVy3_0),.din(w_dff_A_V8PNeLYQ6_0),.clk(gclk));
	jdff dff_A_jx1ARsVy3_0(.dout(w_dff_A_EtJyfVQ54_0),.din(w_dff_A_jx1ARsVy3_0),.clk(gclk));
	jdff dff_A_EtJyfVQ54_0(.dout(w_dff_A_Mtk3Onhd8_0),.din(w_dff_A_EtJyfVQ54_0),.clk(gclk));
	jdff dff_A_Mtk3Onhd8_0(.dout(w_dff_A_DiFH2RKg5_0),.din(w_dff_A_Mtk3Onhd8_0),.clk(gclk));
	jdff dff_A_DiFH2RKg5_0(.dout(w_dff_A_7rYLz2Pt3_0),.din(w_dff_A_DiFH2RKg5_0),.clk(gclk));
	jdff dff_A_7rYLz2Pt3_0(.dout(w_dff_A_7hPpqPks9_0),.din(w_dff_A_7rYLz2Pt3_0),.clk(gclk));
	jdff dff_A_7hPpqPks9_0(.dout(w_dff_A_oz5oGohB1_0),.din(w_dff_A_7hPpqPks9_0),.clk(gclk));
	jdff dff_A_oz5oGohB1_0(.dout(w_dff_A_4z4pNh510_0),.din(w_dff_A_oz5oGohB1_0),.clk(gclk));
	jdff dff_A_4z4pNh510_0(.dout(w_dff_A_hqi8BIDZ9_0),.din(w_dff_A_4z4pNh510_0),.clk(gclk));
	jdff dff_A_hqi8BIDZ9_0(.dout(w_dff_A_Im0opok21_0),.din(w_dff_A_hqi8BIDZ9_0),.clk(gclk));
	jdff dff_A_Im0opok21_0(.dout(w_dff_A_O1IwgoSl3_0),.din(w_dff_A_Im0opok21_0),.clk(gclk));
	jdff dff_A_O1IwgoSl3_0(.dout(G448gat),.din(w_dff_A_O1IwgoSl3_0),.clk(gclk));
	jdff dff_A_pKviZhew7_2(.dout(w_dff_A_WUwHDdlA5_0),.din(w_dff_A_pKviZhew7_2),.clk(gclk));
	jdff dff_A_WUwHDdlA5_0(.dout(w_dff_A_MLBTSbsZ3_0),.din(w_dff_A_WUwHDdlA5_0),.clk(gclk));
	jdff dff_A_MLBTSbsZ3_0(.dout(w_dff_A_rpJgTuYi0_0),.din(w_dff_A_MLBTSbsZ3_0),.clk(gclk));
	jdff dff_A_rpJgTuYi0_0(.dout(w_dff_A_wK7XOcnt3_0),.din(w_dff_A_rpJgTuYi0_0),.clk(gclk));
	jdff dff_A_wK7XOcnt3_0(.dout(w_dff_A_lev5a7F41_0),.din(w_dff_A_wK7XOcnt3_0),.clk(gclk));
	jdff dff_A_lev5a7F41_0(.dout(w_dff_A_UJJdBNSA1_0),.din(w_dff_A_lev5a7F41_0),.clk(gclk));
	jdff dff_A_UJJdBNSA1_0(.dout(w_dff_A_1t61mpq78_0),.din(w_dff_A_UJJdBNSA1_0),.clk(gclk));
	jdff dff_A_1t61mpq78_0(.dout(w_dff_A_Uta5chsW1_0),.din(w_dff_A_1t61mpq78_0),.clk(gclk));
	jdff dff_A_Uta5chsW1_0(.dout(w_dff_A_83cjwK6v0_0),.din(w_dff_A_Uta5chsW1_0),.clk(gclk));
	jdff dff_A_83cjwK6v0_0(.dout(w_dff_A_FH7ENENa4_0),.din(w_dff_A_83cjwK6v0_0),.clk(gclk));
	jdff dff_A_FH7ENENa4_0(.dout(w_dff_A_CaQfbgwv1_0),.din(w_dff_A_FH7ENENa4_0),.clk(gclk));
	jdff dff_A_CaQfbgwv1_0(.dout(w_dff_A_9aTiXfNm9_0),.din(w_dff_A_CaQfbgwv1_0),.clk(gclk));
	jdff dff_A_9aTiXfNm9_0(.dout(w_dff_A_fGAdYluU9_0),.din(w_dff_A_9aTiXfNm9_0),.clk(gclk));
	jdff dff_A_fGAdYluU9_0(.dout(w_dff_A_KFEV1lyz5_0),.din(w_dff_A_fGAdYluU9_0),.clk(gclk));
	jdff dff_A_KFEV1lyz5_0(.dout(w_dff_A_Of2s9mnT3_0),.din(w_dff_A_KFEV1lyz5_0),.clk(gclk));
	jdff dff_A_Of2s9mnT3_0(.dout(w_dff_A_vTgbgUFr0_0),.din(w_dff_A_Of2s9mnT3_0),.clk(gclk));
	jdff dff_A_vTgbgUFr0_0(.dout(w_dff_A_MsihI2xx3_0),.din(w_dff_A_vTgbgUFr0_0),.clk(gclk));
	jdff dff_A_MsihI2xx3_0(.dout(G449gat),.din(w_dff_A_MsihI2xx3_0),.clk(gclk));
	jdff dff_A_DXYPJYMd4_2(.dout(w_dff_A_N7fzxBil4_0),.din(w_dff_A_DXYPJYMd4_2),.clk(gclk));
	jdff dff_A_N7fzxBil4_0(.dout(w_dff_A_LZTHB2zd1_0),.din(w_dff_A_N7fzxBil4_0),.clk(gclk));
	jdff dff_A_LZTHB2zd1_0(.dout(w_dff_A_aVmaBTBD5_0),.din(w_dff_A_LZTHB2zd1_0),.clk(gclk));
	jdff dff_A_aVmaBTBD5_0(.dout(w_dff_A_0RK32nxr3_0),.din(w_dff_A_aVmaBTBD5_0),.clk(gclk));
	jdff dff_A_0RK32nxr3_0(.dout(w_dff_A_XoEkWgyZ5_0),.din(w_dff_A_0RK32nxr3_0),.clk(gclk));
	jdff dff_A_XoEkWgyZ5_0(.dout(w_dff_A_RTHDuTM76_0),.din(w_dff_A_XoEkWgyZ5_0),.clk(gclk));
	jdff dff_A_RTHDuTM76_0(.dout(w_dff_A_eaZyWBaK5_0),.din(w_dff_A_RTHDuTM76_0),.clk(gclk));
	jdff dff_A_eaZyWBaK5_0(.dout(w_dff_A_4FoVSiQL7_0),.din(w_dff_A_eaZyWBaK5_0),.clk(gclk));
	jdff dff_A_4FoVSiQL7_0(.dout(w_dff_A_Loi7ElGu3_0),.din(w_dff_A_4FoVSiQL7_0),.clk(gclk));
	jdff dff_A_Loi7ElGu3_0(.dout(w_dff_A_5Xz8bkrc5_0),.din(w_dff_A_Loi7ElGu3_0),.clk(gclk));
	jdff dff_A_5Xz8bkrc5_0(.dout(w_dff_A_0ksjWoiW1_0),.din(w_dff_A_5Xz8bkrc5_0),.clk(gclk));
	jdff dff_A_0ksjWoiW1_0(.dout(w_dff_A_yS1bS6Kz8_0),.din(w_dff_A_0ksjWoiW1_0),.clk(gclk));
	jdff dff_A_yS1bS6Kz8_0(.dout(w_dff_A_tIx92P8k7_0),.din(w_dff_A_yS1bS6Kz8_0),.clk(gclk));
	jdff dff_A_tIx92P8k7_0(.dout(w_dff_A_5dtrpx958_0),.din(w_dff_A_tIx92P8k7_0),.clk(gclk));
	jdff dff_A_5dtrpx958_0(.dout(w_dff_A_d34oFi6j6_0),.din(w_dff_A_5dtrpx958_0),.clk(gclk));
	jdff dff_A_d34oFi6j6_0(.dout(w_dff_A_NUPHI5O48_0),.din(w_dff_A_d34oFi6j6_0),.clk(gclk));
	jdff dff_A_NUPHI5O48_0(.dout(w_dff_A_z2k2FgAq9_0),.din(w_dff_A_NUPHI5O48_0),.clk(gclk));
	jdff dff_A_z2k2FgAq9_0(.dout(w_dff_A_qE32jqNx9_0),.din(w_dff_A_z2k2FgAq9_0),.clk(gclk));
	jdff dff_A_qE32jqNx9_0(.dout(G450gat),.din(w_dff_A_qE32jqNx9_0),.clk(gclk));
	jdff dff_A_OLTbHvvH0_2(.dout(w_dff_A_7LwcjK0y0_0),.din(w_dff_A_OLTbHvvH0_2),.clk(gclk));
	jdff dff_A_7LwcjK0y0_0(.dout(w_dff_A_XYr7xw2H7_0),.din(w_dff_A_7LwcjK0y0_0),.clk(gclk));
	jdff dff_A_XYr7xw2H7_0(.dout(w_dff_A_QJtNXSHq5_0),.din(w_dff_A_XYr7xw2H7_0),.clk(gclk));
	jdff dff_A_QJtNXSHq5_0(.dout(w_dff_A_OOk4ScND3_0),.din(w_dff_A_QJtNXSHq5_0),.clk(gclk));
	jdff dff_A_OOk4ScND3_0(.dout(w_dff_A_8Fg2Lyhj1_0),.din(w_dff_A_OOk4ScND3_0),.clk(gclk));
	jdff dff_A_8Fg2Lyhj1_0(.dout(w_dff_A_XMianCNc7_0),.din(w_dff_A_8Fg2Lyhj1_0),.clk(gclk));
	jdff dff_A_XMianCNc7_0(.dout(w_dff_A_fNWX4ibp4_0),.din(w_dff_A_XMianCNc7_0),.clk(gclk));
	jdff dff_A_fNWX4ibp4_0(.dout(w_dff_A_oWhyp7Er3_0),.din(w_dff_A_fNWX4ibp4_0),.clk(gclk));
	jdff dff_A_oWhyp7Er3_0(.dout(w_dff_A_RF5GxOWV6_0),.din(w_dff_A_oWhyp7Er3_0),.clk(gclk));
	jdff dff_A_RF5GxOWV6_0(.dout(w_dff_A_zNJCibHF9_0),.din(w_dff_A_RF5GxOWV6_0),.clk(gclk));
	jdff dff_A_zNJCibHF9_0(.dout(w_dff_A_6Bnlvj034_0),.din(w_dff_A_zNJCibHF9_0),.clk(gclk));
	jdff dff_A_6Bnlvj034_0(.dout(w_dff_A_tt1CmXvZ1_0),.din(w_dff_A_6Bnlvj034_0),.clk(gclk));
	jdff dff_A_tt1CmXvZ1_0(.dout(w_dff_A_7BoktcCx1_0),.din(w_dff_A_tt1CmXvZ1_0),.clk(gclk));
	jdff dff_A_7BoktcCx1_0(.dout(w_dff_A_NRtespHK1_0),.din(w_dff_A_7BoktcCx1_0),.clk(gclk));
	jdff dff_A_NRtespHK1_0(.dout(w_dff_A_FScb5QMa7_0),.din(w_dff_A_NRtespHK1_0),.clk(gclk));
	jdff dff_A_FScb5QMa7_0(.dout(w_dff_A_xRMhYuOI2_0),.din(w_dff_A_FScb5QMa7_0),.clk(gclk));
	jdff dff_A_xRMhYuOI2_0(.dout(G767gat),.din(w_dff_A_xRMhYuOI2_0),.clk(gclk));
	jdff dff_A_eFK7LroM1_2(.dout(w_dff_A_sZxFQNy83_0),.din(w_dff_A_eFK7LroM1_2),.clk(gclk));
	jdff dff_A_sZxFQNy83_0(.dout(w_dff_A_X6bNZAtW3_0),.din(w_dff_A_sZxFQNy83_0),.clk(gclk));
	jdff dff_A_X6bNZAtW3_0(.dout(w_dff_A_Oyh92nqn6_0),.din(w_dff_A_X6bNZAtW3_0),.clk(gclk));
	jdff dff_A_Oyh92nqn6_0(.dout(w_dff_A_WKw2PRZy7_0),.din(w_dff_A_Oyh92nqn6_0),.clk(gclk));
	jdff dff_A_WKw2PRZy7_0(.dout(w_dff_A_HKqw4KX41_0),.din(w_dff_A_WKw2PRZy7_0),.clk(gclk));
	jdff dff_A_HKqw4KX41_0(.dout(w_dff_A_v4nydyvP1_0),.din(w_dff_A_HKqw4KX41_0),.clk(gclk));
	jdff dff_A_v4nydyvP1_0(.dout(w_dff_A_VUMnKgYs3_0),.din(w_dff_A_v4nydyvP1_0),.clk(gclk));
	jdff dff_A_VUMnKgYs3_0(.dout(w_dff_A_wlkJxLG59_0),.din(w_dff_A_VUMnKgYs3_0),.clk(gclk));
	jdff dff_A_wlkJxLG59_0(.dout(w_dff_A_SLq7dLTq7_0),.din(w_dff_A_wlkJxLG59_0),.clk(gclk));
	jdff dff_A_SLq7dLTq7_0(.dout(w_dff_A_rK3mPQif7_0),.din(w_dff_A_SLq7dLTq7_0),.clk(gclk));
	jdff dff_A_rK3mPQif7_0(.dout(w_dff_A_vztwDrbc9_0),.din(w_dff_A_rK3mPQif7_0),.clk(gclk));
	jdff dff_A_vztwDrbc9_0(.dout(w_dff_A_cDf4RW9v0_0),.din(w_dff_A_vztwDrbc9_0),.clk(gclk));
	jdff dff_A_cDf4RW9v0_0(.dout(w_dff_A_dmMIlVwQ1_0),.din(w_dff_A_cDf4RW9v0_0),.clk(gclk));
	jdff dff_A_dmMIlVwQ1_0(.dout(w_dff_A_T894taxk0_0),.din(w_dff_A_dmMIlVwQ1_0),.clk(gclk));
	jdff dff_A_T894taxk0_0(.dout(w_dff_A_zSOToXXM2_0),.din(w_dff_A_T894taxk0_0),.clk(gclk));
	jdff dff_A_zSOToXXM2_0(.dout(w_dff_A_s3u7Ckjo0_0),.din(w_dff_A_zSOToXXM2_0),.clk(gclk));
	jdff dff_A_s3u7Ckjo0_0(.dout(G768gat),.din(w_dff_A_s3u7Ckjo0_0),.clk(gclk));
	jdff dff_A_pS0wowaN6_2(.dout(w_dff_A_ks4a92Wh9_0),.din(w_dff_A_pS0wowaN6_2),.clk(gclk));
	jdff dff_A_ks4a92Wh9_0(.dout(w_dff_A_0vVOKW4o9_0),.din(w_dff_A_ks4a92Wh9_0),.clk(gclk));
	jdff dff_A_0vVOKW4o9_0(.dout(w_dff_A_mvXaCdjZ6_0),.din(w_dff_A_0vVOKW4o9_0),.clk(gclk));
	jdff dff_A_mvXaCdjZ6_0(.dout(w_dff_A_b5KCODrM2_0),.din(w_dff_A_mvXaCdjZ6_0),.clk(gclk));
	jdff dff_A_b5KCODrM2_0(.dout(w_dff_A_wL26Jx331_0),.din(w_dff_A_b5KCODrM2_0),.clk(gclk));
	jdff dff_A_wL26Jx331_0(.dout(w_dff_A_hp7UmHj04_0),.din(w_dff_A_wL26Jx331_0),.clk(gclk));
	jdff dff_A_hp7UmHj04_0(.dout(w_dff_A_jfC4LkO81_0),.din(w_dff_A_hp7UmHj04_0),.clk(gclk));
	jdff dff_A_jfC4LkO81_0(.dout(G850gat),.din(w_dff_A_jfC4LkO81_0),.clk(gclk));
	jdff dff_A_uKd4HO2L8_2(.dout(w_dff_A_HgCi46kM4_0),.din(w_dff_A_uKd4HO2L8_2),.clk(gclk));
	jdff dff_A_HgCi46kM4_0(.dout(w_dff_A_YpNUobZl3_0),.din(w_dff_A_HgCi46kM4_0),.clk(gclk));
	jdff dff_A_YpNUobZl3_0(.dout(w_dff_A_rAiVBEsX2_0),.din(w_dff_A_YpNUobZl3_0),.clk(gclk));
	jdff dff_A_rAiVBEsX2_0(.dout(G863gat),.din(w_dff_A_rAiVBEsX2_0),.clk(gclk));
	jdff dff_A_osBm35gL3_2(.dout(w_dff_A_SF9iIUlC6_0),.din(w_dff_A_osBm35gL3_2),.clk(gclk));
	jdff dff_A_SF9iIUlC6_0(.dout(w_dff_A_5JSJaS396_0),.din(w_dff_A_SF9iIUlC6_0),.clk(gclk));
	jdff dff_A_5JSJaS396_0(.dout(w_dff_A_aatVJbvH0_0),.din(w_dff_A_5JSJaS396_0),.clk(gclk));
	jdff dff_A_aatVJbvH0_0(.dout(G864gat),.din(w_dff_A_aatVJbvH0_0),.clk(gclk));
	jdff dff_A_TGjlIEZu5_2(.dout(w_dff_A_OZvexL6z0_0),.din(w_dff_A_TGjlIEZu5_2),.clk(gclk));
	jdff dff_A_OZvexL6z0_0(.dout(w_dff_A_2fore71h0_0),.din(w_dff_A_OZvexL6z0_0),.clk(gclk));
	jdff dff_A_2fore71h0_0(.dout(w_dff_A_hncFd4F85_0),.din(w_dff_A_2fore71h0_0),.clk(gclk));
	jdff dff_A_hncFd4F85_0(.dout(w_dff_A_ZHe4fB7d1_0),.din(w_dff_A_hncFd4F85_0),.clk(gclk));
	jdff dff_A_ZHe4fB7d1_0(.dout(w_dff_A_Hj0sHmmF5_0),.din(w_dff_A_ZHe4fB7d1_0),.clk(gclk));
	jdff dff_A_Hj0sHmmF5_0(.dout(G865gat),.din(w_dff_A_Hj0sHmmF5_0),.clk(gclk));
	jdff dff_A_pjkRVhk99_2(.dout(w_dff_A_Ve8CQfh89_0),.din(w_dff_A_pjkRVhk99_2),.clk(gclk));
	jdff dff_A_Ve8CQfh89_0(.dout(G866gat),.din(w_dff_A_Ve8CQfh89_0),.clk(gclk));
	jdff dff_A_cQvl11VV9_2(.dout(w_dff_A_X7xuBf9F5_0),.din(w_dff_A_cQvl11VV9_2),.clk(gclk));
	jdff dff_A_X7xuBf9F5_0(.dout(G874gat),.din(w_dff_A_X7xuBf9F5_0),.clk(gclk));
endmodule

