module gf_c499(Gic4, Gic2, Gid31, Gid30, Gid28, Gid10, Gic0, Gid8, Gid4, Gid2, Gic6, Gid14, Gid7, Gid15, Gid5, Gid1, Gid6, Gid11, Gic5, Gid9, Gic3, Gid25, Gid12, Gid0, Gr, Gic1, Gid13, Gid29, Gid16, Gid21, Gid17, Gid18, Gid22, Gid3, Gid19, Gic7, Gid23, Gid24, Gid26, Gid20, Gid27, God31, God30, God29, God9, God24, God10, God8, God16, God25, God19, God7, God11, God13, God6, God4, God17, God12, God23, God3, God2, God1, God0, God14, God15, God22, God20, God21, God5, God18, God26, God27, God28);
    input Gic4, Gic2, Gid31, Gid30, Gid28, Gid10, Gic0, Gid8, Gid4, Gid2, Gic6, Gid14, Gid7, Gid15, Gid5, Gid1, Gid6, Gid11, Gic5, Gid9, Gic3, Gid25, Gid12, Gid0, Gr, Gic1, Gid13, Gid29, Gid16, Gid21, Gid17, Gid18, Gid22, Gid3, Gid19, Gic7, Gid23, Gid24, Gid26, Gid20, Gid27;
    output God31, God30, God29, God9, God24, God10, God8, God16, God25, God19, God7, God11, God13, God6, God4, God17, God12, God23, God3, God2, God1, God0, God14, God15, God22, God20, God21, God5, God18, God26, God27, God28;
    wire n76;
    wire n80;
    wire n84;
    wire n88;
    wire n92;
    wire n96;
    wire n100;
    wire n104;
    wire n108;
    wire n112;
    wire n116;
    wire n120;
    wire n124;
    wire n128;
    wire n132;
    wire n136;
    wire n140;
    wire n143;
    wire n147;
    wire n151;
    wire n155;
    wire n159;
    wire n163;
    wire n167;
    wire n171;
    wire n175;
    wire n179;
    wire n183;
    wire n187;
    wire n191;
    wire n195;
    wire n199;
    wire n203;
    wire n207;
    wire n211;
    wire n215;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n243;
    wire n247;
    wire n251;
    wire n255;
    wire n259;
    wire n263;
    wire n267;
    wire n271;
    wire n275;
    wire n279;
    wire n283;
    wire n287;
    wire n291;
    wire n295;
    wire n298;
    wire n302;
    wire n306;
    wire n310;
    wire n314;
    wire n318;
    wire n322;
    wire n326;
    wire n329;
    wire n333;
    wire n337;
    wire n341;
    wire n345;
    wire n349;
    wire n353;
    wire n357;
    wire n361;
    wire n365;
    wire n369;
    wire n373;
    wire n377;
    wire n381;
    wire n384;
    wire n388;
    wire n392;
    wire n395;
    wire n399;
    wire n403;
    wire n407;
    wire n411;
    wire n415;
    wire n419;
    wire n423;
    wire n427;
    wire n431;
    wire n435;
    wire n439;
    wire n443;
    wire n447;
    wire n451;
    wire n455;
    wire n459;
    wire n462;
    wire n466;
    wire n470;
    wire n474;
    wire n478;
    wire n482;
    wire n486;
    wire n490;
    wire n494;
    wire n498;
    wire n502;
    wire n506;
    wire n510;
    wire n514;
    wire n518;
    wire n522;
    wire n526;
    wire n529;
    wire n533;
    wire n537;
    wire n541;
    wire n545;
    wire n549;
    wire n553;
    wire n557;
    wire n561;
    wire n565;
    wire n569;
    wire n573;
    wire n576;
    wire n580;
    wire n584;
    wire n588;
    wire n592;
    wire n596;
    wire n600;
    wire n604;
    wire n608;
    wire n612;
    wire n616;
    wire n620;
    wire n624;
    wire n628;
    wire n632;
    wire n636;
    wire n640;
    wire n644;
    wire n648;
    wire n652;
    wire n656;
    wire n660;
    wire n664;
    wire n668;
    wire n672;
    wire n676;
    wire n680;
    wire n684;
    wire n688;
    wire n692;
    wire n696;
    wire n700;
    wire n704;
    wire n708;
    wire n712;
    wire n720;
    wire n728;
    wire n736;
    wire n744;
    wire n748;
    wire n752;
    wire n760;
    wire n768;
    wire n776;
    wire n784;
    wire n788;
    wire n792;
    wire n796;
    wire n804;
    wire n812;
    wire n820;
    wire n828;
    wire n832;
    wire n840;
    wire n848;
    wire n856;
    wire n1280;
    wire n1284;
    wire n1287;
    wire n1289;
    wire n1293;
    wire n1296;
    wire n1299;
    wire n1302;
    wire n1305;
    wire n1307;
    wire n1310;
    wire n1313;
    wire n1316;
    wire n1319;
    wire n1322;
    wire n1325;
    wire n1328;
    wire n1331;
    wire n1334;
    wire n1337;
    wire n1340;
    wire n1343;
    wire n1346;
    wire n1349;
    wire n1352;
    wire n1355;
    wire n1358;
    wire n1361;
    wire n1364;
    wire n1368;
    wire n1371;
    wire n1374;
    wire n1376;
    wire n1379;
    wire n1382;
    wire n1385;
    wire n1388;
    wire n1392;
    wire n1395;
    wire n1398;
    wire n1401;
    wire n1403;
    wire n1406;
    wire n1409;
    wire n1412;
    wire n1415;
    wire n1419;
    wire n1422;
    wire n1425;
    wire n1427;
    wire n1430;
    wire n1433;
    wire n1436;
    wire n1439;
    wire n1442;
    wire n1445;
    wire n1448;
    wire n1451;
    wire n1454;
    wire n1457;
    wire n1460;
    wire n1463;
    wire n1466;
    wire n1469;
    wire n1472;
    wire n1475;
    wire n1478;
    wire n1481;
    wire n1484;
    wire n1487;
    wire n1490;
    wire n1493;
    wire n1496;
    wire n1499;
    wire n1502;
    wire n1505;
    wire n1509;
    wire n1511;
    wire n1514;
    wire n1517;
    wire n1520;
    wire n1523;
    wire n1526;
    wire n1529;
    wire n1532;
    wire n1535;
    wire n1538;
    wire n1541;
    wire n1544;
    wire n1547;
    wire n1550;
    wire n1553;
    wire n1556;
    wire n1559;
    wire n1562;
    wire n1565;
    wire n1568;
    wire n1571;
    wire n1574;
    wire n1577;
    wire n1580;
    wire n1583;
    wire n1586;
    wire n1589;
    wire n1592;
    wire n1595;
    wire n1599;
    wire n1601;
    wire n1604;
    wire n1607;
    wire n1610;
    wire n1613;
    wire n1616;
    wire n1619;
    wire n1622;
    wire n1625;
    wire n1628;
    wire n1631;
    wire n1634;
    wire n1637;
    wire n1640;
    wire n1643;
    wire n1646;
    wire n1649;
    wire n1652;
    wire n1655;
    wire n1658;
    wire n1661;
    wire n1664;
    wire n1667;
    wire n1670;
    wire n1673;
    wire n1676;
    wire n1679;
    wire n1682;
    wire n1685;
    wire n1688;
    wire n1691;
    wire n1694;
    wire n1697;
    wire n1700;
    wire n1703;
    wire n1706;
    wire n1709;
    wire n1712;
    wire n1715;
    wire n1718;
    wire n1721;
    wire n1724;
    wire n1727;
    wire n1730;
    wire n1733;
    wire n1736;
    wire n1739;
    wire n1742;
    wire n1745;
    wire n1748;
    wire n1751;
    wire n1754;
    wire n1757;
    wire n1760;
    wire n1763;
    wire n1766;
    wire n1769;
    wire n1772;
    wire n1775;
    wire n1778;
    wire n1781;
    wire n1784;
    wire n1787;
    wire n1790;
    wire n1793;
    wire n1796;
    wire n1799;
    wire n1802;
    wire n1805;
    wire n1808;
    wire n1811;
    wire n1814;
    wire n1817;
    wire n1820;
    wire n1823;
    wire n1826;
    wire n1829;
    wire n1832;
    wire n1835;
    wire n1838;
    wire n1841;
    wire n1844;
    wire n1847;
    wire n1850;
    wire n1853;
    wire n1856;
    wire n1859;
    wire n1863;
    wire n1866;
    wire n1869;
    wire n1872;
    wire n1874;
    wire n1877;
    wire n1880;
    wire n1883;
    wire n1886;
    wire n1889;
    wire n1892;
    wire n1895;
    wire n1898;
    wire n1901;
    wire n1904;
    wire n1907;
    wire n1910;
    wire n1913;
    wire n1916;
    wire n1919;
    wire n1922;
    wire n1925;
    wire n1928;
    wire n1931;
    wire n1934;
    wire n1937;
    wire n1940;
    wire n1943;
    wire n1946;
    wire n1949;
    wire n1952;
    wire n1955;
    wire n1958;
    wire n1961;
    wire n1964;
    wire n1967;
    wire n1970;
    wire n1973;
    wire n1976;
    wire n1979;
    wire n1982;
    wire n1985;
    wire n1988;
    wire n1991;
    wire n1994;
    wire n1997;
    wire n2000;
    wire n2003;
    wire n2006;
    wire n2009;
    wire n2012;
    wire n2015;
    wire n2018;
    wire n2021;
    wire n2024;
    wire n2027;
    wire n2030;
    wire n2033;
    wire n2036;
    wire n2039;
    wire n2042;
    wire n2045;
    wire n2048;
    wire n2051;
    wire n2054;
    wire n2057;
    wire n2060;
    wire n2063;
    wire n2066;
    wire n2069;
    wire n2072;
    wire n2075;
    wire n2078;
    wire n2081;
    wire n2084;
    wire n2087;
    wire n2090;
    wire n2093;
    wire n2096;
    wire n2099;
    wire n2102;
    wire n2105;
    wire n2108;
    wire n2111;
    wire n2114;
    wire n2117;
    wire n2120;
    wire n2123;
    wire n2126;
    wire n2129;
    wire n2132;
    wire n2135;
    wire n2138;
    wire n2141;
    wire n2144;
    wire n2147;
    wire n2150;
    wire n2153;
    wire n2156;
    wire n2159;
    wire n2162;
    wire n2165;
    wire n2168;
    wire n2171;
    wire n2174;
    wire n2177;
    wire n2180;
    wire n2183;
    wire n2186;
    wire n2189;
    wire n2192;
    wire n2195;
    wire n2198;
    wire n2201;
    wire n2204;
    wire n2207;
    wire n2210;
    wire n2213;
    wire n2216;
    wire n2219;
    wire n2222;
    wire n2225;
    wire n2228;
    wire n2231;
    wire n2234;
    wire n2237;
    wire n2240;
    wire n2243;
    wire n2246;
    wire n2249;
    wire n2252;
    wire n2255;
    wire n2258;
    wire n2261;
    wire n2264;
    wire n2267;
    wire n2270;
    wire n2273;
    wire n2276;
    wire n2279;
    wire n2282;
    wire n2285;
    wire n2288;
    wire n2291;
    wire n2294;
    wire n2297;
    wire n2300;
    wire n2303;
    wire n2306;
    wire n2309;
    wire n2312;
    wire n2315;
    wire n2318;
    wire n2321;
    wire n2324;
    wire n2327;
    wire n2330;
    wire n2333;
    wire n2336;
    wire n2339;
    wire n2342;
    wire n2345;
    wire n2348;
    wire n2351;
    wire n2354;
    wire n2357;
    wire n2360;
    wire n2363;
    wire n2366;
    wire n2369;
    wire n2372;
    wire n2375;
    wire n2378;
    wire n2381;
    wire n2384;
    wire n2387;
    wire n2390;
    wire n2393;
    wire n2396;
    wire n2399;
    wire n2402;
    wire n2405;
    wire n2408;
    wire n2411;
    wire n2414;
    wire n2417;
    wire n2420;
    wire n2423;
    wire n2426;
    wire n2429;
    wire n2432;
    wire n2435;
    wire n2438;
    wire n2441;
    wire n2444;
    wire n2447;
    wire n2450;
    wire n2453;
    wire n2456;
    wire n2459;
    wire n2462;
    wire n2465;
    wire n2468;
    wire n2471;
    wire n2474;
    wire n2477;
    wire n2480;
    wire n2483;
    wire n2486;
    wire n2489;
    wire n2492;
    wire n2495;
    wire n2498;
    wire n2501;
    wire n2504;
    wire n2507;
    wire n2510;
    wire n2513;
    wire n2516;
    wire n2519;
    wire n2522;
    wire n2525;
    wire n2528;
    wire n2531;
    wire n2534;
    wire n2537;
    wire n2540;
    wire n2543;
    wire n2546;
    wire n2549;
    wire n2552;
    wire n2555;
    wire n2558;
    wire n2561;
    wire n2564;
    wire n2567;
    wire n2570;
    wire n2573;
    wire n2576;
    wire n2579;
    wire n2582;
    wire n2585;
    wire n2588;
    wire n2591;
    wire n2594;
    wire n2597;
    wire n2600;
    wire n2603;
    wire n2606;
    wire n2609;
    wire n2612;
    wire n2615;
    wire n2618;
    wire n2621;
    wire n2624;
    wire n2627;
    wire n2630;
    wire n2633;
    wire n2636;
    wire n2639;
    wire n2642;
    wire n2645;
    wire n2648;
    wire n2651;
    wire n2654;
    wire n2657;
    wire n2660;
    jxor g000(.dinb(Gid8), .dina(Gid12), .dout(n76));
    jxor g001(.dinb(Gid0), .dina(Gid4), .dout(n80));
    jxor g002(.dinb(n76), .dina(n80), .dout(n84));
    jand g003(.dinb(Gic0), .dina(Gr), .dout(n88));
    jxor g004(.dinb(n84), .dina(n1739), .dout(n92));
    jxor g005(.dinb(Gid18), .dina(Gid19), .dout(n96));
    jxor g006(.dinb(Gid16), .dina(Gid17), .dout(n100));
    jxor g007(.dinb(n96), .dina(n100), .dout(n104));
    jxor g008(.dinb(Gid22), .dina(Gid23), .dout(n108));
    jxor g009(.dinb(Gid20), .dina(Gid21), .dout(n112));
    jxor g010(.dinb(n108), .dina(n112), .dout(n116));
    jxor g011(.dinb(n104), .dina(n116), .dout(n120));
    jxor g012(.dinb(n92), .dina(n120), .dout(n124));
    jxor g013(.dinb(Gid27), .dina(Gid31), .dout(n128));
    jxor g014(.dinb(Gid19), .dina(Gid23), .dout(n132));
    jxor g015(.dinb(n128), .dina(n132), .dout(n136));
    jand g016(.dinb(Gic7), .dina(Gr), .dout(n140));
    jnot g017(.din(n140), .dout(n143));
    jxor g018(.dinb(n136), .dina(n143), .dout(n147));
    jxor g019(.dinb(Gid6), .dina(Gid7), .dout(n151));
    jxor g020(.dinb(Gid4), .dina(Gid5), .dout(n155));
    jxor g021(.dinb(n151), .dina(n155), .dout(n159));
    jxor g022(.dinb(Gid14), .dina(Gid15), .dout(n163));
    jxor g023(.dinb(Gid12), .dina(Gid13), .dout(n167));
    jxor g024(.dinb(n163), .dina(n167), .dout(n171));
    jxor g025(.dinb(n159), .dina(n171), .dout(n175));
    jxor g026(.dinb(n147), .dina(n175), .dout(n179));
    jxor g027(.dinb(Gid26), .dina(Gid30), .dout(n183));
    jxor g028(.dinb(Gid18), .dina(Gid22), .dout(n187));
    jxor g029(.dinb(n183), .dina(n187), .dout(n191));
    jand g030(.dinb(Gic6), .dina(Gr), .dout(n195));
    jxor g031(.dinb(n191), .dina(n1509), .dout(n199));
    jxor g032(.dinb(Gid2), .dina(Gid3), .dout(n203));
    jxor g033(.dinb(Gid0), .dina(Gid1), .dout(n207));
    jxor g034(.dinb(n203), .dina(n207), .dout(n211));
    jxor g035(.dinb(Gid10), .dina(Gid11), .dout(n215));
    jxor g036(.dinb(Gid8), .dina(Gid9), .dout(n219));
    jxor g037(.dinb(n215), .dina(n219), .dout(n223));
    jxor g038(.dinb(n211), .dina(n223), .dout(n227));
    jxor g039(.dinb(n199), .dina(n227), .dout(n231));
    jand g040(.dinb(n179), .dina(n231), .dout(n235));
    jxor g041(.dinb(Gid9), .dina(Gid13), .dout(n239));
    jxor g042(.dinb(Gid1), .dina(Gid5), .dout(n243));
    jxor g043(.dinb(n239), .dina(n243), .dout(n247));
    jand g044(.dinb(Gic1), .dina(Gr), .dout(n251));
    jxor g045(.dinb(n247), .dina(n1616), .dout(n255));
    jxor g046(.dinb(Gid30), .dina(Gid31), .dout(n259));
    jxor g047(.dinb(Gid28), .dina(Gid29), .dout(n263));
    jxor g048(.dinb(n259), .dina(n263), .dout(n267));
    jxor g049(.dinb(Gid26), .dina(Gid27), .dout(n271));
    jxor g050(.dinb(Gid24), .dina(Gid25), .dout(n275));
    jxor g051(.dinb(n271), .dina(n275), .dout(n279));
    jxor g052(.dinb(n267), .dina(n279), .dout(n283));
    jxor g053(.dinb(n255), .dina(n283), .dout(n287));
    jxor g054(.dinb(n124), .dina(n287), .dout(n291));
    jand g055(.dinb(Gic3), .dina(Gr), .dout(n295));
    jnot g056(.din(n295), .dout(n298));
    jxor g057(.dinb(n267), .dina(n298), .dout(n302));
    jxor g058(.dinb(Gid11), .dina(Gid15), .dout(n306));
    jxor g059(.dinb(Gid3), .dina(Gid7), .dout(n310));
    jxor g060(.dinb(n306), .dina(n310), .dout(n314));
    jxor g061(.dinb(n116), .dina(n314), .dout(n318));
    jxor g062(.dinb(n302), .dina(n318), .dout(n322));
    jand g063(.dinb(Gic2), .dina(Gr), .dout(n326));
    jnot g064(.din(n326), .dout(n329));
    jxor g065(.dinb(n279), .dina(n329), .dout(n333));
    jxor g066(.dinb(Gid10), .dina(Gid14), .dout(n337));
    jxor g067(.dinb(Gid2), .dina(Gid6), .dout(n341));
    jxor g068(.dinb(n337), .dina(n341), .dout(n345));
    jxor g069(.dinb(n104), .dina(n345), .dout(n349));
    jxor g070(.dinb(n333), .dina(n349), .dout(n353));
    jand g071(.dinb(n322), .dina(n353), .dout(n357));
    jand g072(.dinb(n291), .dina(n357), .dout(n361));
    jxor g073(.dinb(n267), .dina(n2528), .dout(n365));
    jxor g074(.dinb(n365), .dina(n318), .dout(n369));
    jxor g075(.dinb(n279), .dina(n2126), .dout(n373));
    jxor g076(.dinb(n373), .dina(n349), .dout(n377));
    jxor g077(.dinb(n369), .dina(n377), .dout(n381));
    jnot g078(.din(n88), .dout(n384));
    jxor g079(.dinb(n84), .dina(n384), .dout(n388));
    jxor g080(.dinb(n388), .dina(n120), .dout(n392));
    jnot g081(.din(n251), .dout(n395));
    jxor g082(.dinb(n247), .dina(n395), .dout(n399));
    jxor g083(.dinb(n399), .dina(n283), .dout(n403));
    jand g084(.dinb(n392), .dina(n403), .dout(n407));
    jand g085(.dinb(n381), .dina(n407), .dout(n411));
    jor g086(.dinb(n361), .dina(n411), .dout(n415));
    jxor g087(.dinb(Gid24), .dina(Gid28), .dout(n419));
    jxor g088(.dinb(Gid16), .dina(Gid20), .dout(n423));
    jxor g089(.dinb(n419), .dina(n423), .dout(n427));
    jand g090(.dinb(Gic4), .dina(Gr), .dout(n431));
    jxor g091(.dinb(n427), .dina(n1599), .dout(n435));
    jxor g092(.dinb(n159), .dina(n211), .dout(n439));
    jxor g093(.dinb(n435), .dina(n439), .dout(n443));
    jxor g094(.dinb(Gid25), .dina(Gid29), .dout(n447));
    jxor g095(.dinb(Gid17), .dina(Gid21), .dout(n451));
    jxor g096(.dinb(n447), .dina(n451), .dout(n455));
    jand g097(.dinb(Gic5), .dina(Gr), .dout(n459));
    jnot g098(.din(n459), .dout(n462));
    jxor g099(.dinb(n455), .dina(n462), .dout(n466));
    jxor g100(.dinb(n171), .dina(n223), .dout(n470));
    jxor g101(.dinb(n466), .dina(n470), .dout(n474));
    jand g102(.dinb(n443), .dina(n474), .dout(n478));
    jand g103(.dinb(n415), .dina(n1287), .dout(n482));
    jand g104(.dinb(n1289), .dina(n482), .dout(n486));
    jand g105(.dinb(n1352), .dina(n486), .dout(n490));
    jxor g106(.dinb(n1772), .dina(n490), .dout(n494));
    jand g107(.dinb(n1337), .dina(n486), .dout(n498));
    jxor g108(.dinb(n1649), .dina(n498), .dout(n502));
    jand g109(.dinb(n1307), .dina(n486), .dout(n506));
    jxor g110(.dinb(n1904), .dina(n506), .dout(n510));
    jand g111(.dinb(n1322), .dina(n486), .dout(n514));
    jxor g112(.dinb(n2306), .dina(n514), .dout(n518));
    jxor g113(.dinb(n136), .dina(n1550), .dout(n522));
    jxor g114(.dinb(n522), .dina(n175), .dout(n526));
    jnot g115(.din(n231), .dout(n529));
    jand g116(.dinb(n1511), .dina(n529), .dout(n533));
    jand g117(.dinb(n415), .dina(n1305), .dout(n537));
    jand g118(.dinb(n1280), .dina(n537), .dout(n541));
    jand g119(.dinb(n1376), .dina(n541), .dout(n545));
    jxor g120(.dinb(n1742), .dina(n545), .dout(n549));
    jand g121(.dinb(n1601), .dina(n541), .dout(n553));
    jxor g122(.dinb(n1619), .dina(n553), .dout(n557));
    jand g123(.dinb(n1403), .dina(n541), .dout(n561));
    jxor g124(.dinb(n1874), .dina(n561), .dout(n565));
    jand g125(.dinb(n2261), .dina(n541), .dout(n569));
    jxor g126(.dinb(n2276), .dina(n569), .dout(n573));
    jnot g127(.din(n443), .dout(n576));
    jxor g128(.dinb(n455), .dina(n1556), .dout(n580));
    jxor g129(.dinb(n580), .dina(n470), .dout(n584));
    jand g130(.dinb(n576), .dina(n1427), .dout(n588));
    jand g131(.dinb(n1296), .dina(n415), .dout(n592));
    jand g132(.dinb(n1302), .dina(n592), .dout(n596));
    jand g133(.dinb(n1376), .dina(n596), .dout(n600));
    jxor g134(.dinb(n1832), .dina(n600), .dout(n604));
    jand g135(.dinb(n1601), .dina(n596), .dout(n608));
    jxor g136(.dinb(n1709), .dina(n608), .dout(n612));
    jand g137(.dinb(n1403), .dina(n596), .dout(n616));
    jxor g138(.dinb(n1964), .dina(n616), .dout(n620));
    jand g139(.dinb(n2261), .dina(n596), .dout(n624));
    jxor g140(.dinb(n2366), .dina(n624), .dout(n628));
    jand g141(.dinb(n537), .dina(n1302), .dout(n632));
    jand g142(.dinb(n1376), .dina(n632), .dout(n636));
    jxor g143(.dinb(n1802), .dina(n636), .dout(n640));
    jand g144(.dinb(n1601), .dina(n632), .dout(n644));
    jxor g145(.dinb(n1679), .dina(n644), .dout(n648));
    jand g146(.dinb(n1403), .dina(n632), .dout(n652));
    jxor g147(.dinb(n1934), .dina(n652), .dout(n656));
    jand g148(.dinb(n2261), .dina(n632), .dout(n660));
    jxor g149(.dinb(n2336), .dina(n660), .dout(n664));
    jand g150(.dinb(n322), .dina(n377), .dout(n668));
    jand g151(.dinb(n124), .dina(n403), .dout(n672));
    jxor g152(.dinb(n526), .dina(n231), .dout(n676));
    jand g153(.dinb(n1553), .dina(n676), .dout(n680));
    jand g154(.dinb(n1559), .dina(n680), .dout(n684));
    jxor g155(.dinb(n443), .dina(n584), .dout(n688));
    jand g156(.dinb(n1466), .dina(n688), .dout(n692));
    jand g157(.dinb(n1469), .dina(n692), .dout(n696));
    jor g158(.dinb(n684), .dina(n696), .dout(n700));
    jand g159(.dinb(n1374), .dina(n700), .dout(n704));
    jand g160(.dinb(n1401), .dina(n704), .dout(n708));
    jand g161(.dinb(n1562), .dina(n708), .dout(n712));
    jxor g162(.dinb(n2027), .dina(n712), .dout(God16));
    jand g163(.dinb(n1430), .dina(n708), .dout(n720));
    jxor g164(.dinb(n1994), .dina(n720), .dout(God17));
    jand g165(.dinb(n1472), .dina(n708), .dout(n728));
    jxor g166(.dinb(n2093), .dina(n728), .dout(God18));
    jand g167(.dinb(n1514), .dina(n708), .dout(n736));
    jxor g168(.dinb(n2060), .dina(n736), .dout(God19));
    jand g169(.dinb(n369), .dina(n353), .dout(n744));
    jand g170(.dinb(n1872), .dina(n704), .dout(n748));
    jand g171(.dinb(n1562), .dina(n748), .dout(n752));
    jxor g172(.dinb(n2429), .dina(n752), .dout(God20));
    jand g173(.dinb(n1430), .dina(n748), .dout(n760));
    jxor g174(.dinb(n2396), .dina(n760), .dout(God21));
    jand g175(.dinb(n1472), .dina(n748), .dout(n768));
    jxor g176(.dinb(n2495), .dina(n768), .dout(God22));
    jand g177(.dinb(n1514), .dina(n748), .dout(n776));
    jxor g178(.dinb(n2462), .dina(n776), .dout(God23));
    jand g179(.dinb(n392), .dina(n287), .dout(n784));
    jand g180(.dinb(n1425), .dina(n700), .dout(n788));
    jand g181(.dinb(n1401), .dina(n788), .dout(n792));
    jand g182(.dinb(n1562), .dina(n792), .dout(n796));
    jxor g183(.dinb(n2162), .dina(n796), .dout(God24));
    jand g184(.dinb(n1430), .dina(n792), .dout(n804));
    jxor g185(.dinb(n2129), .dina(n804), .dout(God25));
    jand g186(.dinb(n1472), .dina(n792), .dout(n812));
    jxor g187(.dinb(n2228), .dina(n812), .dout(God26));
    jand g188(.dinb(n1514), .dina(n792), .dout(n820));
    jxor g189(.dinb(n2195), .dina(n820), .dout(God27));
    jand g190(.dinb(n1872), .dina(n788), .dout(n828));
    jand g191(.dinb(n1580), .dina(n828), .dout(n832));
    jxor g192(.dinb(n2564), .dina(n832), .dout(God28));
    jand g193(.dinb(n1448), .dina(n828), .dout(n840));
    jxor g194(.dinb(n2531), .dina(n840), .dout(God29));
    jand g195(.dinb(n1490), .dina(n828), .dout(n848));
    jxor g196(.dinb(n2630), .dina(n848), .dout(God30));
    jand g197(.dinb(n1532), .dina(n828), .dout(n856));
    jxor g198(.dinb(n2597), .dina(n856), .dout(God31));
    jdff dff_A_7GIr0kJS3_2(.din(n664), .dout(God15));
    jdff dff_A_UxhabKGn3_2(.din(n656), .dout(God14));
    jdff dff_A_4nkykmME2_2(.din(n648), .dout(God13));
    jdff dff_A_wRRP0kLL9_2(.din(n640), .dout(God12));
    jdff dff_A_gri3Jqev7_2(.din(n628), .dout(God11));
    jdff dff_A_YC1eikXb3_2(.din(n620), .dout(God10));
    jdff dff_A_P1nnemrt1_2(.din(n612), .dout(God9));
    jdff dff_A_SsQEgfrU1_2(.din(n604), .dout(God8));
    jdff dff_A_XgvbmHBM3_2(.din(n573), .dout(God7));
    jdff dff_A_PYCXl0ap5_2(.din(n565), .dout(God6));
    jdff dff_A_n7m9VX7F7_2(.din(n557), .dout(God5));
    jdff dff_A_Fwn0Ij8d6_2(.din(n549), .dout(God4));
    jdff dff_A_VTAVybd45_2(.din(n518), .dout(God3));
    jdff dff_A_34PC55qj0_2(.din(n510), .dout(God2));
    jdff dff_A_5M6o6Ub95_2(.din(n502), .dout(God1));
    jdff dff_A_PMYQK5Tj0_2(.din(n494), .dout(God0));
    jdff dff_A_iJKwPfTv6_0(.din(Gid30), .dout(n2660));
    jdff dff_A_aBvtiYMn9_0(.din(n2660), .dout(n2657));
    jdff dff_A_pDS8zIsB7_0(.din(n2657), .dout(n2654));
    jdff dff_A_yZj45uEo2_0(.din(n2654), .dout(n2651));
    jdff dff_A_vpL9BUYb6_0(.din(n2651), .dout(n2648));
    jdff dff_A_6HlXHswn6_0(.din(n2648), .dout(n2645));
    jdff dff_A_AjSCsUfW6_0(.din(n2645), .dout(n2642));
    jdff dff_A_krNofpEG7_0(.din(n2642), .dout(n2639));
    jdff dff_A_fYFzoGo40_0(.din(n2639), .dout(n2636));
    jdff dff_A_5kiC1pva1_0(.din(n2636), .dout(n2633));
    jdff dff_A_R0VntRor0_0(.din(n2633), .dout(n2630));
    jdff dff_A_ErCKavnX3_0(.din(Gid31), .dout(n2627));
    jdff dff_A_su0c3OnU2_0(.din(n2627), .dout(n2624));
    jdff dff_A_Osg1ps4M8_0(.din(n2624), .dout(n2621));
    jdff dff_A_y0DY56H69_0(.din(n2621), .dout(n2618));
    jdff dff_A_BC7Rpd9W8_0(.din(n2618), .dout(n2615));
    jdff dff_A_4hMMClrs5_0(.din(n2615), .dout(n2612));
    jdff dff_A_tSlxDHv67_0(.din(n2612), .dout(n2609));
    jdff dff_A_dqvs45f62_0(.din(n2609), .dout(n2606));
    jdff dff_A_6cnefFmO1_0(.din(n2606), .dout(n2603));
    jdff dff_A_xEvsVRYM8_0(.din(n2603), .dout(n2600));
    jdff dff_A_xZbhjjVs0_0(.din(n2600), .dout(n2597));
    jdff dff_A_C0FtiK1q2_0(.din(Gid28), .dout(n2594));
    jdff dff_A_zYdL2D6e2_0(.din(n2594), .dout(n2591));
    jdff dff_A_WrbW5WG71_0(.din(n2591), .dout(n2588));
    jdff dff_A_fu0y72oP4_0(.din(n2588), .dout(n2585));
    jdff dff_A_Mad77qnx2_0(.din(n2585), .dout(n2582));
    jdff dff_A_6uFoeYcl2_0(.din(n2582), .dout(n2579));
    jdff dff_A_KTtfpoyp0_0(.din(n2579), .dout(n2576));
    jdff dff_A_uSrkTRLw1_0(.din(n2576), .dout(n2573));
    jdff dff_A_9dhgkiV36_0(.din(n2573), .dout(n2570));
    jdff dff_A_pjxyb87j2_0(.din(n2570), .dout(n2567));
    jdff dff_A_OvFkGplN9_0(.din(n2567), .dout(n2564));
    jdff dff_A_azHUBSfr1_0(.din(Gid29), .dout(n2561));
    jdff dff_A_WBG4S1Ro9_0(.din(n2561), .dout(n2558));
    jdff dff_A_78fXIHfE7_0(.din(n2558), .dout(n2555));
    jdff dff_A_IUELqlgn3_0(.din(n2555), .dout(n2552));
    jdff dff_A_DXADtZmy9_0(.din(n2552), .dout(n2549));
    jdff dff_A_1nL2d3l84_0(.din(n2549), .dout(n2546));
    jdff dff_A_jXpx4bnO2_0(.din(n2546), .dout(n2543));
    jdff dff_A_bLcg0G0I9_0(.din(n2543), .dout(n2540));
    jdff dff_A_GXEKt2T89_0(.din(n2540), .dout(n2537));
    jdff dff_A_1NfHusSD0_0(.din(n2537), .dout(n2534));
    jdff dff_A_I3AI6Ynl2_0(.din(n2534), .dout(n2531));
    jdff dff_A_ieHKHVNB2_0(.din(n295), .dout(n2528));
    jdff dff_A_dDbXMIj37_0(.din(Gid22), .dout(n2525));
    jdff dff_A_Wfivb2Fg1_0(.din(n2525), .dout(n2522));
    jdff dff_A_rEfNOk1Z8_0(.din(n2522), .dout(n2519));
    jdff dff_A_1NjX9CGf4_0(.din(n2519), .dout(n2516));
    jdff dff_A_TA17G0Iy6_0(.din(n2516), .dout(n2513));
    jdff dff_A_npAutbBS9_0(.din(n2513), .dout(n2510));
    jdff dff_A_KB8rMTdo9_0(.din(n2510), .dout(n2507));
    jdff dff_A_kpB5NQOi3_0(.din(n2507), .dout(n2504));
    jdff dff_A_6Ut0vQrG8_0(.din(n2504), .dout(n2501));
    jdff dff_A_T3JgPuRN1_0(.din(n2501), .dout(n2498));
    jdff dff_A_TUXxjpHt8_0(.din(n2498), .dout(n2495));
    jdff dff_A_MdgH81Vo4_0(.din(Gid23), .dout(n2492));
    jdff dff_A_44Qqi6fu9_0(.din(n2492), .dout(n2489));
    jdff dff_A_kXAsLSNA0_0(.din(n2489), .dout(n2486));
    jdff dff_A_oIdN7jbs0_0(.din(n2486), .dout(n2483));
    jdff dff_A_NxDc3Nsk1_0(.din(n2483), .dout(n2480));
    jdff dff_A_HgPP4Jc56_0(.din(n2480), .dout(n2477));
    jdff dff_A_BJiU8Dli1_0(.din(n2477), .dout(n2474));
    jdff dff_A_m0X0DNV68_0(.din(n2474), .dout(n2471));
    jdff dff_A_WvYyWxzg7_0(.din(n2471), .dout(n2468));
    jdff dff_A_xZ34f1IN0_0(.din(n2468), .dout(n2465));
    jdff dff_A_ZZGI2iuE9_0(.din(n2465), .dout(n2462));
    jdff dff_A_QMFA5xbD2_0(.din(Gid20), .dout(n2459));
    jdff dff_A_XW0H1AoH0_0(.din(n2459), .dout(n2456));
    jdff dff_A_SdPtLtkQ1_0(.din(n2456), .dout(n2453));
    jdff dff_A_uUIN0ozZ2_0(.din(n2453), .dout(n2450));
    jdff dff_A_m0p89FOw6_0(.din(n2450), .dout(n2447));
    jdff dff_A_WGwoBsqf6_0(.din(n2447), .dout(n2444));
    jdff dff_A_QVH7nSfG6_0(.din(n2444), .dout(n2441));
    jdff dff_A_QhE8VnNu5_0(.din(n2441), .dout(n2438));
    jdff dff_A_V5zIibt05_0(.din(n2438), .dout(n2435));
    jdff dff_A_lCN1uvi33_0(.din(n2435), .dout(n2432));
    jdff dff_A_X5Pwss0z4_0(.din(n2432), .dout(n2429));
    jdff dff_A_OWywckru0_0(.din(Gid21), .dout(n2426));
    jdff dff_A_Ubj9B6lp2_0(.din(n2426), .dout(n2423));
    jdff dff_A_E28qXkd37_0(.din(n2423), .dout(n2420));
    jdff dff_A_d1OKbcRq4_0(.din(n2420), .dout(n2417));
    jdff dff_A_iNpbyG9T4_0(.din(n2417), .dout(n2414));
    jdff dff_A_X95GqGPh5_0(.din(n2414), .dout(n2411));
    jdff dff_A_FK2uUZDw2_0(.din(n2411), .dout(n2408));
    jdff dff_A_wVx6AIv85_0(.din(n2408), .dout(n2405));
    jdff dff_A_mTG1dvKJ5_0(.din(n2405), .dout(n2402));
    jdff dff_A_EBBf7ufV7_0(.din(n2402), .dout(n2399));
    jdff dff_A_Rp9G3c4u3_0(.din(n2399), .dout(n2396));
    jdff dff_A_DnccThX34_0(.din(Gid11), .dout(n2393));
    jdff dff_A_xbrBFJZR3_0(.din(n2393), .dout(n2390));
    jdff dff_A_xEK5MWRf0_0(.din(n2390), .dout(n2387));
    jdff dff_A_ySQpeBkw8_0(.din(n2387), .dout(n2384));
    jdff dff_A_T4A39mOC7_0(.din(n2384), .dout(n2381));
    jdff dff_A_xmyBsTe45_0(.din(n2381), .dout(n2378));
    jdff dff_A_pBg22DGl9_0(.din(n2378), .dout(n2375));
    jdff dff_A_CBl3IIGX8_0(.din(n2375), .dout(n2372));
    jdff dff_A_QPhhcsxM2_0(.din(n2372), .dout(n2369));
    jdff dff_A_E4hNQIqu8_0(.din(n2369), .dout(n2366));
    jdff dff_A_9kS1c7it8_0(.din(Gid15), .dout(n2363));
    jdff dff_A_e7s5LfX73_0(.din(n2363), .dout(n2360));
    jdff dff_A_JuY88UlQ3_0(.din(n2360), .dout(n2357));
    jdff dff_A_aDdyPWb38_0(.din(n1287), .dout(n1280));
    jdff dff_B_rcJR4sP54_2(.din(n478), .dout(n1284));
    jdff dff_B_QzVgACRg1_2(.din(n1284), .dout(n1287));
    jdff dff_A_6GE9eT2e6_1(.din(n1296), .dout(n1289));
    jdff dff_B_Bv2Pjeql0_2(.din(n235), .dout(n1293));
    jdff dff_B_PvPK2uh24_2(.din(n1293), .dout(n1296));
    jdff dff_B_U6YQwxGQ5_2(.din(n588), .dout(n1299));
    jdff dff_B_u6YsHwn04_2(.din(n1299), .dout(n1302));
    jdff dff_B_K1qUrywU9_0(.din(n533), .dout(n1305));
    jdff dff_A_vYm9ffK76_0(.din(n1310), .dout(n1307));
    jdff dff_A_8m7vKhDh8_0(.din(n1313), .dout(n1310));
    jdff dff_A_jTKP7wBN4_0(.din(n1316), .dout(n1313));
    jdff dff_A_rdAhtn6n6_0(.din(n1319), .dout(n1316));
    jdff dff_A_BpR7RP2O6_0(.din(n377), .dout(n1319));
    jdff dff_A_IaMk4a494_0(.din(n1325), .dout(n1322));
    jdff dff_A_tz9wkayk6_0(.din(n1328), .dout(n1325));
    jdff dff_A_8CAR0Ip75_0(.din(n1331), .dout(n1328));
    jdff dff_A_nA7QdfNz7_0(.din(n1334), .dout(n1331));
    jdff dff_A_zKRcJdAD1_0(.din(n369), .dout(n1334));
    jdff dff_A_0QEC5RPS1_0(.din(n1340), .dout(n1337));
    jdff dff_A_rNaUt7z90_0(.din(n1343), .dout(n1340));
    jdff dff_A_oWVKbCJm2_0(.din(n1346), .dout(n1343));
    jdff dff_A_njpK3b4y3_0(.din(n1349), .dout(n1346));
    jdff dff_A_Yz4tRNK61_0(.din(n287), .dout(n1349));
    jdff dff_A_MXWJnoX17_0(.din(n1355), .dout(n1352));
    jdff dff_A_4XJDLIu03_0(.din(n1358), .dout(n1355));
    jdff dff_A_gz9d8heg8_0(.din(n1361), .dout(n1358));
    jdff dff_A_xlqmfJVf2_0(.din(n1364), .dout(n1361));
    jdff dff_A_AcoMs2LU8_0(.din(n124), .dout(n1364));
    jdff dff_B_aFKaFGhu2_1(.din(n672), .dout(n1368));
    jdff dff_B_eq9fE1rP2_1(.din(n1368), .dout(n1371));
    jdff dff_B_ZnGIKCip6_1(.din(n1371), .dout(n1374));
    jdff dff_A_Lcf74BXH1_0(.din(n1379), .dout(n1376));
    jdff dff_A_yQRXNvKO5_0(.din(n1382), .dout(n1379));
    jdff dff_A_GNcnHxCq3_0(.din(n1385), .dout(n1382));
    jdff dff_A_kTdAH3H60_0(.din(n1388), .dout(n1385));
    jdff dff_A_ItvWWmwT7_0(.din(n124), .dout(n1388));
    jdff dff_B_Ae8t9VTK3_2(.din(n668), .dout(n1392));
    jdff dff_B_dfkZpVnf5_2(.din(n1392), .dout(n1395));
    jdff dff_B_HHc0DKmb7_2(.din(n1395), .dout(n1398));
    jdff dff_B_1bGkhgnf2_2(.din(n1398), .dout(n1401));
    jdff dff_A_y8WsmTur5_0(.din(n1406), .dout(n1403));
    jdff dff_A_B6YCX7mG2_0(.din(n1409), .dout(n1406));
    jdff dff_A_2feKF3Zk2_0(.din(n1412), .dout(n1409));
    jdff dff_A_FK9RJOmj1_0(.din(n1415), .dout(n1412));
    jdff dff_A_Pwr49xPF5_0(.din(n377), .dout(n1415));
    jdff dff_B_hESeV1NC0_1(.din(n784), .dout(n1419));
    jdff dff_B_LSyfilou3_1(.din(n1419), .dout(n1422));
    jdff dff_B_rl6k19680_1(.din(n1422), .dout(n1425));
    jdff dff_A_dRHQyIA50_1(.din(n584), .dout(n1427));
    jdff dff_A_66PxB4UL7_0(.din(n1433), .dout(n1430));
    jdff dff_A_fBWtJRhz3_0(.din(n1436), .dout(n1433));
    jdff dff_A_zuwmcgl61_0(.din(n1439), .dout(n1436));
    jdff dff_A_ZCoSJqDL0_0(.din(n1442), .dout(n1439));
    jdff dff_A_HPvauYvh8_0(.din(n1445), .dout(n1442));
    jdff dff_A_cxvYa9bb2_0(.din(n584), .dout(n1445));
    jdff dff_A_NDutoFw33_2(.din(n1451), .dout(n1448));
    jdff dff_A_e1EDB06P4_2(.din(n1454), .dout(n1451));
    jdff dff_A_4IkPgO2g2_2(.din(n1457), .dout(n1454));
    jdff dff_A_ZzQbgp3B2_2(.din(n1460), .dout(n1457));
    jdff dff_A_ksU8C2KW5_2(.din(n1463), .dout(n1460));
    jdff dff_A_gCAR8UGY4_2(.din(n584), .dout(n1463));
    jdff dff_A_ykLkWruT0_0(.din(n179), .dout(n1466));
    jdff dff_A_QOKelfPT2_0(.din(n529), .dout(n1469));
    jdff dff_A_JyJpomq77_0(.din(n1475), .dout(n1472));
    jdff dff_A_2i641phh3_0(.din(n1478), .dout(n1475));
    jdff dff_A_YPAYDX9B4_0(.din(n1481), .dout(n1478));
    jdff dff_A_jiBeYxFr6_0(.din(n1484), .dout(n1481));
    jdff dff_A_wddZOLmr2_0(.din(n1487), .dout(n1484));
    jdff dff_A_vQpDA4Vz2_0(.din(n231), .dout(n1487));
    jdff dff_A_7REOox3M7_2(.din(n1493), .dout(n1490));
    jdff dff_A_EJ3WYniq1_2(.din(n1496), .dout(n1493));
    jdff dff_A_qqG1XOGj3_2(.din(n1499), .dout(n1496));
    jdff dff_A_Mwo6TomW6_2(.din(n1502), .dout(n1499));
    jdff dff_A_yYXSBgGe6_2(.din(n1505), .dout(n1502));
    jdff dff_A_ohv5oZ1X2_2(.din(n231), .dout(n1505));
    jdff dff_B_Wmn3ofzU8_0(.din(n195), .dout(n1509));
    jdff dff_A_BlxLJbn71_1(.din(n526), .dout(n1511));
    jdff dff_A_DI3JYTHQ3_0(.din(n1517), .dout(n1514));
    jdff dff_A_Hm5n4ftz9_0(.din(n1520), .dout(n1517));
    jdff dff_A_ipGqDGh94_0(.din(n1523), .dout(n1520));
    jdff dff_A_8HehDjDy2_0(.din(n1526), .dout(n1523));
    jdff dff_A_O9Bze4Dq9_0(.din(n1529), .dout(n1526));
    jdff dff_A_HCBrWaSp5_0(.din(n526), .dout(n1529));
    jdff dff_A_x0x1Am6P9_2(.din(n1535), .dout(n1532));
    jdff dff_A_cSpIwoL75_2(.din(n1538), .dout(n1535));
    jdff dff_A_j6NDuhV37_2(.din(n1541), .dout(n1538));
    jdff dff_A_nhBJw5ZR7_2(.din(n1544), .dout(n1541));
    jdff dff_A_uGMXUnrz9_2(.din(n1547), .dout(n1544));
    jdff dff_A_XhUlaSPc8_2(.din(n526), .dout(n1547));
    jdff dff_A_QKvtC1f67_0(.din(n140), .dout(n1550));
    jdff dff_A_mneKHFDU5_0(.din(n474), .dout(n1553));
    jdff dff_A_4kVdwhdl2_0(.din(n459), .dout(n1556));
    jdff dff_A_sDuJvpTu9_0(.din(n576), .dout(n1559));
    jdff dff_A_e4GOGSkB8_0(.din(n1565), .dout(n1562));
    jdff dff_A_HFfemwmf6_0(.din(n1568), .dout(n1565));
    jdff dff_A_KBcOM4Jl7_0(.din(n1571), .dout(n1568));
    jdff dff_A_shjmP9hR0_0(.din(n1574), .dout(n1571));
    jdff dff_A_ZBVWvipt1_0(.din(n1577), .dout(n1574));
    jdff dff_A_FFGOan2N3_0(.din(n443), .dout(n1577));
    jdff dff_A_PrYQ8vk06_2(.din(n1583), .dout(n1580));
    jdff dff_A_HspB0UhW9_2(.din(n1586), .dout(n1583));
    jdff dff_A_Y6koNCAW7_2(.din(n1589), .dout(n1586));
    jdff dff_A_5bUNF2l39_2(.din(n1592), .dout(n1589));
    jdff dff_A_MRD4AoNy9_2(.din(n1595), .dout(n1592));
    jdff dff_A_uzwkQZ2I5_2(.din(n443), .dout(n1595));
    jdff dff_B_u4RzZMEj3_0(.din(n431), .dout(n1599));
    jdff dff_A_JE9A9tqp1_0(.din(n1604), .dout(n1601));
    jdff dff_A_v3ut1IpA9_0(.din(n1607), .dout(n1604));
    jdff dff_A_CwaotxFj9_0(.din(n1610), .dout(n1607));
    jdff dff_A_JATZXH7W9_0(.din(n1613), .dout(n1610));
    jdff dff_A_KkUIyz2i2_0(.din(n287), .dout(n1613));
    jdff dff_A_QSOiowHf1_1(.din(n251), .dout(n1616));
    jdff dff_A_BFwUrL8z7_0(.din(n1622), .dout(n1619));
    jdff dff_A_zXBYBGc16_0(.din(n1625), .dout(n1622));
    jdff dff_A_iFM7iU6v1_0(.din(n1628), .dout(n1625));
    jdff dff_A_Hxu5YBEq6_0(.din(n1631), .dout(n1628));
    jdff dff_A_kx1wugWw2_0(.din(n1634), .dout(n1631));
    jdff dff_A_VvM6vgff7_0(.din(n1637), .dout(n1634));
    jdff dff_A_r58lH3V02_0(.din(n1640), .dout(n1637));
    jdff dff_A_wCD0Yq4R2_0(.din(n1643), .dout(n1640));
    jdff dff_A_UDu7eOFq7_0(.din(n1646), .dout(n1643));
    jdff dff_A_z1gSDu4R5_0(.din(Gid5), .dout(n1646));
    jdff dff_A_TPnZuobl3_0(.din(n1652), .dout(n1649));
    jdff dff_A_GQByEKuD8_0(.din(n1655), .dout(n1652));
    jdff dff_A_jbxrsE4h6_0(.din(n1658), .dout(n1655));
    jdff dff_A_xMBmPMU74_0(.din(n1661), .dout(n1658));
    jdff dff_A_4xZOwaeg3_0(.din(n1664), .dout(n1661));
    jdff dff_A_lJ1zL3Ms5_0(.din(n1667), .dout(n1664));
    jdff dff_A_9CVvwYn06_0(.din(n1670), .dout(n1667));
    jdff dff_A_KRopvc4R2_0(.din(n1673), .dout(n1670));
    jdff dff_A_M4plUTxg3_0(.din(n1676), .dout(n1673));
    jdff dff_A_P5oWNlu53_0(.din(Gid1), .dout(n1676));
    jdff dff_A_i01bXCXd8_0(.din(n1682), .dout(n1679));
    jdff dff_A_P9mIro7b7_0(.din(n1685), .dout(n1682));
    jdff dff_A_Bz7PX8Da4_0(.din(n1688), .dout(n1685));
    jdff dff_A_AqmayLVM3_0(.din(n1691), .dout(n1688));
    jdff dff_A_FCqsPleW6_0(.din(n1694), .dout(n1691));
    jdff dff_A_HoLhvVbY8_0(.din(n1697), .dout(n1694));
    jdff dff_A_sM694yDn0_0(.din(n1700), .dout(n1697));
    jdff dff_A_oAfJG4058_0(.din(n1703), .dout(n1700));
    jdff dff_A_vPyibuVt2_0(.din(n1706), .dout(n1703));
    jdff dff_A_4gDemzTZ7_0(.din(Gid13), .dout(n1706));
    jdff dff_A_wAzpbYQS3_0(.din(n1712), .dout(n1709));
    jdff dff_A_bFF7kmy35_0(.din(n1715), .dout(n1712));
    jdff dff_A_8NOL1TLa2_0(.din(n1718), .dout(n1715));
    jdff dff_A_NPj9osNJ3_0(.din(n1721), .dout(n1718));
    jdff dff_A_XzXrlRO07_0(.din(n1724), .dout(n1721));
    jdff dff_A_yzRbYqvA2_0(.din(n1727), .dout(n1724));
    jdff dff_A_YnV5BC8T0_0(.din(n1730), .dout(n1727));
    jdff dff_A_Wln0iari3_0(.din(n1733), .dout(n1730));
    jdff dff_A_iQnEU6171_0(.din(n1736), .dout(n1733));
    jdff dff_A_Klm57AT37_0(.din(Gid9), .dout(n1736));
    jdff dff_A_nRbvuv8M9_1(.din(n88), .dout(n1739));
    jdff dff_A_hAVEAOku5_0(.din(n1745), .dout(n1742));
    jdff dff_A_GvIgEcnP9_0(.din(n1748), .dout(n1745));
    jdff dff_A_Te3X00v68_0(.din(n1751), .dout(n1748));
    jdff dff_A_q5Yf0Vyz3_0(.din(n1754), .dout(n1751));
    jdff dff_A_8DPc9Uzb7_0(.din(n1757), .dout(n1754));
    jdff dff_A_wUv7iXPn9_0(.din(n1760), .dout(n1757));
    jdff dff_A_9ubRGCaK3_0(.din(n1763), .dout(n1760));
    jdff dff_A_HABd7t814_0(.din(n1766), .dout(n1763));
    jdff dff_A_x9baV45f4_0(.din(n1769), .dout(n1766));
    jdff dff_A_1r2cNNVA0_0(.din(Gid4), .dout(n1769));
    jdff dff_A_vb3rHJys2_0(.din(n1775), .dout(n1772));
    jdff dff_A_pOuc5m0H8_0(.din(n1778), .dout(n1775));
    jdff dff_A_CtZl4NmD8_0(.din(n1781), .dout(n1778));
    jdff dff_A_D6MRQnTe2_0(.din(n1784), .dout(n1781));
    jdff dff_A_6Tt91TuU1_0(.din(n1787), .dout(n1784));
    jdff dff_A_xqW3bDJy5_0(.din(n1790), .dout(n1787));
    jdff dff_A_KtOsEIdM1_0(.din(n1793), .dout(n1790));
    jdff dff_A_FcfR02qE9_0(.din(n1796), .dout(n1793));
    jdff dff_A_uam4Mvpt2_0(.din(n1799), .dout(n1796));
    jdff dff_A_SMk4Rzs98_0(.din(Gid0), .dout(n1799));
    jdff dff_A_6p8rAL8X3_0(.din(n1805), .dout(n1802));
    jdff dff_A_qBIYq7za9_0(.din(n1808), .dout(n1805));
    jdff dff_A_8LMXLivq2_0(.din(n1811), .dout(n1808));
    jdff dff_A_BFZ4Gl6V7_0(.din(n1814), .dout(n1811));
    jdff dff_A_RYeFefF50_0(.din(n1817), .dout(n1814));
    jdff dff_A_wtKv9GSC0_0(.din(n1820), .dout(n1817));
    jdff dff_A_XoTgZfTW8_0(.din(n1823), .dout(n1820));
    jdff dff_A_N1Saaqg35_0(.din(n1826), .dout(n1823));
    jdff dff_A_gu1ax10V9_0(.din(n1829), .dout(n1826));
    jdff dff_A_9wkS9wKr2_0(.din(Gid12), .dout(n1829));
    jdff dff_A_ducNOe8L5_0(.din(n1835), .dout(n1832));
    jdff dff_A_7D9VR66J9_0(.din(n1838), .dout(n1835));
    jdff dff_A_8WQZR0Lo2_0(.din(n1841), .dout(n1838));
    jdff dff_A_hzTifEEj1_0(.din(n1844), .dout(n1841));
    jdff dff_A_kk0O9RQQ1_0(.din(n1847), .dout(n1844));
    jdff dff_A_IiNwgC7z6_0(.din(n1850), .dout(n1847));
    jdff dff_A_ayfZBSiF5_0(.din(n1853), .dout(n1850));
    jdff dff_A_zCH76v066_0(.din(n1856), .dout(n1853));
    jdff dff_A_skjfGmJy5_0(.din(n1859), .dout(n1856));
    jdff dff_A_lLJru4AI4_0(.din(Gid8), .dout(n1859));
    jdff dff_B_i2QgCSY68_2(.din(n744), .dout(n1863));
    jdff dff_B_nLoB99Yf0_2(.din(n1863), .dout(n1866));
    jdff dff_B_5jl0f5es0_2(.din(n1866), .dout(n1869));
    jdff dff_B_d6TFRYE03_2(.din(n1869), .dout(n1872));
    jdff dff_A_UgUr8UBQ2_0(.din(n1877), .dout(n1874));
    jdff dff_A_9vHPGOCY0_0(.din(n1880), .dout(n1877));
    jdff dff_A_TVdCrnvH6_0(.din(n1883), .dout(n1880));
    jdff dff_A_mLuBbqSX2_0(.din(n1886), .dout(n1883));
    jdff dff_A_6RpvnYwd5_0(.din(n1889), .dout(n1886));
    jdff dff_A_8GFgmSi75_0(.din(n1892), .dout(n1889));
    jdff dff_A_uAOKY6xX6_0(.din(n1895), .dout(n1892));
    jdff dff_A_tVccIOZq0_0(.din(n1898), .dout(n1895));
    jdff dff_A_i68Mpp0q3_0(.din(n1901), .dout(n1898));
    jdff dff_A_5pI5wIum6_0(.din(Gid6), .dout(n1901));
    jdff dff_A_fhfL7ZNh2_0(.din(n1907), .dout(n1904));
    jdff dff_A_QtYcn6H17_0(.din(n1910), .dout(n1907));
    jdff dff_A_N5MTlNjS2_0(.din(n1913), .dout(n1910));
    jdff dff_A_j8fZ2d6n1_0(.din(n1916), .dout(n1913));
    jdff dff_A_8RceGFPk9_0(.din(n1919), .dout(n1916));
    jdff dff_A_Azv9j80w7_0(.din(n1922), .dout(n1919));
    jdff dff_A_ws4PACSk6_0(.din(n1925), .dout(n1922));
    jdff dff_A_5PSOEEr27_0(.din(n1928), .dout(n1925));
    jdff dff_A_g93EImtD5_0(.din(n1931), .dout(n1928));
    jdff dff_A_0SJj0lBu8_0(.din(Gid2), .dout(n1931));
    jdff dff_A_HNuj0yP36_0(.din(n1937), .dout(n1934));
    jdff dff_A_zJqql4ae2_0(.din(n1940), .dout(n1937));
    jdff dff_A_oon9BExA8_0(.din(n1943), .dout(n1940));
    jdff dff_A_kABiU4ks4_0(.din(n1946), .dout(n1943));
    jdff dff_A_qzAnkGuX6_0(.din(n1949), .dout(n1946));
    jdff dff_A_t9UoYn2L6_0(.din(n1952), .dout(n1949));
    jdff dff_A_yLqZb8ab4_0(.din(n1955), .dout(n1952));
    jdff dff_A_f1RmbKaB7_0(.din(n1958), .dout(n1955));
    jdff dff_A_fJL16Qb31_0(.din(n1961), .dout(n1958));
    jdff dff_A_LyMrNUTW1_0(.din(Gid14), .dout(n1961));
    jdff dff_A_Rn5TqlOD3_0(.din(n1967), .dout(n1964));
    jdff dff_A_UWXZGQUD1_0(.din(n1970), .dout(n1967));
    jdff dff_A_KtrV4DP85_0(.din(n1973), .dout(n1970));
    jdff dff_A_tRHN7J6B8_0(.din(n1976), .dout(n1973));
    jdff dff_A_EiyU3HGR1_0(.din(n1979), .dout(n1976));
    jdff dff_A_EWmpaWPZ1_0(.din(n1982), .dout(n1979));
    jdff dff_A_CNgnRqxO1_0(.din(n1985), .dout(n1982));
    jdff dff_A_UOdM8lSR2_0(.din(n1988), .dout(n1985));
    jdff dff_A_rOeqALvP1_0(.din(n1991), .dout(n1988));
    jdff dff_A_wYS3BdfW6_0(.din(Gid10), .dout(n1991));
    jdff dff_A_qFWcYLoC7_0(.din(n1997), .dout(n1994));
    jdff dff_A_JmEtiWwd6_0(.din(n2000), .dout(n1997));
    jdff dff_A_GmVmhRdX0_0(.din(n2003), .dout(n2000));
    jdff dff_A_WJUEV0YA2_0(.din(n2006), .dout(n2003));
    jdff dff_A_maGIHF550_0(.din(n2009), .dout(n2006));
    jdff dff_A_rBrydVzj8_0(.din(n2012), .dout(n2009));
    jdff dff_A_Yi4eIttP4_0(.din(n2015), .dout(n2012));
    jdff dff_A_Ab6nBgXj9_0(.din(n2018), .dout(n2015));
    jdff dff_A_Z9o0sFDI8_0(.din(n2021), .dout(n2018));
    jdff dff_A_GZgjHeOx8_0(.din(n2024), .dout(n2021));
    jdff dff_A_kZnL2V1h6_0(.din(Gid17), .dout(n2024));
    jdff dff_A_lGMmi9g90_0(.din(n2030), .dout(n2027));
    jdff dff_A_BAqnZPKJ8_0(.din(n2033), .dout(n2030));
    jdff dff_A_vJQWoq4r7_0(.din(n2036), .dout(n2033));
    jdff dff_A_hQvNw3Qa3_0(.din(n2039), .dout(n2036));
    jdff dff_A_fsyqxTHM3_0(.din(n2042), .dout(n2039));
    jdff dff_A_PH0OJDwd1_0(.din(n2045), .dout(n2042));
    jdff dff_A_k7y2Wtrb7_0(.din(n2048), .dout(n2045));
    jdff dff_A_nnFGBZ531_0(.din(n2051), .dout(n2048));
    jdff dff_A_R9sJ7BM73_0(.din(n2054), .dout(n2051));
    jdff dff_A_nqcVuyQD6_0(.din(n2057), .dout(n2054));
    jdff dff_A_DJEzk7og9_0(.din(Gid16), .dout(n2057));
    jdff dff_A_F8Vfn9dx4_0(.din(n2063), .dout(n2060));
    jdff dff_A_WKlTuUQc7_0(.din(n2066), .dout(n2063));
    jdff dff_A_QMdbRlZh5_0(.din(n2069), .dout(n2066));
    jdff dff_A_drsbM2rL6_0(.din(n2072), .dout(n2069));
    jdff dff_A_APMNqhGG7_0(.din(n2075), .dout(n2072));
    jdff dff_A_UJlRumnJ0_0(.din(n2078), .dout(n2075));
    jdff dff_A_X69MC0nZ4_0(.din(n2081), .dout(n2078));
    jdff dff_A_Zu7sxXR45_0(.din(n2084), .dout(n2081));
    jdff dff_A_7xihvIPF0_0(.din(n2087), .dout(n2084));
    jdff dff_A_ALfTx6m19_0(.din(n2090), .dout(n2087));
    jdff dff_A_culgjWxi5_0(.din(Gid19), .dout(n2090));
    jdff dff_A_Pr0Wo26f8_0(.din(n2096), .dout(n2093));
    jdff dff_A_BCldgjlb5_0(.din(n2099), .dout(n2096));
    jdff dff_A_zFSxSAr91_0(.din(n2102), .dout(n2099));
    jdff dff_A_qOe9KJQn9_0(.din(n2105), .dout(n2102));
    jdff dff_A_mlIfPHH50_0(.din(n2108), .dout(n2105));
    jdff dff_A_gEQ2B0xt9_0(.din(n2111), .dout(n2108));
    jdff dff_A_vWwtNhQM4_0(.din(n2114), .dout(n2111));
    jdff dff_A_qWKTROdI5_0(.din(n2117), .dout(n2114));
    jdff dff_A_eu05rmxx8_0(.din(n2120), .dout(n2117));
    jdff dff_A_T2YkXJPR8_0(.din(n2123), .dout(n2120));
    jdff dff_A_VQhWYieE2_0(.din(Gid18), .dout(n2123));
    jdff dff_A_9ma5OEpZ6_0(.din(n326), .dout(n2126));
    jdff dff_A_8BagOsUg4_0(.din(n2132), .dout(n2129));
    jdff dff_A_HMtBuOwS0_0(.din(n2135), .dout(n2132));
    jdff dff_A_3k77Rm1d7_0(.din(n2138), .dout(n2135));
    jdff dff_A_Rt1Zs4yD5_0(.din(n2141), .dout(n2138));
    jdff dff_A_R6hLT1gF6_0(.din(n2144), .dout(n2141));
    jdff dff_A_Ee2OX39E3_0(.din(n2147), .dout(n2144));
    jdff dff_A_pMjxcQUz9_0(.din(n2150), .dout(n2147));
    jdff dff_A_JH6rEZM93_0(.din(n2153), .dout(n2150));
    jdff dff_A_Ccze5qj86_0(.din(n2156), .dout(n2153));
    jdff dff_A_LX3bRr914_0(.din(n2159), .dout(n2156));
    jdff dff_A_I8rUbnB55_0(.din(Gid25), .dout(n2159));
    jdff dff_A_hJqy3NvD0_0(.din(n2165), .dout(n2162));
    jdff dff_A_LmhYSz0f9_0(.din(n2168), .dout(n2165));
    jdff dff_A_8M1roRHN0_0(.din(n2171), .dout(n2168));
    jdff dff_A_ER1JIcbh4_0(.din(n2174), .dout(n2171));
    jdff dff_A_zEsPKpjQ5_0(.din(n2177), .dout(n2174));
    jdff dff_A_XhjLBntL7_0(.din(n2180), .dout(n2177));
    jdff dff_A_mL1eZsne1_0(.din(n2183), .dout(n2180));
    jdff dff_A_vA3dOAXc9_0(.din(n2186), .dout(n2183));
    jdff dff_A_kbDH5LK66_0(.din(n2189), .dout(n2186));
    jdff dff_A_1uTknrlB2_0(.din(n2192), .dout(n2189));
    jdff dff_A_JDtv5Dbc7_0(.din(Gid24), .dout(n2192));
    jdff dff_A_hAJX8MYo6_0(.din(n2198), .dout(n2195));
    jdff dff_A_SkR9i0C66_0(.din(n2201), .dout(n2198));
    jdff dff_A_nLTRSfP39_0(.din(n2204), .dout(n2201));
    jdff dff_A_IZAKN65i9_0(.din(n2207), .dout(n2204));
    jdff dff_A_fU09Vo9m5_0(.din(n2210), .dout(n2207));
    jdff dff_A_IKH5coRy4_0(.din(n2213), .dout(n2210));
    jdff dff_A_mNK3ulU47_0(.din(n2216), .dout(n2213));
    jdff dff_A_c2ZlCHke9_0(.din(n2219), .dout(n2216));
    jdff dff_A_AXj4PQA77_0(.din(n2222), .dout(n2219));
    jdff dff_A_bDJzTEBM7_0(.din(n2225), .dout(n2222));
    jdff dff_A_VCEw40Ni6_0(.din(Gid27), .dout(n2225));
    jdff dff_A_4XYts8Ih4_0(.din(n2231), .dout(n2228));
    jdff dff_A_OiQ4UZXn2_0(.din(n2234), .dout(n2231));
    jdff dff_A_GEQXTNG92_0(.din(n2237), .dout(n2234));
    jdff dff_A_TrJ5Ua3e6_0(.din(n2240), .dout(n2237));
    jdff dff_A_gi3HS6BD6_0(.din(n2243), .dout(n2240));
    jdff dff_A_i8cqEZ3d1_0(.din(n2246), .dout(n2243));
    jdff dff_A_y7p6YtTU9_0(.din(n2249), .dout(n2246));
    jdff dff_A_Gbttuphg8_0(.din(n2252), .dout(n2249));
    jdff dff_A_Da0CxEfd3_0(.din(n2255), .dout(n2252));
    jdff dff_A_KCBCdx4k0_0(.din(n2258), .dout(n2255));
    jdff dff_A_TQHmocMZ4_0(.din(Gid26), .dout(n2258));
    jdff dff_A_BNTmMqoF1_0(.din(n2264), .dout(n2261));
    jdff dff_A_54N0ugNR8_0(.din(n2267), .dout(n2264));
    jdff dff_A_YiYD7WbE9_0(.din(n2270), .dout(n2267));
    jdff dff_A_NkiZxHnA9_0(.din(n2273), .dout(n2270));
    jdff dff_A_UsLC33ks8_0(.din(n369), .dout(n2273));
    jdff dff_A_XXhkhR7c0_0(.din(n2279), .dout(n2276));
    jdff dff_A_7qIiETBN5_0(.din(n2282), .dout(n2279));
    jdff dff_A_yCSWFzxC4_0(.din(n2285), .dout(n2282));
    jdff dff_A_z0xVy3rQ8_0(.din(n2288), .dout(n2285));
    jdff dff_A_Fl31Y6cF4_0(.din(n2291), .dout(n2288));
    jdff dff_A_XBN8ZKPt8_0(.din(n2294), .dout(n2291));
    jdff dff_A_hZtC0qdE5_0(.din(n2297), .dout(n2294));
    jdff dff_A_qTZFW09T6_0(.din(n2300), .dout(n2297));
    jdff dff_A_WYgKLuSK9_0(.din(n2303), .dout(n2300));
    jdff dff_A_ipJAZuyO5_0(.din(Gid7), .dout(n2303));
    jdff dff_A_Shhlcgov3_0(.din(n2309), .dout(n2306));
    jdff dff_A_8BknCDYj9_0(.din(n2312), .dout(n2309));
    jdff dff_A_bfr27rka7_0(.din(n2315), .dout(n2312));
    jdff dff_A_t2CEq2bh9_0(.din(n2318), .dout(n2315));
    jdff dff_A_xqUB5j9J1_0(.din(n2321), .dout(n2318));
    jdff dff_A_60zMKwgT3_0(.din(n2324), .dout(n2321));
    jdff dff_A_FYOqB6Jq1_0(.din(n2327), .dout(n2324));
    jdff dff_A_PuMsEJvb8_0(.din(n2330), .dout(n2327));
    jdff dff_A_vupwB64w1_0(.din(n2333), .dout(n2330));
    jdff dff_A_vn5rWJvX4_0(.din(Gid3), .dout(n2333));
    jdff dff_A_L7uZj2Jn7_0(.din(n2339), .dout(n2336));
    jdff dff_A_lG6GjrXS9_0(.din(n2342), .dout(n2339));
    jdff dff_A_7gIX5W2F1_0(.din(n2345), .dout(n2342));
    jdff dff_A_40U1t4ak5_0(.din(n2348), .dout(n2345));
    jdff dff_A_yaObO7Ng2_0(.din(n2351), .dout(n2348));
    jdff dff_A_D0kKTEau4_0(.din(n2354), .dout(n2351));
    jdff dff_A_gQzXy2BT0_0(.din(n2357), .dout(n2354));
endmodule

