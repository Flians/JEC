/*

c3540:
	jxor: 48
	jspl: 222
	jspl3: 321
	jnot: 175
	jcb: 349
	jdff: 1517
	jand: 495

Summary:
	jxor: 48
	jspl: 222
	jspl3: 321
	jnot: 175
	jcb: 349
	jdff: 1517
	jand: 495
*/

module c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G13_0;
	wire [2:0] w_G13_1;
	wire [1:0] w_G13_2;
	wire [2:0] w_G20_0;
	wire [2:0] w_G20_1;
	wire [2:0] w_G20_2;
	wire [2:0] w_G20_3;
	wire [2:0] w_G20_4;
	wire [2:0] w_G20_5;
	wire [2:0] w_G20_6;
	wire [1:0] w_G20_7;
	wire [2:0] w_G33_0;
	wire [2:0] w_G33_1;
	wire [2:0] w_G33_2;
	wire [2:0] w_G33_3;
	wire [2:0] w_G33_4;
	wire [2:0] w_G33_5;
	wire [2:0] w_G33_6;
	wire [2:0] w_G33_7;
	wire [2:0] w_G33_8;
	wire [2:0] w_G33_9;
	wire [2:0] w_G33_10;
	wire [1:0] w_G33_11;
	wire [2:0] w_G41_0;
	wire [2:0] w_G45_0;
	wire [1:0] w_G45_1;
	wire [2:0] w_G50_0;
	wire [2:0] w_G50_1;
	wire [2:0] w_G50_2;
	wire [2:0] w_G50_3;
	wire [2:0] w_G50_4;
	wire [2:0] w_G50_5;
	wire [2:0] w_G50_6;
	wire [2:0] w_G58_0;
	wire [2:0] w_G58_1;
	wire [2:0] w_G58_2;
	wire [2:0] w_G58_3;
	wire [2:0] w_G58_4;
	wire [2:0] w_G58_5;
	wire [2:0] w_G58_6;
	wire [2:0] w_G68_0;
	wire [2:0] w_G68_1;
	wire [2:0] w_G68_2;
	wire [2:0] w_G68_3;
	wire [2:0] w_G68_4;
	wire [2:0] w_G68_5;
	wire [2:0] w_G77_0;
	wire [2:0] w_G77_1;
	wire [2:0] w_G77_2;
	wire [2:0] w_G77_3;
	wire [2:0] w_G77_4;
	wire [2:0] w_G87_0;
	wire [2:0] w_G87_1;
	wire [2:0] w_G87_2;
	wire [2:0] w_G87_3;
	wire [1:0] w_G87_4;
	wire [2:0] w_G97_0;
	wire [2:0] w_G97_1;
	wire [2:0] w_G97_2;
	wire [2:0] w_G97_3;
	wire [2:0] w_G97_4;
	wire [1:0] w_G97_5;
	wire [2:0] w_G107_0;
	wire [2:0] w_G107_1;
	wire [2:0] w_G107_2;
	wire [2:0] w_G107_3;
	wire [2:0] w_G116_0;
	wire [2:0] w_G116_1;
	wire [2:0] w_G116_2;
	wire [2:0] w_G116_3;
	wire [2:0] w_G116_4;
	wire [1:0] w_G116_5;
	wire [1:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G132_0;
	wire [1:0] w_G132_1;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G143_0;
	wire [2:0] w_G143_1;
	wire [1:0] w_G143_2;
	wire [2:0] w_G150_0;
	wire [2:0] w_G150_1;
	wire [2:0] w_G150_2;
	wire [1:0] w_G150_3;
	wire [2:0] w_G159_0;
	wire [2:0] w_G159_1;
	wire [2:0] w_G159_2;
	wire [2:0] w_G159_3;
	wire [2:0] w_G169_0;
	wire [2:0] w_G169_1;
	wire [1:0] w_G169_2;
	wire [2:0] w_G179_0;
	wire [1:0] w_G179_1;
	wire [2:0] w_G190_0;
	wire [2:0] w_G190_1;
	wire [2:0] w_G190_2;
	wire [2:0] w_G190_3;
	wire [2:0] w_G190_4;
	wire [2:0] w_G200_0;
	wire [2:0] w_G200_1;
	wire [1:0] w_G200_2;
	wire [1:0] w_G213_0;
	wire [1:0] w_G223_0;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [2:0] w_G232_0;
	wire [1:0] w_G232_1;
	wire [2:0] w_G238_0;
	wire [1:0] w_G238_1;
	wire [2:0] w_G244_0;
	wire [1:0] w_G244_1;
	wire [2:0] w_G250_0;
	wire [2:0] w_G250_1;
	wire [2:0] w_G257_0;
	wire [1:0] w_G257_1;
	wire [1:0] w_G264_0;
	wire [1:0] w_G270_0;
	wire [2:0] w_G274_0;
	wire [2:0] w_G283_0;
	wire [2:0] w_G283_1;
	wire [2:0] w_G283_2;
	wire [2:0] w_G283_3;
	wire [2:0] w_G294_0;
	wire [2:0] w_G294_1;
	wire [2:0] w_G294_2;
	wire [1:0] w_G294_3;
	wire [2:0] w_G303_0;
	wire [2:0] w_G303_1;
	wire [2:0] w_G303_2;
	wire [2:0] w_G311_0;
	wire [2:0] w_G311_1;
	wire [2:0] w_G317_0;
	wire [1:0] w_G317_1;
	wire [2:0] w_G322_0;
	wire [1:0] w_G326_0;
	wire [2:0] w_G330_0;
	wire [1:0] w_G343_0;
	wire [2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire [1:0] w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire [2:0] w_n73_0;
	wire [1:0] w_n73_1;
	wire [1:0] w_n74_0;
	wire [1:0] w_n75_0;
	wire [2:0] w_n78_0;
	wire [1:0] w_n78_1;
	wire [2:0] w_n79_0;
	wire [1:0] w_n79_1;
	wire [2:0] w_n80_0;
	wire [2:0] w_n80_1;
	wire [2:0] w_n80_2;
	wire [2:0] w_n83_0;
	wire [2:0] w_n84_0;
	wire [1:0] w_n84_1;
	wire [2:0] w_n85_0;
	wire [1:0] w_n85_1;
	wire [1:0] w_n88_0;
	wire [2:0] w_n89_0;
	wire [2:0] w_n90_0;
	wire [2:0] w_n90_1;
	wire [2:0] w_n92_0;
	wire [2:0] w_n94_0;
	wire [1:0] w_n95_0;
	wire [2:0] w_n99_0;
	wire [2:0] w_n99_1;
	wire [2:0] w_n103_0;
	wire [2:0] w_n103_1;
	wire [1:0] w_n104_0;
	wire [2:0] w_n107_0;
	wire [2:0] w_n108_0;
	wire [1:0] w_n108_1;
	wire [1:0] w_n109_0;
	wire [2:0] w_n112_0;
	wire [2:0] w_n112_1;
	wire [1:0] w_n113_0;
	wire [1:0] w_n118_0;
	wire [1:0] w_n127_0;
	wire [1:0] w_n131_0;
	wire [1:0] w_n135_0;
	wire [1:0] w_n138_0;
	wire [2:0] w_n140_0;
	wire [2:0] w_n140_1;
	wire [1:0] w_n141_0;
	wire [2:0] w_n142_0;
	wire [2:0] w_n142_1;
	wire [2:0] w_n142_2;
	wire [2:0] w_n142_3;
	wire [1:0] w_n142_4;
	wire [2:0] w_n143_0;
	wire [2:0] w_n143_1;
	wire [1:0] w_n143_2;
	wire [1:0] w_n144_0;
	wire [2:0] w_n145_0;
	wire [2:0] w_n145_1;
	wire [1:0] w_n145_2;
	wire [2:0] w_n148_0;
	wire [2:0] w_n151_0;
	wire [2:0] w_n151_1;
	wire [2:0] w_n151_2;
	wire [2:0] w_n151_3;
	wire [1:0] w_n151_4;
	wire [1:0] w_n152_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n153_1;
	wire [2:0] w_n153_2;
	wire [2:0] w_n153_3;
	wire [2:0] w_n153_4;
	wire [2:0] w_n153_5;
	wire [2:0] w_n153_6;
	wire [2:0] w_n153_7;
	wire [2:0] w_n153_8;
	wire [1:0] w_n162_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n163_1;
	wire [1:0] w_n165_0;
	wire [2:0] w_n167_0;
	wire [2:0] w_n167_1;
	wire [2:0] w_n167_2;
	wire [2:0] w_n167_3;
	wire [1:0] w_n167_4;
	wire [1:0] w_n168_0;
	wire [2:0] w_n169_0;
	wire [1:0] w_n169_1;
	wire [2:0] w_n170_0;
	wire [2:0] w_n171_0;
	wire [1:0] w_n171_1;
	wire [1:0] w_n172_0;
	wire [2:0] w_n173_0;
	wire [2:0] w_n175_0;
	wire [2:0] w_n175_1;
	wire [2:0] w_n175_2;
	wire [1:0] w_n175_3;
	wire [2:0] w_n176_0;
	wire [2:0] w_n176_1;
	wire [2:0] w_n176_2;
	wire [1:0] w_n176_3;
	wire [1:0] w_n177_0;
	wire [2:0] w_n181_0;
	wire [1:0] w_n181_1;
	wire [1:0] w_n183_0;
	wire [1:0] w_n187_0;
	wire [1:0] w_n189_0;
	wire [2:0] w_n191_0;
	wire [2:0] w_n191_1;
	wire [2:0] w_n191_2;
	wire [2:0] w_n191_3;
	wire [2:0] w_n193_0;
	wire [2:0] w_n199_0;
	wire [1:0] w_n200_0;
	wire [2:0] w_n202_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n208_0;
	wire [1:0] w_n210_0;
	wire [1:0] w_n211_0;
	wire [1:0] w_n214_0;
	wire [2:0] w_n221_0;
	wire [1:0] w_n221_1;
	wire [1:0] w_n223_0;
	wire [1:0] w_n225_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n233_0;
	wire [1:0] w_n234_0;
	wire [2:0] w_n237_0;
	wire [2:0] w_n237_1;
	wire [1:0] w_n243_0;
	wire [2:0] w_n246_0;
	wire [2:0] w_n251_0;
	wire [2:0] w_n251_1;
	wire [2:0] w_n251_2;
	wire [2:0] w_n255_0;
	wire [1:0] w_n255_1;
	wire [2:0] w_n267_0;
	wire [2:0] w_n267_1;
	wire [1:0] w_n268_0;
	wire [1:0] w_n269_0;
	wire [1:0] w_n272_0;
	wire [1:0] w_n275_0;
	wire [2:0] w_n283_0;
	wire [1:0] w_n283_1;
	wire [2:0] w_n284_0;
	wire [2:0] w_n284_1;
	wire [1:0] w_n285_0;
	wire [1:0] w_n289_0;
	wire [1:0] w_n290_0;
	wire [1:0] w_n291_0;
	wire [1:0] w_n292_0;
	wire [1:0] w_n294_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n297_0;
	wire [1:0] w_n298_0;
	wire [1:0] w_n301_0;
	wire [2:0] w_n306_0;
	wire [1:0] w_n306_1;
	wire [1:0] w_n307_0;
	wire [1:0] w_n309_0;
	wire [1:0] w_n312_0;
	wire [2:0] w_n320_0;
	wire [1:0] w_n320_1;
	wire [1:0] w_n321_0;
	wire [2:0] w_n327_0;
	wire [1:0] w_n327_1;
	wire [1:0] w_n330_0;
	wire [1:0] w_n331_0;
	wire [1:0] w_n334_0;
	wire [1:0] w_n335_0;
	wire [1:0] w_n338_0;
	wire [2:0] w_n339_0;
	wire [1:0] w_n339_1;
	wire [1:0] w_n341_0;
	wire [1:0] w_n342_0;
	wire [2:0] w_n350_0;
	wire [1:0] w_n350_1;
	wire [2:0] w_n354_0;
	wire [1:0] w_n354_1;
	wire [1:0] w_n357_0;
	wire [1:0] w_n362_0;
	wire [1:0] w_n364_0;
	wire [1:0] w_n370_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n374_0;
	wire [1:0] w_n375_0;
	wire [2:0] w_n381_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n391_0;
	wire [1:0] w_n391_1;
	wire [1:0] w_n394_0;
	wire [2:0] w_n403_0;
	wire [2:0] w_n406_0;
	wire [1:0] w_n409_0;
	wire [1:0] w_n414_0;
	wire [2:0] w_n415_0;
	wire [1:0] w_n415_1;
	wire [2:0] w_n424_0;
	wire [1:0] w_n424_1;
	wire [1:0] w_n427_0;
	wire [1:0] w_n430_0;
	wire [1:0] w_n436_0;
	wire [2:0] w_n440_0;
	wire [1:0] w_n443_0;
	wire [1:0] w_n448_0;
	wire [1:0] w_n449_0;
	wire [2:0] w_n458_0;
	wire [1:0] w_n458_1;
	wire [1:0] w_n472_0;
	wire [2:0] w_n476_0;
	wire [1:0] w_n478_0;
	wire [1:0] w_n483_0;
	wire [1:0] w_n484_0;
	wire [1:0] w_n486_0;
	wire [2:0] w_n487_0;
	wire [1:0] w_n491_0;
	wire [1:0] w_n497_0;
	wire [1:0] w_n501_0;
	wire [1:0] w_n506_0;
	wire [1:0] w_n510_0;
	wire [1:0] w_n513_0;
	wire [1:0] w_n514_0;
	wire [1:0] w_n520_0;
	wire [1:0] w_n525_0;
	wire [2:0] w_n530_0;
	wire [1:0] w_n530_1;
	wire [2:0] w_n531_0;
	wire [2:0] w_n531_1;
	wire [2:0] w_n531_2;
	wire [2:0] w_n531_3;
	wire [2:0] w_n531_4;
	wire [1:0] w_n533_0;
	wire [1:0] w_n534_0;
	wire [1:0] w_n535_0;
	wire [1:0] w_n537_0;
	wire [2:0] w_n538_0;
	wire [2:0] w_n539_0;
	wire [2:0] w_n541_0;
	wire [2:0] w_n541_1;
	wire [1:0] w_n542_0;
	wire [2:0] w_n544_0;
	wire [2:0] w_n546_0;
	wire [1:0] w_n546_1;
	wire [2:0] w_n559_0;
	wire [2:0] w_n559_1;
	wire [2:0] w_n561_0;
	wire [1:0] w_n561_1;
	wire [2:0] w_n564_0;
	wire [2:0] w_n564_1;
	wire [2:0] w_n565_0;
	wire [2:0] w_n573_0;
	wire [2:0] w_n573_1;
	wire [2:0] w_n574_0;
	wire [2:0] w_n574_1;
	wire [2:0] w_n574_2;
	wire [2:0] w_n574_3;
	wire [1:0] w_n574_4;
	wire [2:0] w_n575_0;
	wire [2:0] w_n578_0;
	wire [2:0] w_n578_1;
	wire [1:0] w_n578_2;
	wire [2:0] w_n579_0;
	wire [2:0] w_n579_1;
	wire [1:0] w_n582_0;
	wire [1:0] w_n583_0;
	wire [2:0] w_n584_0;
	wire [2:0] w_n584_1;
	wire [2:0] w_n584_2;
	wire [2:0] w_n584_3;
	wire [1:0] w_n584_4;
	wire [1:0] w_n585_0;
	wire [2:0] w_n586_0;
	wire [1:0] w_n587_0;
	wire [2:0] w_n588_0;
	wire [2:0] w_n588_1;
	wire [2:0] w_n588_2;
	wire [2:0] w_n588_3;
	wire [2:0] w_n588_4;
	wire [2:0] w_n588_5;
	wire [2:0] w_n588_6;
	wire [1:0] w_n588_7;
	wire [2:0] w_n592_0;
	wire [2:0] w_n592_1;
	wire [2:0] w_n592_2;
	wire [2:0] w_n592_3;
	wire [2:0] w_n592_4;
	wire [2:0] w_n592_5;
	wire [2:0] w_n592_6;
	wire [1:0] w_n592_7;
	wire [2:0] w_n594_0;
	wire [2:0] w_n594_1;
	wire [2:0] w_n594_2;
	wire [2:0] w_n594_3;
	wire [2:0] w_n594_4;
	wire [2:0] w_n594_5;
	wire [1:0] w_n594_6;
	wire [1:0] w_n595_0;
	wire [1:0] w_n597_0;
	wire [2:0] w_n598_0;
	wire [2:0] w_n598_1;
	wire [2:0] w_n598_2;
	wire [2:0] w_n598_3;
	wire [2:0] w_n598_4;
	wire [2:0] w_n598_5;
	wire [2:0] w_n598_6;
	wire [1:0] w_n598_7;
	wire [1:0] w_n600_0;
	wire [1:0] w_n601_0;
	wire [2:0] w_n603_0;
	wire [2:0] w_n603_1;
	wire [2:0] w_n603_2;
	wire [2:0] w_n603_3;
	wire [2:0] w_n603_4;
	wire [2:0] w_n603_5;
	wire [2:0] w_n603_6;
	wire [1:0] w_n603_7;
	wire [2:0] w_n607_0;
	wire [2:0] w_n607_1;
	wire [2:0] w_n607_2;
	wire [2:0] w_n607_3;
	wire [2:0] w_n607_4;
	wire [1:0] w_n607_5;
	wire [1:0] w_n608_0;
	wire [2:0] w_n609_0;
	wire [2:0] w_n609_1;
	wire [2:0] w_n609_2;
	wire [2:0] w_n609_3;
	wire [2:0] w_n609_4;
	wire [2:0] w_n609_5;
	wire [2:0] w_n609_6;
	wire [1:0] w_n609_7;
	wire [2:0] w_n634_0;
	wire [2:0] w_n634_1;
	wire [2:0] w_n634_2;
	wire [2:0] w_n634_3;
	wire [1:0] w_n634_4;
	wire [1:0] w_n637_0;
	wire [2:0] w_n639_0;
	wire [1:0] w_n640_0;
	wire [2:0] w_n645_0;
	wire [1:0] w_n645_1;
	wire [1:0] w_n647_0;
	wire [2:0] w_n658_0;
	wire [2:0] w_n662_0;
	wire [1:0] w_n662_1;
	wire [1:0] w_n674_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n701_0;
	wire [2:0] w_n703_0;
	wire [2:0] w_n714_0;
	wire [1:0] w_n715_0;
	wire [1:0] w_n717_0;
	wire [2:0] w_n718_0;
	wire [2:0] w_n721_0;
	wire [1:0] w_n721_1;
	wire [1:0] w_n725_0;
	wire [1:0] w_n726_0;
	wire [2:0] w_n727_0;
	wire [1:0] w_n729_0;
	wire [1:0] w_n731_0;
	wire [1:0] w_n734_0;
	wire [1:0] w_n738_0;
	wire [2:0] w_n755_0;
	wire [1:0] w_n760_0;
	wire [1:0] w_n764_0;
	wire [1:0] w_n768_0;
	wire [1:0] w_n771_0;
	wire [1:0] w_n778_0;
	wire [1:0] w_n780_0;
	wire [1:0] w_n801_0;
	wire [2:0] w_n810_0;
	wire [1:0] w_n819_0;
	wire [2:0] w_n824_0;
	wire [1:0] w_n825_0;
	wire [2:0] w_n827_0;
	wire [2:0] w_n832_0;
	wire [1:0] w_n834_0;
	wire [1:0] w_n839_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n866_0;
	wire [2:0] w_n897_0;
	wire [1:0] w_n913_0;
	wire [2:0] w_n946_0;
	wire [2:0] w_n948_0;
	wire [2:0] w_n949_0;
	wire [1:0] w_n952_0;
	wire [2:0] w_n961_0;
	wire [1:0] w_n965_0;
	wire [1:0] w_n966_0;
	wire [2:0] w_n1008_0;
	wire [1:0] w_n1011_0;
	wire [1:0] w_n1018_0;
	wire [1:0] w_n1028_0;
	wire [2:0] w_n1065_0;
	wire [2:0] w_n1111_0;
	wire [1:0] w_n1113_0;
	wire [1:0] w_n1114_0;
	wire [1:0] w_n1121_0;
	wire [1:0] w_n1123_0;
	wire [1:0] w_n1124_0;
	wire [1:0] w_n1125_0;
	wire [1:0] w_n1133_0;
	wire [1:0] w_n1134_0;
	wire w_dff_B_r3kRAIpQ2_1;
	wire w_dff_B_jGjlJCd88_1;
	wire w_dff_B_dPcDd7Q30_0;
	wire w_dff_B_bj3H9JTn3_0;
	wire w_dff_B_waQ3RwkB3_0;
	wire w_dff_B_S49LDRpI9_1;
	wire w_dff_B_6QtizgNK7_0;
	wire w_dff_B_NTDd2y4p9_1;
	wire w_dff_B_YpTj6EKW6_1;
	wire w_dff_B_pURHap6Y8_1;
	wire w_dff_B_DClWGZvT8_1;
	wire w_dff_B_Qmhn8zsG1_1;
	wire w_dff_B_lUhdfPXP3_1;
	wire w_dff_B_iBVGmfQV5_1;
	wire w_dff_B_qie6ORYr8_1;
	wire w_dff_B_O822c8kH0_1;
	wire w_dff_B_h8b3xB5Q6_1;
	wire w_dff_B_UrEtn1Rm5_1;
	wire w_dff_B_JycR5cH96_1;
	wire w_dff_B_KZyMGIYv2_1;
	wire w_dff_B_3w172eFQ5_1;
	wire w_dff_B_TL65JbtS7_0;
	wire w_dff_B_r8qjqQ3n3_0;
	wire w_dff_B_OS2rrGMa4_0;
	wire w_dff_B_CbMaE2zY9_0;
	wire w_dff_B_ptaXhLjm1_0;
	wire w_dff_B_jDtbR5Jj2_0;
	wire w_dff_B_N1Ub3KP60_0;
	wire w_dff_B_cCosgA6U3_0;
	wire w_dff_B_8S1vNq1b8_0;
	wire w_dff_B_s8NVsuFV5_0;
	wire w_dff_B_PHJb2qWP2_0;
	wire w_dff_B_Jqbswo0l1_0;
	wire w_dff_B_8R83VQXs5_0;
	wire w_dff_B_ibgIVVWs3_0;
	wire w_dff_B_LYav221B2_0;
	wire w_dff_B_BBx7zaFd7_0;
	wire w_dff_B_ajjuE9LJ1_0;
	wire w_dff_B_7Lk5itsx4_0;
	wire w_dff_B_YFABmYhq7_0;
	wire w_dff_B_1fHMWvHf6_0;
	wire w_dff_B_ATa868hN3_0;
	wire w_dff_B_H9XDiLOP9_0;
	wire w_dff_B_UXJUApCm4_0;
	wire w_dff_B_B7zaxIUB3_0;
	wire w_dff_B_sHpu8Rdi2_0;
	wire w_dff_B_gJEemIMr6_0;
	wire w_dff_B_P2GbtctS6_0;
	wire w_dff_B_UrjTCb297_0;
	wire w_dff_B_Eb7ZkVKn9_0;
	wire w_dff_B_rSUdwkVl7_0;
	wire w_dff_B_LzkS9f5x3_1;
	wire w_dff_B_fX66LWDV4_0;
	wire w_dff_B_DV69GAnb8_1;
	wire w_dff_B_mXpOadW13_1;
	wire w_dff_B_DVIPRSJw1_1;
	wire w_dff_B_CmOGlC6W4_1;
	wire w_dff_B_QBvwxmlc9_1;
	wire w_dff_B_GlkVDUc64_1;
	wire w_dff_B_OerIHMfS6_1;
	wire w_dff_B_I0C8CyNJ4_1;
	wire w_dff_B_BBdJqaQv5_1;
	wire w_dff_B_6nMD3evY1_1;
	wire w_dff_B_sWmRlXx04_1;
	wire w_dff_B_tQ76jetn4_1;
	wire w_dff_B_c8QKqT2q2_1;
	wire w_dff_B_s71eIqgP3_1;
	wire w_dff_B_7wNTkWxA6_1;
	wire w_dff_B_C0KWpf0w3_1;
	wire w_dff_B_kGrMpqO54_0;
	wire w_dff_B_A9hHRejn5_0;
	wire w_dff_B_HxkD4b9J1_0;
	wire w_dff_B_X9idg66l4_0;
	wire w_dff_B_WY3neuGy6_0;
	wire w_dff_B_ADgAvYvc2_0;
	wire w_dff_B_tIvGYJEx6_1;
	wire w_dff_B_9wjLRXn98_0;
	wire w_dff_B_A1EWhcBU9_0;
	wire w_dff_B_yHsBKicb7_1;
	wire w_dff_B_SapRLWNS5_1;
	wire w_dff_B_OWuBgYMA9_1;
	wire w_dff_B_VneAKUWQ0_1;
	wire w_dff_B_ABBEEnfy1_1;
	wire w_dff_A_CQmIbAnm1_1;
	wire w_dff_A_Le8kUKpP8_1;
	wire w_dff_A_DbV8GDW21_1;
	wire w_dff_B_f9ngZ1SD7_0;
	wire w_dff_B_CzT4pdQb5_0;
	wire w_dff_B_R4v33W5T8_0;
	wire w_dff_B_LnBZBnHP3_0;
	wire w_dff_B_qOXUUY664_0;
	wire w_dff_B_14jL4H7C1_0;
	wire w_dff_B_Sg4nGMbq9_0;
	wire w_dff_B_q6OC8l0N7_0;
	wire w_dff_B_HBXTYAzj3_0;
	wire w_dff_B_lGAfzhEC2_0;
	wire w_dff_B_4MFQ0rBK2_0;
	wire w_dff_B_UUZaD1jK0_0;
	wire w_dff_B_dOZtQB3m0_0;
	wire w_dff_B_CIqPzpgN0_0;
	wire w_dff_B_r3jfSRTx8_0;
	wire w_dff_B_gMTsxEsl0_0;
	wire w_dff_B_QpmcwTas3_0;
	wire w_dff_B_wxhLeqir4_0;
	wire w_dff_B_wZ0uvnqf6_0;
	wire w_dff_B_LTeDXujm0_0;
	wire w_dff_B_snArqUtM4_0;
	wire w_dff_B_zP5YUKbg9_0;
	wire w_dff_B_m1rbH33D4_0;
	wire w_dff_B_F7opRmds6_0;
	wire w_dff_B_OqV6vmQM6_1;
	wire w_dff_B_47RNrqGq8_2;
	wire w_dff_B_5Tpf33HU8_2;
	wire w_dff_B_OA7DF1Bj6_2;
	wire w_dff_B_Jgi8miKW4_2;
	wire w_dff_B_5mrVt7GO1_2;
	wire w_dff_B_9EW4iv9v6_2;
	wire w_dff_B_9Aix1DWN2_2;
	wire w_dff_B_nWbrj5Xq9_2;
	wire w_dff_B_L1ggevO54_2;
	wire w_dff_B_uKvOAJjL1_2;
	wire w_dff_B_KGeqL9GY7_2;
	wire w_dff_B_54XVvIGB2_2;
	wire w_dff_B_OKcuJluz3_2;
	wire w_dff_B_sgl3PZ2n2_2;
	wire w_dff_B_RY46vdQ46_2;
	wire w_dff_B_0U4xSHlJ0_2;
	wire w_dff_B_h5tQU98Z2_2;
	wire w_dff_B_jvRKEBnT5_2;
	wire w_dff_B_Dt9CRmEA6_2;
	wire w_dff_B_SYhdm9Wo2_2;
	wire w_dff_B_HwM3TxD34_2;
	wire w_dff_A_uFH8kqJz5_0;
	wire w_dff_A_zPreM2Rj7_0;
	wire w_dff_A_R7m49jkZ5_0;
	wire w_dff_A_CUwa98da6_0;
	wire w_dff_A_c7dW74vt0_0;
	wire w_dff_A_WJqEKpoo6_0;
	wire w_dff_A_ybUbKBm75_0;
	wire w_dff_A_uRkVU4529_0;
	wire w_dff_A_QfGNPeLp2_0;
	wire w_dff_A_j6Lurujp3_0;
	wire w_dff_A_zIbyO1mU6_0;
	wire w_dff_A_xUZBvXgV6_0;
	wire w_dff_A_oKYmP77o2_0;
	wire w_dff_A_t5JRguzs0_0;
	wire w_dff_A_XvidrjEG4_0;
	wire w_dff_A_fTWY8M770_0;
	wire w_dff_A_DbbxjWhF7_0;
	wire w_dff_A_qc4snaze3_0;
	wire w_dff_A_boRgIYP70_0;
	wire w_dff_A_lsCXNBZX3_0;
	wire w_dff_A_3PytOADh8_0;
	wire w_dff_A_QhKTE00P1_0;
	wire w_dff_A_WHOdOuRe0_0;
	wire w_dff_A_ljyVV2Qy8_0;
	wire w_dff_A_dl8KQIxb6_0;
	wire w_dff_A_kQQvnavx6_0;
	wire w_dff_A_w5xjl9lA6_0;
	wire w_dff_A_0Q6EldbN6_1;
	wire w_dff_B_S8WVM1hS3_0;
	wire w_dff_B_UZtwq4PO0_0;
	wire w_dff_B_3GSQrYB29_0;
	wire w_dff_B_mxH9uoAT4_0;
	wire w_dff_B_AXvvbDg23_0;
	wire w_dff_B_RK1iR2RE8_0;
	wire w_dff_B_DTWfMLSi6_0;
	wire w_dff_B_U1ktPB0e7_0;
	wire w_dff_B_WS7OFj0P0_0;
	wire w_dff_B_nKk6nYl89_0;
	wire w_dff_B_vCa5fqnJ1_1;
	wire w_dff_B_i6UbJX2C4_1;
	wire w_dff_B_y37tZ4Lc5_1;
	wire w_dff_B_9HOrcZI27_1;
	wire w_dff_B_Oqeoyf9n3_1;
	wire w_dff_B_zU2R2PzE4_1;
	wire w_dff_B_kC2ssVMQ9_1;
	wire w_dff_B_cWQFdEAc9_1;
	wire w_dff_B_5cZ1O0xr1_0;
	wire w_dff_B_2JA7K7KZ0_0;
	wire w_dff_A_OR4B7QlQ7_1;
	wire w_dff_A_vGyWv8B62_1;
	wire w_dff_A_eUpbv59v7_1;
	wire w_dff_A_pz73L3iA4_1;
	wire w_dff_A_pYr5Q0wG0_1;
	wire w_dff_A_ICV7M9LY9_1;
	wire w_dff_A_K3YCUiXo4_1;
	wire w_dff_A_BfDQ3R3W4_1;
	wire w_dff_A_kwK8aTq29_1;
	wire w_dff_A_Dowq88ls1_1;
	wire w_dff_B_uchyO9Lh0_1;
	wire w_dff_B_edmWya649_1;
	wire w_dff_B_vUDW9NkC7_1;
	wire w_dff_B_EV8IBihK4_1;
	wire w_dff_B_EbJKsm921_1;
	wire w_dff_B_Keavc4sM0_1;
	wire w_dff_A_2kvRam4i1_0;
	wire w_dff_A_Zp6vcKg74_0;
	wire w_dff_B_ElAcdpYs0_2;
	wire w_dff_B_HtTIFEwZ6_2;
	wire w_dff_B_XckPm41r1_1;
	wire w_dff_B_f5m4rwjz6_0;
	wire w_dff_B_smSuVHDx3_0;
	wire w_dff_B_8mjbPghj8_0;
	wire w_dff_B_mBpWAGl59_0;
	wire w_dff_B_BlWMooR57_0;
	wire w_dff_B_s905FG0E6_0;
	wire w_dff_B_IgFdMaRH6_0;
	wire w_dff_B_EGBK8yHP2_0;
	wire w_dff_B_u08wbZlj7_0;
	wire w_dff_B_HvPTZidA6_0;
	wire w_dff_B_bvJN8E9G5_1;
	wire w_dff_B_f35JV3Ep9_2;
	wire w_dff_B_hrXs8Eb47_2;
	wire w_dff_B_3ciWDK0f1_2;
	wire w_dff_B_LciRUnhA4_0;
	wire w_dff_A_dadJwbjL5_1;
	wire w_dff_A_v9rMCZ7a8_1;
	wire w_dff_B_H1vwYt9V7_0;
	wire w_dff_B_vZGGj2Qm5_0;
	wire w_dff_A_gdJhmvkv7_1;
	wire w_dff_A_ADenmync1_1;
	wire w_dff_B_DkZ3iT6Y7_2;
	wire w_dff_B_oCNxCbQi4_2;
	wire w_dff_B_8HkJADyj7_2;
	wire w_dff_B_UeLHqPQg9_0;
	wire w_dff_B_b2BqNUgk9_0;
	wire w_dff_A_EQI4XA034_0;
	wire w_dff_A_5eegF3ti5_0;
	wire w_dff_A_BrlEhjNb0_0;
	wire w_dff_A_097lohcG9_2;
	wire w_dff_A_fYNL4EM06_2;
	wire w_dff_A_ma02ySPw1_2;
	wire w_dff_A_3eRvBS125_2;
	wire w_dff_A_dOiBy7mD3_2;
	wire w_dff_B_kWlhMqib3_0;
	wire w_dff_B_RbEAYj8h2_0;
	wire w_dff_B_58Zn26et7_0;
	wire w_dff_B_5Kh7yM324_0;
	wire w_dff_B_oqr6lieX7_0;
	wire w_dff_B_XBbiO69Z5_0;
	wire w_dff_B_Fu5xcM1d2_0;
	wire w_dff_B_NEbCJ37P3_0;
	wire w_dff_B_U1vlPODo9_0;
	wire w_dff_B_vrgbrAzy6_0;
	wire w_dff_B_M3as2jdR2_0;
	wire w_dff_B_L7D1CmnO6_0;
	wire w_dff_B_vWvobxQE9_1;
	wire w_dff_B_1iIe0ggf8_1;
	wire w_dff_B_mjwmoLdh9_1;
	wire w_dff_B_LkLvAd1X5_0;
	wire w_dff_B_fq1EQPkL3_0;
	wire w_dff_B_Kt8Pkl8Y8_3;
	wire w_dff_B_3snf7RKg4_3;
	wire w_dff_B_LoEDOQo05_3;
	wire w_dff_A_5FM9sSZX4_0;
	wire w_dff_A_2HSi2V1s9_0;
	wire w_dff_A_zBJPXltE3_0;
	wire w_dff_A_JXUbd1bh4_2;
	wire w_dff_A_nfeQYIfl6_2;
	wire w_dff_A_c0hMX5Af4_2;
	wire w_dff_A_PXNzbcOa8_0;
	wire w_dff_A_LngoYsIR5_0;
	wire w_dff_A_gKySxZzv8_0;
	wire w_dff_A_US7ki9f44_0;
	wire w_dff_A_vwztvN8M5_0;
	wire w_dff_A_W8tnGj2F9_0;
	wire w_dff_A_19aJx0qV7_0;
	wire w_dff_A_3HDi1XbW8_1;
	wire w_dff_A_0qUpa6Nl8_1;
	wire w_dff_A_dO770lKP4_1;
	wire w_dff_A_POjjuOXP3_1;
	wire w_dff_A_pcYsestV9_1;
	wire w_dff_B_3DM4Z68X4_3;
	wire w_dff_A_y0rI58hY0_1;
	wire w_dff_A_phUlYsr64_1;
	wire w_dff_A_WYqfzLwj0_1;
	wire w_dff_A_Ohcw8xeW9_1;
	wire w_dff_A_gOIn9MML3_1;
	wire w_dff_A_I5Tqi5Xu2_2;
	wire w_dff_A_os8MM3Za8_2;
	wire w_dff_A_0LaYx7rt6_2;
	wire w_dff_A_nsu0JxYL4_2;
	wire w_dff_A_vR5rV29I9_2;
	wire w_dff_A_wvhqducA2_2;
	wire w_dff_A_MMgmZvqe4_2;
	wire w_dff_A_FxRl3JTB6_0;
	wire w_dff_A_MA0rPdw98_0;
	wire w_dff_A_Zb2QFsoF3_0;
	wire w_dff_A_Dl6pYAmz1_1;
	wire w_dff_A_yaO282oz6_1;
	wire w_dff_A_GhUoLhoJ8_1;
	wire w_dff_A_IsgXaCh32_1;
	wire w_dff_A_9Bk1bKCu0_0;
	wire w_dff_A_QKVqJgMz7_0;
	wire w_dff_A_JU99Oa223_0;
	wire w_dff_A_MRR3uDbp7_0;
	wire w_dff_A_dUpis0yX9_0;
	wire w_dff_A_qj9iYWu55_0;
	wire w_dff_A_miCrs79F0_0;
	wire w_dff_A_6htQD5nO4_0;
	wire w_dff_A_t6jLmTvA9_0;
	wire w_dff_A_ycXKvQzM5_0;
	wire w_dff_A_AFBer5jh7_0;
	wire w_dff_A_gsVQJr0B7_2;
	wire w_dff_A_tBWwSSqg8_2;
	wire w_dff_A_vH9QyFAH4_0;
	wire w_dff_B_OJKARMjA2_1;
	wire w_dff_A_t45hlgsX8_0;
	wire w_dff_A_sS1Clive5_0;
	wire w_dff_A_o8MNwIAq7_1;
	wire w_dff_A_wp8QsmI95_1;
	wire w_dff_A_6qQ0zdwa5_1;
	wire w_dff_A_F8KG0rd27_1;
	wire w_dff_B_JwVbT8Ib5_3;
	wire w_dff_B_AHRCaxL13_3;
	wire w_dff_A_5FAdf8by2_0;
	wire w_dff_A_Ph6wgQJk7_0;
	wire w_dff_A_FNp8w6bp1_0;
	wire w_dff_B_bXb4hhhe3_0;
	wire w_dff_A_vQK9rPe47_0;
	wire w_dff_B_mRGVovu76_1;
	wire w_dff_B_XKI9VZ5k9_1;
	wire w_dff_B_H0JpnCjm0_1;
	wire w_dff_B_2tHWsNiR9_0;
	wire w_dff_A_Hfd7It0H9_1;
	wire w_dff_A_B46Hbzmp1_2;
	wire w_dff_B_R08Ih9bi6_1;
	wire w_dff_B_N05izYLT1_1;
	wire w_dff_B_azvrYdGl8_0;
	wire w_dff_B_2c7q3EWk1_0;
	wire w_dff_A_J1Hp3aej6_0;
	wire w_dff_A_ar5rILi53_0;
	wire w_dff_A_Z4bHatZS4_0;
	wire w_dff_A_WDdd8SeS3_1;
	wire w_dff_A_XYjb7VEd5_1;
	wire w_dff_A_73UYEdBJ2_1;
	wire w_dff_B_8MCw01Rg0_1;
	wire w_dff_A_yDkvygq41_1;
	wire w_dff_B_XI3alUZC5_1;
	wire w_dff_B_wG9g4L8p8_1;
	wire w_dff_B_UU5jplzl4_0;
	wire w_dff_B_AMvP1x4O6_0;
	wire w_dff_B_YoXN2Ew11_0;
	wire w_dff_A_zZbqqVKJ0_0;
	wire w_dff_A_TLdDlbQB2_1;
	wire w_dff_A_3KBrRDM28_1;
	wire w_dff_A_3z5vq90N2_1;
	wire w_dff_B_fCpVejhE2_1;
	wire w_dff_B_dbxYtjsB5_1;
	wire w_dff_B_1i9JVmsm0_1;
	wire w_dff_B_wO9YYGgD8_1;
	wire w_dff_B_GJ5XoSC99_2;
	wire w_dff_B_HboFerw58_2;
	wire w_dff_A_UXK1BWGK5_0;
	wire w_dff_A_WGFVMaPx8_1;
	wire w_dff_A_FW53Yhps1_1;
	wire w_dff_A_akqUpS582_1;
	wire w_dff_B_0I7edd237_1;
	wire w_dff_B_z3fMj7fk0_1;
	wire w_dff_A_3iuqr9z28_0;
	wire w_dff_A_wSx9gRti9_0;
	wire w_dff_A_DS0kuLJX4_0;
	wire w_dff_A_L5ZUWAUW0_0;
	wire w_dff_B_vud1sdUj5_0;
	wire w_dff_B_yWflXVes1_0;
	wire w_dff_B_msIF60Dn0_0;
	wire w_dff_A_FwUPWvLI2_0;
	wire w_dff_A_W2Ki44GS9_1;
	wire w_dff_A_8anq8RjV4_1;
	wire w_dff_A_p26f3lRV2_1;
	wire w_dff_A_W091tQYi5_0;
	wire w_dff_B_b5ePqyXQ6_2;
	wire w_dff_B_kYwFt9Yr7_2;
	wire w_dff_B_btql5Epw5_2;
	wire w_dff_B_gmp3csBQ2_2;
	wire w_dff_B_FZ4kgAJ67_2;
	wire w_dff_B_HLIqN8EU8_2;
	wire w_dff_A_UxchZKH33_1;
	wire w_dff_B_xHpBB69J6_1;
	wire w_dff_B_yE92zG6r5_1;
	wire w_dff_B_UqFtJkCs7_1;
	wire w_dff_A_LJrLFR8L9_0;
	wire w_dff_A_Jwcz2mmN1_0;
	wire w_dff_A_Vr0d0vvE7_0;
	wire w_dff_A_VWO1Fd9K5_2;
	wire w_dff_A_DIwyCqDw2_2;
	wire w_dff_A_5TScZkiy6_1;
	wire w_dff_B_gN2NqprP1_0;
	wire w_dff_B_nM1Ib5xW8_0;
	wire w_dff_B_WXPU0Eer4_0;
	wire w_dff_B_ThjMCZdC7_0;
	wire w_dff_B_lorWBVYy3_0;
	wire w_dff_B_n51VEqSr3_0;
	wire w_dff_A_fDXdL3SA3_0;
	wire w_dff_B_DBRdK7Kn4_3;
	wire w_dff_B_VW85mSJm6_3;
	wire w_dff_B_RxdeFCrb9_3;
	wire w_dff_A_lq1gdekD5_0;
	wire w_dff_A_fzmmIHUK9_0;
	wire w_dff_A_Arvo39BC6_0;
	wire w_dff_A_kHuGlsUy6_0;
	wire w_dff_A_7z3M0q8G9_0;
	wire w_dff_A_XnzcFuZW6_0;
	wire w_dff_A_ptrud9cU5_0;
	wire w_dff_A_yUptmQBo9_1;
	wire w_dff_A_BaDMvh899_1;
	wire w_dff_A_gAyzsRWo3_1;
	wire w_dff_A_6IkSOGA19_1;
	wire w_dff_A_siOXgMss2_1;
	wire w_dff_A_SSDiQdoU2_1;
	wire w_dff_A_P7Rv0l8F9_1;
	wire w_dff_A_afHsN3HE2_1;
	wire w_dff_B_qegTJfwP3_0;
	wire w_dff_B_2VSmEWrt8_0;
	wire w_dff_B_HMjhaAFe1_0;
	wire w_dff_B_yXkkCsrs6_0;
	wire w_dff_A_XWryLDgY7_0;
	wire w_dff_A_qDMZAbvO3_0;
	wire w_dff_A_DoPik7nl2_0;
	wire w_dff_B_2lravuW69_0;
	wire w_dff_B_afLhG7oH1_0;
	wire w_dff_A_zfRA3oVw7_2;
	wire w_dff_A_27yDXbBi6_2;
	wire w_dff_A_41I9nSRK2_1;
	wire w_dff_B_klgUUWDg7_2;
	wire w_dff_B_CwEn7Y6z2_1;
	wire w_dff_B_DXhI0XcQ3_0;
	wire w_dff_A_iOpRD2AB1_1;
	wire w_dff_A_ra2ovdSy7_1;
	wire w_dff_A_XCor1GRt1_1;
	wire w_dff_A_VKlXmtLv3_2;
	wire w_dff_A_n1rNZ6VJ4_2;
	wire w_dff_B_Yxob6LeF8_1;
	wire w_dff_A_xRweCtHC4_1;
	wire w_dff_A_HRH4bXPe7_1;
	wire w_dff_A_gLmHOx7C6_2;
	wire w_dff_A_kXI2QyuQ6_0;
	wire w_dff_B_90XzA1Er2_2;
	wire w_dff_A_zOeZyDd71_2;
	wire w_dff_B_fPnJjukF7_0;
	wire w_dff_B_cjLmZ3eg8_0;
	wire w_dff_A_qKWFEasm0_1;
	wire w_dff_A_WB9p8lUe4_1;
	wire w_dff_A_4kvJkFvK4_1;
	wire w_dff_A_SaZw2CP78_1;
	wire w_dff_B_z6hjKqff5_1;
	wire w_dff_B_BAtwaBZ78_1;
	wire w_dff_B_ZZIZqtV64_1;
	wire w_dff_B_V6zxnBaT1_1;
	wire w_dff_B_Ed9eR1hD6_1;
	wire w_dff_B_JMR7Jm0s6_1;
	wire w_dff_B_Z5oLgYEv9_1;
	wire w_dff_B_WcwNvsPZ5_1;
	wire w_dff_B_d37Ewm1F7_1;
	wire w_dff_B_7ogxw4qH9_1;
	wire w_dff_B_O54W1JxW3_0;
	wire w_dff_B_uQHEYYsw4_0;
	wire w_dff_B_eGPjewSt7_0;
	wire w_dff_B_tNfVI2BL3_0;
	wire w_dff_B_LtshSjJE2_0;
	wire w_dff_B_ALmO11cs1_0;
	wire w_dff_B_ShVlZ9431_1;
	wire w_dff_B_SzLMeSQE7_0;
	wire w_dff_B_QSPc2gnM7_1;
	wire w_dff_B_D5X8rJBq2_0;
	wire w_dff_A_s2WD0Y0I5_0;
	wire w_dff_B_56hO7Xjw7_0;
	wire w_dff_A_EBAejq0L1_2;
	wire w_dff_A_auJTCT6x6_0;
	wire w_dff_A_7qDifxOM7_0;
	wire w_dff_A_BuIzhQVL9_0;
	wire w_dff_A_u1JnJXQ80_0;
	wire w_dff_A_Eh9zIp8q1_1;
	wire w_dff_A_CgbQ7OTl9_1;
	wire w_dff_A_cuvHcPcG3_1;
	wire w_dff_A_JciXvHZn2_1;
	wire w_dff_B_iPrd9TeX5_0;
	wire w_dff_A_vodGdxag8_0;
	wire w_dff_A_f96N0cPC9_0;
	wire w_dff_A_nR4R98C65_1;
	wire w_dff_A_ANdly2E41_1;
	wire w_dff_A_jdBXqUPm7_1;
	wire w_dff_B_hbgj2NQa0_2;
	wire w_dff_B_t1HLMZXK2_2;
	wire w_dff_B_c9IpNzOX5_0;
	wire w_dff_B_7uTgNvTx3_0;
	wire w_dff_B_gZvYO2tJ3_0;
	wire w_dff_B_JZwssl0w9_0;
	wire w_dff_B_6mI38QDp5_0;
	wire w_dff_B_7RaG3MoD4_0;
	wire w_dff_B_erdOwoPR9_0;
	wire w_dff_B_CX9qtM3w1_1;
	wire w_dff_B_3DYUwprA2_1;
	wire w_dff_B_7nbBkGuI5_0;
	wire w_dff_A_XIOaokYB8_0;
	wire w_dff_B_HMDYWvaT5_0;
	wire w_dff_B_nHjT9ivE9_3;
	wire w_dff_B_7jNdzNhw0_3;
	wire w_dff_B_DnzrD0rl8_3;
	wire w_dff_B_2MkF5Ibi1_3;
	wire w_dff_B_FJ0yVpZr8_3;
	wire w_dff_B_zrwlyaUU3_3;
	wire w_dff_A_Th4JHEbi6_0;
	wire w_dff_A_nSuweLyS0_0;
	wire w_dff_A_BLmq1XbH5_1;
	wire w_dff_A_Ih9jq9Sa3_1;
	wire w_dff_A_2ylipEtU7_0;
	wire w_dff_B_gj7NzOOx8_1;
	wire w_dff_B_gyCkCVW80_0;
	wire w_dff_A_1oitqJRV5_1;
	wire w_dff_A_7RI8VtIk1_1;
	wire w_dff_A_l6PcCziw9_1;
	wire w_dff_A_hlWLWior1_1;
	wire w_dff_B_Tgc52uHY7_0;
	wire w_dff_B_bZqFMHI27_0;
	wire w_dff_B_rqhWIE9n5_1;
	wire w_dff_B_v658yW0u7_1;
	wire w_dff_B_iYrA9RZ57_1;
	wire w_dff_B_lJMPZ3y32_0;
	wire w_dff_A_tV0FgGOD4_1;
	wire w_dff_A_MxRcqYg14_1;
	wire w_dff_A_5OB9D1s01_1;
	wire w_dff_B_QHGupD9O5_0;
	wire w_dff_B_CYKxdWpc3_0;
	wire w_dff_B_7FoqHNTg6_0;
	wire w_dff_B_enwv1RSk2_0;
	wire w_dff_B_fRfLC7wP3_0;
	wire w_dff_B_naovNozt1_0;
	wire w_dff_B_kSPUY3b25_0;
	wire w_dff_B_30CLogu30_0;
	wire w_dff_B_nyCuQUXp5_0;
	wire w_dff_B_popybWGT3_0;
	wire w_dff_B_EoVue6r71_0;
	wire w_dff_B_uVYZmFoa2_0;
	wire w_dff_B_jUyMRLqf9_1;
	wire w_dff_B_HxXAlIrC8_1;
	wire w_dff_B_6QpDm6ob6_1;
	wire w_dff_B_ELOV9xVH7_1;
	wire w_dff_B_1OG4qX6U7_1;
	wire w_dff_B_LlUIFToS7_1;
	wire w_dff_B_Fc1BDKqS9_0;
	wire w_dff_B_F3XZmJmq0_0;
	wire w_dff_B_rVv7XDPP0_0;
	wire w_dff_A_lKgum9Dc3_0;
	wire w_dff_A_M2LnEw7Y9_0;
	wire w_dff_A_Zv3tUhWl4_1;
	wire w_dff_A_zFPCULDU7_1;
	wire w_dff_A_5amnptMJ8_1;
	wire w_dff_A_9QSiTYBb6_1;
	wire w_dff_A_LPCp8wUi4_1;
	wire w_dff_B_FmJuE4933_0;
	wire w_dff_B_zJiB3lEY7_0;
	wire w_dff_B_YqXng1Tl4_0;
	wire w_dff_A_DaGiIoEz7_1;
	wire w_dff_B_Cvdy09qm7_0;
	wire w_dff_A_ILbNzyuE6_1;
	wire w_dff_A_TNYJ7iBL0_1;
	wire w_dff_A_XQmfFHEB3_1;
	wire w_dff_A_PHS2RXKV3_2;
	wire w_dff_A_bXd2SWAe9_2;
	wire w_dff_A_LX63CiXg6_0;
	wire w_dff_A_MFW7rTmx9_0;
	wire w_dff_A_CqdVymKg8_1;
	wire w_dff_A_Pw3VdEjM4_1;
	wire w_dff_A_zIsp6HRb7_2;
	wire w_dff_A_6cENp0FW9_2;
	wire w_dff_A_bgcYkwPV5_2;
	wire w_dff_A_c577wqMH2_1;
	wire w_dff_A_5RTE3ISJ7_1;
	wire w_dff_A_nZ7gWBPL1_1;
	wire w_dff_A_guwEpJeY9_0;
	wire w_dff_A_nvKubPcz8_1;
	wire w_dff_B_tyhBi3LE7_3;
	wire w_dff_B_KH0k5irM5_3;
	wire w_dff_A_TkmKvSnH5_0;
	wire w_dff_A_6rWT0e2E1_0;
	wire w_dff_A_4OZnzc347_1;
	wire w_dff_A_3PFdd2zu2_1;
	wire w_dff_A_tdhUzLrN3_0;
	wire w_dff_A_ksnOaavp9_0;
	wire w_dff_A_3vO6REX67_0;
	wire w_dff_A_LHtDBGoa3_1;
	wire w_dff_A_J0e7aXRe2_1;
	wire w_dff_A_VhN3Y8XQ5_1;
	wire w_dff_A_dSupes7L3_1;
	wire w_dff_A_Vs8BAEzk3_1;
	wire w_dff_A_NipjuKUi1_1;
	wire w_dff_A_FC3MZrhx5_2;
	wire w_dff_A_v9gX4OE79_2;
	wire w_dff_A_AlWz1lJ56_2;
	wire w_dff_A_kcHBLyaI9_0;
	wire w_dff_A_3YfeII840_2;
	wire w_dff_A_X8XzmPe39_2;
	wire w_dff_A_e2PL1fzF4_2;
	wire w_dff_A_BwHLonLY8_2;
	wire w_dff_A_XN7tJbQv3_2;
	wire w_dff_A_9dFVMJ195_2;
	wire w_dff_A_kdVNOwJ95_2;
	wire w_dff_A_jnql4Twp1_1;
	wire w_dff_A_Dz2EHSEq0_0;
	wire w_dff_A_zofU3MdX8_0;
	wire w_dff_A_NmVd0pp08_0;
	wire w_dff_A_m2v9p7Rr3_0;
	wire w_dff_A_a0n21v4d7_0;
	wire w_dff_A_KRynQWo53_0;
	wire w_dff_A_vlFA9Oth2_0;
	wire w_dff_A_M5l0UahZ2_0;
	wire w_dff_A_IDNEl2ZS0_0;
	wire w_dff_A_bD87Onbr9_0;
	wire w_dff_A_dAgqKiCL4_0;
	wire w_dff_A_Mb1QoJJ16_0;
	wire w_dff_A_XxpKgWzr6_1;
	wire w_dff_A_qouqHV0E4_1;
	wire w_dff_A_XJ1WFJjT2_1;
	wire w_dff_A_SAOtFZLC4_1;
	wire w_dff_A_IQ4shD001_1;
	wire w_dff_A_nQyxS2Ra9_1;
	wire w_dff_B_nuLMXo2V1_1;
	wire w_dff_B_8Xb02A4E5_1;
	wire w_dff_B_w0igAweX8_1;
	wire w_dff_B_m2KEuw7G7_1;
	wire w_dff_A_sOt7iCiN6_0;
	wire w_dff_B_a9Bq9Jbt6_0;
	wire w_dff_B_92Xyjyt49_0;
	wire w_dff_A_HP1SQecO2_0;
	wire w_dff_A_IrqUSM7k7_0;
	wire w_dff_A_7LwcJ7e83_0;
	wire w_dff_A_uDBMBd6j5_0;
	wire w_dff_A_8ak2UWrj6_0;
	wire w_dff_B_weVp08Pp5_2;
	wire w_dff_B_irG8Eo2N2_2;
	wire w_dff_B_2sX8viCE6_1;
	wire w_dff_B_K5kPQRym6_1;
	wire w_dff_B_a3L0F4cM6_1;
	wire w_dff_B_Xsx7zUaF5_1;
	wire w_dff_B_jqYBxtNK9_1;
	wire w_dff_B_WHMoBw497_1;
	wire w_dff_B_SW1uqonc9_0;
	wire w_dff_A_u1iOwQ3o1_2;
	wire w_dff_A_7LZyPDqT9_1;
	wire w_dff_A_ATjqoJSG6_1;
	wire w_dff_A_nKpt3kIN3_1;
	wire w_dff_A_OuUDbJ9h6_1;
	wire w_dff_A_iHzsrRMf2_1;
	wire w_dff_A_dFeogwBV2_1;
	wire w_dff_A_koRkDfe93_1;
	wire w_dff_A_v45iXzmy9_1;
	wire w_dff_A_DuVn1rsK2_1;
	wire w_dff_A_qRSk5vFg3_1;
	wire w_dff_A_WWbyJ8n71_1;
	wire w_dff_A_HUiclmJB9_2;
	wire w_dff_A_Lqffpbav6_2;
	wire w_dff_A_TiiSdpQG7_2;
	wire w_dff_A_YEyTH6s70_2;
	wire w_dff_A_rFwZtK179_2;
	wire w_dff_A_OOnSfLez6_2;
	wire w_dff_A_aIFlGAtg5_2;
	wire w_dff_A_0o0f1lf62_2;
	wire w_dff_B_1BNxiPH74_1;
	wire w_dff_B_zK9Y8eAx8_1;
	wire w_dff_B_PXQbvnM88_1;
	wire w_dff_A_kzR7u1TD1_1;
	wire w_dff_B_yOM4cw0L7_1;
	wire w_dff_B_VxFm5xip0_0;
	wire w_dff_A_2W7L7zYy3_0;
	wire w_dff_A_rXfHdOZq3_0;
	wire w_dff_A_Lvok6WBq7_0;
	wire w_dff_A_7KWpzyRE0_1;
	wire w_dff_A_0ZhmkXJ00_1;
	wire w_dff_A_gWN7ECOm3_2;
	wire w_dff_A_gmDsf9ec5_2;
	wire w_dff_A_kYJkszQe9_2;
	wire w_dff_A_ex4bYEwq2_1;
	wire w_dff_B_IOoAVviH4_2;
	wire w_dff_B_MNhyYSQm0_0;
	wire w_dff_A_dpknuFx02_1;
	wire w_dff_A_6nQF6u7s9_1;
	wire w_dff_A_nuUKsgjt7_0;
	wire w_dff_A_bMVuxE5G0_0;
	wire w_dff_A_ZHa1CROU4_0;
	wire w_dff_A_GXpsoGnT9_0;
	wire w_dff_A_h3ncExe39_1;
	wire w_dff_B_xlKVheb49_0;
	wire w_dff_A_WQyxfCM38_1;
	wire w_dff_A_DZ7VIiJY5_1;
	wire w_dff_A_s5KBHbYF5_1;
	wire w_dff_A_t5mJqnh39_2;
	wire w_dff_A_F51UaCPE1_2;
	wire w_dff_A_Vt7nZ2km2_2;
	wire w_dff_A_efSbgbCQ2_1;
	wire w_dff_B_bsd1qens3_2;
	wire w_dff_B_Fvc9IbLX9_2;
	wire w_dff_A_Tg48kJFf3_0;
	wire w_dff_A_GgI2SKKZ4_0;
	wire w_dff_A_VYQW2B8n1_2;
	wire w_dff_B_6hZTUKfw7_0;
	wire w_dff_A_mBQNp16G1_1;
	wire w_dff_A_qI8LMykU9_0;
	wire w_dff_A_Ivahdf7R9_1;
	wire w_dff_A_NyYRzj6E9_1;
	wire w_dff_A_1NcBMjnV7_1;
	wire w_dff_B_BZ4DsGxm4_0;
	wire w_dff_A_Rc1cOJEn9_0;
	wire w_dff_B_Su4cP8Us5_0;
	wire w_dff_A_xdO5RVy33_0;
	wire w_dff_A_SLgBHqgl5_1;
	wire w_dff_B_qdGSDyRC3_1;
	wire w_dff_A_Jq39jHdr6_0;
	wire w_dff_A_4ZkRuOox8_0;
	wire w_dff_A_Jb85nn0H4_2;
	wire w_dff_B_NMpI85nN2_1;
	wire w_dff_B_lLNwMGRH2_0;
	wire w_dff_B_yxtZg7tQ0_0;
	wire w_dff_B_EiP3ThKA5_0;
	wire w_dff_B_52PmUoso1_0;
	wire w_dff_A_2YVx9pA02_0;
	wire w_dff_A_3qsiCGA71_0;
	wire w_dff_A_GoKqyPRw1_2;
	wire w_dff_A_ak5WnuVE9_0;
	wire w_dff_B_ak8NJgpB3_2;
	wire w_dff_B_vu9Wbdxq9_1;
	wire w_dff_B_nOF57Ihc9_0;
	wire w_dff_A_7yVOR6bZ8_1;
	wire w_dff_A_Z4RwFHax0_2;
	wire w_dff_A_1pEbSX8l2_0;
	wire w_dff_A_ER2hJ8O59_0;
	wire w_dff_A_n87Vl5Io4_1;
	wire w_dff_A_6dK1w0MQ3_1;
	wire w_dff_A_B6Vs1lec3_1;
	wire w_dff_A_deBmJCFF2_2;
	wire w_dff_A_zd486uqH3_2;
	wire w_dff_A_3hxgHbCD4_1;
	wire w_dff_A_hh55e6nh0_1;
	wire w_dff_A_5F61E4JD0_1;
	wire w_dff_A_KjkG0oBM0_2;
	wire w_dff_A_agEXFetD7_2;
	wire w_dff_A_et9S8n2w5_0;
	wire w_dff_A_au7JGJKz5_0;
	wire w_dff_A_nyLEkgiy9_0;
	wire w_dff_B_RTHaLB9P4_2;
	wire w_dff_A_USzALghU5_0;
	wire w_dff_A_TDDQKBda6_0;
	wire w_dff_A_zupOeHI68_0;
	wire w_dff_A_pFE1Frdz6_0;
	wire w_dff_A_OppAy5Zf5_0;
	wire w_dff_A_XN6l2aJN6_1;
	wire w_dff_A_S99EpfW01_1;
	wire w_dff_A_Y5gNh7m69_1;
	wire w_dff_B_zkwCK5Dw6_0;
	wire w_dff_A_IgTa6ZNf1_1;
	wire w_dff_A_sqJjZZ9z9_0;
	wire w_dff_A_ghJ8wUVE0_2;
	wire w_dff_A_HN76owjW0_2;
	wire w_dff_A_2xUdHjSB5_2;
	wire w_dff_A_f28f5INd7_2;
	wire w_dff_B_w13kkr5n3_3;
	wire w_dff_B_DuujXMuX4_3;
	wire w_dff_B_6JNF1BfV2_3;
	wire w_dff_B_mQ5ZAuB85_3;
	wire w_dff_A_8lR3zUvc4_1;
	wire w_dff_A_W7gmO0gB4_1;
	wire w_dff_A_prKTJLcj5_1;
	wire w_dff_A_6IsqXu5a7_2;
	wire w_dff_A_dK2rfGwR3_2;
	wire w_dff_B_s1MZ71WS2_0;
	wire w_dff_B_Sc8WFc9M4_0;
	wire w_dff_B_witi1zg83_0;
	wire w_dff_B_MMoY9aKr6_0;
	wire w_dff_A_nnK8K6Yd5_1;
	wire w_dff_A_jEkaSazK0_1;
	wire w_dff_B_OlWs8Heb2_0;
	wire w_dff_A_Y6eoVmlR8_1;
	wire w_dff_A_WgCxRYDW1_1;
	wire w_dff_A_vUBv06Fc3_2;
	wire w_dff_A_RfNyO60m7_0;
	wire w_dff_A_2kHRESU46_0;
	wire w_dff_A_9jfPiPj04_2;
	wire w_dff_A_GsXmotwF4_2;
	wire w_dff_B_QtalDuBA3_0;
	wire w_dff_A_5cPOZy7q5_0;
	wire w_dff_B_K7Pdc8mo9_1;
	wire w_dff_A_ZvC7meZE3_1;
	wire w_dff_A_hzv3AJbH0_1;
	wire w_dff_A_Z9sZP4ti6_1;
	wire w_dff_A_K5fo6cxL0_1;
	wire w_dff_A_aAnbTL744_2;
	wire w_dff_A_SPflITre2_0;
	wire w_dff_B_IluYWD2B6_2;
	wire w_dff_A_bERrxIDg1_0;
	wire w_dff_A_zXkfapMO8_1;
	wire w_dff_A_iXH7P5d46_1;
	wire w_dff_A_tGIwWPc98_0;
	wire w_dff_A_x836GCzJ0_0;
	wire w_dff_A_yLyYwaU37_0;
	wire w_dff_A_5AF34kqV1_2;
	wire w_dff_A_54pfsnNL9_2;
	wire w_dff_B_Bas7vXo25_1;
	wire w_dff_B_oLqY92ZG7_1;
	wire w_dff_B_WafiYv6g5_0;
	wire w_dff_A_Xkk2p6Kp8_2;
	wire w_dff_A_oTrsiTn54_0;
	wire w_dff_A_4itEZmO81_0;
	wire w_dff_A_8SbsIMPh6_1;
	wire w_dff_A_EnmipDdM3_1;
	wire w_dff_A_yuQOSCFe1_2;
	wire w_dff_A_It1b8Apm1_2;
	wire w_dff_A_NYiak4bQ0_2;
	wire w_dff_A_d4neQDxl2_0;
	wire w_dff_A_Mguwjh3Y5_0;
	wire w_dff_A_xPlFSzND5_0;
	wire w_dff_A_J8Xrpnru1_0;
	wire w_dff_A_MfTlVsaB8_2;
	wire w_dff_A_8sSiV2zs4_1;
	wire w_dff_A_GzGL9BU06_1;
	wire w_dff_A_6ynn85cg3_1;
	wire w_dff_A_3raSrlKE7_1;
	wire w_dff_A_NingPJJr5_0;
	wire w_dff_A_FrefPK8O5_0;
	wire w_dff_A_THdACRsx7_0;
	wire w_dff_A_zihQz6gZ9_0;
	wire w_dff_A_5No72I6T6_0;
	wire w_dff_A_L227eugT4_0;
	wire w_dff_A_8YmVFp8d9_2;
	wire w_dff_B_k3R0GRDO1_1;
	wire w_dff_B_9AtbX24Q1_0;
	wire w_dff_B_bqSrjtx16_0;
	wire w_dff_B_aPDOq9fw2_0;
	wire w_dff_B_tiVVBsFY0_1;
	wire w_dff_B_0vRxV8tn7_1;
	wire w_dff_B_zJLrF8qo5_1;
	wire w_dff_B_vNQOvYjL3_1;
	wire w_dff_B_BkPSlq8z9_0;
	wire w_dff_B_Y9mIcjJJ2_0;
	wire w_dff_A_9DOAq5WU0_0;
	wire w_dff_A_Yp6EBFDp7_0;
	wire w_dff_B_JxW6VFUK4_2;
	wire w_dff_A_ytxfUw0E9_2;
	wire w_dff_A_p1wf4wwP0_2;
	wire w_dff_A_iMa7f0N08_2;
	wire w_dff_A_Uxiv7mDf4_1;
	wire w_dff_A_KOPMjFeF6_1;
	wire w_dff_A_DUwZdRKu2_1;
	wire w_dff_A_ml3cqTxh8_1;
	wire w_dff_A_sucufshR2_1;
	wire w_dff_A_47GHoTMv4_1;
	wire w_dff_A_ERpOTMRg7_1;
	wire w_dff_A_YZd3ftvQ7_1;
	wire w_dff_A_AosIMfix1_2;
	wire w_dff_A_lt8TWJel9_2;
	wire w_dff_A_vEhoGedL2_2;
	wire w_dff_B_3ZrYfTLl2_1;
	wire w_dff_B_7cKiESw98_1;
	wire w_dff_B_coLmqX0w8_1;
	wire w_dff_B_3i0omfmu0_1;
	wire w_dff_B_EJaLm2yo5_0;
	wire w_dff_B_Cv0jdZhY0_0;
	wire w_dff_B_frWjfpCC8_0;
	wire w_dff_A_HGiHmRHa9_1;
	wire w_dff_A_YssGkI0D9_1;
	wire w_dff_A_Q6r6O0Ff9_1;
	wire w_dff_A_q76h1Grp0_1;
	wire w_dff_A_ZNWPlGT61_0;
	wire w_dff_A_L324XXoF0_1;
	wire w_dff_A_wDEjfRe06_1;
	wire w_dff_A_nLvSUpGX2_1;
	wire w_dff_A_6zURVSFX1_2;
	wire w_dff_A_BuFQ7ENo7_2;
	wire w_dff_A_NtRs0Lns7_2;
	wire w_dff_A_ZUAPrBEK6_0;
	wire w_dff_A_b9GROpJW2_0;
	wire w_dff_A_G2slVSIU2_1;
	wire w_dff_A_O14BRBRi1_0;
	wire w_dff_A_4Ip61xn62_1;
	wire w_dff_A_P2k1ZYb97_1;
	wire w_dff_A_VcM5NMVd3_1;
	wire w_dff_A_9mcLTUWd1_1;
	wire w_dff_A_8wdWQmrJ2_1;
	wire w_dff_A_x3cqZVrK0_1;
	wire w_dff_A_mwQXrT2J4_1;
	wire w_dff_A_qC7rVrwi6_1;
	wire w_dff_A_QqpC6r7Z8_2;
	wire w_dff_A_HH7vxqTT1_2;
	wire w_dff_A_NpB3G7Bq5_0;
	wire w_dff_A_lavui2pd4_1;
	wire w_dff_A_nZFqLcox7_1;
	wire w_dff_A_qcS1sfZV7_0;
	wire w_dff_A_AdIubfXa6_0;
	wire w_dff_A_OO7uJMLQ3_2;
	wire w_dff_B_4Gh0fwtc9_2;
	wire w_dff_B_856zJ3iP1_2;
	wire w_dff_B_C9KSGfsQ0_2;
	wire w_dff_B_EO90XBws6_3;
	wire w_dff_B_aWlbAKyW4_3;
	wire w_dff_B_pIQiSaGZ0_3;
	wire w_dff_B_Ty1SYtPV1_3;
	wire w_dff_B_mXNucLYp9_3;
	wire w_dff_B_Pa74sO4r2_3;
	wire w_dff_B_Zcm9hBc21_1;
	wire w_dff_B_JVJHfrUM2_1;
	wire w_dff_B_GXaL3ZsG0_1;
	wire w_dff_A_g0CTxuN66_0;
	wire w_dff_A_WkIZ9Ipi3_0;
	wire w_dff_A_QktPgrCA7_0;
	wire w_dff_A_35I4PX3a1_0;
	wire w_dff_A_LjQXjsAQ4_0;
	wire w_dff_A_g8b3qWfZ8_0;
	wire w_dff_A_b02XpM220_1;
	wire w_dff_A_ZvST1GIK2_1;
	wire w_dff_A_qeqK6uzc8_1;
	wire w_dff_B_5lXSsvLL5_3;
	wire w_dff_B_JUdPVsRX7_3;
	wire w_dff_B_kZ0fZPgi3_3;
	wire w_dff_A_OqvBEi9O5_0;
	wire w_dff_A_EDjJCaEM3_0;
	wire w_dff_A_9xqjFTvx0_0;
	wire w_dff_A_6QIZpNEc4_2;
	wire w_dff_A_hMiY208a9_2;
	wire w_dff_A_iUBzaUNc4_2;
	wire w_dff_A_5hCaIDoL6_1;
	wire w_dff_A_WW8we5c08_0;
	wire w_dff_A_Npus9YKO8_0;
	wire w_dff_A_FhAe9Zg75_0;
	wire w_dff_A_cuGTOmQg6_1;
	wire w_dff_A_Oa27SE9W4_1;
	wire w_dff_A_fXEdsmQ75_1;
	wire w_dff_A_iKTNXKZc3_0;
	wire w_dff_A_tikgggIb4_0;
	wire w_dff_A_69Qogbok1_1;
	wire w_dff_A_uCZnG92N2_0;
	wire w_dff_A_ynTVZFdy6_1;
	wire w_dff_B_8VStsy0h7_3;
	wire w_dff_B_6tq39FvZ8_3;
	wire w_dff_A_VWmwSnvD7_0;
	wire w_dff_A_d4tngxdW3_0;
	wire w_dff_A_LSZJC3xa5_0;
	wire w_dff_A_0WdZJnEe2_0;
	wire w_dff_A_fXfdB0lU2_1;
	wire w_dff_A_9mtb9rSS4_1;
	wire w_dff_A_yQd0I7028_1;
	wire w_dff_A_ZOM03yNy5_1;
	wire w_dff_A_iNETUz0D5_0;
	wire w_dff_A_NqtSGlXd4_1;
	wire w_dff_A_mESEmxt54_0;
	wire w_dff_A_T0huWdzQ2_0;
	wire w_dff_A_k3uNQ6l93_1;
	wire w_dff_A_Y8g8JBsj4_0;
	wire w_dff_A_hRrX8oGS5_1;
	wire w_dff_A_YfqCN7g38_1;
	wire w_dff_A_Cb6U7dYo9_1;
	wire w_dff_A_SY8jVMB27_1;
	wire w_dff_A_fMQD3J5V6_1;
	wire w_dff_A_zPbPefOx5_2;
	wire w_dff_A_c26WNJs30_2;
	wire w_dff_A_XB9u5wBA3_2;
	wire w_dff_A_WQ9NFfDz5_1;
	wire w_dff_A_tK2tHP670_1;
	wire w_dff_A_YC9e3UYf0_1;
	wire w_dff_A_tz4ezU1Z1_2;
	wire w_dff_A_qt1oHG395_2;
	wire w_dff_A_wyqwC8n39_2;
	wire w_dff_A_zc5L4iXU9_1;
	wire w_dff_A_w10T9dZ60_1;
	wire w_dff_A_OKTHj1IG9_1;
	wire w_dff_A_ybXPjCr49_2;
	wire w_dff_A_x1ZLCVR54_2;
	wire w_dff_A_7IDlMxKm4_2;
	wire w_dff_A_UhOdz5az7_2;
	wire w_dff_A_3YOwGcrz0_2;
	wire w_dff_A_XteHk1YD6_2;
	wire w_dff_A_OoJdkKVT5_1;
	wire w_dff_A_V3ZYA3xF7_1;
	wire w_dff_A_WATa9lbd5_1;
	wire w_dff_A_ca7ACg321_1;
	wire w_dff_A_PiKjDvWl7_1;
	wire w_dff_A_RsJcQgEB6_1;
	wire w_dff_A_0wkcZKDD1_2;
	wire w_dff_A_vETwgtEH4_2;
	wire w_dff_A_5AcsddxH0_2;
	wire w_dff_A_z83nPjcq3_2;
	wire w_dff_A_Eme40qrN6_2;
	wire w_dff_A_BHi2T2dg0_2;
	wire w_dff_A_xIcLbesx1_1;
	wire w_dff_A_Ue9sukoG5_1;
	wire w_dff_A_3LU1iai92_1;
	wire w_dff_A_XEtSx5NJ2_1;
	wire w_dff_A_CLNDS7V07_1;
	wire w_dff_A_KTSnkItS2_2;
	wire w_dff_A_F1j5wBK80_2;
	wire w_dff_A_OH7CtWHC1_2;
	wire w_dff_A_BxkjGqqB8_2;
	wire w_dff_A_vh7UCrih5_2;
	wire w_dff_A_CKJkWGGl9_2;
	wire w_dff_A_1TN1V6Zt4_2;
	wire w_dff_A_0sn6RaSv1_0;
	wire w_dff_A_XlLw9ZLW4_1;
	wire w_dff_A_t19azNHw0_0;
	wire w_dff_A_5B2x4W2w6_0;
	wire w_dff_A_CwrNi5cu0_0;
	wire w_dff_A_QWWvgvKW9_1;
	wire w_dff_A_2mcTbHyJ7_1;
	wire w_dff_A_AeYLXE9H6_1;
	wire w_dff_A_Mt88KHO83_0;
	wire w_dff_A_1wDiKAeu7_0;
	wire w_dff_A_0V8mqk7o9_1;
	wire w_dff_A_uVpjaaK94_1;
	wire w_dff_A_czSiPcGG6_1;
	wire w_dff_A_HEG50RAb2_0;
	wire w_dff_A_d4tqvVTr0_0;
	wire w_dff_A_hsbDY3rh5_0;
	wire w_dff_A_xFE0W88I6_1;
	wire w_dff_A_PouHlUSh2_1;
	wire w_dff_A_Earr44st9_1;
	wire w_dff_A_U81WuUBA8_0;
	wire w_dff_A_kPdL6L0q5_0;
	wire w_dff_A_a4bonOBI8_0;
	wire w_dff_A_6lhPNLrv1_0;
	wire w_dff_A_iV1NPdKu0_0;
	wire w_dff_A_iH1O1xLw5_0;
	wire w_dff_A_YQ8M2Mcf1_0;
	wire w_dff_A_UrjXRtc59_2;
	wire w_dff_A_cAOo0EWf3_2;
	wire w_dff_A_dKytGgwp2_2;
	wire w_dff_A_eNB2q96Y2_2;
	wire w_dff_A_LSMCeX8K1_2;
	wire w_dff_A_zJh6XiLg1_2;
	wire w_dff_A_epqVj9Gl4_2;
	wire w_dff_A_Sf5n20R13_2;
	wire w_dff_A_3OQCcMXd8_1;
	wire w_dff_A_29Z0gz3k4_1;
	wire w_dff_A_0TjFo9LS7_1;
	wire w_dff_A_QNqpnw0L2_1;
	wire w_dff_A_TiC7mZPB2_1;
	wire w_dff_A_JQ5IT0bb7_1;
	wire w_dff_A_uDlIdtm69_1;
	wire w_dff_A_OqOZjD7v9_1;
	wire w_dff_A_Tc0cGRKe8_1;
	wire w_dff_A_7WM1I46y6_2;
	wire w_dff_A_oOwsZbF53_2;
	wire w_dff_A_gXxOmiAh1_2;
	wire w_dff_A_isXvbwmC7_2;
	wire w_dff_A_YEKzohOc6_2;
	wire w_dff_A_ypt91aZp8_2;
	wire w_dff_A_3VbCZcko9_2;
	wire w_dff_A_vQcL9gd23_0;
	wire w_dff_A_7ODBYoAU0_0;
	wire w_dff_A_aJkDY9jT9_0;
	wire w_dff_A_xoPW5xzo0_0;
	wire w_dff_A_1VmBzJMq9_0;
	wire w_dff_A_KNWpJ1814_0;
	wire w_dff_A_ognYgis48_0;
	wire w_dff_A_qoKVMUri9_0;
	wire w_dff_A_FK04W79i4_0;
	wire w_dff_A_JILh3T5A3_2;
	wire w_dff_A_Rb6AHIed4_2;
	wire w_dff_A_0jl5l4hp5_2;
	wire w_dff_A_6MEQgBni0_2;
	wire w_dff_A_ymmBDbG78_2;
	wire w_dff_A_dH2z5x6g4_2;
	wire w_dff_A_DbuiHhS49_2;
	wire w_dff_A_Kh0W7LJm7_0;
	wire w_dff_A_9qTpjvg52_0;
	wire w_dff_A_BrtoE2Cx9_1;
	wire w_dff_A_RzBvpja00_1;
	wire w_dff_A_8PiacHDd5_1;
	wire w_dff_A_SpgKQ8sL4_0;
	wire w_dff_A_9cZizQgL7_0;
	wire w_dff_A_la4Lg7iy3_0;
	wire w_dff_B_8219FGGN1_0;
	wire w_dff_B_qv6ztYWL1_0;
	wire w_dff_A_fAgM6g8M2_2;
	wire w_dff_A_N4SXkTLS6_2;
	wire w_dff_A_2jLXFuQv9_2;
	wire w_dff_A_KAwmpeJO5_1;
	wire w_dff_A_bDA0GVVs0_1;
	wire w_dff_A_9E02IJP68_2;
	wire w_dff_A_BllAhk3v7_1;
	wire w_dff_A_Jx4UkCvz0_1;
	wire w_dff_A_lSEecwiY4_1;
	wire w_dff_A_4gOG3Ltk0_2;
	wire w_dff_A_zi7A3axm0_0;
	wire w_dff_A_xDdIks2k5_0;
	wire w_dff_A_YLiZrEYK7_0;
	wire w_dff_A_HbCePM388_0;
	wire w_dff_A_f3NzufjE0_0;
	wire w_dff_A_9S3vw8Ew3_0;
	wire w_dff_A_VpS1disS9_1;
	wire w_dff_A_XWODCJk37_1;
	wire w_dff_A_hkOcqSpi0_1;
	wire w_dff_A_f9fPes1r4_1;
	wire w_dff_A_KPYgOAhA6_2;
	wire w_dff_A_SDOExKsY0_2;
	wire w_dff_A_tc25riLF0_2;
	wire w_dff_A_emKsr4Fg6_2;
	wire w_dff_A_0tYGGUoq8_1;
	wire w_dff_A_j1hc41OV4_1;
	wire w_dff_A_paEEYKD64_1;
	wire w_dff_B_t80UjEDy7_2;
	wire w_dff_A_xfzRTbUX5_1;
	wire w_dff_A_Cc185wxx8_1;
	wire w_dff_A_QKpOV3Co8_1;
	wire w_dff_B_lZ0KuJ4o5_1;
	wire w_dff_B_Di3rUeFI3_1;
	wire w_dff_A_Y8hYC2IV0_1;
	wire w_dff_A_RA89g64K2_1;
	wire w_dff_A_DnLvpEAF5_1;
	wire w_dff_A_xIPSMYqF5_1;
	wire w_dff_A_x5iny7C70_1;
	wire w_dff_A_hRzyRzXw2_1;
	wire w_dff_A_AZKHoWiQ4_2;
	wire w_dff_A_36D7eIJr5_2;
	wire w_dff_A_Yym9ARtr7_2;
	wire w_dff_A_Q8nlyQ1Z4_2;
	wire w_dff_A_xYaBeaJI4_2;
	wire w_dff_A_gwt26j987_2;
	wire w_dff_A_a5fQVTzg2_2;
	wire w_dff_A_eNK4R6Wc2_1;
	wire w_dff_A_9znQbK8K4_1;
	wire w_dff_A_Pjipn1Bh4_2;
	wire w_dff_A_VnHop4lI8_2;
	wire w_dff_A_YReyY20D5_1;
	wire w_dff_A_zFoFmfc91_1;
	wire w_dff_A_HA43TPzI4_2;
	wire w_dff_A_cVCIdqAS5_2;
	wire w_dff_A_fEYszTsu9_2;
	wire w_dff_A_YCFcJsKT1_2;
	wire w_dff_A_pvLVCwaM3_2;
	wire w_dff_A_3eBytgpX4_1;
	wire w_dff_A_3usa37dt1_1;
	wire w_dff_A_e0xAzYEy0_1;
	wire w_dff_A_Byv1Yxey2_1;
	wire w_dff_A_yDQKd7iq0_1;
	wire w_dff_A_AdX3ri1D4_1;
	wire w_dff_A_8rPchjsM9_2;
	wire w_dff_A_qvasqyZf6_1;
	wire w_dff_A_ABYWI6VE8_1;
	wire w_dff_A_fvx1FcJL2_1;
	wire w_dff_A_0ywe8Y0j3_0;
	wire w_dff_B_gF9WsJ4t1_0;
	wire w_dff_A_hSILwcqq7_2;
	wire w_dff_A_fj4txxlY0_0;
	wire w_dff_A_czs1bfAp0_2;
	wire w_dff_A_XCdy0zIb4_0;
	wire w_dff_A_0IZjeug70_0;
	wire w_dff_A_zyKZmBA41_0;
	wire w_dff_A_v5J5apna9_1;
	wire w_dff_A_DV6vWHAV8_1;
	wire w_dff_A_yfwxKucK7_1;
	wire w_dff_A_aqfcMpWq8_1;
	wire w_dff_A_KpbIBopu1_1;
	wire w_dff_A_VCMu02xU2_2;
	wire w_dff_A_CTDjGbnj1_2;
	wire w_dff_A_GKRYpEuA5_2;
	wire w_dff_A_DSBvx0Ah3_2;
	wire w_dff_A_JS0tIAsY3_0;
	wire w_dff_A_dzOtopaT8_0;
	wire w_dff_A_drWM7Ylr6_0;
	wire w_dff_A_hPZj13FQ6_0;
	wire w_dff_A_0wL0cO0E4_2;
	wire w_dff_A_fe3aKREo2_2;
	wire w_dff_A_KMDWpFI76_2;
	wire w_dff_A_I11MkcQE4_2;
	wire w_dff_A_1ehwWKnk4_2;
	wire w_dff_A_1pMPP5rW9_2;
	wire w_dff_A_0S5FIjkv8_1;
	wire w_dff_A_KO3ZZ86d4_1;
	wire w_dff_A_RJv6eMpf7_0;
	wire w_dff_A_7GZeRR1V0_0;
	wire w_dff_A_L1LfM2zG9_0;
	wire w_dff_A_fOVcn0cu7_1;
	wire w_dff_B_h7yKL39l2_0;
	wire w_dff_B_DAC8bilL0_3;
	wire w_dff_A_jDCWKkcP8_1;
	wire w_dff_A_VzEBntKb0_1;
	wire w_dff_A_uivRfVn56_1;
	wire w_dff_A_g5fnT28m4_1;
	wire w_dff_A_5LXrVV437_2;
	wire w_dff_A_1ZCCUhkB4_2;
	wire w_dff_A_oQN1rgso3_0;
	wire w_dff_A_rJTuoJ295_0;
	wire w_dff_A_zIemMhgn9_0;
	wire w_dff_A_IMmRtMZE4_1;
	wire w_dff_A_FG0ioKLT5_1;
	wire w_dff_A_WRB8si7u2_1;
	wire w_dff_A_XPicNu6b4_0;
	wire w_dff_A_ynPFlVee7_0;
	wire w_dff_A_u9ZGdr624_0;
	wire w_dff_A_oYsg2RoG3_2;
	wire w_dff_A_iH77Os1e9_2;
	wire w_dff_A_gHd0RMZ40_2;
	wire w_dff_A_w31GkA329_0;
	wire w_dff_A_Jh9CEhWh9_0;
	wire w_dff_A_iBXhMxwh8_2;
	wire w_dff_A_t7bk5ory4_0;
	wire w_dff_A_c1JWmLH73_0;
	wire w_dff_A_qWmm4XBe9_1;
	wire w_dff_A_JyVyhI943_1;
	wire w_dff_A_B5Q1wpPz9_1;
	wire w_dff_A_vatFgBln0_1;
	wire w_dff_A_Aj3lUnKW1_0;
	wire w_dff_A_VrttsOYA9_2;
	wire w_dff_A_kQnQgSOO9_2;
	wire w_dff_A_s8fqRlFn4_1;
	wire w_dff_A_2myHAoyQ6_0;
	wire w_dff_A_1Du0ZaHl4_0;
	wire w_dff_A_oyhlAvoM2_0;
	wire w_dff_A_Mwwm7nIY8_0;
	wire w_dff_A_Uz9cwlyk5_0;
	wire w_dff_A_7Wmj5fAf5_0;
	wire w_dff_A_eBfeswso1_0;
	wire w_dff_A_U6vvSeoE1_0;
	wire w_dff_A_SyUTfx7y4_0;
	wire w_dff_A_dH9Yogdq5_0;
	wire w_dff_A_CDWKKud07_0;
	wire w_dff_A_EdceNqbx6_0;
	wire w_dff_A_XgFv67y14_0;
	wire w_dff_A_0sdUi2d00_0;
	wire w_dff_A_ucWjFwd26_0;
	wire w_dff_A_s2Qb03pe3_0;
	wire w_dff_A_3ismzyuC2_0;
	wire w_dff_A_ByMvWYW64_1;
	wire w_dff_A_JElLs7Gx3_1;
	wire w_dff_B_rwldEtvG9_1;
	wire w_dff_B_JapuFSpL8_1;
	wire w_dff_A_9J1j9XG43_0;
	wire w_dff_A_THLLKRTA2_0;
	wire w_dff_A_UOhAl3AG6_0;
	wire w_dff_A_L3IOk9wr4_1;
	wire w_dff_A_hXLqg86h2_1;
	wire w_dff_A_iP9w2g1g0_1;
	wire w_dff_A_Wjps8uhV2_1;
	wire w_dff_A_rWES0KiL5_1;
	wire w_dff_A_NWQxB7k92_1;
	wire w_dff_A_kIGrJzaO2_1;
	wire w_dff_A_01IyBm3r8_2;
	wire w_dff_B_os1UX2Uh9_3;
	wire w_dff_B_zd5dVfUd6_3;
	wire w_dff_B_K5rKf5gl6_3;
	wire w_dff_B_988m3ij01_3;
	wire w_dff_A_lbKQYAN26_0;
	wire w_dff_A_t4aTUrN55_0;
	wire w_dff_A_enyAnlgb9_0;
	wire w_dff_A_MBfHdSgu8_0;
	wire w_dff_A_ce9dhZGO4_0;
	wire w_dff_A_jIv7nspd0_0;
	wire w_dff_A_7bDZaXzh3_0;
	wire w_dff_A_v7mod6Fz3_0;
	wire w_dff_A_YQABj98p0_0;
	wire w_dff_A_Nhg0tDvh7_0;
	wire w_dff_A_cKU9WJCE0_0;
	wire w_dff_A_OacZVhaD0_2;
	wire w_dff_A_Tjp1h7dN3_1;
	wire w_dff_A_s1ptZKpM2_1;
	wire w_dff_B_9wQpPHUb9_1;
	wire w_dff_B_wuSjxGMb3_1;
	wire w_dff_B_aUzpgTQD2_1;
	wire w_dff_B_saO59Fmz8_1;
	wire w_dff_A_Tqry09g46_0;
	wire w_dff_A_ZSDab67S5_0;
	wire w_dff_A_vV64sr3w8_0;
	wire w_dff_A_0DUZvNbg9_0;
	wire w_dff_A_XTGG9y8x7_2;
	wire w_dff_A_qP9inbNF1_2;
	wire w_dff_A_9ud1mzav9_2;
	wire w_dff_A_Xa25Z2Up3_2;
	wire w_dff_A_cSHrJns84_1;
	wire w_dff_A_jSiJcNSL3_1;
	wire w_dff_A_HDfvmbSy5_1;
	wire w_dff_A_VwcYS28T1_2;
	wire w_dff_A_OdCd76oN4_2;
	wire w_dff_A_skgac2vk4_2;
	wire w_dff_A_6aYC8LGG7_2;
	wire w_dff_A_WntodRxc7_2;
	wire w_dff_A_An85pV1v5_2;
	wire w_dff_A_DytGePDb4_1;
	wire w_dff_A_6WaQmQZx7_0;
	wire w_dff_A_Fha37d1V2_0;
	wire w_dff_A_OgmqfJ9Y9_0;
	wire w_dff_A_zBAtWpy87_1;
	wire w_dff_A_t7ycE5da5_1;
	wire w_dff_A_japh8m6f2_1;
	wire w_dff_A_BNN3rqAD9_0;
	wire w_dff_A_kWk1fZDO7_0;
	wire w_dff_A_Z4gpDrdV4_0;
	wire w_dff_A_Y6N4dNAR7_1;
	wire w_dff_A_9WKlBnfF9_1;
	wire w_dff_A_6Nv8glqm8_1;
	wire w_dff_A_Ytt10nUx2_0;
	wire w_dff_A_kOWn8T0U2_0;
	wire w_dff_A_Y7vdIFIK6_1;
	wire w_dff_A_si3cUgSf0_0;
	wire w_dff_A_A4rf8QyB8_0;
	wire w_dff_A_FEZpIib27_0;
	wire w_dff_B_jviK8z9P0_0;
	wire w_dff_A_qTqAcC4z7_2;
	wire w_dff_A_xBj5cX0X9_2;
	wire w_dff_A_PneygkG64_0;
	wire w_dff_A_RsTLAMxA9_1;
	wire w_dff_A_L8RaPNdA8_0;
	wire w_dff_A_OTVES8wK6_1;
	wire w_dff_A_Gvez15wZ2_2;
	wire w_dff_A_ym6S5rR28_2;
	wire w_dff_A_0lhVdymT3_2;
	wire w_dff_A_L7ZuTVMZ3_2;
	wire w_dff_A_1AiiHIgY1_0;
	wire w_dff_A_R7XW4HVH1_1;
	wire w_dff_A_MlDAFvhn9_2;
	wire w_dff_A_DzYTHKxa5_0;
	wire w_dff_A_QxIYbuhb7_0;
	wire w_dff_A_QvlrAJJ99_1;
	wire w_dff_A_kfyvtHr53_0;
	wire w_dff_A_J6dLmODg2_0;
	wire w_dff_A_JBh6SnlL3_1;
	wire w_dff_A_wQiY8xZZ6_1;
	wire w_dff_A_6jGnGUuh6_1;
	wire w_dff_A_4AZOtCLP3_1;
	wire w_dff_A_P28HTxyQ2_1;
	wire w_dff_A_ueunDt7R6_2;
	wire w_dff_A_iOyGJcSv8_2;
	wire w_dff_A_AYHq6CK15_0;
	wire w_dff_A_uFxFIb6L8_2;
	wire w_dff_A_vFeSx1O01_2;
	wire w_dff_A_7r9CT32r7_2;
	wire w_dff_A_HIJ7ju3t0_1;
	wire w_dff_A_qs52CrPS9_1;
	wire w_dff_A_Nsl13udB4_1;
	wire w_dff_A_UT885Zls5_2;
	wire w_dff_A_HWqYXczf8_2;
	wire w_dff_A_399Kevc33_2;
	wire w_dff_A_hFnmCp9o6_1;
	wire w_dff_A_yhCoLZdL9_1;
	wire w_dff_B_HpxBCUdY2_3;
	wire w_dff_B_VuWeNsBL3_3;
	wire w_dff_B_hkgUZhFI7_3;
	wire w_dff_B_LS61dqx66_3;
	wire w_dff_B_tXsgcTSw2_3;
	wire w_dff_B_BwWvCrM99_3;
	wire w_dff_B_YlrImd1e3_3;
	wire w_dff_B_qR0nOs1x3_3;
	wire w_dff_B_OEg4m9xA1_3;
	wire w_dff_B_ZhZ4D0zS4_3;
	wire w_dff_B_0dXxVJuE3_3;
	wire w_dff_B_hWTaQiHW1_3;
	wire w_dff_A_wq17tauH8_1;
	wire w_dff_A_odPI4HrQ6_1;
	wire w_dff_A_eq5YLhq75_1;
	wire w_dff_A_o6mjsxuy0_1;
	wire w_dff_A_8QnkC18e8_1;
	wire w_dff_A_ChNSborp8_1;
	wire w_dff_A_G3muGB1A2_1;
	wire w_dff_A_PJflLZpI6_1;
	wire w_dff_A_LK58E5yq2_1;
	wire w_dff_A_HcC95OHT5_2;
	wire w_dff_A_bRIPMCeQ2_2;
	wire w_dff_A_BSCoWUSj4_2;
	wire w_dff_A_2i7L6yMM1_2;
	wire w_dff_A_LkQJ7Yen8_2;
	wire w_dff_A_4bcMFsIz0_2;
	wire w_dff_A_FwqPq3SO6_0;
	wire w_dff_A_MIMMLezA6_0;
	wire w_dff_A_n4OUThTi6_0;
	wire w_dff_A_8ENOy4QH8_0;
	wire w_dff_A_xbKGV8NW7_0;
	wire w_dff_A_U62r0qJs5_0;
	wire w_dff_A_2xtU7aLo1_0;
	wire w_dff_A_kMWFvHvv5_0;
	wire w_dff_A_6HVwM8yu0_1;
	wire w_dff_A_3dyDH51V9_1;
	wire w_dff_A_NrhTesYA0_1;
	wire w_dff_A_T7h3xX7x7_1;
	wire w_dff_A_qUZtGVCA1_1;
	wire w_dff_A_EI3WYb5P3_1;
	wire w_dff_A_j6WSIunK5_2;
	wire w_dff_A_1ySQcKkI4_2;
	wire w_dff_A_xlQbREQG7_2;
	wire w_dff_A_wT7z0BGQ2_2;
	wire w_dff_A_LshbYJWD0_2;
	wire w_dff_A_dsPI1f6d0_2;
	wire w_dff_A_CjqlpFYP9_2;
	wire w_dff_A_bull1NsZ7_2;
	wire w_dff_A_bGLM5hDN8_2;
	wire w_dff_A_XhX0mBD51_2;
	wire w_dff_A_IBtBOk9U7_2;
	wire w_dff_A_O9lR93Wb3_2;
	wire w_dff_A_Z1wyCwtZ5_2;
	wire w_dff_A_1AnaTcwN1_2;
	wire w_dff_A_rntIr00f0_2;
	wire w_dff_A_Jf5yIcVn3_0;
	wire w_dff_A_wb0wzZSE9_0;
	wire w_dff_A_jKgZNIMu7_0;
	wire w_dff_A_xDPBuZb37_0;
	wire w_dff_A_ZISYk3go7_0;
	wire w_dff_A_0ZTjpXni3_0;
	wire w_dff_A_8lkKjvOA5_0;
	wire w_dff_A_xnnJk6NX3_0;
	wire w_dff_A_F8Wh3OG13_0;
	wire w_dff_A_O9Hvuued7_0;
	wire w_dff_A_qLPUx0zY9_0;
	wire w_dff_A_JAjcmLmg2_0;
	wire w_dff_A_UdbYpxOn5_0;
	wire w_dff_A_jR0uzgHd6_1;
	wire w_dff_A_fP9zkEzN6_1;
	wire w_dff_A_28pLuohY1_1;
	wire w_dff_A_Z6I2cObm2_1;
	wire w_dff_A_qNisaUU57_1;
	wire w_dff_A_Q5cVGGPa3_1;
	wire w_dff_A_8X2wSEvH9_1;
	wire w_dff_A_LSBen3VT6_1;
	wire w_dff_A_IKY4WGqU3_1;
	wire w_dff_A_eZTnycEY0_1;
	wire w_dff_A_PwS40WEr4_1;
	wire w_dff_A_suiCb5en8_1;
	wire w_dff_A_PKBNQTrc3_1;
	wire w_dff_A_Zj2o4NDI8_1;
	wire w_dff_A_LSVW6T4U5_1;
	wire w_dff_A_QMz9OikZ6_1;
	wire w_dff_A_KWPFfSFI3_1;
	wire w_dff_A_sepS8pSO6_1;
	wire w_dff_A_NaxjPiNG0_1;
	wire w_dff_A_qtlOBJgE6_1;
	wire w_dff_A_rYEg0xQW4_1;
	wire w_dff_A_CQ9if87m6_1;
	wire w_dff_A_DervnNSt4_1;
	wire w_dff_A_GFjYngmS2_1;
	wire w_dff_A_KCXX7tRl7_1;
	wire w_dff_A_6P2bOYnB9_1;
	wire w_dff_A_C8D6vxpD9_2;
	wire w_dff_A_Vt8mm9Rn7_2;
	wire w_dff_A_v9RSeGlc2_2;
	wire w_dff_A_8AiQklu46_2;
	wire w_dff_A_duFtBtYo7_2;
	wire w_dff_A_jyxrqg485_2;
	wire w_dff_A_HHn99T6W3_2;
	wire w_dff_A_rBNz9LNg5_2;
	wire w_dff_A_WrHiGEOx6_2;
	wire w_dff_A_JV2OWS1j2_2;
	wire w_dff_A_KPaBokur1_2;
	wire w_dff_A_QtGdZ2P71_2;
	wire w_dff_A_QsyBmHKn1_2;
	wire w_dff_A_oF0G75GT9_2;
	wire w_dff_B_TbB8LnBB0_3;
	wire w_dff_B_Sj4KfGWI2_0;
	wire w_dff_A_NINlQxwq3_1;
	wire w_dff_A_NwbguLHv3_1;
	wire w_dff_A_kC2B1HrP3_1;
	wire w_dff_A_S0swvLc28_0;
	wire w_dff_A_V2sEVFqm3_0;
	wire w_dff_A_4DbpvSP54_0;
	wire w_dff_A_jyntGYM43_0;
	wire w_dff_A_n5LQbdfq2_0;
	wire w_dff_A_c25JhkaE2_0;
	wire w_dff_A_vVl1w5EO7_0;
	wire w_dff_A_ZxSMuo5S0_0;
	wire w_dff_A_GpSmMdZv1_0;
	wire w_dff_A_T185TyPJ9_0;
	wire w_dff_A_6ThDI6n79_0;
	wire w_dff_A_2Z5DWBrz8_0;
	wire w_dff_A_TUeKvJNr8_0;
	wire w_dff_A_HHOYeyMC1_0;
	wire w_dff_A_qIOZQG3K4_0;
	wire w_dff_A_yZfjNgZR7_0;
	wire w_dff_A_k1RkcxC58_1;
	wire w_dff_A_5iromuUB8_1;
	wire w_dff_A_Eplzsdje0_1;
	wire w_dff_A_D6wIkQq63_1;
	wire w_dff_A_dvKQ3T2E6_1;
	wire w_dff_A_3OvbDbXf2_1;
	wire w_dff_A_0ku9FXH22_1;
	wire w_dff_A_l9l4KR9Q6_1;
	wire w_dff_A_3C2r4G7N4_1;
	wire w_dff_A_fgjGIS8G1_1;
	wire w_dff_A_zyTKAbuF7_1;
	wire w_dff_A_Bcu0894d5_1;
	wire w_dff_A_QUJzufsG6_1;
	wire w_dff_A_oX0tGj6o2_1;
	wire w_dff_A_Q3oncG7x6_2;
	wire w_dff_A_WCpF15mb9_2;
	wire w_dff_A_siDBz2mL7_2;
	wire w_dff_A_sibQJt2b4_2;
	wire w_dff_A_4hiLJwyr0_2;
	wire w_dff_A_C1RyuKyV3_2;
	wire w_dff_A_rqsCTgRs1_2;
	wire w_dff_A_ShMnqvVX2_2;
	wire w_dff_A_38seGSQL2_2;
	wire w_dff_A_uRrYSUoL8_2;
	wire w_dff_A_21Sx4Cu24_2;
	wire w_dff_A_86ZLDcDD8_2;
	wire w_dff_A_A3K07Dcc6_2;
	wire w_dff_A_JmiBRX3w8_2;
	wire w_dff_A_4UcCWp4o5_0;
	wire w_dff_A_KdbihPk27_0;
	wire w_dff_A_LqgYjfVH8_0;
	wire w_dff_A_9tX7QRMf3_0;
	wire w_dff_A_ChUb69I77_0;
	wire w_dff_A_ludhWNJg3_0;
	wire w_dff_A_xtPru4fd9_0;
	wire w_dff_A_ywt0VBYD4_0;
	wire w_dff_A_Huq76DsN7_0;
	wire w_dff_A_vvTiUY1m5_0;
	wire w_dff_A_ZOX8m0mE2_0;
	wire w_dff_A_vMztpKWN1_0;
	wire w_dff_A_OKKURVhr0_0;
	wire w_dff_A_LPh7b7Kr5_0;
	wire w_dff_A_VEUEFbh67_1;
	wire w_dff_A_e87aQQn08_2;
	wire w_dff_A_YvlyyIbO2_2;
	wire w_dff_A_6o6zkLh70_2;
	wire w_dff_A_bfz3X9zz6_2;
	wire w_dff_A_B7DRBSMe4_1;
	wire w_dff_A_d7G0uZeB0_1;
	wire w_dff_A_B75geTHS5_1;
	wire w_dff_A_97fE0sGQ5_1;
	wire w_dff_A_YTabs3iB8_1;
	wire w_dff_A_mmvX0yiL9_1;
	wire w_dff_A_Jqsgc3Ot4_1;
	wire w_dff_A_eUpDNywa0_2;
	wire w_dff_A_WqVsXXA43_2;
	jnot g0000(.din(w_G77_4[2]),.dout(n73),.clk(gclk));
	jcb g0001(.dina(w_G68_5[2]),.dinb(w_G58_6[2]),.dout(n74));
	jcb g0002(.dina(w_n74_0[1]),.dinb(w_G50_6[2]),.dout(n75));
	jnot g0003(.din(w_n75_0[1]),.dout(n76),.clk(gclk));
	jand g0004(.dina(n76),.dinb(w_n73_1[1]),.dout(G353),.clk(gclk));
	jnot g0005(.din(w_G87_4[1]),.dout(n78),.clk(gclk));
	jnot g0006(.din(w_G97_5[1]),.dout(n79),.clk(gclk));
	jnot g0007(.din(w_G107_3[2]),.dout(n80),.clk(gclk));
	jand g0008(.dina(w_n80_2[2]),.dinb(w_n79_1[1]),.dout(n81),.clk(gclk));
	jcb g0009(.dina(n81),.dinb(w_n78_1[1]),.dout(G355_fa_));
	jnot g0010(.din(w_G250_1[2]),.dout(n83),.clk(gclk));
	jnot g0011(.din(w_G257_1[1]),.dout(n84),.clk(gclk));
	jnot g0012(.din(w_G264_0[1]),.dout(n85),.clk(gclk));
	jand g0013(.dina(w_n85_1[1]),.dinb(w_n84_1[1]),.dout(n86),.clk(gclk));
	jcb g0014(.dina(n86),.dinb(w_n83_0[2]),.dout(n87));
	jnot g0015(.din(w_G13_2[1]),.dout(n88),.clk(gclk));
	jand g0016(.dina(w_n88_0[1]),.dinb(w_G1_2[1]),.dout(n89),.clk(gclk));
	jand g0017(.dina(w_n89_0[2]),.dinb(w_G20_7[1]),.dout(n90),.clk(gclk));
	jand g0018(.dina(w_n90_1[2]),.dinb(w_dff_B_S49LDRpI9_1),.dout(n91),.clk(gclk));
	jand g0019(.dina(w_n74_0[0]),.dinb(w_G50_6[1]),.dout(n92),.clk(gclk));
	jnot g0020(.din(w_n92_0[2]),.dout(n93),.clk(gclk));
	jand g0021(.dina(w_G20_7[0]),.dinb(w_G1_2[0]),.dout(n94),.clk(gclk));
	jand g0022(.dina(w_n94_0[2]),.dinb(w_G13_2[0]),.dout(n95),.clk(gclk));
	jand g0023(.dina(w_n95_0[1]),.dinb(n93),.dout(n96),.clk(gclk));
	jcb g0024(.dina(w_dff_B_waQ3RwkB3_0),.dinb(n91),.dout(n97));
	jcb g0025(.dina(w_n83_0[1]),.dinb(w_n78_1[0]),.dout(n98));
	jnot g0026(.din(w_G50_6[0]),.dout(n99),.clk(gclk));
	jnot g0027(.din(w_G226_1[2]),.dout(n100),.clk(gclk));
	jcb g0028(.dina(n100),.dinb(w_n99_1[2]),.dout(n101));
	jand g0029(.dina(n101),.dinb(n98),.dout(n102),.clk(gclk));
	jnot g0030(.din(w_G68_5[1]),.dout(n103),.clk(gclk));
	jnot g0031(.din(w_G238_1[1]),.dout(n104),.clk(gclk));
	jcb g0032(.dina(w_n104_0[1]),.dinb(w_n103_1[2]),.dout(n105));
	jand g0033(.dina(w_dff_B_bj3H9JTn3_0),.dinb(n102),.dout(n106),.clk(gclk));
	jnot g0034(.din(w_n94_0[1]),.dout(n107),.clk(gclk));
	jnot g0035(.din(w_G58_6[1]),.dout(n108),.clk(gclk));
	jnot g0036(.din(w_G232_1[1]),.dout(n109),.clk(gclk));
	jcb g0037(.dina(w_n109_0[1]),.dinb(w_n108_1[1]),.dout(n110));
	jand g0038(.dina(w_dff_B_dPcDd7Q30_0),.dinb(w_n107_0[2]),.dout(n111),.clk(gclk));
	jnot g0039(.din(w_G116_5[1]),.dout(n112),.clk(gclk));
	jnot g0040(.din(w_G270_0[1]),.dout(n113),.clk(gclk));
	jcb g0041(.dina(w_n113_0[1]),.dinb(w_n112_1[2]),.dout(n114));
	jcb g0042(.dina(w_n85_1[0]),.dinb(w_n80_2[1]),.dout(n115));
	jand g0043(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jcb g0044(.dina(w_n84_1[0]),.dinb(w_n79_1[0]),.dout(n117));
	jnot g0045(.din(w_G244_1[1]),.dout(n118),.clk(gclk));
	jcb g0046(.dina(w_n118_0[1]),.dinb(w_n73_1[0]),.dout(n119));
	jand g0047(.dina(n119),.dinb(n117),.dout(n120),.clk(gclk));
	jand g0048(.dina(n120),.dinb(n116),.dout(n121),.clk(gclk));
	jand g0049(.dina(n121),.dinb(n111),.dout(n122),.clk(gclk));
	jand g0050(.dina(n122),.dinb(w_dff_B_jGjlJCd88_1),.dout(n123),.clk(gclk));
	jcb g0051(.dina(n123),.dinb(w_dff_B_r3kRAIpQ2_1),.dout(G361));
	jxor g0052(.dina(w_G270_0[0]),.dinb(w_n85_0[2]),.dout(n125),.clk(gclk));
	jxor g0053(.dina(w_G257_1[0]),.dinb(w_G250_1[1]),.dout(n126),.clk(gclk));
	jxor g0054(.dina(w_dff_B_HMDYWvaT5_0),.dinb(n125),.dout(n127),.clk(gclk));
	jnot g0055(.din(w_n127_0[1]),.dout(n128),.clk(gclk));
	jxor g0056(.dina(w_G244_1[0]),.dinb(w_n104_0[0]),.dout(n129),.clk(gclk));
	jxor g0057(.dina(w_G232_1[0]),.dinb(w_G226_1[1]),.dout(n130),.clk(gclk));
	jxor g0058(.dina(w_dff_B_Cvdy09qm7_0),.dinb(n129),.dout(n131),.clk(gclk));
	jxor g0059(.dina(w_n131_0[1]),.dinb(n128),.dout(G358),.clk(gclk));
	jxor g0060(.dina(w_G58_6[0]),.dinb(w_G50_5[2]),.dout(n133),.clk(gclk));
	jxor g0061(.dina(w_G77_4[1]),.dinb(w_G68_5[0]),.dout(n134),.clk(gclk));
	jxor g0062(.dina(n134),.dinb(n133),.dout(n135),.clk(gclk));
	jxor g0063(.dina(w_G116_5[0]),.dinb(w_n80_2[0]),.dout(n136),.clk(gclk));
	jxor g0064(.dina(w_G97_5[0]),.dinb(w_G87_4[0]),.dout(n137),.clk(gclk));
	jxor g0065(.dina(w_dff_B_56hO7Xjw7_0),.dinb(n136),.dout(n138),.clk(gclk));
	jxor g0066(.dina(w_n138_0[1]),.dinb(w_n135_0[1]),.dout(G351),.clk(gclk));
	jand g0067(.dina(w_G13_1[2]),.dinb(w_G1_1[2]),.dout(n140),.clk(gclk));
	jand g0068(.dina(w_n94_0[0]),.dinb(w_G33_11[1]),.dout(n141),.clk(gclk));
	jcb g0069(.dina(w_n141_0[1]),.dinb(w_n140_1[2]),.dout(n142));
	jnot g0070(.din(w_G1_1[1]),.dout(n143),.clk(gclk));
	jand g0071(.dina(w_G13_1[1]),.dinb(w_n143_2[1]),.dout(n144),.clk(gclk));
	jand g0072(.dina(w_n144_0[1]),.dinb(w_G20_6[2]),.dout(n145),.clk(gclk));
	jcb g0073(.dina(w_n145_2[1]),.dinb(w_n142_4[1]),.dout(n146));
	jand g0074(.dina(w_G33_11[0]),.dinb(w_n143_2[0]),.dout(n147),.clk(gclk));
	jcb g0075(.dina(w_dff_B_jviK8z9P0_0),.dinb(n146),.dout(n148));
	jcb g0076(.dina(w_n148_0[2]),.dinb(w_n112_1[1]),.dout(n149));
	jand g0077(.dina(w_G116_4[2]),.dinb(w_G20_6[1]),.dout(n150),.clk(gclk));
	jnot g0078(.din(w_G20_6[0]),.dout(n151),.clk(gclk));
	jand g0079(.dina(w_G283_3[2]),.dinb(w_G33_10[2]),.dout(n152),.clk(gclk));
	jnot g0080(.din(w_G33_10[1]),.dout(n153),.clk(gclk));
	jand g0081(.dina(w_G97_4[2]),.dinb(w_n153_8[2]),.dout(n154),.clk(gclk));
	jcb g0082(.dina(n154),.dinb(w_n152_0[1]),.dout(n155));
	jand g0083(.dina(n155),.dinb(w_n151_4[1]),.dout(n156),.clk(gclk));
	jcb g0084(.dina(n156),.dinb(w_dff_B_saO59Fmz8_1),.dout(n157));
	jand g0085(.dina(n157),.dinb(w_n142_4[0]),.dout(n158),.clk(gclk));
	jand g0086(.dina(w_n145_2[0]),.dinb(w_n112_1[0]),.dout(n159),.clk(gclk));
	jcb g0087(.dina(n159),.dinb(n158),.dout(n160));
	jnot g0088(.din(n160),.dout(n161),.clk(gclk));
	jand g0089(.dina(n161),.dinb(w_dff_B_wuSjxGMb3_1),.dout(n162),.clk(gclk));
	jnot g0090(.din(w_G169_2[1]),.dout(n163),.clk(gclk));
	jnot g0091(.din(w_G274_0[2]),.dout(n164),.clk(gclk));
	jand g0092(.dina(w_G41_0[2]),.dinb(w_G33_10[0]),.dout(n165),.clk(gclk));
	jnot g0093(.din(w_n165_0[1]),.dout(n166),.clk(gclk));
	jand g0094(.dina(n166),.dinb(w_n140_1[1]),.dout(n167),.clk(gclk));
	jcb g0095(.dina(w_n167_4[1]),.dinb(w_dff_B_JapuFSpL8_1),.dout(n168));
	jnot g0096(.din(w_G41_0[1]),.dout(n169),.clk(gclk));
	jand g0097(.dina(w_G45_1[1]),.dinb(w_n143_1[2]),.dout(n170),.clk(gclk));
	jand g0098(.dina(w_n170_0[2]),.dinb(w_n169_1[1]),.dout(n171),.clk(gclk));
	jnot g0099(.din(w_n171_1[1]),.dout(n172),.clk(gclk));
	jcb g0100(.dina(w_n172_0[1]),.dinb(w_n168_0[1]),.dout(n173));
	jnot g0101(.din(w_n140_1[0]),.dout(n174),.clk(gclk));
	jcb g0102(.dina(w_n165_0[0]),.dinb(n174),.dout(n175));
	jand g0103(.dina(w_G1698_0[2]),.dinb(w_n153_8[1]),.dout(n176),.clk(gclk));
	jand g0104(.dina(w_n176_3[1]),.dinb(w_G264_0[0]),.dout(n177),.clk(gclk));
	jnot g0105(.din(w_n177_0[1]),.dout(n178),.clk(gclk));
	jand g0106(.dina(w_G303_2[2]),.dinb(w_G33_9[2]),.dout(n179),.clk(gclk));
	jnot g0107(.din(n179),.dout(n180),.clk(gclk));
	jcb g0108(.dina(w_G1698_0[1]),.dinb(w_G33_9[1]),.dout(n181));
	jcb g0109(.dina(w_n181_1[1]),.dinb(w_n84_0[2]),.dout(n182));
	jand g0110(.dina(w_dff_B_h7yKL39l2_0),.dinb(n180),.dout(n183),.clk(gclk));
	jand g0111(.dina(w_n183_0[1]),.dinb(n178),.dout(n184),.clk(gclk));
	jcb g0112(.dina(n184),.dinb(w_n175_3[1]),.dout(n185));
	jcb g0113(.dina(w_n171_1[0]),.dinb(w_n113_0[0]),.dout(n186));
	jcb g0114(.dina(n186),.dinb(w_n167_4[0]),.dout(n187));
	jand g0115(.dina(w_n187_0[1]),.dinb(n185),.dout(n188),.clk(gclk));
	jand g0116(.dina(n188),.dinb(w_n173_0[2]),.dout(n189),.clk(gclk));
	jcb g0117(.dina(w_n189_0[1]),.dinb(w_n163_1[1]),.dout(n190));
	jnot g0118(.din(w_G179_1[1]),.dout(n191),.clk(gclk));
	jand g0119(.dina(w_n175_3[0]),.dinb(w_G274_0[1]),.dout(n192),.clk(gclk));
	jand g0120(.dina(w_n171_0[2]),.dinb(n192),.dout(n193),.clk(gclk));
	jnot g0121(.din(w_n183_0[0]),.dout(n194),.clk(gclk));
	jcb g0122(.dina(n194),.dinb(w_n177_0[0]),.dout(n195));
	jand g0123(.dina(n195),.dinb(w_n167_3[2]),.dout(n196),.clk(gclk));
	jnot g0124(.din(w_n187_0[0]),.dout(n197),.clk(gclk));
	jcb g0125(.dina(w_dff_B_gF9WsJ4t1_0),.dinb(n196),.dout(n198));
	jcb g0126(.dina(n198),.dinb(w_n193_0[2]),.dout(n199));
	jcb g0127(.dina(w_n199_0[2]),.dinb(w_n191_3[2]),.dout(n200));
	jand g0128(.dina(w_n200_0[1]),.dinb(n190),.dout(n201),.clk(gclk));
	jcb g0129(.dina(n201),.dinb(w_n162_0[1]),.dout(n202));
	jand g0130(.dina(w_n199_0[1]),.dinb(w_G200_2[1]),.dout(n203),.clk(gclk));
	jnot g0131(.din(w_n162_0[0]),.dout(n204),.clk(gclk));
	jand g0132(.dina(w_n189_0[0]),.dinb(w_G190_4[2]),.dout(n205),.clk(gclk));
	jcb g0133(.dina(n205),.dinb(w_n204_0[1]),.dout(n206));
	jcb g0134(.dina(n206),.dinb(w_dff_B_Di3rUeFI3_1),.dout(n207));
	jand g0135(.dina(n207),.dinb(w_n202_0[2]),.dout(n208),.clk(gclk));
	jcb g0136(.dina(w_n171_0[1]),.dinb(w_n85_0[1]),.dout(n209));
	jcb g0137(.dina(n209),.dinb(w_n167_3[1]),.dout(n210));
	jnot g0138(.din(w_G1698_0[0]),.dout(n211),.clk(gclk));
	jcb g0139(.dina(w_n211_0[1]),.dinb(w_G33_9[0]),.dout(n212));
	jcb g0140(.dina(n212),.dinb(w_n84_0[1]),.dout(n213));
	jand g0141(.dina(w_G294_3[1]),.dinb(w_G33_8[2]),.dout(n214),.clk(gclk));
	jnot g0142(.din(w_n214_0[1]),.dout(n215),.clk(gclk));
	jcb g0143(.dina(w_n181_1[0]),.dinb(w_n83_0[0]),.dout(n216));
	jand g0144(.dina(w_dff_B_WafiYv6g5_0),.dinb(n215),.dout(n217),.clk(gclk));
	jand g0145(.dina(n217),.dinb(w_dff_B_oLqY92ZG7_1),.dout(n218),.clk(gclk));
	jcb g0146(.dina(n218),.dinb(w_n175_2[2]),.dout(n219));
	jand g0147(.dina(n219),.dinb(w_n173_0[1]),.dout(n220),.clk(gclk));
	jand g0148(.dina(n220),.dinb(w_n210_0[1]),.dout(n221),.clk(gclk));
	jcb g0149(.dina(w_n221_1[1]),.dinb(w_G169_2[0]),.dout(n222));
	jcb g0150(.dina(w_n148_0[1]),.dinb(w_n80_1[2]),.dout(n223));
	jnot g0151(.din(w_n223_0[1]),.dout(n224),.clk(gclk));
	jcb g0152(.dina(w_n141_0[0]),.dinb(w_G13_1[0]),.dout(n225));
	jand g0153(.dina(w_n80_1[1]),.dinb(w_G20_5[2]),.dout(n226),.clk(gclk));
	jand g0154(.dina(n226),.dinb(w_n225_0[1]),.dout(n227),.clk(gclk));
	jand g0155(.dina(w_G116_4[1]),.dinb(w_G33_8[1]),.dout(n228),.clk(gclk));
	jand g0156(.dina(w_G87_3[2]),.dinb(w_n153_8[0]),.dout(n229),.clk(gclk));
	jcb g0157(.dina(n229),.dinb(w_n228_0[1]),.dout(n230));
	jand g0158(.dina(n230),.dinb(w_n142_3[2]),.dout(n231),.clk(gclk));
	jand g0159(.dina(n231),.dinb(w_n151_4[0]),.dout(n232),.clk(gclk));
	jcb g0160(.dina(n232),.dinb(w_dff_B_K7Pdc8mo9_1),.dout(n233));
	jcb g0161(.dina(w_n233_0[1]),.dinb(n224),.dout(n234));
	jnot g0162(.din(w_n210_0[0]),.dout(n235),.clk(gclk));
	jand g0163(.dina(w_n176_3[0]),.dinb(w_G257_0[2]),.dout(n236),.clk(gclk));
	jand g0164(.dina(w_n211_0[0]),.dinb(w_n153_7[2]),.dout(n237),.clk(gclk));
	jand g0165(.dina(w_n237_1[2]),.dinb(w_G250_1[0]),.dout(n238),.clk(gclk));
	jcb g0166(.dina(n238),.dinb(w_n214_0[0]),.dout(n239));
	jcb g0167(.dina(n239),.dinb(n236),.dout(n240));
	jand g0168(.dina(n240),.dinb(w_n167_3[0]),.dout(n241),.clk(gclk));
	jcb g0169(.dina(n241),.dinb(w_n193_0[1]),.dout(n242));
	jcb g0170(.dina(n242),.dinb(n235),.dout(n243));
	jcb g0171(.dina(w_n243_0[1]),.dinb(w_G179_1[0]),.dout(n244));
	jand g0172(.dina(n244),.dinb(w_n234_0[1]),.dout(n245),.clk(gclk));
	jand g0173(.dina(w_dff_B_QtalDuBA3_0),.dinb(n222),.dout(n246),.clk(gclk));
	jand g0174(.dina(w_n221_1[0]),.dinb(w_G190_4[1]),.dout(n247),.clk(gclk));
	jnot g0175(.din(n247),.dout(n248),.clk(gclk));
	jnot g0176(.din(w_n233_0[0]),.dout(n249),.clk(gclk));
	jand g0177(.dina(n249),.dinb(w_n223_0[0]),.dout(n250),.clk(gclk));
	jnot g0178(.din(w_G200_2[0]),.dout(n251),.clk(gclk));
	jcb g0179(.dina(w_n221_0[2]),.dinb(w_n251_2[2]),.dout(n252));
	jand g0180(.dina(n252),.dinb(n250),.dout(n253),.clk(gclk));
	jand g0181(.dina(w_dff_B_OlWs8Heb2_0),.dinb(n248),.dout(n254),.clk(gclk));
	jcb g0182(.dina(n254),.dinb(w_n246_0[2]),.dout(n255));
	jnot g0183(.din(w_n255_1[1]),.dout(n256),.clk(gclk));
	jand g0184(.dina(w_n176_2[2]),.dinb(w_G244_0[2]),.dout(n257),.clk(gclk));
	jand g0185(.dina(w_n237_1[1]),.dinb(w_G238_1[0]),.dout(n258),.clk(gclk));
	jcb g0186(.dina(n258),.dinb(w_n228_0[0]),.dout(n259));
	jcb g0187(.dina(n259),.dinb(n257),.dout(n260));
	jcb g0188(.dina(n260),.dinb(w_n175_2[1]),.dout(n261));
	jnot g0189(.din(w_n170_0[1]),.dout(n262),.clk(gclk));
	jand g0190(.dina(n262),.dinb(w_G250_0[2]),.dout(n263),.clk(gclk));
	jand g0191(.dina(w_n170_0[0]),.dinb(w_G274_0[0]),.dout(n264),.clk(gclk));
	jcb g0192(.dina(w_dff_B_nOF57Ihc9_0),.dinb(n263),.dout(n265));
	jcb g0193(.dina(n265),.dinb(w_n167_2[2]),.dout(n266));
	jand g0194(.dina(n266),.dinb(w_dff_B_vu9Wbdxq9_1),.dout(n267),.clk(gclk));
	jand g0195(.dina(w_n267_1[2]),.dinb(w_G200_1[2]),.dout(n268),.clk(gclk));
	jnot g0196(.din(w_n148_0[0]),.dout(n269),.clk(gclk));
	jand g0197(.dina(w_n269_0[1]),.dinb(w_G87_3[1]),.dout(n270),.clk(gclk));
	jand g0198(.dina(w_n79_0[2]),.dinb(w_n78_0[2]),.dout(n271),.clk(gclk));
	jand g0199(.dina(n271),.dinb(w_n80_1[0]),.dout(n272),.clk(gclk));
	jand g0200(.dina(w_n272_0[1]),.dinb(w_G20_5[1]),.dout(n273),.clk(gclk));
	jnot g0201(.din(n273),.dout(n274),.clk(gclk));
	jand g0202(.dina(w_G97_4[1]),.dinb(w_G33_8[0]),.dout(n275),.clk(gclk));
	jand g0203(.dina(w_G68_4[2]),.dinb(w_n153_7[1]),.dout(n276),.clk(gclk));
	jcb g0204(.dina(n276),.dinb(w_G20_5[0]),.dout(n277));
	jcb g0205(.dina(n277),.dinb(w_n275_0[1]),.dout(n278));
	jand g0206(.dina(n278),.dinb(w_n142_3[1]),.dout(n279),.clk(gclk));
	jand g0207(.dina(w_dff_B_52PmUoso1_0),.dinb(n274),.dout(n280),.clk(gclk));
	jand g0208(.dina(w_n145_1[2]),.dinb(w_n78_0[1]),.dout(n281),.clk(gclk));
	jcb g0209(.dina(w_dff_B_yxtZg7tQ0_0),.dinb(n280),.dout(n282));
	jcb g0210(.dina(n282),.dinb(w_dff_B_NMpI85nN2_1),.dout(n283));
	jnot g0211(.din(w_G190_4[0]),.dout(n284),.clk(gclk));
	jcb g0212(.dina(w_n267_1[1]),.dinb(w_n284_1[2]),.dout(n285));
	jnot g0213(.din(w_n285_0[1]),.dout(n286),.clk(gclk));
	jcb g0214(.dina(n286),.dinb(w_n283_1[1]),.dout(n287));
	jcb g0215(.dina(n287),.dinb(w_n268_0[1]),.dout(n288));
	jnot g0216(.din(w_n267_1[0]),.dout(n289),.clk(gclk));
	jand g0217(.dina(w_n289_0[1]),.dinb(w_n191_3[1]),.dout(n290),.clk(gclk));
	jnot g0218(.din(w_n283_1[0]),.dout(n291),.clk(gclk));
	jand g0219(.dina(w_n267_0[2]),.dinb(w_n163_1[0]),.dout(n292),.clk(gclk));
	jcb g0220(.dina(w_n292_0[1]),.dinb(w_n291_0[1]),.dout(n293));
	jcb g0221(.dina(n293),.dinb(w_n290_0[1]),.dout(n294));
	jand g0222(.dina(w_n294_0[1]),.dinb(w_dff_B_2sX8viCE6_1),.dout(n295),.clk(gclk));
	jand g0223(.dina(w_n172_0[0]),.dinb(w_G257_0[1]),.dout(n296),.clk(gclk));
	jand g0224(.dina(n296),.dinb(w_n175_2[0]),.dout(n297),.clk(gclk));
	jand g0225(.dina(w_n176_2[1]),.dinb(w_G250_0[1]),.dout(n298),.clk(gclk));
	jnot g0226(.din(w_n152_0[0]),.dout(n299),.clk(gclk));
	jcb g0227(.dina(w_n181_0[2]),.dinb(w_n118_0[0]),.dout(n300));
	jand g0228(.dina(w_dff_B_Su4cP8Us5_0),.dinb(n299),.dout(n301),.clk(gclk));
	jnot g0229(.din(w_n301_0[1]),.dout(n302),.clk(gclk));
	jcb g0230(.dina(n302),.dinb(w_n298_0[1]),.dout(n303));
	jand g0231(.dina(n303),.dinb(w_n167_2[1]),.dout(n304),.clk(gclk));
	jcb g0232(.dina(n304),.dinb(w_n193_0[0]),.dout(n305));
	jcb g0233(.dina(w_dff_B_BZ4DsGxm4_0),.dinb(w_n297_0[1]),.dout(n306));
	jand g0234(.dina(w_n306_1[1]),.dinb(w_n163_0[2]),.dout(n307),.clk(gclk));
	jand g0235(.dina(w_n269_0[0]),.dinb(w_G97_4[0]),.dout(n308),.clk(gclk));
	jxor g0236(.dina(w_G107_3[1]),.dinb(w_G97_3[2]),.dout(n309),.clk(gclk));
	jand g0237(.dina(w_n309_0[1]),.dinb(w_G20_4[2]),.dout(n310),.clk(gclk));
	jnot g0238(.din(n310),.dout(n311),.clk(gclk));
	jand g0239(.dina(w_G107_3[0]),.dinb(w_G33_7[2]),.dout(n312),.clk(gclk));
	jand g0240(.dina(w_G77_4[0]),.dinb(w_n153_7[0]),.dout(n313),.clk(gclk));
	jcb g0241(.dina(n313),.dinb(w_G20_4[1]),.dout(n314));
	jcb g0242(.dina(n314),.dinb(w_n312_0[1]),.dout(n315));
	jand g0243(.dina(n315),.dinb(w_n142_3[0]),.dout(n316),.clk(gclk));
	jand g0244(.dina(n316),.dinb(n311),.dout(n317),.clk(gclk));
	jand g0245(.dina(w_n145_1[1]),.dinb(w_n79_0[1]),.dout(n318),.clk(gclk));
	jcb g0246(.dina(n318),.dinb(n317),.dout(n319));
	jcb g0247(.dina(w_dff_B_6hZTUKfw7_0),.dinb(n308),.dout(n320));
	jnot g0248(.din(w_n320_1[1]),.dout(n321),.clk(gclk));
	jnot g0249(.din(w_n297_0[0]),.dout(n322),.clk(gclk));
	jnot g0250(.din(w_n298_0[0]),.dout(n323),.clk(gclk));
	jand g0251(.dina(w_n301_0[0]),.dinb(n323),.dout(n324),.clk(gclk));
	jcb g0252(.dina(n324),.dinb(w_n175_1[2]),.dout(n325));
	jand g0253(.dina(n325),.dinb(w_n173_0[0]),.dout(n326),.clk(gclk));
	jand g0254(.dina(w_dff_B_xlKVheb49_0),.dinb(n322),.dout(n327),.clk(gclk));
	jand g0255(.dina(w_n327_1[1]),.dinb(w_n191_3[0]),.dout(n328),.clk(gclk));
	jcb g0256(.dina(n328),.dinb(w_n321_0[1]),.dout(n329));
	jcb g0257(.dina(n329),.dinb(w_n307_0[1]),.dout(n330));
	jand g0258(.dina(w_n327_1[0]),.dinb(w_G190_3[2]),.dout(n331),.clk(gclk));
	jand g0259(.dina(w_n306_1[0]),.dinb(w_G200_1[1]),.dout(n332),.clk(gclk));
	jcb g0260(.dina(n332),.dinb(w_n320_1[0]),.dout(n333));
	jcb g0261(.dina(w_dff_B_92Xyjyt49_0),.dinb(w_n331_0[1]),.dout(n334));
	jand g0262(.dina(w_n334_0[1]),.dinb(w_n330_0[1]),.dout(n335),.clk(gclk));
	jand g0263(.dina(w_n335_0[1]),.dinb(w_n295_0[1]),.dout(n336),.clk(gclk));
	jand g0264(.dina(n336),.dinb(w_dff_B_m2KEuw7G7_1),.dout(n337),.clk(gclk));
	jand g0265(.dina(n337),.dinb(w_n208_0[1]),.dout(n338),.clk(gclk));
	jnot g0266(.din(w_G45_1[0]),.dout(n339),.clk(gclk));
	jand g0267(.dina(w_n339_1[1]),.dinb(w_n169_1[0]),.dout(n340),.clk(gclk));
	jcb g0268(.dina(n340),.dinb(w_G1_1[0]),.dout(n341));
	jcb g0269(.dina(w_n341_0[1]),.dinb(w_n168_0[0]),.dout(n342));
	jand g0270(.dina(w_n176_2[0]),.dinb(w_G238_0[2]),.dout(n343),.clk(gclk));
	jnot g0271(.din(n343),.dout(n344),.clk(gclk));
	jnot g0272(.din(w_n312_0[0]),.dout(n345),.clk(gclk));
	jcb g0273(.dina(w_n181_0[1]),.dinb(w_n109_0[0]),.dout(n346));
	jand g0274(.dina(w_dff_B_cjLmZ3eg8_0),.dinb(n345),.dout(n347),.clk(gclk));
	jand g0275(.dina(w_dff_B_fPnJjukF7_0),.dinb(n344),.dout(n348),.clk(gclk));
	jcb g0276(.dina(n348),.dinb(w_n175_1[1]),.dout(n349));
	jand g0277(.dina(w_n341_0[0]),.dinb(w_n175_1[0]),.dout(n350),.clk(gclk));
	jand g0278(.dina(w_n350_1[1]),.dinb(w_G244_0[1]),.dout(n351),.clk(gclk));
	jnot g0279(.din(n351),.dout(n352),.clk(gclk));
	jand g0280(.dina(n352),.dinb(n349),.dout(n353),.clk(gclk));
	jand g0281(.dina(n353),.dinb(w_n342_0[1]),.dout(n354),.clk(gclk));
	jnot g0282(.din(w_n354_1[1]),.dout(n355),.clk(gclk));
	jand g0283(.dina(n355),.dinb(w_n163_0[1]),.dout(n356),.clk(gclk));
	jand g0284(.dina(w_G87_3[0]),.dinb(w_G33_7[1]),.dout(n357),.clk(gclk));
	jand g0285(.dina(w_G58_5[2]),.dinb(w_n153_6[2]),.dout(n358),.clk(gclk));
	jcb g0286(.dina(n358),.dinb(w_n357_0[1]),.dout(n359));
	jand g0287(.dina(n359),.dinb(w_n151_3[2]),.dout(n360),.clk(gclk));
	jand g0288(.dina(n360),.dinb(w_n142_2[2]),.dout(n361),.clk(gclk));
	jand g0289(.dina(w_n140_0[2]),.dinb(w_n151_3[1]),.dout(n362),.clk(gclk));
	jnot g0290(.din(w_n362_0[1]),.dout(n363),.clk(gclk));
	jand g0291(.dina(w_G20_4[0]),.dinb(w_n143_1[1]),.dout(n364),.clk(gclk));
	jnot g0292(.din(w_n364_0[1]),.dout(n365),.clk(gclk));
	jand g0293(.dina(n365),.dinb(w_G77_3[2]),.dout(n366),.clk(gclk));
	jand g0294(.dina(n366),.dinb(w_dff_B_Yxob6LeF8_1),.dout(n367),.clk(gclk));
	jand g0295(.dina(w_n145_1[0]),.dinb(w_n73_0[2]),.dout(n368),.clk(gclk));
	jcb g0296(.dina(w_dff_B_DXhI0XcQ3_0),.dinb(n367),.dout(n369));
	jcb g0297(.dina(n369),.dinb(w_dff_B_CwEn7Y6z2_1),.dout(n370));
	jnot g0298(.din(w_n370_0[1]),.dout(n371),.clk(gclk));
	jand g0299(.dina(w_n354_1[0]),.dinb(w_n191_2[2]),.dout(n372),.clk(gclk));
	jcb g0300(.dina(n372),.dinb(w_n371_0[1]),.dout(n373));
	jcb g0301(.dina(w_dff_B_afLhG7oH1_0),.dinb(n356),.dout(n374));
	jnot g0302(.din(w_n374_0[1]),.dout(n375),.clk(gclk));
	jand g0303(.dina(w_n354_0[2]),.dinb(w_G190_3[1]),.dout(n376),.clk(gclk));
	jnot g0304(.din(n376),.dout(n377),.clk(gclk));
	jcb g0305(.dina(w_n354_0[1]),.dinb(w_n251_2[1]),.dout(n378));
	jand g0306(.dina(n378),.dinb(w_n371_0[0]),.dout(n379),.clk(gclk));
	jand g0307(.dina(w_dff_B_2lravuW69_0),.dinb(n377),.dout(n380),.clk(gclk));
	jcb g0308(.dina(n380),.dinb(w_n375_0[1]),.dout(n381));
	jand g0309(.dina(w_n350_1[0]),.dinb(w_G238_0[1]),.dout(n382),.clk(gclk));
	jnot g0310(.din(w_n342_0[0]),.dout(n383),.clk(gclk));
	jand g0311(.dina(w_n176_1[2]),.dinb(w_G232_0[2]),.dout(n384),.clk(gclk));
	jand g0312(.dina(w_n237_1[0]),.dinb(w_G226_1[0]),.dout(n385),.clk(gclk));
	jcb g0313(.dina(n385),.dinb(w_n275_0[0]),.dout(n386));
	jcb g0314(.dina(n386),.dinb(n384),.dout(n387));
	jand g0315(.dina(n387),.dinb(w_n167_2[0]),.dout(n388),.clk(gclk));
	jcb g0316(.dina(n388),.dinb(w_n383_0[2]),.dout(n389));
	jcb g0317(.dina(n389),.dinb(n382),.dout(n390));
	jnot g0318(.din(n390),.dout(n391),.clk(gclk));
	jand g0319(.dina(w_n391_1[1]),.dinb(w_G190_3[0]),.dout(n392),.clk(gclk));
	jnot g0320(.din(n392),.dout(n393),.clk(gclk));
	jand g0321(.dina(w_G77_3[1]),.dinb(w_G33_7[0]),.dout(n394),.clk(gclk));
	jand g0322(.dina(w_G50_5[1]),.dinb(w_n153_6[1]),.dout(n395),.clk(gclk));
	jcb g0323(.dina(n395),.dinb(w_n394_0[1]),.dout(n396));
	jand g0324(.dina(n396),.dinb(w_n142_2[1]),.dout(n397),.clk(gclk));
	jand g0325(.dina(n397),.dinb(w_n151_3[0]),.dout(n398),.clk(gclk));
	jnot g0326(.din(n398),.dout(n399),.clk(gclk));
	jand g0327(.dina(w_n103_1[1]),.dinb(w_G20_3[2]),.dout(n400),.clk(gclk));
	jand g0328(.dina(n400),.dinb(w_n225_0[0]),.dout(n401),.clk(gclk));
	jnot g0329(.din(n401),.dout(n402),.clk(gclk));
	jcb g0330(.dina(w_n364_0[0]),.dinb(w_n142_2[0]),.dout(n403));
	jcb g0331(.dina(w_n403_0[2]),.dinb(w_n103_1[0]),.dout(n404));
	jand g0332(.dina(w_dff_B_msIF60Dn0_0),.dinb(n402),.dout(n405),.clk(gclk));
	jand g0333(.dina(n405),.dinb(n399),.dout(n406),.clk(gclk));
	jcb g0334(.dina(w_n391_1[0]),.dinb(w_n251_2[0]),.dout(n407));
	jand g0335(.dina(w_dff_B_vud1sdUj5_0),.dinb(w_n406_0[2]),.dout(n408),.clk(gclk));
	jand g0336(.dina(n408),.dinb(n393),.dout(n409),.clk(gclk));
	jcb g0337(.dina(w_n391_0[2]),.dinb(w_G169_1[2]),.dout(n410));
	jand g0338(.dina(w_n391_0[1]),.dinb(w_n191_2[1]),.dout(n411),.clk(gclk));
	jcb g0339(.dina(n411),.dinb(w_n406_0[1]),.dout(n412));
	jnot g0340(.din(n412),.dout(n413),.clk(gclk));
	jand g0341(.dina(n413),.dinb(w_dff_B_z3fMj7fk0_1),.dout(n414),.clk(gclk));
	jcb g0342(.dina(w_n414_0[1]),.dinb(w_n409_0[1]),.dout(n415));
	jand g0343(.dina(w_n350_0[2]),.dinb(w_G226_0[2]),.dout(n416),.clk(gclk));
	jand g0344(.dina(w_n176_1[1]),.dinb(w_G223_0[1]),.dout(n417),.clk(gclk));
	jand g0345(.dina(w_n237_0[2]),.dinb(w_dff_B_wO9YYGgD8_1),.dout(n418),.clk(gclk));
	jcb g0346(.dina(n418),.dinb(w_n394_0[0]),.dout(n419));
	jcb g0347(.dina(n419),.dinb(n417),.dout(n420));
	jand g0348(.dina(n420),.dinb(w_n167_1[2]),.dout(n421),.clk(gclk));
	jcb g0349(.dina(n421),.dinb(w_n383_0[1]),.dout(n422));
	jcb g0350(.dina(n422),.dinb(n416),.dout(n423));
	jnot g0351(.din(n423),.dout(n424),.clk(gclk));
	jand g0352(.dina(w_n424_1[1]),.dinb(w_G190_2[2]),.dout(n425),.clk(gclk));
	jnot g0353(.din(n425),.dout(n426),.clk(gclk));
	jand g0354(.dina(w_G33_6[2]),.dinb(w_n151_2[2]),.dout(n427),.clk(gclk));
	jand g0355(.dina(w_n427_0[1]),.dinb(w_G58_5[1]),.dout(n428),.clk(gclk));
	jand g0356(.dina(w_n75_0[0]),.dinb(w_G20_3[1]),.dout(n429),.clk(gclk));
	jand g0357(.dina(w_n153_6[0]),.dinb(w_n151_2[1]),.dout(n430),.clk(gclk));
	jand g0358(.dina(w_n430_0[1]),.dinb(w_G150_3[1]),.dout(n431),.clk(gclk));
	jcb g0359(.dina(n431),.dinb(w_dff_B_dbxYtjsB5_1),.dout(n432));
	jcb g0360(.dina(n432),.dinb(n428),.dout(n433));
	jand g0361(.dina(n433),.dinb(w_n142_1[2]),.dout(n434),.clk(gclk));
	jnot g0362(.din(n434),.dout(n435),.clk(gclk));
	jnot g0363(.din(w_n145_0[2]),.dout(n436),.clk(gclk));
	jand g0364(.dina(w_n436_0[1]),.dinb(w_n99_1[1]),.dout(n437),.clk(gclk));
	jand g0365(.dina(w_n403_0[1]),.dinb(w_G50_5[0]),.dout(n438),.clk(gclk));
	jcb g0366(.dina(w_dff_B_YoXN2Ew11_0),.dinb(n437),.dout(n439));
	jand g0367(.dina(n439),.dinb(n435),.dout(n440),.clk(gclk));
	jcb g0368(.dina(w_n424_1[0]),.dinb(w_n251_1[2]),.dout(n441));
	jand g0369(.dina(w_dff_B_UU5jplzl4_0),.dinb(w_n440_0[2]),.dout(n442),.clk(gclk));
	jand g0370(.dina(n442),.dinb(n426),.dout(n443),.clk(gclk));
	jcb g0371(.dina(w_n424_0[2]),.dinb(w_G169_1[1]),.dout(n444));
	jand g0372(.dina(w_n424_0[1]),.dinb(w_n191_2[0]),.dout(n445),.clk(gclk));
	jcb g0373(.dina(n445),.dinb(w_n440_0[1]),.dout(n446));
	jnot g0374(.din(n446),.dout(n447),.clk(gclk));
	jand g0375(.dina(n447),.dinb(w_dff_B_wG9g4L8p8_1),.dout(n448),.clk(gclk));
	jcb g0376(.dina(w_n448_0[1]),.dinb(w_n443_0[1]),.dout(n449));
	jand g0377(.dina(w_n350_0[1]),.dinb(w_G232_0[1]),.dout(n450),.clk(gclk));
	jand g0378(.dina(w_n176_1[0]),.dinb(w_G226_0[1]),.dout(n451),.clk(gclk));
	jand g0379(.dina(w_n237_0[1]),.dinb(w_G223_0[0]),.dout(n452),.clk(gclk));
	jcb g0380(.dina(n452),.dinb(w_n357_0[0]),.dout(n453));
	jcb g0381(.dina(n453),.dinb(n451),.dout(n454));
	jand g0382(.dina(n454),.dinb(w_n167_1[1]),.dout(n455),.clk(gclk));
	jcb g0383(.dina(n455),.dinb(w_n383_0[0]),.dout(n456));
	jcb g0384(.dina(n456),.dinb(n450),.dout(n457));
	jnot g0385(.din(n457),.dout(n458),.clk(gclk));
	jcb g0386(.dina(w_n458_1[1]),.dinb(w_G169_1[0]),.dout(n459));
	jand g0387(.dina(w_n430_0[0]),.dinb(w_G159_3[2]),.dout(n460),.clk(gclk));
	jxor g0388(.dina(w_G68_4[1]),.dinb(w_G58_5[0]),.dout(n461),.clk(gclk));
	jcb g0389(.dina(n461),.dinb(w_n151_2[0]),.dout(n462));
	jnot g0390(.din(n462),.dout(n463),.clk(gclk));
	jand g0391(.dina(w_n427_0[0]),.dinb(w_G68_4[0]),.dout(n464),.clk(gclk));
	jcb g0392(.dina(n464),.dinb(w_dff_B_8MCw01Rg0_1),.dout(n465));
	jcb g0393(.dina(n465),.dinb(n460),.dout(n466));
	jand g0394(.dina(n466),.dinb(w_n142_1[1]),.dout(n467),.clk(gclk));
	jnot g0395(.din(n467),.dout(n468),.clk(gclk));
	jand g0396(.dina(w_n436_0[0]),.dinb(w_n108_1[0]),.dout(n469),.clk(gclk));
	jand g0397(.dina(w_n403_0[0]),.dinb(w_G58_4[2]),.dout(n470),.clk(gclk));
	jcb g0398(.dina(w_dff_B_2c7q3EWk1_0),.dinb(n469),.dout(n471));
	jand g0399(.dina(n471),.dinb(n468),.dout(n472),.clk(gclk));
	jand g0400(.dina(w_n458_1[0]),.dinb(w_n191_1[2]),.dout(n473),.clk(gclk));
	jcb g0401(.dina(n473),.dinb(w_n472_0[1]),.dout(n474));
	jnot g0402(.din(n474),.dout(n475),.clk(gclk));
	jand g0403(.dina(n475),.dinb(w_dff_B_N05izYLT1_1),.dout(n476),.clk(gclk));
	jcb g0404(.dina(w_n458_0[2]),.dinb(w_n251_1[1]),.dout(n477));
	jnot g0405(.din(w_n472_0[0]),.dout(n478),.clk(gclk));
	jand g0406(.dina(w_n458_0[1]),.dinb(w_G190_2[1]),.dout(n479),.clk(gclk));
	jcb g0407(.dina(w_dff_B_2tHWsNiR9_0),.dinb(w_n478_0[1]),.dout(n480));
	jnot g0408(.din(n480),.dout(n481),.clk(gclk));
	jand g0409(.dina(n481),.dinb(w_dff_B_H0JpnCjm0_1),.dout(n482),.clk(gclk));
	jcb g0410(.dina(n482),.dinb(w_n476_0[2]),.dout(n483));
	jcb g0411(.dina(w_n483_0[1]),.dinb(w_n449_0[1]),.dout(n484));
	jcb g0412(.dina(w_n484_0[1]),.dinb(w_n415_1[1]),.dout(n485));
	jcb g0413(.dina(w_dff_B_bXb4hhhe3_0),.dinb(w_n381_0[2]),.dout(n486));
	jnot g0414(.din(w_n486_0[1]),.dout(n487),.clk(gclk));
	jand g0415(.dina(w_n487_0[2]),.dinb(w_n338_0[1]),.dout(G372),.clk(gclk));
	jnot g0416(.din(w_n268_0[0]),.dout(n489),.clk(gclk));
	jand g0417(.dina(w_n285_0[0]),.dinb(w_n291_0[0]),.dout(n490),.clk(gclk));
	jand g0418(.dina(n490),.dinb(w_dff_B_qdGSDyRC3_1),.dout(n491),.clk(gclk));
	jcb g0419(.dina(w_n330_0[0]),.dinb(w_n491_0[1]),.dout(n492));
	jnot g0420(.din(w_n290_0[0]),.dout(n493),.clk(gclk));
	jnot g0421(.din(w_n292_0[0]),.dout(n494),.clk(gclk));
	jand g0422(.dina(n494),.dinb(w_n283_0[2]),.dout(n495),.clk(gclk));
	jand g0423(.dina(n495),.dinb(n493),.dout(n496),.clk(gclk));
	jcb g0424(.dina(n496),.dinb(w_n491_0[0]),.dout(n497));
	jnot g0425(.din(w_n307_0[0]),.dout(n498),.clk(gclk));
	jcb g0426(.dina(w_n306_0[2]),.dinb(w_G179_0[2]),.dout(n499));
	jand g0427(.dina(n499),.dinb(w_n320_0[2]),.dout(n500),.clk(gclk));
	jand g0428(.dina(w_dff_B_MNhyYSQm0_0),.dinb(n498),.dout(n501),.clk(gclk));
	jnot g0429(.din(w_n331_0[0]),.dout(n502),.clk(gclk));
	jcb g0430(.dina(w_n327_0[2]),.dinb(w_n251_1[0]),.dout(n503));
	jand g0431(.dina(n503),.dinb(w_n321_0[0]),.dout(n504),.clk(gclk));
	jand g0432(.dina(w_dff_B_VxFm5xip0_0),.dinb(n502),.dout(n505),.clk(gclk));
	jcb g0433(.dina(n505),.dinb(w_n501_0[1]),.dout(n506));
	jcb g0434(.dina(w_n506_0[1]),.dinb(w_n497_0[1]),.dout(n507));
	jnot g0435(.din(w_n246_0[1]),.dout(n508),.clk(gclk));
	jcb g0436(.dina(w_n255_1[0]),.dinb(w_n202_0[1]),.dout(n509));
	jand g0437(.dina(n509),.dinb(w_dff_B_yOM4cw0L7_1),.dout(n510),.clk(gclk));
	jcb g0438(.dina(w_n510_0[1]),.dinb(n507),.dout(n511));
	jand g0439(.dina(n511),.dinb(w_n294_0[0]),.dout(n512),.clk(gclk));
	jand g0440(.dina(n512),.dinb(w_dff_B_PXQbvnM88_1),.dout(n513),.clk(gclk));
	jcb g0441(.dina(w_n513_0[1]),.dinb(w_n486_0[0]),.dout(n514));
	jnot g0442(.din(w_n514_0[1]),.dout(n515),.clk(gclk));
	jnot g0443(.din(w_n443_0[0]),.dout(n516),.clk(gclk));
	jand g0444(.dina(w_n476_0[1]),.dinb(n516),.dout(n517),.clk(gclk));
	jnot g0445(.din(n517),.dout(n518),.clk(gclk));
	jnot g0446(.din(w_n448_0[0]),.dout(n519),.clk(gclk));
	jnot g0447(.din(w_n414_0[0]),.dout(n520),.clk(gclk));
	jcb g0448(.dina(w_n415_1[0]),.dinb(w_n374_0[0]),.dout(n521));
	jand g0449(.dina(n521),.dinb(w_n520_0[1]),.dout(n522),.clk(gclk));
	jcb g0450(.dina(n522),.dinb(w_n484_0[0]),.dout(n523));
	jand g0451(.dina(n523),.dinb(w_dff_B_OJKARMjA2_1),.dout(n524),.clk(gclk));
	jand g0452(.dina(n524),.dinb(n518),.dout(n525),.clk(gclk));
	jnot g0453(.din(w_n525_0[1]),.dout(n526),.clk(gclk));
	jcb g0454(.dina(w_dff_B_6QtizgNK7_0),.dinb(n515),.dout(G369));
	jnot g0455(.din(w_n208_0[0]),.dout(n528),.clk(gclk));
	jand g0456(.dina(w_G213_0[1]),.dinb(w_n151_1[2]),.dout(n529),.clk(gclk));
	jand g0457(.dina(n529),.dinb(w_n144_0[0]),.dout(n530),.clk(gclk));
	jand g0458(.dina(w_n530_1[1]),.dinb(w_G343_0[1]),.dout(n531),.clk(gclk));
	jand g0459(.dina(w_n531_4[2]),.dinb(w_n204_0[0]),.dout(n532),.clk(gclk));
	jxor g0460(.dina(w_dff_B_qv6ztYWL1_0),.dinb(n528),.dout(n533),.clk(gclk));
	jnot g0461(.din(w_n533_0[1]),.dout(n534),.clk(gclk));
	jand g0462(.dina(w_n534_0[1]),.dinb(w_G330_0[2]),.dout(n535),.clk(gclk));
	jand g0463(.dina(w_n531_4[1]),.dinb(w_n234_0[0]),.dout(n536),.clk(gclk));
	jxor g0464(.dina(w_dff_B_MMoY9aKr6_0),.dinb(w_n255_0[2]),.dout(n537),.clk(gclk));
	jnot g0465(.din(w_n537_0[1]),.dout(n538),.clk(gclk));
	jand g0466(.dina(w_n538_0[2]),.dinb(w_n535_0[1]),.dout(n539),.clk(gclk));
	jnot g0467(.din(w_n510_0[0]),.dout(n540),.clk(gclk));
	jnot g0468(.din(w_n531_4[0]),.dout(n541),.clk(gclk));
	jand g0469(.dina(w_n541_1[2]),.dinb(n540),.dout(n542),.clk(gclk));
	jcb g0470(.dina(w_n542_0[1]),.dinb(w_n539_0[2]),.dout(G399));
	jand g0471(.dina(w_n90_1[1]),.dinb(w_n169_0[2]),.dout(n544),.clk(gclk));
	jand g0472(.dina(w_n544_0[2]),.dinb(w_n92_0[1]),.dout(n545),.clk(gclk));
	jcb g0473(.dina(w_n531_3[2]),.dinb(w_n513_0[0]),.dout(n546));
	jand g0474(.dina(w_n306_0[1]),.dinb(w_n191_1[1]),.dout(n547),.clk(gclk));
	jand g0475(.dina(w_n267_0[1]),.dinb(w_n243_0[0]),.dout(n548),.clk(gclk));
	jand g0476(.dina(n548),.dinb(w_n199_0[0]),.dout(n549),.clk(gclk));
	jand g0477(.dina(n549),.dinb(n547),.dout(n550),.clk(gclk));
	jnot g0478(.din(w_n200_0[0]),.dout(n551),.clk(gclk));
	jand g0479(.dina(w_n289_0[0]),.dinb(w_n221_0[1]),.dout(n552),.clk(gclk));
	jand g0480(.dina(w_dff_B_SW1uqonc9_0),.dinb(w_n327_0[1]),.dout(n553),.clk(gclk));
	jand g0481(.dina(n553),.dinb(w_dff_B_WHMoBw497_1),.dout(n554),.clk(gclk));
	jcb g0482(.dina(n554),.dinb(w_dff_B_a3L0F4cM6_1),.dout(n555));
	jcb g0483(.dina(n555),.dinb(w_n541_1[1]),.dout(n556));
	jcb g0484(.dina(w_n531_3[1]),.dinb(w_n338_0[0]),.dout(n557));
	jand g0485(.dina(n557),.dinb(w_dff_B_w0igAweX8_1),.dout(n558),.clk(gclk));
	jand g0486(.dina(n558),.dinb(w_G330_0[1]),.dout(n559),.clk(gclk));
	jnot g0487(.din(w_n559_1[2]),.dout(n560),.clk(gclk));
	jand g0488(.dina(n560),.dinb(w_n546_1[1]),.dout(n561),.clk(gclk));
	jnot g0489(.din(w_n561_1[1]),.dout(n562),.clk(gclk));
	jand g0490(.dina(n562),.dinb(w_n143_1[0]),.dout(n563),.clk(gclk));
	jnot g0491(.din(w_n544_0[1]),.dout(n564),.clk(gclk));
	jand g0492(.dina(w_n272_0[0]),.dinb(w_n112_0[2]),.dout(n565),.clk(gclk));
	jand g0493(.dina(w_n565_0[2]),.dinb(w_G1_0[2]),.dout(n566),.clk(gclk));
	jand g0494(.dina(n566),.dinb(w_n564_1[2]),.dout(n567),.clk(gclk));
	jcb g0495(.dina(w_dff_B_8R83VQXs5_0),.dinb(n563),.dout(n568));
	jcb g0496(.dina(n568),.dinb(w_dff_B_3w172eFQ5_1),.dout(G364));
	jand g0497(.dina(w_G45_0[2]),.dinb(w_G13_0[2]),.dout(n570),.clk(gclk));
	jcb g0498(.dina(n570),.dinb(w_n143_0[2]),.dout(n571));
	jand g0499(.dina(w_dff_B_Sj4KfGWI2_0),.dinb(w_n107_0[1]),.dout(n572),.clk(gclk));
	jnot g0500(.din(n572),.dout(n573),.clk(gclk));
	jand g0501(.dina(w_n573_1[2]),.dinb(w_n564_1[1]),.dout(n574),.clk(gclk));
	jnot g0502(.din(w_n574_4[1]),.dout(n575),.clk(gclk));
	jxor g0503(.dina(w_n534_0[0]),.dinb(w_G330_0[0]),.dout(n576),.clk(gclk));
	jand g0504(.dina(n576),.dinb(w_n575_0[2]),.dout(n577),.clk(gclk));
	jand g0505(.dina(w_n153_5[2]),.dinb(w_n88_0[0]),.dout(n578),.clk(gclk));
	jand g0506(.dina(w_n578_2[1]),.dinb(w_n151_1[1]),.dout(n579),.clk(gclk));
	jand g0507(.dina(w_n579_1[2]),.dinb(w_n533_0[0]),.dout(n580),.clk(gclk));
	jnot g0508(.din(n580),.dout(n581),.clk(gclk));
	jand g0509(.dina(w_G200_1[0]),.dinb(w_G20_3[0]),.dout(n582),.clk(gclk));
	jand g0510(.dina(w_n582_0[1]),.dinb(w_n191_1[0]),.dout(n583),.clk(gclk));
	jand g0511(.dina(w_n583_0[1]),.dinb(w_n284_1[1]),.dout(n584),.clk(gclk));
	jand g0512(.dina(w_n584_4[1]),.dinb(w_G107_2[2]),.dout(n585),.clk(gclk));
	jand g0513(.dina(w_G179_0[1]),.dinb(w_G20_2[2]),.dout(n586),.clk(gclk));
	jand g0514(.dina(w_n586_0[2]),.dinb(w_G200_0[2]),.dout(n587),.clk(gclk));
	jand g0515(.dina(w_n587_0[1]),.dinb(w_G190_2[0]),.dout(n588),.clk(gclk));
	jand g0516(.dina(w_n588_7[1]),.dinb(w_G50_4[2]),.dout(n589),.clk(gclk));
	jcb g0517(.dina(n589),.dinb(w_n585_0[1]),.dout(n590));
	jcb g0518(.dina(n590),.dinb(w_G33_6[1]),.dout(n591));
	jand g0519(.dina(w_n587_0[0]),.dinb(w_n284_1[0]),.dout(n592),.clk(gclk));
	jand g0520(.dina(w_n592_7[1]),.dinb(w_G68_3[2]),.dout(n593),.clk(gclk));
	jand g0521(.dina(w_n583_0[0]),.dinb(w_G190_1[2]),.dout(n594),.clk(gclk));
	jand g0522(.dina(w_n594_6[1]),.dinb(w_G87_2[2]),.dout(n595),.clk(gclk));
	jcb g0523(.dina(w_n595_0[1]),.dinb(n593),.dout(n596));
	jand g0524(.dina(w_n586_0[1]),.dinb(w_n251_0[2]),.dout(n597),.clk(gclk));
	jand g0525(.dina(w_n597_0[1]),.dinb(w_G190_1[1]),.dout(n598),.clk(gclk));
	jand g0526(.dina(w_n598_7[1]),.dinb(w_G58_4[1]),.dout(n599),.clk(gclk));
	jand g0527(.dina(w_n284_0[2]),.dinb(w_G20_2[1]),.dout(n600),.clk(gclk));
	jcb g0528(.dina(w_n586_0[0]),.dinb(w_n582_0[0]),.dout(n601));
	jnot g0529(.din(w_n601_0[1]),.dout(n602),.clk(gclk));
	jand g0530(.dina(n602),.dinb(w_n600_0[1]),.dout(n603),.clk(gclk));
	jand g0531(.dina(w_n603_7[1]),.dinb(w_G159_3[1]),.dout(n604),.clk(gclk));
	jcb g0532(.dina(n604),.dinb(n599),.dout(n605));
	jcb g0533(.dina(w_n601_0[0]),.dinb(w_n600_0[0]),.dout(n606));
	jnot g0534(.din(n606),.dout(n607),.clk(gclk));
	jand g0535(.dina(w_n607_5[1]),.dinb(w_G97_3[1]),.dout(n608),.clk(gclk));
	jand g0536(.dina(w_n597_0[0]),.dinb(w_n284_0[1]),.dout(n609),.clk(gclk));
	jand g0537(.dina(w_n609_7[1]),.dinb(w_G77_3[0]),.dout(n610),.clk(gclk));
	jcb g0538(.dina(n610),.dinb(w_n608_0[1]),.dout(n611));
	jcb g0539(.dina(n611),.dinb(n605),.dout(n612));
	jcb g0540(.dina(n612),.dinb(n596),.dout(n613));
	jcb g0541(.dina(n613),.dinb(n591),.dout(n614));
	jand g0542(.dina(w_n594_6[0]),.dinb(w_G303_2[1]),.dout(n615),.clk(gclk));
	jand g0543(.dina(w_n584_4[0]),.dinb(w_G283_3[1]),.dout(n616),.clk(gclk));
	jand g0544(.dina(w_n609_7[0]),.dinb(w_G311_1[2]),.dout(n617),.clk(gclk));
	jcb g0545(.dina(n617),.dinb(n616),.dout(n618));
	jand g0546(.dina(w_n607_5[0]),.dinb(w_G294_3[0]),.dout(n619),.clk(gclk));
	jcb g0547(.dina(n619),.dinb(n618),.dout(n620));
	jand g0548(.dina(w_n603_7[0]),.dinb(w_dff_B_GXaL3ZsG0_1),.dout(n621),.clk(gclk));
	jand g0549(.dina(w_n598_7[0]),.dinb(w_G322_0[2]),.dout(n622),.clk(gclk));
	jand g0550(.dina(w_n592_7[0]),.dinb(w_G317_1[1]),.dout(n623),.clk(gclk));
	jcb g0551(.dina(n623),.dinb(n622),.dout(n624));
	jand g0552(.dina(w_n588_7[0]),.dinb(w_G326_0[1]),.dout(n625),.clk(gclk));
	jcb g0553(.dina(n625),.dinb(w_n153_5[1]),.dout(n626));
	jcb g0554(.dina(n626),.dinb(n624),.dout(n627));
	jcb g0555(.dina(n627),.dinb(n621),.dout(n628));
	jcb g0556(.dina(n628),.dinb(n620),.dout(n629));
	jcb g0557(.dina(n629),.dinb(n615),.dout(n630));
	jand g0558(.dina(n630),.dinb(n614),.dout(n631),.clk(gclk));
	jand g0559(.dina(w_n140_0[1]),.dinb(w_G169_0[2]),.dout(n632),.clk(gclk));
	jcb g0560(.dina(n632),.dinb(w_n362_0[0]),.dout(n633));
	jnot g0561(.din(n633),.dout(n634),.clk(gclk));
	jcb g0562(.dina(w_n634_4[1]),.dinb(n631),.dout(n635));
	jnot g0563(.din(w_n579_1[1]),.dout(n636),.clk(gclk));
	jand g0564(.dina(w_n634_4[0]),.dinb(n636),.dout(n637),.clk(gclk));
	jcb g0565(.dina(w_n135_0[0]),.dinb(w_n339_1[0]),.dout(n638));
	jand g0566(.dina(w_n90_1[0]),.dinb(w_G33_6[0]),.dout(n639),.clk(gclk));
	jnot g0567(.din(w_n639_0[2]),.dout(n640),.clk(gclk));
	jand g0568(.dina(w_n92_0[0]),.dinb(w_n339_0[2]),.dout(n641),.clk(gclk));
	jcb g0569(.dina(w_dff_B_frWjfpCC8_0),.dinb(w_n640_0[1]),.dout(n642));
	jnot g0570(.din(n642),.dout(n643),.clk(gclk));
	jand g0571(.dina(n643),.dinb(w_dff_B_3i0omfmu0_1),.dout(n644),.clk(gclk));
	jnot g0572(.din(w_n90_0[2]),.dout(n645),.clk(gclk));
	jand g0573(.dina(w_n645_1[1]),.dinb(w_n112_0[1]),.dout(n646),.clk(gclk));
	jand g0574(.dina(w_n90_0[1]),.dinb(w_n153_5[0]),.dout(n647),.clk(gclk));
	jand g0575(.dina(w_n647_0[1]),.dinb(w_G355_0),.dout(n648),.clk(gclk));
	jcb g0576(.dina(n648),.dinb(n646),.dout(n649));
	jcb g0577(.dina(w_dff_B_Y9mIcjJJ2_0),.dinb(n644),.dout(n650));
	jand g0578(.dina(n650),.dinb(w_n637_0[1]),.dout(n651),.clk(gclk));
	jnot g0579(.din(n651),.dout(n652),.clk(gclk));
	jand g0580(.dina(n652),.dinb(w_dff_B_vNQOvYjL3_1),.dout(n653),.clk(gclk));
	jand g0581(.dina(w_dff_B_aPDOq9fw2_0),.dinb(n581),.dout(n654),.clk(gclk));
	jand g0582(.dina(n654),.dinb(w_n574_4[0]),.dout(n655),.clk(gclk));
	jcb g0583(.dina(n655),.dinb(w_dff_B_k3R0GRDO1_1),.dout(G396_fa_));
	jand g0584(.dina(w_n531_3[0]),.dinb(w_n370_0[0]),.dout(n657),.clk(gclk));
	jxor g0585(.dina(w_dff_B_yXkkCsrs6_0),.dinb(w_n381_0[1]),.dout(n658),.clk(gclk));
	jand g0586(.dina(w_n658_0[2]),.dinb(w_n578_2[0]),.dout(n659),.clk(gclk));
	jnot g0587(.din(n659),.dout(n660),.clk(gclk));
	jnot g0588(.din(w_n578_1[2]),.dout(n661),.clk(gclk));
	jand g0589(.dina(w_n634_3[2]),.dinb(n661),.dout(n662),.clk(gclk));
	jand g0590(.dina(w_n662_1[1]),.dinb(w_n73_0[1]),.dout(n663),.clk(gclk));
	jnot g0591(.din(n663),.dout(n664),.clk(gclk));
	jand g0592(.dina(w_n588_6[2]),.dinb(w_G303_2[0]),.dout(n665),.clk(gclk));
	jand g0593(.dina(w_n598_6[2]),.dinb(w_G294_2[2]),.dout(n666),.clk(gclk));
	jcb g0594(.dina(n666),.dinb(n665),.dout(n667));
	jand g0595(.dina(w_n592_6[2]),.dinb(w_G283_3[0]),.dout(n668),.clk(gclk));
	jcb g0596(.dina(n668),.dinb(n667),.dout(n669));
	jand g0597(.dina(w_n594_5[2]),.dinb(w_G107_2[1]),.dout(n670),.clk(gclk));
	jcb g0598(.dina(n670),.dinb(w_n153_4[2]),.dout(n671));
	jcb g0599(.dina(n671),.dinb(w_n608_0[0]),.dout(n672));
	jand g0600(.dina(w_n609_6[2]),.dinb(w_G116_4[0]),.dout(n673),.clk(gclk));
	jand g0601(.dina(w_n584_3[2]),.dinb(w_G87_2[1]),.dout(n674),.clk(gclk));
	jcb g0602(.dina(w_n674_0[1]),.dinb(n673),.dout(n675));
	jand g0603(.dina(w_n603_6[2]),.dinb(w_G311_1[1]),.dout(n676),.clk(gclk));
	jcb g0604(.dina(n676),.dinb(n675),.dout(n677));
	jcb g0605(.dina(n677),.dinb(n672),.dout(n678));
	jcb g0606(.dina(n678),.dinb(n669),.dout(n679));
	jand g0607(.dina(w_n598_6[1]),.dinb(w_G143_2[1]),.dout(n680),.clk(gclk));
	jand g0608(.dina(w_n603_6[1]),.dinb(w_G132_1[1]),.dout(n681),.clk(gclk));
	jcb g0609(.dina(n681),.dinb(n680),.dout(n682));
	jand g0610(.dina(w_n592_6[1]),.dinb(w_G150_3[0]),.dout(n683),.clk(gclk));
	jand g0611(.dina(w_n607_4[2]),.dinb(w_G58_4[0]),.dout(n684),.clk(gclk));
	jcb g0612(.dina(n684),.dinb(n683),.dout(n685));
	jcb g0613(.dina(n685),.dinb(n682),.dout(n686));
	jand g0614(.dina(w_n584_3[1]),.dinb(w_G68_3[1]),.dout(n687),.clk(gclk));
	jand g0615(.dina(w_n588_6[1]),.dinb(w_G137_1[2]),.dout(n688),.clk(gclk));
	jcb g0616(.dina(n688),.dinb(w_n687_0[1]),.dout(n689));
	jand g0617(.dina(w_n594_5[1]),.dinb(w_G50_4[1]),.dout(n690),.clk(gclk));
	jand g0618(.dina(w_n609_6[1]),.dinb(w_G159_3[0]),.dout(n691),.clk(gclk));
	jcb g0619(.dina(n691),.dinb(n690),.dout(n692));
	jcb g0620(.dina(n692),.dinb(w_G33_5[2]),.dout(n693));
	jcb g0621(.dina(n693),.dinb(n689),.dout(n694));
	jcb g0622(.dina(n694),.dinb(n686),.dout(n695));
	jand g0623(.dina(n695),.dinb(n679),.dout(n696),.clk(gclk));
	jcb g0624(.dina(n696),.dinb(w_n634_3[1]),.dout(n697));
	jand g0625(.dina(w_dff_B_n51VEqSr3_0),.dinb(n664),.dout(n698),.clk(gclk));
	jand g0626(.dina(n698),.dinb(w_n574_3[2]),.dout(n699),.clk(gclk));
	jand g0627(.dina(w_dff_B_lorWBVYy3_0),.dinb(n660),.dout(n700),.clk(gclk));
	jcb g0628(.dina(w_n546_1[0]),.dinb(w_n381_0[0]),.dout(n701));
	jnot g0629(.din(w_n546_0[2]),.dout(n702),.clk(gclk));
	jnot g0630(.din(w_n658_0[1]),.dout(n703),.clk(gclk));
	jcb g0631(.dina(w_n703_0[2]),.dinb(n702),.dout(n704));
	jand g0632(.dina(n704),.dinb(w_n701_0[1]),.dout(n705),.clk(gclk));
	jxor g0633(.dina(n705),.dinb(w_n559_1[1]),.dout(n706),.clk(gclk));
	jand g0634(.dina(n706),.dinb(w_n575_0[1]),.dout(n707),.clk(gclk));
	jcb g0635(.dina(n707),.dinb(w_dff_B_UqFtJkCs7_1),.dout(G384_fa_));
	jnot g0636(.din(w_n89_0[1]),.dout(n709),.clk(gclk));
	jand g0637(.dina(w_n107_0[0]),.dinb(n709),.dout(n710),.clk(gclk));
	jnot g0638(.din(w_n476_0[0]),.dout(n711),.clk(gclk));
	jcb g0639(.dina(w_n530_1[0]),.dinb(n711),.dout(n712));
	jand g0640(.dina(w_n530_0[2]),.dinb(w_n478_0[0]),.dout(n713),.clk(gclk));
	jxor g0641(.dina(w_dff_B_kWlhMqib3_0),.dinb(w_n483_0[0]),.dout(n714),.clk(gclk));
	jcb g0642(.dina(w_n531_2[2]),.dinb(w_n520_0[0]),.dout(n715));
	jand g0643(.dina(w_n541_1[0]),.dinb(w_n375_0[0]),.dout(n716),.clk(gclk));
	jnot g0644(.din(n716),.dout(n717),.clk(gclk));
	jand g0645(.dina(w_n717_0[1]),.dinb(w_n701_0[0]),.dout(n718),.clk(gclk));
	jnot g0646(.din(w_n406_0[0]),.dout(n719),.clk(gclk));
	jand g0647(.dina(w_n531_2[1]),.dinb(n719),.dout(n720),.clk(gclk));
	jxor g0648(.dina(n720),.dinb(w_n415_0[2]),.dout(n721),.clk(gclk));
	jcb g0649(.dina(w_n721_1[1]),.dinb(w_n718_0[2]),.dout(n722));
	jand g0650(.dina(n722),.dinb(w_n715_0[1]),.dout(n723),.clk(gclk));
	jcb g0651(.dina(n723),.dinb(w_n714_0[2]),.dout(n724));
	jand g0652(.dina(n724),.dinb(w_dff_B_Keavc4sM0_1),.dout(n725),.clk(gclk));
	jnot g0653(.din(w_n714_0[1]),.dout(n726),.clk(gclk));
	jnot g0654(.din(w_n721_1[0]),.dout(n727),.clk(gclk));
	jand g0655(.dina(w_n727_0[2]),.dinb(w_n726_0[1]),.dout(n728),.clk(gclk));
	jand g0656(.dina(n728),.dinb(w_n703_0[1]),.dout(n729),.clk(gclk));
	jand g0657(.dina(w_n729_0[1]),.dinb(w_n559_1[0]),.dout(n730),.clk(gclk));
	jnot g0658(.din(n730),.dout(n731),.clk(gclk));
	jcb g0659(.dina(w_n731_0[1]),.dinb(w_n487_0[1]),.dout(n732));
	jand g0660(.dina(w_n559_0[2]),.dinb(w_n487_0[0]),.dout(n733),.clk(gclk));
	jnot g0661(.din(n733),.dout(n734),.clk(gclk));
	jcb g0662(.dina(w_n734_0[1]),.dinb(w_n729_0[0]),.dout(n735));
	jand g0663(.dina(n735),.dinb(n732),.dout(n736),.clk(gclk));
	jcb g0664(.dina(w_n531_2[0]),.dinb(w_n514_0[0]),.dout(n737));
	jand g0665(.dina(n737),.dinb(w_n525_0[0]),.dout(n738),.clk(gclk));
	jnot g0666(.din(w_n738_0[1]),.dout(n739),.clk(gclk));
	jxor g0667(.dina(w_dff_B_HxkD4b9J1_0),.dinb(n736),.dout(n740),.clk(gclk));
	jxor g0668(.dina(n740),.dinb(w_n725_0[1]),.dout(n741),.clk(gclk));
	jand g0669(.dina(n741),.dinb(w_dff_B_C0KWpf0w3_1),.dout(n742),.clk(gclk));
	jcb g0670(.dina(w_n103_0[2]),.dinb(w_n108_0[2]),.dout(n743));
	jand g0671(.dina(n743),.dinb(w_G77_2[2]),.dout(n744),.clk(gclk));
	jcb g0672(.dina(n744),.dinb(w_n99_1[0]),.dout(n745));
	jand g0673(.dina(w_G58_3[2]),.dinb(w_G50_4[0]),.dout(n746),.clk(gclk));
	jcb g0674(.dina(n746),.dinb(w_G68_3[0]),.dout(n747));
	jand g0675(.dina(w_dff_B_fX66LWDV4_0),.dinb(w_n89_0[0]),.dout(n748),.clk(gclk));
	jand g0676(.dina(n748),.dinb(w_dff_B_LzkS9f5x3_1),.dout(n749),.clk(gclk));
	jand g0677(.dina(w_n309_0[0]),.dinb(w_n95_0[0]),.dout(n750),.clk(gclk));
	jand g0678(.dina(n750),.dinb(w_G116_3[2]),.dout(n751),.clk(gclk));
	jcb g0679(.dina(n751),.dinb(n749),.dout(n752));
	jcb g0680(.dina(w_dff_B_rSUdwkVl7_0),.dinb(n742),.dout(G367));
	jand g0681(.dina(w_n531_1[2]),.dinb(w_n320_0[1]),.dout(n754),.clk(gclk));
	jxor g0682(.dina(w_dff_B_fRfLC7wP3_0),.dinb(w_n506_0[0]),.dout(n755),.clk(gclk));
	jnot g0683(.din(w_n755_0[2]),.dout(n756),.clk(gclk));
	jand g0684(.dina(w_dff_B_lJMPZ3y32_0),.dinb(w_n539_0[1]),.dout(n757),.clk(gclk));
	jand g0685(.dina(w_n334_0[0]),.dinb(w_n246_0[0]),.dout(n758),.clk(gclk));
	jcb g0686(.dina(n758),.dinb(w_n501_0[0]),.dout(n759));
	jnot g0687(.din(w_n202_0[0]),.dout(n760),.clk(gclk));
	jand g0688(.dina(w_n538_0[1]),.dinb(w_n335_0[0]),.dout(n761),.clk(gclk));
	jand g0689(.dina(n761),.dinb(w_n760_0[1]),.dout(n762),.clk(gclk));
	jcb g0690(.dina(n762),.dinb(w_dff_B_iYrA9RZ57_1),.dout(n763));
	jand g0691(.dina(n763),.dinb(w_n541_0[2]),.dout(n764),.clk(gclk));
	jnot g0692(.din(w_n764_0[1]),.dout(n765),.clk(gclk));
	jcb g0693(.dina(n765),.dinb(w_n295_0[0]),.dout(n766));
	jand g0694(.dina(w_n531_1[1]),.dinb(w_n283_0[1]),.dout(n767),.clk(gclk));
	jxor g0695(.dina(w_dff_B_bZqFMHI27_0),.dinb(w_n497_0[0]),.dout(n768),.clk(gclk));
	jcb g0696(.dina(w_n768_0[1]),.dinb(w_n764_0[0]),.dout(n769));
	jand g0697(.dina(w_dff_B_gyCkCVW80_0),.dinb(n766),.dout(n770),.clk(gclk));
	jxor g0698(.dina(n770),.dinb(w_dff_B_gj7NzOOx8_1),.dout(n771),.clk(gclk));
	jcb g0699(.dina(w_n771_0[1]),.dinb(w_n573_1[1]),.dout(n772));
	jand g0700(.dina(w_n768_0[0]),.dinb(w_n579_1[0]),.dout(n773),.clk(gclk));
	jnot g0701(.din(n773),.dout(n774),.clk(gclk));
	jand g0702(.dina(w_n609_6[0]),.dinb(w_G50_3[2]),.dout(n775),.clk(gclk));
	jand g0703(.dina(w_n592_6[0]),.dinb(w_G159_2[2]),.dout(n776),.clk(gclk));
	jcb g0704(.dina(n776),.dinb(n775),.dout(n777));
	jand g0705(.dina(w_n607_4[1]),.dinb(w_G68_2[2]),.dout(n778),.clk(gclk));
	jand g0706(.dina(w_n598_6[0]),.dinb(w_G150_2[2]),.dout(n779),.clk(gclk));
	jand g0707(.dina(w_n584_3[0]),.dinb(w_G77_2[1]),.dout(n780),.clk(gclk));
	jcb g0708(.dina(w_n780_0[1]),.dinb(n779),.dout(n781));
	jcb g0709(.dina(n781),.dinb(w_n778_0[1]),.dout(n782));
	jand g0710(.dina(w_n603_6[0]),.dinb(w_G137_1[1]),.dout(n783),.clk(gclk));
	jand g0711(.dina(w_n588_6[0]),.dinb(w_G143_2[0]),.dout(n784),.clk(gclk));
	jcb g0712(.dina(n784),.dinb(n783),.dout(n785));
	jand g0713(.dina(w_n594_5[0]),.dinb(w_G58_3[1]),.dout(n786),.clk(gclk));
	jcb g0714(.dina(n786),.dinb(w_G33_5[1]),.dout(n787));
	jcb g0715(.dina(n787),.dinb(n785),.dout(n788));
	jcb g0716(.dina(n788),.dinb(n782),.dout(n789));
	jcb g0717(.dina(n789),.dinb(n777),.dout(n790));
	jand g0718(.dina(w_n607_4[0]),.dinb(w_G107_2[0]),.dout(n791),.clk(gclk));
	jand g0719(.dina(w_n588_5[2]),.dinb(w_G311_1[0]),.dout(n792),.clk(gclk));
	jcb g0720(.dina(n792),.dinb(w_n153_4[1]),.dout(n793));
	jcb g0721(.dina(n793),.dinb(n791),.dout(n794));
	jand g0722(.dina(w_n598_5[2]),.dinb(w_G303_1[2]),.dout(n795),.clk(gclk));
	jand g0723(.dina(w_n592_5[2]),.dinb(w_G294_2[1]),.dout(n796),.clk(gclk));
	jcb g0724(.dina(n796),.dinb(n795),.dout(n797));
	jand g0725(.dina(w_n609_5[2]),.dinb(w_G283_2[2]),.dout(n798),.clk(gclk));
	jcb g0726(.dina(n798),.dinb(n797),.dout(n799));
	jand g0727(.dina(w_n594_4[2]),.dinb(w_G116_3[1]),.dout(n800),.clk(gclk));
	jand g0728(.dina(w_n584_2[2]),.dinb(w_G97_3[0]),.dout(n801),.clk(gclk));
	jcb g0729(.dina(w_n801_0[1]),.dinb(n800),.dout(n802));
	jand g0730(.dina(w_n603_5[2]),.dinb(w_G317_1[0]),.dout(n803),.clk(gclk));
	jcb g0731(.dina(n803),.dinb(n802),.dout(n804));
	jcb g0732(.dina(n804),.dinb(n799),.dout(n805));
	jcb g0733(.dina(n805),.dinb(n794),.dout(n806));
	jand g0734(.dina(n806),.dinb(n790),.dout(n807),.clk(gclk));
	jcb g0735(.dina(n807),.dinb(w_n634_3[0]),.dout(n808));
	jand g0736(.dina(w_n645_1[0]),.dinb(w_G87_2[0]),.dout(n809),.clk(gclk));
	jnot g0737(.din(w_n637_0[0]),.dout(n810),.clk(gclk));
	jand g0738(.dina(w_n639_0[1]),.dinb(w_n127_0[0]),.dout(n811),.clk(gclk));
	jcb g0739(.dina(w_dff_B_7nbBkGuI5_0),.dinb(w_n810_0[2]),.dout(n812));
	jcb g0740(.dina(n812),.dinb(w_dff_B_3DYUwprA2_1),.dout(n813));
	jand g0741(.dina(n813),.dinb(w_dff_B_CX9qtM3w1_1),.dout(n814),.clk(gclk));
	jand g0742(.dina(w_dff_B_erdOwoPR9_0),.dinb(n774),.dout(n815),.clk(gclk));
	jand g0743(.dina(n815),.dinb(w_n574_3[1]),.dout(n816),.clk(gclk));
	jnot g0744(.din(n816),.dout(n817),.clk(gclk));
	jand g0745(.dina(w_dff_B_7uTgNvTx3_0),.dinb(n772),.dout(n818),.clk(gclk));
	jand g0746(.dina(w_n541_0[1]),.dinb(w_n760_0[0]),.dout(n819),.clk(gclk));
	jcb g0747(.dina(w_n819_0[1]),.dinb(w_n538_0[0]),.dout(n820));
	jnot g0748(.din(w_n819_0[0]),.dout(n821),.clk(gclk));
	jcb g0749(.dina(n821),.dinb(w_n255_0[1]),.dout(n822));
	jand g0750(.dina(n822),.dinb(n820),.dout(n823),.clk(gclk));
	jxor g0751(.dina(w_dff_B_zkwCK5Dw6_0),.dinb(w_n535_0[0]),.dout(n824),.clk(gclk));
	jnot g0752(.din(w_n824_0[2]),.dout(n825),.clk(gclk));
	jxor g0753(.dina(w_n542_0[0]),.dinb(w_n539_0[0]),.dout(n826),.clk(gclk));
	jxor g0754(.dina(n826),.dinb(w_n755_0[1]),.dout(n827),.clk(gclk));
	jcb g0755(.dina(w_n827_0[2]),.dinb(w_n825_0[1]),.dout(n828));
	jand g0756(.dina(w_dff_B_iPrd9TeX5_0),.dinb(w_n561_1[0]),.dout(n829),.clk(gclk));
	jcb g0757(.dina(n829),.dinb(w_n564_1[0]),.dout(n830));
	jcb g0758(.dina(n830),.dinb(w_n771_0[0]),.dout(n831));
	jand g0759(.dina(n831),.dinb(n818),.dout(n832),.clk(gclk));
	jnot g0760(.din(w_n832_0[2]),.dout(G387),.clk(gclk));
	jand g0761(.dina(w_n561_0[2]),.dinb(w_n544_0[0]),.dout(n834),.clk(gclk));
	jnot g0762(.din(w_n834_0[1]),.dout(n835),.clk(gclk));
	jand g0763(.dina(n835),.dinb(w_n825_0[0]),.dout(n836),.clk(gclk));
	jand g0764(.dina(w_n824_0[1]),.dinb(w_n561_0[1]),.dout(n837),.clk(gclk));
	jand g0765(.dina(n837),.dinb(w_n573_1[0]),.dout(n838),.clk(gclk));
	jcb g0766(.dina(n838),.dinb(w_n574_3[0]),.dout(n839));
	jcb g0767(.dina(w_n839_0[1]),.dinb(n836),.dout(n840));
	jand g0768(.dina(w_n579_0[2]),.dinb(w_n537_0[0]),.dout(n841),.clk(gclk));
	jnot g0769(.din(n841),.dout(n842),.clk(gclk));
	jand g0770(.dina(w_n603_5[1]),.dinb(w_G326_0[0]),.dout(n843),.clk(gclk));
	jand g0771(.dina(w_n584_2[1]),.dinb(w_G116_3[0]),.dout(n844),.clk(gclk));
	jand g0772(.dina(w_n594_4[1]),.dinb(w_G294_2[0]),.dout(n845),.clk(gclk));
	jcb g0773(.dina(n845),.dinb(n844),.dout(n846));
	jand g0774(.dina(w_n607_3[2]),.dinb(w_G283_2[1]),.dout(n847),.clk(gclk));
	jcb g0775(.dina(n847),.dinb(n846),.dout(n848));
	jcb g0776(.dina(n848),.dinb(n843),.dout(n849));
	jand g0777(.dina(w_n588_5[1]),.dinb(w_G322_0[1]),.dout(n850),.clk(gclk));
	jcb g0778(.dina(n850),.dinb(w_n153_4[0]),.dout(n851));
	jand g0779(.dina(w_n598_5[1]),.dinb(w_G317_0[2]),.dout(n852),.clk(gclk));
	jand g0780(.dina(w_n592_5[1]),.dinb(w_G311_0[2]),.dout(n853),.clk(gclk));
	jcb g0781(.dina(n853),.dinb(n852),.dout(n854));
	jand g0782(.dina(w_n609_5[1]),.dinb(w_G303_1[1]),.dout(n855),.clk(gclk));
	jcb g0783(.dina(n855),.dinb(n854),.dout(n856));
	jcb g0784(.dina(n856),.dinb(n851),.dout(n857));
	jcb g0785(.dina(n857),.dinb(n849),.dout(n858));
	jand g0786(.dina(w_n607_3[1]),.dinb(w_G87_1[2]),.dout(n859),.clk(gclk));
	jand g0787(.dina(w_n609_5[0]),.dinb(w_G68_2[1]),.dout(n860),.clk(gclk));
	jand g0788(.dina(w_n598_5[0]),.dinb(w_G50_3[1]),.dout(n861),.clk(gclk));
	jcb g0789(.dina(n861),.dinb(n860),.dout(n862));
	jand g0790(.dina(w_n592_5[0]),.dinb(w_G58_3[0]),.dout(n863),.clk(gclk));
	jcb g0791(.dina(n863),.dinb(w_G33_5[0]),.dout(n864));
	jcb g0792(.dina(n864),.dinb(n862),.dout(n865));
	jand g0793(.dina(w_n594_4[0]),.dinb(w_G77_2[0]),.dout(n866),.clk(gclk));
	jcb g0794(.dina(w_n866_0[1]),.dinb(w_n801_0[0]),.dout(n867));
	jand g0795(.dina(w_n588_5[0]),.dinb(w_G159_2[1]),.dout(n868),.clk(gclk));
	jand g0796(.dina(w_n603_5[0]),.dinb(w_G150_2[1]),.dout(n869),.clk(gclk));
	jcb g0797(.dina(n869),.dinb(n868),.dout(n870));
	jcb g0798(.dina(n870),.dinb(n867),.dout(n871));
	jcb g0799(.dina(n871),.dinb(n865),.dout(n872));
	jcb g0800(.dina(n872),.dinb(w_n859_0[1]),.dout(n873));
	jand g0801(.dina(n873),.dinb(n858),.dout(n874),.clk(gclk));
	jcb g0802(.dina(n874),.dinb(w_n634_2[2]),.dout(n875));
	jand g0803(.dina(w_n645_0[2]),.dinb(w_n80_0[2]),.dout(n876),.clk(gclk));
	jnot g0804(.din(n876),.dout(n877),.clk(gclk));
	jnot g0805(.din(w_n565_0[1]),.dout(n878),.clk(gclk));
	jand g0806(.dina(w_n647_0[0]),.dinb(n878),.dout(n879),.clk(gclk));
	jnot g0807(.din(n879),.dout(n880),.clk(gclk));
	jand g0808(.dina(w_n131_0[0]),.dinb(w_G45_0[1]),.dout(n881),.clk(gclk));
	jcb g0809(.dina(w_dff_B_YqXng1Tl4_0),.dinb(w_n640_0[0]),.dout(n882));
	jand g0810(.dina(w_dff_B_zJiB3lEY7_0),.dinb(n880),.dout(n883),.clk(gclk));
	jand g0811(.dina(w_G77_1[2]),.dinb(w_G68_2[0]),.dout(n884),.clk(gclk));
	jnot g0812(.din(n884),.dout(n885),.clk(gclk));
	jand g0813(.dina(w_G58_2[2]),.dinb(w_n99_0[2]),.dout(n886),.clk(gclk));
	jand g0814(.dina(n886),.dinb(n885),.dout(n887),.clk(gclk));
	jand g0815(.dina(w_dff_B_rVv7XDPP0_0),.dinb(w_n565_0[0]),.dout(n888),.clk(gclk));
	jand g0816(.dina(n888),.dinb(w_n339_0[1]),.dout(n889),.clk(gclk));
	jcb g0817(.dina(w_dff_B_F3XZmJmq0_0),.dinb(n883),.dout(n890));
	jand g0818(.dina(n890),.dinb(w_dff_B_LlUIFToS7_1),.dout(n891),.clk(gclk));
	jcb g0819(.dina(n891),.dinb(w_n810_0[1]),.dout(n892));
	jand g0820(.dina(n892),.dinb(w_dff_B_ELOV9xVH7_1),.dout(n893),.clk(gclk));
	jand g0821(.dina(w_dff_B_uVYZmFoa2_0),.dinb(n842),.dout(n894),.clk(gclk));
	jand g0822(.dina(n894),.dinb(w_n574_2[2]),.dout(n895),.clk(gclk));
	jnot g0823(.din(n895),.dout(n896),.clk(gclk));
	jand g0824(.dina(w_dff_B_popybWGT3_0),.dinb(n840),.dout(n897),.clk(gclk));
	jnot g0825(.din(w_n897_0[2]),.dout(G393),.clk(gclk));
	jand g0826(.dina(w_n755_0[0]),.dinb(w_n579_0[1]),.dout(n899),.clk(gclk));
	jnot g0827(.din(n899),.dout(n900),.clk(gclk));
	jand g0828(.dina(w_n645_0[1]),.dinb(w_G97_2[2]),.dout(n901),.clk(gclk));
	jand g0829(.dina(w_n639_0[0]),.dinb(w_n138_0[0]),.dout(n902),.clk(gclk));
	jcb g0830(.dina(w_dff_B_D5X8rJBq2_0),.dinb(w_n810_0[0]),.dout(n903));
	jcb g0831(.dina(n903),.dinb(w_dff_B_QSPc2gnM7_1),.dout(n904));
	jand g0832(.dina(w_n609_4[2]),.dinb(w_G58_2[1]),.dout(n905),.clk(gclk));
	jand g0833(.dina(w_n598_4[2]),.dinb(w_G159_2[0]),.dout(n906),.clk(gclk));
	jcb g0834(.dina(n906),.dinb(n905),.dout(n907));
	jand g0835(.dina(w_n594_3[2]),.dinb(w_G68_1[2]),.dout(n908),.clk(gclk));
	jand g0836(.dina(w_n588_4[2]),.dinb(w_G150_2[0]),.dout(n909),.clk(gclk));
	jand g0837(.dina(w_n603_4[2]),.dinb(w_G143_1[2]),.dout(n910),.clk(gclk));
	jcb g0838(.dina(n910),.dinb(n909),.dout(n911));
	jcb g0839(.dina(n911),.dinb(n908),.dout(n912));
	jand g0840(.dina(w_n607_3[0]),.dinb(w_G77_1[1]),.dout(n913),.clk(gclk));
	jcb g0841(.dina(w_n913_0[1]),.dinb(w_n674_0[0]),.dout(n914));
	jand g0842(.dina(w_n592_4[2]),.dinb(w_G50_3[0]),.dout(n915),.clk(gclk));
	jcb g0843(.dina(n915),.dinb(w_G33_4[2]),.dout(n916));
	jcb g0844(.dina(n916),.dinb(n914),.dout(n917));
	jcb g0845(.dina(n917),.dinb(n912),.dout(n918));
	jcb g0846(.dina(n918),.dinb(n907),.dout(n919));
	jand g0847(.dina(w_n594_3[1]),.dinb(w_G283_2[0]),.dout(n920),.clk(gclk));
	jcb g0848(.dina(n920),.dinb(w_n153_3[2]),.dout(n921));
	jcb g0849(.dina(n921),.dinb(w_n585_0[0]),.dout(n922));
	jand g0850(.dina(w_n588_4[1]),.dinb(w_G317_0[1]),.dout(n923),.clk(gclk));
	jand g0851(.dina(w_n598_4[1]),.dinb(w_G311_0[1]),.dout(n924),.clk(gclk));
	jcb g0852(.dina(n924),.dinb(n923),.dout(n925));
	jand g0853(.dina(w_n603_4[1]),.dinb(w_G322_0[0]),.dout(n926),.clk(gclk));
	jcb g0854(.dina(n926),.dinb(n925),.dout(n927));
	jand g0855(.dina(w_n592_4[1]),.dinb(w_G303_1[0]),.dout(n928),.clk(gclk));
	jand g0856(.dina(w_n607_2[2]),.dinb(w_G116_2[2]),.dout(n929),.clk(gclk));
	jcb g0857(.dina(n929),.dinb(n928),.dout(n930));
	jand g0858(.dina(w_n609_4[1]),.dinb(w_G294_1[2]),.dout(n931),.clk(gclk));
	jcb g0859(.dina(n931),.dinb(n930),.dout(n932));
	jcb g0860(.dina(n932),.dinb(n927),.dout(n933));
	jcb g0861(.dina(n933),.dinb(n922),.dout(n934));
	jand g0862(.dina(n934),.dinb(n919),.dout(n935),.clk(gclk));
	jcb g0863(.dina(n935),.dinb(w_n634_2[1]),.dout(n936));
	jand g0864(.dina(w_dff_B_SzLMeSQE7_0),.dinb(w_n574_2[1]),.dout(n937),.clk(gclk));
	jand g0865(.dina(n937),.dinb(w_dff_B_ShVlZ9431_1),.dout(n938),.clk(gclk));
	jand g0866(.dina(w_dff_B_ALmO11cs1_0),.dinb(n900),.dout(n939),.clk(gclk));
	jnot g0867(.din(n939),.dout(n940),.clk(gclk));
	jcb g0868(.dina(w_n839_0[0]),.dinb(w_n827_0[1]),.dout(n941));
	jand g0869(.dina(w_n834_0[0]),.dinb(w_n827_0[0]),.dout(n942),.clk(gclk));
	jand g0870(.dina(n942),.dinb(w_n824_0[0]),.dout(n943),.clk(gclk));
	jnot g0871(.din(n943),.dout(n944),.clk(gclk));
	jand g0872(.dina(n944),.dinb(w_dff_B_7ogxw4qH9_1),.dout(n945),.clk(gclk));
	jand g0873(.dina(n945),.dinb(w_dff_B_WcwNvsPZ5_1),.dout(n946),.clk(gclk));
	jnot g0874(.din(w_n946_0[2]),.dout(G390),.clk(gclk));
	jand g0875(.dina(w_n738_0[0]),.dinb(w_n734_0[0]),.dout(n948),.clk(gclk));
	jand g0876(.dina(w_n703_0[0]),.dinb(w_n559_0[1]),.dout(n949),.clk(gclk));
	jxor g0877(.dina(w_n949_0[2]),.dinb(w_n721_0[2]),.dout(n950),.clk(gclk));
	jxor g0878(.dina(n950),.dinb(w_n718_0[1]),.dout(n951),.clk(gclk));
	jand g0879(.dina(n951),.dinb(w_n948_0[2]),.dout(n952),.clk(gclk));
	jnot g0880(.din(w_n952_0[1]),.dout(n953),.clk(gclk));
	jand g0881(.dina(w_n949_0[1]),.dinb(w_n727_0[1]),.dout(n954),.clk(gclk));
	jcb g0882(.dina(w_n658_0[0]),.dinb(w_n415_0[1]),.dout(n955));
	jcb g0883(.dina(w_dff_B_b2BqNUgk9_0),.dinb(w_n546_0[1]),.dout(n956));
	jcb g0884(.dina(w_n717_0[0]),.dinb(w_n409_0[0]),.dout(n957));
	jand g0885(.dina(n957),.dinb(w_n715_0[0]),.dout(n958),.clk(gclk));
	jand g0886(.dina(n958),.dinb(n956),.dout(n959),.clk(gclk));
	jxor g0887(.dina(n959),.dinb(w_n726_0[0]),.dout(n960),.clk(gclk));
	jxor g0888(.dina(w_dff_B_vZGGj2Qm5_0),.dinb(n954),.dout(n961),.clk(gclk));
	jnot g0889(.din(w_n961_0[2]),.dout(n962),.clk(gclk));
	jcb g0890(.dina(n962),.dinb(w_n564_0[2]),.dout(n963));
	jcb g0891(.dina(w_dff_B_LciRUnhA4_0),.dinb(n953),.dout(n964));
	jcb g0892(.dina(w_n952_0[0]),.dinb(w_n564_0[1]),.dout(n965));
	jand g0893(.dina(w_n965_0[1]),.dinb(w_n573_0[2]),.dout(n966),.clk(gclk));
	jcb g0894(.dina(w_n966_0[1]),.dinb(w_n961_0[1]),.dout(n967));
	jand g0895(.dina(w_n714_0[0]),.dinb(w_n578_1[1]),.dout(n968),.clk(gclk));
	jnot g0896(.din(n968),.dout(n969),.clk(gclk));
	jand g0897(.dina(w_n584_2[0]),.dinb(w_G50_2[2]),.dout(n970),.clk(gclk));
	jand g0898(.dina(w_n598_4[0]),.dinb(w_G132_1[0]),.dout(n971),.clk(gclk));
	jand g0899(.dina(w_n603_4[0]),.dinb(w_G125_0[1]),.dout(n972),.clk(gclk));
	jcb g0900(.dina(n972),.dinb(n971),.dout(n973));
	jcb g0901(.dina(n973),.dinb(n970),.dout(n974));
	jand g0902(.dina(w_n588_4[0]),.dinb(w_G128_0[2]),.dout(n975),.clk(gclk));
	jand g0903(.dina(w_n592_4[0]),.dinb(w_G137_1[0]),.dout(n976),.clk(gclk));
	jand g0904(.dina(w_n607_2[1]),.dinb(w_G159_1[2]),.dout(n977),.clk(gclk));
	jcb g0905(.dina(n977),.dinb(n976),.dout(n978));
	jcb g0906(.dina(n978),.dinb(n975),.dout(n979));
	jand g0907(.dina(w_n609_4[0]),.dinb(w_G143_1[1]),.dout(n980),.clk(gclk));
	jand g0908(.dina(w_n594_3[0]),.dinb(w_G150_1[2]),.dout(n981),.clk(gclk));
	jcb g0909(.dina(n981),.dinb(n980),.dout(n982));
	jcb g0910(.dina(n982),.dinb(w_G33_4[1]),.dout(n983));
	jcb g0911(.dina(n983),.dinb(n979),.dout(n984));
	jcb g0912(.dina(n984),.dinb(n974),.dout(n985));
	jand g0913(.dina(w_n588_3[2]),.dinb(w_G283_1[2]),.dout(n986),.clk(gclk));
	jand g0914(.dina(w_n609_3[2]),.dinb(w_G97_2[1]),.dout(n987),.clk(gclk));
	jcb g0915(.dina(n987),.dinb(n986),.dout(n988));
	jand g0916(.dina(w_n598_3[2]),.dinb(w_G116_2[1]),.dout(n989),.clk(gclk));
	jcb g0917(.dina(n989),.dinb(w_n913_0[0]),.dout(n990));
	jcb g0918(.dina(n990),.dinb(n988),.dout(n991));
	jcb g0919(.dina(w_n687_0[0]),.dinb(w_n595_0[0]),.dout(n992));
	jand g0920(.dina(w_n592_3[2]),.dinb(w_G107_1[2]),.dout(n993),.clk(gclk));
	jand g0921(.dina(w_n603_3[2]),.dinb(w_G294_1[1]),.dout(n994),.clk(gclk));
	jcb g0922(.dina(n994),.dinb(n993),.dout(n995));
	jcb g0923(.dina(n995),.dinb(n992),.dout(n996));
	jcb g0924(.dina(n996),.dinb(n991),.dout(n997));
	jcb g0925(.dina(n997),.dinb(w_n153_3[1]),.dout(n998));
	jand g0926(.dina(n998),.dinb(n985),.dout(n999),.clk(gclk));
	jcb g0927(.dina(n999),.dinb(w_n634_2[0]),.dout(n1000));
	jand g0928(.dina(w_n662_1[0]),.dinb(w_n108_0[1]),.dout(n1001),.clk(gclk));
	jnot g0929(.din(n1001),.dout(n1002),.clk(gclk));
	jand g0930(.dina(n1002),.dinb(w_dff_B_bvJN8E9G5_1),.dout(n1003),.clk(gclk));
	jand g0931(.dina(n1003),.dinb(w_n574_2[0]),.dout(n1004),.clk(gclk));
	jand g0932(.dina(w_dff_B_HvPTZidA6_0),.dinb(n969),.dout(n1005),.clk(gclk));
	jnot g0933(.din(n1005),.dout(n1006),.clk(gclk));
	jand g0934(.dina(w_dff_B_s905FG0E6_0),.dinb(n967),.dout(n1007),.clk(gclk));
	jand g0935(.dina(n1007),.dinb(w_dff_B_XckPm41r1_1),.dout(n1008),.clk(gclk));
	jnot g0936(.din(w_n1008_0[2]),.dout(G378),.clk(gclk));
	jxor g0937(.dina(w_n949_0[0]),.dinb(w_n727_0[0]),.dout(n1010),.clk(gclk));
	jxor g0938(.dina(n1010),.dinb(w_n718_0[0]),.dout(n1011),.clk(gclk));
	jcb g0939(.dina(w_n961_0[0]),.dinb(w_n1011_0[1]),.dout(n1012));
	jand g0940(.dina(n1012),.dinb(w_n948_0[1]),.dout(n1013),.clk(gclk));
	jand g0941(.dina(n1013),.dinb(w_n573_0[1]),.dout(n1014),.clk(gclk));
	jcb g0942(.dina(n1014),.dinb(w_n574_1[2]),.dout(n1015));
	jnot g0943(.din(w_n440_0[0]),.dout(n1016),.clk(gclk));
	jand g0944(.dina(w_n530_0[1]),.dinb(n1016),.dout(n1017),.clk(gclk));
	jxor g0945(.dina(n1017),.dinb(w_n449_0[0]),.dout(n1018),.clk(gclk));
	jxor g0946(.dina(w_n1018_0[1]),.dinb(w_n725_0[0]),.dout(n1019),.clk(gclk));
	jxor g0947(.dina(n1019),.dinb(w_n731_0[0]),.dout(n1020),.clk(gclk));
	jcb g0948(.dina(w_dff_B_2JA7K7KZ0_0),.dinb(n1015),.dout(n1021));
	jand g0949(.dina(w_n1018_0[0]),.dinb(w_n578_1[0]),.dout(n1022),.clk(gclk));
	jnot g0950(.din(n1022),.dout(n1023),.clk(gclk));
	jand g0951(.dina(w_n662_0[2]),.dinb(w_n99_0[1]),.dout(n1024),.clk(gclk));
	jnot g0952(.din(n1024),.dout(n1025),.clk(gclk));
	jand g0953(.dina(w_G50_2[1]),.dinb(w_G41_0[0]),.dout(n1026),.clk(gclk));
	jand g0954(.dina(w_n598_3[1]),.dinb(w_G107_1[1]),.dout(n1027),.clk(gclk));
	jand g0955(.dina(w_n584_1[2]),.dinb(w_G58_2[0]),.dout(n1028),.clk(gclk));
	jcb g0956(.dina(w_n1028_0[1]),.dinb(n1027),.dout(n1029));
	jand g0957(.dina(w_n609_3[1]),.dinb(w_G87_1[1]),.dout(n1030),.clk(gclk));
	jand g0958(.dina(w_n603_3[1]),.dinb(w_G283_1[1]),.dout(n1031),.clk(gclk));
	jcb g0959(.dina(n1031),.dinb(w_n153_3[0]),.dout(n1032));
	jcb g0960(.dina(n1032),.dinb(n1030),.dout(n1033));
	jcb g0961(.dina(w_n866_0[0]),.dinb(w_n778_0[0]),.dout(n1034));
	jand g0962(.dina(w_n588_3[1]),.dinb(w_G116_2[0]),.dout(n1035),.clk(gclk));
	jand g0963(.dina(w_n592_3[1]),.dinb(w_G97_2[0]),.dout(n1036),.clk(gclk));
	jcb g0964(.dina(n1036),.dinb(n1035),.dout(n1037));
	jcb g0965(.dina(n1037),.dinb(n1034),.dout(n1038));
	jcb g0966(.dina(n1038),.dinb(n1033),.dout(n1039));
	jcb g0967(.dina(n1039),.dinb(n1029),.dout(n1040));
	jand g0968(.dina(w_n594_2[2]),.dinb(w_G143_1[0]),.dout(n1041),.clk(gclk));
	jand g0969(.dina(w_n609_3[0]),.dinb(w_G137_0[2]),.dout(n1042),.clk(gclk));
	jcb g0970(.dina(n1042),.dinb(w_G33_4[0]),.dout(n1043));
	jcb g0971(.dina(n1043),.dinb(n1041),.dout(n1044));
	jand g0972(.dina(w_n598_3[0]),.dinb(w_G128_0[1]),.dout(n1045),.clk(gclk));
	jand g0973(.dina(w_n584_1[1]),.dinb(w_G159_1[1]),.dout(n1046),.clk(gclk));
	jcb g0974(.dina(n1046),.dinb(n1045),.dout(n1047));
	jand g0975(.dina(w_n592_3[0]),.dinb(w_G132_0[2]),.dout(n1048),.clk(gclk));
	jand g0976(.dina(w_n588_3[0]),.dinb(w_G125_0[0]),.dout(n1049),.clk(gclk));
	jcb g0977(.dina(n1049),.dinb(n1048),.dout(n1050));
	jand g0978(.dina(w_n603_3[0]),.dinb(w_dff_B_cWQFdEAc9_1),.dout(n1051),.clk(gclk));
	jand g0979(.dina(w_n607_2[0]),.dinb(w_G150_1[1]),.dout(n1052),.clk(gclk));
	jcb g0980(.dina(n1052),.dinb(n1051),.dout(n1053));
	jcb g0981(.dina(n1053),.dinb(n1050),.dout(n1054));
	jcb g0982(.dina(n1054),.dinb(n1047),.dout(n1055));
	jcb g0983(.dina(n1055),.dinb(n1044),.dout(n1056));
	jand g0984(.dina(n1056),.dinb(n1040),.dout(n1057),.clk(gclk));
	jand g0985(.dina(n1057),.dinb(w_n169_0[1]),.dout(n1058),.clk(gclk));
	jcb g0986(.dina(n1058),.dinb(w_n634_1[2]),.dout(n1059));
	jcb g0987(.dina(n1059),.dinb(w_dff_B_Oqeoyf9n3_1),.dout(n1060));
	jand g0988(.dina(n1060),.dinb(n1025),.dout(n1061),.clk(gclk));
	jand g0989(.dina(w_dff_B_nKk6nYl89_0),.dinb(n1023),.dout(n1062),.clk(gclk));
	jand g0990(.dina(n1062),.dinb(w_n574_1[1]),.dout(n1063),.clk(gclk));
	jnot g0991(.din(n1063),.dout(n1064),.clk(gclk));
	jand g0992(.dina(w_dff_B_RK1iR2RE8_0),.dinb(n1021),.dout(n1065),.clk(gclk));
	jnot g0993(.din(w_n1065_0[2]),.dout(G375),.clk(gclk));
	jnot g0994(.din(w_n965_0[0]),.dout(n1067),.clk(gclk));
	jand g0995(.dina(n1067),.dinb(w_n948_0[0]),.dout(n1068),.clk(gclk));
	jnot g0996(.din(n1068),.dout(n1069),.clk(gclk));
	jcb g0997(.dina(w_n966_0[0]),.dinb(w_n1011_0[0]),.dout(n1070));
	jand g0998(.dina(w_n721_0[1]),.dinb(w_n578_0[2]),.dout(n1071),.clk(gclk));
	jnot g0999(.din(n1071),.dout(n1072),.clk(gclk));
	jand g1000(.dina(w_n607_1[2]),.dinb(w_G50_2[0]),.dout(n1073),.clk(gclk));
	jcb g1001(.dina(n1073),.dinb(w_n1028_0[0]),.dout(n1074));
	jand g1002(.dina(w_n592_2[2]),.dinb(w_G143_0[2]),.dout(n1075),.clk(gclk));
	jand g1003(.dina(w_n609_2[2]),.dinb(w_G150_1[0]),.dout(n1076),.clk(gclk));
	jcb g1004(.dina(n1076),.dinb(n1075),.dout(n1077));
	jcb g1005(.dina(n1077),.dinb(w_G33_3[2]),.dout(n1078));
	jcb g1006(.dina(n1078),.dinb(n1074),.dout(n1079));
	jand g1007(.dina(w_n594_2[1]),.dinb(w_G159_1[0]),.dout(n1080),.clk(gclk));
	jand g1008(.dina(w_n588_2[2]),.dinb(w_G132_0[1]),.dout(n1081),.clk(gclk));
	jand g1009(.dina(w_n598_2[2]),.dinb(w_G137_0[1]),.dout(n1082),.clk(gclk));
	jand g1010(.dina(w_n603_2[2]),.dinb(w_G128_0[0]),.dout(n1083),.clk(gclk));
	jcb g1011(.dina(n1083),.dinb(n1082),.dout(n1084));
	jcb g1012(.dina(n1084),.dinb(n1081),.dout(n1085));
	jcb g1013(.dina(n1085),.dinb(n1080),.dout(n1086));
	jcb g1014(.dina(n1086),.dinb(n1079),.dout(n1087));
	jand g1015(.dina(w_n588_2[1]),.dinb(w_G294_1[0]),.dout(n1088),.clk(gclk));
	jand g1016(.dina(w_n609_2[1]),.dinb(w_G107_1[0]),.dout(n1089),.clk(gclk));
	jand g1017(.dina(w_n603_2[1]),.dinb(w_G303_0[2]),.dout(n1090),.clk(gclk));
	jcb g1018(.dina(n1090),.dinb(w_n153_2[2]),.dout(n1091));
	jcb g1019(.dina(n1091),.dinb(n1089),.dout(n1092));
	jand g1020(.dina(w_n594_2[0]),.dinb(w_G97_1[2]),.dout(n1093),.clk(gclk));
	jand g1021(.dina(w_n592_2[1]),.dinb(w_G116_1[2]),.dout(n1094),.clk(gclk));
	jcb g1022(.dina(n1094),.dinb(n1093),.dout(n1095));
	jand g1023(.dina(w_n598_2[1]),.dinb(w_G283_1[0]),.dout(n1096),.clk(gclk));
	jcb g1024(.dina(n1096),.dinb(w_n780_0[0]),.dout(n1097));
	jcb g1025(.dina(n1097),.dinb(n1095),.dout(n1098));
	jcb g1026(.dina(n1098),.dinb(n1092),.dout(n1099));
	jcb g1027(.dina(n1099),.dinb(n1088),.dout(n1100));
	jcb g1028(.dina(n1100),.dinb(w_n859_0[0]),.dout(n1101));
	jand g1029(.dina(n1101),.dinb(n1087),.dout(n1102),.clk(gclk));
	jcb g1030(.dina(n1102),.dinb(w_n634_1[1]),.dout(n1103));
	jand g1031(.dina(w_n662_0[1]),.dinb(w_n103_0[1]),.dout(n1104),.clk(gclk));
	jcb g1032(.dina(w_dff_B_fq1EQPkL3_0),.dinb(w_n575_0[0]),.dout(n1105));
	jnot g1033(.din(n1105),.dout(n1106),.clk(gclk));
	jand g1034(.dina(n1106),.dinb(w_dff_B_mjwmoLdh9_1),.dout(n1107),.clk(gclk));
	jand g1035(.dina(w_dff_B_L7D1CmnO6_0),.dinb(n1072),.dout(n1108),.clk(gclk));
	jnot g1036(.din(n1108),.dout(n1109),.clk(gclk));
	jand g1037(.dina(w_dff_B_vrgbrAzy6_0),.dinb(n1070),.dout(n1110),.clk(gclk));
	jand g1038(.dina(w_dff_B_58Zn26et7_0),.dinb(n1069),.dout(n1111),.clk(gclk));
	jnot g1039(.din(w_n1111_0[2]),.dout(G381),.clk(gclk));
	jand g1040(.dina(w_n1065_0[1]),.dinb(w_n1008_0[1]),.dout(n1113),.clk(gclk));
	jnot g1041(.din(w_G384_0),.dout(n1114),.clk(gclk));
	jand g1042(.dina(w_n1111_0[1]),.dinb(w_n1114_0[1]),.dout(n1115),.clk(gclk));
	jand g1043(.dina(w_n946_0[1]),.dinb(w_n832_0[1]),.dout(n1116),.clk(gclk));
	jnot g1044(.din(w_G396_0[1]),.dout(n1117),.clk(gclk));
	jand g1045(.dina(w_n897_0[1]),.dinb(w_dff_B_ABBEEnfy1_1),.dout(n1118),.clk(gclk));
	jand g1046(.dina(w_dff_B_A1EWhcBU9_0),.dinb(n1116),.dout(n1119),.clk(gclk));
	jand g1047(.dina(n1119),.dinb(w_dff_B_tIvGYJEx6_1),.dout(n1120),.clk(gclk));
	jand g1048(.dina(n1120),.dinb(w_n1113_0[1]),.dout(n1121),.clk(gclk));
	jnot g1049(.din(w_n1121_0[1]),.dout(G407),.clk(gclk));
	jnot g1050(.din(w_G213_0[0]),.dout(n1123),.clk(gclk));
	jcb g1051(.dina(w_G343_0[0]),.dinb(w_n1123_0[1]),.dout(n1124));
	jnot g1052(.din(w_n1124_0[1]),.dout(n1125),.clk(gclk));
	jand g1053(.dina(w_n1125_0[1]),.dinb(w_n1113_0[0]),.dout(n1126),.clk(gclk));
	jcb g1054(.dina(n1126),.dinb(w_n1123_0[0]),.dout(n1127));
	jcb g1055(.dina(w_dff_B_ADgAvYvc2_0),.dinb(w_n1121_0[0]),.dout(G409));
	jxor g1056(.dina(w_n897_0[0]),.dinb(w_G396_0[0]),.dout(n1129),.clk(gclk));
	jxor g1057(.dina(w_n946_0[0]),.dinb(w_n832_0[0]),.dout(n1130),.clk(gclk));
	jxor g1058(.dina(n1130),.dinb(w_dff_B_BAtwaBZ78_1),.dout(n1131),.clk(gclk));
	jxor g1059(.dina(w_n1111_0[0]),.dinb(w_n1114_0[0]),.dout(n1132),.clk(gclk));
	jxor g1060(.dina(w_dff_B_RbEAYj8h2_0),.dinb(n1131),.dout(n1133),.clk(gclk));
	jxor g1061(.dina(w_n1065_0[0]),.dinb(w_n1008_0[0]),.dout(n1134),.clk(gclk));
	jcb g1062(.dina(w_n1134_0[1]),.dinb(w_n1125_0[0]),.dout(n1135));
	jcb g1063(.dina(w_n1124_0[0]),.dinb(w_dff_B_OqV6vmQM6_1),.dout(n1136));
	jand g1064(.dina(w_dff_B_F7opRmds6_0),.dinb(n1135),.dout(n1137),.clk(gclk));
	jxor g1065(.dina(w_dff_B_CzT4pdQb5_0),.dinb(w_n1133_0[1]),.dout(G405),.clk(gclk));
	jxor g1066(.dina(w_n1134_0[0]),.dinb(w_n1133_0[0]),.dout(G402),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_dff_A_bfz3X9zz6_2),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_dff_A_V2sEVFqm3_0),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_dff_A_VEUEFbh67_1),.din(w_G1_0[1]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_G13_0[1]),.doutc(w_G13_0[2]),.din(G13));
	jspl3 jspl3_w_G13_1(.douta(w_dff_A_QxIYbuhb7_0),.doutb(w_dff_A_QvlrAJJ99_1),.doutc(w_G13_1[2]),.din(w_G13_0[0]));
	jspl jspl_w_G13_2(.douta(w_dff_A_LPh7b7Kr5_0),.doutb(w_G13_2[1]),.din(w_G13_0[1]));
	jspl3 jspl3_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.doutc(w_G20_0[2]),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_dff_A_PneygkG64_0),.doutb(w_dff_A_RsTLAMxA9_1),.doutc(w_G20_1[2]),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_dff_A_B75geTHS5_1),.doutc(w_G20_2[2]),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_G20_3[1]),.doutc(w_dff_A_BHi2T2dg0_2),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_G20_4[0]),.doutb(w_dff_A_Ivahdf7R9_1),.doutc(w_G20_4[2]),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_dff_A_bERrxIDg1_0),.doutb(w_dff_A_iXH7P5d46_1),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_G20_6[0]),.doutb(w_G20_6[1]),.doutc(w_dff_A_xBj5cX0X9_2),.din(w_G20_1[2]));
	jspl jspl_w_G20_7(.douta(w_G20_7[0]),.doutb(w_dff_A_d7G0uZeB0_1),.din(w_G20_2[0]));
	jspl3 jspl3_w_G33_0(.douta(w_dff_A_1AiiHIgY1_0),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_dff_A_hsbDY3rh5_0),.doutb(w_dff_A_Earr44st9_1),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_dff_A_OTVES8wK6_1),.doutc(w_dff_A_L7ZuTVMZ3_2),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_G33_4[0]),.doutb(w_G33_4[1]),.doutc(w_G33_4[2]),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_G33_5[0]),.doutb(w_G33_5[1]),.doutc(w_G33_5[2]),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_dff_A_1wDiKAeu7_0),.doutb(w_dff_A_czSiPcGG6_1),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_G33_7[0]),.doutb(w_G33_7[1]),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_G33_8[0]),.doutb(w_G33_8[1]),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_dff_A_w31GkA329_0),.doutb(w_G33_9[1]),.doutc(w_G33_9[2]),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_G33_10[0]),.doutb(w_G33_10[1]),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl jspl_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_G41_0[1]),.doutc(w_G41_0[2]),.din(G41));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_dff_A_kC2B1HrP3_1),.doutc(w_G45_0[2]),.din(G45));
	jspl jspl_w_G45_1(.douta(w_G45_1[0]),.doutb(w_dff_A_s8fqRlFn4_1),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_G50_0[1]),.doutc(w_dff_A_XteHk1YD6_2),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_G50_1[0]),.doutb(w_G50_1[1]),.doutc(w_G50_1[2]),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_dff_A_zBJPXltE3_0),.doutb(w_G50_2[1]),.doutc(w_dff_A_c0hMX5Af4_2),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_G50_3[0]),.doutb(w_G50_3[1]),.doutc(w_G50_3[2]),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_G50_4[0]),.doutb(w_dff_A_OKTHj1IG9_1),.doutc(w_dff_A_7IDlMxKm4_2),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_dff_A_b9GROpJW2_0),.doutb(w_dff_A_G2slVSIU2_1),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G50_6(.douta(w_G50_6[0]),.doutb(w_G50_6[1]),.doutc(w_G50_6[2]),.din(w_G50_1[2]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_dff_A_k3uNQ6l93_1),.doutc(w_G58_0[2]),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_dff_A_T0huWdzQ2_0),.doutb(w_G58_1[1]),.doutc(w_G58_1[2]),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_dff_A_M2LnEw7Y9_0),.doutb(w_dff_A_zFPCULDU7_1),.doutc(w_G58_2[2]),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_dff_A_3vO6REX67_0),.doutb(w_dff_A_VhN3Y8XQ5_1),.doutc(w_G58_3[2]),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_dff_A_iNETUz0D5_0),.doutb(w_dff_A_NqtSGlXd4_1),.doutc(w_G58_4[2]),.din(w_G58_1[0]));
	jspl3 jspl3_w_G58_5(.douta(w_G58_5[0]),.doutb(w_dff_A_HRH4bXPe7_1),.doutc(w_dff_A_gLmHOx7C6_2),.din(w_G58_1[1]));
	jspl3 jspl3_w_G58_6(.douta(w_G58_6[0]),.doutb(w_G58_6[1]),.doutc(w_G58_6[2]),.din(w_G58_1[2]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_dff_A_XB9u5wBA3_2),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_G68_1[0]),.doutb(w_G68_1[1]),.doutc(w_dff_A_NtRs0Lns7_2),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_dff_A_NipjuKUi1_1),.doutc(w_dff_A_AlWz1lJ56_2),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_dff_A_fMQD3J5V6_1),.doutc(w_dff_A_c26WNJs30_2),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_dff_A_3qsiCGA71_0),.doutb(w_G68_4[1]),.doutc(w_dff_A_GoKqyPRw1_2),.din(w_G68_1[0]));
	jspl3 jspl3_w_G68_5(.douta(w_G68_5[0]),.doutb(w_G68_5[1]),.doutc(w_G68_5[2]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_dff_A_5hCaIDoL6_1),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_G77_1[0]),.doutb(w_dff_A_nLvSUpGX2_1),.doutc(w_G77_1[2]),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_dff_A_6rWT0e2E1_0),.doutb(w_dff_A_3PFdd2zu2_1),.doutc(w_G77_2[2]),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_dff_A_9xqjFTvx0_0),.doutb(w_G77_3[1]),.doutc(w_dff_A_iUBzaUNc4_2),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_dff_A_ZNWPlGT61_0),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl3 jspl3_w_G87_0(.douta(w_G87_0[0]),.doutb(w_dff_A_Cb6U7dYo9_1),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_dff_A_YZd3ftvQ7_1),.doutc(w_dff_A_vEhoGedL2_2),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_dff_A_Y8g8JBsj4_0),.doutb(w_G87_2[1]),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_G87_3[0]),.doutb(w_dff_A_K5fo6cxL0_1),.doutc(w_dff_A_aAnbTL744_2),.din(w_G87_0[2]));
	jspl jspl_w_G87_4(.douta(w_G87_4[0]),.doutb(w_G87_4[1]),.din(w_G87_1[0]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_dff_A_HDfvmbSy5_1),.doutc(w_G97_0[2]),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_G97_1[1]),.doutc(w_dff_A_Xa25Z2Up3_2),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_G97_2[1]),.doutc(w_dff_A_EBAejq0L1_2),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_dff_A_FhAe9Zg75_0),.doutb(w_dff_A_fXEdsmQ75_1),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_dff_A_0DUZvNbg9_0),.doutb(w_G97_4[1]),.doutc(w_dff_A_XTGG9y8x7_2),.din(w_G97_1[0]));
	jspl jspl_w_G97_5(.douta(w_G97_5[0]),.doutb(w_G97_5[1]),.din(w_G97_1[1]));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_CwrNi5cu0_0),.doutb(w_dff_A_AeYLXE9H6_1),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_G107_1[1]),.doutc(w_G107_1[2]),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_G107_2[1]),.doutc(w_G107_2[2]),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_G107_3[0]),.doutb(w_G107_3[1]),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_dff_A_Nsl13udB4_1),.doutc(w_dff_A_399Kevc33_2),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_G116_1[1]),.doutc(w_dff_A_7r9CT32r7_2),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_G116_2[1]),.doutc(w_G116_2[2]),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_G116_3[0]),.doutb(w_G116_3[1]),.doutc(w_G116_3[2]),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_dff_A_FEZpIib27_0),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl jspl_w_G116_5(.douta(w_dff_A_AYHq6CK15_0),.doutb(w_G116_5[1]),.din(w_G116_1[1]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_G125_0[1]),.din(w_dff_B_3ciWDK0f1_2));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(w_dff_B_LoEDOQo05_3));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(w_dff_B_RxdeFCrb9_3));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_G132_1[1]),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(w_dff_B_zrwlyaUU3_3));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_G137_1[1]),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(w_dff_B_DnzrD0rl8_3));
	jspl3 jspl3_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.doutc(w_G143_1[2]),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_dff_A_guwEpJeY9_0),.doutb(w_dff_A_nvKubPcz8_1),.doutc(w_G150_0[2]),.din(w_dff_B_KH0k5irM5_3));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_G150_1[1]),.doutc(w_G150_1[2]),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_G150_2[1]),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_dff_A_fDXdL3SA3_0),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_dff_A_uCZnG92N2_0),.doutb(w_dff_A_ynTVZFdy6_1),.doutc(w_G159_0[2]),.din(w_dff_B_6tq39FvZ8_3));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_G159_1[2]),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_dff_A_tikgggIb4_0),.doutb(w_dff_A_69Qogbok1_1),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_dff_A_cKU9WJCE0_0),.doutb(w_G169_0[1]),.doutc(w_dff_A_OacZVhaD0_2),.din(G169));
	jspl3 jspl3_w_G169_1(.douta(w_G169_1[0]),.doutb(w_G169_1[1]),.doutc(w_G169_1[2]),.din(w_G169_0[0]));
	jspl jspl_w_G169_2(.douta(w_dff_A_jIv7nspd0_0),.doutb(w_G169_2[1]),.din(w_G169_0[1]));
	jspl3 jspl3_w_G179_0(.douta(w_G179_0[0]),.doutb(w_G179_0[1]),.doutc(w_dff_A_1pMPP5rW9_2),.din(G179));
	jspl jspl_w_G179_1(.douta(w_dff_A_hPZj13FQ6_0),.doutb(w_G179_1[1]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G190_0(.douta(w_G190_0[0]),.doutb(w_dff_A_zFoFmfc91_1),.doutc(w_dff_A_pvLVCwaM3_2),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_G190_1[0]),.doutb(w_dff_A_9znQbK8K4_1),.doutc(w_dff_A_VnHop4lI8_2),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_G190_2[0]),.doutb(w_dff_A_YC9e3UYf0_1),.doutc(w_dff_A_wyqwC8n39_2),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_G190_3[0]),.doutb(w_dff_A_0ZhmkXJ00_1),.doutc(w_dff_A_kYJkszQe9_2),.din(w_G190_0[2]));
	jspl3 jspl3_w_G190_4(.douta(w_G190_4[0]),.doutb(w_dff_A_hRzyRzXw2_1),.doutc(w_dff_A_a5fQVTzg2_2),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_dff_A_8rPchjsM9_2),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_G200_1[0]),.doutb(w_dff_A_RsJcQgEB6_1),.doutc(w_dff_A_Eme40qrN6_2),.din(w_G200_0[0]));
	jspl jspl_w_G200_2(.douta(w_G200_2[0]),.doutb(w_dff_A_AdX3ri1D4_1),.din(w_G200_0[1]));
	jspl jspl_w_G213_0(.douta(w_G213_0[0]),.doutb(w_dff_A_0tYGGUoq8_1),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(w_dff_B_HboFerw58_2));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_dff_A_Pw3VdEjM4_1),.doutc(w_dff_A_bgcYkwPV5_2),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_dff_A_MFW7rTmx9_0),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_dff_A_XQmfFHEB3_1),.doutc(w_dff_A_bXd2SWAe9_2),.din(G232));
	jspl jspl_w_G232_1(.douta(w_G232_1[0]),.doutb(w_G232_1[1]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_G238_0[0]),.doutb(w_dff_A_B6Vs1lec3_1),.doutc(w_dff_A_zd486uqH3_2),.din(G238));
	jspl jspl_w_G238_1(.douta(w_dff_A_ER2hJ8O59_0),.doutb(w_G238_1[1]),.din(w_G238_0[0]));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_dff_A_5F61E4JD0_1),.doutc(w_dff_A_agEXFetD7_2),.din(G244));
	jspl jspl_w_G244_1(.douta(w_dff_A_xdO5RVy33_0),.doutb(w_G244_1[1]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_G250_0[0]),.doutb(w_dff_A_EnmipDdM3_1),.doutc(w_dff_A_NYiak4bQ0_2),.din(G250));
	jspl3 jspl3_w_G250_1(.douta(w_dff_A_4itEZmO81_0),.doutb(w_G250_1[1]),.doutc(w_G250_1[2]),.din(w_G250_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_dff_A_g5fnT28m4_1),.doutc(w_dff_A_1ZCCUhkB4_2),.din(G257));
	jspl jspl_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.din(w_G257_0[0]));
	jspl jspl_w_G264_0(.douta(w_dff_A_c1JWmLH73_0),.doutb(w_G264_0[1]),.din(G264));
	jspl jspl_w_G270_0(.douta(w_dff_A_L1LfM2zG9_0),.doutb(w_G270_0[1]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_dff_A_UOhAl3AG6_0),.doutb(w_dff_A_hXLqg86h2_1),.doutc(w_G274_0[2]),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_dff_A_Z4gpDrdV4_0),.doutb(w_dff_A_6Nv8glqm8_1),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_G283_1[1]),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_G283_2[0]),.doutb(w_G283_2[1]),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_dff_A_OgmqfJ9Y9_0),.doutb(w_dff_A_japh8m6f2_1),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_dff_A_g8b3qWfZ8_0),.doutb(w_dff_A_qeqK6uzc8_1),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_G294_1[1]),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_G294_2[0]),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_dff_A_QktPgrCA7_0),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_dff_A_u9ZGdr624_0),.doutb(w_G303_0[1]),.doutc(w_dff_A_gHd0RMZ40_2),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_dff_A_zIemMhgn9_0),.doutb(w_dff_A_WRB8si7u2_1),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(w_dff_B_kZ0fZPgi3_3));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_G311_1[1]),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(w_dff_B_pIQiSaGZ0_3));
	jspl jspl_w_G317_1(.douta(w_G317_1[0]),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_G322_0[0]),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(w_dff_B_Pa74sO4r2_3));
	jspl jspl_w_G326_0(.douta(w_G326_0[0]),.doutb(w_G326_0[1]),.din(w_dff_B_C9KSGfsQ0_2));
	jspl3 jspl3_w_G330_0(.douta(w_G330_0[0]),.doutb(w_dff_A_yhCoLZdL9_1),.doutc(w_G330_0[2]),.din(w_dff_B_hWTaQiHW1_3));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_dff_A_paEEYKD64_1),.din(w_dff_B_t80UjEDy7_2));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_dff_A_iBXhMxwh8_2),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_dff_A_Yp6EBFDp7_0),.doutb(G355),.din(w_dff_B_JxW6VFUK4_2));
	jspl3 jspl3_w_G396_0(.douta(w_dff_A_L227eugT4_0),.doutb(w_G396_0[1]),.doutc(w_dff_A_8YmVFp8d9_2),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_G384_0),.doutb(w_dff_A_UxchZKH33_1),.din(G384_fa_));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_dff_A_XCor1GRt1_1),.doutc(w_dff_A_n1rNZ6VJ4_2),.din(n73));
	jspl jspl_w_n73_1(.douta(w_n73_1[0]),.doutb(w_n73_1[1]),.din(w_n73_0[0]));
	jspl jspl_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.din(n74));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl3 jspl3_w_n78_0(.douta(w_n78_0[0]),.doutb(w_dff_A_sucufshR2_1),.doutc(w_n78_0[2]),.din(n78));
	jspl jspl_w_n78_1(.douta(w_n78_1[0]),.doutb(w_dff_A_DUwZdRKu2_1),.din(w_n78_0[0]));
	jspl3 jspl3_w_n79_0(.douta(w_n79_0[0]),.doutb(w_dff_A_KOPMjFeF6_1),.doutc(w_n79_0[2]),.din(n79));
	jspl jspl_w_n79_1(.douta(w_n79_1[0]),.doutb(w_n79_1[1]),.din(w_n79_0[0]));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.doutc(w_dff_A_iMa7f0N08_2),.din(n80));
	jspl3 jspl3_w_n80_1(.douta(w_dff_A_yLyYwaU37_0),.doutb(w_n80_1[1]),.doutc(w_dff_A_54pfsnNL9_2),.din(w_n80_0[0]));
	jspl3 jspl3_w_n80_2(.douta(w_n80_2[0]),.doutb(w_n80_2[1]),.doutc(w_n80_2[2]),.din(w_n80_0[1]));
	jspl3 jspl3_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.doutc(w_dff_A_Xkk2p6Kp8_2),.din(n83));
	jspl3 jspl3_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.doutc(w_n84_0[2]),.din(n84));
	jspl jspl_w_n84_1(.douta(w_n84_1[0]),.doutb(w_n84_1[1]),.din(w_n84_0[0]));
	jspl3 jspl3_w_n85_0(.douta(w_n85_0[0]),.doutb(w_dff_A_3raSrlKE7_1),.doutc(w_n85_0[2]),.din(n85));
	jspl jspl_w_n85_1(.douta(w_n85_1[0]),.doutb(w_n85_1[1]),.din(w_n85_0[0]));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n89_0(.douta(w_n89_0[0]),.doutb(w_n89_0[1]),.doutc(w_n89_0[2]),.din(n89));
	jspl3 jspl3_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n90_1(.douta(w_n90_1[0]),.doutb(w_n90_1[1]),.doutc(w_n90_1[2]),.din(w_n90_0[0]));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_dff_A_Q6r6O0Ff9_1),.doutc(w_n92_0[2]),.din(n92));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl jspl_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.din(n95));
	jspl3 jspl3_w_n99_0(.douta(w_n99_0[0]),.doutb(w_dff_A_LPCp8wUi4_1),.doutc(w_n99_0[2]),.din(n99));
	jspl3 jspl3_w_n99_1(.douta(w_dff_A_zZbqqVKJ0_0),.doutb(w_dff_A_3z5vq90N2_1),.doutc(w_n99_1[2]),.din(w_n99_0[0]));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_p26f3lRV2_1),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n103_1(.douta(w_dff_A_FwUPWvLI2_0),.doutb(w_n103_1[1]),.doutc(w_n103_1[2]),.din(w_n103_0[0]));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl3 jspl3_w_n107_0(.douta(w_dff_A_4DbpvSP54_0),.doutb(w_n107_0[1]),.doutc(w_n107_0[2]),.din(n107));
	jspl3 jspl3_w_n108_0(.douta(w_n108_0[0]),.doutb(w_dff_A_73UYEdBJ2_1),.doutc(w_n108_0[2]),.din(n108));
	jspl jspl_w_n108_1(.douta(w_dff_A_Z4bHatZS4_0),.doutb(w_n108_1[1]),.din(w_n108_0[0]));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_dff_A_P28HTxyQ2_1),.doutc(w_dff_A_iOyGJcSv8_2),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_dff_A_J6dLmODg2_0),.doutb(w_dff_A_wQiY8xZZ6_1),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl jspl_w_n113_0(.douta(w_dff_A_7GZeRR1V0_0),.doutb(w_n113_0[1]),.din(n113));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n127_0(.douta(w_dff_A_XIOaokYB8_0),.doutb(w_n127_0[1]),.din(n127));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_dff_A_DaGiIoEz7_1),.din(n131));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_dff_A_q76h1Grp0_1),.din(n135));
	jspl jspl_w_n138_0(.douta(w_dff_A_s2WD0Y0I5_0),.doutb(w_n138_0[1]),.din(n138));
	jspl3 jspl3_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.doutc(w_n140_0[2]),.din(n140));
	jspl3 jspl3_w_n140_1(.douta(w_n140_1[0]),.doutb(w_dff_A_R7XW4HVH1_1),.doutc(w_dff_A_MlDAFvhn9_2),.din(w_n140_0[0]));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl3 jspl3_w_n142_0(.douta(w_dff_A_L8RaPNdA8_0),.doutb(w_n142_0[1]),.doutc(w_n142_0[2]),.din(n142));
	jspl3 jspl3_w_n142_1(.douta(w_n142_1[0]),.doutb(w_n142_1[1]),.doutc(w_n142_1[2]),.din(w_n142_0[0]));
	jspl3 jspl3_w_n142_2(.douta(w_n142_2[0]),.doutb(w_n142_2[1]),.doutc(w_dff_A_zOeZyDd71_2),.din(w_n142_0[1]));
	jspl3 jspl3_w_n142_3(.douta(w_n142_3[0]),.doutb(w_n142_3[1]),.doutc(w_n142_3[2]),.din(w_n142_0[2]));
	jspl jspl_w_n142_4(.douta(w_n142_4[0]),.doutb(w_n142_4[1]),.din(w_n142_1[0]));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl3 jspl3_w_n143_1(.douta(w_dff_A_3ismzyuC2_0),.doutb(w_n143_1[1]),.doutc(w_n143_1[2]),.din(w_n143_0[0]));
	jspl jspl_w_n143_2(.douta(w_n143_2[0]),.doutb(w_n143_2[1]),.din(w_n143_0[1]));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(n144));
	jspl3 jspl3_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.doutc(w_n145_0[2]),.din(n145));
	jspl3 jspl3_w_n145_1(.douta(w_n145_1[0]),.doutb(w_n145_1[1]),.doutc(w_n145_1[2]),.din(w_n145_0[0]));
	jspl jspl_w_n145_2(.douta(w_n145_2[0]),.doutb(w_n145_2[1]),.din(w_n145_0[1]));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_dff_A_kOWn8T0U2_0),.doutb(w_dff_A_Y7vdIFIK6_1),.doutc(w_n151_1[2]),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_dff_A_AdIubfXa6_0),.doutb(w_n151_3[1]),.doutc(w_dff_A_OO7uJMLQ3_2),.din(w_n151_0[2]));
	jspl jspl_w_n151_4(.douta(w_dff_A_Ytt10nUx2_0),.doutb(w_n151_4[1]),.din(w_n151_1[0]));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_dff_A_DytGePDb4_1),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_dff_A_An85pV1v5_2),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_dff_A_la4Lg7iy3_0),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_dff_A_skgac2vk4_2),.din(w_n153_0[1]));
	jspl3 jspl3_w_n153_3(.douta(w_n153_3[0]),.doutb(w_n153_3[1]),.doutc(w_n153_3[2]),.din(w_n153_0[2]));
	jspl3 jspl3_w_n153_4(.douta(w_n153_4[0]),.doutb(w_n153_4[1]),.doutc(w_n153_4[2]),.din(w_n153_1[0]));
	jspl3 jspl3_w_n153_5(.douta(w_dff_A_9qTpjvg52_0),.doutb(w_dff_A_8PiacHDd5_1),.doutc(w_n153_5[2]),.din(w_n153_1[1]));
	jspl3 jspl3_w_n153_6(.douta(w_n153_6[0]),.doutb(w_n153_6[1]),.doutc(w_n153_6[2]),.din(w_n153_1[2]));
	jspl3 jspl3_w_n153_7(.douta(w_n153_7[0]),.doutb(w_n153_7[1]),.doutc(w_n153_7[2]),.din(w_n153_2[0]));
	jspl3 jspl3_w_n153_8(.douta(w_n153_8[0]),.doutb(w_n153_8[1]),.doutc(w_n153_8[2]),.din(w_n153_2[1]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_dff_A_s1ptZKpM2_1),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_dff_A_kIGrJzaO2_1),.doutc(w_dff_A_01IyBm3r8_2),.din(w_dff_B_988m3ij01_3));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_dff_A_Wjps8uhV2_1),.din(w_n163_0[0]));
	jspl jspl_w_n165_0(.douta(w_dff_A_9J1j9XG43_0),.doutb(w_n165_0[1]),.din(n165));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl3 jspl3_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.doutc(w_n167_1[2]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n167_2(.douta(w_n167_2[0]),.doutb(w_dff_A_7yVOR6bZ8_1),.doutc(w_dff_A_Z4RwFHax0_2),.din(w_n167_0[1]));
	jspl3 jspl3_w_n167_3(.douta(w_n167_3[0]),.doutb(w_n167_3[1]),.doutc(w_dff_A_hSILwcqq7_2),.din(w_n167_0[2]));
	jspl jspl_w_n167_4(.douta(w_n167_4[0]),.doutb(w_n167_4[1]),.din(w_n167_1[0]));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_dff_A_JElLs7Gx3_1),.din(n168));
	jspl3 jspl3_w_n169_0(.douta(w_n169_0[0]),.doutb(w_dff_A_Jqsgc3Ot4_1),.doutc(w_dff_A_WqVsXXA43_2),.din(n169));
	jspl jspl_w_n169_1(.douta(w_n169_1[0]),.doutb(w_dff_A_ByMvWYW64_1),.din(w_n169_0[0]));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl3 jspl3_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.doutc(w_n171_0[2]),.din(n171));
	jspl jspl_w_n171_1(.douta(w_n171_1[0]),.doutb(w_n171_1[1]),.din(w_n171_0[0]));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n173_0(.douta(w_dff_A_Aj3lUnKW1_0),.doutb(w_n173_0[1]),.doutc(w_dff_A_kQnQgSOO9_2),.din(n173));
	jspl3 jspl3_w_n175_0(.douta(w_n175_0[0]),.doutb(w_dff_A_vatFgBln0_1),.doutc(w_n175_0[2]),.din(n175));
	jspl3 jspl3_w_n175_1(.douta(w_n175_1[0]),.doutb(w_dff_A_s5KBHbYF5_1),.doutc(w_dff_A_Vt7nZ2km2_2),.din(w_n175_0[0]));
	jspl3 jspl3_w_n175_2(.douta(w_dff_A_J8Xrpnru1_0),.doutb(w_n175_2[1]),.doutc(w_dff_A_MfTlVsaB8_2),.din(w_n175_0[1]));
	jspl jspl_w_n175_3(.douta(w_n175_3[0]),.doutb(w_dff_A_B5Q1wpPz9_1),.din(w_n175_0[2]));
	jspl3 jspl3_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.doutc(w_n176_0[2]),.din(n176));
	jspl3 jspl3_w_n176_1(.douta(w_n176_1[0]),.doutb(w_n176_1[1]),.doutc(w_n176_1[2]),.din(w_n176_0[0]));
	jspl3 jspl3_w_n176_2(.douta(w_n176_2[0]),.doutb(w_n176_2[1]),.doutc(w_n176_2[2]),.din(w_n176_0[1]));
	jspl jspl_w_n176_3(.douta(w_n176_3[0]),.doutb(w_n176_3[1]),.din(w_n176_0[2]));
	jspl jspl_w_n177_0(.douta(w_dff_A_Jh9CEhWh9_0),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(w_dff_B_DAC8bilL0_3));
	jspl jspl_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.din(w_n181_0[0]));
	jspl jspl_w_n183_0(.douta(w_n183_0[0]),.doutb(w_dff_A_fOVcn0cu7_1),.din(n183));
	jspl jspl_w_n187_0(.douta(w_n187_0[0]),.doutb(w_dff_A_KO3ZZ86d4_1),.din(n187));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_dff_A_KpbIBopu1_1),.doutc(w_dff_A_DSBvx0Ah3_2),.din(n191));
	jspl3 jspl3_w_n191_1(.douta(w_n191_1[0]),.doutb(w_dff_A_CLNDS7V07_1),.doutc(w_dff_A_BxkjGqqB8_2),.din(w_n191_0[0]));
	jspl3 jspl3_w_n191_2(.douta(w_n191_2[0]),.doutb(w_n191_2[1]),.doutc(w_dff_A_27yDXbBi6_2),.din(w_n191_0[1]));
	jspl3 jspl3_w_n191_3(.douta(w_dff_A_zyKZmBA41_0),.doutb(w_dff_A_v5J5apna9_1),.doutc(w_n191_3[2]),.din(w_n191_0[2]));
	jspl3 jspl3_w_n193_0(.douta(w_dff_A_fj4txxlY0_0),.doutb(w_n193_0[1]),.doutc(w_dff_A_czs1bfAp0_2),.din(n193));
	jspl3 jspl3_w_n199_0(.douta(w_dff_A_0ywe8Y0j3_0),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_dff_A_fvx1FcJL2_1),.din(n200));
	jspl3 jspl3_w_n202_0(.douta(w_n202_0[0]),.doutb(w_dff_A_qvasqyZf6_1),.doutc(w_n202_0[2]),.din(n202));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_dff_A_3eBytgpX4_1),.din(n204));
	jspl jspl_w_n208_0(.douta(w_n208_0[0]),.doutb(w_dff_A_QKpOV3Co8_1),.din(n208));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_dff_A_GzGL9BU06_1),.din(n210));
	jspl jspl_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.din(n211));
	jspl jspl_w_n214_0(.douta(w_dff_A_Mguwjh3Y5_0),.doutb(w_n214_0[1]),.din(n214));
	jspl3 jspl3_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.doutc(w_n221_0[2]),.din(n221));
	jspl jspl_w_n221_1(.douta(w_n221_1[0]),.doutb(w_n221_1[1]),.din(w_n221_0[0]));
	jspl jspl_w_n223_0(.douta(w_dff_A_x836GCzJ0_0),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(n225));
	jspl jspl_w_n228_0(.douta(w_dff_A_SPflITre2_0),.doutb(w_n228_0[1]),.din(w_dff_B_IluYWD2B6_2));
	jspl jspl_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.din(n233));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.din(n234));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_n237_0[1]),.doutc(w_n237_0[2]),.din(n237));
	jspl3 jspl3_w_n237_1(.douta(w_n237_1[0]),.doutb(w_n237_1[1]),.doutc(w_n237_1[2]),.din(w_n237_0[0]));
	jspl jspl_w_n243_0(.douta(w_dff_A_5cPOZy7q5_0),.doutb(w_n243_0[1]),.din(n243));
	jspl3 jspl3_w_n246_0(.douta(w_dff_A_2kHRESU46_0),.doutb(w_n246_0[1]),.doutc(w_dff_A_GsXmotwF4_2),.din(n246));
	jspl3 jspl3_w_n251_0(.douta(w_dff_A_0WdZJnEe2_0),.doutb(w_dff_A_ZOM03yNy5_1),.doutc(w_n251_0[2]),.din(n251));
	jspl3 jspl3_w_n251_1(.douta(w_dff_A_Lvok6WBq7_0),.doutb(w_n251_1[1]),.doutc(w_n251_1[2]),.din(w_n251_0[0]));
	jspl3 jspl3_w_n251_2(.douta(w_n251_2[0]),.doutb(w_dff_A_WgCxRYDW1_1),.doutc(w_dff_A_vUBv06Fc3_2),.din(w_n251_0[1]));
	jspl3 jspl3_w_n255_0(.douta(w_n255_0[0]),.doutb(w_dff_A_jEkaSazK0_1),.doutc(w_n255_0[2]),.din(n255));
	jspl jspl_w_n255_1(.douta(w_n255_1[0]),.doutb(w_n255_1[1]),.din(w_n255_0[0]));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n267_1(.douta(w_n267_1[0]),.doutb(w_n267_1[1]),.doutc(w_n267_1[2]),.din(w_n267_0[0]));
	jspl jspl_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.din(n268));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(n269));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n275_0(.douta(w_dff_A_ak5WnuVE9_0),.doutb(w_n275_0[1]),.din(w_dff_B_ak8NJgpB3_2));
	jspl3 jspl3_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.doutc(w_dff_A_Jb85nn0H4_2),.din(n283));
	jspl jspl_w_n283_1(.douta(w_n283_1[0]),.doutb(w_n283_1[1]),.din(w_n283_0[0]));
	jspl3 jspl3_w_n284_0(.douta(w_dff_A_0sn6RaSv1_0),.doutb(w_dff_A_XlLw9ZLW4_1),.doutc(w_n284_0[2]),.din(n284));
	jspl3 jspl3_w_n284_1(.douta(w_n284_1[0]),.doutb(w_n284_1[1]),.doutc(w_dff_A_1TN1V6Zt4_2),.din(w_n284_0[0]));
	jspl jspl_w_n285_0(.douta(w_dff_A_4ZkRuOox8_0),.doutb(w_n285_0[1]),.din(n285));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(n289));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(n290));
	jspl jspl_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.din(n291));
	jspl jspl_w_n292_0(.douta(w_n292_0[0]),.doutb(w_dff_A_h3ncExe39_1),.din(n292));
	jspl jspl_w_n294_0(.douta(w_dff_A_GXpsoGnT9_0),.doutb(w_n294_0[1]),.din(n294));
	jspl jspl_w_n295_0(.douta(w_dff_A_8ak2UWrj6_0),.doutb(w_n295_0[1]),.din(w_dff_B_irG8Eo2N2_2));
	jspl jspl_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.din(n297));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_dff_A_SLgBHqgl5_1),.din(n298));
	jspl jspl_w_n301_0(.douta(w_dff_A_Rc1cOJEn9_0),.doutb(w_n301_0[1]),.din(n301));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.doutc(w_n306_0[2]),.din(n306));
	jspl jspl_w_n306_1(.douta(w_n306_1[0]),.doutb(w_n306_1[1]),.din(w_n306_0[0]));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_dff_A_1NcBMjnV7_1),.din(n307));
	jspl jspl_w_n309_0(.douta(w_dff_A_qI8LMykU9_0),.doutb(w_n309_0[1]),.din(n309));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_dff_A_mBQNp16G1_1),.din(n312));
	jspl3 jspl3_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.doutc(w_dff_A_VYQW2B8n1_2),.din(n320));
	jspl jspl_w_n320_1(.douta(w_dff_A_GgI2SKKZ4_0),.doutb(w_n320_1[1]),.din(w_n320_0[0]));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_efSbgbCQ2_1),.din(w_dff_B_Fvc9IbLX9_2));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl jspl_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.din(w_n327_0[0]));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n331_0(.douta(w_n331_0[0]),.doutb(w_n331_0[1]),.din(n331));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n335_0(.douta(w_dff_A_sOt7iCiN6_0),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl3 jspl3_w_n339_0(.douta(w_n339_0[0]),.doutb(w_dff_A_9mcLTUWd1_1),.doutc(w_n339_0[2]),.din(n339));
	jspl jspl_w_n339_1(.douta(w_dff_A_O14BRBRi1_0),.doutb(w_n339_1[1]),.din(w_n339_0[0]));
	jspl jspl_w_n341_0(.douta(w_n341_0[0]),.doutb(w_dff_A_SaZw2CP78_1),.din(n341));
	jspl jspl_w_n342_0(.douta(w_n342_0[0]),.doutb(w_dff_A_4kvJkFvK4_1),.din(n342));
	jspl3 jspl3_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.doutc(w_n350_0[2]),.din(n350));
	jspl jspl_w_n350_1(.douta(w_n350_1[0]),.doutb(w_n350_1[1]),.din(w_n350_0[0]));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(n354));
	jspl jspl_w_n354_1(.douta(w_n354_1[0]),.doutb(w_n354_1[1]),.din(w_n354_0[0]));
	jspl jspl_w_n357_0(.douta(w_dff_A_kXI2QyuQ6_0),.doutb(w_n357_0[1]),.din(w_dff_B_90XzA1Er2_2));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_dff_A_41I9nSRK2_1),.din(w_dff_B_klgUUWDg7_2));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl3 jspl3_w_n381_0(.douta(w_dff_A_DoPik7nl2_0),.doutb(w_n381_0[1]),.doutc(w_n381_0[2]),.din(n381));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl jspl_w_n391_1(.douta(w_n391_1[0]),.doutb(w_n391_1[1]),.din(w_n391_0[0]));
	jspl jspl_w_n394_0(.douta(w_dff_A_W091tQYi5_0),.doutb(w_n394_0[1]),.din(w_dff_B_b5ePqyXQ6_2));
	jspl3 jspl3_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.doutc(w_n403_0[2]),.din(n403));
	jspl3 jspl3_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.doutc(w_n406_0[2]),.din(n406));
	jspl jspl_w_n409_0(.douta(w_dff_A_L5ZUWAUW0_0),.doutb(w_n409_0[1]),.din(n409));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl3 jspl3_w_n415_0(.douta(w_dff_A_UXK1BWGK5_0),.doutb(w_dff_A_akqUpS582_1),.doutc(w_n415_0[2]),.din(n415));
	jspl jspl_w_n415_1(.douta(w_n415_1[0]),.doutb(w_n415_1[1]),.din(w_n415_0[0]));
	jspl3 jspl3_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.doutc(w_n424_0[2]),.din(n424));
	jspl jspl_w_n424_1(.douta(w_n424_1[0]),.doutb(w_n424_1[1]),.din(w_n424_0[0]));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(n427));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl3 jspl3_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.doutc(w_n440_0[2]),.din(n440));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl jspl_w_n449_0(.douta(w_n449_0[0]),.doutb(w_dff_A_yDkvygq41_1),.din(n449));
	jspl3 jspl3_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.doutc(w_n458_0[2]),.din(n458));
	jspl jspl_w_n458_1(.douta(w_n458_1[0]),.doutb(w_n458_1[1]),.din(w_n458_0[0]));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl3 jspl3_w_n476_0(.douta(w_n476_0[0]),.doutb(w_dff_A_Hfd7It0H9_1),.doutc(w_dff_A_B46Hbzmp1_2),.din(n476));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n484_0(.douta(w_dff_A_vQK9rPe47_0),.doutb(w_n484_0[1]),.din(n484));
	jspl jspl_w_n486_0(.douta(w_dff_A_FNp8w6bp1_0),.doutb(w_n486_0[1]),.din(n486));
	jspl3 jspl3_w_n487_0(.douta(w_dff_A_sS1Clive5_0),.doutb(w_dff_A_F8KG0rd27_1),.doutc(w_n487_0[2]),.din(w_dff_B_AHRCaxL13_3));
	jspl jspl_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.din(n491));
	jspl jspl_w_n497_0(.douta(w_n497_0[0]),.doutb(w_dff_A_6nQF6u7s9_1),.din(n497));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_dff_A_ex4bYEwq2_1),.din(w_dff_B_IOoAVviH4_2));
	jspl jspl_w_n506_0(.douta(w_n506_0[0]),.doutb(w_n506_0[1]),.din(n506));
	jspl jspl_w_n510_0(.douta(w_n510_0[0]),.doutb(w_dff_A_kzR7u1TD1_1),.din(n510));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n525_0(.douta(w_dff_A_vH9QyFAH4_0),.doutb(w_n525_0[1]),.din(n525));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_dff_A_f9fPes1r4_1),.doutc(w_dff_A_emKsr4Fg6_2),.din(n530));
	jspl jspl_w_n530_1(.douta(w_dff_A_9S3vw8Ew3_0),.doutb(w_n530_1[1]),.din(w_n530_0[0]));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_dff_A_lSEecwiY4_1),.doutc(w_dff_A_4gOG3Ltk0_2),.din(n531));
	jspl3 jspl3_w_n531_1(.douta(w_n531_1[0]),.doutb(w_dff_A_bDA0GVVs0_1),.doutc(w_dff_A_9E02IJP68_2),.din(w_n531_0[0]));
	jspl3 jspl3_w_n531_2(.douta(w_dff_A_AFBer5jh7_0),.doutb(w_n531_2[1]),.doutc(w_dff_A_tBWwSSqg8_2),.din(w_n531_0[1]));
	jspl3 jspl3_w_n531_3(.douta(w_n531_3[0]),.doutb(w_dff_A_WWbyJ8n71_1),.doutc(w_dff_A_0o0f1lf62_2),.din(w_n531_0[2]));
	jspl3 jspl3_w_n531_4(.douta(w_n531_4[0]),.doutb(w_n531_4[1]),.doutc(w_dff_A_2jLXFuQv9_2),.din(w_n531_1[0]));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl3 jspl3_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.doutc(w_dff_A_dK2rfGwR3_2),.din(n538));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl3 jspl3_w_n541_0(.douta(w_dff_A_sqJjZZ9z9_0),.doutb(w_n541_0[1]),.doutc(w_dff_A_f28f5INd7_2),.din(w_dff_B_mQ5ZAuB85_3));
	jspl3 jspl3_w_n541_1(.douta(w_n541_1[0]),.doutb(w_n541_1[1]),.doutc(w_dff_A_u1iOwQ3o1_2),.din(w_n541_0[0]));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_t1HLMZXK2_2));
	jspl3 jspl3_w_n544_0(.douta(w_dff_A_OKKURVhr0_0),.doutb(w_n544_0[1]),.doutc(w_n544_0[2]),.din(n544));
	jspl3 jspl3_w_n546_0(.douta(w_n546_0[0]),.doutb(w_n546_0[1]),.doutc(w_n546_0[2]),.din(n546));
	jspl jspl_w_n546_1(.douta(w_n546_1[0]),.doutb(w_dff_A_nKpt3kIN3_1),.din(w_n546_0[0]));
	jspl3 jspl3_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.doutc(w_n559_0[2]),.din(n559));
	jspl3 jspl3_w_n559_1(.douta(w_n559_1[0]),.doutb(w_n559_1[1]),.doutc(w_n559_1[2]),.din(w_n559_0[0]));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.din(w_n561_0[0]));
	jspl3 jspl3_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_oX0tGj6o2_1),.doutc(w_dff_A_JmiBRX3w8_2),.din(n564));
	jspl3 jspl3_w_n564_1(.douta(w_dff_A_yZfjNgZR7_0),.doutb(w_n564_1[1]),.doutc(w_n564_1[2]),.din(w_n564_0[0]));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_dff_A_6P2bOYnB9_1),.doutc(w_dff_A_oF0G75GT9_2),.din(w_dff_B_TbB8LnBB0_3));
	jspl3 jspl3_w_n573_1(.douta(w_dff_A_UdbYpxOn5_0),.doutb(w_dff_A_suiCb5en8_1),.doutc(w_n573_1[2]),.din(w_n573_0[0]));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_dff_A_rntIr00f0_2),.din(n574));
	jspl3 jspl3_w_n574_1(.douta(w_n574_1[0]),.doutb(w_dff_A_EI3WYb5P3_1),.doutc(w_dff_A_1AnaTcwN1_2),.din(w_n574_0[0]));
	jspl3 jspl3_w_n574_2(.douta(w_dff_A_kcHBLyaI9_0),.doutb(w_n574_2[1]),.doutc(w_dff_A_kdVNOwJ95_2),.din(w_n574_0[1]));
	jspl3 jspl3_w_n574_3(.douta(w_dff_A_Mb1QoJJ16_0),.doutb(w_dff_A_nQyxS2Ra9_1),.doutc(w_n574_3[2]),.din(w_n574_0[2]));
	jspl jspl_w_n574_4(.douta(w_dff_A_kMWFvHvv5_0),.doutb(w_n574_4[1]),.din(w_n574_1[0]));
	jspl3 jspl3_w_n575_0(.douta(w_n575_0[0]),.doutb(w_dff_A_LK58E5yq2_1),.doutc(w_dff_A_4bcMFsIz0_2),.din(n575));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_dff_A_DbuiHhS49_2),.din(n578));
	jspl3 jspl3_w_n578_1(.douta(w_dff_A_ptrud9cU5_0),.doutb(w_dff_A_afHsN3HE2_1),.doutc(w_n578_1[2]),.din(w_n578_0[0]));
	jspl jspl_w_n578_2(.douta(w_dff_A_FK04W79i4_0),.doutb(w_n578_2[1]),.din(w_n578_0[1]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_dff_A_Tc0cGRKe8_1),.doutc(w_dff_A_3VbCZcko9_2),.din(n579));
	jspl3 jspl3_w_n579_1(.douta(w_dff_A_YQ8M2Mcf1_0),.doutb(w_n579_1[1]),.doutc(w_dff_A_Sf5n20R13_2),.din(w_n579_0[0]));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(n583));
	jspl3 jspl3_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.doutc(w_n584_0[2]),.din(n584));
	jspl3 jspl3_w_n584_1(.douta(w_n584_1[0]),.doutb(w_n584_1[1]),.doutc(w_n584_1[2]),.din(w_n584_0[0]));
	jspl3 jspl3_w_n584_2(.douta(w_n584_2[0]),.doutb(w_n584_2[1]),.doutc(w_n584_2[2]),.din(w_n584_0[1]));
	jspl3 jspl3_w_n584_3(.douta(w_n584_3[0]),.doutb(w_n584_3[1]),.doutc(w_n584_3[2]),.din(w_n584_0[2]));
	jspl jspl_w_n584_4(.douta(w_n584_4[0]),.doutb(w_n584_4[1]),.din(w_n584_1[0]));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.din(n587));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl3 jspl3_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.doutc(w_n588_1[2]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n588_2(.douta(w_n588_2[0]),.doutb(w_n588_2[1]),.doutc(w_n588_2[2]),.din(w_n588_0[1]));
	jspl3 jspl3_w_n588_3(.douta(w_n588_3[0]),.doutb(w_n588_3[1]),.doutc(w_n588_3[2]),.din(w_n588_0[2]));
	jspl3 jspl3_w_n588_4(.douta(w_n588_4[0]),.doutb(w_n588_4[1]),.doutc(w_n588_4[2]),.din(w_n588_1[0]));
	jspl3 jspl3_w_n588_5(.douta(w_n588_5[0]),.doutb(w_n588_5[1]),.doutc(w_n588_5[2]),.din(w_n588_1[1]));
	jspl3 jspl3_w_n588_6(.douta(w_n588_6[0]),.doutb(w_n588_6[1]),.doutc(w_n588_6[2]),.din(w_n588_1[2]));
	jspl jspl_w_n588_7(.douta(w_n588_7[0]),.doutb(w_n588_7[1]),.din(w_n588_2[0]));
	jspl3 jspl3_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.doutc(w_n592_0[2]),.din(n592));
	jspl3 jspl3_w_n592_1(.douta(w_n592_1[0]),.doutb(w_n592_1[1]),.doutc(w_n592_1[2]),.din(w_n592_0[0]));
	jspl3 jspl3_w_n592_2(.douta(w_n592_2[0]),.doutb(w_n592_2[1]),.doutc(w_n592_2[2]),.din(w_n592_0[1]));
	jspl3 jspl3_w_n592_3(.douta(w_n592_3[0]),.doutb(w_n592_3[1]),.doutc(w_n592_3[2]),.din(w_n592_0[2]));
	jspl3 jspl3_w_n592_4(.douta(w_n592_4[0]),.doutb(w_n592_4[1]),.doutc(w_n592_4[2]),.din(w_n592_1[0]));
	jspl3 jspl3_w_n592_5(.douta(w_n592_5[0]),.doutb(w_n592_5[1]),.doutc(w_n592_5[2]),.din(w_n592_1[1]));
	jspl3 jspl3_w_n592_6(.douta(w_n592_6[0]),.doutb(w_n592_6[1]),.doutc(w_n592_6[2]),.din(w_n592_1[2]));
	jspl jspl_w_n592_7(.douta(w_n592_7[0]),.doutb(w_n592_7[1]),.din(w_n592_2[0]));
	jspl3 jspl3_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.doutc(w_n594_0[2]),.din(n594));
	jspl3 jspl3_w_n594_1(.douta(w_n594_1[0]),.doutb(w_n594_1[1]),.doutc(w_n594_1[2]),.din(w_n594_0[0]));
	jspl3 jspl3_w_n594_2(.douta(w_n594_2[0]),.doutb(w_n594_2[1]),.doutc(w_n594_2[2]),.din(w_n594_0[1]));
	jspl3 jspl3_w_n594_3(.douta(w_n594_3[0]),.doutb(w_n594_3[1]),.doutc(w_n594_3[2]),.din(w_n594_0[2]));
	jspl3 jspl3_w_n594_4(.douta(w_n594_4[0]),.doutb(w_n594_4[1]),.doutc(w_n594_4[2]),.din(w_n594_1[0]));
	jspl3 jspl3_w_n594_5(.douta(w_n594_5[0]),.doutb(w_n594_5[1]),.doutc(w_n594_5[2]),.din(w_n594_1[1]));
	jspl jspl_w_n594_6(.douta(w_n594_6[0]),.doutb(w_n594_6[1]),.din(w_n594_1[2]));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl3 jspl3_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.doutc(w_n598_0[2]),.din(n598));
	jspl3 jspl3_w_n598_1(.douta(w_n598_1[0]),.doutb(w_n598_1[1]),.doutc(w_n598_1[2]),.din(w_n598_0[0]));
	jspl3 jspl3_w_n598_2(.douta(w_n598_2[0]),.doutb(w_n598_2[1]),.doutc(w_n598_2[2]),.din(w_n598_0[1]));
	jspl3 jspl3_w_n598_3(.douta(w_n598_3[0]),.doutb(w_n598_3[1]),.doutc(w_n598_3[2]),.din(w_n598_0[2]));
	jspl3 jspl3_w_n598_4(.douta(w_n598_4[0]),.doutb(w_n598_4[1]),.doutc(w_n598_4[2]),.din(w_n598_1[0]));
	jspl3 jspl3_w_n598_5(.douta(w_n598_5[0]),.doutb(w_n598_5[1]),.doutc(w_n598_5[2]),.din(w_n598_1[1]));
	jspl3 jspl3_w_n598_6(.douta(w_n598_6[0]),.doutb(w_n598_6[1]),.doutc(w_n598_6[2]),.din(w_n598_1[2]));
	jspl jspl_w_n598_7(.douta(w_n598_7[0]),.doutb(w_n598_7[1]),.din(w_n598_2[0]));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl jspl_w_n601_0(.douta(w_dff_A_iKTNXKZc3_0),.doutb(w_n601_0[1]),.din(n601));
	jspl3 jspl3_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.doutc(w_n603_0[2]),.din(n603));
	jspl3 jspl3_w_n603_1(.douta(w_n603_1[0]),.doutb(w_n603_1[1]),.doutc(w_n603_1[2]),.din(w_n603_0[0]));
	jspl3 jspl3_w_n603_2(.douta(w_n603_2[0]),.doutb(w_n603_2[1]),.doutc(w_n603_2[2]),.din(w_n603_0[1]));
	jspl3 jspl3_w_n603_3(.douta(w_n603_3[0]),.doutb(w_n603_3[1]),.doutc(w_n603_3[2]),.din(w_n603_0[2]));
	jspl3 jspl3_w_n603_4(.douta(w_n603_4[0]),.doutb(w_n603_4[1]),.doutc(w_n603_4[2]),.din(w_n603_1[0]));
	jspl3 jspl3_w_n603_5(.douta(w_n603_5[0]),.doutb(w_n603_5[1]),.doutc(w_n603_5[2]),.din(w_n603_1[1]));
	jspl3 jspl3_w_n603_6(.douta(w_n603_6[0]),.doutb(w_n603_6[1]),.doutc(w_n603_6[2]),.din(w_n603_1[2]));
	jspl jspl_w_n603_7(.douta(w_n603_7[0]),.doutb(w_n603_7[1]),.din(w_n603_2[0]));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl3 jspl3_w_n607_1(.douta(w_n607_1[0]),.doutb(w_n607_1[1]),.doutc(w_n607_1[2]),.din(w_n607_0[0]));
	jspl3 jspl3_w_n607_2(.douta(w_n607_2[0]),.doutb(w_n607_2[1]),.doutc(w_n607_2[2]),.din(w_n607_0[1]));
	jspl3 jspl3_w_n607_3(.douta(w_n607_3[0]),.doutb(w_n607_3[1]),.doutc(w_n607_3[2]),.din(w_n607_0[2]));
	jspl3 jspl3_w_n607_4(.douta(w_n607_4[0]),.doutb(w_n607_4[1]),.doutc(w_n607_4[2]),.din(w_n607_1[0]));
	jspl jspl_w_n607_5(.douta(w_n607_5[0]),.doutb(w_n607_5[1]),.din(w_n607_1[1]));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n609_1(.douta(w_n609_1[0]),.doutb(w_n609_1[1]),.doutc(w_n609_1[2]),.din(w_n609_0[0]));
	jspl3 jspl3_w_n609_2(.douta(w_n609_2[0]),.doutb(w_n609_2[1]),.doutc(w_n609_2[2]),.din(w_n609_0[1]));
	jspl3 jspl3_w_n609_3(.douta(w_n609_3[0]),.doutb(w_n609_3[1]),.doutc(w_n609_3[2]),.din(w_n609_0[2]));
	jspl3 jspl3_w_n609_4(.douta(w_n609_4[0]),.doutb(w_n609_4[1]),.doutc(w_n609_4[2]),.din(w_n609_1[0]));
	jspl3 jspl3_w_n609_5(.douta(w_n609_5[0]),.doutb(w_n609_5[1]),.doutc(w_n609_5[2]),.din(w_n609_1[1]));
	jspl3 jspl3_w_n609_6(.douta(w_n609_6[0]),.doutb(w_n609_6[1]),.doutc(w_n609_6[2]),.din(w_n609_1[2]));
	jspl jspl_w_n609_7(.douta(w_n609_7[0]),.doutb(w_n609_7[1]),.din(w_n609_2[0]));
	jspl3 jspl3_w_n634_0(.douta(w_dff_A_NpB3G7Bq5_0),.doutb(w_dff_A_nZFqLcox7_1),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n634_1(.douta(w_n634_1[0]),.doutb(w_dff_A_qC7rVrwi6_1),.doutc(w_dff_A_HH7vxqTT1_2),.din(w_n634_0[0]));
	jspl3 jspl3_w_n634_2(.douta(w_n634_2[0]),.doutb(w_n634_2[1]),.doutc(w_n634_2[2]),.din(w_n634_0[1]));
	jspl3 jspl3_w_n634_3(.douta(w_dff_A_nSuweLyS0_0),.doutb(w_dff_A_Ih9jq9Sa3_1),.doutc(w_n634_3[2]),.din(w_n634_0[2]));
	jspl jspl_w_n634_4(.douta(w_n634_4[0]),.doutb(w_dff_A_mwQXrT2J4_1),.din(w_n634_1[0]));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_dff_A_x3cqZVrK0_1),.din(n637));
	jspl3 jspl3_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.doutc(w_n639_0[2]),.din(n639));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl jspl_w_n645_1(.douta(w_n645_1[0]),.doutb(w_n645_1[1]),.din(w_n645_0[0]));
	jspl jspl_w_n647_0(.douta(w_dff_A_9DOAq5WU0_0),.doutb(w_n647_0[1]),.din(n647));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(n658));
	jspl3 jspl3_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.doutc(w_n662_0[2]),.din(n662));
	jspl jspl_w_n662_1(.douta(w_n662_1[0]),.doutb(w_n662_1[1]),.din(w_n662_0[0]));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(n674));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_dff_A_5TScZkiy6_1),.din(n701));
	jspl3 jspl3_w_n703_0(.douta(w_dff_A_Vr0d0vvE7_0),.doutb(w_n703_0[1]),.doutc(w_dff_A_DIwyCqDw2_2),.din(n703));
	jspl3 jspl3_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.doutc(w_dff_A_dOiBy7mD3_2),.din(n714));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_dff_A_ADenmync1_1),.din(w_dff_B_8HkJADyj7_2));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_dff_A_IsgXaCh32_1),.din(n717));
	jspl3 jspl3_w_n718_0(.douta(w_dff_A_Zb2QFsoF3_0),.doutb(w_dff_A_GhUoLhoJ8_1),.doutc(w_n718_0[2]),.din(n718));
	jspl3 jspl3_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.doutc(w_dff_A_MMgmZvqe4_2),.din(n721));
	jspl jspl_w_n721_1(.douta(w_n721_1[0]),.doutb(w_dff_A_gOIn9MML3_1),.din(w_n721_0[0]));
	jspl jspl_w_n725_0(.douta(w_n725_0[0]),.doutb(w_dff_A_Dowq88ls1_1),.din(n725));
	jspl jspl_w_n726_0(.douta(w_dff_A_BrlEhjNb0_0),.doutb(w_n726_0[1]),.din(n726));
	jspl3 jspl3_w_n727_0(.douta(w_dff_A_19aJx0qV7_0),.doutb(w_dff_A_pcYsestV9_1),.doutc(w_n727_0[2]),.din(w_dff_B_3DM4Z68X4_3));
	jspl jspl_w_n729_0(.douta(w_dff_A_Zp6vcKg74_0),.doutb(w_n729_0[1]),.din(w_dff_B_HtTIFEwZ6_2));
	jspl jspl_w_n731_0(.douta(w_n731_0[0]),.doutb(w_n731_0[1]),.din(n731));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n738_0(.douta(w_dff_A_dUpis0yX9_0),.doutb(w_n738_0[1]),.din(n738));
	jspl3 jspl3_w_n755_0(.douta(w_n755_0[0]),.doutb(w_dff_A_5OB9D1s01_1),.doutc(w_n755_0[2]),.din(n755));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_dff_A_prKTJLcj5_1),.din(n760));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(n764));
	jspl jspl_w_n768_0(.douta(w_n768_0[0]),.doutb(w_dff_A_hlWLWior1_1),.din(n768));
	jspl jspl_w_n771_0(.douta(w_dff_A_2ylipEtU7_0),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.din(n801));
	jspl3 jspl3_w_n810_0(.douta(w_n810_0[0]),.doutb(w_dff_A_nZ7gWBPL1_1),.doutc(w_n810_0[2]),.din(n810));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_dff_A_IgTa6ZNf1_1),.din(n819));
	jspl3 jspl3_w_n824_0(.douta(w_dff_A_OppAy5Zf5_0),.doutb(w_dff_A_Y5gNh7m69_1),.doutc(w_n824_0[2]),.din(n824));
	jspl jspl_w_n825_0(.douta(w_dff_A_nyLEkgiy9_0),.doutb(w_n825_0[1]),.din(w_dff_B_RTHaLB9P4_2));
	jspl3 jspl3_w_n827_0(.douta(w_dff_A_f96N0cPC9_0),.doutb(w_dff_A_jdBXqUPm7_1),.doutc(w_n827_0[2]),.din(n827));
	jspl3 jspl3_w_n832_0(.douta(w_dff_A_u1JnJXQ80_0),.doutb(w_dff_A_JciXvHZn2_1),.doutc(w_n832_0[2]),.din(n832));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_dff_A_jnql4Twp1_1),.din(n839));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(n866));
	jspl3 jspl3_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.doutc(w_n897_0[2]),.din(n897));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl3 jspl3_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.doutc(w_n946_0[2]),.din(n946));
	jspl3 jspl3_w_n948_0(.douta(w_dff_A_QKVqJgMz7_0),.doutb(w_n948_0[1]),.doutc(w_n948_0[2]),.din(n948));
	jspl3 jspl3_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.doutc(w_n949_0[2]),.din(n949));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl3 jspl3_w_n961_0(.douta(w_n961_0[0]),.doutb(w_dff_A_v9rMCZ7a8_1),.doutc(w_n961_0[2]),.din(n961));
	jspl jspl_w_n965_0(.douta(w_n965_0[0]),.doutb(w_n965_0[1]),.din(n965));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(n966));
	jspl3 jspl3_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.doutc(w_n1008_0[2]),.din(n1008));
	jspl jspl_w_n1011_0(.douta(w_dff_A_LngoYsIR5_0),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_dff_A_K3YCUiXo4_1),.din(n1018));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(n1028));
	jspl3 jspl3_w_n1065_0(.douta(w_dff_A_w5xjl9lA6_0),.doutb(w_dff_A_0Q6EldbN6_1),.doutc(w_n1065_0[2]),.din(n1065));
	jspl3 jspl3_w_n1111_0(.douta(w_n1111_0[0]),.doutb(w_n1111_0[1]),.doutc(w_n1111_0[2]),.din(n1111));
	jspl jspl_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_dff_A_DbV8GDW21_1),.din(n1113));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(w_dff_B_HLIqN8EU8_2));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(n1121));
	jspl jspl_w_n1123_0(.douta(w_dff_A_WHOdOuRe0_0),.doutb(w_n1123_0[1]),.din(n1123));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.din(w_dff_B_HwM3TxD34_2));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(n1133));
	jspl jspl_w_n1134_0(.douta(w_dff_A_kQQvnavx6_0),.doutb(w_n1134_0[1]),.din(n1134));
	jdff dff_B_r3kRAIpQ2_1(.din(n97),.dout(w_dff_B_r3kRAIpQ2_1),.clk(gclk));
	jdff dff_B_jGjlJCd88_1(.din(n106),.dout(w_dff_B_jGjlJCd88_1),.clk(gclk));
	jdff dff_B_dPcDd7Q30_0(.din(n110),.dout(w_dff_B_dPcDd7Q30_0),.clk(gclk));
	jdff dff_B_bj3H9JTn3_0(.din(n105),.dout(w_dff_B_bj3H9JTn3_0),.clk(gclk));
	jdff dff_B_waQ3RwkB3_0(.din(n96),.dout(w_dff_B_waQ3RwkB3_0),.clk(gclk));
	jdff dff_B_S49LDRpI9_1(.din(n87),.dout(w_dff_B_S49LDRpI9_1),.clk(gclk));
	jdff dff_B_6QtizgNK7_0(.din(n526),.dout(w_dff_B_6QtizgNK7_0),.clk(gclk));
	jdff dff_B_NTDd2y4p9_1(.din(n545),.dout(w_dff_B_NTDd2y4p9_1),.clk(gclk));
	jdff dff_B_YpTj6EKW6_1(.din(w_dff_B_NTDd2y4p9_1),.dout(w_dff_B_YpTj6EKW6_1),.clk(gclk));
	jdff dff_B_pURHap6Y8_1(.din(w_dff_B_YpTj6EKW6_1),.dout(w_dff_B_pURHap6Y8_1),.clk(gclk));
	jdff dff_B_DClWGZvT8_1(.din(w_dff_B_pURHap6Y8_1),.dout(w_dff_B_DClWGZvT8_1),.clk(gclk));
	jdff dff_B_Qmhn8zsG1_1(.din(w_dff_B_DClWGZvT8_1),.dout(w_dff_B_Qmhn8zsG1_1),.clk(gclk));
	jdff dff_B_lUhdfPXP3_1(.din(w_dff_B_Qmhn8zsG1_1),.dout(w_dff_B_lUhdfPXP3_1),.clk(gclk));
	jdff dff_B_iBVGmfQV5_1(.din(w_dff_B_lUhdfPXP3_1),.dout(w_dff_B_iBVGmfQV5_1),.clk(gclk));
	jdff dff_B_qie6ORYr8_1(.din(w_dff_B_iBVGmfQV5_1),.dout(w_dff_B_qie6ORYr8_1),.clk(gclk));
	jdff dff_B_O822c8kH0_1(.din(w_dff_B_qie6ORYr8_1),.dout(w_dff_B_O822c8kH0_1),.clk(gclk));
	jdff dff_B_h8b3xB5Q6_1(.din(w_dff_B_O822c8kH0_1),.dout(w_dff_B_h8b3xB5Q6_1),.clk(gclk));
	jdff dff_B_UrEtn1Rm5_1(.din(w_dff_B_h8b3xB5Q6_1),.dout(w_dff_B_UrEtn1Rm5_1),.clk(gclk));
	jdff dff_B_JycR5cH96_1(.din(w_dff_B_UrEtn1Rm5_1),.dout(w_dff_B_JycR5cH96_1),.clk(gclk));
	jdff dff_B_KZyMGIYv2_1(.din(w_dff_B_JycR5cH96_1),.dout(w_dff_B_KZyMGIYv2_1),.clk(gclk));
	jdff dff_B_3w172eFQ5_1(.din(w_dff_B_KZyMGIYv2_1),.dout(w_dff_B_3w172eFQ5_1),.clk(gclk));
	jdff dff_B_TL65JbtS7_0(.din(n567),.dout(w_dff_B_TL65JbtS7_0),.clk(gclk));
	jdff dff_B_r8qjqQ3n3_0(.din(w_dff_B_TL65JbtS7_0),.dout(w_dff_B_r8qjqQ3n3_0),.clk(gclk));
	jdff dff_B_OS2rrGMa4_0(.din(w_dff_B_r8qjqQ3n3_0),.dout(w_dff_B_OS2rrGMa4_0),.clk(gclk));
	jdff dff_B_CbMaE2zY9_0(.din(w_dff_B_OS2rrGMa4_0),.dout(w_dff_B_CbMaE2zY9_0),.clk(gclk));
	jdff dff_B_ptaXhLjm1_0(.din(w_dff_B_CbMaE2zY9_0),.dout(w_dff_B_ptaXhLjm1_0),.clk(gclk));
	jdff dff_B_jDtbR5Jj2_0(.din(w_dff_B_ptaXhLjm1_0),.dout(w_dff_B_jDtbR5Jj2_0),.clk(gclk));
	jdff dff_B_N1Ub3KP60_0(.din(w_dff_B_jDtbR5Jj2_0),.dout(w_dff_B_N1Ub3KP60_0),.clk(gclk));
	jdff dff_B_cCosgA6U3_0(.din(w_dff_B_N1Ub3KP60_0),.dout(w_dff_B_cCosgA6U3_0),.clk(gclk));
	jdff dff_B_8S1vNq1b8_0(.din(w_dff_B_cCosgA6U3_0),.dout(w_dff_B_8S1vNq1b8_0),.clk(gclk));
	jdff dff_B_s8NVsuFV5_0(.din(w_dff_B_8S1vNq1b8_0),.dout(w_dff_B_s8NVsuFV5_0),.clk(gclk));
	jdff dff_B_PHJb2qWP2_0(.din(w_dff_B_s8NVsuFV5_0),.dout(w_dff_B_PHJb2qWP2_0),.clk(gclk));
	jdff dff_B_Jqbswo0l1_0(.din(w_dff_B_PHJb2qWP2_0),.dout(w_dff_B_Jqbswo0l1_0),.clk(gclk));
	jdff dff_B_8R83VQXs5_0(.din(w_dff_B_Jqbswo0l1_0),.dout(w_dff_B_8R83VQXs5_0),.clk(gclk));
	jdff dff_B_ibgIVVWs3_0(.din(n752),.dout(w_dff_B_ibgIVVWs3_0),.clk(gclk));
	jdff dff_B_LYav221B2_0(.din(w_dff_B_ibgIVVWs3_0),.dout(w_dff_B_LYav221B2_0),.clk(gclk));
	jdff dff_B_BBx7zaFd7_0(.din(w_dff_B_LYav221B2_0),.dout(w_dff_B_BBx7zaFd7_0),.clk(gclk));
	jdff dff_B_ajjuE9LJ1_0(.din(w_dff_B_BBx7zaFd7_0),.dout(w_dff_B_ajjuE9LJ1_0),.clk(gclk));
	jdff dff_B_7Lk5itsx4_0(.din(w_dff_B_ajjuE9LJ1_0),.dout(w_dff_B_7Lk5itsx4_0),.clk(gclk));
	jdff dff_B_YFABmYhq7_0(.din(w_dff_B_7Lk5itsx4_0),.dout(w_dff_B_YFABmYhq7_0),.clk(gclk));
	jdff dff_B_1fHMWvHf6_0(.din(w_dff_B_YFABmYhq7_0),.dout(w_dff_B_1fHMWvHf6_0),.clk(gclk));
	jdff dff_B_ATa868hN3_0(.din(w_dff_B_1fHMWvHf6_0),.dout(w_dff_B_ATa868hN3_0),.clk(gclk));
	jdff dff_B_H9XDiLOP9_0(.din(w_dff_B_ATa868hN3_0),.dout(w_dff_B_H9XDiLOP9_0),.clk(gclk));
	jdff dff_B_UXJUApCm4_0(.din(w_dff_B_H9XDiLOP9_0),.dout(w_dff_B_UXJUApCm4_0),.clk(gclk));
	jdff dff_B_B7zaxIUB3_0(.din(w_dff_B_UXJUApCm4_0),.dout(w_dff_B_B7zaxIUB3_0),.clk(gclk));
	jdff dff_B_sHpu8Rdi2_0(.din(w_dff_B_B7zaxIUB3_0),.dout(w_dff_B_sHpu8Rdi2_0),.clk(gclk));
	jdff dff_B_gJEemIMr6_0(.din(w_dff_B_sHpu8Rdi2_0),.dout(w_dff_B_gJEemIMr6_0),.clk(gclk));
	jdff dff_B_P2GbtctS6_0(.din(w_dff_B_gJEemIMr6_0),.dout(w_dff_B_P2GbtctS6_0),.clk(gclk));
	jdff dff_B_UrjTCb297_0(.din(w_dff_B_P2GbtctS6_0),.dout(w_dff_B_UrjTCb297_0),.clk(gclk));
	jdff dff_B_Eb7ZkVKn9_0(.din(w_dff_B_UrjTCb297_0),.dout(w_dff_B_Eb7ZkVKn9_0),.clk(gclk));
	jdff dff_B_rSUdwkVl7_0(.din(w_dff_B_Eb7ZkVKn9_0),.dout(w_dff_B_rSUdwkVl7_0),.clk(gclk));
	jdff dff_B_LzkS9f5x3_1(.din(n745),.dout(w_dff_B_LzkS9f5x3_1),.clk(gclk));
	jdff dff_B_fX66LWDV4_0(.din(n747),.dout(w_dff_B_fX66LWDV4_0),.clk(gclk));
	jdff dff_B_DV69GAnb8_1(.din(n710),.dout(w_dff_B_DV69GAnb8_1),.clk(gclk));
	jdff dff_B_mXpOadW13_1(.din(w_dff_B_DV69GAnb8_1),.dout(w_dff_B_mXpOadW13_1),.clk(gclk));
	jdff dff_B_DVIPRSJw1_1(.din(w_dff_B_mXpOadW13_1),.dout(w_dff_B_DVIPRSJw1_1),.clk(gclk));
	jdff dff_B_CmOGlC6W4_1(.din(w_dff_B_DVIPRSJw1_1),.dout(w_dff_B_CmOGlC6W4_1),.clk(gclk));
	jdff dff_B_QBvwxmlc9_1(.din(w_dff_B_CmOGlC6W4_1),.dout(w_dff_B_QBvwxmlc9_1),.clk(gclk));
	jdff dff_B_GlkVDUc64_1(.din(w_dff_B_QBvwxmlc9_1),.dout(w_dff_B_GlkVDUc64_1),.clk(gclk));
	jdff dff_B_OerIHMfS6_1(.din(w_dff_B_GlkVDUc64_1),.dout(w_dff_B_OerIHMfS6_1),.clk(gclk));
	jdff dff_B_I0C8CyNJ4_1(.din(w_dff_B_OerIHMfS6_1),.dout(w_dff_B_I0C8CyNJ4_1),.clk(gclk));
	jdff dff_B_BBdJqaQv5_1(.din(w_dff_B_I0C8CyNJ4_1),.dout(w_dff_B_BBdJqaQv5_1),.clk(gclk));
	jdff dff_B_6nMD3evY1_1(.din(w_dff_B_BBdJqaQv5_1),.dout(w_dff_B_6nMD3evY1_1),.clk(gclk));
	jdff dff_B_sWmRlXx04_1(.din(w_dff_B_6nMD3evY1_1),.dout(w_dff_B_sWmRlXx04_1),.clk(gclk));
	jdff dff_B_tQ76jetn4_1(.din(w_dff_B_sWmRlXx04_1),.dout(w_dff_B_tQ76jetn4_1),.clk(gclk));
	jdff dff_B_c8QKqT2q2_1(.din(w_dff_B_tQ76jetn4_1),.dout(w_dff_B_c8QKqT2q2_1),.clk(gclk));
	jdff dff_B_s71eIqgP3_1(.din(w_dff_B_c8QKqT2q2_1),.dout(w_dff_B_s71eIqgP3_1),.clk(gclk));
	jdff dff_B_7wNTkWxA6_1(.din(w_dff_B_s71eIqgP3_1),.dout(w_dff_B_7wNTkWxA6_1),.clk(gclk));
	jdff dff_B_C0KWpf0w3_1(.din(w_dff_B_7wNTkWxA6_1),.dout(w_dff_B_C0KWpf0w3_1),.clk(gclk));
	jdff dff_B_kGrMpqO54_0(.din(n739),.dout(w_dff_B_kGrMpqO54_0),.clk(gclk));
	jdff dff_B_A9hHRejn5_0(.din(w_dff_B_kGrMpqO54_0),.dout(w_dff_B_A9hHRejn5_0),.clk(gclk));
	jdff dff_B_HxkD4b9J1_0(.din(w_dff_B_A9hHRejn5_0),.dout(w_dff_B_HxkD4b9J1_0),.clk(gclk));
	jdff dff_B_X9idg66l4_0(.din(n1127),.dout(w_dff_B_X9idg66l4_0),.clk(gclk));
	jdff dff_B_WY3neuGy6_0(.din(w_dff_B_X9idg66l4_0),.dout(w_dff_B_WY3neuGy6_0),.clk(gclk));
	jdff dff_B_ADgAvYvc2_0(.din(w_dff_B_WY3neuGy6_0),.dout(w_dff_B_ADgAvYvc2_0),.clk(gclk));
	jdff dff_B_tIvGYJEx6_1(.din(n1115),.dout(w_dff_B_tIvGYJEx6_1),.clk(gclk));
	jdff dff_B_9wjLRXn98_0(.din(n1118),.dout(w_dff_B_9wjLRXn98_0),.clk(gclk));
	jdff dff_B_A1EWhcBU9_0(.din(w_dff_B_9wjLRXn98_0),.dout(w_dff_B_A1EWhcBU9_0),.clk(gclk));
	jdff dff_B_yHsBKicb7_1(.din(n1117),.dout(w_dff_B_yHsBKicb7_1),.clk(gclk));
	jdff dff_B_SapRLWNS5_1(.din(w_dff_B_yHsBKicb7_1),.dout(w_dff_B_SapRLWNS5_1),.clk(gclk));
	jdff dff_B_OWuBgYMA9_1(.din(w_dff_B_SapRLWNS5_1),.dout(w_dff_B_OWuBgYMA9_1),.clk(gclk));
	jdff dff_B_VneAKUWQ0_1(.din(w_dff_B_OWuBgYMA9_1),.dout(w_dff_B_VneAKUWQ0_1),.clk(gclk));
	jdff dff_B_ABBEEnfy1_1(.din(w_dff_B_VneAKUWQ0_1),.dout(w_dff_B_ABBEEnfy1_1),.clk(gclk));
	jdff dff_A_CQmIbAnm1_1(.dout(w_n1113_0[1]),.din(w_dff_A_CQmIbAnm1_1),.clk(gclk));
	jdff dff_A_Le8kUKpP8_1(.dout(w_dff_A_CQmIbAnm1_1),.din(w_dff_A_Le8kUKpP8_1),.clk(gclk));
	jdff dff_A_DbV8GDW21_1(.dout(w_dff_A_Le8kUKpP8_1),.din(w_dff_A_DbV8GDW21_1),.clk(gclk));
	jdff dff_B_f9ngZ1SD7_0(.din(n1137),.dout(w_dff_B_f9ngZ1SD7_0),.clk(gclk));
	jdff dff_B_CzT4pdQb5_0(.din(w_dff_B_f9ngZ1SD7_0),.dout(w_dff_B_CzT4pdQb5_0),.clk(gclk));
	jdff dff_B_R4v33W5T8_0(.din(n1136),.dout(w_dff_B_R4v33W5T8_0),.clk(gclk));
	jdff dff_B_LnBZBnHP3_0(.din(w_dff_B_R4v33W5T8_0),.dout(w_dff_B_LnBZBnHP3_0),.clk(gclk));
	jdff dff_B_qOXUUY664_0(.din(w_dff_B_LnBZBnHP3_0),.dout(w_dff_B_qOXUUY664_0),.clk(gclk));
	jdff dff_B_14jL4H7C1_0(.din(w_dff_B_qOXUUY664_0),.dout(w_dff_B_14jL4H7C1_0),.clk(gclk));
	jdff dff_B_Sg4nGMbq9_0(.din(w_dff_B_14jL4H7C1_0),.dout(w_dff_B_Sg4nGMbq9_0),.clk(gclk));
	jdff dff_B_q6OC8l0N7_0(.din(w_dff_B_Sg4nGMbq9_0),.dout(w_dff_B_q6OC8l0N7_0),.clk(gclk));
	jdff dff_B_HBXTYAzj3_0(.din(w_dff_B_q6OC8l0N7_0),.dout(w_dff_B_HBXTYAzj3_0),.clk(gclk));
	jdff dff_B_lGAfzhEC2_0(.din(w_dff_B_HBXTYAzj3_0),.dout(w_dff_B_lGAfzhEC2_0),.clk(gclk));
	jdff dff_B_4MFQ0rBK2_0(.din(w_dff_B_lGAfzhEC2_0),.dout(w_dff_B_4MFQ0rBK2_0),.clk(gclk));
	jdff dff_B_UUZaD1jK0_0(.din(w_dff_B_4MFQ0rBK2_0),.dout(w_dff_B_UUZaD1jK0_0),.clk(gclk));
	jdff dff_B_dOZtQB3m0_0(.din(w_dff_B_UUZaD1jK0_0),.dout(w_dff_B_dOZtQB3m0_0),.clk(gclk));
	jdff dff_B_CIqPzpgN0_0(.din(w_dff_B_dOZtQB3m0_0),.dout(w_dff_B_CIqPzpgN0_0),.clk(gclk));
	jdff dff_B_r3jfSRTx8_0(.din(w_dff_B_CIqPzpgN0_0),.dout(w_dff_B_r3jfSRTx8_0),.clk(gclk));
	jdff dff_B_gMTsxEsl0_0(.din(w_dff_B_r3jfSRTx8_0),.dout(w_dff_B_gMTsxEsl0_0),.clk(gclk));
	jdff dff_B_QpmcwTas3_0(.din(w_dff_B_gMTsxEsl0_0),.dout(w_dff_B_QpmcwTas3_0),.clk(gclk));
	jdff dff_B_wxhLeqir4_0(.din(w_dff_B_QpmcwTas3_0),.dout(w_dff_B_wxhLeqir4_0),.clk(gclk));
	jdff dff_B_wZ0uvnqf6_0(.din(w_dff_B_wxhLeqir4_0),.dout(w_dff_B_wZ0uvnqf6_0),.clk(gclk));
	jdff dff_B_LTeDXujm0_0(.din(w_dff_B_wZ0uvnqf6_0),.dout(w_dff_B_LTeDXujm0_0),.clk(gclk));
	jdff dff_B_snArqUtM4_0(.din(w_dff_B_LTeDXujm0_0),.dout(w_dff_B_snArqUtM4_0),.clk(gclk));
	jdff dff_B_zP5YUKbg9_0(.din(w_dff_B_snArqUtM4_0),.dout(w_dff_B_zP5YUKbg9_0),.clk(gclk));
	jdff dff_B_m1rbH33D4_0(.din(w_dff_B_zP5YUKbg9_0),.dout(w_dff_B_m1rbH33D4_0),.clk(gclk));
	jdff dff_B_F7opRmds6_0(.din(w_dff_B_m1rbH33D4_0),.dout(w_dff_B_F7opRmds6_0),.clk(gclk));
	jdff dff_B_OqV6vmQM6_1(.din(G2897),.dout(w_dff_B_OqV6vmQM6_1),.clk(gclk));
	jdff dff_B_47RNrqGq8_2(.din(n1125),.dout(w_dff_B_47RNrqGq8_2),.clk(gclk));
	jdff dff_B_5Tpf33HU8_2(.din(w_dff_B_47RNrqGq8_2),.dout(w_dff_B_5Tpf33HU8_2),.clk(gclk));
	jdff dff_B_OA7DF1Bj6_2(.din(w_dff_B_5Tpf33HU8_2),.dout(w_dff_B_OA7DF1Bj6_2),.clk(gclk));
	jdff dff_B_Jgi8miKW4_2(.din(w_dff_B_OA7DF1Bj6_2),.dout(w_dff_B_Jgi8miKW4_2),.clk(gclk));
	jdff dff_B_5mrVt7GO1_2(.din(w_dff_B_Jgi8miKW4_2),.dout(w_dff_B_5mrVt7GO1_2),.clk(gclk));
	jdff dff_B_9EW4iv9v6_2(.din(w_dff_B_5mrVt7GO1_2),.dout(w_dff_B_9EW4iv9v6_2),.clk(gclk));
	jdff dff_B_9Aix1DWN2_2(.din(w_dff_B_9EW4iv9v6_2),.dout(w_dff_B_9Aix1DWN2_2),.clk(gclk));
	jdff dff_B_nWbrj5Xq9_2(.din(w_dff_B_9Aix1DWN2_2),.dout(w_dff_B_nWbrj5Xq9_2),.clk(gclk));
	jdff dff_B_L1ggevO54_2(.din(w_dff_B_nWbrj5Xq9_2),.dout(w_dff_B_L1ggevO54_2),.clk(gclk));
	jdff dff_B_uKvOAJjL1_2(.din(w_dff_B_L1ggevO54_2),.dout(w_dff_B_uKvOAJjL1_2),.clk(gclk));
	jdff dff_B_KGeqL9GY7_2(.din(w_dff_B_uKvOAJjL1_2),.dout(w_dff_B_KGeqL9GY7_2),.clk(gclk));
	jdff dff_B_54XVvIGB2_2(.din(w_dff_B_KGeqL9GY7_2),.dout(w_dff_B_54XVvIGB2_2),.clk(gclk));
	jdff dff_B_OKcuJluz3_2(.din(w_dff_B_54XVvIGB2_2),.dout(w_dff_B_OKcuJluz3_2),.clk(gclk));
	jdff dff_B_sgl3PZ2n2_2(.din(w_dff_B_OKcuJluz3_2),.dout(w_dff_B_sgl3PZ2n2_2),.clk(gclk));
	jdff dff_B_RY46vdQ46_2(.din(w_dff_B_sgl3PZ2n2_2),.dout(w_dff_B_RY46vdQ46_2),.clk(gclk));
	jdff dff_B_0U4xSHlJ0_2(.din(w_dff_B_RY46vdQ46_2),.dout(w_dff_B_0U4xSHlJ0_2),.clk(gclk));
	jdff dff_B_h5tQU98Z2_2(.din(w_dff_B_0U4xSHlJ0_2),.dout(w_dff_B_h5tQU98Z2_2),.clk(gclk));
	jdff dff_B_jvRKEBnT5_2(.din(w_dff_B_h5tQU98Z2_2),.dout(w_dff_B_jvRKEBnT5_2),.clk(gclk));
	jdff dff_B_Dt9CRmEA6_2(.din(w_dff_B_jvRKEBnT5_2),.dout(w_dff_B_Dt9CRmEA6_2),.clk(gclk));
	jdff dff_B_SYhdm9Wo2_2(.din(w_dff_B_Dt9CRmEA6_2),.dout(w_dff_B_SYhdm9Wo2_2),.clk(gclk));
	jdff dff_B_HwM3TxD34_2(.din(w_dff_B_SYhdm9Wo2_2),.dout(w_dff_B_HwM3TxD34_2),.clk(gclk));
	jdff dff_A_uFH8kqJz5_0(.dout(w_n1123_0[0]),.din(w_dff_A_uFH8kqJz5_0),.clk(gclk));
	jdff dff_A_zPreM2Rj7_0(.dout(w_dff_A_uFH8kqJz5_0),.din(w_dff_A_zPreM2Rj7_0),.clk(gclk));
	jdff dff_A_R7m49jkZ5_0(.dout(w_dff_A_zPreM2Rj7_0),.din(w_dff_A_R7m49jkZ5_0),.clk(gclk));
	jdff dff_A_CUwa98da6_0(.dout(w_dff_A_R7m49jkZ5_0),.din(w_dff_A_CUwa98da6_0),.clk(gclk));
	jdff dff_A_c7dW74vt0_0(.dout(w_dff_A_CUwa98da6_0),.din(w_dff_A_c7dW74vt0_0),.clk(gclk));
	jdff dff_A_WJqEKpoo6_0(.dout(w_dff_A_c7dW74vt0_0),.din(w_dff_A_WJqEKpoo6_0),.clk(gclk));
	jdff dff_A_ybUbKBm75_0(.dout(w_dff_A_WJqEKpoo6_0),.din(w_dff_A_ybUbKBm75_0),.clk(gclk));
	jdff dff_A_uRkVU4529_0(.dout(w_dff_A_ybUbKBm75_0),.din(w_dff_A_uRkVU4529_0),.clk(gclk));
	jdff dff_A_QfGNPeLp2_0(.dout(w_dff_A_uRkVU4529_0),.din(w_dff_A_QfGNPeLp2_0),.clk(gclk));
	jdff dff_A_j6Lurujp3_0(.dout(w_dff_A_QfGNPeLp2_0),.din(w_dff_A_j6Lurujp3_0),.clk(gclk));
	jdff dff_A_zIbyO1mU6_0(.dout(w_dff_A_j6Lurujp3_0),.din(w_dff_A_zIbyO1mU6_0),.clk(gclk));
	jdff dff_A_xUZBvXgV6_0(.dout(w_dff_A_zIbyO1mU6_0),.din(w_dff_A_xUZBvXgV6_0),.clk(gclk));
	jdff dff_A_oKYmP77o2_0(.dout(w_dff_A_xUZBvXgV6_0),.din(w_dff_A_oKYmP77o2_0),.clk(gclk));
	jdff dff_A_t5JRguzs0_0(.dout(w_dff_A_oKYmP77o2_0),.din(w_dff_A_t5JRguzs0_0),.clk(gclk));
	jdff dff_A_XvidrjEG4_0(.dout(w_dff_A_t5JRguzs0_0),.din(w_dff_A_XvidrjEG4_0),.clk(gclk));
	jdff dff_A_fTWY8M770_0(.dout(w_dff_A_XvidrjEG4_0),.din(w_dff_A_fTWY8M770_0),.clk(gclk));
	jdff dff_A_DbbxjWhF7_0(.dout(w_dff_A_fTWY8M770_0),.din(w_dff_A_DbbxjWhF7_0),.clk(gclk));
	jdff dff_A_qc4snaze3_0(.dout(w_dff_A_DbbxjWhF7_0),.din(w_dff_A_qc4snaze3_0),.clk(gclk));
	jdff dff_A_boRgIYP70_0(.dout(w_dff_A_qc4snaze3_0),.din(w_dff_A_boRgIYP70_0),.clk(gclk));
	jdff dff_A_lsCXNBZX3_0(.dout(w_dff_A_boRgIYP70_0),.din(w_dff_A_lsCXNBZX3_0),.clk(gclk));
	jdff dff_A_3PytOADh8_0(.dout(w_dff_A_lsCXNBZX3_0),.din(w_dff_A_3PytOADh8_0),.clk(gclk));
	jdff dff_A_QhKTE00P1_0(.dout(w_dff_A_3PytOADh8_0),.din(w_dff_A_QhKTE00P1_0),.clk(gclk));
	jdff dff_A_WHOdOuRe0_0(.dout(w_dff_A_QhKTE00P1_0),.din(w_dff_A_WHOdOuRe0_0),.clk(gclk));
	jdff dff_A_ljyVV2Qy8_0(.dout(w_n1134_0[0]),.din(w_dff_A_ljyVV2Qy8_0),.clk(gclk));
	jdff dff_A_dl8KQIxb6_0(.dout(w_dff_A_ljyVV2Qy8_0),.din(w_dff_A_dl8KQIxb6_0),.clk(gclk));
	jdff dff_A_kQQvnavx6_0(.dout(w_dff_A_dl8KQIxb6_0),.din(w_dff_A_kQQvnavx6_0),.clk(gclk));
	jdff dff_A_w5xjl9lA6_0(.dout(w_n1065_0[0]),.din(w_dff_A_w5xjl9lA6_0),.clk(gclk));
	jdff dff_A_0Q6EldbN6_1(.dout(w_n1065_0[1]),.din(w_dff_A_0Q6EldbN6_1),.clk(gclk));
	jdff dff_B_S8WVM1hS3_0(.din(n1064),.dout(w_dff_B_S8WVM1hS3_0),.clk(gclk));
	jdff dff_B_UZtwq4PO0_0(.din(w_dff_B_S8WVM1hS3_0),.dout(w_dff_B_UZtwq4PO0_0),.clk(gclk));
	jdff dff_B_3GSQrYB29_0(.din(w_dff_B_UZtwq4PO0_0),.dout(w_dff_B_3GSQrYB29_0),.clk(gclk));
	jdff dff_B_mxH9uoAT4_0(.din(w_dff_B_3GSQrYB29_0),.dout(w_dff_B_mxH9uoAT4_0),.clk(gclk));
	jdff dff_B_AXvvbDg23_0(.din(w_dff_B_mxH9uoAT4_0),.dout(w_dff_B_AXvvbDg23_0),.clk(gclk));
	jdff dff_B_RK1iR2RE8_0(.din(w_dff_B_AXvvbDg23_0),.dout(w_dff_B_RK1iR2RE8_0),.clk(gclk));
	jdff dff_B_DTWfMLSi6_0(.din(n1061),.dout(w_dff_B_DTWfMLSi6_0),.clk(gclk));
	jdff dff_B_U1ktPB0e7_0(.din(w_dff_B_DTWfMLSi6_0),.dout(w_dff_B_U1ktPB0e7_0),.clk(gclk));
	jdff dff_B_WS7OFj0P0_0(.din(w_dff_B_U1ktPB0e7_0),.dout(w_dff_B_WS7OFj0P0_0),.clk(gclk));
	jdff dff_B_nKk6nYl89_0(.din(w_dff_B_WS7OFj0P0_0),.dout(w_dff_B_nKk6nYl89_0),.clk(gclk));
	jdff dff_B_vCa5fqnJ1_1(.din(n1026),.dout(w_dff_B_vCa5fqnJ1_1),.clk(gclk));
	jdff dff_B_i6UbJX2C4_1(.din(w_dff_B_vCa5fqnJ1_1),.dout(w_dff_B_i6UbJX2C4_1),.clk(gclk));
	jdff dff_B_y37tZ4Lc5_1(.din(w_dff_B_i6UbJX2C4_1),.dout(w_dff_B_y37tZ4Lc5_1),.clk(gclk));
	jdff dff_B_9HOrcZI27_1(.din(w_dff_B_y37tZ4Lc5_1),.dout(w_dff_B_9HOrcZI27_1),.clk(gclk));
	jdff dff_B_Oqeoyf9n3_1(.din(w_dff_B_9HOrcZI27_1),.dout(w_dff_B_Oqeoyf9n3_1),.clk(gclk));
	jdff dff_B_zU2R2PzE4_1(.din(G124),.dout(w_dff_B_zU2R2PzE4_1),.clk(gclk));
	jdff dff_B_kC2ssVMQ9_1(.din(w_dff_B_zU2R2PzE4_1),.dout(w_dff_B_kC2ssVMQ9_1),.clk(gclk));
	jdff dff_B_cWQFdEAc9_1(.din(w_dff_B_kC2ssVMQ9_1),.dout(w_dff_B_cWQFdEAc9_1),.clk(gclk));
	jdff dff_B_5cZ1O0xr1_0(.din(n1020),.dout(w_dff_B_5cZ1O0xr1_0),.clk(gclk));
	jdff dff_B_2JA7K7KZ0_0(.din(w_dff_B_5cZ1O0xr1_0),.dout(w_dff_B_2JA7K7KZ0_0),.clk(gclk));
	jdff dff_A_OR4B7QlQ7_1(.dout(w_n1018_0[1]),.din(w_dff_A_OR4B7QlQ7_1),.clk(gclk));
	jdff dff_A_vGyWv8B62_1(.dout(w_dff_A_OR4B7QlQ7_1),.din(w_dff_A_vGyWv8B62_1),.clk(gclk));
	jdff dff_A_eUpbv59v7_1(.dout(w_dff_A_vGyWv8B62_1),.din(w_dff_A_eUpbv59v7_1),.clk(gclk));
	jdff dff_A_pz73L3iA4_1(.dout(w_dff_A_eUpbv59v7_1),.din(w_dff_A_pz73L3iA4_1),.clk(gclk));
	jdff dff_A_pYr5Q0wG0_1(.dout(w_dff_A_pz73L3iA4_1),.din(w_dff_A_pYr5Q0wG0_1),.clk(gclk));
	jdff dff_A_ICV7M9LY9_1(.dout(w_dff_A_pYr5Q0wG0_1),.din(w_dff_A_ICV7M9LY9_1),.clk(gclk));
	jdff dff_A_K3YCUiXo4_1(.dout(w_dff_A_ICV7M9LY9_1),.din(w_dff_A_K3YCUiXo4_1),.clk(gclk));
	jdff dff_A_BfDQ3R3W4_1(.dout(w_n725_0[1]),.din(w_dff_A_BfDQ3R3W4_1),.clk(gclk));
	jdff dff_A_kwK8aTq29_1(.dout(w_dff_A_BfDQ3R3W4_1),.din(w_dff_A_kwK8aTq29_1),.clk(gclk));
	jdff dff_A_Dowq88ls1_1(.dout(w_dff_A_kwK8aTq29_1),.din(w_dff_A_Dowq88ls1_1),.clk(gclk));
	jdff dff_B_uchyO9Lh0_1(.din(n712),.dout(w_dff_B_uchyO9Lh0_1),.clk(gclk));
	jdff dff_B_edmWya649_1(.din(w_dff_B_uchyO9Lh0_1),.dout(w_dff_B_edmWya649_1),.clk(gclk));
	jdff dff_B_vUDW9NkC7_1(.din(w_dff_B_edmWya649_1),.dout(w_dff_B_vUDW9NkC7_1),.clk(gclk));
	jdff dff_B_EV8IBihK4_1(.din(w_dff_B_vUDW9NkC7_1),.dout(w_dff_B_EV8IBihK4_1),.clk(gclk));
	jdff dff_B_EbJKsm921_1(.din(w_dff_B_EV8IBihK4_1),.dout(w_dff_B_EbJKsm921_1),.clk(gclk));
	jdff dff_B_Keavc4sM0_1(.din(w_dff_B_EbJKsm921_1),.dout(w_dff_B_Keavc4sM0_1),.clk(gclk));
	jdff dff_A_2kvRam4i1_0(.dout(w_n729_0[0]),.din(w_dff_A_2kvRam4i1_0),.clk(gclk));
	jdff dff_A_Zp6vcKg74_0(.dout(w_dff_A_2kvRam4i1_0),.din(w_dff_A_Zp6vcKg74_0),.clk(gclk));
	jdff dff_B_ElAcdpYs0_2(.din(n729),.dout(w_dff_B_ElAcdpYs0_2),.clk(gclk));
	jdff dff_B_HtTIFEwZ6_2(.din(w_dff_B_ElAcdpYs0_2),.dout(w_dff_B_HtTIFEwZ6_2),.clk(gclk));
	jdff dff_B_XckPm41r1_1(.din(n964),.dout(w_dff_B_XckPm41r1_1),.clk(gclk));
	jdff dff_B_f5m4rwjz6_0(.din(n1006),.dout(w_dff_B_f5m4rwjz6_0),.clk(gclk));
	jdff dff_B_smSuVHDx3_0(.din(w_dff_B_f5m4rwjz6_0),.dout(w_dff_B_smSuVHDx3_0),.clk(gclk));
	jdff dff_B_8mjbPghj8_0(.din(w_dff_B_smSuVHDx3_0),.dout(w_dff_B_8mjbPghj8_0),.clk(gclk));
	jdff dff_B_mBpWAGl59_0(.din(w_dff_B_8mjbPghj8_0),.dout(w_dff_B_mBpWAGl59_0),.clk(gclk));
	jdff dff_B_BlWMooR57_0(.din(w_dff_B_mBpWAGl59_0),.dout(w_dff_B_BlWMooR57_0),.clk(gclk));
	jdff dff_B_s905FG0E6_0(.din(w_dff_B_BlWMooR57_0),.dout(w_dff_B_s905FG0E6_0),.clk(gclk));
	jdff dff_B_IgFdMaRH6_0(.din(n1004),.dout(w_dff_B_IgFdMaRH6_0),.clk(gclk));
	jdff dff_B_EGBK8yHP2_0(.din(w_dff_B_IgFdMaRH6_0),.dout(w_dff_B_EGBK8yHP2_0),.clk(gclk));
	jdff dff_B_u08wbZlj7_0(.din(w_dff_B_EGBK8yHP2_0),.dout(w_dff_B_u08wbZlj7_0),.clk(gclk));
	jdff dff_B_HvPTZidA6_0(.din(w_dff_B_u08wbZlj7_0),.dout(w_dff_B_HvPTZidA6_0),.clk(gclk));
	jdff dff_B_bvJN8E9G5_1(.din(n1000),.dout(w_dff_B_bvJN8E9G5_1),.clk(gclk));
	jdff dff_B_f35JV3Ep9_2(.din(G125),.dout(w_dff_B_f35JV3Ep9_2),.clk(gclk));
	jdff dff_B_hrXs8Eb47_2(.din(w_dff_B_f35JV3Ep9_2),.dout(w_dff_B_hrXs8Eb47_2),.clk(gclk));
	jdff dff_B_3ciWDK0f1_2(.din(w_dff_B_hrXs8Eb47_2),.dout(w_dff_B_3ciWDK0f1_2),.clk(gclk));
	jdff dff_B_LciRUnhA4_0(.din(n963),.dout(w_dff_B_LciRUnhA4_0),.clk(gclk));
	jdff dff_A_dadJwbjL5_1(.dout(w_n961_0[1]),.din(w_dff_A_dadJwbjL5_1),.clk(gclk));
	jdff dff_A_v9rMCZ7a8_1(.dout(w_dff_A_dadJwbjL5_1),.din(w_dff_A_v9rMCZ7a8_1),.clk(gclk));
	jdff dff_B_H1vwYt9V7_0(.din(n960),.dout(w_dff_B_H1vwYt9V7_0),.clk(gclk));
	jdff dff_B_vZGGj2Qm5_0(.din(w_dff_B_H1vwYt9V7_0),.dout(w_dff_B_vZGGj2Qm5_0),.clk(gclk));
	jdff dff_A_gdJhmvkv7_1(.dout(w_n715_0[1]),.din(w_dff_A_gdJhmvkv7_1),.clk(gclk));
	jdff dff_A_ADenmync1_1(.dout(w_dff_A_gdJhmvkv7_1),.din(w_dff_A_ADenmync1_1),.clk(gclk));
	jdff dff_B_DkZ3iT6Y7_2(.din(n715),.dout(w_dff_B_DkZ3iT6Y7_2),.clk(gclk));
	jdff dff_B_oCNxCbQi4_2(.din(w_dff_B_DkZ3iT6Y7_2),.dout(w_dff_B_oCNxCbQi4_2),.clk(gclk));
	jdff dff_B_8HkJADyj7_2(.din(w_dff_B_oCNxCbQi4_2),.dout(w_dff_B_8HkJADyj7_2),.clk(gclk));
	jdff dff_B_UeLHqPQg9_0(.din(n955),.dout(w_dff_B_UeLHqPQg9_0),.clk(gclk));
	jdff dff_B_b2BqNUgk9_0(.din(w_dff_B_UeLHqPQg9_0),.dout(w_dff_B_b2BqNUgk9_0),.clk(gclk));
	jdff dff_A_EQI4XA034_0(.dout(w_n726_0[0]),.din(w_dff_A_EQI4XA034_0),.clk(gclk));
	jdff dff_A_5eegF3ti5_0(.dout(w_dff_A_EQI4XA034_0),.din(w_dff_A_5eegF3ti5_0),.clk(gclk));
	jdff dff_A_BrlEhjNb0_0(.dout(w_dff_A_5eegF3ti5_0),.din(w_dff_A_BrlEhjNb0_0),.clk(gclk));
	jdff dff_A_097lohcG9_2(.dout(w_n714_0[2]),.din(w_dff_A_097lohcG9_2),.clk(gclk));
	jdff dff_A_fYNL4EM06_2(.dout(w_dff_A_097lohcG9_2),.din(w_dff_A_fYNL4EM06_2),.clk(gclk));
	jdff dff_A_ma02ySPw1_2(.dout(w_dff_A_fYNL4EM06_2),.din(w_dff_A_ma02ySPw1_2),.clk(gclk));
	jdff dff_A_3eRvBS125_2(.dout(w_dff_A_ma02ySPw1_2),.din(w_dff_A_3eRvBS125_2),.clk(gclk));
	jdff dff_A_dOiBy7mD3_2(.dout(w_dff_A_3eRvBS125_2),.din(w_dff_A_dOiBy7mD3_2),.clk(gclk));
	jdff dff_B_kWlhMqib3_0(.din(n713),.dout(w_dff_B_kWlhMqib3_0),.clk(gclk));
	jdff dff_B_RbEAYj8h2_0(.din(n1132),.dout(w_dff_B_RbEAYj8h2_0),.clk(gclk));
	jdff dff_B_58Zn26et7_0(.din(n1110),.dout(w_dff_B_58Zn26et7_0),.clk(gclk));
	jdff dff_B_5Kh7yM324_0(.din(n1109),.dout(w_dff_B_5Kh7yM324_0),.clk(gclk));
	jdff dff_B_oqr6lieX7_0(.din(w_dff_B_5Kh7yM324_0),.dout(w_dff_B_oqr6lieX7_0),.clk(gclk));
	jdff dff_B_XBbiO69Z5_0(.din(w_dff_B_oqr6lieX7_0),.dout(w_dff_B_XBbiO69Z5_0),.clk(gclk));
	jdff dff_B_Fu5xcM1d2_0(.din(w_dff_B_XBbiO69Z5_0),.dout(w_dff_B_Fu5xcM1d2_0),.clk(gclk));
	jdff dff_B_NEbCJ37P3_0(.din(w_dff_B_Fu5xcM1d2_0),.dout(w_dff_B_NEbCJ37P3_0),.clk(gclk));
	jdff dff_B_U1vlPODo9_0(.din(w_dff_B_NEbCJ37P3_0),.dout(w_dff_B_U1vlPODo9_0),.clk(gclk));
	jdff dff_B_vrgbrAzy6_0(.din(w_dff_B_U1vlPODo9_0),.dout(w_dff_B_vrgbrAzy6_0),.clk(gclk));
	jdff dff_B_M3as2jdR2_0(.din(n1107),.dout(w_dff_B_M3as2jdR2_0),.clk(gclk));
	jdff dff_B_L7D1CmnO6_0(.din(w_dff_B_M3as2jdR2_0),.dout(w_dff_B_L7D1CmnO6_0),.clk(gclk));
	jdff dff_B_vWvobxQE9_1(.din(n1103),.dout(w_dff_B_vWvobxQE9_1),.clk(gclk));
	jdff dff_B_1iIe0ggf8_1(.din(w_dff_B_vWvobxQE9_1),.dout(w_dff_B_1iIe0ggf8_1),.clk(gclk));
	jdff dff_B_mjwmoLdh9_1(.din(w_dff_B_1iIe0ggf8_1),.dout(w_dff_B_mjwmoLdh9_1),.clk(gclk));
	jdff dff_B_LkLvAd1X5_0(.din(n1104),.dout(w_dff_B_LkLvAd1X5_0),.clk(gclk));
	jdff dff_B_fq1EQPkL3_0(.din(w_dff_B_LkLvAd1X5_0),.dout(w_dff_B_fq1EQPkL3_0),.clk(gclk));
	jdff dff_B_Kt8Pkl8Y8_3(.din(G128),.dout(w_dff_B_Kt8Pkl8Y8_3),.clk(gclk));
	jdff dff_B_3snf7RKg4_3(.din(w_dff_B_Kt8Pkl8Y8_3),.dout(w_dff_B_3snf7RKg4_3),.clk(gclk));
	jdff dff_B_LoEDOQo05_3(.din(w_dff_B_3snf7RKg4_3),.dout(w_dff_B_LoEDOQo05_3),.clk(gclk));
	jdff dff_A_5FM9sSZX4_0(.dout(w_G50_2[0]),.din(w_dff_A_5FM9sSZX4_0),.clk(gclk));
	jdff dff_A_2HSi2V1s9_0(.dout(w_dff_A_5FM9sSZX4_0),.din(w_dff_A_2HSi2V1s9_0),.clk(gclk));
	jdff dff_A_zBJPXltE3_0(.dout(w_dff_A_2HSi2V1s9_0),.din(w_dff_A_zBJPXltE3_0),.clk(gclk));
	jdff dff_A_JXUbd1bh4_2(.dout(w_G50_2[2]),.din(w_dff_A_JXUbd1bh4_2),.clk(gclk));
	jdff dff_A_nfeQYIfl6_2(.dout(w_dff_A_JXUbd1bh4_2),.din(w_dff_A_nfeQYIfl6_2),.clk(gclk));
	jdff dff_A_c0hMX5Af4_2(.dout(w_dff_A_nfeQYIfl6_2),.din(w_dff_A_c0hMX5Af4_2),.clk(gclk));
	jdff dff_A_PXNzbcOa8_0(.dout(w_n1011_0[0]),.din(w_dff_A_PXNzbcOa8_0),.clk(gclk));
	jdff dff_A_LngoYsIR5_0(.dout(w_dff_A_PXNzbcOa8_0),.din(w_dff_A_LngoYsIR5_0),.clk(gclk));
	jdff dff_A_gKySxZzv8_0(.dout(w_n727_0[0]),.din(w_dff_A_gKySxZzv8_0),.clk(gclk));
	jdff dff_A_US7ki9f44_0(.dout(w_dff_A_gKySxZzv8_0),.din(w_dff_A_US7ki9f44_0),.clk(gclk));
	jdff dff_A_vwztvN8M5_0(.dout(w_dff_A_US7ki9f44_0),.din(w_dff_A_vwztvN8M5_0),.clk(gclk));
	jdff dff_A_W8tnGj2F9_0(.dout(w_dff_A_vwztvN8M5_0),.din(w_dff_A_W8tnGj2F9_0),.clk(gclk));
	jdff dff_A_19aJx0qV7_0(.dout(w_dff_A_W8tnGj2F9_0),.din(w_dff_A_19aJx0qV7_0),.clk(gclk));
	jdff dff_A_3HDi1XbW8_1(.dout(w_n727_0[1]),.din(w_dff_A_3HDi1XbW8_1),.clk(gclk));
	jdff dff_A_0qUpa6Nl8_1(.dout(w_dff_A_3HDi1XbW8_1),.din(w_dff_A_0qUpa6Nl8_1),.clk(gclk));
	jdff dff_A_dO770lKP4_1(.dout(w_dff_A_0qUpa6Nl8_1),.din(w_dff_A_dO770lKP4_1),.clk(gclk));
	jdff dff_A_POjjuOXP3_1(.dout(w_dff_A_dO770lKP4_1),.din(w_dff_A_POjjuOXP3_1),.clk(gclk));
	jdff dff_A_pcYsestV9_1(.dout(w_dff_A_POjjuOXP3_1),.din(w_dff_A_pcYsestV9_1),.clk(gclk));
	jdff dff_B_3DM4Z68X4_3(.din(n727),.dout(w_dff_B_3DM4Z68X4_3),.clk(gclk));
	jdff dff_A_y0rI58hY0_1(.dout(w_n721_1[1]),.din(w_dff_A_y0rI58hY0_1),.clk(gclk));
	jdff dff_A_phUlYsr64_1(.dout(w_dff_A_y0rI58hY0_1),.din(w_dff_A_phUlYsr64_1),.clk(gclk));
	jdff dff_A_WYqfzLwj0_1(.dout(w_dff_A_phUlYsr64_1),.din(w_dff_A_WYqfzLwj0_1),.clk(gclk));
	jdff dff_A_Ohcw8xeW9_1(.dout(w_dff_A_WYqfzLwj0_1),.din(w_dff_A_Ohcw8xeW9_1),.clk(gclk));
	jdff dff_A_gOIn9MML3_1(.dout(w_dff_A_Ohcw8xeW9_1),.din(w_dff_A_gOIn9MML3_1),.clk(gclk));
	jdff dff_A_I5Tqi5Xu2_2(.dout(w_n721_0[2]),.din(w_dff_A_I5Tqi5Xu2_2),.clk(gclk));
	jdff dff_A_os8MM3Za8_2(.dout(w_dff_A_I5Tqi5Xu2_2),.din(w_dff_A_os8MM3Za8_2),.clk(gclk));
	jdff dff_A_0LaYx7rt6_2(.dout(w_dff_A_os8MM3Za8_2),.din(w_dff_A_0LaYx7rt6_2),.clk(gclk));
	jdff dff_A_nsu0JxYL4_2(.dout(w_dff_A_0LaYx7rt6_2),.din(w_dff_A_nsu0JxYL4_2),.clk(gclk));
	jdff dff_A_vR5rV29I9_2(.dout(w_dff_A_nsu0JxYL4_2),.din(w_dff_A_vR5rV29I9_2),.clk(gclk));
	jdff dff_A_wvhqducA2_2(.dout(w_dff_A_vR5rV29I9_2),.din(w_dff_A_wvhqducA2_2),.clk(gclk));
	jdff dff_A_MMgmZvqe4_2(.dout(w_dff_A_wvhqducA2_2),.din(w_dff_A_MMgmZvqe4_2),.clk(gclk));
	jdff dff_A_FxRl3JTB6_0(.dout(w_n718_0[0]),.din(w_dff_A_FxRl3JTB6_0),.clk(gclk));
	jdff dff_A_MA0rPdw98_0(.dout(w_dff_A_FxRl3JTB6_0),.din(w_dff_A_MA0rPdw98_0),.clk(gclk));
	jdff dff_A_Zb2QFsoF3_0(.dout(w_dff_A_MA0rPdw98_0),.din(w_dff_A_Zb2QFsoF3_0),.clk(gclk));
	jdff dff_A_Dl6pYAmz1_1(.dout(w_n718_0[1]),.din(w_dff_A_Dl6pYAmz1_1),.clk(gclk));
	jdff dff_A_yaO282oz6_1(.dout(w_dff_A_Dl6pYAmz1_1),.din(w_dff_A_yaO282oz6_1),.clk(gclk));
	jdff dff_A_GhUoLhoJ8_1(.dout(w_dff_A_yaO282oz6_1),.din(w_dff_A_GhUoLhoJ8_1),.clk(gclk));
	jdff dff_A_IsgXaCh32_1(.dout(w_n717_0[1]),.din(w_dff_A_IsgXaCh32_1),.clk(gclk));
	jdff dff_A_9Bk1bKCu0_0(.dout(w_n948_0[0]),.din(w_dff_A_9Bk1bKCu0_0),.clk(gclk));
	jdff dff_A_QKVqJgMz7_0(.dout(w_dff_A_9Bk1bKCu0_0),.din(w_dff_A_QKVqJgMz7_0),.clk(gclk));
	jdff dff_A_JU99Oa223_0(.dout(w_n738_0[0]),.din(w_dff_A_JU99Oa223_0),.clk(gclk));
	jdff dff_A_MRR3uDbp7_0(.dout(w_dff_A_JU99Oa223_0),.din(w_dff_A_MRR3uDbp7_0),.clk(gclk));
	jdff dff_A_dUpis0yX9_0(.dout(w_dff_A_MRR3uDbp7_0),.din(w_dff_A_dUpis0yX9_0),.clk(gclk));
	jdff dff_A_qj9iYWu55_0(.dout(w_n531_2[0]),.din(w_dff_A_qj9iYWu55_0),.clk(gclk));
	jdff dff_A_miCrs79F0_0(.dout(w_dff_A_qj9iYWu55_0),.din(w_dff_A_miCrs79F0_0),.clk(gclk));
	jdff dff_A_6htQD5nO4_0(.dout(w_dff_A_miCrs79F0_0),.din(w_dff_A_6htQD5nO4_0),.clk(gclk));
	jdff dff_A_t6jLmTvA9_0(.dout(w_dff_A_6htQD5nO4_0),.din(w_dff_A_t6jLmTvA9_0),.clk(gclk));
	jdff dff_A_ycXKvQzM5_0(.dout(w_dff_A_t6jLmTvA9_0),.din(w_dff_A_ycXKvQzM5_0),.clk(gclk));
	jdff dff_A_AFBer5jh7_0(.dout(w_dff_A_ycXKvQzM5_0),.din(w_dff_A_AFBer5jh7_0),.clk(gclk));
	jdff dff_A_gsVQJr0B7_2(.dout(w_n531_2[2]),.din(w_dff_A_gsVQJr0B7_2),.clk(gclk));
	jdff dff_A_tBWwSSqg8_2(.dout(w_dff_A_gsVQJr0B7_2),.din(w_dff_A_tBWwSSqg8_2),.clk(gclk));
	jdff dff_A_vH9QyFAH4_0(.dout(w_n525_0[0]),.din(w_dff_A_vH9QyFAH4_0),.clk(gclk));
	jdff dff_B_OJKARMjA2_1(.din(n519),.dout(w_dff_B_OJKARMjA2_1),.clk(gclk));
	jdff dff_A_t45hlgsX8_0(.dout(w_n487_0[0]),.din(w_dff_A_t45hlgsX8_0),.clk(gclk));
	jdff dff_A_sS1Clive5_0(.dout(w_dff_A_t45hlgsX8_0),.din(w_dff_A_sS1Clive5_0),.clk(gclk));
	jdff dff_A_o8MNwIAq7_1(.dout(w_n487_0[1]),.din(w_dff_A_o8MNwIAq7_1),.clk(gclk));
	jdff dff_A_wp8QsmI95_1(.dout(w_dff_A_o8MNwIAq7_1),.din(w_dff_A_wp8QsmI95_1),.clk(gclk));
	jdff dff_A_6qQ0zdwa5_1(.dout(w_dff_A_wp8QsmI95_1),.din(w_dff_A_6qQ0zdwa5_1),.clk(gclk));
	jdff dff_A_F8KG0rd27_1(.dout(w_dff_A_6qQ0zdwa5_1),.din(w_dff_A_F8KG0rd27_1),.clk(gclk));
	jdff dff_B_JwVbT8Ib5_3(.din(n487),.dout(w_dff_B_JwVbT8Ib5_3),.clk(gclk));
	jdff dff_B_AHRCaxL13_3(.din(w_dff_B_JwVbT8Ib5_3),.dout(w_dff_B_AHRCaxL13_3),.clk(gclk));
	jdff dff_A_5FAdf8by2_0(.dout(w_n486_0[0]),.din(w_dff_A_5FAdf8by2_0),.clk(gclk));
	jdff dff_A_Ph6wgQJk7_0(.dout(w_dff_A_5FAdf8by2_0),.din(w_dff_A_Ph6wgQJk7_0),.clk(gclk));
	jdff dff_A_FNp8w6bp1_0(.dout(w_dff_A_Ph6wgQJk7_0),.din(w_dff_A_FNp8w6bp1_0),.clk(gclk));
	jdff dff_B_bXb4hhhe3_0(.din(n485),.dout(w_dff_B_bXb4hhhe3_0),.clk(gclk));
	jdff dff_A_vQK9rPe47_0(.dout(w_n484_0[0]),.din(w_dff_A_vQK9rPe47_0),.clk(gclk));
	jdff dff_B_mRGVovu76_1(.din(n477),.dout(w_dff_B_mRGVovu76_1),.clk(gclk));
	jdff dff_B_XKI9VZ5k9_1(.din(w_dff_B_mRGVovu76_1),.dout(w_dff_B_XKI9VZ5k9_1),.clk(gclk));
	jdff dff_B_H0JpnCjm0_1(.din(w_dff_B_XKI9VZ5k9_1),.dout(w_dff_B_H0JpnCjm0_1),.clk(gclk));
	jdff dff_B_2tHWsNiR9_0(.din(n479),.dout(w_dff_B_2tHWsNiR9_0),.clk(gclk));
	jdff dff_A_Hfd7It0H9_1(.dout(w_n476_0[1]),.din(w_dff_A_Hfd7It0H9_1),.clk(gclk));
	jdff dff_A_B46Hbzmp1_2(.dout(w_n476_0[2]),.din(w_dff_A_B46Hbzmp1_2),.clk(gclk));
	jdff dff_B_R08Ih9bi6_1(.din(n459),.dout(w_dff_B_R08Ih9bi6_1),.clk(gclk));
	jdff dff_B_N05izYLT1_1(.din(w_dff_B_R08Ih9bi6_1),.dout(w_dff_B_N05izYLT1_1),.clk(gclk));
	jdff dff_B_azvrYdGl8_0(.din(n470),.dout(w_dff_B_azvrYdGl8_0),.clk(gclk));
	jdff dff_B_2c7q3EWk1_0(.din(w_dff_B_azvrYdGl8_0),.dout(w_dff_B_2c7q3EWk1_0),.clk(gclk));
	jdff dff_A_J1Hp3aej6_0(.dout(w_n108_1[0]),.din(w_dff_A_J1Hp3aej6_0),.clk(gclk));
	jdff dff_A_ar5rILi53_0(.dout(w_dff_A_J1Hp3aej6_0),.din(w_dff_A_ar5rILi53_0),.clk(gclk));
	jdff dff_A_Z4bHatZS4_0(.dout(w_dff_A_ar5rILi53_0),.din(w_dff_A_Z4bHatZS4_0),.clk(gclk));
	jdff dff_A_WDdd8SeS3_1(.dout(w_n108_0[1]),.din(w_dff_A_WDdd8SeS3_1),.clk(gclk));
	jdff dff_A_XYjb7VEd5_1(.dout(w_dff_A_WDdd8SeS3_1),.din(w_dff_A_XYjb7VEd5_1),.clk(gclk));
	jdff dff_A_73UYEdBJ2_1(.dout(w_dff_A_XYjb7VEd5_1),.din(w_dff_A_73UYEdBJ2_1),.clk(gclk));
	jdff dff_B_8MCw01Rg0_1(.din(n463),.dout(w_dff_B_8MCw01Rg0_1),.clk(gclk));
	jdff dff_A_yDkvygq41_1(.dout(w_n449_0[1]),.din(w_dff_A_yDkvygq41_1),.clk(gclk));
	jdff dff_B_XI3alUZC5_1(.din(n444),.dout(w_dff_B_XI3alUZC5_1),.clk(gclk));
	jdff dff_B_wG9g4L8p8_1(.din(w_dff_B_XI3alUZC5_1),.dout(w_dff_B_wG9g4L8p8_1),.clk(gclk));
	jdff dff_B_UU5jplzl4_0(.din(n441),.dout(w_dff_B_UU5jplzl4_0),.clk(gclk));
	jdff dff_B_AMvP1x4O6_0(.din(n438),.dout(w_dff_B_AMvP1x4O6_0),.clk(gclk));
	jdff dff_B_YoXN2Ew11_0(.din(w_dff_B_AMvP1x4O6_0),.dout(w_dff_B_YoXN2Ew11_0),.clk(gclk));
	jdff dff_A_zZbqqVKJ0_0(.dout(w_n99_1[0]),.din(w_dff_A_zZbqqVKJ0_0),.clk(gclk));
	jdff dff_A_TLdDlbQB2_1(.dout(w_n99_1[1]),.din(w_dff_A_TLdDlbQB2_1),.clk(gclk));
	jdff dff_A_3KBrRDM28_1(.dout(w_dff_A_TLdDlbQB2_1),.din(w_dff_A_3KBrRDM28_1),.clk(gclk));
	jdff dff_A_3z5vq90N2_1(.dout(w_dff_A_3KBrRDM28_1),.din(w_dff_A_3z5vq90N2_1),.clk(gclk));
	jdff dff_B_fCpVejhE2_1(.din(n429),.dout(w_dff_B_fCpVejhE2_1),.clk(gclk));
	jdff dff_B_dbxYtjsB5_1(.din(w_dff_B_fCpVejhE2_1),.dout(w_dff_B_dbxYtjsB5_1),.clk(gclk));
	jdff dff_B_1i9JVmsm0_1(.din(G222),.dout(w_dff_B_1i9JVmsm0_1),.clk(gclk));
	jdff dff_B_wO9YYGgD8_1(.din(w_dff_B_1i9JVmsm0_1),.dout(w_dff_B_wO9YYGgD8_1),.clk(gclk));
	jdff dff_B_GJ5XoSC99_2(.din(G223),.dout(w_dff_B_GJ5XoSC99_2),.clk(gclk));
	jdff dff_B_HboFerw58_2(.din(w_dff_B_GJ5XoSC99_2),.dout(w_dff_B_HboFerw58_2),.clk(gclk));
	jdff dff_A_UXK1BWGK5_0(.dout(w_n415_0[0]),.din(w_dff_A_UXK1BWGK5_0),.clk(gclk));
	jdff dff_A_WGFVMaPx8_1(.dout(w_n415_0[1]),.din(w_dff_A_WGFVMaPx8_1),.clk(gclk));
	jdff dff_A_FW53Yhps1_1(.dout(w_dff_A_WGFVMaPx8_1),.din(w_dff_A_FW53Yhps1_1),.clk(gclk));
	jdff dff_A_akqUpS582_1(.dout(w_dff_A_FW53Yhps1_1),.din(w_dff_A_akqUpS582_1),.clk(gclk));
	jdff dff_B_0I7edd237_1(.din(n410),.dout(w_dff_B_0I7edd237_1),.clk(gclk));
	jdff dff_B_z3fMj7fk0_1(.din(w_dff_B_0I7edd237_1),.dout(w_dff_B_z3fMj7fk0_1),.clk(gclk));
	jdff dff_A_3iuqr9z28_0(.dout(w_n409_0[0]),.din(w_dff_A_3iuqr9z28_0),.clk(gclk));
	jdff dff_A_wSx9gRti9_0(.dout(w_dff_A_3iuqr9z28_0),.din(w_dff_A_wSx9gRti9_0),.clk(gclk));
	jdff dff_A_DS0kuLJX4_0(.dout(w_dff_A_wSx9gRti9_0),.din(w_dff_A_DS0kuLJX4_0),.clk(gclk));
	jdff dff_A_L5ZUWAUW0_0(.dout(w_dff_A_DS0kuLJX4_0),.din(w_dff_A_L5ZUWAUW0_0),.clk(gclk));
	jdff dff_B_vud1sdUj5_0(.din(n407),.dout(w_dff_B_vud1sdUj5_0),.clk(gclk));
	jdff dff_B_yWflXVes1_0(.din(n404),.dout(w_dff_B_yWflXVes1_0),.clk(gclk));
	jdff dff_B_msIF60Dn0_0(.din(w_dff_B_yWflXVes1_0),.dout(w_dff_B_msIF60Dn0_0),.clk(gclk));
	jdff dff_A_FwUPWvLI2_0(.dout(w_n103_1[0]),.din(w_dff_A_FwUPWvLI2_0),.clk(gclk));
	jdff dff_A_W2Ki44GS9_1(.dout(w_n103_0[1]),.din(w_dff_A_W2Ki44GS9_1),.clk(gclk));
	jdff dff_A_8anq8RjV4_1(.dout(w_dff_A_W2Ki44GS9_1),.din(w_dff_A_8anq8RjV4_1),.clk(gclk));
	jdff dff_A_p26f3lRV2_1(.dout(w_dff_A_8anq8RjV4_1),.din(w_dff_A_p26f3lRV2_1),.clk(gclk));
	jdff dff_A_W091tQYi5_0(.dout(w_n394_0[0]),.din(w_dff_A_W091tQYi5_0),.clk(gclk));
	jdff dff_B_b5ePqyXQ6_2(.din(n394),.dout(w_dff_B_b5ePqyXQ6_2),.clk(gclk));
	jdff dff_B_kYwFt9Yr7_2(.din(n1114),.dout(w_dff_B_kYwFt9Yr7_2),.clk(gclk));
	jdff dff_B_btql5Epw5_2(.din(w_dff_B_kYwFt9Yr7_2),.dout(w_dff_B_btql5Epw5_2),.clk(gclk));
	jdff dff_B_gmp3csBQ2_2(.din(w_dff_B_btql5Epw5_2),.dout(w_dff_B_gmp3csBQ2_2),.clk(gclk));
	jdff dff_B_FZ4kgAJ67_2(.din(w_dff_B_gmp3csBQ2_2),.dout(w_dff_B_FZ4kgAJ67_2),.clk(gclk));
	jdff dff_B_HLIqN8EU8_2(.din(w_dff_B_FZ4kgAJ67_2),.dout(w_dff_B_HLIqN8EU8_2),.clk(gclk));
	jdff dff_A_UxchZKH33_1(.dout(G384),.din(w_dff_A_UxchZKH33_1),.clk(gclk));
	jdff dff_B_xHpBB69J6_1(.din(n700),.dout(w_dff_B_xHpBB69J6_1),.clk(gclk));
	jdff dff_B_yE92zG6r5_1(.din(w_dff_B_xHpBB69J6_1),.dout(w_dff_B_yE92zG6r5_1),.clk(gclk));
	jdff dff_B_UqFtJkCs7_1(.din(w_dff_B_yE92zG6r5_1),.dout(w_dff_B_UqFtJkCs7_1),.clk(gclk));
	jdff dff_A_LJrLFR8L9_0(.dout(w_n703_0[0]),.din(w_dff_A_LJrLFR8L9_0),.clk(gclk));
	jdff dff_A_Jwcz2mmN1_0(.dout(w_dff_A_LJrLFR8L9_0),.din(w_dff_A_Jwcz2mmN1_0),.clk(gclk));
	jdff dff_A_Vr0d0vvE7_0(.dout(w_dff_A_Jwcz2mmN1_0),.din(w_dff_A_Vr0d0vvE7_0),.clk(gclk));
	jdff dff_A_VWO1Fd9K5_2(.dout(w_n703_0[2]),.din(w_dff_A_VWO1Fd9K5_2),.clk(gclk));
	jdff dff_A_DIwyCqDw2_2(.dout(w_dff_A_VWO1Fd9K5_2),.din(w_dff_A_DIwyCqDw2_2),.clk(gclk));
	jdff dff_A_5TScZkiy6_1(.dout(w_n701_0[1]),.din(w_dff_A_5TScZkiy6_1),.clk(gclk));
	jdff dff_B_gN2NqprP1_0(.din(n699),.dout(w_dff_B_gN2NqprP1_0),.clk(gclk));
	jdff dff_B_nM1Ib5xW8_0(.din(w_dff_B_gN2NqprP1_0),.dout(w_dff_B_nM1Ib5xW8_0),.clk(gclk));
	jdff dff_B_WXPU0Eer4_0(.din(w_dff_B_nM1Ib5xW8_0),.dout(w_dff_B_WXPU0Eer4_0),.clk(gclk));
	jdff dff_B_ThjMCZdC7_0(.din(w_dff_B_WXPU0Eer4_0),.dout(w_dff_B_ThjMCZdC7_0),.clk(gclk));
	jdff dff_B_lorWBVYy3_0(.din(w_dff_B_ThjMCZdC7_0),.dout(w_dff_B_lorWBVYy3_0),.clk(gclk));
	jdff dff_B_n51VEqSr3_0(.din(n697),.dout(w_dff_B_n51VEqSr3_0),.clk(gclk));
	jdff dff_A_fDXdL3SA3_0(.dout(w_G150_3[0]),.din(w_dff_A_fDXdL3SA3_0),.clk(gclk));
	jdff dff_B_DBRdK7Kn4_3(.din(G132),.dout(w_dff_B_DBRdK7Kn4_3),.clk(gclk));
	jdff dff_B_VW85mSJm6_3(.din(w_dff_B_DBRdK7Kn4_3),.dout(w_dff_B_VW85mSJm6_3),.clk(gclk));
	jdff dff_B_RxdeFCrb9_3(.din(w_dff_B_VW85mSJm6_3),.dout(w_dff_B_RxdeFCrb9_3),.clk(gclk));
	jdff dff_A_lq1gdekD5_0(.dout(w_n578_1[0]),.din(w_dff_A_lq1gdekD5_0),.clk(gclk));
	jdff dff_A_fzmmIHUK9_0(.dout(w_dff_A_lq1gdekD5_0),.din(w_dff_A_fzmmIHUK9_0),.clk(gclk));
	jdff dff_A_Arvo39BC6_0(.dout(w_dff_A_fzmmIHUK9_0),.din(w_dff_A_Arvo39BC6_0),.clk(gclk));
	jdff dff_A_kHuGlsUy6_0(.dout(w_dff_A_Arvo39BC6_0),.din(w_dff_A_kHuGlsUy6_0),.clk(gclk));
	jdff dff_A_7z3M0q8G9_0(.dout(w_dff_A_kHuGlsUy6_0),.din(w_dff_A_7z3M0q8G9_0),.clk(gclk));
	jdff dff_A_XnzcFuZW6_0(.dout(w_dff_A_7z3M0q8G9_0),.din(w_dff_A_XnzcFuZW6_0),.clk(gclk));
	jdff dff_A_ptrud9cU5_0(.dout(w_dff_A_XnzcFuZW6_0),.din(w_dff_A_ptrud9cU5_0),.clk(gclk));
	jdff dff_A_yUptmQBo9_1(.dout(w_n578_1[1]),.din(w_dff_A_yUptmQBo9_1),.clk(gclk));
	jdff dff_A_BaDMvh899_1(.dout(w_dff_A_yUptmQBo9_1),.din(w_dff_A_BaDMvh899_1),.clk(gclk));
	jdff dff_A_gAyzsRWo3_1(.dout(w_dff_A_BaDMvh899_1),.din(w_dff_A_gAyzsRWo3_1),.clk(gclk));
	jdff dff_A_6IkSOGA19_1(.dout(w_dff_A_gAyzsRWo3_1),.din(w_dff_A_6IkSOGA19_1),.clk(gclk));
	jdff dff_A_siOXgMss2_1(.dout(w_dff_A_6IkSOGA19_1),.din(w_dff_A_siOXgMss2_1),.clk(gclk));
	jdff dff_A_SSDiQdoU2_1(.dout(w_dff_A_siOXgMss2_1),.din(w_dff_A_SSDiQdoU2_1),.clk(gclk));
	jdff dff_A_P7Rv0l8F9_1(.dout(w_dff_A_SSDiQdoU2_1),.din(w_dff_A_P7Rv0l8F9_1),.clk(gclk));
	jdff dff_A_afHsN3HE2_1(.dout(w_dff_A_P7Rv0l8F9_1),.din(w_dff_A_afHsN3HE2_1),.clk(gclk));
	jdff dff_B_qegTJfwP3_0(.din(n657),.dout(w_dff_B_qegTJfwP3_0),.clk(gclk));
	jdff dff_B_2VSmEWrt8_0(.din(w_dff_B_qegTJfwP3_0),.dout(w_dff_B_2VSmEWrt8_0),.clk(gclk));
	jdff dff_B_HMjhaAFe1_0(.din(w_dff_B_2VSmEWrt8_0),.dout(w_dff_B_HMjhaAFe1_0),.clk(gclk));
	jdff dff_B_yXkkCsrs6_0(.din(w_dff_B_HMjhaAFe1_0),.dout(w_dff_B_yXkkCsrs6_0),.clk(gclk));
	jdff dff_A_XWryLDgY7_0(.dout(w_n381_0[0]),.din(w_dff_A_XWryLDgY7_0),.clk(gclk));
	jdff dff_A_qDMZAbvO3_0(.dout(w_dff_A_XWryLDgY7_0),.din(w_dff_A_qDMZAbvO3_0),.clk(gclk));
	jdff dff_A_DoPik7nl2_0(.dout(w_dff_A_qDMZAbvO3_0),.din(w_dff_A_DoPik7nl2_0),.clk(gclk));
	jdff dff_B_2lravuW69_0(.din(n379),.dout(w_dff_B_2lravuW69_0),.clk(gclk));
	jdff dff_B_afLhG7oH1_0(.din(n373),.dout(w_dff_B_afLhG7oH1_0),.clk(gclk));
	jdff dff_A_zfRA3oVw7_2(.dout(w_n191_2[2]),.din(w_dff_A_zfRA3oVw7_2),.clk(gclk));
	jdff dff_A_27yDXbBi6_2(.dout(w_dff_A_zfRA3oVw7_2),.din(w_dff_A_27yDXbBi6_2),.clk(gclk));
	jdff dff_A_41I9nSRK2_1(.dout(w_n371_0[1]),.din(w_dff_A_41I9nSRK2_1),.clk(gclk));
	jdff dff_B_klgUUWDg7_2(.din(n371),.dout(w_dff_B_klgUUWDg7_2),.clk(gclk));
	jdff dff_B_CwEn7Y6z2_1(.din(n361),.dout(w_dff_B_CwEn7Y6z2_1),.clk(gclk));
	jdff dff_B_DXhI0XcQ3_0(.din(n368),.dout(w_dff_B_DXhI0XcQ3_0),.clk(gclk));
	jdff dff_A_iOpRD2AB1_1(.dout(w_n73_0[1]),.din(w_dff_A_iOpRD2AB1_1),.clk(gclk));
	jdff dff_A_ra2ovdSy7_1(.dout(w_dff_A_iOpRD2AB1_1),.din(w_dff_A_ra2ovdSy7_1),.clk(gclk));
	jdff dff_A_XCor1GRt1_1(.dout(w_dff_A_ra2ovdSy7_1),.din(w_dff_A_XCor1GRt1_1),.clk(gclk));
	jdff dff_A_VKlXmtLv3_2(.dout(w_n73_0[2]),.din(w_dff_A_VKlXmtLv3_2),.clk(gclk));
	jdff dff_A_n1rNZ6VJ4_2(.dout(w_dff_A_VKlXmtLv3_2),.din(w_dff_A_n1rNZ6VJ4_2),.clk(gclk));
	jdff dff_B_Yxob6LeF8_1(.din(n363),.dout(w_dff_B_Yxob6LeF8_1),.clk(gclk));
	jdff dff_A_xRweCtHC4_1(.dout(w_G58_5[1]),.din(w_dff_A_xRweCtHC4_1),.clk(gclk));
	jdff dff_A_HRH4bXPe7_1(.dout(w_dff_A_xRweCtHC4_1),.din(w_dff_A_HRH4bXPe7_1),.clk(gclk));
	jdff dff_A_gLmHOx7C6_2(.dout(w_G58_5[2]),.din(w_dff_A_gLmHOx7C6_2),.clk(gclk));
	jdff dff_A_kXI2QyuQ6_0(.dout(w_n357_0[0]),.din(w_dff_A_kXI2QyuQ6_0),.clk(gclk));
	jdff dff_B_90XzA1Er2_2(.din(n357),.dout(w_dff_B_90XzA1Er2_2),.clk(gclk));
	jdff dff_A_zOeZyDd71_2(.dout(w_n142_2[2]),.din(w_dff_A_zOeZyDd71_2),.clk(gclk));
	jdff dff_B_fPnJjukF7_0(.din(n347),.dout(w_dff_B_fPnJjukF7_0),.clk(gclk));
	jdff dff_B_cjLmZ3eg8_0(.din(n346),.dout(w_dff_B_cjLmZ3eg8_0),.clk(gclk));
	jdff dff_A_qKWFEasm0_1(.dout(w_n342_0[1]),.din(w_dff_A_qKWFEasm0_1),.clk(gclk));
	jdff dff_A_WB9p8lUe4_1(.dout(w_dff_A_qKWFEasm0_1),.din(w_dff_A_WB9p8lUe4_1),.clk(gclk));
	jdff dff_A_4kvJkFvK4_1(.dout(w_dff_A_WB9p8lUe4_1),.din(w_dff_A_4kvJkFvK4_1),.clk(gclk));
	jdff dff_A_SaZw2CP78_1(.dout(w_n341_0[1]),.din(w_dff_A_SaZw2CP78_1),.clk(gclk));
	jdff dff_B_z6hjKqff5_1(.din(n1129),.dout(w_dff_B_z6hjKqff5_1),.clk(gclk));
	jdff dff_B_BAtwaBZ78_1(.din(w_dff_B_z6hjKqff5_1),.dout(w_dff_B_BAtwaBZ78_1),.clk(gclk));
	jdff dff_B_ZZIZqtV64_1(.din(n940),.dout(w_dff_B_ZZIZqtV64_1),.clk(gclk));
	jdff dff_B_V6zxnBaT1_1(.din(w_dff_B_ZZIZqtV64_1),.dout(w_dff_B_V6zxnBaT1_1),.clk(gclk));
	jdff dff_B_Ed9eR1hD6_1(.din(w_dff_B_V6zxnBaT1_1),.dout(w_dff_B_Ed9eR1hD6_1),.clk(gclk));
	jdff dff_B_JMR7Jm0s6_1(.din(w_dff_B_Ed9eR1hD6_1),.dout(w_dff_B_JMR7Jm0s6_1),.clk(gclk));
	jdff dff_B_Z5oLgYEv9_1(.din(w_dff_B_JMR7Jm0s6_1),.dout(w_dff_B_Z5oLgYEv9_1),.clk(gclk));
	jdff dff_B_WcwNvsPZ5_1(.din(w_dff_B_Z5oLgYEv9_1),.dout(w_dff_B_WcwNvsPZ5_1),.clk(gclk));
	jdff dff_B_d37Ewm1F7_1(.din(n941),.dout(w_dff_B_d37Ewm1F7_1),.clk(gclk));
	jdff dff_B_7ogxw4qH9_1(.din(w_dff_B_d37Ewm1F7_1),.dout(w_dff_B_7ogxw4qH9_1),.clk(gclk));
	jdff dff_B_O54W1JxW3_0(.din(n938),.dout(w_dff_B_O54W1JxW3_0),.clk(gclk));
	jdff dff_B_uQHEYYsw4_0(.din(w_dff_B_O54W1JxW3_0),.dout(w_dff_B_uQHEYYsw4_0),.clk(gclk));
	jdff dff_B_eGPjewSt7_0(.din(w_dff_B_uQHEYYsw4_0),.dout(w_dff_B_eGPjewSt7_0),.clk(gclk));
	jdff dff_B_tNfVI2BL3_0(.din(w_dff_B_eGPjewSt7_0),.dout(w_dff_B_tNfVI2BL3_0),.clk(gclk));
	jdff dff_B_LtshSjJE2_0(.din(w_dff_B_tNfVI2BL3_0),.dout(w_dff_B_LtshSjJE2_0),.clk(gclk));
	jdff dff_B_ALmO11cs1_0(.din(w_dff_B_LtshSjJE2_0),.dout(w_dff_B_ALmO11cs1_0),.clk(gclk));
	jdff dff_B_ShVlZ9431_1(.din(n904),.dout(w_dff_B_ShVlZ9431_1),.clk(gclk));
	jdff dff_B_SzLMeSQE7_0(.din(n936),.dout(w_dff_B_SzLMeSQE7_0),.clk(gclk));
	jdff dff_B_QSPc2gnM7_1(.din(n901),.dout(w_dff_B_QSPc2gnM7_1),.clk(gclk));
	jdff dff_B_D5X8rJBq2_0(.din(n902),.dout(w_dff_B_D5X8rJBq2_0),.clk(gclk));
	jdff dff_A_s2WD0Y0I5_0(.dout(w_n138_0[0]),.din(w_dff_A_s2WD0Y0I5_0),.clk(gclk));
	jdff dff_B_56hO7Xjw7_0(.din(n137),.dout(w_dff_B_56hO7Xjw7_0),.clk(gclk));
	jdff dff_A_EBAejq0L1_2(.dout(w_G97_2[2]),.din(w_dff_A_EBAejq0L1_2),.clk(gclk));
	jdff dff_A_auJTCT6x6_0(.dout(w_n832_0[0]),.din(w_dff_A_auJTCT6x6_0),.clk(gclk));
	jdff dff_A_7qDifxOM7_0(.dout(w_dff_A_auJTCT6x6_0),.din(w_dff_A_7qDifxOM7_0),.clk(gclk));
	jdff dff_A_BuIzhQVL9_0(.dout(w_dff_A_7qDifxOM7_0),.din(w_dff_A_BuIzhQVL9_0),.clk(gclk));
	jdff dff_A_u1JnJXQ80_0(.dout(w_dff_A_BuIzhQVL9_0),.din(w_dff_A_u1JnJXQ80_0),.clk(gclk));
	jdff dff_A_Eh9zIp8q1_1(.dout(w_n832_0[1]),.din(w_dff_A_Eh9zIp8q1_1),.clk(gclk));
	jdff dff_A_CgbQ7OTl9_1(.dout(w_dff_A_Eh9zIp8q1_1),.din(w_dff_A_CgbQ7OTl9_1),.clk(gclk));
	jdff dff_A_cuvHcPcG3_1(.dout(w_dff_A_CgbQ7OTl9_1),.din(w_dff_A_cuvHcPcG3_1),.clk(gclk));
	jdff dff_A_JciXvHZn2_1(.dout(w_dff_A_cuvHcPcG3_1),.din(w_dff_A_JciXvHZn2_1),.clk(gclk));
	jdff dff_B_iPrd9TeX5_0(.din(n828),.dout(w_dff_B_iPrd9TeX5_0),.clk(gclk));
	jdff dff_A_vodGdxag8_0(.dout(w_n827_0[0]),.din(w_dff_A_vodGdxag8_0),.clk(gclk));
	jdff dff_A_f96N0cPC9_0(.dout(w_dff_A_vodGdxag8_0),.din(w_dff_A_f96N0cPC9_0),.clk(gclk));
	jdff dff_A_nR4R98C65_1(.dout(w_n827_0[1]),.din(w_dff_A_nR4R98C65_1),.clk(gclk));
	jdff dff_A_ANdly2E41_1(.dout(w_dff_A_nR4R98C65_1),.din(w_dff_A_ANdly2E41_1),.clk(gclk));
	jdff dff_A_jdBXqUPm7_1(.dout(w_dff_A_ANdly2E41_1),.din(w_dff_A_jdBXqUPm7_1),.clk(gclk));
	jdff dff_B_hbgj2NQa0_2(.din(n542),.dout(w_dff_B_hbgj2NQa0_2),.clk(gclk));
	jdff dff_B_t1HLMZXK2_2(.din(w_dff_B_hbgj2NQa0_2),.dout(w_dff_B_t1HLMZXK2_2),.clk(gclk));
	jdff dff_B_c9IpNzOX5_0(.din(n817),.dout(w_dff_B_c9IpNzOX5_0),.clk(gclk));
	jdff dff_B_7uTgNvTx3_0(.din(w_dff_B_c9IpNzOX5_0),.dout(w_dff_B_7uTgNvTx3_0),.clk(gclk));
	jdff dff_B_gZvYO2tJ3_0(.din(n814),.dout(w_dff_B_gZvYO2tJ3_0),.clk(gclk));
	jdff dff_B_JZwssl0w9_0(.din(w_dff_B_gZvYO2tJ3_0),.dout(w_dff_B_JZwssl0w9_0),.clk(gclk));
	jdff dff_B_6mI38QDp5_0(.din(w_dff_B_JZwssl0w9_0),.dout(w_dff_B_6mI38QDp5_0),.clk(gclk));
	jdff dff_B_7RaG3MoD4_0(.din(w_dff_B_6mI38QDp5_0),.dout(w_dff_B_7RaG3MoD4_0),.clk(gclk));
	jdff dff_B_erdOwoPR9_0(.din(w_dff_B_7RaG3MoD4_0),.dout(w_dff_B_erdOwoPR9_0),.clk(gclk));
	jdff dff_B_CX9qtM3w1_1(.din(n808),.dout(w_dff_B_CX9qtM3w1_1),.clk(gclk));
	jdff dff_B_3DYUwprA2_1(.din(n809),.dout(w_dff_B_3DYUwprA2_1),.clk(gclk));
	jdff dff_B_7nbBkGuI5_0(.din(n811),.dout(w_dff_B_7nbBkGuI5_0),.clk(gclk));
	jdff dff_A_XIOaokYB8_0(.dout(w_n127_0[0]),.din(w_dff_A_XIOaokYB8_0),.clk(gclk));
	jdff dff_B_HMDYWvaT5_0(.din(n126),.dout(w_dff_B_HMDYWvaT5_0),.clk(gclk));
	jdff dff_B_nHjT9ivE9_3(.din(G143),.dout(w_dff_B_nHjT9ivE9_3),.clk(gclk));
	jdff dff_B_7jNdzNhw0_3(.din(w_dff_B_nHjT9ivE9_3),.dout(w_dff_B_7jNdzNhw0_3),.clk(gclk));
	jdff dff_B_DnzrD0rl8_3(.din(w_dff_B_7jNdzNhw0_3),.dout(w_dff_B_DnzrD0rl8_3),.clk(gclk));
	jdff dff_B_2MkF5Ibi1_3(.din(G137),.dout(w_dff_B_2MkF5Ibi1_3),.clk(gclk));
	jdff dff_B_FJ0yVpZr8_3(.din(w_dff_B_2MkF5Ibi1_3),.dout(w_dff_B_FJ0yVpZr8_3),.clk(gclk));
	jdff dff_B_zrwlyaUU3_3(.din(w_dff_B_FJ0yVpZr8_3),.dout(w_dff_B_zrwlyaUU3_3),.clk(gclk));
	jdff dff_A_Th4JHEbi6_0(.dout(w_n634_3[0]),.din(w_dff_A_Th4JHEbi6_0),.clk(gclk));
	jdff dff_A_nSuweLyS0_0(.dout(w_dff_A_Th4JHEbi6_0),.din(w_dff_A_nSuweLyS0_0),.clk(gclk));
	jdff dff_A_BLmq1XbH5_1(.dout(w_n634_3[1]),.din(w_dff_A_BLmq1XbH5_1),.clk(gclk));
	jdff dff_A_Ih9jq9Sa3_1(.dout(w_dff_A_BLmq1XbH5_1),.din(w_dff_A_Ih9jq9Sa3_1),.clk(gclk));
	jdff dff_A_2ylipEtU7_0(.dout(w_n771_0[0]),.din(w_dff_A_2ylipEtU7_0),.clk(gclk));
	jdff dff_B_gj7NzOOx8_1(.din(n757),.dout(w_dff_B_gj7NzOOx8_1),.clk(gclk));
	jdff dff_B_gyCkCVW80_0(.din(n769),.dout(w_dff_B_gyCkCVW80_0),.clk(gclk));
	jdff dff_A_1oitqJRV5_1(.dout(w_n768_0[1]),.din(w_dff_A_1oitqJRV5_1),.clk(gclk));
	jdff dff_A_7RI8VtIk1_1(.dout(w_dff_A_1oitqJRV5_1),.din(w_dff_A_7RI8VtIk1_1),.clk(gclk));
	jdff dff_A_l6PcCziw9_1(.dout(w_dff_A_7RI8VtIk1_1),.din(w_dff_A_l6PcCziw9_1),.clk(gclk));
	jdff dff_A_hlWLWior1_1(.dout(w_dff_A_l6PcCziw9_1),.din(w_dff_A_hlWLWior1_1),.clk(gclk));
	jdff dff_B_Tgc52uHY7_0(.din(n767),.dout(w_dff_B_Tgc52uHY7_0),.clk(gclk));
	jdff dff_B_bZqFMHI27_0(.din(w_dff_B_Tgc52uHY7_0),.dout(w_dff_B_bZqFMHI27_0),.clk(gclk));
	jdff dff_B_rqhWIE9n5_1(.din(n759),.dout(w_dff_B_rqhWIE9n5_1),.clk(gclk));
	jdff dff_B_v658yW0u7_1(.din(w_dff_B_rqhWIE9n5_1),.dout(w_dff_B_v658yW0u7_1),.clk(gclk));
	jdff dff_B_iYrA9RZ57_1(.din(w_dff_B_v658yW0u7_1),.dout(w_dff_B_iYrA9RZ57_1),.clk(gclk));
	jdff dff_B_lJMPZ3y32_0(.din(n756),.dout(w_dff_B_lJMPZ3y32_0),.clk(gclk));
	jdff dff_A_tV0FgGOD4_1(.dout(w_n755_0[1]),.din(w_dff_A_tV0FgGOD4_1),.clk(gclk));
	jdff dff_A_MxRcqYg14_1(.dout(w_dff_A_tV0FgGOD4_1),.din(w_dff_A_MxRcqYg14_1),.clk(gclk));
	jdff dff_A_5OB9D1s01_1(.dout(w_dff_A_MxRcqYg14_1),.din(w_dff_A_5OB9D1s01_1),.clk(gclk));
	jdff dff_B_QHGupD9O5_0(.din(n754),.dout(w_dff_B_QHGupD9O5_0),.clk(gclk));
	jdff dff_B_CYKxdWpc3_0(.din(w_dff_B_QHGupD9O5_0),.dout(w_dff_B_CYKxdWpc3_0),.clk(gclk));
	jdff dff_B_7FoqHNTg6_0(.din(w_dff_B_CYKxdWpc3_0),.dout(w_dff_B_7FoqHNTg6_0),.clk(gclk));
	jdff dff_B_enwv1RSk2_0(.din(w_dff_B_7FoqHNTg6_0),.dout(w_dff_B_enwv1RSk2_0),.clk(gclk));
	jdff dff_B_fRfLC7wP3_0(.din(w_dff_B_enwv1RSk2_0),.dout(w_dff_B_fRfLC7wP3_0),.clk(gclk));
	jdff dff_B_naovNozt1_0(.din(n896),.dout(w_dff_B_naovNozt1_0),.clk(gclk));
	jdff dff_B_kSPUY3b25_0(.din(w_dff_B_naovNozt1_0),.dout(w_dff_B_kSPUY3b25_0),.clk(gclk));
	jdff dff_B_30CLogu30_0(.din(w_dff_B_kSPUY3b25_0),.dout(w_dff_B_30CLogu30_0),.clk(gclk));
	jdff dff_B_nyCuQUXp5_0(.din(w_dff_B_30CLogu30_0),.dout(w_dff_B_nyCuQUXp5_0),.clk(gclk));
	jdff dff_B_popybWGT3_0(.din(w_dff_B_nyCuQUXp5_0),.dout(w_dff_B_popybWGT3_0),.clk(gclk));
	jdff dff_B_EoVue6r71_0(.din(n893),.dout(w_dff_B_EoVue6r71_0),.clk(gclk));
	jdff dff_B_uVYZmFoa2_0(.din(w_dff_B_EoVue6r71_0),.dout(w_dff_B_uVYZmFoa2_0),.clk(gclk));
	jdff dff_B_jUyMRLqf9_1(.din(n875),.dout(w_dff_B_jUyMRLqf9_1),.clk(gclk));
	jdff dff_B_HxXAlIrC8_1(.din(w_dff_B_jUyMRLqf9_1),.dout(w_dff_B_HxXAlIrC8_1),.clk(gclk));
	jdff dff_B_6QpDm6ob6_1(.din(w_dff_B_HxXAlIrC8_1),.dout(w_dff_B_6QpDm6ob6_1),.clk(gclk));
	jdff dff_B_ELOV9xVH7_1(.din(w_dff_B_6QpDm6ob6_1),.dout(w_dff_B_ELOV9xVH7_1),.clk(gclk));
	jdff dff_B_1OG4qX6U7_1(.din(n877),.dout(w_dff_B_1OG4qX6U7_1),.clk(gclk));
	jdff dff_B_LlUIFToS7_1(.din(w_dff_B_1OG4qX6U7_1),.dout(w_dff_B_LlUIFToS7_1),.clk(gclk));
	jdff dff_B_Fc1BDKqS9_0(.din(n889),.dout(w_dff_B_Fc1BDKqS9_0),.clk(gclk));
	jdff dff_B_F3XZmJmq0_0(.din(w_dff_B_Fc1BDKqS9_0),.dout(w_dff_B_F3XZmJmq0_0),.clk(gclk));
	jdff dff_B_rVv7XDPP0_0(.din(n887),.dout(w_dff_B_rVv7XDPP0_0),.clk(gclk));
	jdff dff_A_lKgum9Dc3_0(.dout(w_G58_2[0]),.din(w_dff_A_lKgum9Dc3_0),.clk(gclk));
	jdff dff_A_M2LnEw7Y9_0(.dout(w_dff_A_lKgum9Dc3_0),.din(w_dff_A_M2LnEw7Y9_0),.clk(gclk));
	jdff dff_A_Zv3tUhWl4_1(.dout(w_G58_2[1]),.din(w_dff_A_Zv3tUhWl4_1),.clk(gclk));
	jdff dff_A_zFPCULDU7_1(.dout(w_dff_A_Zv3tUhWl4_1),.din(w_dff_A_zFPCULDU7_1),.clk(gclk));
	jdff dff_A_5amnptMJ8_1(.dout(w_n99_0[1]),.din(w_dff_A_5amnptMJ8_1),.clk(gclk));
	jdff dff_A_9QSiTYBb6_1(.dout(w_dff_A_5amnptMJ8_1),.din(w_dff_A_9QSiTYBb6_1),.clk(gclk));
	jdff dff_A_LPCp8wUi4_1(.dout(w_dff_A_9QSiTYBb6_1),.din(w_dff_A_LPCp8wUi4_1),.clk(gclk));
	jdff dff_B_FmJuE4933_0(.din(n882),.dout(w_dff_B_FmJuE4933_0),.clk(gclk));
	jdff dff_B_zJiB3lEY7_0(.din(w_dff_B_FmJuE4933_0),.dout(w_dff_B_zJiB3lEY7_0),.clk(gclk));
	jdff dff_B_YqXng1Tl4_0(.din(n881),.dout(w_dff_B_YqXng1Tl4_0),.clk(gclk));
	jdff dff_A_DaGiIoEz7_1(.dout(w_n131_0[1]),.din(w_dff_A_DaGiIoEz7_1),.clk(gclk));
	jdff dff_B_Cvdy09qm7_0(.din(n130),.dout(w_dff_B_Cvdy09qm7_0),.clk(gclk));
	jdff dff_A_ILbNzyuE6_1(.dout(w_G232_0[1]),.din(w_dff_A_ILbNzyuE6_1),.clk(gclk));
	jdff dff_A_TNYJ7iBL0_1(.dout(w_dff_A_ILbNzyuE6_1),.din(w_dff_A_TNYJ7iBL0_1),.clk(gclk));
	jdff dff_A_XQmfFHEB3_1(.dout(w_dff_A_TNYJ7iBL0_1),.din(w_dff_A_XQmfFHEB3_1),.clk(gclk));
	jdff dff_A_PHS2RXKV3_2(.dout(w_G232_0[2]),.din(w_dff_A_PHS2RXKV3_2),.clk(gclk));
	jdff dff_A_bXd2SWAe9_2(.dout(w_dff_A_PHS2RXKV3_2),.din(w_dff_A_bXd2SWAe9_2),.clk(gclk));
	jdff dff_A_LX63CiXg6_0(.dout(w_G226_1[0]),.din(w_dff_A_LX63CiXg6_0),.clk(gclk));
	jdff dff_A_MFW7rTmx9_0(.dout(w_dff_A_LX63CiXg6_0),.din(w_dff_A_MFW7rTmx9_0),.clk(gclk));
	jdff dff_A_CqdVymKg8_1(.dout(w_G226_0[1]),.din(w_dff_A_CqdVymKg8_1),.clk(gclk));
	jdff dff_A_Pw3VdEjM4_1(.dout(w_dff_A_CqdVymKg8_1),.din(w_dff_A_Pw3VdEjM4_1),.clk(gclk));
	jdff dff_A_zIsp6HRb7_2(.dout(w_G226_0[2]),.din(w_dff_A_zIsp6HRb7_2),.clk(gclk));
	jdff dff_A_6cENp0FW9_2(.dout(w_dff_A_zIsp6HRb7_2),.din(w_dff_A_6cENp0FW9_2),.clk(gclk));
	jdff dff_A_bgcYkwPV5_2(.dout(w_dff_A_6cENp0FW9_2),.din(w_dff_A_bgcYkwPV5_2),.clk(gclk));
	jdff dff_A_c577wqMH2_1(.dout(w_n810_0[1]),.din(w_dff_A_c577wqMH2_1),.clk(gclk));
	jdff dff_A_5RTE3ISJ7_1(.dout(w_dff_A_c577wqMH2_1),.din(w_dff_A_5RTE3ISJ7_1),.clk(gclk));
	jdff dff_A_nZ7gWBPL1_1(.dout(w_dff_A_5RTE3ISJ7_1),.din(w_dff_A_nZ7gWBPL1_1),.clk(gclk));
	jdff dff_A_guwEpJeY9_0(.dout(w_G150_0[0]),.din(w_dff_A_guwEpJeY9_0),.clk(gclk));
	jdff dff_A_nvKubPcz8_1(.dout(w_G150_0[1]),.din(w_dff_A_nvKubPcz8_1),.clk(gclk));
	jdff dff_B_tyhBi3LE7_3(.din(G150),.dout(w_dff_B_tyhBi3LE7_3),.clk(gclk));
	jdff dff_B_KH0k5irM5_3(.din(w_dff_B_tyhBi3LE7_3),.dout(w_dff_B_KH0k5irM5_3),.clk(gclk));
	jdff dff_A_TkmKvSnH5_0(.dout(w_G77_2[0]),.din(w_dff_A_TkmKvSnH5_0),.clk(gclk));
	jdff dff_A_6rWT0e2E1_0(.dout(w_dff_A_TkmKvSnH5_0),.din(w_dff_A_6rWT0e2E1_0),.clk(gclk));
	jdff dff_A_4OZnzc347_1(.dout(w_G77_2[1]),.din(w_dff_A_4OZnzc347_1),.clk(gclk));
	jdff dff_A_3PFdd2zu2_1(.dout(w_dff_A_4OZnzc347_1),.din(w_dff_A_3PFdd2zu2_1),.clk(gclk));
	jdff dff_A_tdhUzLrN3_0(.dout(w_G58_3[0]),.din(w_dff_A_tdhUzLrN3_0),.clk(gclk));
	jdff dff_A_ksnOaavp9_0(.dout(w_dff_A_tdhUzLrN3_0),.din(w_dff_A_ksnOaavp9_0),.clk(gclk));
	jdff dff_A_3vO6REX67_0(.dout(w_dff_A_ksnOaavp9_0),.din(w_dff_A_3vO6REX67_0),.clk(gclk));
	jdff dff_A_LHtDBGoa3_1(.dout(w_G58_3[1]),.din(w_dff_A_LHtDBGoa3_1),.clk(gclk));
	jdff dff_A_J0e7aXRe2_1(.dout(w_dff_A_LHtDBGoa3_1),.din(w_dff_A_J0e7aXRe2_1),.clk(gclk));
	jdff dff_A_VhN3Y8XQ5_1(.dout(w_dff_A_J0e7aXRe2_1),.din(w_dff_A_VhN3Y8XQ5_1),.clk(gclk));
	jdff dff_A_dSupes7L3_1(.dout(w_G68_2[1]),.din(w_dff_A_dSupes7L3_1),.clk(gclk));
	jdff dff_A_Vs8BAEzk3_1(.dout(w_dff_A_dSupes7L3_1),.din(w_dff_A_Vs8BAEzk3_1),.clk(gclk));
	jdff dff_A_NipjuKUi1_1(.dout(w_dff_A_Vs8BAEzk3_1),.din(w_dff_A_NipjuKUi1_1),.clk(gclk));
	jdff dff_A_FC3MZrhx5_2(.dout(w_G68_2[2]),.din(w_dff_A_FC3MZrhx5_2),.clk(gclk));
	jdff dff_A_v9gX4OE79_2(.dout(w_dff_A_FC3MZrhx5_2),.din(w_dff_A_v9gX4OE79_2),.clk(gclk));
	jdff dff_A_AlWz1lJ56_2(.dout(w_dff_A_v9gX4OE79_2),.din(w_dff_A_AlWz1lJ56_2),.clk(gclk));
	jdff dff_A_kcHBLyaI9_0(.dout(w_n574_2[0]),.din(w_dff_A_kcHBLyaI9_0),.clk(gclk));
	jdff dff_A_3YfeII840_2(.dout(w_n574_2[2]),.din(w_dff_A_3YfeII840_2),.clk(gclk));
	jdff dff_A_X8XzmPe39_2(.dout(w_dff_A_3YfeII840_2),.din(w_dff_A_X8XzmPe39_2),.clk(gclk));
	jdff dff_A_e2PL1fzF4_2(.dout(w_dff_A_X8XzmPe39_2),.din(w_dff_A_e2PL1fzF4_2),.clk(gclk));
	jdff dff_A_BwHLonLY8_2(.dout(w_dff_A_e2PL1fzF4_2),.din(w_dff_A_BwHLonLY8_2),.clk(gclk));
	jdff dff_A_XN7tJbQv3_2(.dout(w_dff_A_BwHLonLY8_2),.din(w_dff_A_XN7tJbQv3_2),.clk(gclk));
	jdff dff_A_9dFVMJ195_2(.dout(w_dff_A_XN7tJbQv3_2),.din(w_dff_A_9dFVMJ195_2),.clk(gclk));
	jdff dff_A_kdVNOwJ95_2(.dout(w_dff_A_9dFVMJ195_2),.din(w_dff_A_kdVNOwJ95_2),.clk(gclk));
	jdff dff_A_jnql4Twp1_1(.dout(w_n839_0[1]),.din(w_dff_A_jnql4Twp1_1),.clk(gclk));
	jdff dff_A_Dz2EHSEq0_0(.dout(w_n574_3[0]),.din(w_dff_A_Dz2EHSEq0_0),.clk(gclk));
	jdff dff_A_zofU3MdX8_0(.dout(w_dff_A_Dz2EHSEq0_0),.din(w_dff_A_zofU3MdX8_0),.clk(gclk));
	jdff dff_A_NmVd0pp08_0(.dout(w_dff_A_zofU3MdX8_0),.din(w_dff_A_NmVd0pp08_0),.clk(gclk));
	jdff dff_A_m2v9p7Rr3_0(.dout(w_dff_A_NmVd0pp08_0),.din(w_dff_A_m2v9p7Rr3_0),.clk(gclk));
	jdff dff_A_a0n21v4d7_0(.dout(w_dff_A_m2v9p7Rr3_0),.din(w_dff_A_a0n21v4d7_0),.clk(gclk));
	jdff dff_A_KRynQWo53_0(.dout(w_dff_A_a0n21v4d7_0),.din(w_dff_A_KRynQWo53_0),.clk(gclk));
	jdff dff_A_vlFA9Oth2_0(.dout(w_dff_A_KRynQWo53_0),.din(w_dff_A_vlFA9Oth2_0),.clk(gclk));
	jdff dff_A_M5l0UahZ2_0(.dout(w_dff_A_vlFA9Oth2_0),.din(w_dff_A_M5l0UahZ2_0),.clk(gclk));
	jdff dff_A_IDNEl2ZS0_0(.dout(w_dff_A_M5l0UahZ2_0),.din(w_dff_A_IDNEl2ZS0_0),.clk(gclk));
	jdff dff_A_bD87Onbr9_0(.dout(w_dff_A_IDNEl2ZS0_0),.din(w_dff_A_bD87Onbr9_0),.clk(gclk));
	jdff dff_A_dAgqKiCL4_0(.dout(w_dff_A_bD87Onbr9_0),.din(w_dff_A_dAgqKiCL4_0),.clk(gclk));
	jdff dff_A_Mb1QoJJ16_0(.dout(w_dff_A_dAgqKiCL4_0),.din(w_dff_A_Mb1QoJJ16_0),.clk(gclk));
	jdff dff_A_XxpKgWzr6_1(.dout(w_n574_3[1]),.din(w_dff_A_XxpKgWzr6_1),.clk(gclk));
	jdff dff_A_qouqHV0E4_1(.dout(w_dff_A_XxpKgWzr6_1),.din(w_dff_A_qouqHV0E4_1),.clk(gclk));
	jdff dff_A_XJ1WFJjT2_1(.dout(w_dff_A_qouqHV0E4_1),.din(w_dff_A_XJ1WFJjT2_1),.clk(gclk));
	jdff dff_A_SAOtFZLC4_1(.dout(w_dff_A_XJ1WFJjT2_1),.din(w_dff_A_SAOtFZLC4_1),.clk(gclk));
	jdff dff_A_IQ4shD001_1(.dout(w_dff_A_SAOtFZLC4_1),.din(w_dff_A_IQ4shD001_1),.clk(gclk));
	jdff dff_A_nQyxS2Ra9_1(.dout(w_dff_A_IQ4shD001_1),.din(w_dff_A_nQyxS2Ra9_1),.clk(gclk));
	jdff dff_B_nuLMXo2V1_1(.din(n556),.dout(w_dff_B_nuLMXo2V1_1),.clk(gclk));
	jdff dff_B_8Xb02A4E5_1(.din(w_dff_B_nuLMXo2V1_1),.dout(w_dff_B_8Xb02A4E5_1),.clk(gclk));
	jdff dff_B_w0igAweX8_1(.din(w_dff_B_8Xb02A4E5_1),.dout(w_dff_B_w0igAweX8_1),.clk(gclk));
	jdff dff_B_m2KEuw7G7_1(.din(n256),.dout(w_dff_B_m2KEuw7G7_1),.clk(gclk));
	jdff dff_A_sOt7iCiN6_0(.dout(w_n335_0[0]),.din(w_dff_A_sOt7iCiN6_0),.clk(gclk));
	jdff dff_B_a9Bq9Jbt6_0(.din(n333),.dout(w_dff_B_a9Bq9Jbt6_0),.clk(gclk));
	jdff dff_B_92Xyjyt49_0(.din(w_dff_B_a9Bq9Jbt6_0),.dout(w_dff_B_92Xyjyt49_0),.clk(gclk));
	jdff dff_A_HP1SQecO2_0(.dout(w_n295_0[0]),.din(w_dff_A_HP1SQecO2_0),.clk(gclk));
	jdff dff_A_IrqUSM7k7_0(.dout(w_dff_A_HP1SQecO2_0),.din(w_dff_A_IrqUSM7k7_0),.clk(gclk));
	jdff dff_A_7LwcJ7e83_0(.dout(w_dff_A_IrqUSM7k7_0),.din(w_dff_A_7LwcJ7e83_0),.clk(gclk));
	jdff dff_A_uDBMBd6j5_0(.dout(w_dff_A_7LwcJ7e83_0),.din(w_dff_A_uDBMBd6j5_0),.clk(gclk));
	jdff dff_A_8ak2UWrj6_0(.dout(w_dff_A_uDBMBd6j5_0),.din(w_dff_A_8ak2UWrj6_0),.clk(gclk));
	jdff dff_B_weVp08Pp5_2(.din(n295),.dout(w_dff_B_weVp08Pp5_2),.clk(gclk));
	jdff dff_B_irG8Eo2N2_2(.din(w_dff_B_weVp08Pp5_2),.dout(w_dff_B_irG8Eo2N2_2),.clk(gclk));
	jdff dff_B_2sX8viCE6_1(.din(n288),.dout(w_dff_B_2sX8viCE6_1),.clk(gclk));
	jdff dff_B_K5kPQRym6_1(.din(n550),.dout(w_dff_B_K5kPQRym6_1),.clk(gclk));
	jdff dff_B_a3L0F4cM6_1(.din(w_dff_B_K5kPQRym6_1),.dout(w_dff_B_a3L0F4cM6_1),.clk(gclk));
	jdff dff_B_Xsx7zUaF5_1(.din(n551),.dout(w_dff_B_Xsx7zUaF5_1),.clk(gclk));
	jdff dff_B_jqYBxtNK9_1(.din(w_dff_B_Xsx7zUaF5_1),.dout(w_dff_B_jqYBxtNK9_1),.clk(gclk));
	jdff dff_B_WHMoBw497_1(.din(w_dff_B_jqYBxtNK9_1),.dout(w_dff_B_WHMoBw497_1),.clk(gclk));
	jdff dff_B_SW1uqonc9_0(.din(n552),.dout(w_dff_B_SW1uqonc9_0),.clk(gclk));
	jdff dff_A_u1iOwQ3o1_2(.dout(w_n541_1[2]),.din(w_dff_A_u1iOwQ3o1_2),.clk(gclk));
	jdff dff_A_7LZyPDqT9_1(.dout(w_n546_1[1]),.din(w_dff_A_7LZyPDqT9_1),.clk(gclk));
	jdff dff_A_ATjqoJSG6_1(.dout(w_dff_A_7LZyPDqT9_1),.din(w_dff_A_ATjqoJSG6_1),.clk(gclk));
	jdff dff_A_nKpt3kIN3_1(.dout(w_dff_A_ATjqoJSG6_1),.din(w_dff_A_nKpt3kIN3_1),.clk(gclk));
	jdff dff_A_OuUDbJ9h6_1(.dout(w_n531_3[1]),.din(w_dff_A_OuUDbJ9h6_1),.clk(gclk));
	jdff dff_A_iHzsrRMf2_1(.dout(w_dff_A_OuUDbJ9h6_1),.din(w_dff_A_iHzsrRMf2_1),.clk(gclk));
	jdff dff_A_dFeogwBV2_1(.dout(w_dff_A_iHzsrRMf2_1),.din(w_dff_A_dFeogwBV2_1),.clk(gclk));
	jdff dff_A_koRkDfe93_1(.dout(w_dff_A_dFeogwBV2_1),.din(w_dff_A_koRkDfe93_1),.clk(gclk));
	jdff dff_A_v45iXzmy9_1(.dout(w_dff_A_koRkDfe93_1),.din(w_dff_A_v45iXzmy9_1),.clk(gclk));
	jdff dff_A_DuVn1rsK2_1(.dout(w_dff_A_v45iXzmy9_1),.din(w_dff_A_DuVn1rsK2_1),.clk(gclk));
	jdff dff_A_qRSk5vFg3_1(.dout(w_dff_A_DuVn1rsK2_1),.din(w_dff_A_qRSk5vFg3_1),.clk(gclk));
	jdff dff_A_WWbyJ8n71_1(.dout(w_dff_A_qRSk5vFg3_1),.din(w_dff_A_WWbyJ8n71_1),.clk(gclk));
	jdff dff_A_HUiclmJB9_2(.dout(w_n531_3[2]),.din(w_dff_A_HUiclmJB9_2),.clk(gclk));
	jdff dff_A_Lqffpbav6_2(.dout(w_dff_A_HUiclmJB9_2),.din(w_dff_A_Lqffpbav6_2),.clk(gclk));
	jdff dff_A_TiiSdpQG7_2(.dout(w_dff_A_Lqffpbav6_2),.din(w_dff_A_TiiSdpQG7_2),.clk(gclk));
	jdff dff_A_YEyTH6s70_2(.dout(w_dff_A_TiiSdpQG7_2),.din(w_dff_A_YEyTH6s70_2),.clk(gclk));
	jdff dff_A_rFwZtK179_2(.dout(w_dff_A_YEyTH6s70_2),.din(w_dff_A_rFwZtK179_2),.clk(gclk));
	jdff dff_A_OOnSfLez6_2(.dout(w_dff_A_rFwZtK179_2),.din(w_dff_A_OOnSfLez6_2),.clk(gclk));
	jdff dff_A_aIFlGAtg5_2(.dout(w_dff_A_OOnSfLez6_2),.din(w_dff_A_aIFlGAtg5_2),.clk(gclk));
	jdff dff_A_0o0f1lf62_2(.dout(w_dff_A_aIFlGAtg5_2),.din(w_dff_A_0o0f1lf62_2),.clk(gclk));
	jdff dff_B_1BNxiPH74_1(.din(n492),.dout(w_dff_B_1BNxiPH74_1),.clk(gclk));
	jdff dff_B_zK9Y8eAx8_1(.din(w_dff_B_1BNxiPH74_1),.dout(w_dff_B_zK9Y8eAx8_1),.clk(gclk));
	jdff dff_B_PXQbvnM88_1(.din(w_dff_B_zK9Y8eAx8_1),.dout(w_dff_B_PXQbvnM88_1),.clk(gclk));
	jdff dff_A_kzR7u1TD1_1(.dout(w_n510_0[1]),.din(w_dff_A_kzR7u1TD1_1),.clk(gclk));
	jdff dff_B_yOM4cw0L7_1(.din(n508),.dout(w_dff_B_yOM4cw0L7_1),.clk(gclk));
	jdff dff_B_VxFm5xip0_0(.din(n504),.dout(w_dff_B_VxFm5xip0_0),.clk(gclk));
	jdff dff_A_2W7L7zYy3_0(.dout(w_n251_1[0]),.din(w_dff_A_2W7L7zYy3_0),.clk(gclk));
	jdff dff_A_rXfHdOZq3_0(.dout(w_dff_A_2W7L7zYy3_0),.din(w_dff_A_rXfHdOZq3_0),.clk(gclk));
	jdff dff_A_Lvok6WBq7_0(.dout(w_dff_A_rXfHdOZq3_0),.din(w_dff_A_Lvok6WBq7_0),.clk(gclk));
	jdff dff_A_7KWpzyRE0_1(.dout(w_G190_3[1]),.din(w_dff_A_7KWpzyRE0_1),.clk(gclk));
	jdff dff_A_0ZhmkXJ00_1(.dout(w_dff_A_7KWpzyRE0_1),.din(w_dff_A_0ZhmkXJ00_1),.clk(gclk));
	jdff dff_A_gWN7ECOm3_2(.dout(w_G190_3[2]),.din(w_dff_A_gWN7ECOm3_2),.clk(gclk));
	jdff dff_A_gmDsf9ec5_2(.dout(w_dff_A_gWN7ECOm3_2),.din(w_dff_A_gmDsf9ec5_2),.clk(gclk));
	jdff dff_A_kYJkszQe9_2(.dout(w_dff_A_gmDsf9ec5_2),.din(w_dff_A_kYJkszQe9_2),.clk(gclk));
	jdff dff_A_ex4bYEwq2_1(.dout(w_n501_0[1]),.din(w_dff_A_ex4bYEwq2_1),.clk(gclk));
	jdff dff_B_IOoAVviH4_2(.din(n501),.dout(w_dff_B_IOoAVviH4_2),.clk(gclk));
	jdff dff_B_MNhyYSQm0_0(.din(n500),.dout(w_dff_B_MNhyYSQm0_0),.clk(gclk));
	jdff dff_A_dpknuFx02_1(.dout(w_n497_0[1]),.din(w_dff_A_dpknuFx02_1),.clk(gclk));
	jdff dff_A_6nQF6u7s9_1(.dout(w_dff_A_dpknuFx02_1),.din(w_dff_A_6nQF6u7s9_1),.clk(gclk));
	jdff dff_A_nuUKsgjt7_0(.dout(w_n294_0[0]),.din(w_dff_A_nuUKsgjt7_0),.clk(gclk));
	jdff dff_A_bMVuxE5G0_0(.dout(w_dff_A_nuUKsgjt7_0),.din(w_dff_A_bMVuxE5G0_0),.clk(gclk));
	jdff dff_A_ZHa1CROU4_0(.dout(w_dff_A_bMVuxE5G0_0),.din(w_dff_A_ZHa1CROU4_0),.clk(gclk));
	jdff dff_A_GXpsoGnT9_0(.dout(w_dff_A_ZHa1CROU4_0),.din(w_dff_A_GXpsoGnT9_0),.clk(gclk));
	jdff dff_A_h3ncExe39_1(.dout(w_n292_0[1]),.din(w_dff_A_h3ncExe39_1),.clk(gclk));
	jdff dff_B_xlKVheb49_0(.din(n326),.dout(w_dff_B_xlKVheb49_0),.clk(gclk));
	jdff dff_A_WQyxfCM38_1(.dout(w_n175_1[1]),.din(w_dff_A_WQyxfCM38_1),.clk(gclk));
	jdff dff_A_DZ7VIiJY5_1(.dout(w_dff_A_WQyxfCM38_1),.din(w_dff_A_DZ7VIiJY5_1),.clk(gclk));
	jdff dff_A_s5KBHbYF5_1(.dout(w_dff_A_DZ7VIiJY5_1),.din(w_dff_A_s5KBHbYF5_1),.clk(gclk));
	jdff dff_A_t5mJqnh39_2(.dout(w_n175_1[2]),.din(w_dff_A_t5mJqnh39_2),.clk(gclk));
	jdff dff_A_F51UaCPE1_2(.dout(w_dff_A_t5mJqnh39_2),.din(w_dff_A_F51UaCPE1_2),.clk(gclk));
	jdff dff_A_Vt7nZ2km2_2(.dout(w_dff_A_F51UaCPE1_2),.din(w_dff_A_Vt7nZ2km2_2),.clk(gclk));
	jdff dff_A_efSbgbCQ2_1(.dout(w_n321_0[1]),.din(w_dff_A_efSbgbCQ2_1),.clk(gclk));
	jdff dff_B_bsd1qens3_2(.din(n321),.dout(w_dff_B_bsd1qens3_2),.clk(gclk));
	jdff dff_B_Fvc9IbLX9_2(.din(w_dff_B_bsd1qens3_2),.dout(w_dff_B_Fvc9IbLX9_2),.clk(gclk));
	jdff dff_A_Tg48kJFf3_0(.dout(w_n320_1[0]),.din(w_dff_A_Tg48kJFf3_0),.clk(gclk));
	jdff dff_A_GgI2SKKZ4_0(.dout(w_dff_A_Tg48kJFf3_0),.din(w_dff_A_GgI2SKKZ4_0),.clk(gclk));
	jdff dff_A_VYQW2B8n1_2(.dout(w_n320_0[2]),.din(w_dff_A_VYQW2B8n1_2),.clk(gclk));
	jdff dff_B_6hZTUKfw7_0(.din(n319),.dout(w_dff_B_6hZTUKfw7_0),.clk(gclk));
	jdff dff_A_mBQNp16G1_1(.dout(w_n312_0[1]),.din(w_dff_A_mBQNp16G1_1),.clk(gclk));
	jdff dff_A_qI8LMykU9_0(.dout(w_n309_0[0]),.din(w_dff_A_qI8LMykU9_0),.clk(gclk));
	jdff dff_A_Ivahdf7R9_1(.dout(w_G20_4[1]),.din(w_dff_A_Ivahdf7R9_1),.clk(gclk));
	jdff dff_A_NyYRzj6E9_1(.dout(w_n307_0[1]),.din(w_dff_A_NyYRzj6E9_1),.clk(gclk));
	jdff dff_A_1NcBMjnV7_1(.dout(w_dff_A_NyYRzj6E9_1),.din(w_dff_A_1NcBMjnV7_1),.clk(gclk));
	jdff dff_B_BZ4DsGxm4_0(.din(n305),.dout(w_dff_B_BZ4DsGxm4_0),.clk(gclk));
	jdff dff_A_Rc1cOJEn9_0(.dout(w_n301_0[0]),.din(w_dff_A_Rc1cOJEn9_0),.clk(gclk));
	jdff dff_B_Su4cP8Us5_0(.din(n300),.dout(w_dff_B_Su4cP8Us5_0),.clk(gclk));
	jdff dff_A_xdO5RVy33_0(.dout(w_G244_1[0]),.din(w_dff_A_xdO5RVy33_0),.clk(gclk));
	jdff dff_A_SLgBHqgl5_1(.dout(w_n298_0[1]),.din(w_dff_A_SLgBHqgl5_1),.clk(gclk));
	jdff dff_B_qdGSDyRC3_1(.din(n489),.dout(w_dff_B_qdGSDyRC3_1),.clk(gclk));
	jdff dff_A_Jq39jHdr6_0(.dout(w_n285_0[0]),.din(w_dff_A_Jq39jHdr6_0),.clk(gclk));
	jdff dff_A_4ZkRuOox8_0(.dout(w_dff_A_Jq39jHdr6_0),.din(w_dff_A_4ZkRuOox8_0),.clk(gclk));
	jdff dff_A_Jb85nn0H4_2(.dout(w_n283_0[2]),.din(w_dff_A_Jb85nn0H4_2),.clk(gclk));
	jdff dff_B_NMpI85nN2_1(.din(n270),.dout(w_dff_B_NMpI85nN2_1),.clk(gclk));
	jdff dff_B_lLNwMGRH2_0(.din(n281),.dout(w_dff_B_lLNwMGRH2_0),.clk(gclk));
	jdff dff_B_yxtZg7tQ0_0(.din(w_dff_B_lLNwMGRH2_0),.dout(w_dff_B_yxtZg7tQ0_0),.clk(gclk));
	jdff dff_B_EiP3ThKA5_0(.din(n279),.dout(w_dff_B_EiP3ThKA5_0),.clk(gclk));
	jdff dff_B_52PmUoso1_0(.din(w_dff_B_EiP3ThKA5_0),.dout(w_dff_B_52PmUoso1_0),.clk(gclk));
	jdff dff_A_2YVx9pA02_0(.dout(w_G68_4[0]),.din(w_dff_A_2YVx9pA02_0),.clk(gclk));
	jdff dff_A_3qsiCGA71_0(.dout(w_dff_A_2YVx9pA02_0),.din(w_dff_A_3qsiCGA71_0),.clk(gclk));
	jdff dff_A_GoKqyPRw1_2(.dout(w_G68_4[2]),.din(w_dff_A_GoKqyPRw1_2),.clk(gclk));
	jdff dff_A_ak5WnuVE9_0(.dout(w_n275_0[0]),.din(w_dff_A_ak5WnuVE9_0),.clk(gclk));
	jdff dff_B_ak8NJgpB3_2(.din(n275),.dout(w_dff_B_ak8NJgpB3_2),.clk(gclk));
	jdff dff_B_vu9Wbdxq9_1(.din(n261),.dout(w_dff_B_vu9Wbdxq9_1),.clk(gclk));
	jdff dff_B_nOF57Ihc9_0(.din(n264),.dout(w_dff_B_nOF57Ihc9_0),.clk(gclk));
	jdff dff_A_7yVOR6bZ8_1(.dout(w_n167_2[1]),.din(w_dff_A_7yVOR6bZ8_1),.clk(gclk));
	jdff dff_A_Z4RwFHax0_2(.dout(w_n167_2[2]),.din(w_dff_A_Z4RwFHax0_2),.clk(gclk));
	jdff dff_A_1pEbSX8l2_0(.dout(w_G238_1[0]),.din(w_dff_A_1pEbSX8l2_0),.clk(gclk));
	jdff dff_A_ER2hJ8O59_0(.dout(w_dff_A_1pEbSX8l2_0),.din(w_dff_A_ER2hJ8O59_0),.clk(gclk));
	jdff dff_A_n87Vl5Io4_1(.dout(w_G238_0[1]),.din(w_dff_A_n87Vl5Io4_1),.clk(gclk));
	jdff dff_A_6dK1w0MQ3_1(.dout(w_dff_A_n87Vl5Io4_1),.din(w_dff_A_6dK1w0MQ3_1),.clk(gclk));
	jdff dff_A_B6Vs1lec3_1(.dout(w_dff_A_6dK1w0MQ3_1),.din(w_dff_A_B6Vs1lec3_1),.clk(gclk));
	jdff dff_A_deBmJCFF2_2(.dout(w_G238_0[2]),.din(w_dff_A_deBmJCFF2_2),.clk(gclk));
	jdff dff_A_zd486uqH3_2(.dout(w_dff_A_deBmJCFF2_2),.din(w_dff_A_zd486uqH3_2),.clk(gclk));
	jdff dff_A_3hxgHbCD4_1(.dout(w_G244_0[1]),.din(w_dff_A_3hxgHbCD4_1),.clk(gclk));
	jdff dff_A_hh55e6nh0_1(.dout(w_dff_A_3hxgHbCD4_1),.din(w_dff_A_hh55e6nh0_1),.clk(gclk));
	jdff dff_A_5F61E4JD0_1(.dout(w_dff_A_hh55e6nh0_1),.din(w_dff_A_5F61E4JD0_1),.clk(gclk));
	jdff dff_A_KjkG0oBM0_2(.dout(w_G244_0[2]),.din(w_dff_A_KjkG0oBM0_2),.clk(gclk));
	jdff dff_A_agEXFetD7_2(.dout(w_dff_A_KjkG0oBM0_2),.din(w_dff_A_agEXFetD7_2),.clk(gclk));
	jdff dff_A_et9S8n2w5_0(.dout(w_n825_0[0]),.din(w_dff_A_et9S8n2w5_0),.clk(gclk));
	jdff dff_A_au7JGJKz5_0(.dout(w_dff_A_et9S8n2w5_0),.din(w_dff_A_au7JGJKz5_0),.clk(gclk));
	jdff dff_A_nyLEkgiy9_0(.dout(w_dff_A_au7JGJKz5_0),.din(w_dff_A_nyLEkgiy9_0),.clk(gclk));
	jdff dff_B_RTHaLB9P4_2(.din(n825),.dout(w_dff_B_RTHaLB9P4_2),.clk(gclk));
	jdff dff_A_USzALghU5_0(.dout(w_n824_0[0]),.din(w_dff_A_USzALghU5_0),.clk(gclk));
	jdff dff_A_TDDQKBda6_0(.dout(w_dff_A_USzALghU5_0),.din(w_dff_A_TDDQKBda6_0),.clk(gclk));
	jdff dff_A_zupOeHI68_0(.dout(w_dff_A_TDDQKBda6_0),.din(w_dff_A_zupOeHI68_0),.clk(gclk));
	jdff dff_A_pFE1Frdz6_0(.dout(w_dff_A_zupOeHI68_0),.din(w_dff_A_pFE1Frdz6_0),.clk(gclk));
	jdff dff_A_OppAy5Zf5_0(.dout(w_dff_A_pFE1Frdz6_0),.din(w_dff_A_OppAy5Zf5_0),.clk(gclk));
	jdff dff_A_XN6l2aJN6_1(.dout(w_n824_0[1]),.din(w_dff_A_XN6l2aJN6_1),.clk(gclk));
	jdff dff_A_S99EpfW01_1(.dout(w_dff_A_XN6l2aJN6_1),.din(w_dff_A_S99EpfW01_1),.clk(gclk));
	jdff dff_A_Y5gNh7m69_1(.dout(w_dff_A_S99EpfW01_1),.din(w_dff_A_Y5gNh7m69_1),.clk(gclk));
	jdff dff_B_zkwCK5Dw6_0(.din(n823),.dout(w_dff_B_zkwCK5Dw6_0),.clk(gclk));
	jdff dff_A_IgTa6ZNf1_1(.dout(w_n819_0[1]),.din(w_dff_A_IgTa6ZNf1_1),.clk(gclk));
	jdff dff_A_sqJjZZ9z9_0(.dout(w_n541_0[0]),.din(w_dff_A_sqJjZZ9z9_0),.clk(gclk));
	jdff dff_A_ghJ8wUVE0_2(.dout(w_n541_0[2]),.din(w_dff_A_ghJ8wUVE0_2),.clk(gclk));
	jdff dff_A_HN76owjW0_2(.dout(w_dff_A_ghJ8wUVE0_2),.din(w_dff_A_HN76owjW0_2),.clk(gclk));
	jdff dff_A_2xUdHjSB5_2(.dout(w_dff_A_HN76owjW0_2),.din(w_dff_A_2xUdHjSB5_2),.clk(gclk));
	jdff dff_A_f28f5INd7_2(.dout(w_dff_A_2xUdHjSB5_2),.din(w_dff_A_f28f5INd7_2),.clk(gclk));
	jdff dff_B_w13kkr5n3_3(.din(n541),.dout(w_dff_B_w13kkr5n3_3),.clk(gclk));
	jdff dff_B_DuujXMuX4_3(.din(w_dff_B_w13kkr5n3_3),.dout(w_dff_B_DuujXMuX4_3),.clk(gclk));
	jdff dff_B_6JNF1BfV2_3(.din(w_dff_B_DuujXMuX4_3),.dout(w_dff_B_6JNF1BfV2_3),.clk(gclk));
	jdff dff_B_mQ5ZAuB85_3(.din(w_dff_B_6JNF1BfV2_3),.dout(w_dff_B_mQ5ZAuB85_3),.clk(gclk));
	jdff dff_A_8lR3zUvc4_1(.dout(w_n760_0[1]),.din(w_dff_A_8lR3zUvc4_1),.clk(gclk));
	jdff dff_A_W7gmO0gB4_1(.dout(w_dff_A_8lR3zUvc4_1),.din(w_dff_A_W7gmO0gB4_1),.clk(gclk));
	jdff dff_A_prKTJLcj5_1(.dout(w_dff_A_W7gmO0gB4_1),.din(w_dff_A_prKTJLcj5_1),.clk(gclk));
	jdff dff_A_6IsqXu5a7_2(.dout(w_n538_0[2]),.din(w_dff_A_6IsqXu5a7_2),.clk(gclk));
	jdff dff_A_dK2rfGwR3_2(.dout(w_dff_A_6IsqXu5a7_2),.din(w_dff_A_dK2rfGwR3_2),.clk(gclk));
	jdff dff_B_s1MZ71WS2_0(.din(n536),.dout(w_dff_B_s1MZ71WS2_0),.clk(gclk));
	jdff dff_B_Sc8WFc9M4_0(.din(w_dff_B_s1MZ71WS2_0),.dout(w_dff_B_Sc8WFc9M4_0),.clk(gclk));
	jdff dff_B_witi1zg83_0(.din(w_dff_B_Sc8WFc9M4_0),.dout(w_dff_B_witi1zg83_0),.clk(gclk));
	jdff dff_B_MMoY9aKr6_0(.din(w_dff_B_witi1zg83_0),.dout(w_dff_B_MMoY9aKr6_0),.clk(gclk));
	jdff dff_A_nnK8K6Yd5_1(.dout(w_n255_0[1]),.din(w_dff_A_nnK8K6Yd5_1),.clk(gclk));
	jdff dff_A_jEkaSazK0_1(.dout(w_dff_A_nnK8K6Yd5_1),.din(w_dff_A_jEkaSazK0_1),.clk(gclk));
	jdff dff_B_OlWs8Heb2_0(.din(n253),.dout(w_dff_B_OlWs8Heb2_0),.clk(gclk));
	jdff dff_A_Y6eoVmlR8_1(.dout(w_n251_2[1]),.din(w_dff_A_Y6eoVmlR8_1),.clk(gclk));
	jdff dff_A_WgCxRYDW1_1(.dout(w_dff_A_Y6eoVmlR8_1),.din(w_dff_A_WgCxRYDW1_1),.clk(gclk));
	jdff dff_A_vUBv06Fc3_2(.dout(w_n251_2[2]),.din(w_dff_A_vUBv06Fc3_2),.clk(gclk));
	jdff dff_A_RfNyO60m7_0(.dout(w_n246_0[0]),.din(w_dff_A_RfNyO60m7_0),.clk(gclk));
	jdff dff_A_2kHRESU46_0(.dout(w_dff_A_RfNyO60m7_0),.din(w_dff_A_2kHRESU46_0),.clk(gclk));
	jdff dff_A_9jfPiPj04_2(.dout(w_n246_0[2]),.din(w_dff_A_9jfPiPj04_2),.clk(gclk));
	jdff dff_A_GsXmotwF4_2(.dout(w_dff_A_9jfPiPj04_2),.din(w_dff_A_GsXmotwF4_2),.clk(gclk));
	jdff dff_B_QtalDuBA3_0(.din(n245),.dout(w_dff_B_QtalDuBA3_0),.clk(gclk));
	jdff dff_A_5cPOZy7q5_0(.dout(w_n243_0[0]),.din(w_dff_A_5cPOZy7q5_0),.clk(gclk));
	jdff dff_B_K7Pdc8mo9_1(.din(n227),.dout(w_dff_B_K7Pdc8mo9_1),.clk(gclk));
	jdff dff_A_ZvC7meZE3_1(.dout(w_G87_3[1]),.din(w_dff_A_ZvC7meZE3_1),.clk(gclk));
	jdff dff_A_hzv3AJbH0_1(.dout(w_dff_A_ZvC7meZE3_1),.din(w_dff_A_hzv3AJbH0_1),.clk(gclk));
	jdff dff_A_Z9sZP4ti6_1(.dout(w_dff_A_hzv3AJbH0_1),.din(w_dff_A_Z9sZP4ti6_1),.clk(gclk));
	jdff dff_A_K5fo6cxL0_1(.dout(w_dff_A_Z9sZP4ti6_1),.din(w_dff_A_K5fo6cxL0_1),.clk(gclk));
	jdff dff_A_aAnbTL744_2(.dout(w_G87_3[2]),.din(w_dff_A_aAnbTL744_2),.clk(gclk));
	jdff dff_A_SPflITre2_0(.dout(w_n228_0[0]),.din(w_dff_A_SPflITre2_0),.clk(gclk));
	jdff dff_B_IluYWD2B6_2(.din(n228),.dout(w_dff_B_IluYWD2B6_2),.clk(gclk));
	jdff dff_A_bERrxIDg1_0(.dout(w_G20_5[0]),.din(w_dff_A_bERrxIDg1_0),.clk(gclk));
	jdff dff_A_zXkfapMO8_1(.dout(w_G20_5[1]),.din(w_dff_A_zXkfapMO8_1),.clk(gclk));
	jdff dff_A_iXH7P5d46_1(.dout(w_dff_A_zXkfapMO8_1),.din(w_dff_A_iXH7P5d46_1),.clk(gclk));
	jdff dff_A_tGIwWPc98_0(.dout(w_n223_0[0]),.din(w_dff_A_tGIwWPc98_0),.clk(gclk));
	jdff dff_A_x836GCzJ0_0(.dout(w_dff_A_tGIwWPc98_0),.din(w_dff_A_x836GCzJ0_0),.clk(gclk));
	jdff dff_A_yLyYwaU37_0(.dout(w_n80_1[0]),.din(w_dff_A_yLyYwaU37_0),.clk(gclk));
	jdff dff_A_5AF34kqV1_2(.dout(w_n80_1[2]),.din(w_dff_A_5AF34kqV1_2),.clk(gclk));
	jdff dff_A_54pfsnNL9_2(.dout(w_dff_A_5AF34kqV1_2),.din(w_dff_A_54pfsnNL9_2),.clk(gclk));
	jdff dff_B_Bas7vXo25_1(.din(n213),.dout(w_dff_B_Bas7vXo25_1),.clk(gclk));
	jdff dff_B_oLqY92ZG7_1(.din(w_dff_B_Bas7vXo25_1),.dout(w_dff_B_oLqY92ZG7_1),.clk(gclk));
	jdff dff_B_WafiYv6g5_0(.din(n216),.dout(w_dff_B_WafiYv6g5_0),.clk(gclk));
	jdff dff_A_Xkk2p6Kp8_2(.dout(w_n83_0[2]),.din(w_dff_A_Xkk2p6Kp8_2),.clk(gclk));
	jdff dff_A_oTrsiTn54_0(.dout(w_G250_1[0]),.din(w_dff_A_oTrsiTn54_0),.clk(gclk));
	jdff dff_A_4itEZmO81_0(.dout(w_dff_A_oTrsiTn54_0),.din(w_dff_A_4itEZmO81_0),.clk(gclk));
	jdff dff_A_8SbsIMPh6_1(.dout(w_G250_0[1]),.din(w_dff_A_8SbsIMPh6_1),.clk(gclk));
	jdff dff_A_EnmipDdM3_1(.dout(w_dff_A_8SbsIMPh6_1),.din(w_dff_A_EnmipDdM3_1),.clk(gclk));
	jdff dff_A_yuQOSCFe1_2(.dout(w_G250_0[2]),.din(w_dff_A_yuQOSCFe1_2),.clk(gclk));
	jdff dff_A_It1b8Apm1_2(.dout(w_dff_A_yuQOSCFe1_2),.din(w_dff_A_It1b8Apm1_2),.clk(gclk));
	jdff dff_A_NYiak4bQ0_2(.dout(w_dff_A_It1b8Apm1_2),.din(w_dff_A_NYiak4bQ0_2),.clk(gclk));
	jdff dff_A_d4neQDxl2_0(.dout(w_n214_0[0]),.din(w_dff_A_d4neQDxl2_0),.clk(gclk));
	jdff dff_A_Mguwjh3Y5_0(.dout(w_dff_A_d4neQDxl2_0),.din(w_dff_A_Mguwjh3Y5_0),.clk(gclk));
	jdff dff_A_xPlFSzND5_0(.dout(w_n175_2[0]),.din(w_dff_A_xPlFSzND5_0),.clk(gclk));
	jdff dff_A_J8Xrpnru1_0(.dout(w_dff_A_xPlFSzND5_0),.din(w_dff_A_J8Xrpnru1_0),.clk(gclk));
	jdff dff_A_MfTlVsaB8_2(.dout(w_n175_2[2]),.din(w_dff_A_MfTlVsaB8_2),.clk(gclk));
	jdff dff_A_8sSiV2zs4_1(.dout(w_n210_0[1]),.din(w_dff_A_8sSiV2zs4_1),.clk(gclk));
	jdff dff_A_GzGL9BU06_1(.dout(w_dff_A_8sSiV2zs4_1),.din(w_dff_A_GzGL9BU06_1),.clk(gclk));
	jdff dff_A_6ynn85cg3_1(.dout(w_n85_0[1]),.din(w_dff_A_6ynn85cg3_1),.clk(gclk));
	jdff dff_A_3raSrlKE7_1(.dout(w_dff_A_6ynn85cg3_1),.din(w_dff_A_3raSrlKE7_1),.clk(gclk));
	jdff dff_A_NingPJJr5_0(.dout(w_G396_0[0]),.din(w_dff_A_NingPJJr5_0),.clk(gclk));
	jdff dff_A_FrefPK8O5_0(.dout(w_dff_A_NingPJJr5_0),.din(w_dff_A_FrefPK8O5_0),.clk(gclk));
	jdff dff_A_THdACRsx7_0(.dout(w_dff_A_FrefPK8O5_0),.din(w_dff_A_THdACRsx7_0),.clk(gclk));
	jdff dff_A_zihQz6gZ9_0(.dout(w_dff_A_THdACRsx7_0),.din(w_dff_A_zihQz6gZ9_0),.clk(gclk));
	jdff dff_A_5No72I6T6_0(.dout(w_dff_A_zihQz6gZ9_0),.din(w_dff_A_5No72I6T6_0),.clk(gclk));
	jdff dff_A_L227eugT4_0(.dout(w_dff_A_5No72I6T6_0),.din(w_dff_A_L227eugT4_0),.clk(gclk));
	jdff dff_A_8YmVFp8d9_2(.dout(G396),.din(w_dff_A_8YmVFp8d9_2),.clk(gclk));
	jdff dff_B_k3R0GRDO1_1(.din(n577),.dout(w_dff_B_k3R0GRDO1_1),.clk(gclk));
	jdff dff_B_9AtbX24Q1_0(.din(n653),.dout(w_dff_B_9AtbX24Q1_0),.clk(gclk));
	jdff dff_B_bqSrjtx16_0(.din(w_dff_B_9AtbX24Q1_0),.dout(w_dff_B_bqSrjtx16_0),.clk(gclk));
	jdff dff_B_aPDOq9fw2_0(.din(w_dff_B_bqSrjtx16_0),.dout(w_dff_B_aPDOq9fw2_0),.clk(gclk));
	jdff dff_B_tiVVBsFY0_1(.din(n635),.dout(w_dff_B_tiVVBsFY0_1),.clk(gclk));
	jdff dff_B_0vRxV8tn7_1(.din(w_dff_B_tiVVBsFY0_1),.dout(w_dff_B_0vRxV8tn7_1),.clk(gclk));
	jdff dff_B_zJLrF8qo5_1(.din(w_dff_B_0vRxV8tn7_1),.dout(w_dff_B_zJLrF8qo5_1),.clk(gclk));
	jdff dff_B_vNQOvYjL3_1(.din(w_dff_B_zJLrF8qo5_1),.dout(w_dff_B_vNQOvYjL3_1),.clk(gclk));
	jdff dff_B_BkPSlq8z9_0(.din(n649),.dout(w_dff_B_BkPSlq8z9_0),.clk(gclk));
	jdff dff_B_Y9mIcjJJ2_0(.din(w_dff_B_BkPSlq8z9_0),.dout(w_dff_B_Y9mIcjJJ2_0),.clk(gclk));
	jdff dff_A_9DOAq5WU0_0(.dout(w_n647_0[0]),.din(w_dff_A_9DOAq5WU0_0),.clk(gclk));
	jdff dff_A_Yp6EBFDp7_0(.dout(w_G355_0),.din(w_dff_A_Yp6EBFDp7_0),.clk(gclk));
	jdff dff_B_JxW6VFUK4_2(.din(G355_fa_),.dout(w_dff_B_JxW6VFUK4_2),.clk(gclk));
	jdff dff_A_ytxfUw0E9_2(.dout(w_n80_0[2]),.din(w_dff_A_ytxfUw0E9_2),.clk(gclk));
	jdff dff_A_p1wf4wwP0_2(.dout(w_dff_A_ytxfUw0E9_2),.din(w_dff_A_p1wf4wwP0_2),.clk(gclk));
	jdff dff_A_iMa7f0N08_2(.dout(w_dff_A_p1wf4wwP0_2),.din(w_dff_A_iMa7f0N08_2),.clk(gclk));
	jdff dff_A_Uxiv7mDf4_1(.dout(w_n79_0[1]),.din(w_dff_A_Uxiv7mDf4_1),.clk(gclk));
	jdff dff_A_KOPMjFeF6_1(.dout(w_dff_A_Uxiv7mDf4_1),.din(w_dff_A_KOPMjFeF6_1),.clk(gclk));
	jdff dff_A_DUwZdRKu2_1(.dout(w_n78_1[1]),.din(w_dff_A_DUwZdRKu2_1),.clk(gclk));
	jdff dff_A_ml3cqTxh8_1(.dout(w_n78_0[1]),.din(w_dff_A_ml3cqTxh8_1),.clk(gclk));
	jdff dff_A_sucufshR2_1(.dout(w_dff_A_ml3cqTxh8_1),.din(w_dff_A_sucufshR2_1),.clk(gclk));
	jdff dff_A_47GHoTMv4_1(.dout(w_G87_1[1]),.din(w_dff_A_47GHoTMv4_1),.clk(gclk));
	jdff dff_A_ERpOTMRg7_1(.dout(w_dff_A_47GHoTMv4_1),.din(w_dff_A_ERpOTMRg7_1),.clk(gclk));
	jdff dff_A_YZd3ftvQ7_1(.dout(w_dff_A_ERpOTMRg7_1),.din(w_dff_A_YZd3ftvQ7_1),.clk(gclk));
	jdff dff_A_AosIMfix1_2(.dout(w_G87_1[2]),.din(w_dff_A_AosIMfix1_2),.clk(gclk));
	jdff dff_A_lt8TWJel9_2(.dout(w_dff_A_AosIMfix1_2),.din(w_dff_A_lt8TWJel9_2),.clk(gclk));
	jdff dff_A_vEhoGedL2_2(.dout(w_dff_A_lt8TWJel9_2),.din(w_dff_A_vEhoGedL2_2),.clk(gclk));
	jdff dff_B_3ZrYfTLl2_1(.din(n638),.dout(w_dff_B_3ZrYfTLl2_1),.clk(gclk));
	jdff dff_B_7cKiESw98_1(.din(w_dff_B_3ZrYfTLl2_1),.dout(w_dff_B_7cKiESw98_1),.clk(gclk));
	jdff dff_B_coLmqX0w8_1(.din(w_dff_B_7cKiESw98_1),.dout(w_dff_B_coLmqX0w8_1),.clk(gclk));
	jdff dff_B_3i0omfmu0_1(.din(w_dff_B_coLmqX0w8_1),.dout(w_dff_B_3i0omfmu0_1),.clk(gclk));
	jdff dff_B_EJaLm2yo5_0(.din(n641),.dout(w_dff_B_EJaLm2yo5_0),.clk(gclk));
	jdff dff_B_Cv0jdZhY0_0(.din(w_dff_B_EJaLm2yo5_0),.dout(w_dff_B_Cv0jdZhY0_0),.clk(gclk));
	jdff dff_B_frWjfpCC8_0(.din(w_dff_B_Cv0jdZhY0_0),.dout(w_dff_B_frWjfpCC8_0),.clk(gclk));
	jdff dff_A_HGiHmRHa9_1(.dout(w_n92_0[1]),.din(w_dff_A_HGiHmRHa9_1),.clk(gclk));
	jdff dff_A_YssGkI0D9_1(.dout(w_dff_A_HGiHmRHa9_1),.din(w_dff_A_YssGkI0D9_1),.clk(gclk));
	jdff dff_A_Q6r6O0Ff9_1(.dout(w_dff_A_YssGkI0D9_1),.din(w_dff_A_Q6r6O0Ff9_1),.clk(gclk));
	jdff dff_A_q76h1Grp0_1(.dout(w_n135_0[1]),.din(w_dff_A_q76h1Grp0_1),.clk(gclk));
	jdff dff_A_ZNWPlGT61_0(.dout(w_G77_4[0]),.din(w_dff_A_ZNWPlGT61_0),.clk(gclk));
	jdff dff_A_L324XXoF0_1(.dout(w_G77_1[1]),.din(w_dff_A_L324XXoF0_1),.clk(gclk));
	jdff dff_A_wDEjfRe06_1(.dout(w_dff_A_L324XXoF0_1),.din(w_dff_A_wDEjfRe06_1),.clk(gclk));
	jdff dff_A_nLvSUpGX2_1(.dout(w_dff_A_wDEjfRe06_1),.din(w_dff_A_nLvSUpGX2_1),.clk(gclk));
	jdff dff_A_6zURVSFX1_2(.dout(w_G68_1[2]),.din(w_dff_A_6zURVSFX1_2),.clk(gclk));
	jdff dff_A_BuFQ7ENo7_2(.dout(w_dff_A_6zURVSFX1_2),.din(w_dff_A_BuFQ7ENo7_2),.clk(gclk));
	jdff dff_A_NtRs0Lns7_2(.dout(w_dff_A_BuFQ7ENo7_2),.din(w_dff_A_NtRs0Lns7_2),.clk(gclk));
	jdff dff_A_ZUAPrBEK6_0(.dout(w_G50_5[0]),.din(w_dff_A_ZUAPrBEK6_0),.clk(gclk));
	jdff dff_A_b9GROpJW2_0(.dout(w_dff_A_ZUAPrBEK6_0),.din(w_dff_A_b9GROpJW2_0),.clk(gclk));
	jdff dff_A_G2slVSIU2_1(.dout(w_G50_5[1]),.din(w_dff_A_G2slVSIU2_1),.clk(gclk));
	jdff dff_A_O14BRBRi1_0(.dout(w_n339_1[0]),.din(w_dff_A_O14BRBRi1_0),.clk(gclk));
	jdff dff_A_4Ip61xn62_1(.dout(w_n339_0[1]),.din(w_dff_A_4Ip61xn62_1),.clk(gclk));
	jdff dff_A_P2k1ZYb97_1(.dout(w_dff_A_4Ip61xn62_1),.din(w_dff_A_P2k1ZYb97_1),.clk(gclk));
	jdff dff_A_VcM5NMVd3_1(.dout(w_dff_A_P2k1ZYb97_1),.din(w_dff_A_VcM5NMVd3_1),.clk(gclk));
	jdff dff_A_9mcLTUWd1_1(.dout(w_dff_A_VcM5NMVd3_1),.din(w_dff_A_9mcLTUWd1_1),.clk(gclk));
	jdff dff_A_8wdWQmrJ2_1(.dout(w_n637_0[1]),.din(w_dff_A_8wdWQmrJ2_1),.clk(gclk));
	jdff dff_A_x3cqZVrK0_1(.dout(w_dff_A_8wdWQmrJ2_1),.din(w_dff_A_x3cqZVrK0_1),.clk(gclk));
	jdff dff_A_mwQXrT2J4_1(.dout(w_n634_4[1]),.din(w_dff_A_mwQXrT2J4_1),.clk(gclk));
	jdff dff_A_qC7rVrwi6_1(.dout(w_n634_1[1]),.din(w_dff_A_qC7rVrwi6_1),.clk(gclk));
	jdff dff_A_QqpC6r7Z8_2(.dout(w_n634_1[2]),.din(w_dff_A_QqpC6r7Z8_2),.clk(gclk));
	jdff dff_A_HH7vxqTT1_2(.dout(w_dff_A_QqpC6r7Z8_2),.din(w_dff_A_HH7vxqTT1_2),.clk(gclk));
	jdff dff_A_NpB3G7Bq5_0(.dout(w_n634_0[0]),.din(w_dff_A_NpB3G7Bq5_0),.clk(gclk));
	jdff dff_A_lavui2pd4_1(.dout(w_n634_0[1]),.din(w_dff_A_lavui2pd4_1),.clk(gclk));
	jdff dff_A_nZFqLcox7_1(.dout(w_dff_A_lavui2pd4_1),.din(w_dff_A_nZFqLcox7_1),.clk(gclk));
	jdff dff_A_qcS1sfZV7_0(.dout(w_n151_3[0]),.din(w_dff_A_qcS1sfZV7_0),.clk(gclk));
	jdff dff_A_AdIubfXa6_0(.dout(w_dff_A_qcS1sfZV7_0),.din(w_dff_A_AdIubfXa6_0),.clk(gclk));
	jdff dff_A_OO7uJMLQ3_2(.dout(w_n151_3[2]),.din(w_dff_A_OO7uJMLQ3_2),.clk(gclk));
	jdff dff_B_4Gh0fwtc9_2(.din(G326),.dout(w_dff_B_4Gh0fwtc9_2),.clk(gclk));
	jdff dff_B_856zJ3iP1_2(.din(w_dff_B_4Gh0fwtc9_2),.dout(w_dff_B_856zJ3iP1_2),.clk(gclk));
	jdff dff_B_C9KSGfsQ0_2(.din(w_dff_B_856zJ3iP1_2),.dout(w_dff_B_C9KSGfsQ0_2),.clk(gclk));
	jdff dff_B_EO90XBws6_3(.din(G317),.dout(w_dff_B_EO90XBws6_3),.clk(gclk));
	jdff dff_B_aWlbAKyW4_3(.din(w_dff_B_EO90XBws6_3),.dout(w_dff_B_aWlbAKyW4_3),.clk(gclk));
	jdff dff_B_pIQiSaGZ0_3(.din(w_dff_B_aWlbAKyW4_3),.dout(w_dff_B_pIQiSaGZ0_3),.clk(gclk));
	jdff dff_B_Ty1SYtPV1_3(.din(G322),.dout(w_dff_B_Ty1SYtPV1_3),.clk(gclk));
	jdff dff_B_mXNucLYp9_3(.din(w_dff_B_Ty1SYtPV1_3),.dout(w_dff_B_mXNucLYp9_3),.clk(gclk));
	jdff dff_B_Pa74sO4r2_3(.din(w_dff_B_mXNucLYp9_3),.dout(w_dff_B_Pa74sO4r2_3),.clk(gclk));
	jdff dff_B_Zcm9hBc21_1(.din(G329),.dout(w_dff_B_Zcm9hBc21_1),.clk(gclk));
	jdff dff_B_JVJHfrUM2_1(.din(w_dff_B_Zcm9hBc21_1),.dout(w_dff_B_JVJHfrUM2_1),.clk(gclk));
	jdff dff_B_GXaL3ZsG0_1(.din(w_dff_B_JVJHfrUM2_1),.dout(w_dff_B_GXaL3ZsG0_1),.clk(gclk));
	jdff dff_A_g0CTxuN66_0(.dout(w_G294_3[0]),.din(w_dff_A_g0CTxuN66_0),.clk(gclk));
	jdff dff_A_WkIZ9Ipi3_0(.dout(w_dff_A_g0CTxuN66_0),.din(w_dff_A_WkIZ9Ipi3_0),.clk(gclk));
	jdff dff_A_QktPgrCA7_0(.dout(w_dff_A_WkIZ9Ipi3_0),.din(w_dff_A_QktPgrCA7_0),.clk(gclk));
	jdff dff_A_35I4PX3a1_0(.dout(w_G294_0[0]),.din(w_dff_A_35I4PX3a1_0),.clk(gclk));
	jdff dff_A_LjQXjsAQ4_0(.dout(w_dff_A_35I4PX3a1_0),.din(w_dff_A_LjQXjsAQ4_0),.clk(gclk));
	jdff dff_A_g8b3qWfZ8_0(.dout(w_dff_A_LjQXjsAQ4_0),.din(w_dff_A_g8b3qWfZ8_0),.clk(gclk));
	jdff dff_A_b02XpM220_1(.dout(w_G294_0[1]),.din(w_dff_A_b02XpM220_1),.clk(gclk));
	jdff dff_A_ZvST1GIK2_1(.dout(w_dff_A_b02XpM220_1),.din(w_dff_A_ZvST1GIK2_1),.clk(gclk));
	jdff dff_A_qeqK6uzc8_1(.dout(w_dff_A_ZvST1GIK2_1),.din(w_dff_A_qeqK6uzc8_1),.clk(gclk));
	jdff dff_B_5lXSsvLL5_3(.din(G311),.dout(w_dff_B_5lXSsvLL5_3),.clk(gclk));
	jdff dff_B_JUdPVsRX7_3(.din(w_dff_B_5lXSsvLL5_3),.dout(w_dff_B_JUdPVsRX7_3),.clk(gclk));
	jdff dff_B_kZ0fZPgi3_3(.din(w_dff_B_JUdPVsRX7_3),.dout(w_dff_B_kZ0fZPgi3_3),.clk(gclk));
	jdff dff_A_OqvBEi9O5_0(.dout(w_G77_3[0]),.din(w_dff_A_OqvBEi9O5_0),.clk(gclk));
	jdff dff_A_EDjJCaEM3_0(.dout(w_dff_A_OqvBEi9O5_0),.din(w_dff_A_EDjJCaEM3_0),.clk(gclk));
	jdff dff_A_9xqjFTvx0_0(.dout(w_dff_A_EDjJCaEM3_0),.din(w_dff_A_9xqjFTvx0_0),.clk(gclk));
	jdff dff_A_6QIZpNEc4_2(.dout(w_G77_3[2]),.din(w_dff_A_6QIZpNEc4_2),.clk(gclk));
	jdff dff_A_hMiY208a9_2(.dout(w_dff_A_6QIZpNEc4_2),.din(w_dff_A_hMiY208a9_2),.clk(gclk));
	jdff dff_A_iUBzaUNc4_2(.dout(w_dff_A_hMiY208a9_2),.din(w_dff_A_iUBzaUNc4_2),.clk(gclk));
	jdff dff_A_5hCaIDoL6_1(.dout(w_G77_0[1]),.din(w_dff_A_5hCaIDoL6_1),.clk(gclk));
	jdff dff_A_WW8we5c08_0(.dout(w_G97_3[0]),.din(w_dff_A_WW8we5c08_0),.clk(gclk));
	jdff dff_A_Npus9YKO8_0(.dout(w_dff_A_WW8we5c08_0),.din(w_dff_A_Npus9YKO8_0),.clk(gclk));
	jdff dff_A_FhAe9Zg75_0(.dout(w_dff_A_Npus9YKO8_0),.din(w_dff_A_FhAe9Zg75_0),.clk(gclk));
	jdff dff_A_cuGTOmQg6_1(.dout(w_G97_3[1]),.din(w_dff_A_cuGTOmQg6_1),.clk(gclk));
	jdff dff_A_Oa27SE9W4_1(.dout(w_dff_A_cuGTOmQg6_1),.din(w_dff_A_Oa27SE9W4_1),.clk(gclk));
	jdff dff_A_fXEdsmQ75_1(.dout(w_dff_A_Oa27SE9W4_1),.din(w_dff_A_fXEdsmQ75_1),.clk(gclk));
	jdff dff_A_iKTNXKZc3_0(.dout(w_n601_0[0]),.din(w_dff_A_iKTNXKZc3_0),.clk(gclk));
	jdff dff_A_tikgggIb4_0(.dout(w_G159_3[0]),.din(w_dff_A_tikgggIb4_0),.clk(gclk));
	jdff dff_A_69Qogbok1_1(.dout(w_G159_3[1]),.din(w_dff_A_69Qogbok1_1),.clk(gclk));
	jdff dff_A_uCZnG92N2_0(.dout(w_G159_0[0]),.din(w_dff_A_uCZnG92N2_0),.clk(gclk));
	jdff dff_A_ynTVZFdy6_1(.dout(w_G159_0[1]),.din(w_dff_A_ynTVZFdy6_1),.clk(gclk));
	jdff dff_B_8VStsy0h7_3(.din(G159),.dout(w_dff_B_8VStsy0h7_3),.clk(gclk));
	jdff dff_B_6tq39FvZ8_3(.din(w_dff_B_8VStsy0h7_3),.dout(w_dff_B_6tq39FvZ8_3),.clk(gclk));
	jdff dff_A_VWmwSnvD7_0(.dout(w_n251_0[0]),.din(w_dff_A_VWmwSnvD7_0),.clk(gclk));
	jdff dff_A_d4tngxdW3_0(.dout(w_dff_A_VWmwSnvD7_0),.din(w_dff_A_d4tngxdW3_0),.clk(gclk));
	jdff dff_A_LSZJC3xa5_0(.dout(w_dff_A_d4tngxdW3_0),.din(w_dff_A_LSZJC3xa5_0),.clk(gclk));
	jdff dff_A_0WdZJnEe2_0(.dout(w_dff_A_LSZJC3xa5_0),.din(w_dff_A_0WdZJnEe2_0),.clk(gclk));
	jdff dff_A_fXfdB0lU2_1(.dout(w_n251_0[1]),.din(w_dff_A_fXfdB0lU2_1),.clk(gclk));
	jdff dff_A_9mtb9rSS4_1(.dout(w_dff_A_fXfdB0lU2_1),.din(w_dff_A_9mtb9rSS4_1),.clk(gclk));
	jdff dff_A_yQd0I7028_1(.dout(w_dff_A_9mtb9rSS4_1),.din(w_dff_A_yQd0I7028_1),.clk(gclk));
	jdff dff_A_ZOM03yNy5_1(.dout(w_dff_A_yQd0I7028_1),.din(w_dff_A_ZOM03yNy5_1),.clk(gclk));
	jdff dff_A_iNETUz0D5_0(.dout(w_G58_4[0]),.din(w_dff_A_iNETUz0D5_0),.clk(gclk));
	jdff dff_A_NqtSGlXd4_1(.dout(w_G58_4[1]),.din(w_dff_A_NqtSGlXd4_1),.clk(gclk));
	jdff dff_A_mESEmxt54_0(.dout(w_G58_1[0]),.din(w_dff_A_mESEmxt54_0),.clk(gclk));
	jdff dff_A_T0huWdzQ2_0(.dout(w_dff_A_mESEmxt54_0),.din(w_dff_A_T0huWdzQ2_0),.clk(gclk));
	jdff dff_A_k3uNQ6l93_1(.dout(w_G58_0[1]),.din(w_dff_A_k3uNQ6l93_1),.clk(gclk));
	jdff dff_A_Y8g8JBsj4_0(.dout(w_G87_2[0]),.din(w_dff_A_Y8g8JBsj4_0),.clk(gclk));
	jdff dff_A_hRrX8oGS5_1(.dout(w_G87_0[1]),.din(w_dff_A_hRrX8oGS5_1),.clk(gclk));
	jdff dff_A_YfqCN7g38_1(.dout(w_dff_A_hRrX8oGS5_1),.din(w_dff_A_YfqCN7g38_1),.clk(gclk));
	jdff dff_A_Cb6U7dYo9_1(.dout(w_dff_A_YfqCN7g38_1),.din(w_dff_A_Cb6U7dYo9_1),.clk(gclk));
	jdff dff_A_SY8jVMB27_1(.dout(w_G68_3[1]),.din(w_dff_A_SY8jVMB27_1),.clk(gclk));
	jdff dff_A_fMQD3J5V6_1(.dout(w_dff_A_SY8jVMB27_1),.din(w_dff_A_fMQD3J5V6_1),.clk(gclk));
	jdff dff_A_zPbPefOx5_2(.dout(w_G68_3[2]),.din(w_dff_A_zPbPefOx5_2),.clk(gclk));
	jdff dff_A_c26WNJs30_2(.dout(w_dff_A_zPbPefOx5_2),.din(w_dff_A_c26WNJs30_2),.clk(gclk));
	jdff dff_A_XB9u5wBA3_2(.dout(w_G68_0[2]),.din(w_dff_A_XB9u5wBA3_2),.clk(gclk));
	jdff dff_A_WQ9NFfDz5_1(.dout(w_G190_2[1]),.din(w_dff_A_WQ9NFfDz5_1),.clk(gclk));
	jdff dff_A_tK2tHP670_1(.dout(w_dff_A_WQ9NFfDz5_1),.din(w_dff_A_tK2tHP670_1),.clk(gclk));
	jdff dff_A_YC9e3UYf0_1(.dout(w_dff_A_tK2tHP670_1),.din(w_dff_A_YC9e3UYf0_1),.clk(gclk));
	jdff dff_A_tz4ezU1Z1_2(.dout(w_G190_2[2]),.din(w_dff_A_tz4ezU1Z1_2),.clk(gclk));
	jdff dff_A_qt1oHG395_2(.dout(w_dff_A_tz4ezU1Z1_2),.din(w_dff_A_qt1oHG395_2),.clk(gclk));
	jdff dff_A_wyqwC8n39_2(.dout(w_dff_A_qt1oHG395_2),.din(w_dff_A_wyqwC8n39_2),.clk(gclk));
	jdff dff_A_zc5L4iXU9_1(.dout(w_G50_4[1]),.din(w_dff_A_zc5L4iXU9_1),.clk(gclk));
	jdff dff_A_w10T9dZ60_1(.dout(w_dff_A_zc5L4iXU9_1),.din(w_dff_A_w10T9dZ60_1),.clk(gclk));
	jdff dff_A_OKTHj1IG9_1(.dout(w_dff_A_w10T9dZ60_1),.din(w_dff_A_OKTHj1IG9_1),.clk(gclk));
	jdff dff_A_ybXPjCr49_2(.dout(w_G50_4[2]),.din(w_dff_A_ybXPjCr49_2),.clk(gclk));
	jdff dff_A_x1ZLCVR54_2(.dout(w_dff_A_ybXPjCr49_2),.din(w_dff_A_x1ZLCVR54_2),.clk(gclk));
	jdff dff_A_7IDlMxKm4_2(.dout(w_dff_A_x1ZLCVR54_2),.din(w_dff_A_7IDlMxKm4_2),.clk(gclk));
	jdff dff_A_UhOdz5az7_2(.dout(w_G50_0[2]),.din(w_dff_A_UhOdz5az7_2),.clk(gclk));
	jdff dff_A_3YOwGcrz0_2(.dout(w_dff_A_UhOdz5az7_2),.din(w_dff_A_3YOwGcrz0_2),.clk(gclk));
	jdff dff_A_XteHk1YD6_2(.dout(w_dff_A_3YOwGcrz0_2),.din(w_dff_A_XteHk1YD6_2),.clk(gclk));
	jdff dff_A_OoJdkKVT5_1(.dout(w_G200_1[1]),.din(w_dff_A_OoJdkKVT5_1),.clk(gclk));
	jdff dff_A_V3ZYA3xF7_1(.dout(w_dff_A_OoJdkKVT5_1),.din(w_dff_A_V3ZYA3xF7_1),.clk(gclk));
	jdff dff_A_WATa9lbd5_1(.dout(w_dff_A_V3ZYA3xF7_1),.din(w_dff_A_WATa9lbd5_1),.clk(gclk));
	jdff dff_A_ca7ACg321_1(.dout(w_dff_A_WATa9lbd5_1),.din(w_dff_A_ca7ACg321_1),.clk(gclk));
	jdff dff_A_PiKjDvWl7_1(.dout(w_dff_A_ca7ACg321_1),.din(w_dff_A_PiKjDvWl7_1),.clk(gclk));
	jdff dff_A_RsJcQgEB6_1(.dout(w_dff_A_PiKjDvWl7_1),.din(w_dff_A_RsJcQgEB6_1),.clk(gclk));
	jdff dff_A_0wkcZKDD1_2(.dout(w_G200_1[2]),.din(w_dff_A_0wkcZKDD1_2),.clk(gclk));
	jdff dff_A_vETwgtEH4_2(.dout(w_dff_A_0wkcZKDD1_2),.din(w_dff_A_vETwgtEH4_2),.clk(gclk));
	jdff dff_A_5AcsddxH0_2(.dout(w_dff_A_vETwgtEH4_2),.din(w_dff_A_5AcsddxH0_2),.clk(gclk));
	jdff dff_A_z83nPjcq3_2(.dout(w_dff_A_5AcsddxH0_2),.din(w_dff_A_z83nPjcq3_2),.clk(gclk));
	jdff dff_A_Eme40qrN6_2(.dout(w_dff_A_z83nPjcq3_2),.din(w_dff_A_Eme40qrN6_2),.clk(gclk));
	jdff dff_A_BHi2T2dg0_2(.dout(w_G20_3[2]),.din(w_dff_A_BHi2T2dg0_2),.clk(gclk));
	jdff dff_A_xIcLbesx1_1(.dout(w_n191_1[1]),.din(w_dff_A_xIcLbesx1_1),.clk(gclk));
	jdff dff_A_Ue9sukoG5_1(.dout(w_dff_A_xIcLbesx1_1),.din(w_dff_A_Ue9sukoG5_1),.clk(gclk));
	jdff dff_A_3LU1iai92_1(.dout(w_dff_A_Ue9sukoG5_1),.din(w_dff_A_3LU1iai92_1),.clk(gclk));
	jdff dff_A_XEtSx5NJ2_1(.dout(w_dff_A_3LU1iai92_1),.din(w_dff_A_XEtSx5NJ2_1),.clk(gclk));
	jdff dff_A_CLNDS7V07_1(.dout(w_dff_A_XEtSx5NJ2_1),.din(w_dff_A_CLNDS7V07_1),.clk(gclk));
	jdff dff_A_KTSnkItS2_2(.dout(w_n191_1[2]),.din(w_dff_A_KTSnkItS2_2),.clk(gclk));
	jdff dff_A_F1j5wBK80_2(.dout(w_dff_A_KTSnkItS2_2),.din(w_dff_A_F1j5wBK80_2),.clk(gclk));
	jdff dff_A_OH7CtWHC1_2(.dout(w_dff_A_F1j5wBK80_2),.din(w_dff_A_OH7CtWHC1_2),.clk(gclk));
	jdff dff_A_BxkjGqqB8_2(.dout(w_dff_A_OH7CtWHC1_2),.din(w_dff_A_BxkjGqqB8_2),.clk(gclk));
	jdff dff_A_vh7UCrih5_2(.dout(w_n284_1[2]),.din(w_dff_A_vh7UCrih5_2),.clk(gclk));
	jdff dff_A_CKJkWGGl9_2(.dout(w_dff_A_vh7UCrih5_2),.din(w_dff_A_CKJkWGGl9_2),.clk(gclk));
	jdff dff_A_1TN1V6Zt4_2(.dout(w_dff_A_CKJkWGGl9_2),.din(w_dff_A_1TN1V6Zt4_2),.clk(gclk));
	jdff dff_A_0sn6RaSv1_0(.dout(w_n284_0[0]),.din(w_dff_A_0sn6RaSv1_0),.clk(gclk));
	jdff dff_A_XlLw9ZLW4_1(.dout(w_n284_0[1]),.din(w_dff_A_XlLw9ZLW4_1),.clk(gclk));
	jdff dff_A_t19azNHw0_0(.dout(w_G107_0[0]),.din(w_dff_A_t19azNHw0_0),.clk(gclk));
	jdff dff_A_5B2x4W2w6_0(.dout(w_dff_A_t19azNHw0_0),.din(w_dff_A_5B2x4W2w6_0),.clk(gclk));
	jdff dff_A_CwrNi5cu0_0(.dout(w_dff_A_5B2x4W2w6_0),.din(w_dff_A_CwrNi5cu0_0),.clk(gclk));
	jdff dff_A_QWWvgvKW9_1(.dout(w_G107_0[1]),.din(w_dff_A_QWWvgvKW9_1),.clk(gclk));
	jdff dff_A_2mcTbHyJ7_1(.dout(w_dff_A_QWWvgvKW9_1),.din(w_dff_A_2mcTbHyJ7_1),.clk(gclk));
	jdff dff_A_AeYLXE9H6_1(.dout(w_dff_A_2mcTbHyJ7_1),.din(w_dff_A_AeYLXE9H6_1),.clk(gclk));
	jdff dff_A_Mt88KHO83_0(.dout(w_G33_6[0]),.din(w_dff_A_Mt88KHO83_0),.clk(gclk));
	jdff dff_A_1wDiKAeu7_0(.dout(w_dff_A_Mt88KHO83_0),.din(w_dff_A_1wDiKAeu7_0),.clk(gclk));
	jdff dff_A_0V8mqk7o9_1(.dout(w_G33_6[1]),.din(w_dff_A_0V8mqk7o9_1),.clk(gclk));
	jdff dff_A_uVpjaaK94_1(.dout(w_dff_A_0V8mqk7o9_1),.din(w_dff_A_uVpjaaK94_1),.clk(gclk));
	jdff dff_A_czSiPcGG6_1(.dout(w_dff_A_uVpjaaK94_1),.din(w_dff_A_czSiPcGG6_1),.clk(gclk));
	jdff dff_A_HEG50RAb2_0(.dout(w_G33_1[0]),.din(w_dff_A_HEG50RAb2_0),.clk(gclk));
	jdff dff_A_d4tqvVTr0_0(.dout(w_dff_A_HEG50RAb2_0),.din(w_dff_A_d4tqvVTr0_0),.clk(gclk));
	jdff dff_A_hsbDY3rh5_0(.dout(w_dff_A_d4tqvVTr0_0),.din(w_dff_A_hsbDY3rh5_0),.clk(gclk));
	jdff dff_A_xFE0W88I6_1(.dout(w_G33_1[1]),.din(w_dff_A_xFE0W88I6_1),.clk(gclk));
	jdff dff_A_PouHlUSh2_1(.dout(w_dff_A_xFE0W88I6_1),.din(w_dff_A_PouHlUSh2_1),.clk(gclk));
	jdff dff_A_Earr44st9_1(.dout(w_dff_A_PouHlUSh2_1),.din(w_dff_A_Earr44st9_1),.clk(gclk));
	jdff dff_A_U81WuUBA8_0(.dout(w_n579_1[0]),.din(w_dff_A_U81WuUBA8_0),.clk(gclk));
	jdff dff_A_kPdL6L0q5_0(.dout(w_dff_A_U81WuUBA8_0),.din(w_dff_A_kPdL6L0q5_0),.clk(gclk));
	jdff dff_A_a4bonOBI8_0(.dout(w_dff_A_kPdL6L0q5_0),.din(w_dff_A_a4bonOBI8_0),.clk(gclk));
	jdff dff_A_6lhPNLrv1_0(.dout(w_dff_A_a4bonOBI8_0),.din(w_dff_A_6lhPNLrv1_0),.clk(gclk));
	jdff dff_A_iV1NPdKu0_0(.dout(w_dff_A_6lhPNLrv1_0),.din(w_dff_A_iV1NPdKu0_0),.clk(gclk));
	jdff dff_A_iH1O1xLw5_0(.dout(w_dff_A_iV1NPdKu0_0),.din(w_dff_A_iH1O1xLw5_0),.clk(gclk));
	jdff dff_A_YQ8M2Mcf1_0(.dout(w_dff_A_iH1O1xLw5_0),.din(w_dff_A_YQ8M2Mcf1_0),.clk(gclk));
	jdff dff_A_UrjXRtc59_2(.dout(w_n579_1[2]),.din(w_dff_A_UrjXRtc59_2),.clk(gclk));
	jdff dff_A_cAOo0EWf3_2(.dout(w_dff_A_UrjXRtc59_2),.din(w_dff_A_cAOo0EWf3_2),.clk(gclk));
	jdff dff_A_dKytGgwp2_2(.dout(w_dff_A_cAOo0EWf3_2),.din(w_dff_A_dKytGgwp2_2),.clk(gclk));
	jdff dff_A_eNB2q96Y2_2(.dout(w_dff_A_dKytGgwp2_2),.din(w_dff_A_eNB2q96Y2_2),.clk(gclk));
	jdff dff_A_LSMCeX8K1_2(.dout(w_dff_A_eNB2q96Y2_2),.din(w_dff_A_LSMCeX8K1_2),.clk(gclk));
	jdff dff_A_zJh6XiLg1_2(.dout(w_dff_A_LSMCeX8K1_2),.din(w_dff_A_zJh6XiLg1_2),.clk(gclk));
	jdff dff_A_epqVj9Gl4_2(.dout(w_dff_A_zJh6XiLg1_2),.din(w_dff_A_epqVj9Gl4_2),.clk(gclk));
	jdff dff_A_Sf5n20R13_2(.dout(w_dff_A_epqVj9Gl4_2),.din(w_dff_A_Sf5n20R13_2),.clk(gclk));
	jdff dff_A_3OQCcMXd8_1(.dout(w_n579_0[1]),.din(w_dff_A_3OQCcMXd8_1),.clk(gclk));
	jdff dff_A_29Z0gz3k4_1(.dout(w_dff_A_3OQCcMXd8_1),.din(w_dff_A_29Z0gz3k4_1),.clk(gclk));
	jdff dff_A_0TjFo9LS7_1(.dout(w_dff_A_29Z0gz3k4_1),.din(w_dff_A_0TjFo9LS7_1),.clk(gclk));
	jdff dff_A_QNqpnw0L2_1(.dout(w_dff_A_0TjFo9LS7_1),.din(w_dff_A_QNqpnw0L2_1),.clk(gclk));
	jdff dff_A_TiC7mZPB2_1(.dout(w_dff_A_QNqpnw0L2_1),.din(w_dff_A_TiC7mZPB2_1),.clk(gclk));
	jdff dff_A_JQ5IT0bb7_1(.dout(w_dff_A_TiC7mZPB2_1),.din(w_dff_A_JQ5IT0bb7_1),.clk(gclk));
	jdff dff_A_uDlIdtm69_1(.dout(w_dff_A_JQ5IT0bb7_1),.din(w_dff_A_uDlIdtm69_1),.clk(gclk));
	jdff dff_A_OqOZjD7v9_1(.dout(w_dff_A_uDlIdtm69_1),.din(w_dff_A_OqOZjD7v9_1),.clk(gclk));
	jdff dff_A_Tc0cGRKe8_1(.dout(w_dff_A_OqOZjD7v9_1),.din(w_dff_A_Tc0cGRKe8_1),.clk(gclk));
	jdff dff_A_7WM1I46y6_2(.dout(w_n579_0[2]),.din(w_dff_A_7WM1I46y6_2),.clk(gclk));
	jdff dff_A_oOwsZbF53_2(.dout(w_dff_A_7WM1I46y6_2),.din(w_dff_A_oOwsZbF53_2),.clk(gclk));
	jdff dff_A_gXxOmiAh1_2(.dout(w_dff_A_oOwsZbF53_2),.din(w_dff_A_gXxOmiAh1_2),.clk(gclk));
	jdff dff_A_isXvbwmC7_2(.dout(w_dff_A_gXxOmiAh1_2),.din(w_dff_A_isXvbwmC7_2),.clk(gclk));
	jdff dff_A_YEKzohOc6_2(.dout(w_dff_A_isXvbwmC7_2),.din(w_dff_A_YEKzohOc6_2),.clk(gclk));
	jdff dff_A_ypt91aZp8_2(.dout(w_dff_A_YEKzohOc6_2),.din(w_dff_A_ypt91aZp8_2),.clk(gclk));
	jdff dff_A_3VbCZcko9_2(.dout(w_dff_A_ypt91aZp8_2),.din(w_dff_A_3VbCZcko9_2),.clk(gclk));
	jdff dff_A_vQcL9gd23_0(.dout(w_n578_2[0]),.din(w_dff_A_vQcL9gd23_0),.clk(gclk));
	jdff dff_A_7ODBYoAU0_0(.dout(w_dff_A_vQcL9gd23_0),.din(w_dff_A_7ODBYoAU0_0),.clk(gclk));
	jdff dff_A_aJkDY9jT9_0(.dout(w_dff_A_7ODBYoAU0_0),.din(w_dff_A_aJkDY9jT9_0),.clk(gclk));
	jdff dff_A_xoPW5xzo0_0(.dout(w_dff_A_aJkDY9jT9_0),.din(w_dff_A_xoPW5xzo0_0),.clk(gclk));
	jdff dff_A_1VmBzJMq9_0(.dout(w_dff_A_xoPW5xzo0_0),.din(w_dff_A_1VmBzJMq9_0),.clk(gclk));
	jdff dff_A_KNWpJ1814_0(.dout(w_dff_A_1VmBzJMq9_0),.din(w_dff_A_KNWpJ1814_0),.clk(gclk));
	jdff dff_A_ognYgis48_0(.dout(w_dff_A_KNWpJ1814_0),.din(w_dff_A_ognYgis48_0),.clk(gclk));
	jdff dff_A_qoKVMUri9_0(.dout(w_dff_A_ognYgis48_0),.din(w_dff_A_qoKVMUri9_0),.clk(gclk));
	jdff dff_A_FK04W79i4_0(.dout(w_dff_A_qoKVMUri9_0),.din(w_dff_A_FK04W79i4_0),.clk(gclk));
	jdff dff_A_JILh3T5A3_2(.dout(w_n578_0[2]),.din(w_dff_A_JILh3T5A3_2),.clk(gclk));
	jdff dff_A_Rb6AHIed4_2(.dout(w_dff_A_JILh3T5A3_2),.din(w_dff_A_Rb6AHIed4_2),.clk(gclk));
	jdff dff_A_0jl5l4hp5_2(.dout(w_dff_A_Rb6AHIed4_2),.din(w_dff_A_0jl5l4hp5_2),.clk(gclk));
	jdff dff_A_6MEQgBni0_2(.dout(w_dff_A_0jl5l4hp5_2),.din(w_dff_A_6MEQgBni0_2),.clk(gclk));
	jdff dff_A_ymmBDbG78_2(.dout(w_dff_A_6MEQgBni0_2),.din(w_dff_A_ymmBDbG78_2),.clk(gclk));
	jdff dff_A_dH2z5x6g4_2(.dout(w_dff_A_ymmBDbG78_2),.din(w_dff_A_dH2z5x6g4_2),.clk(gclk));
	jdff dff_A_DbuiHhS49_2(.dout(w_dff_A_dH2z5x6g4_2),.din(w_dff_A_DbuiHhS49_2),.clk(gclk));
	jdff dff_A_Kh0W7LJm7_0(.dout(w_n153_5[0]),.din(w_dff_A_Kh0W7LJm7_0),.clk(gclk));
	jdff dff_A_9qTpjvg52_0(.dout(w_dff_A_Kh0W7LJm7_0),.din(w_dff_A_9qTpjvg52_0),.clk(gclk));
	jdff dff_A_BrtoE2Cx9_1(.dout(w_n153_5[1]),.din(w_dff_A_BrtoE2Cx9_1),.clk(gclk));
	jdff dff_A_RzBvpja00_1(.dout(w_dff_A_BrtoE2Cx9_1),.din(w_dff_A_RzBvpja00_1),.clk(gclk));
	jdff dff_A_8PiacHDd5_1(.dout(w_dff_A_RzBvpja00_1),.din(w_dff_A_8PiacHDd5_1),.clk(gclk));
	jdff dff_A_SpgKQ8sL4_0(.dout(w_n153_1[0]),.din(w_dff_A_SpgKQ8sL4_0),.clk(gclk));
	jdff dff_A_9cZizQgL7_0(.dout(w_dff_A_SpgKQ8sL4_0),.din(w_dff_A_9cZizQgL7_0),.clk(gclk));
	jdff dff_A_la4Lg7iy3_0(.dout(w_dff_A_9cZizQgL7_0),.din(w_dff_A_la4Lg7iy3_0),.clk(gclk));
	jdff dff_B_8219FGGN1_0(.din(n532),.dout(w_dff_B_8219FGGN1_0),.clk(gclk));
	jdff dff_B_qv6ztYWL1_0(.din(w_dff_B_8219FGGN1_0),.dout(w_dff_B_qv6ztYWL1_0),.clk(gclk));
	jdff dff_A_fAgM6g8M2_2(.dout(w_n531_4[2]),.din(w_dff_A_fAgM6g8M2_2),.clk(gclk));
	jdff dff_A_N4SXkTLS6_2(.dout(w_dff_A_fAgM6g8M2_2),.din(w_dff_A_N4SXkTLS6_2),.clk(gclk));
	jdff dff_A_2jLXFuQv9_2(.dout(w_dff_A_N4SXkTLS6_2),.din(w_dff_A_2jLXFuQv9_2),.clk(gclk));
	jdff dff_A_KAwmpeJO5_1(.dout(w_n531_1[1]),.din(w_dff_A_KAwmpeJO5_1),.clk(gclk));
	jdff dff_A_bDA0GVVs0_1(.dout(w_dff_A_KAwmpeJO5_1),.din(w_dff_A_bDA0GVVs0_1),.clk(gclk));
	jdff dff_A_9E02IJP68_2(.dout(w_n531_1[2]),.din(w_dff_A_9E02IJP68_2),.clk(gclk));
	jdff dff_A_BllAhk3v7_1(.dout(w_n531_0[1]),.din(w_dff_A_BllAhk3v7_1),.clk(gclk));
	jdff dff_A_Jx4UkCvz0_1(.dout(w_dff_A_BllAhk3v7_1),.din(w_dff_A_Jx4UkCvz0_1),.clk(gclk));
	jdff dff_A_lSEecwiY4_1(.dout(w_dff_A_Jx4UkCvz0_1),.din(w_dff_A_lSEecwiY4_1),.clk(gclk));
	jdff dff_A_4gOG3Ltk0_2(.dout(w_n531_0[2]),.din(w_dff_A_4gOG3Ltk0_2),.clk(gclk));
	jdff dff_A_zi7A3axm0_0(.dout(w_n530_1[0]),.din(w_dff_A_zi7A3axm0_0),.clk(gclk));
	jdff dff_A_xDdIks2k5_0(.dout(w_dff_A_zi7A3axm0_0),.din(w_dff_A_xDdIks2k5_0),.clk(gclk));
	jdff dff_A_YLiZrEYK7_0(.dout(w_dff_A_xDdIks2k5_0),.din(w_dff_A_YLiZrEYK7_0),.clk(gclk));
	jdff dff_A_HbCePM388_0(.dout(w_dff_A_YLiZrEYK7_0),.din(w_dff_A_HbCePM388_0),.clk(gclk));
	jdff dff_A_f3NzufjE0_0(.dout(w_dff_A_HbCePM388_0),.din(w_dff_A_f3NzufjE0_0),.clk(gclk));
	jdff dff_A_9S3vw8Ew3_0(.dout(w_dff_A_f3NzufjE0_0),.din(w_dff_A_9S3vw8Ew3_0),.clk(gclk));
	jdff dff_A_VpS1disS9_1(.dout(w_n530_0[1]),.din(w_dff_A_VpS1disS9_1),.clk(gclk));
	jdff dff_A_XWODCJk37_1(.dout(w_dff_A_VpS1disS9_1),.din(w_dff_A_XWODCJk37_1),.clk(gclk));
	jdff dff_A_hkOcqSpi0_1(.dout(w_dff_A_XWODCJk37_1),.din(w_dff_A_hkOcqSpi0_1),.clk(gclk));
	jdff dff_A_f9fPes1r4_1(.dout(w_dff_A_hkOcqSpi0_1),.din(w_dff_A_f9fPes1r4_1),.clk(gclk));
	jdff dff_A_KPYgOAhA6_2(.dout(w_n530_0[2]),.din(w_dff_A_KPYgOAhA6_2),.clk(gclk));
	jdff dff_A_SDOExKsY0_2(.dout(w_dff_A_KPYgOAhA6_2),.din(w_dff_A_SDOExKsY0_2),.clk(gclk));
	jdff dff_A_tc25riLF0_2(.dout(w_dff_A_SDOExKsY0_2),.din(w_dff_A_tc25riLF0_2),.clk(gclk));
	jdff dff_A_emKsr4Fg6_2(.dout(w_dff_A_tc25riLF0_2),.din(w_dff_A_emKsr4Fg6_2),.clk(gclk));
	jdff dff_A_0tYGGUoq8_1(.dout(w_G213_0[1]),.din(w_dff_A_0tYGGUoq8_1),.clk(gclk));
	jdff dff_A_j1hc41OV4_1(.dout(w_G343_0[1]),.din(w_dff_A_j1hc41OV4_1),.clk(gclk));
	jdff dff_A_paEEYKD64_1(.dout(w_dff_A_j1hc41OV4_1),.din(w_dff_A_paEEYKD64_1),.clk(gclk));
	jdff dff_B_t80UjEDy7_2(.din(G343),.dout(w_dff_B_t80UjEDy7_2),.clk(gclk));
	jdff dff_A_xfzRTbUX5_1(.dout(w_n208_0[1]),.din(w_dff_A_xfzRTbUX5_1),.clk(gclk));
	jdff dff_A_Cc185wxx8_1(.dout(w_dff_A_xfzRTbUX5_1),.din(w_dff_A_Cc185wxx8_1),.clk(gclk));
	jdff dff_A_QKpOV3Co8_1(.dout(w_dff_A_Cc185wxx8_1),.din(w_dff_A_QKpOV3Co8_1),.clk(gclk));
	jdff dff_B_lZ0KuJ4o5_1(.din(n203),.dout(w_dff_B_lZ0KuJ4o5_1),.clk(gclk));
	jdff dff_B_Di3rUeFI3_1(.din(w_dff_B_lZ0KuJ4o5_1),.dout(w_dff_B_Di3rUeFI3_1),.clk(gclk));
	jdff dff_A_Y8hYC2IV0_1(.dout(w_G190_4[1]),.din(w_dff_A_Y8hYC2IV0_1),.clk(gclk));
	jdff dff_A_RA89g64K2_1(.dout(w_dff_A_Y8hYC2IV0_1),.din(w_dff_A_RA89g64K2_1),.clk(gclk));
	jdff dff_A_DnLvpEAF5_1(.dout(w_dff_A_RA89g64K2_1),.din(w_dff_A_DnLvpEAF5_1),.clk(gclk));
	jdff dff_A_xIPSMYqF5_1(.dout(w_dff_A_DnLvpEAF5_1),.din(w_dff_A_xIPSMYqF5_1),.clk(gclk));
	jdff dff_A_x5iny7C70_1(.dout(w_dff_A_xIPSMYqF5_1),.din(w_dff_A_x5iny7C70_1),.clk(gclk));
	jdff dff_A_hRzyRzXw2_1(.dout(w_dff_A_x5iny7C70_1),.din(w_dff_A_hRzyRzXw2_1),.clk(gclk));
	jdff dff_A_AZKHoWiQ4_2(.dout(w_G190_4[2]),.din(w_dff_A_AZKHoWiQ4_2),.clk(gclk));
	jdff dff_A_36D7eIJr5_2(.dout(w_dff_A_AZKHoWiQ4_2),.din(w_dff_A_36D7eIJr5_2),.clk(gclk));
	jdff dff_A_Yym9ARtr7_2(.dout(w_dff_A_36D7eIJr5_2),.din(w_dff_A_Yym9ARtr7_2),.clk(gclk));
	jdff dff_A_Q8nlyQ1Z4_2(.dout(w_dff_A_Yym9ARtr7_2),.din(w_dff_A_Q8nlyQ1Z4_2),.clk(gclk));
	jdff dff_A_xYaBeaJI4_2(.dout(w_dff_A_Q8nlyQ1Z4_2),.din(w_dff_A_xYaBeaJI4_2),.clk(gclk));
	jdff dff_A_gwt26j987_2(.dout(w_dff_A_xYaBeaJI4_2),.din(w_dff_A_gwt26j987_2),.clk(gclk));
	jdff dff_A_a5fQVTzg2_2(.dout(w_dff_A_gwt26j987_2),.din(w_dff_A_a5fQVTzg2_2),.clk(gclk));
	jdff dff_A_eNK4R6Wc2_1(.dout(w_G190_1[1]),.din(w_dff_A_eNK4R6Wc2_1),.clk(gclk));
	jdff dff_A_9znQbK8K4_1(.dout(w_dff_A_eNK4R6Wc2_1),.din(w_dff_A_9znQbK8K4_1),.clk(gclk));
	jdff dff_A_Pjipn1Bh4_2(.dout(w_G190_1[2]),.din(w_dff_A_Pjipn1Bh4_2),.clk(gclk));
	jdff dff_A_VnHop4lI8_2(.dout(w_dff_A_Pjipn1Bh4_2),.din(w_dff_A_VnHop4lI8_2),.clk(gclk));
	jdff dff_A_YReyY20D5_1(.dout(w_G190_0[1]),.din(w_dff_A_YReyY20D5_1),.clk(gclk));
	jdff dff_A_zFoFmfc91_1(.dout(w_dff_A_YReyY20D5_1),.din(w_dff_A_zFoFmfc91_1),.clk(gclk));
	jdff dff_A_HA43TPzI4_2(.dout(w_G190_0[2]),.din(w_dff_A_HA43TPzI4_2),.clk(gclk));
	jdff dff_A_cVCIdqAS5_2(.dout(w_dff_A_HA43TPzI4_2),.din(w_dff_A_cVCIdqAS5_2),.clk(gclk));
	jdff dff_A_fEYszTsu9_2(.dout(w_dff_A_cVCIdqAS5_2),.din(w_dff_A_fEYszTsu9_2),.clk(gclk));
	jdff dff_A_YCFcJsKT1_2(.dout(w_dff_A_fEYszTsu9_2),.din(w_dff_A_YCFcJsKT1_2),.clk(gclk));
	jdff dff_A_pvLVCwaM3_2(.dout(w_dff_A_YCFcJsKT1_2),.din(w_dff_A_pvLVCwaM3_2),.clk(gclk));
	jdff dff_A_3eBytgpX4_1(.dout(w_n204_0[1]),.din(w_dff_A_3eBytgpX4_1),.clk(gclk));
	jdff dff_A_3usa37dt1_1(.dout(w_G200_2[1]),.din(w_dff_A_3usa37dt1_1),.clk(gclk));
	jdff dff_A_e0xAzYEy0_1(.dout(w_dff_A_3usa37dt1_1),.din(w_dff_A_e0xAzYEy0_1),.clk(gclk));
	jdff dff_A_Byv1Yxey2_1(.dout(w_dff_A_e0xAzYEy0_1),.din(w_dff_A_Byv1Yxey2_1),.clk(gclk));
	jdff dff_A_yDQKd7iq0_1(.dout(w_dff_A_Byv1Yxey2_1),.din(w_dff_A_yDQKd7iq0_1),.clk(gclk));
	jdff dff_A_AdX3ri1D4_1(.dout(w_dff_A_yDQKd7iq0_1),.din(w_dff_A_AdX3ri1D4_1),.clk(gclk));
	jdff dff_A_8rPchjsM9_2(.dout(w_G200_0[2]),.din(w_dff_A_8rPchjsM9_2),.clk(gclk));
	jdff dff_A_qvasqyZf6_1(.dout(w_n202_0[1]),.din(w_dff_A_qvasqyZf6_1),.clk(gclk));
	jdff dff_A_ABYWI6VE8_1(.dout(w_n200_0[1]),.din(w_dff_A_ABYWI6VE8_1),.clk(gclk));
	jdff dff_A_fvx1FcJL2_1(.dout(w_dff_A_ABYWI6VE8_1),.din(w_dff_A_fvx1FcJL2_1),.clk(gclk));
	jdff dff_A_0ywe8Y0j3_0(.dout(w_n199_0[0]),.din(w_dff_A_0ywe8Y0j3_0),.clk(gclk));
	jdff dff_B_gF9WsJ4t1_0(.din(n197),.dout(w_dff_B_gF9WsJ4t1_0),.clk(gclk));
	jdff dff_A_hSILwcqq7_2(.dout(w_n167_3[2]),.din(w_dff_A_hSILwcqq7_2),.clk(gclk));
	jdff dff_A_fj4txxlY0_0(.dout(w_n193_0[0]),.din(w_dff_A_fj4txxlY0_0),.clk(gclk));
	jdff dff_A_czs1bfAp0_2(.dout(w_n193_0[2]),.din(w_dff_A_czs1bfAp0_2),.clk(gclk));
	jdff dff_A_XCdy0zIb4_0(.dout(w_n191_3[0]),.din(w_dff_A_XCdy0zIb4_0),.clk(gclk));
	jdff dff_A_0IZjeug70_0(.dout(w_dff_A_XCdy0zIb4_0),.din(w_dff_A_0IZjeug70_0),.clk(gclk));
	jdff dff_A_zyKZmBA41_0(.dout(w_dff_A_0IZjeug70_0),.din(w_dff_A_zyKZmBA41_0),.clk(gclk));
	jdff dff_A_v5J5apna9_1(.dout(w_n191_3[1]),.din(w_dff_A_v5J5apna9_1),.clk(gclk));
	jdff dff_A_DV6vWHAV8_1(.dout(w_n191_0[1]),.din(w_dff_A_DV6vWHAV8_1),.clk(gclk));
	jdff dff_A_yfwxKucK7_1(.dout(w_dff_A_DV6vWHAV8_1),.din(w_dff_A_yfwxKucK7_1),.clk(gclk));
	jdff dff_A_aqfcMpWq8_1(.dout(w_dff_A_yfwxKucK7_1),.din(w_dff_A_aqfcMpWq8_1),.clk(gclk));
	jdff dff_A_KpbIBopu1_1(.dout(w_dff_A_aqfcMpWq8_1),.din(w_dff_A_KpbIBopu1_1),.clk(gclk));
	jdff dff_A_VCMu02xU2_2(.dout(w_n191_0[2]),.din(w_dff_A_VCMu02xU2_2),.clk(gclk));
	jdff dff_A_CTDjGbnj1_2(.dout(w_dff_A_VCMu02xU2_2),.din(w_dff_A_CTDjGbnj1_2),.clk(gclk));
	jdff dff_A_GKRYpEuA5_2(.dout(w_dff_A_CTDjGbnj1_2),.din(w_dff_A_GKRYpEuA5_2),.clk(gclk));
	jdff dff_A_DSBvx0Ah3_2(.dout(w_dff_A_GKRYpEuA5_2),.din(w_dff_A_DSBvx0Ah3_2),.clk(gclk));
	jdff dff_A_JS0tIAsY3_0(.dout(w_G179_1[0]),.din(w_dff_A_JS0tIAsY3_0),.clk(gclk));
	jdff dff_A_dzOtopaT8_0(.dout(w_dff_A_JS0tIAsY3_0),.din(w_dff_A_dzOtopaT8_0),.clk(gclk));
	jdff dff_A_drWM7Ylr6_0(.dout(w_dff_A_dzOtopaT8_0),.din(w_dff_A_drWM7Ylr6_0),.clk(gclk));
	jdff dff_A_hPZj13FQ6_0(.dout(w_dff_A_drWM7Ylr6_0),.din(w_dff_A_hPZj13FQ6_0),.clk(gclk));
	jdff dff_A_0wL0cO0E4_2(.dout(w_G179_0[2]),.din(w_dff_A_0wL0cO0E4_2),.clk(gclk));
	jdff dff_A_fe3aKREo2_2(.dout(w_dff_A_0wL0cO0E4_2),.din(w_dff_A_fe3aKREo2_2),.clk(gclk));
	jdff dff_A_KMDWpFI76_2(.dout(w_dff_A_fe3aKREo2_2),.din(w_dff_A_KMDWpFI76_2),.clk(gclk));
	jdff dff_A_I11MkcQE4_2(.dout(w_dff_A_KMDWpFI76_2),.din(w_dff_A_I11MkcQE4_2),.clk(gclk));
	jdff dff_A_1ehwWKnk4_2(.dout(w_dff_A_I11MkcQE4_2),.din(w_dff_A_1ehwWKnk4_2),.clk(gclk));
	jdff dff_A_1pMPP5rW9_2(.dout(w_dff_A_1ehwWKnk4_2),.din(w_dff_A_1pMPP5rW9_2),.clk(gclk));
	jdff dff_A_0S5FIjkv8_1(.dout(w_n187_0[1]),.din(w_dff_A_0S5FIjkv8_1),.clk(gclk));
	jdff dff_A_KO3ZZ86d4_1(.dout(w_dff_A_0S5FIjkv8_1),.din(w_dff_A_KO3ZZ86d4_1),.clk(gclk));
	jdff dff_A_RJv6eMpf7_0(.dout(w_n113_0[0]),.din(w_dff_A_RJv6eMpf7_0),.clk(gclk));
	jdff dff_A_7GZeRR1V0_0(.dout(w_dff_A_RJv6eMpf7_0),.din(w_dff_A_7GZeRR1V0_0),.clk(gclk));
	jdff dff_A_L1LfM2zG9_0(.dout(w_G270_0[0]),.din(w_dff_A_L1LfM2zG9_0),.clk(gclk));
	jdff dff_A_fOVcn0cu7_1(.dout(w_n183_0[1]),.din(w_dff_A_fOVcn0cu7_1),.clk(gclk));
	jdff dff_B_h7yKL39l2_0(.din(n182),.dout(w_dff_B_h7yKL39l2_0),.clk(gclk));
	jdff dff_B_DAC8bilL0_3(.din(n181),.dout(w_dff_B_DAC8bilL0_3),.clk(gclk));
	jdff dff_A_jDCWKkcP8_1(.dout(w_G257_0[1]),.din(w_dff_A_jDCWKkcP8_1),.clk(gclk));
	jdff dff_A_VzEBntKb0_1(.dout(w_dff_A_jDCWKkcP8_1),.din(w_dff_A_VzEBntKb0_1),.clk(gclk));
	jdff dff_A_uivRfVn56_1(.dout(w_dff_A_VzEBntKb0_1),.din(w_dff_A_uivRfVn56_1),.clk(gclk));
	jdff dff_A_g5fnT28m4_1(.dout(w_dff_A_uivRfVn56_1),.din(w_dff_A_g5fnT28m4_1),.clk(gclk));
	jdff dff_A_5LXrVV437_2(.dout(w_G257_0[2]),.din(w_dff_A_5LXrVV437_2),.clk(gclk));
	jdff dff_A_1ZCCUhkB4_2(.dout(w_dff_A_5LXrVV437_2),.din(w_dff_A_1ZCCUhkB4_2),.clk(gclk));
	jdff dff_A_oQN1rgso3_0(.dout(w_G303_2[0]),.din(w_dff_A_oQN1rgso3_0),.clk(gclk));
	jdff dff_A_rJTuoJ295_0(.dout(w_dff_A_oQN1rgso3_0),.din(w_dff_A_rJTuoJ295_0),.clk(gclk));
	jdff dff_A_zIemMhgn9_0(.dout(w_dff_A_rJTuoJ295_0),.din(w_dff_A_zIemMhgn9_0),.clk(gclk));
	jdff dff_A_IMmRtMZE4_1(.dout(w_G303_2[1]),.din(w_dff_A_IMmRtMZE4_1),.clk(gclk));
	jdff dff_A_FG0ioKLT5_1(.dout(w_dff_A_IMmRtMZE4_1),.din(w_dff_A_FG0ioKLT5_1),.clk(gclk));
	jdff dff_A_WRB8si7u2_1(.dout(w_dff_A_FG0ioKLT5_1),.din(w_dff_A_WRB8si7u2_1),.clk(gclk));
	jdff dff_A_XPicNu6b4_0(.dout(w_G303_0[0]),.din(w_dff_A_XPicNu6b4_0),.clk(gclk));
	jdff dff_A_ynPFlVee7_0(.dout(w_dff_A_XPicNu6b4_0),.din(w_dff_A_ynPFlVee7_0),.clk(gclk));
	jdff dff_A_u9ZGdr624_0(.dout(w_dff_A_ynPFlVee7_0),.din(w_dff_A_u9ZGdr624_0),.clk(gclk));
	jdff dff_A_oYsg2RoG3_2(.dout(w_G303_0[2]),.din(w_dff_A_oYsg2RoG3_2),.clk(gclk));
	jdff dff_A_iH77Os1e9_2(.dout(w_dff_A_oYsg2RoG3_2),.din(w_dff_A_iH77Os1e9_2),.clk(gclk));
	jdff dff_A_gHd0RMZ40_2(.dout(w_dff_A_iH77Os1e9_2),.din(w_dff_A_gHd0RMZ40_2),.clk(gclk));
	jdff dff_A_w31GkA329_0(.dout(w_G33_9[0]),.din(w_dff_A_w31GkA329_0),.clk(gclk));
	jdff dff_A_Jh9CEhWh9_0(.dout(w_n177_0[0]),.din(w_dff_A_Jh9CEhWh9_0),.clk(gclk));
	jdff dff_A_iBXhMxwh8_2(.dout(w_G1698_0[2]),.din(w_dff_A_iBXhMxwh8_2),.clk(gclk));
	jdff dff_A_t7bk5ory4_0(.dout(w_G264_0[0]),.din(w_dff_A_t7bk5ory4_0),.clk(gclk));
	jdff dff_A_c1JWmLH73_0(.dout(w_dff_A_t7bk5ory4_0),.din(w_dff_A_c1JWmLH73_0),.clk(gclk));
	jdff dff_A_qWmm4XBe9_1(.dout(w_n175_3[1]),.din(w_dff_A_qWmm4XBe9_1),.clk(gclk));
	jdff dff_A_JyVyhI943_1(.dout(w_dff_A_qWmm4XBe9_1),.din(w_dff_A_JyVyhI943_1),.clk(gclk));
	jdff dff_A_B5Q1wpPz9_1(.dout(w_dff_A_JyVyhI943_1),.din(w_dff_A_B5Q1wpPz9_1),.clk(gclk));
	jdff dff_A_vatFgBln0_1(.dout(w_n175_0[1]),.din(w_dff_A_vatFgBln0_1),.clk(gclk));
	jdff dff_A_Aj3lUnKW1_0(.dout(w_n173_0[0]),.din(w_dff_A_Aj3lUnKW1_0),.clk(gclk));
	jdff dff_A_VrttsOYA9_2(.dout(w_n173_0[2]),.din(w_dff_A_VrttsOYA9_2),.clk(gclk));
	jdff dff_A_kQnQgSOO9_2(.dout(w_dff_A_VrttsOYA9_2),.din(w_dff_A_kQnQgSOO9_2),.clk(gclk));
	jdff dff_A_s8fqRlFn4_1(.dout(w_G45_1[1]),.din(w_dff_A_s8fqRlFn4_1),.clk(gclk));
	jdff dff_A_2myHAoyQ6_0(.dout(w_n143_1[0]),.din(w_dff_A_2myHAoyQ6_0),.clk(gclk));
	jdff dff_A_1Du0ZaHl4_0(.dout(w_dff_A_2myHAoyQ6_0),.din(w_dff_A_1Du0ZaHl4_0),.clk(gclk));
	jdff dff_A_oyhlAvoM2_0(.dout(w_dff_A_1Du0ZaHl4_0),.din(w_dff_A_oyhlAvoM2_0),.clk(gclk));
	jdff dff_A_Mwwm7nIY8_0(.dout(w_dff_A_oyhlAvoM2_0),.din(w_dff_A_Mwwm7nIY8_0),.clk(gclk));
	jdff dff_A_Uz9cwlyk5_0(.dout(w_dff_A_Mwwm7nIY8_0),.din(w_dff_A_Uz9cwlyk5_0),.clk(gclk));
	jdff dff_A_7Wmj5fAf5_0(.dout(w_dff_A_Uz9cwlyk5_0),.din(w_dff_A_7Wmj5fAf5_0),.clk(gclk));
	jdff dff_A_eBfeswso1_0(.dout(w_dff_A_7Wmj5fAf5_0),.din(w_dff_A_eBfeswso1_0),.clk(gclk));
	jdff dff_A_U6vvSeoE1_0(.dout(w_dff_A_eBfeswso1_0),.din(w_dff_A_U6vvSeoE1_0),.clk(gclk));
	jdff dff_A_SyUTfx7y4_0(.dout(w_dff_A_U6vvSeoE1_0),.din(w_dff_A_SyUTfx7y4_0),.clk(gclk));
	jdff dff_A_dH9Yogdq5_0(.dout(w_dff_A_SyUTfx7y4_0),.din(w_dff_A_dH9Yogdq5_0),.clk(gclk));
	jdff dff_A_CDWKKud07_0(.dout(w_dff_A_dH9Yogdq5_0),.din(w_dff_A_CDWKKud07_0),.clk(gclk));
	jdff dff_A_EdceNqbx6_0(.dout(w_dff_A_CDWKKud07_0),.din(w_dff_A_EdceNqbx6_0),.clk(gclk));
	jdff dff_A_XgFv67y14_0(.dout(w_dff_A_EdceNqbx6_0),.din(w_dff_A_XgFv67y14_0),.clk(gclk));
	jdff dff_A_0sdUi2d00_0(.dout(w_dff_A_XgFv67y14_0),.din(w_dff_A_0sdUi2d00_0),.clk(gclk));
	jdff dff_A_ucWjFwd26_0(.dout(w_dff_A_0sdUi2d00_0),.din(w_dff_A_ucWjFwd26_0),.clk(gclk));
	jdff dff_A_s2Qb03pe3_0(.dout(w_dff_A_ucWjFwd26_0),.din(w_dff_A_s2Qb03pe3_0),.clk(gclk));
	jdff dff_A_3ismzyuC2_0(.dout(w_dff_A_s2Qb03pe3_0),.din(w_dff_A_3ismzyuC2_0),.clk(gclk));
	jdff dff_A_ByMvWYW64_1(.dout(w_n169_1[1]),.din(w_dff_A_ByMvWYW64_1),.clk(gclk));
	jdff dff_A_JElLs7Gx3_1(.dout(w_n168_0[1]),.din(w_dff_A_JElLs7Gx3_1),.clk(gclk));
	jdff dff_B_rwldEtvG9_1(.din(n164),.dout(w_dff_B_rwldEtvG9_1),.clk(gclk));
	jdff dff_B_JapuFSpL8_1(.din(w_dff_B_rwldEtvG9_1),.dout(w_dff_B_JapuFSpL8_1),.clk(gclk));
	jdff dff_A_9J1j9XG43_0(.dout(w_n165_0[0]),.din(w_dff_A_9J1j9XG43_0),.clk(gclk));
	jdff dff_A_THLLKRTA2_0(.dout(w_G274_0[0]),.din(w_dff_A_THLLKRTA2_0),.clk(gclk));
	jdff dff_A_UOhAl3AG6_0(.dout(w_dff_A_THLLKRTA2_0),.din(w_dff_A_UOhAl3AG6_0),.clk(gclk));
	jdff dff_A_L3IOk9wr4_1(.dout(w_G274_0[1]),.din(w_dff_A_L3IOk9wr4_1),.clk(gclk));
	jdff dff_A_hXLqg86h2_1(.dout(w_dff_A_L3IOk9wr4_1),.din(w_dff_A_hXLqg86h2_1),.clk(gclk));
	jdff dff_A_iP9w2g1g0_1(.dout(w_n163_1[1]),.din(w_dff_A_iP9w2g1g0_1),.clk(gclk));
	jdff dff_A_Wjps8uhV2_1(.dout(w_dff_A_iP9w2g1g0_1),.din(w_dff_A_Wjps8uhV2_1),.clk(gclk));
	jdff dff_A_rWES0KiL5_1(.dout(w_n163_0[1]),.din(w_dff_A_rWES0KiL5_1),.clk(gclk));
	jdff dff_A_NWQxB7k92_1(.dout(w_dff_A_rWES0KiL5_1),.din(w_dff_A_NWQxB7k92_1),.clk(gclk));
	jdff dff_A_kIGrJzaO2_1(.dout(w_dff_A_NWQxB7k92_1),.din(w_dff_A_kIGrJzaO2_1),.clk(gclk));
	jdff dff_A_01IyBm3r8_2(.dout(w_n163_0[2]),.din(w_dff_A_01IyBm3r8_2),.clk(gclk));
	jdff dff_B_os1UX2Uh9_3(.din(n163),.dout(w_dff_B_os1UX2Uh9_3),.clk(gclk));
	jdff dff_B_zd5dVfUd6_3(.din(w_dff_B_os1UX2Uh9_3),.dout(w_dff_B_zd5dVfUd6_3),.clk(gclk));
	jdff dff_B_K5rKf5gl6_3(.din(w_dff_B_zd5dVfUd6_3),.dout(w_dff_B_K5rKf5gl6_3),.clk(gclk));
	jdff dff_B_988m3ij01_3(.din(w_dff_B_K5rKf5gl6_3),.dout(w_dff_B_988m3ij01_3),.clk(gclk));
	jdff dff_A_lbKQYAN26_0(.dout(w_G169_2[0]),.din(w_dff_A_lbKQYAN26_0),.clk(gclk));
	jdff dff_A_t4aTUrN55_0(.dout(w_dff_A_lbKQYAN26_0),.din(w_dff_A_t4aTUrN55_0),.clk(gclk));
	jdff dff_A_enyAnlgb9_0(.dout(w_dff_A_t4aTUrN55_0),.din(w_dff_A_enyAnlgb9_0),.clk(gclk));
	jdff dff_A_MBfHdSgu8_0(.dout(w_dff_A_enyAnlgb9_0),.din(w_dff_A_MBfHdSgu8_0),.clk(gclk));
	jdff dff_A_ce9dhZGO4_0(.dout(w_dff_A_MBfHdSgu8_0),.din(w_dff_A_ce9dhZGO4_0),.clk(gclk));
	jdff dff_A_jIv7nspd0_0(.dout(w_dff_A_ce9dhZGO4_0),.din(w_dff_A_jIv7nspd0_0),.clk(gclk));
	jdff dff_A_7bDZaXzh3_0(.dout(w_G169_0[0]),.din(w_dff_A_7bDZaXzh3_0),.clk(gclk));
	jdff dff_A_v7mod6Fz3_0(.dout(w_dff_A_7bDZaXzh3_0),.din(w_dff_A_v7mod6Fz3_0),.clk(gclk));
	jdff dff_A_YQABj98p0_0(.dout(w_dff_A_v7mod6Fz3_0),.din(w_dff_A_YQABj98p0_0),.clk(gclk));
	jdff dff_A_Nhg0tDvh7_0(.dout(w_dff_A_YQABj98p0_0),.din(w_dff_A_Nhg0tDvh7_0),.clk(gclk));
	jdff dff_A_cKU9WJCE0_0(.dout(w_dff_A_Nhg0tDvh7_0),.din(w_dff_A_cKU9WJCE0_0),.clk(gclk));
	jdff dff_A_OacZVhaD0_2(.dout(w_G169_0[2]),.din(w_dff_A_OacZVhaD0_2),.clk(gclk));
	jdff dff_A_Tjp1h7dN3_1(.dout(w_n162_0[1]),.din(w_dff_A_Tjp1h7dN3_1),.clk(gclk));
	jdff dff_A_s1ptZKpM2_1(.dout(w_dff_A_Tjp1h7dN3_1),.din(w_dff_A_s1ptZKpM2_1),.clk(gclk));
	jdff dff_B_9wQpPHUb9_1(.din(n149),.dout(w_dff_B_9wQpPHUb9_1),.clk(gclk));
	jdff dff_B_wuSjxGMb3_1(.din(w_dff_B_9wQpPHUb9_1),.dout(w_dff_B_wuSjxGMb3_1),.clk(gclk));
	jdff dff_B_aUzpgTQD2_1(.din(n150),.dout(w_dff_B_aUzpgTQD2_1),.clk(gclk));
	jdff dff_B_saO59Fmz8_1(.din(w_dff_B_aUzpgTQD2_1),.dout(w_dff_B_saO59Fmz8_1),.clk(gclk));
	jdff dff_A_Tqry09g46_0(.dout(w_G97_4[0]),.din(w_dff_A_Tqry09g46_0),.clk(gclk));
	jdff dff_A_ZSDab67S5_0(.dout(w_dff_A_Tqry09g46_0),.din(w_dff_A_ZSDab67S5_0),.clk(gclk));
	jdff dff_A_vV64sr3w8_0(.dout(w_dff_A_ZSDab67S5_0),.din(w_dff_A_vV64sr3w8_0),.clk(gclk));
	jdff dff_A_0DUZvNbg9_0(.dout(w_dff_A_vV64sr3w8_0),.din(w_dff_A_0DUZvNbg9_0),.clk(gclk));
	jdff dff_A_XTGG9y8x7_2(.dout(w_G97_4[2]),.din(w_dff_A_XTGG9y8x7_2),.clk(gclk));
	jdff dff_A_qP9inbNF1_2(.dout(w_G97_1[2]),.din(w_dff_A_qP9inbNF1_2),.clk(gclk));
	jdff dff_A_9ud1mzav9_2(.dout(w_dff_A_qP9inbNF1_2),.din(w_dff_A_9ud1mzav9_2),.clk(gclk));
	jdff dff_A_Xa25Z2Up3_2(.dout(w_dff_A_9ud1mzav9_2),.din(w_dff_A_Xa25Z2Up3_2),.clk(gclk));
	jdff dff_A_cSHrJns84_1(.dout(w_G97_0[1]),.din(w_dff_A_cSHrJns84_1),.clk(gclk));
	jdff dff_A_jSiJcNSL3_1(.dout(w_dff_A_cSHrJns84_1),.din(w_dff_A_jSiJcNSL3_1),.clk(gclk));
	jdff dff_A_HDfvmbSy5_1(.dout(w_dff_A_jSiJcNSL3_1),.din(w_dff_A_HDfvmbSy5_1),.clk(gclk));
	jdff dff_A_VwcYS28T1_2(.dout(w_n153_2[2]),.din(w_dff_A_VwcYS28T1_2),.clk(gclk));
	jdff dff_A_OdCd76oN4_2(.dout(w_dff_A_VwcYS28T1_2),.din(w_dff_A_OdCd76oN4_2),.clk(gclk));
	jdff dff_A_skgac2vk4_2(.dout(w_dff_A_OdCd76oN4_2),.din(w_dff_A_skgac2vk4_2),.clk(gclk));
	jdff dff_A_6aYC8LGG7_2(.dout(w_n153_0[2]),.din(w_dff_A_6aYC8LGG7_2),.clk(gclk));
	jdff dff_A_WntodRxc7_2(.dout(w_dff_A_6aYC8LGG7_2),.din(w_dff_A_WntodRxc7_2),.clk(gclk));
	jdff dff_A_An85pV1v5_2(.dout(w_dff_A_WntodRxc7_2),.din(w_dff_A_An85pV1v5_2),.clk(gclk));
	jdff dff_A_DytGePDb4_1(.dout(w_n152_0[1]),.din(w_dff_A_DytGePDb4_1),.clk(gclk));
	jdff dff_A_6WaQmQZx7_0(.dout(w_G283_3[0]),.din(w_dff_A_6WaQmQZx7_0),.clk(gclk));
	jdff dff_A_Fha37d1V2_0(.dout(w_dff_A_6WaQmQZx7_0),.din(w_dff_A_Fha37d1V2_0),.clk(gclk));
	jdff dff_A_OgmqfJ9Y9_0(.dout(w_dff_A_Fha37d1V2_0),.din(w_dff_A_OgmqfJ9Y9_0),.clk(gclk));
	jdff dff_A_zBAtWpy87_1(.dout(w_G283_3[1]),.din(w_dff_A_zBAtWpy87_1),.clk(gclk));
	jdff dff_A_t7ycE5da5_1(.dout(w_dff_A_zBAtWpy87_1),.din(w_dff_A_t7ycE5da5_1),.clk(gclk));
	jdff dff_A_japh8m6f2_1(.dout(w_dff_A_t7ycE5da5_1),.din(w_dff_A_japh8m6f2_1),.clk(gclk));
	jdff dff_A_BNN3rqAD9_0(.dout(w_G283_0[0]),.din(w_dff_A_BNN3rqAD9_0),.clk(gclk));
	jdff dff_A_kWk1fZDO7_0(.dout(w_dff_A_BNN3rqAD9_0),.din(w_dff_A_kWk1fZDO7_0),.clk(gclk));
	jdff dff_A_Z4gpDrdV4_0(.dout(w_dff_A_kWk1fZDO7_0),.din(w_dff_A_Z4gpDrdV4_0),.clk(gclk));
	jdff dff_A_Y6N4dNAR7_1(.dout(w_G283_0[1]),.din(w_dff_A_Y6N4dNAR7_1),.clk(gclk));
	jdff dff_A_9WKlBnfF9_1(.dout(w_dff_A_Y6N4dNAR7_1),.din(w_dff_A_9WKlBnfF9_1),.clk(gclk));
	jdff dff_A_6Nv8glqm8_1(.dout(w_dff_A_9WKlBnfF9_1),.din(w_dff_A_6Nv8glqm8_1),.clk(gclk));
	jdff dff_A_Ytt10nUx2_0(.dout(w_n151_4[0]),.din(w_dff_A_Ytt10nUx2_0),.clk(gclk));
	jdff dff_A_kOWn8T0U2_0(.dout(w_n151_1[0]),.din(w_dff_A_kOWn8T0U2_0),.clk(gclk));
	jdff dff_A_Y7vdIFIK6_1(.dout(w_n151_1[1]),.din(w_dff_A_Y7vdIFIK6_1),.clk(gclk));
	jdff dff_A_si3cUgSf0_0(.dout(w_G116_4[0]),.din(w_dff_A_si3cUgSf0_0),.clk(gclk));
	jdff dff_A_A4rf8QyB8_0(.dout(w_dff_A_si3cUgSf0_0),.din(w_dff_A_A4rf8QyB8_0),.clk(gclk));
	jdff dff_A_FEZpIib27_0(.dout(w_dff_A_A4rf8QyB8_0),.din(w_dff_A_FEZpIib27_0),.clk(gclk));
	jdff dff_B_jviK8z9P0_0(.din(n147),.dout(w_dff_B_jviK8z9P0_0),.clk(gclk));
	jdff dff_A_qTqAcC4z7_2(.dout(w_G20_6[2]),.din(w_dff_A_qTqAcC4z7_2),.clk(gclk));
	jdff dff_A_xBj5cX0X9_2(.dout(w_dff_A_qTqAcC4z7_2),.din(w_dff_A_xBj5cX0X9_2),.clk(gclk));
	jdff dff_A_PneygkG64_0(.dout(w_G20_1[0]),.din(w_dff_A_PneygkG64_0),.clk(gclk));
	jdff dff_A_RsTLAMxA9_1(.dout(w_G20_1[1]),.din(w_dff_A_RsTLAMxA9_1),.clk(gclk));
	jdff dff_A_L8RaPNdA8_0(.dout(w_n142_0[0]),.din(w_dff_A_L8RaPNdA8_0),.clk(gclk));
	jdff dff_A_OTVES8wK6_1(.dout(w_G33_3[1]),.din(w_dff_A_OTVES8wK6_1),.clk(gclk));
	jdff dff_A_Gvez15wZ2_2(.dout(w_G33_3[2]),.din(w_dff_A_Gvez15wZ2_2),.clk(gclk));
	jdff dff_A_ym6S5rR28_2(.dout(w_dff_A_Gvez15wZ2_2),.din(w_dff_A_ym6S5rR28_2),.clk(gclk));
	jdff dff_A_0lhVdymT3_2(.dout(w_dff_A_ym6S5rR28_2),.din(w_dff_A_0lhVdymT3_2),.clk(gclk));
	jdff dff_A_L7ZuTVMZ3_2(.dout(w_dff_A_0lhVdymT3_2),.din(w_dff_A_L7ZuTVMZ3_2),.clk(gclk));
	jdff dff_A_1AiiHIgY1_0(.dout(w_G33_0[0]),.din(w_dff_A_1AiiHIgY1_0),.clk(gclk));
	jdff dff_A_R7XW4HVH1_1(.dout(w_n140_1[1]),.din(w_dff_A_R7XW4HVH1_1),.clk(gclk));
	jdff dff_A_MlDAFvhn9_2(.dout(w_n140_1[2]),.din(w_dff_A_MlDAFvhn9_2),.clk(gclk));
	jdff dff_A_DzYTHKxa5_0(.dout(w_G13_1[0]),.din(w_dff_A_DzYTHKxa5_0),.clk(gclk));
	jdff dff_A_QxIYbuhb7_0(.dout(w_dff_A_DzYTHKxa5_0),.din(w_dff_A_QxIYbuhb7_0),.clk(gclk));
	jdff dff_A_QvlrAJJ99_1(.dout(w_G13_1[1]),.din(w_dff_A_QvlrAJJ99_1),.clk(gclk));
	jdff dff_A_kfyvtHr53_0(.dout(w_n112_1[0]),.din(w_dff_A_kfyvtHr53_0),.clk(gclk));
	jdff dff_A_J6dLmODg2_0(.dout(w_dff_A_kfyvtHr53_0),.din(w_dff_A_J6dLmODg2_0),.clk(gclk));
	jdff dff_A_JBh6SnlL3_1(.dout(w_n112_1[1]),.din(w_dff_A_JBh6SnlL3_1),.clk(gclk));
	jdff dff_A_wQiY8xZZ6_1(.dout(w_dff_A_JBh6SnlL3_1),.din(w_dff_A_wQiY8xZZ6_1),.clk(gclk));
	jdff dff_A_6jGnGUuh6_1(.dout(w_n112_0[1]),.din(w_dff_A_6jGnGUuh6_1),.clk(gclk));
	jdff dff_A_4AZOtCLP3_1(.dout(w_dff_A_6jGnGUuh6_1),.din(w_dff_A_4AZOtCLP3_1),.clk(gclk));
	jdff dff_A_P28HTxyQ2_1(.dout(w_dff_A_4AZOtCLP3_1),.din(w_dff_A_P28HTxyQ2_1),.clk(gclk));
	jdff dff_A_ueunDt7R6_2(.dout(w_n112_0[2]),.din(w_dff_A_ueunDt7R6_2),.clk(gclk));
	jdff dff_A_iOyGJcSv8_2(.dout(w_dff_A_ueunDt7R6_2),.din(w_dff_A_iOyGJcSv8_2),.clk(gclk));
	jdff dff_A_AYHq6CK15_0(.dout(w_G116_5[0]),.din(w_dff_A_AYHq6CK15_0),.clk(gclk));
	jdff dff_A_uFxFIb6L8_2(.dout(w_G116_1[2]),.din(w_dff_A_uFxFIb6L8_2),.clk(gclk));
	jdff dff_A_vFeSx1O01_2(.dout(w_dff_A_uFxFIb6L8_2),.din(w_dff_A_vFeSx1O01_2),.clk(gclk));
	jdff dff_A_7r9CT32r7_2(.dout(w_dff_A_vFeSx1O01_2),.din(w_dff_A_7r9CT32r7_2),.clk(gclk));
	jdff dff_A_HIJ7ju3t0_1(.dout(w_G116_0[1]),.din(w_dff_A_HIJ7ju3t0_1),.clk(gclk));
	jdff dff_A_qs52CrPS9_1(.dout(w_dff_A_HIJ7ju3t0_1),.din(w_dff_A_qs52CrPS9_1),.clk(gclk));
	jdff dff_A_Nsl13udB4_1(.dout(w_dff_A_qs52CrPS9_1),.din(w_dff_A_Nsl13udB4_1),.clk(gclk));
	jdff dff_A_UT885Zls5_2(.dout(w_G116_0[2]),.din(w_dff_A_UT885Zls5_2),.clk(gclk));
	jdff dff_A_HWqYXczf8_2(.dout(w_dff_A_UT885Zls5_2),.din(w_dff_A_HWqYXczf8_2),.clk(gclk));
	jdff dff_A_399Kevc33_2(.dout(w_dff_A_HWqYXczf8_2),.din(w_dff_A_399Kevc33_2),.clk(gclk));
	jdff dff_A_hFnmCp9o6_1(.dout(w_G330_0[1]),.din(w_dff_A_hFnmCp9o6_1),.clk(gclk));
	jdff dff_A_yhCoLZdL9_1(.dout(w_dff_A_hFnmCp9o6_1),.din(w_dff_A_yhCoLZdL9_1),.clk(gclk));
	jdff dff_B_HpxBCUdY2_3(.din(G330),.dout(w_dff_B_HpxBCUdY2_3),.clk(gclk));
	jdff dff_B_VuWeNsBL3_3(.din(w_dff_B_HpxBCUdY2_3),.dout(w_dff_B_VuWeNsBL3_3),.clk(gclk));
	jdff dff_B_hkgUZhFI7_3(.din(w_dff_B_VuWeNsBL3_3),.dout(w_dff_B_hkgUZhFI7_3),.clk(gclk));
	jdff dff_B_LS61dqx66_3(.din(w_dff_B_hkgUZhFI7_3),.dout(w_dff_B_LS61dqx66_3),.clk(gclk));
	jdff dff_B_tXsgcTSw2_3(.din(w_dff_B_LS61dqx66_3),.dout(w_dff_B_tXsgcTSw2_3),.clk(gclk));
	jdff dff_B_BwWvCrM99_3(.din(w_dff_B_tXsgcTSw2_3),.dout(w_dff_B_BwWvCrM99_3),.clk(gclk));
	jdff dff_B_YlrImd1e3_3(.din(w_dff_B_BwWvCrM99_3),.dout(w_dff_B_YlrImd1e3_3),.clk(gclk));
	jdff dff_B_qR0nOs1x3_3(.din(w_dff_B_YlrImd1e3_3),.dout(w_dff_B_qR0nOs1x3_3),.clk(gclk));
	jdff dff_B_OEg4m9xA1_3(.din(w_dff_B_qR0nOs1x3_3),.dout(w_dff_B_OEg4m9xA1_3),.clk(gclk));
	jdff dff_B_ZhZ4D0zS4_3(.din(w_dff_B_OEg4m9xA1_3),.dout(w_dff_B_ZhZ4D0zS4_3),.clk(gclk));
	jdff dff_B_0dXxVJuE3_3(.din(w_dff_B_ZhZ4D0zS4_3),.dout(w_dff_B_0dXxVJuE3_3),.clk(gclk));
	jdff dff_B_hWTaQiHW1_3(.din(w_dff_B_0dXxVJuE3_3),.dout(w_dff_B_hWTaQiHW1_3),.clk(gclk));
	jdff dff_A_wq17tauH8_1(.dout(w_n575_0[1]),.din(w_dff_A_wq17tauH8_1),.clk(gclk));
	jdff dff_A_odPI4HrQ6_1(.dout(w_dff_A_wq17tauH8_1),.din(w_dff_A_odPI4HrQ6_1),.clk(gclk));
	jdff dff_A_eq5YLhq75_1(.dout(w_dff_A_odPI4HrQ6_1),.din(w_dff_A_eq5YLhq75_1),.clk(gclk));
	jdff dff_A_o6mjsxuy0_1(.dout(w_dff_A_eq5YLhq75_1),.din(w_dff_A_o6mjsxuy0_1),.clk(gclk));
	jdff dff_A_8QnkC18e8_1(.dout(w_dff_A_o6mjsxuy0_1),.din(w_dff_A_8QnkC18e8_1),.clk(gclk));
	jdff dff_A_ChNSborp8_1(.dout(w_dff_A_8QnkC18e8_1),.din(w_dff_A_ChNSborp8_1),.clk(gclk));
	jdff dff_A_G3muGB1A2_1(.dout(w_dff_A_ChNSborp8_1),.din(w_dff_A_G3muGB1A2_1),.clk(gclk));
	jdff dff_A_PJflLZpI6_1(.dout(w_dff_A_G3muGB1A2_1),.din(w_dff_A_PJflLZpI6_1),.clk(gclk));
	jdff dff_A_LK58E5yq2_1(.dout(w_dff_A_PJflLZpI6_1),.din(w_dff_A_LK58E5yq2_1),.clk(gclk));
	jdff dff_A_HcC95OHT5_2(.dout(w_n575_0[2]),.din(w_dff_A_HcC95OHT5_2),.clk(gclk));
	jdff dff_A_bRIPMCeQ2_2(.dout(w_dff_A_HcC95OHT5_2),.din(w_dff_A_bRIPMCeQ2_2),.clk(gclk));
	jdff dff_A_BSCoWUSj4_2(.dout(w_dff_A_bRIPMCeQ2_2),.din(w_dff_A_BSCoWUSj4_2),.clk(gclk));
	jdff dff_A_2i7L6yMM1_2(.dout(w_dff_A_BSCoWUSj4_2),.din(w_dff_A_2i7L6yMM1_2),.clk(gclk));
	jdff dff_A_LkQJ7Yen8_2(.dout(w_dff_A_2i7L6yMM1_2),.din(w_dff_A_LkQJ7Yen8_2),.clk(gclk));
	jdff dff_A_4bcMFsIz0_2(.dout(w_dff_A_LkQJ7Yen8_2),.din(w_dff_A_4bcMFsIz0_2),.clk(gclk));
	jdff dff_A_FwqPq3SO6_0(.dout(w_n574_4[0]),.din(w_dff_A_FwqPq3SO6_0),.clk(gclk));
	jdff dff_A_MIMMLezA6_0(.dout(w_dff_A_FwqPq3SO6_0),.din(w_dff_A_MIMMLezA6_0),.clk(gclk));
	jdff dff_A_n4OUThTi6_0(.dout(w_dff_A_MIMMLezA6_0),.din(w_dff_A_n4OUThTi6_0),.clk(gclk));
	jdff dff_A_8ENOy4QH8_0(.dout(w_dff_A_n4OUThTi6_0),.din(w_dff_A_8ENOy4QH8_0),.clk(gclk));
	jdff dff_A_xbKGV8NW7_0(.dout(w_dff_A_8ENOy4QH8_0),.din(w_dff_A_xbKGV8NW7_0),.clk(gclk));
	jdff dff_A_U62r0qJs5_0(.dout(w_dff_A_xbKGV8NW7_0),.din(w_dff_A_U62r0qJs5_0),.clk(gclk));
	jdff dff_A_2xtU7aLo1_0(.dout(w_dff_A_U62r0qJs5_0),.din(w_dff_A_2xtU7aLo1_0),.clk(gclk));
	jdff dff_A_kMWFvHvv5_0(.dout(w_dff_A_2xtU7aLo1_0),.din(w_dff_A_kMWFvHvv5_0),.clk(gclk));
	jdff dff_A_6HVwM8yu0_1(.dout(w_n574_1[1]),.din(w_dff_A_6HVwM8yu0_1),.clk(gclk));
	jdff dff_A_3dyDH51V9_1(.dout(w_dff_A_6HVwM8yu0_1),.din(w_dff_A_3dyDH51V9_1),.clk(gclk));
	jdff dff_A_NrhTesYA0_1(.dout(w_dff_A_3dyDH51V9_1),.din(w_dff_A_NrhTesYA0_1),.clk(gclk));
	jdff dff_A_T7h3xX7x7_1(.dout(w_dff_A_NrhTesYA0_1),.din(w_dff_A_T7h3xX7x7_1),.clk(gclk));
	jdff dff_A_qUZtGVCA1_1(.dout(w_dff_A_T7h3xX7x7_1),.din(w_dff_A_qUZtGVCA1_1),.clk(gclk));
	jdff dff_A_EI3WYb5P3_1(.dout(w_dff_A_qUZtGVCA1_1),.din(w_dff_A_EI3WYb5P3_1),.clk(gclk));
	jdff dff_A_j6WSIunK5_2(.dout(w_n574_1[2]),.din(w_dff_A_j6WSIunK5_2),.clk(gclk));
	jdff dff_A_1ySQcKkI4_2(.dout(w_dff_A_j6WSIunK5_2),.din(w_dff_A_1ySQcKkI4_2),.clk(gclk));
	jdff dff_A_xlQbREQG7_2(.dout(w_dff_A_1ySQcKkI4_2),.din(w_dff_A_xlQbREQG7_2),.clk(gclk));
	jdff dff_A_wT7z0BGQ2_2(.dout(w_dff_A_xlQbREQG7_2),.din(w_dff_A_wT7z0BGQ2_2),.clk(gclk));
	jdff dff_A_LshbYJWD0_2(.dout(w_dff_A_wT7z0BGQ2_2),.din(w_dff_A_LshbYJWD0_2),.clk(gclk));
	jdff dff_A_dsPI1f6d0_2(.dout(w_dff_A_LshbYJWD0_2),.din(w_dff_A_dsPI1f6d0_2),.clk(gclk));
	jdff dff_A_CjqlpFYP9_2(.dout(w_dff_A_dsPI1f6d0_2),.din(w_dff_A_CjqlpFYP9_2),.clk(gclk));
	jdff dff_A_bull1NsZ7_2(.dout(w_dff_A_CjqlpFYP9_2),.din(w_dff_A_bull1NsZ7_2),.clk(gclk));
	jdff dff_A_bGLM5hDN8_2(.dout(w_dff_A_bull1NsZ7_2),.din(w_dff_A_bGLM5hDN8_2),.clk(gclk));
	jdff dff_A_XhX0mBD51_2(.dout(w_dff_A_bGLM5hDN8_2),.din(w_dff_A_XhX0mBD51_2),.clk(gclk));
	jdff dff_A_IBtBOk9U7_2(.dout(w_dff_A_XhX0mBD51_2),.din(w_dff_A_IBtBOk9U7_2),.clk(gclk));
	jdff dff_A_O9lR93Wb3_2(.dout(w_dff_A_IBtBOk9U7_2),.din(w_dff_A_O9lR93Wb3_2),.clk(gclk));
	jdff dff_A_Z1wyCwtZ5_2(.dout(w_dff_A_O9lR93Wb3_2),.din(w_dff_A_Z1wyCwtZ5_2),.clk(gclk));
	jdff dff_A_1AnaTcwN1_2(.dout(w_dff_A_Z1wyCwtZ5_2),.din(w_dff_A_1AnaTcwN1_2),.clk(gclk));
	jdff dff_A_rntIr00f0_2(.dout(w_n574_0[2]),.din(w_dff_A_rntIr00f0_2),.clk(gclk));
	jdff dff_A_Jf5yIcVn3_0(.dout(w_n573_1[0]),.din(w_dff_A_Jf5yIcVn3_0),.clk(gclk));
	jdff dff_A_wb0wzZSE9_0(.dout(w_dff_A_Jf5yIcVn3_0),.din(w_dff_A_wb0wzZSE9_0),.clk(gclk));
	jdff dff_A_jKgZNIMu7_0(.dout(w_dff_A_wb0wzZSE9_0),.din(w_dff_A_jKgZNIMu7_0),.clk(gclk));
	jdff dff_A_xDPBuZb37_0(.dout(w_dff_A_jKgZNIMu7_0),.din(w_dff_A_xDPBuZb37_0),.clk(gclk));
	jdff dff_A_ZISYk3go7_0(.dout(w_dff_A_xDPBuZb37_0),.din(w_dff_A_ZISYk3go7_0),.clk(gclk));
	jdff dff_A_0ZTjpXni3_0(.dout(w_dff_A_ZISYk3go7_0),.din(w_dff_A_0ZTjpXni3_0),.clk(gclk));
	jdff dff_A_8lkKjvOA5_0(.dout(w_dff_A_0ZTjpXni3_0),.din(w_dff_A_8lkKjvOA5_0),.clk(gclk));
	jdff dff_A_xnnJk6NX3_0(.dout(w_dff_A_8lkKjvOA5_0),.din(w_dff_A_xnnJk6NX3_0),.clk(gclk));
	jdff dff_A_F8Wh3OG13_0(.dout(w_dff_A_xnnJk6NX3_0),.din(w_dff_A_F8Wh3OG13_0),.clk(gclk));
	jdff dff_A_O9Hvuued7_0(.dout(w_dff_A_F8Wh3OG13_0),.din(w_dff_A_O9Hvuued7_0),.clk(gclk));
	jdff dff_A_qLPUx0zY9_0(.dout(w_dff_A_O9Hvuued7_0),.din(w_dff_A_qLPUx0zY9_0),.clk(gclk));
	jdff dff_A_JAjcmLmg2_0(.dout(w_dff_A_qLPUx0zY9_0),.din(w_dff_A_JAjcmLmg2_0),.clk(gclk));
	jdff dff_A_UdbYpxOn5_0(.dout(w_dff_A_JAjcmLmg2_0),.din(w_dff_A_UdbYpxOn5_0),.clk(gclk));
	jdff dff_A_jR0uzgHd6_1(.dout(w_n573_1[1]),.din(w_dff_A_jR0uzgHd6_1),.clk(gclk));
	jdff dff_A_fP9zkEzN6_1(.dout(w_dff_A_jR0uzgHd6_1),.din(w_dff_A_fP9zkEzN6_1),.clk(gclk));
	jdff dff_A_28pLuohY1_1(.dout(w_dff_A_fP9zkEzN6_1),.din(w_dff_A_28pLuohY1_1),.clk(gclk));
	jdff dff_A_Z6I2cObm2_1(.dout(w_dff_A_28pLuohY1_1),.din(w_dff_A_Z6I2cObm2_1),.clk(gclk));
	jdff dff_A_qNisaUU57_1(.dout(w_dff_A_Z6I2cObm2_1),.din(w_dff_A_qNisaUU57_1),.clk(gclk));
	jdff dff_A_Q5cVGGPa3_1(.dout(w_dff_A_qNisaUU57_1),.din(w_dff_A_Q5cVGGPa3_1),.clk(gclk));
	jdff dff_A_8X2wSEvH9_1(.dout(w_dff_A_Q5cVGGPa3_1),.din(w_dff_A_8X2wSEvH9_1),.clk(gclk));
	jdff dff_A_LSBen3VT6_1(.dout(w_dff_A_8X2wSEvH9_1),.din(w_dff_A_LSBen3VT6_1),.clk(gclk));
	jdff dff_A_IKY4WGqU3_1(.dout(w_dff_A_LSBen3VT6_1),.din(w_dff_A_IKY4WGqU3_1),.clk(gclk));
	jdff dff_A_eZTnycEY0_1(.dout(w_dff_A_IKY4WGqU3_1),.din(w_dff_A_eZTnycEY0_1),.clk(gclk));
	jdff dff_A_PwS40WEr4_1(.dout(w_dff_A_eZTnycEY0_1),.din(w_dff_A_PwS40WEr4_1),.clk(gclk));
	jdff dff_A_suiCb5en8_1(.dout(w_dff_A_PwS40WEr4_1),.din(w_dff_A_suiCb5en8_1),.clk(gclk));
	jdff dff_A_PKBNQTrc3_1(.dout(w_n573_0[1]),.din(w_dff_A_PKBNQTrc3_1),.clk(gclk));
	jdff dff_A_Zj2o4NDI8_1(.dout(w_dff_A_PKBNQTrc3_1),.din(w_dff_A_Zj2o4NDI8_1),.clk(gclk));
	jdff dff_A_LSVW6T4U5_1(.dout(w_dff_A_Zj2o4NDI8_1),.din(w_dff_A_LSVW6T4U5_1),.clk(gclk));
	jdff dff_A_QMz9OikZ6_1(.dout(w_dff_A_LSVW6T4U5_1),.din(w_dff_A_QMz9OikZ6_1),.clk(gclk));
	jdff dff_A_KWPFfSFI3_1(.dout(w_dff_A_QMz9OikZ6_1),.din(w_dff_A_KWPFfSFI3_1),.clk(gclk));
	jdff dff_A_sepS8pSO6_1(.dout(w_dff_A_KWPFfSFI3_1),.din(w_dff_A_sepS8pSO6_1),.clk(gclk));
	jdff dff_A_NaxjPiNG0_1(.dout(w_dff_A_sepS8pSO6_1),.din(w_dff_A_NaxjPiNG0_1),.clk(gclk));
	jdff dff_A_qtlOBJgE6_1(.dout(w_dff_A_NaxjPiNG0_1),.din(w_dff_A_qtlOBJgE6_1),.clk(gclk));
	jdff dff_A_rYEg0xQW4_1(.dout(w_dff_A_qtlOBJgE6_1),.din(w_dff_A_rYEg0xQW4_1),.clk(gclk));
	jdff dff_A_CQ9if87m6_1(.dout(w_dff_A_rYEg0xQW4_1),.din(w_dff_A_CQ9if87m6_1),.clk(gclk));
	jdff dff_A_DervnNSt4_1(.dout(w_dff_A_CQ9if87m6_1),.din(w_dff_A_DervnNSt4_1),.clk(gclk));
	jdff dff_A_GFjYngmS2_1(.dout(w_dff_A_DervnNSt4_1),.din(w_dff_A_GFjYngmS2_1),.clk(gclk));
	jdff dff_A_KCXX7tRl7_1(.dout(w_dff_A_GFjYngmS2_1),.din(w_dff_A_KCXX7tRl7_1),.clk(gclk));
	jdff dff_A_6P2bOYnB9_1(.dout(w_dff_A_KCXX7tRl7_1),.din(w_dff_A_6P2bOYnB9_1),.clk(gclk));
	jdff dff_A_C8D6vxpD9_2(.dout(w_n573_0[2]),.din(w_dff_A_C8D6vxpD9_2),.clk(gclk));
	jdff dff_A_Vt8mm9Rn7_2(.dout(w_dff_A_C8D6vxpD9_2),.din(w_dff_A_Vt8mm9Rn7_2),.clk(gclk));
	jdff dff_A_v9RSeGlc2_2(.dout(w_dff_A_Vt8mm9Rn7_2),.din(w_dff_A_v9RSeGlc2_2),.clk(gclk));
	jdff dff_A_8AiQklu46_2(.dout(w_dff_A_v9RSeGlc2_2),.din(w_dff_A_8AiQklu46_2),.clk(gclk));
	jdff dff_A_duFtBtYo7_2(.dout(w_dff_A_8AiQklu46_2),.din(w_dff_A_duFtBtYo7_2),.clk(gclk));
	jdff dff_A_jyxrqg485_2(.dout(w_dff_A_duFtBtYo7_2),.din(w_dff_A_jyxrqg485_2),.clk(gclk));
	jdff dff_A_HHn99T6W3_2(.dout(w_dff_A_jyxrqg485_2),.din(w_dff_A_HHn99T6W3_2),.clk(gclk));
	jdff dff_A_rBNz9LNg5_2(.dout(w_dff_A_HHn99T6W3_2),.din(w_dff_A_rBNz9LNg5_2),.clk(gclk));
	jdff dff_A_WrHiGEOx6_2(.dout(w_dff_A_rBNz9LNg5_2),.din(w_dff_A_WrHiGEOx6_2),.clk(gclk));
	jdff dff_A_JV2OWS1j2_2(.dout(w_dff_A_WrHiGEOx6_2),.din(w_dff_A_JV2OWS1j2_2),.clk(gclk));
	jdff dff_A_KPaBokur1_2(.dout(w_dff_A_JV2OWS1j2_2),.din(w_dff_A_KPaBokur1_2),.clk(gclk));
	jdff dff_A_QtGdZ2P71_2(.dout(w_dff_A_KPaBokur1_2),.din(w_dff_A_QtGdZ2P71_2),.clk(gclk));
	jdff dff_A_QsyBmHKn1_2(.dout(w_dff_A_QtGdZ2P71_2),.din(w_dff_A_QsyBmHKn1_2),.clk(gclk));
	jdff dff_A_oF0G75GT9_2(.dout(w_dff_A_QsyBmHKn1_2),.din(w_dff_A_oF0G75GT9_2),.clk(gclk));
	jdff dff_B_TbB8LnBB0_3(.din(n573),.dout(w_dff_B_TbB8LnBB0_3),.clk(gclk));
	jdff dff_B_Sj4KfGWI2_0(.din(n571),.dout(w_dff_B_Sj4KfGWI2_0),.clk(gclk));
	jdff dff_A_NINlQxwq3_1(.dout(w_G45_0[1]),.din(w_dff_A_NINlQxwq3_1),.clk(gclk));
	jdff dff_A_NwbguLHv3_1(.dout(w_dff_A_NINlQxwq3_1),.din(w_dff_A_NwbguLHv3_1),.clk(gclk));
	jdff dff_A_kC2B1HrP3_1(.dout(w_dff_A_NwbguLHv3_1),.din(w_dff_A_kC2B1HrP3_1),.clk(gclk));
	jdff dff_A_S0swvLc28_0(.dout(w_G1_1[0]),.din(w_dff_A_S0swvLc28_0),.clk(gclk));
	jdff dff_A_V2sEVFqm3_0(.dout(w_dff_A_S0swvLc28_0),.din(w_dff_A_V2sEVFqm3_0),.clk(gclk));
	jdff dff_A_4DbpvSP54_0(.dout(w_n107_0[0]),.din(w_dff_A_4DbpvSP54_0),.clk(gclk));
	jdff dff_A_jyntGYM43_0(.dout(w_n564_1[0]),.din(w_dff_A_jyntGYM43_0),.clk(gclk));
	jdff dff_A_n5LQbdfq2_0(.dout(w_dff_A_jyntGYM43_0),.din(w_dff_A_n5LQbdfq2_0),.clk(gclk));
	jdff dff_A_c25JhkaE2_0(.dout(w_dff_A_n5LQbdfq2_0),.din(w_dff_A_c25JhkaE2_0),.clk(gclk));
	jdff dff_A_vVl1w5EO7_0(.dout(w_dff_A_c25JhkaE2_0),.din(w_dff_A_vVl1w5EO7_0),.clk(gclk));
	jdff dff_A_ZxSMuo5S0_0(.dout(w_dff_A_vVl1w5EO7_0),.din(w_dff_A_ZxSMuo5S0_0),.clk(gclk));
	jdff dff_A_GpSmMdZv1_0(.dout(w_dff_A_ZxSMuo5S0_0),.din(w_dff_A_GpSmMdZv1_0),.clk(gclk));
	jdff dff_A_T185TyPJ9_0(.dout(w_dff_A_GpSmMdZv1_0),.din(w_dff_A_T185TyPJ9_0),.clk(gclk));
	jdff dff_A_6ThDI6n79_0(.dout(w_dff_A_T185TyPJ9_0),.din(w_dff_A_6ThDI6n79_0),.clk(gclk));
	jdff dff_A_2Z5DWBrz8_0(.dout(w_dff_A_6ThDI6n79_0),.din(w_dff_A_2Z5DWBrz8_0),.clk(gclk));
	jdff dff_A_TUeKvJNr8_0(.dout(w_dff_A_2Z5DWBrz8_0),.din(w_dff_A_TUeKvJNr8_0),.clk(gclk));
	jdff dff_A_HHOYeyMC1_0(.dout(w_dff_A_TUeKvJNr8_0),.din(w_dff_A_HHOYeyMC1_0),.clk(gclk));
	jdff dff_A_qIOZQG3K4_0(.dout(w_dff_A_HHOYeyMC1_0),.din(w_dff_A_qIOZQG3K4_0),.clk(gclk));
	jdff dff_A_yZfjNgZR7_0(.dout(w_dff_A_qIOZQG3K4_0),.din(w_dff_A_yZfjNgZR7_0),.clk(gclk));
	jdff dff_A_k1RkcxC58_1(.dout(w_n564_0[1]),.din(w_dff_A_k1RkcxC58_1),.clk(gclk));
	jdff dff_A_5iromuUB8_1(.dout(w_dff_A_k1RkcxC58_1),.din(w_dff_A_5iromuUB8_1),.clk(gclk));
	jdff dff_A_Eplzsdje0_1(.dout(w_dff_A_5iromuUB8_1),.din(w_dff_A_Eplzsdje0_1),.clk(gclk));
	jdff dff_A_D6wIkQq63_1(.dout(w_dff_A_Eplzsdje0_1),.din(w_dff_A_D6wIkQq63_1),.clk(gclk));
	jdff dff_A_dvKQ3T2E6_1(.dout(w_dff_A_D6wIkQq63_1),.din(w_dff_A_dvKQ3T2E6_1),.clk(gclk));
	jdff dff_A_3OvbDbXf2_1(.dout(w_dff_A_dvKQ3T2E6_1),.din(w_dff_A_3OvbDbXf2_1),.clk(gclk));
	jdff dff_A_0ku9FXH22_1(.dout(w_dff_A_3OvbDbXf2_1),.din(w_dff_A_0ku9FXH22_1),.clk(gclk));
	jdff dff_A_l9l4KR9Q6_1(.dout(w_dff_A_0ku9FXH22_1),.din(w_dff_A_l9l4KR9Q6_1),.clk(gclk));
	jdff dff_A_3C2r4G7N4_1(.dout(w_dff_A_l9l4KR9Q6_1),.din(w_dff_A_3C2r4G7N4_1),.clk(gclk));
	jdff dff_A_fgjGIS8G1_1(.dout(w_dff_A_3C2r4G7N4_1),.din(w_dff_A_fgjGIS8G1_1),.clk(gclk));
	jdff dff_A_zyTKAbuF7_1(.dout(w_dff_A_fgjGIS8G1_1),.din(w_dff_A_zyTKAbuF7_1),.clk(gclk));
	jdff dff_A_Bcu0894d5_1(.dout(w_dff_A_zyTKAbuF7_1),.din(w_dff_A_Bcu0894d5_1),.clk(gclk));
	jdff dff_A_QUJzufsG6_1(.dout(w_dff_A_Bcu0894d5_1),.din(w_dff_A_QUJzufsG6_1),.clk(gclk));
	jdff dff_A_oX0tGj6o2_1(.dout(w_dff_A_QUJzufsG6_1),.din(w_dff_A_oX0tGj6o2_1),.clk(gclk));
	jdff dff_A_Q3oncG7x6_2(.dout(w_n564_0[2]),.din(w_dff_A_Q3oncG7x6_2),.clk(gclk));
	jdff dff_A_WCpF15mb9_2(.dout(w_dff_A_Q3oncG7x6_2),.din(w_dff_A_WCpF15mb9_2),.clk(gclk));
	jdff dff_A_siDBz2mL7_2(.dout(w_dff_A_WCpF15mb9_2),.din(w_dff_A_siDBz2mL7_2),.clk(gclk));
	jdff dff_A_sibQJt2b4_2(.dout(w_dff_A_siDBz2mL7_2),.din(w_dff_A_sibQJt2b4_2),.clk(gclk));
	jdff dff_A_4hiLJwyr0_2(.dout(w_dff_A_sibQJt2b4_2),.din(w_dff_A_4hiLJwyr0_2),.clk(gclk));
	jdff dff_A_C1RyuKyV3_2(.dout(w_dff_A_4hiLJwyr0_2),.din(w_dff_A_C1RyuKyV3_2),.clk(gclk));
	jdff dff_A_rqsCTgRs1_2(.dout(w_dff_A_C1RyuKyV3_2),.din(w_dff_A_rqsCTgRs1_2),.clk(gclk));
	jdff dff_A_ShMnqvVX2_2(.dout(w_dff_A_rqsCTgRs1_2),.din(w_dff_A_ShMnqvVX2_2),.clk(gclk));
	jdff dff_A_38seGSQL2_2(.dout(w_dff_A_ShMnqvVX2_2),.din(w_dff_A_38seGSQL2_2),.clk(gclk));
	jdff dff_A_uRrYSUoL8_2(.dout(w_dff_A_38seGSQL2_2),.din(w_dff_A_uRrYSUoL8_2),.clk(gclk));
	jdff dff_A_21Sx4Cu24_2(.dout(w_dff_A_uRrYSUoL8_2),.din(w_dff_A_21Sx4Cu24_2),.clk(gclk));
	jdff dff_A_86ZLDcDD8_2(.dout(w_dff_A_21Sx4Cu24_2),.din(w_dff_A_86ZLDcDD8_2),.clk(gclk));
	jdff dff_A_A3K07Dcc6_2(.dout(w_dff_A_86ZLDcDD8_2),.din(w_dff_A_A3K07Dcc6_2),.clk(gclk));
	jdff dff_A_JmiBRX3w8_2(.dout(w_dff_A_A3K07Dcc6_2),.din(w_dff_A_JmiBRX3w8_2),.clk(gclk));
	jdff dff_A_4UcCWp4o5_0(.dout(w_n544_0[0]),.din(w_dff_A_4UcCWp4o5_0),.clk(gclk));
	jdff dff_A_KdbihPk27_0(.dout(w_dff_A_4UcCWp4o5_0),.din(w_dff_A_KdbihPk27_0),.clk(gclk));
	jdff dff_A_LqgYjfVH8_0(.dout(w_dff_A_KdbihPk27_0),.din(w_dff_A_LqgYjfVH8_0),.clk(gclk));
	jdff dff_A_9tX7QRMf3_0(.dout(w_dff_A_LqgYjfVH8_0),.din(w_dff_A_9tX7QRMf3_0),.clk(gclk));
	jdff dff_A_ChUb69I77_0(.dout(w_dff_A_9tX7QRMf3_0),.din(w_dff_A_ChUb69I77_0),.clk(gclk));
	jdff dff_A_ludhWNJg3_0(.dout(w_dff_A_ChUb69I77_0),.din(w_dff_A_ludhWNJg3_0),.clk(gclk));
	jdff dff_A_xtPru4fd9_0(.dout(w_dff_A_ludhWNJg3_0),.din(w_dff_A_xtPru4fd9_0),.clk(gclk));
	jdff dff_A_ywt0VBYD4_0(.dout(w_dff_A_xtPru4fd9_0),.din(w_dff_A_ywt0VBYD4_0),.clk(gclk));
	jdff dff_A_Huq76DsN7_0(.dout(w_dff_A_ywt0VBYD4_0),.din(w_dff_A_Huq76DsN7_0),.clk(gclk));
	jdff dff_A_vvTiUY1m5_0(.dout(w_dff_A_Huq76DsN7_0),.din(w_dff_A_vvTiUY1m5_0),.clk(gclk));
	jdff dff_A_ZOX8m0mE2_0(.dout(w_dff_A_vvTiUY1m5_0),.din(w_dff_A_ZOX8m0mE2_0),.clk(gclk));
	jdff dff_A_vMztpKWN1_0(.dout(w_dff_A_ZOX8m0mE2_0),.din(w_dff_A_vMztpKWN1_0),.clk(gclk));
	jdff dff_A_OKKURVhr0_0(.dout(w_dff_A_vMztpKWN1_0),.din(w_dff_A_OKKURVhr0_0),.clk(gclk));
	jdff dff_A_LPh7b7Kr5_0(.dout(w_G13_2[0]),.din(w_dff_A_LPh7b7Kr5_0),.clk(gclk));
	jdff dff_A_VEUEFbh67_1(.dout(w_G1_2[1]),.din(w_dff_A_VEUEFbh67_1),.clk(gclk));
	jdff dff_A_e87aQQn08_2(.dout(w_G1_0[2]),.din(w_dff_A_e87aQQn08_2),.clk(gclk));
	jdff dff_A_YvlyyIbO2_2(.dout(w_dff_A_e87aQQn08_2),.din(w_dff_A_YvlyyIbO2_2),.clk(gclk));
	jdff dff_A_6o6zkLh70_2(.dout(w_dff_A_YvlyyIbO2_2),.din(w_dff_A_6o6zkLh70_2),.clk(gclk));
	jdff dff_A_bfz3X9zz6_2(.dout(w_dff_A_6o6zkLh70_2),.din(w_dff_A_bfz3X9zz6_2),.clk(gclk));
	jdff dff_A_B7DRBSMe4_1(.dout(w_G20_7[1]),.din(w_dff_A_B7DRBSMe4_1),.clk(gclk));
	jdff dff_A_d7G0uZeB0_1(.dout(w_dff_A_B7DRBSMe4_1),.din(w_dff_A_d7G0uZeB0_1),.clk(gclk));
	jdff dff_A_B75geTHS5_1(.dout(w_G20_2[1]),.din(w_dff_A_B75geTHS5_1),.clk(gclk));
	jdff dff_A_97fE0sGQ5_1(.dout(w_n169_0[1]),.din(w_dff_A_97fE0sGQ5_1),.clk(gclk));
	jdff dff_A_YTabs3iB8_1(.dout(w_dff_A_97fE0sGQ5_1),.din(w_dff_A_YTabs3iB8_1),.clk(gclk));
	jdff dff_A_mmvX0yiL9_1(.dout(w_dff_A_YTabs3iB8_1),.din(w_dff_A_mmvX0yiL9_1),.clk(gclk));
	jdff dff_A_Jqsgc3Ot4_1(.dout(w_dff_A_mmvX0yiL9_1),.din(w_dff_A_Jqsgc3Ot4_1),.clk(gclk));
	jdff dff_A_eUpDNywa0_2(.dout(w_n169_0[2]),.din(w_dff_A_eUpDNywa0_2),.clk(gclk));
	jdff dff_A_WqVsXXA43_2(.dout(w_dff_A_eUpDNywa0_2),.din(w_dff_A_WqVsXXA43_2),.clk(gclk));
endmodule

