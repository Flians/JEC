/*

c880:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jcb: 122
	jdff: 823
	jand: 151

Summary:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jcb: 122
	jdff: 823
	jand: 151
*/

module c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n103;
	wire n104;
	wire n105;
	wire n107;
	wire n108;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n119;
	wire n120;
	wire n122;
	wire n123;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire [2:0] w_G1gat_0;
	wire [1:0] w_G1gat_1;
	wire [1:0] w_G8gat_0;
	wire [1:0] w_G13gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G17gat_1;
	wire [2:0] w_G17gat_2;
	wire [1:0] w_G26gat_0;
	wire [2:0] w_G29gat_0;
	wire [1:0] w_G36gat_0;
	wire [2:0] w_G42gat_0;
	wire [2:0] w_G42gat_1;
	wire [1:0] w_G42gat_2;
	wire [2:0] w_G51gat_0;
	wire [1:0] w_G51gat_1;
	wire [2:0] w_G55gat_0;
	wire [2:0] w_G59gat_0;
	wire [1:0] w_G59gat_1;
	wire [1:0] w_G68gat_0;
	wire [1:0] w_G75gat_0;
	wire [2:0] w_G80gat_0;
	wire [2:0] w_G91gat_0;
	wire [2:0] w_G96gat_0;
	wire [2:0] w_G101gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G111gat_0;
	wire [2:0] w_G116gat_0;
	wire [2:0] w_G121gat_0;
	wire [2:0] w_G126gat_0;
	wire [1:0] w_G130gat_0;
	wire [2:0] w_G138gat_0;
	wire [1:0] w_G138gat_1;
	wire [1:0] w_G143gat_0;
	wire [1:0] w_G146gat_0;
	wire [1:0] w_G149gat_0;
	wire [2:0] w_G153gat_0;
	wire [1:0] w_G156gat_0;
	wire [2:0] w_G159gat_0;
	wire [2:0] w_G159gat_1;
	wire [2:0] w_G165gat_0;
	wire [2:0] w_G165gat_1;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G177gat_0;
	wire [2:0] w_G177gat_1;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G183gat_1;
	wire [2:0] w_G189gat_0;
	wire [2:0] w_G189gat_1;
	wire [1:0] w_G189gat_2;
	wire [2:0] w_G195gat_0;
	wire [2:0] w_G195gat_1;
	wire [1:0] w_G195gat_2;
	wire [2:0] w_G201gat_0;
	wire [1:0] w_G201gat_1;
	wire [2:0] w_G210gat_0;
	wire [2:0] w_G210gat_1;
	wire [2:0] w_G210gat_2;
	wire [1:0] w_G210gat_3;
	wire [2:0] w_G219gat_0;
	wire [2:0] w_G219gat_1;
	wire [2:0] w_G219gat_2;
	wire [2:0] w_G219gat_3;
	wire [2:0] w_G228gat_0;
	wire [2:0] w_G228gat_1;
	wire [2:0] w_G228gat_2;
	wire [1:0] w_G228gat_3;
	wire [2:0] w_G237gat_0;
	wire [2:0] w_G237gat_1;
	wire [2:0] w_G237gat_2;
	wire [1:0] w_G237gat_3;
	wire [2:0] w_G246gat_0;
	wire [2:0] w_G246gat_1;
	wire [2:0] w_G246gat_2;
	wire [1:0] w_G246gat_3;
	wire [2:0] w_G255gat_0;
	wire [2:0] w_G261gat_0;
	wire [1:0] w_G268gat_0;
	wire [1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire [2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [1:0] w_n92_0;
	wire [1:0] w_n93_0;
	wire [2:0] w_n95_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n113_0;
	wire [2:0] w_n119_0;
	wire [1:0] w_n122_0;
	wire [1:0] w_n144_0;
	wire [1:0] w_n146_0;
	wire [2:0] w_n148_0;
	wire [2:0] w_n148_1;
	wire [1:0] w_n149_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n164_0;
	wire [2:0] w_n164_1;
	wire [2:0] w_n164_2;
	wire [1:0] w_n164_3;
	wire [1:0] w_n167_0;
	wire [1:0] w_n168_0;
	wire [2:0] w_n170_0;
	wire [1:0] w_n170_1;
	wire [1:0] w_n173_0;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n178_2;
	wire [1:0] w_n178_3;
	wire [2:0] w_n181_0;
	wire [1:0] w_n185_0;
	wire [2:0] w_n197_0;
	wire [2:0] w_n198_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n209_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [2:0] w_n219_0;
	wire [2:0] w_n222_0;
	wire [2:0] w_n233_0;
	wire [1:0] w_n233_1;
	wire [1:0] w_n234_0;
	wire [1:0] w_n235_0;
	wire [2:0] w_n239_0;
	wire [1:0] w_n239_1;
	wire [1:0] w_n240_0;
	wire [1:0] w_n241_0;
	wire [1:0] w_n242_0;
	wire [1:0] w_n245_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n258_0;
	wire [1:0] w_n260_0;
	wire [1:0] w_n262_0;
	wire [2:0] w_n267_0;
	wire [2:0] w_n285_0;
	wire [2:0] w_n303_0;
	wire [1:0] w_n303_1;
	wire [2:0] w_n306_0;
	wire [1:0] w_n306_1;
	wire [2:0] w_n311_0;
	wire [2:0] w_n311_1;
	wire [2:0] w_n319_0;
	wire [2:0] w_n319_1;
	wire [1:0] w_n320_0;
	wire [1:0] w_n321_0;
	wire [2:0] w_n327_0;
	wire [2:0] w_n327_1;
	wire [1:0] w_n328_0;
	wire [1:0] w_n329_0;
	wire [2:0] w_n335_0;
	wire [1:0] w_n335_1;
	wire [2:0] w_n336_0;
	wire [1:0] w_n339_0;
	wire [1:0] w_n343_0;
	wire [1:0] w_n346_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n352_0;
	wire [1:0] w_n355_0;
	wire [1:0] w_n361_0;
	wire [2:0] w_n377_0;
	wire [1:0] w_n391_0;
	wire [1:0] w_n393_0;
	wire [2:0] w_n404_0;
	wire [2:0] w_n420_0;
	wire w_dff_A_CGqpf3Ic4_1;
	wire w_dff_A_GrE8512v4_0;
	wire w_dff_B_Kxz2Dri24_2;
	wire w_dff_B_MUHJqlsa3_1;
	wire w_dff_B_D5KQVx4N8_1;
	wire w_dff_B_IMJTrLm56_1;
	wire w_dff_B_kltv1uDD9_1;
	wire w_dff_B_SWsBNjgP5_1;
	wire w_dff_B_SwAJvB7p8_1;
	wire w_dff_A_cdbfX95G2_1;
	wire w_dff_B_TPcV03838_1;
	wire w_dff_B_8q5RoEtf6_1;
	wire w_dff_B_5ygL2A6b4_1;
	wire w_dff_B_atjGC3YD0_1;
	wire w_dff_B_mOxQql009_1;
	wire w_dff_B_HNfNVR8z4_1;
	wire w_dff_B_sYsY2Xrd2_1;
	wire w_dff_B_JNhqm3lS9_1;
	wire w_dff_B_Tc3tWnSk6_0;
	wire w_dff_B_9AOImXTe6_0;
	wire w_dff_B_18Whazdq0_0;
	wire w_dff_B_mmVXoTq22_0;
	wire w_dff_B_9clIZ1G66_0;
	wire w_dff_B_i4hGdTD60_0;
	wire w_dff_B_x2sN5suX5_0;
	wire w_dff_B_mSd8cxZv9_0;
	wire w_dff_B_JkHntt2U0_0;
	wire w_dff_B_nzh4t6dO4_0;
	wire w_dff_B_KDBSoOv51_0;
	wire w_dff_A_kcSaOgBj7_0;
	wire w_dff_A_eOmbkkKK7_0;
	wire w_dff_A_ZJAKB7245_0;
	wire w_dff_A_l2oQh35B4_0;
	wire w_dff_B_c76GNu681_1;
	wire w_dff_B_VXEXTzTa3_1;
	wire w_dff_B_twHoBtLm8_1;
	wire w_dff_B_G23ZZq9F9_1;
	wire w_dff_B_mPC2hAMR7_1;
	wire w_dff_B_swztmzOe3_1;
	wire w_dff_B_iVi9uWFn7_0;
	wire w_dff_B_vd8DefqJ3_1;
	wire w_dff_B_FEjPi52X4_1;
	wire w_dff_B_kw8OM5yr9_1;
	wire w_dff_B_mdY2YZjG4_1;
	wire w_dff_B_4sjJETFE3_1;
	wire w_dff_B_FSdXD1d11_1;
	wire w_dff_B_abiyQRox7_0;
	wire w_dff_B_nUltx7Tg2_0;
	wire w_dff_B_sMTwHmq87_0;
	wire w_dff_B_BM4PMVxL2_0;
	wire w_dff_B_XYVWrlwg0_0;
	wire w_dff_B_peq3b0pW1_0;
	wire w_dff_B_TciQSPIr2_0;
	wire w_dff_A_RTB5cNrH8_1;
	wire w_dff_A_lT5BDjlx9_1;
	wire w_dff_A_7L9LTNAp1_1;
	wire w_dff_A_JhTgU0BS8_1;
	wire w_dff_A_ag8uLg3T9_1;
	wire w_dff_A_AkCmnQQX5_1;
	wire w_dff_A_TQi4cZKh2_0;
	wire w_dff_A_dg5UlAL93_0;
	wire w_dff_A_6qMOCYBK6_0;
	wire w_dff_A_0kLhHTXP1_0;
	wire w_dff_A_cbz4fwcC7_1;
	wire w_dff_A_YtPcYc5j3_1;
	wire w_dff_A_3EFehQgQ5_1;
	wire w_dff_A_QPAVvka71_1;
	wire w_dff_A_fHSpneZv5_1;
	wire w_dff_A_l1YZ2Gd11_1;
	wire w_dff_A_GZUfWPL59_1;
	wire w_dff_A_8YjeJZ702_1;
	wire w_dff_B_vfrcgtj62_1;
	wire w_dff_B_hpvNr7mY4_1;
	wire w_dff_B_Qc5Ep4Et7_1;
	wire w_dff_B_mSYXw8eD5_1;
	wire w_dff_B_KYyTr8kZ9_1;
	wire w_dff_B_9AB076ns0_0;
	wire w_dff_B_4IHM62Q08_0;
	wire w_dff_B_eRAyobKB9_0;
	wire w_dff_A_wWjTsjEO8_1;
	wire w_dff_B_w8J3QZD11_0;
	wire w_dff_B_6pBXQl0J0_0;
	wire w_dff_B_i5rM6Lyh2_0;
	wire w_dff_B_8bO6AFix8_1;
	wire w_dff_B_Mhj4yigo2_1;
	wire w_dff_B_5vQ5oGUA7_1;
	wire w_dff_B_GPFA6cjJ3_1;
	wire w_dff_B_qcuLo3QQ8_1;
	wire w_dff_B_7UHTb3y94_1;
	wire w_dff_B_z8ELfjDw5_1;
	wire w_dff_B_OpAWbcsq9_1;
	wire w_dff_B_Fg1Gbfcy3_1;
	wire w_dff_B_cbzNglHz5_1;
	wire w_dff_B_tLVV8sgM8_0;
	wire w_dff_B_ty9Yyy5w2_0;
	wire w_dff_B_AOlezAnq9_0;
	wire w_dff_B_D1nOBTit1_0;
	wire w_dff_B_YtZGeX4D6_0;
	wire w_dff_A_DzFSMGnM2_1;
	wire w_dff_A_s39czw265_1;
	wire w_dff_A_7O3U6y6e2_1;
	wire w_dff_A_QFejvGR19_1;
	wire w_dff_A_R43HBhu72_1;
	wire w_dff_B_cAjIsP5b6_1;
	wire w_dff_B_Ger2NZoh9_1;
	wire w_dff_B_fGvbyBJA5_1;
	wire w_dff_B_FX7SA9iW4_1;
	wire w_dff_B_LWzEiq9O1_0;
	wire w_dff_B_oFKigCyb2_0;
	wire w_dff_B_0iPckTON6_0;
	wire w_dff_B_5tk9Ng485_0;
	wire w_dff_B_4bUShkSf5_0;
	wire w_dff_B_QeLuuleW6_0;
	wire w_dff_B_ZfyCljN99_0;
	wire w_dff_B_jshBZBSI7_0;
	wire w_dff_B_cxlGlZI51_0;
	wire w_dff_B_qoyXegVq0_1;
	wire w_dff_B_IVrEZG6f2_1;
	wire w_dff_B_B3ass3li8_1;
	wire w_dff_B_pHz2bQjf1_1;
	wire w_dff_B_28Pg7Chg7_1;
	wire w_dff_B_oZ2mumHy2_1;
	wire w_dff_B_gLxFFouQ5_0;
	wire w_dff_B_KUqZWgip8_0;
	wire w_dff_B_FssnNeB03_0;
	wire w_dff_B_F7CSIpNA6_0;
	wire w_dff_B_NElr3muP5_0;
	wire w_dff_A_d7Xsperi1_1;
	wire w_dff_A_hjd6GLBh9_1;
	wire w_dff_A_Bf1tSGQD0_1;
	wire w_dff_A_vSxnLJ9U6_1;
	wire w_dff_B_9qzIs8wg5_1;
	wire w_dff_B_3a3WQmmx7_1;
	wire w_dff_B_q0XmMZTp5_1;
	wire w_dff_B_f4uRBHLF5_1;
	wire w_dff_B_ulRN76xC9_1;
	wire w_dff_B_nduxFZnu9_1;
	wire w_dff_B_t3ezegcD5_1;
	wire w_dff_B_UNokS3si3_1;
	wire w_dff_B_CBRBtQeq6_1;
	wire w_dff_B_WlG0mSKq4_1;
	wire w_dff_B_q2WYnYNi0_1;
	wire w_dff_B_FGgtUkCF1_1;
	wire w_dff_B_Dsin8gAB5_1;
	wire w_dff_B_0kJwRmP97_1;
	wire w_dff_B_iGT7ybQT9_1;
	wire w_dff_B_OcC37nY42_1;
	wire w_dff_B_dCPzLgYM7_1;
	wire w_dff_B_Aji7Bi1B0_1;
	wire w_dff_B_iOYwoYdk4_1;
	wire w_dff_B_dRqKBnj94_1;
	wire w_dff_B_o1wsCmzP6_1;
	wire w_dff_B_TDFpNZwg1_1;
	wire w_dff_A_dCMo2yu14_0;
	wire w_dff_A_HNKnGvbD6_0;
	wire w_dff_A_w1A9S7e51_0;
	wire w_dff_A_LwAixRhC6_0;
	wire w_dff_A_EuFvweOY7_0;
	wire w_dff_A_K3St2tcO9_0;
	wire w_dff_A_qIS9NgnR5_1;
	wire w_dff_A_CDGiNcbs7_1;
	wire w_dff_A_0VuttSU13_1;
	wire w_dff_A_rCUEQCJY8_1;
	wire w_dff_A_Y0wwgnqY3_1;
	wire w_dff_A_ZUppNKUk6_1;
	wire w_dff_B_9LrSJ0Kr3_0;
	wire w_dff_B_FuP7dzmg7_0;
	wire w_dff_B_Mdi0xSTC6_0;
	wire w_dff_B_FLIDAsOS3_0;
	wire w_dff_B_mvBzfZ2u9_0;
	wire w_dff_B_Nfcr0bzR3_0;
	wire w_dff_B_kSGpyvbW1_0;
	wire w_dff_B_y7IukNiW4_0;
	wire w_dff_B_xJNQDe2B7_0;
	wire w_dff_B_5e3LN8Mb1_0;
	wire w_dff_B_Q9e22nuI2_0;
	wire w_dff_B_W8HFDH5P9_1;
	wire w_dff_B_1JMh91Xp6_1;
	wire w_dff_B_jbJW216R2_1;
	wire w_dff_B_aeJyEo2r6_1;
	wire w_dff_A_982UkWgj0_0;
	wire w_dff_A_0RAZQmfo6_0;
	wire w_dff_A_VcS46n8X2_0;
	wire w_dff_A_7MmasVGu5_0;
	wire w_dff_A_CGl3dEfJ4_0;
	wire w_dff_A_LbkBKiXU0_0;
	wire w_dff_A_SaVK1kLN8_0;
	wire w_dff_A_rNMfhchC8_0;
	wire w_dff_A_S7Avvjfk1_0;
	wire w_dff_A_dy2TlCbN1_0;
	wire w_dff_A_c1NVpzwA2_0;
	wire w_dff_A_JfoasXjw1_0;
	wire w_dff_A_loYMBPnY5_0;
	wire w_dff_A_OQxJnndM3_0;
	wire w_dff_A_FMMyHLc56_0;
	wire w_dff_A_hLNHqSZs7_0;
	wire w_dff_A_Z5EfJoiX1_0;
	wire w_dff_A_SEYXpYpz4_0;
	wire w_dff_B_Pgydenyu2_1;
	wire w_dff_B_kigoaMPV8_1;
	wire w_dff_B_ua5mdZHW7_1;
	wire w_dff_B_tIB9YUQI7_1;
	wire w_dff_B_Gryezse61_1;
	wire w_dff_B_wHdF1m8M7_1;
	wire w_dff_B_4d6awUTU5_1;
	wire w_dff_A_NWvFy5Hw2_0;
	wire w_dff_A_Sdlj9REF0_0;
	wire w_dff_A_RcBFuB6l7_0;
	wire w_dff_A_lFqBu8ff3_1;
	wire w_dff_A_CIR6gLEO2_1;
	wire w_dff_A_yyLGguNy6_1;
	wire w_dff_A_nKSADduP4_1;
	wire w_dff_A_jOiGhT7j7_1;
	wire w_dff_A_dN2iwtJG6_0;
	wire w_dff_A_tuWIrX232_0;
	wire w_dff_A_3nDModQ05_0;
	wire w_dff_A_6uVQRxkF7_0;
	wire w_dff_A_xCGh9Dik9_0;
	wire w_dff_A_bDGdhnR76_0;
	wire w_dff_B_LdfayXuk2_1;
	wire w_dff_B_0zEf7tRx3_1;
	wire w_dff_B_idbxuYqm5_1;
	wire w_dff_B_QB7OndPV7_1;
	wire w_dff_B_fZ38KBMZ0_1;
	wire w_dff_B_HFDlZuMX4_1;
	wire w_dff_B_1JMPf21u8_1;
	wire w_dff_B_r008HAdm7_1;
	wire w_dff_B_qMihiaua6_1;
	wire w_dff_B_WIoMev244_1;
	wire w_dff_B_a7I7qVPu9_0;
	wire w_dff_B_ADo2BB3P8_0;
	wire w_dff_B_hjgrIZ3j7_0;
	wire w_dff_B_qjgcuFW77_0;
	wire w_dff_B_yiPhGhBJ3_0;
	wire w_dff_B_0h0mUdec1_0;
	wire w_dff_B_zTmpkxaA7_0;
	wire w_dff_B_l3ntDq6M2_0;
	wire w_dff_B_WzdsCEQ61_1;
	wire w_dff_B_wOXiouiC2_1;
	wire w_dff_B_1LLCSq9R4_1;
	wire w_dff_B_rNEezTIS7_1;
	wire w_dff_B_ZwnIq4qE3_1;
	wire w_dff_B_TReuXL9t2_1;
	wire w_dff_B_VAcRZKeS7_1;
	wire w_dff_B_WIKRwLFC7_1;
	wire w_dff_B_Fv3rBYbU3_1;
	wire w_dff_B_tR9RhVxv1_1;
	wire w_dff_B_oWFtll3n6_1;
	wire w_dff_B_MQp7jTcs0_1;
	wire w_dff_B_kQCU9bhP1_1;
	wire w_dff_A_Lw2nkXRA7_1;
	wire w_dff_A_2psb8fgB0_1;
	wire w_dff_A_ZW9u7zkC4_1;
	wire w_dff_A_VsPrxV389_1;
	wire w_dff_A_ntaRptit4_1;
	wire w_dff_A_Ixj01O2b5_1;
	wire w_dff_A_1EgNIh4p0_1;
	wire w_dff_A_SHhAVmmh8_1;
	wire w_dff_A_T11TeQpQ0_1;
	wire w_dff_A_FEZopSkl9_1;
	wire w_dff_A_Vfj7nTLU6_1;
	wire w_dff_A_uGUfn8pZ9_1;
	wire w_dff_A_OZAPhxzk8_1;
	wire w_dff_A_xsg5iuCv3_1;
	wire w_dff_A_58KaghXt5_1;
	wire w_dff_A_QSLRiiCz1_1;
	wire w_dff_A_2iUk5Bju8_1;
	wire w_dff_A_Jc707j8k5_1;
	wire w_dff_A_sopswqjr8_1;
	wire w_dff_A_tSEJwimh4_1;
	wire w_dff_A_WWdNkkQo7_0;
	wire w_dff_A_6aj3ALzR6_0;
	wire w_dff_A_WKqgjHLf1_0;
	wire w_dff_A_mGkyNChX3_0;
	wire w_dff_A_wJ0ToPjs9_0;
	wire w_dff_A_RIOFRY1c3_1;
	wire w_dff_A_61SjS4mf6_1;
	wire w_dff_A_UJ4GzRM53_1;
	wire w_dff_A_VznsKQfu4_1;
	wire w_dff_A_565O5jmn6_1;
	wire w_dff_B_tQydU9YP5_0;
	wire w_dff_B_Dkm7EISG0_0;
	wire w_dff_B_KD5l42ko3_0;
	wire w_dff_B_f5EXtC6H9_0;
	wire w_dff_B_Zb0KeNRc4_0;
	wire w_dff_B_XlqSPRHB8_0;
	wire w_dff_B_ykhVGkkf7_0;
	wire w_dff_B_6wNC4TZh8_0;
	wire w_dff_A_oDjmOo787_1;
	wire w_dff_A_4YXFuWR95_1;
	wire w_dff_A_Rtb4ygeS1_1;
	wire w_dff_A_5dzD6IV28_1;
	wire w_dff_A_Sti2pNHY4_1;
	wire w_dff_A_0gJUaOWj9_1;
	wire w_dff_A_UpJRFN434_1;
	wire w_dff_A_LOMqImEe6_1;
	wire w_dff_A_c1UHsm5x5_1;
	wire w_dff_A_J9C4nb5O7_1;
	wire w_dff_B_yanJwCB44_0;
	wire w_dff_B_c6refnxp3_0;
	wire w_dff_B_LUQVtbp02_0;
	wire w_dff_B_cI2qUmAb1_0;
	wire w_dff_B_aI0lAFX63_0;
	wire w_dff_B_OZFlQu3P9_1;
	wire w_dff_A_sF7pYkdu3_1;
	wire w_dff_A_36UdQolH2_1;
	wire w_dff_A_ZSdgoZUi4_1;
	wire w_dff_A_8WD9Ab1h0_1;
	wire w_dff_A_cXx4m2f19_1;
	wire w_dff_A_R3hqFTFh7_1;
	wire w_dff_A_07ktnM4N1_2;
	wire w_dff_A_p7sELI7H8_2;
	wire w_dff_A_sKT9uFrm1_2;
	wire w_dff_A_LYRp8ABC4_2;
	wire w_dff_A_MdwO1Gv75_2;
	wire w_dff_A_OYECsV1Y5_2;
	wire w_dff_A_upcNwBLK1_2;
	wire w_dff_B_rW1EU6Te4_1;
	wire w_dff_B_EyTziCDF9_1;
	wire w_dff_B_OBzCZk2W9_1;
	wire w_dff_B_wEdu6AHF8_1;
	wire w_dff_B_MssoguAC5_1;
	wire w_dff_B_72sKcRBa7_1;
	wire w_dff_B_BqekfUUL7_1;
	wire w_dff_B_woM3vRP19_1;
	wire w_dff_B_5EfUWnzb2_1;
	wire w_dff_B_E5KRjqAt4_0;
	wire w_dff_B_PpYIByju5_0;
	wire w_dff_B_DjiXcTp32_0;
	wire w_dff_B_qrNMyGa71_0;
	wire w_dff_B_bsbK8xZW9_0;
	wire w_dff_B_Zbk6Cu6J0_0;
	wire w_dff_B_cG3Xjw698_0;
	wire w_dff_B_mOUJgLFa0_1;
	wire w_dff_B_bNUevt1G2_1;
	wire w_dff_B_dXgHK3Yp3_1;
	wire w_dff_B_cZMYYE268_1;
	wire w_dff_B_vHnDE2rC4_1;
	wire w_dff_B_QkKGhZt22_1;
	wire w_dff_B_rk1a4uK05_1;
	wire w_dff_B_h1z0VhRv5_1;
	wire w_dff_B_7R8VIzpJ5_1;
	wire w_dff_B_IfJ9V8Iv0_1;
	wire w_dff_B_03IvlBp05_1;
	wire w_dff_A_SPHf5gbO2_1;
	wire w_dff_A_mS5cLRA47_1;
	wire w_dff_A_mGtiqhbr3_1;
	wire w_dff_A_zbMvYBGP4_1;
	wire w_dff_A_hHCAGVJo6_1;
	wire w_dff_A_CTbhVQDo6_1;
	wire w_dff_A_9ObARDXq4_1;
	wire w_dff_A_zJIgK1Bg2_1;
	wire w_dff_A_zqrSmoA51_1;
	wire w_dff_A_DedMGlCN7_1;
	wire w_dff_A_y6plcCYG4_1;
	wire w_dff_A_MkH3xeQL1_1;
	wire w_dff_A_r0cTBsIR1_1;
	wire w_dff_A_IuZ5LARV5_1;
	wire w_dff_A_6HCHyGQQ9_1;
	wire w_dff_A_TSZsjlpV1_1;
	wire w_dff_A_DlXKxutM3_1;
	wire w_dff_A_fQNP7HS99_1;
	wire w_dff_A_bD5zvcQ85_0;
	wire w_dff_A_HYozMjNj5_0;
	wire w_dff_A_o90QN0yh6_0;
	wire w_dff_A_ePc1xQin2_0;
	wire w_dff_A_7UQSFdWA5_0;
	wire w_dff_A_YmakPBz43_0;
	wire w_dff_A_uSBCJs0L2_1;
	wire w_dff_A_CJVIKroK9_1;
	wire w_dff_A_jiVdyjUa6_1;
	wire w_dff_A_dfbKhmrs3_1;
	wire w_dff_A_B16m9Pz97_1;
	wire w_dff_A_xrAKoSCS0_1;
	wire w_dff_B_vZpFLVwD0_0;
	wire w_dff_B_DrDOqf6g9_0;
	wire w_dff_B_ZLQlakEG2_0;
	wire w_dff_B_C0eZyB142_0;
	wire w_dff_B_JjyBe0Tl7_0;
	wire w_dff_B_Rhue5dRa1_0;
	wire w_dff_B_i3zowgiz9_0;
	wire w_dff_B_AXPtbETS2_0;
	wire w_dff_A_0IQAcb3k1_1;
	wire w_dff_A_SmWtqAwe8_1;
	wire w_dff_A_s16vtcMS6_1;
	wire w_dff_A_uiFXOIqy7_1;
	wire w_dff_A_tVvGk56O2_1;
	wire w_dff_A_ehnFyZms5_1;
	wire w_dff_A_2H2vucLm3_1;
	wire w_dff_A_esZKSQfr0_1;
	wire w_dff_A_n2wj0pkY2_1;
	wire w_dff_A_fKX7qDbX4_1;
	wire w_dff_A_AXBQXbDI0_1;
	wire w_dff_A_MKvadVPG1_1;
	wire w_dff_A_SOubNi2I9_1;
	wire w_dff_A_QBszpqbZ2_1;
	wire w_dff_B_zVjBrFHL1_0;
	wire w_dff_B_og1wBcb82_0;
	wire w_dff_B_ydvYg7mL0_0;
	wire w_dff_B_bQDqAH6q8_0;
	wire w_dff_B_9JrxwEvH3_0;
	wire w_dff_A_J3nc7o1c4_1;
	wire w_dff_A_Qe7FKe0u8_1;
	wire w_dff_A_cOvZmYvq4_1;
	wire w_dff_A_ovxeSliI1_1;
	wire w_dff_A_Tm74dXJS5_1;
	wire w_dff_A_IqRzScHt9_2;
	wire w_dff_A_cUN7fqHM0_2;
	wire w_dff_A_9DkCoM124_2;
	wire w_dff_A_eCraVxkm0_2;
	wire w_dff_A_Vt9q6fv93_2;
	wire w_dff_A_yqRDbJJ93_2;
	wire w_dff_B_jhSL01uD2_3;
	wire w_dff_B_KJXC6WmS8_1;
	wire w_dff_B_dOaZpg373_1;
	wire w_dff_B_TlNcn5Pv4_1;
	wire w_dff_B_uJlR2KdT4_1;
	wire w_dff_B_aeYg415G4_1;
	wire w_dff_B_sMyLpKxq2_1;
	wire w_dff_B_3eVLZlkj4_1;
	wire w_dff_B_YSwBDnKS8_1;
	wire w_dff_B_Jmt0lTr00_1;
	wire w_dff_B_6FS7ywOQ1_1;
	wire w_dff_B_aKQvAoRF6_1;
	wire w_dff_B_74NRWyks0_1;
	wire w_dff_B_xuosGLmR3_1;
	wire w_dff_B_SZO2vpfW5_1;
	wire w_dff_B_vctFiGWx8_1;
	wire w_dff_B_oWJGObSn8_1;
	wire w_dff_B_fnNvb5kg5_1;
	wire w_dff_B_XXM4xDtG9_1;
	wire w_dff_B_NxF3yOF08_1;
	wire w_dff_B_eyRduMUH2_1;
	wire w_dff_B_CFs5Y1xx7_1;
	wire w_dff_B_yMHv5IkB9_0;
	wire w_dff_B_zXYD6iSI0_0;
	wire w_dff_B_DWlw1QNO9_0;
	wire w_dff_B_S3sYJPcS1_0;
	wire w_dff_A_Wf2H0hlY2_0;
	wire w_dff_A_ZjTjFceJ6_2;
	wire w_dff_A_IAiiqf3i6_0;
	wire w_dff_A_o97X8kgB7_0;
	wire w_dff_A_Kbnq7u2O1_0;
	wire w_dff_A_Z46QNUuo2_0;
	wire w_dff_A_zS1JG0L90_0;
	wire w_dff_A_trNkA0at5_2;
	wire w_dff_B_NFJP6KVg8_3;
	wire w_dff_B_zjjYFn9h6_3;
	wire w_dff_B_8A0IAFZs3_3;
	wire w_dff_B_TzjtyDDp6_3;
	wire w_dff_B_17y8TwHh1_3;
	wire w_dff_B_1nGfh1w22_3;
	wire w_dff_B_qusmwgnb2_3;
	wire w_dff_B_lh7zMWQ93_3;
	wire w_dff_B_wDGhJLLo9_3;
	wire w_dff_B_SWnVk3fM4_0;
	wire w_dff_B_faK5CgCR4_0;
	wire w_dff_B_OpAQCHQY5_0;
	wire w_dff_B_mVVOJtFA1_0;
	wire w_dff_B_mYze1cyB0_0;
	wire w_dff_B_HgvTrgrE4_1;
	wire w_dff_B_9LoH4KPU1_1;
	wire w_dff_B_aTDe0dh08_1;
	wire w_dff_B_CfTfS9m79_1;
	wire w_dff_B_odkAes6T3_1;
	wire w_dff_B_fFMHPjKW7_1;
	wire w_dff_B_iQF2qdDc8_1;
	wire w_dff_B_iAbdEwOF6_1;
	wire w_dff_B_174OM27a1_1;
	wire w_dff_B_vhh45I5e9_1;
	wire w_dff_B_TOWDjmT62_1;
	wire w_dff_B_qbt2vy6h2_1;
	wire w_dff_B_mlaOqiYt2_1;
	wire w_dff_B_AEHREUcU6_1;
	wire w_dff_B_KHqf8zhh8_1;
	wire w_dff_A_dXaXVj1q0_1;
	wire w_dff_A_ksjfY7GK7_1;
	wire w_dff_B_XdtsCMJR9_2;
	wire w_dff_B_SiCG6sbq2_2;
	wire w_dff_B_v0KGXehj0_2;
	wire w_dff_B_JyUnwTMj7_2;
	wire w_dff_B_8CLSBiVb8_2;
	wire w_dff_B_4SBoA1ic7_2;
	wire w_dff_B_tgNJEoev1_2;
	wire w_dff_A_1IBYGsO18_0;
	wire w_dff_A_D4woEsY74_0;
	wire w_dff_A_jB1P23PB0_0;
	wire w_dff_A_SiiAtopi7_0;
	wire w_dff_A_gWlp2XUR5_0;
	wire w_dff_A_CHDEXkLs0_0;
	wire w_dff_A_7wpFEAVr2_0;
	wire w_dff_A_6gRVB6vU5_2;
	wire w_dff_A_oD1PAPfr0_2;
	wire w_dff_A_nnfEkIhN5_2;
	wire w_dff_A_UkosGhHV9_2;
	wire w_dff_A_kLSexX1o4_2;
	wire w_dff_A_sL0toZFT4_2;
	wire w_dff_A_nqQkIykf5_2;
	wire w_dff_A_alRdQcG84_2;
	wire w_dff_A_Xvcckb5q5_2;
	wire w_dff_B_EEo6iHmn8_0;
	wire w_dff_B_QHzuWFgV4_0;
	wire w_dff_B_yWnPKxVu2_0;
	wire w_dff_B_8rvGSJTv5_0;
	wire w_dff_B_LXHGXDS25_1;
	wire w_dff_B_rjEnrd192_1;
	wire w_dff_B_VNrkrfuU0_1;
	wire w_dff_B_yzra5jcw6_0;
	wire w_dff_A_UBalm7Lv3_1;
	wire w_dff_A_pD37gmHI4_1;
	wire w_dff_A_RBhIt13U0_1;
	wire w_dff_A_sOLrYTH73_1;
	wire w_dff_A_zkfDkXYw9_1;
	wire w_dff_B_06ecEtg02_3;
	wire w_dff_B_oq7NxDPX3_3;
	wire w_dff_B_UEkLvT6m8_3;
	wire w_dff_B_yFgtCBhi9_3;
	wire w_dff_B_z5Smd1ad6_3;
	wire w_dff_B_rmc1moKw7_3;
	wire w_dff_B_aeLYM4i55_3;
	wire w_dff_A_suOJKDa05_1;
	wire w_dff_A_YZ83nlWG2_1;
	wire w_dff_A_IPvx8p3y3_1;
	wire w_dff_A_b2awXjOu8_1;
	wire w_dff_A_H8RsPoNV2_1;
	wire w_dff_A_wB7S1cRe7_1;
	wire w_dff_A_ULAE3HpL3_1;
	wire w_dff_A_DpahGmAm1_1;
	wire w_dff_A_d11fSYTr4_1;
	wire w_dff_A_ESlTA6IA9_1;
	wire w_dff_A_OPWn0AdZ8_1;
	wire w_dff_A_YSF8Dwbr8_1;
	wire w_dff_A_q5LsXBCT6_1;
	wire w_dff_A_Zl6fLIM01_1;
	wire w_dff_A_5I7d8ltg5_1;
	wire w_dff_A_uvNG0BQX1_1;
	wire w_dff_A_U1w57x487_1;
	wire w_dff_A_nEtWniCD5_2;
	wire w_dff_A_PZTH6ZlS0_2;
	wire w_dff_A_w7mMJzuS1_2;
	wire w_dff_A_myQyaN844_2;
	wire w_dff_A_oyiRnW668_2;
	wire w_dff_A_SYPybmbJ0_2;
	wire w_dff_A_OQsddf6b0_1;
	wire w_dff_A_EQ06nY0c5_1;
	wire w_dff_A_BONjA3LD0_1;
	wire w_dff_A_JeGlmZaJ4_1;
	wire w_dff_A_gblR4WM46_1;
	wire w_dff_B_GZeGIeJg7_0;
	wire w_dff_A_dCB7B7Mt5_0;
	wire w_dff_A_p8ekeHrl2_0;
	wire w_dff_A_jyotcOTw4_0;
	wire w_dff_A_XwizvcJe4_0;
	wire w_dff_A_KyQsSQ0E2_0;
	wire w_dff_A_r2rIaCPk6_0;
	wire w_dff_A_8RPEXi2V4_0;
	wire w_dff_A_nWYoHk6q9_0;
	wire w_dff_A_CblQHe8Z2_0;
	wire w_dff_A_AugJmRfe2_0;
	wire w_dff_A_nYxAQpCt9_0;
	wire w_dff_A_mph99VEh3_2;
	wire w_dff_A_E2JqAQvl6_2;
	wire w_dff_A_v8QyBFIZ8_2;
	wire w_dff_A_hB4lQznq7_2;
	wire w_dff_A_nWno1Wal2_1;
	wire w_dff_A_re5dLjmD7_1;
	wire w_dff_A_sgBEVCZO9_1;
	wire w_dff_A_fT2zX8mp0_1;
	wire w_dff_A_Cd0ItszR6_1;
	wire w_dff_A_LqsTnaKk6_1;
	wire w_dff_A_FObxGTHh5_1;
	wire w_dff_A_ktS4YwME7_1;
	wire w_dff_A_8u6x1zgP9_1;
	wire w_dff_A_Y14E0BAy5_1;
	wire w_dff_A_CP88kakA0_1;
	wire w_dff_A_3VLFMT3U3_1;
	wire w_dff_A_Nhp5KMZX9_2;
	wire w_dff_A_MFyv88hl6_2;
	wire w_dff_A_d5bGZOk15_2;
	wire w_dff_A_vtQCxj908_2;
	wire w_dff_A_87qMAd0C7_2;
	wire w_dff_A_8cuxrSrU0_2;
	wire w_dff_A_bXXcMXfy8_1;
	wire w_dff_A_0lAv7VJc6_1;
	wire w_dff_A_2XhZqoQH4_1;
	wire w_dff_A_2iJHIspx2_1;
	wire w_dff_A_2agpt3LK1_1;
	wire w_dff_A_vVTloqkZ2_1;
	wire w_dff_B_FqU1p9qq9_0;
	wire w_dff_B_0ilOWy2G4_2;
	wire w_dff_B_MRjS1Njp8_2;
	wire w_dff_B_gRcPpe5u6_2;
	wire w_dff_B_NSpcUwYz7_2;
	wire w_dff_A_oZmKzSsl3_1;
	wire w_dff_A_97LCpHz03_1;
	wire w_dff_A_crK0N7Vs8_1;
	wire w_dff_A_c1N16EQg6_1;
	wire w_dff_A_bWkaAc2M5_1;
	wire w_dff_A_tXEFaYxt1_0;
	wire w_dff_A_tS9FdZ5z7_0;
	wire w_dff_A_CwYXyIC57_0;
	wire w_dff_A_UzEpeajt9_0;
	wire w_dff_A_IHAUkHO70_0;
	wire w_dff_A_otoplOJD7_0;
	wire w_dff_A_GI8UFyGU1_2;
	wire w_dff_A_zDQ4ax1z6_2;
	wire w_dff_A_MX0Zr1Yw4_2;
	wire w_dff_A_Lb4784C42_2;
	wire w_dff_A_PotDqNv55_0;
	wire w_dff_A_vcxIwZ0Q9_0;
	wire w_dff_A_Uex1Sy8D9_0;
	wire w_dff_B_BFM5aiq04_1;
	wire w_dff_B_aPH4xSno0_1;
	wire w_dff_B_LHtW3sfA3_1;
	wire w_dff_B_1Wcb2P884_1;
	wire w_dff_B_eiKI6U6S8_1;
	wire w_dff_B_HC1jVCeB8_1;
	wire w_dff_A_5cxBnz5X5_1;
	wire w_dff_A_fLnI7T5g4_1;
	wire w_dff_A_VOjLmj5e3_1;
	wire w_dff_A_YOt3qKd65_1;
	wire w_dff_A_qjpVXUau6_1;
	wire w_dff_A_BVH0VYLg1_1;
	wire w_dff_A_gnhZkBHY0_1;
	wire w_dff_B_tExV6k4Y7_0;
	wire w_dff_A_zQVbo4Md0_0;
	wire w_dff_A_KthTLXre9_0;
	wire w_dff_A_AwLQZzfH2_0;
	wire w_dff_B_YcLKcsg87_2;
	wire w_dff_B_MT7eeJA04_2;
	wire w_dff_B_DgHKgcrT3_2;
	wire w_dff_B_9ieTWPER3_2;
	wire w_dff_A_YkoPwWJI0_1;
	wire w_dff_A_QhNNhfQG7_1;
	wire w_dff_A_zYDUrmcf6_1;
	wire w_dff_A_H8oosr1I6_1;
	wire w_dff_A_wbINvpvQ9_1;
	wire w_dff_A_ibJ16uri5_2;
	wire w_dff_A_USHhy8Zp4_2;
	wire w_dff_A_pUoGMm6J3_2;
	wire w_dff_A_y0tuKOT93_2;
	wire w_dff_A_EnOzxcB10_2;
	wire w_dff_A_SOYVUpiV3_2;
	wire w_dff_A_ofK71HAU6_0;
	wire w_dff_A_oNxFUwe10_0;
	wire w_dff_A_xyIK1zVJ4_0;
	wire w_dff_A_6ChR3N6F0_0;
	wire w_dff_B_PEHi7lLT7_1;
	wire w_dff_B_5pYlq4ee6_1;
	wire w_dff_B_OhZtvwu41_1;
	wire w_dff_B_BuP4IWfi8_1;
	wire w_dff_B_uT4SdLTS5_1;
	wire w_dff_B_6NKaHX122_1;
	wire w_dff_A_xSUtLzvB8_2;
	wire w_dff_A_PkRi1psv1_2;
	wire w_dff_A_QzUVvIL82_2;
	wire w_dff_A_a8LNnxp19_2;
	wire w_dff_A_4jYozLls1_2;
	wire w_dff_A_svH6yMxW8_2;
	wire w_dff_A_Rr19MyhV6_2;
	wire w_dff_A_8pmlUdXC8_2;
	wire w_dff_B_Fdm4RsM11_0;
	wire w_dff_B_s1Db8RCQ1_0;
	wire w_dff_B_EdJFt1En8_0;
	wire w_dff_B_jIabbdRv7_0;
	wire w_dff_B_xfwW9Hcw6_0;
	wire w_dff_A_fvIu41ZS9_0;
	wire w_dff_A_My0mWd8l0_0;
	wire w_dff_A_cac9qL9k1_0;
	wire w_dff_A_xpiSFEr42_0;
	wire w_dff_A_tVlgc52J8_2;
	wire w_dff_A_SoFnZV9s5_2;
	wire w_dff_A_lFsG8WrJ4_2;
	wire w_dff_A_5PsbKJ721_2;
	wire w_dff_A_TyLSCsX71_0;
	wire w_dff_A_jHSDHRod4_0;
	wire w_dff_A_29S4EfEs0_0;
	wire w_dff_A_tDyp7s3m2_0;
	wire w_dff_A_7RxM1HFo4_0;
	wire w_dff_A_Q5tBt3Dt9_1;
	wire w_dff_A_E1zMHKly0_1;
	wire w_dff_A_giy5uNC20_1;
	wire w_dff_A_VzVE7bFf2_1;
	wire w_dff_A_i1d2TrVF8_1;
	wire w_dff_A_lUNGMeER4_1;
	wire w_dff_A_2tKN5lYi4_1;
	wire w_dff_A_2rwWqu043_1;
	wire w_dff_A_hFupe5IP8_1;
	wire w_dff_A_HocxKQJ23_1;
	wire w_dff_A_01X2N3y46_2;
	wire w_dff_A_UGQgXXv72_2;
	wire w_dff_A_eflLSDKj8_2;
	wire w_dff_A_VddeiRVt5_2;
	wire w_dff_A_9voGgNWk1_2;
	wire w_dff_A_rKopKHok9_2;
	wire w_dff_B_viTRVlxQ2_0;
	wire w_dff_A_jBnBKk4m9_0;
	wire w_dff_A_J4srjupc3_0;
	wire w_dff_A_me8cEVlX2_0;
	wire w_dff_A_m2fWDuOw9_0;
	wire w_dff_A_XvYe7sEs4_0;
	wire w_dff_A_hSenj8Fx6_2;
	wire w_dff_A_pEiVFWVm5_2;
	wire w_dff_A_cWUMsuP71_2;
	wire w_dff_A_XTSl5f3d1_2;
	wire w_dff_A_dio62ymb4_2;
	wire w_dff_B_ML60B5756_3;
	wire w_dff_B_Bgn1qL6f9_0;
	wire w_dff_B_YSglphc89_0;
	wire w_dff_B_0gGQ4aty2_0;
	wire w_dff_B_DowX2YEs5_0;
	wire w_dff_B_dFK2gmNP0_0;
	wire w_dff_B_UyXzk69G3_0;
	wire w_dff_B_sKQwZKGO0_0;
	wire w_dff_A_3S1ZAduI2_1;
	wire w_dff_A_6NDJ6yQb2_1;
	wire w_dff_A_eTmUPtl63_1;
	wire w_dff_A_aJpXrbLV9_1;
	wire w_dff_A_jJ3Agiua5_1;
	wire w_dff_A_0cWndKis9_0;
	wire w_dff_A_819gHp0h9_0;
	wire w_dff_A_Oac5nl3V1_0;
	wire w_dff_A_dfgJzSTR9_0;
	wire w_dff_A_oZNfvIV19_0;
	wire w_dff_A_pv6Llxho5_0;
	wire w_dff_A_NZNGj85j5_0;
	wire w_dff_A_pXiBHGgW9_0;
	wire w_dff_B_Zz8qS1RX9_3;
	wire w_dff_B_zYXFjQ8f0_3;
	wire w_dff_B_FCpXZ9jE2_3;
	wire w_dff_B_yayIqxlm6_3;
	wire w_dff_B_6N5lYVNw8_3;
	wire w_dff_B_AqJWYsQB9_3;
	wire w_dff_B_PKDSliMz0_3;
	wire w_dff_B_aSMCM9EO5_0;
	wire w_dff_B_4QqzGzgF3_0;
	wire w_dff_B_O7heLr722_0;
	wire w_dff_B_rR21cPeg6_0;
	wire w_dff_B_MSQsjCHr1_0;
	wire w_dff_A_dOndz9hd4_1;
	wire w_dff_B_cxQVaFZO1_2;
	wire w_dff_B_Ts7w3xfM1_2;
	wire w_dff_B_PZTWlNOE1_2;
	wire w_dff_B_yWvWJbNP7_2;
	wire w_dff_B_S6JGZ4BK1_0;
	wire w_dff_B_3Mit8GXY2_0;
	wire w_dff_B_uBWyZ4wu8_1;
	wire w_dff_A_EuLMJAVz8_1;
	wire w_dff_A_XDrhQoL33_0;
	wire w_dff_A_svFjUYC56_2;
	wire w_dff_A_8o2GDxRU3_2;
	wire w_dff_A_HBKRtCN28_1;
	wire w_dff_A_CGNMA64Z8_1;
	wire w_dff_A_sojqwtga4_1;
	wire w_dff_A_kIJH5AZc0_1;
	wire w_dff_A_5QQC5bE49_1;
	wire w_dff_A_GzPcAlQd1_2;
	wire w_dff_A_tZhBeJBZ3_1;
	wire w_dff_A_rMq5VKvg8_0;
	wire w_dff_A_75Zmf9AN2_0;
	wire w_dff_A_2b6CFqz22_2;
	wire w_dff_A_HumMNYpW3_0;
	wire w_dff_A_8YW7iErV4_0;
	wire w_dff_A_oWqVhi8U0_0;
	wire w_dff_A_k2hAoUcH6_0;
	wire w_dff_A_U5kbN1Si1_0;
	wire w_dff_A_F5JMnWxN1_0;
	wire w_dff_A_OYHwywK25_0;
	wire w_dff_A_ra75qUdI7_0;
	wire w_dff_A_kGD97uD18_0;
	wire w_dff_A_s4RucgmH5_1;
	wire w_dff_A_F6szztgT6_1;
	wire w_dff_A_R3mMVGf93_1;
	wire w_dff_B_6a7pafLu0_2;
	wire w_dff_B_Z6YaJEQ33_2;
	wire w_dff_B_SNIlPIe11_2;
	wire w_dff_B_nqtVZAax0_2;
	wire w_dff_A_nKhPqxsF5_0;
	wire w_dff_A_TfErT3cr0_0;
	wire w_dff_A_7P5OOGI81_0;
	wire w_dff_A_wN3TuHHf4_0;
	wire w_dff_A_eD2zl0ft8_0;
	wire w_dff_A_3StBpSnb5_0;
	wire w_dff_A_Ms4I4KGx6_2;
	wire w_dff_A_j3KPQP6N1_2;
	wire w_dff_A_QXsUzNsy5_2;
	wire w_dff_A_zz3gx5pR3_2;
	wire w_dff_A_aD3vSyb00_2;
	wire w_dff_A_YjhNPzNL6_2;
	wire w_dff_A_DwycHNr98_2;
	wire w_dff_A_JpqlyuDb6_0;
	wire w_dff_A_LTmUMlhz6_0;
	wire w_dff_A_xHTspfHT1_0;
	wire w_dff_B_MqzXXQpS0_0;
	wire w_dff_A_5mOXuFtE3_1;
	wire w_dff_A_uX1ST8167_1;
	wire w_dff_A_Cw9lnBBc6_1;
	wire w_dff_A_z6M065IR9_1;
	wire w_dff_A_IxRrFqPx2_1;
	wire w_dff_A_uUTggaeS6_1;
	wire w_dff_A_7uPyF1rD4_1;
	wire w_dff_A_Okid8rW94_1;
	wire w_dff_A_tuOdJaz41_2;
	wire w_dff_A_iCl7TOn50_1;
	wire w_dff_A_hw9j201Q8_1;
	wire w_dff_A_YW6fEiix2_0;
	wire w_dff_A_z1Q9CbA68_1;
	wire w_dff_A_nmfxa6Js2_1;
	wire w_dff_B_mL6ahJM19_3;
	wire w_dff_B_i5JhTpjB3_3;
	wire w_dff_A_5NJTiXpF1_1;
	wire w_dff_A_nKiX7A6H8_1;
	wire w_dff_A_sBEqGzWZ3_1;
	wire w_dff_A_AWASG99i6_1;
	wire w_dff_A_Q5vtmiXM1_1;
	wire w_dff_A_pkWdKiuy2_1;
	wire w_dff_A_qgJr1mYT1_2;
	wire w_dff_A_UlNQ7CI57_2;
	wire w_dff_A_WoO4NXHP1_2;
	wire w_dff_A_ZSdoUlp44_2;
	wire w_dff_A_1aAZXfux4_2;
	wire w_dff_A_iscgakJ79_2;
	wire w_dff_A_4MhYOLGE7_2;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(G388gat),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(G389gat),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(G391gat),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_n92_0[1]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_G17gat_2[2]),.dout(G418gat),.clk(gclk));
	jnot g009(.din(w_G17gat_2[1]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G13gat_0[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G1gat_1[0]),.dout(n97),.clk(gclk));
	jnot g012(.din(w_G26gat_0[1]),.dout(n98),.clk(gclk));
	jcb g013(.dina(n98),.dinb(w_n97_0[1]),.dout(n99));
	jcb g014(.dina(w_n99_0[1]),.dinb(n96),.dout(n100));
	jcb g015(.dina(n100),.dinb(w_n95_0[2]),.dout(n101));
	jcb g016(.dina(w_n101_0[1]),.dinb(w_G390gat_0[1]),.dout(G419gat));
	jnot g017(.din(w_G80gat_0[1]),.dout(n103),.clk(gclk));
	jand g018(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n104),.clk(gclk));
	jnot g019(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jcb g020(.dina(n105),.dinb(w_n103_0[1]),.dout(G420gat));
	jnot g021(.din(w_G36gat_0[0]),.dout(n107),.clk(gclk));
	jnot g022(.din(w_G59gat_1[0]),.dout(n108),.clk(gclk));
	jcb g023(.dina(w_n108_0[1]),.dinb(n107),.dout(n109));
	jcb g024(.dina(w_n109_0[1]),.dinb(w_n103_0[0]),.dout(G421gat));
	jnot g025(.din(w_G42gat_1[2]),.dout(n111),.clk(gclk));
	jcb g026(.dina(w_n109_0[0]),.dinb(w_n111_0[1]),.dout(G422gat));
	jcb g027(.dina(G88gat),.dinb(G87gat),.dout(n113));
	jand g028(.dina(w_n113_0[1]),.dinb(G90gat),.dout(G423gat),.clk(gclk));
	jnot g029(.din(w_G390gat_0[0]),.dout(n115),.clk(gclk));
	jcb g030(.dina(w_n101_0[0]),.dinb(n115),.dout(G446gat));
	jand g031(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g033(.dina(w_n93_0[0]),.dinb(w_G55gat_0[2]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_n119_0[2]),.dinb(w_G29gat_0[0]),.dout(n120),.clk(gclk));
	jand g035(.dina(n120),.dinb(w_G68gat_0[1]),.dout(G448gat),.clk(gclk));
	jand g036(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n122),.clk(gclk));
	jand g037(.dina(w_n119_0[1]),.dinb(w_dff_B_IMJTrLm56_1),.dout(n123),.clk(gclk));
	jand g038(.dina(n123),.dinb(w_n122_0[1]),.dout(G449gat),.clk(gclk));
	jand g039(.dina(w_n113_0[0]),.dinb(G89gat),.dout(G450gat),.clk(gclk));
	jxor g040(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n126),.clk(gclk));
	jxor g041(.dina(n126),.dinb(w_dff_B_SWsBNjgP5_1),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n128),.clk(gclk));
	jxor g043(.dina(n128),.dinb(w_G130gat_0[1]),.dout(n129),.clk(gclk));
	jxor g044(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G126gat_0[2]),.dinb(w_G121gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(n131),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n129),.dout(n133),.clk(gclk));
	jxor g048(.dina(n133),.dinb(w_dff_B_kltv1uDD9_1),.dout(G767gat),.clk(gclk));
	jxor g049(.dina(w_G189gat_2[1]),.dinb(w_G183gat_1[2]),.dout(n135),.clk(gclk));
	jxor g050(.dina(n135),.dinb(w_dff_B_TPcV03838_1),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_G159gat_1[2]),.dinb(w_G130gat_0[0]),.dout(n137),.clk(gclk));
	jxor g052(.dina(n137),.dinb(w_G165gat_1[2]),.dout(n138),.clk(gclk));
	jxor g053(.dina(w_G177gat_1[2]),.dinb(w_G171gat_1[2]),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G201gat_1[1]),.dinb(w_G195gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g057(.dina(n142),.dinb(w_dff_B_SwAJvB7p8_1),.dout(G768gat),.clk(gclk));
	jnot g058(.din(w_G268gat_0[1]),.dout(n144),.clk(gclk));
	jand g059(.dina(w_G447gat_1),.dinb(w_G80gat_0[0]),.dout(n145),.clk(gclk));
	jand g060(.dina(n145),.dinb(w_n86_0[0]),.dout(n146),.clk(gclk));
	jand g061(.dina(w_n146_0[1]),.dinb(w_G55gat_0[1]),.dout(n147),.clk(gclk));
	jand g062(.dina(n147),.dinb(w_n144_0[1]),.dout(n148),.clk(gclk));
	jand g063(.dina(w_n111_0[0]),.dinb(w_n95_0[1]),.dout(n149),.clk(gclk));
	jnot g064(.din(w_n149_0[1]),.dout(n150),.clk(gclk));
	jand g065(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(w_G42gat_1[1]),.dinb(w_G17gat_2[0]),.dout(n152),.clk(gclk));
	jnot g067(.din(w_n152_0[1]),.dout(n153),.clk(gclk));
	jand g068(.dina(n153),.dinb(w_n151_0[1]),.dout(n154),.clk(gclk));
	jand g069(.dina(n154),.dinb(w_G447gat_0[2]),.dout(n155),.clk(gclk));
	jand g070(.dina(n155),.dinb(w_dff_B_uBWyZ4wu8_1),.dout(n156),.clk(gclk));
	jnot g071(.din(w_n92_0[0]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n104_0[0]),.dinb(w_G42gat_1[0]),.dout(n158),.clk(gclk));
	jand g073(.dina(w_G51gat_1[0]),.dinb(w_G17gat_1[2]),.dout(n159),.clk(gclk));
	jnot g074(.din(n159),.dout(n160),.clk(gclk));
	jcb g075(.dina(n160),.dinb(n158),.dout(n161));
	jcb g076(.dina(n161),.dinb(n157),.dout(n162));
	jnot g077(.din(w_n162_0[1]),.dout(n163),.clk(gclk));
	jcb g078(.dina(w_dff_B_3Mit8GXY2_0),.dinb(n156),.dout(n164));
	jand g079(.dina(w_n164_3[1]),.dinb(w_G126gat_0[1]),.dout(n165),.clk(gclk));
	jnot g080(.din(w_G156gat_0[0]),.dout(n166),.clk(gclk));
	jcb g081(.dina(n166),.dinb(w_n108_0[0]),.dout(n167));
	jand g082(.dina(w_n167_0[1]),.dinb(w_G447gat_0[1]),.dout(n168),.clk(gclk));
	jand g083(.dina(w_n168_0[1]),.dinb(w_G17gat_1[1]),.dout(n169),.clk(gclk));
	jcb g084(.dina(n169),.dinb(w_n97_0[0]),.dout(n170));
	jand g085(.dina(w_n170_1[1]),.dinb(w_G153gat_0[2]),.dout(n171),.clk(gclk));
	jcb g086(.dina(w_dff_B_S3sYJPcS1_0),.dinb(n165),.dout(n172));
	jcb g087(.dina(n172),.dinb(w_n148_1[2]),.dout(n173));
	jand g088(.dina(w_n173_0[1]),.dinb(w_G246gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_n122_0[0]),.dinb(w_G42gat_0[2]),.dout(n175),.clk(gclk));
	jand g090(.dina(G73gat),.dinb(G72gat),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_MqzXXQpS0_0),.dinb(n175),.dout(n177),.clk(gclk));
	jand g092(.dina(n177),.dinb(w_n119_0[0]),.dout(n178),.clk(gclk));
	jand g093(.dina(w_n178_3[1]),.dinb(w_G201gat_1[0]),.dout(n179),.clk(gclk));
	jcb g094(.dina(w_dff_B_KDBSoOv51_0),.dinb(n174),.dout(n180));
	jnot g095(.din(w_G201gat_0[2]),.dout(n181),.clk(gclk));
	jnot g096(.din(w_n148_1[1]),.dout(n182),.clk(gclk));
	jnot g097(.din(w_G126gat_0[0]),.dout(n183),.clk(gclk));
	jnot g098(.din(w_G51gat_0[2]),.dout(n184),.clk(gclk));
	jcb g099(.dina(w_n99_0[0]),.dinb(n184),.dout(n185));
	jcb g100(.dina(w_n152_0[0]),.dinb(w_n167_0[0]),.dout(n186));
	jcb g101(.dina(n186),.dinb(w_n185_0[1]),.dout(n187));
	jcb g102(.dina(w_dff_B_yzra5jcw6_0),.dinb(w_n149_0[0]),.dout(n188));
	jand g103(.dina(w_n162_0[0]),.dinb(n188),.dout(n189),.clk(gclk));
	jcb g104(.dina(n189),.dinb(w_dff_B_VNrkrfuU0_1),.dout(n190));
	jnot g105(.din(w_G153gat_0[1]),.dout(n191),.clk(gclk));
	jcb g106(.dina(w_n151_0[0]),.dinb(w_n185_0[0]),.dout(n192));
	jcb g107(.dina(n192),.dinb(w_n95_0[0]),.dout(n193));
	jand g108(.dina(n193),.dinb(w_G1gat_0[1]),.dout(n194),.clk(gclk));
	jcb g109(.dina(n194),.dinb(w_dff_B_LXHGXDS25_1),.dout(n195));
	jand g110(.dina(w_dff_B_8rvGSJTv5_0),.dinb(n190),.dout(n196),.clk(gclk));
	jand g111(.dina(w_dff_B_yWnPKxVu2_0),.dinb(n182),.dout(n197),.clk(gclk));
	jxor g112(.dina(w_n197_0[2]),.dinb(w_n181_0[2]),.dout(n198),.clk(gclk));
	jand g113(.dina(w_n198_0[2]),.dinb(w_G228gat_3[1]),.dout(n199),.clk(gclk));
	jand g114(.dina(w_n173_0[0]),.dinb(w_G201gat_0[1]),.dout(n200),.clk(gclk));
	jand g115(.dina(w_n200_0[1]),.dinb(w_G237gat_3[1]),.dout(n201),.clk(gclk));
	jand g116(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n202),.clk(gclk));
	jand g117(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n203),.clk(gclk));
	jcb g118(.dina(n203),.dinb(n202),.dout(n204));
	jcb g119(.dina(w_dff_B_JkHntt2U0_0),.dinb(n201),.dout(n205));
	jcb g120(.dina(w_dff_B_9AOImXTe6_0),.dinb(n199),.dout(n206));
	jcb g121(.dina(n206),.dinb(w_dff_B_JNhqm3lS9_1),.dout(n207));
	jcb g122(.dina(w_n198_0[1]),.dinb(w_G261gat_0[2]),.dout(n208));
	jnot g123(.din(w_G261gat_0[1]),.dout(n209),.clk(gclk));
	jnot g124(.din(w_n198_0[0]),.dout(n210),.clk(gclk));
	jcb g125(.dina(n210),.dinb(w_n209_0[1]),.dout(n211));
	jand g126(.dina(n211),.dinb(w_G219gat_3[2]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_mOxQql009_1),.dout(n213),.clk(gclk));
	jcb g128(.dina(n213),.dinb(w_dff_B_5ygL2A6b4_1),.dout(G850gat));
	jand g129(.dina(w_n164_3[0]),.dinb(w_G111gat_0[1]),.dout(n215),.clk(gclk));
	jand g130(.dina(w_n170_1[0]),.dinb(w_G143gat_0[1]),.dout(n216),.clk(gclk));
	jcb g131(.dina(w_dff_B_tExV6k4Y7_0),.dinb(w_n148_1[0]),.dout(n217));
	jcb g132(.dina(n217),.dinb(n215),.dout(n218));
	jxor g133(.dina(w_n218_1[1]),.dinb(w_G183gat_1[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n219_0[2]),.dinb(w_G228gat_3[0]),.dout(n220),.clk(gclk));
	jand g135(.dina(w_n178_3[0]),.dinb(w_G183gat_1[0]),.dout(n221),.clk(gclk));
	jand g136(.dina(w_n218_1[0]),.dinb(w_G183gat_0[2]),.dout(n222),.clk(gclk));
	jand g137(.dina(w_n222_0[2]),.dinb(w_G237gat_3[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n218_0[2]),.dinb(w_G246gat_3[0]),.dout(n224),.clk(gclk));
	jand g139(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n225),.clk(gclk));
	jcb g140(.dina(w_dff_B_TciQSPIr2_0),.dinb(n224),.dout(n226));
	jcb g141(.dina(w_dff_B_abiyQRox7_0),.dinb(n223),.dout(n227));
	jcb g142(.dina(n227),.dinb(w_dff_B_FSdXD1d11_1),.dout(n228));
	jcb g143(.dina(n228),.dinb(n220),.dout(n229));
	jand g144(.dina(w_n164_2[2]),.dinb(w_G116gat_0[1]),.dout(n230),.clk(gclk));
	jand g145(.dina(w_n170_0[2]),.dinb(w_G146gat_0[1]),.dout(n231),.clk(gclk));
	jcb g146(.dina(w_dff_B_FqU1p9qq9_0),.dinb(w_n148_0[2]),.dout(n232));
	jcb g147(.dina(n232),.dinb(n230),.dout(n233));
	jand g148(.dina(w_n233_1[1]),.dinb(w_G189gat_2[0]),.dout(n234),.clk(gclk));
	jcb g149(.dina(w_n233_1[0]),.dinb(w_G189gat_1[2]),.dout(n235));
	jand g150(.dina(w_n164_2[1]),.dinb(w_G121gat_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n170_0[1]),.dinb(w_G149gat_0[1]),.dout(n237),.clk(gclk));
	jcb g152(.dina(w_dff_B_GZeGIeJg7_0),.dinb(w_n148_0[1]),.dout(n238));
	jcb g153(.dina(n238),.dinb(n236),.dout(n239));
	jand g154(.dina(w_n239_1[1]),.dinb(w_G195gat_2[0]),.dout(n240),.clk(gclk));
	jcb g155(.dina(w_n239_1[0]),.dinb(w_G195gat_1[2]),.dout(n241));
	jand g156(.dina(w_n197_0[1]),.dinb(w_n181_0[1]),.dout(n242),.clk(gclk));
	jnot g157(.din(w_n242_0[1]),.dout(n243),.clk(gclk));
	jcb g158(.dina(w_n200_0[0]),.dinb(w_G261gat_0[0]),.dout(n244));
	jand g159(.dina(w_dff_B_DWlw1QNO9_0),.dinb(n243),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n245_0[1]),.dinb(w_n241_0[1]),.dout(n246),.clk(gclk));
	jcb g161(.dina(n246),.dinb(w_n240_0[1]),.dout(n247));
	jand g162(.dina(w_n247_0[1]),.dinb(w_n235_0[1]),.dout(n248),.clk(gclk));
	jcb g163(.dina(n248),.dinb(w_n234_0[1]),.dout(n249));
	jcb g164(.dina(w_n249_0[1]),.dinb(w_n219_0[1]),.dout(n250));
	jnot g165(.din(w_n219_0[0]),.dout(n251),.clk(gclk));
	jnot g166(.din(w_n234_0[0]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n235_0[0]),.dout(n253),.clk(gclk));
	jnot g168(.din(w_n240_0[0]),.dout(n254),.clk(gclk));
	jnot g169(.din(w_n241_0[0]),.dout(n255),.clk(gclk));
	jcb g170(.dina(w_n197_0[0]),.dinb(w_n181_0[0]),.dout(n256));
	jand g171(.dina(n256),.dinb(w_n209_0[0]),.dout(n257),.clk(gclk));
	jcb g172(.dina(n257),.dinb(w_n242_0[0]),.dout(n258));
	jcb g173(.dina(w_n258_0[1]),.dinb(w_dff_B_KHqf8zhh8_1),.dout(n259));
	jand g174(.dina(n259),.dinb(w_dff_B_mlaOqiYt2_1),.dout(n260),.clk(gclk));
	jcb g175(.dina(w_n260_0[1]),.dinb(w_dff_B_qbt2vy6h2_1),.dout(n261));
	jand g176(.dina(n261),.dinb(w_dff_B_174OM27a1_1),.dout(n262),.clk(gclk));
	jcb g177(.dina(w_n262_0[1]),.dinb(w_dff_B_kw8OM5yr9_1),.dout(n263));
	jand g178(.dina(n263),.dinb(w_G219gat_3[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(w_dff_B_iVi9uWFn7_0),.dinb(n250),.dout(n265),.clk(gclk));
	jcb g180(.dina(n265),.dinb(w_dff_B_swztmzOe3_1),.dout(G863gat));
	jxor g181(.dina(w_n233_0[2]),.dinb(w_G189gat_1[1]),.dout(n267),.clk(gclk));
	jand g182(.dina(w_n267_0[2]),.dinb(w_G228gat_2[2]),.dout(n268),.clk(gclk));
	jand g183(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n269),.clk(gclk));
	jand g184(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n270),.clk(gclk));
	jcb g185(.dina(n270),.dinb(w_G246gat_2[2]),.dout(n271));
	jand g186(.dina(w_dff_B_YtZGeX4D6_0),.dinb(w_n233_0[1]),.dout(n272),.clk(gclk));
	jcb g187(.dina(n272),.dinb(w_dff_B_cbzNglHz5_1),.dout(n273));
	jand g188(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n274),.clk(gclk));
	jand g189(.dina(w_n178_2[2]),.dinb(w_G189gat_0[2]),.dout(n275),.clk(gclk));
	jcb g190(.dina(n275),.dinb(w_dff_B_GPFA6cjJ3_1),.dout(n276));
	jcb g191(.dina(w_dff_B_i5rM6Lyh2_0),.dinb(n273),.dout(n277));
	jcb g192(.dina(w_dff_B_w8J3QZD11_0),.dinb(n268),.dout(n278));
	jcb g193(.dina(w_n267_0[1]),.dinb(w_n247_0[0]),.dout(n279));
	jnot g194(.din(w_n267_0[0]),.dout(n280),.clk(gclk));
	jcb g195(.dina(w_dff_B_eRAyobKB9_0),.dinb(w_n260_0[0]),.dout(n281));
	jand g196(.dina(n281),.dinb(w_G219gat_3[0]),.dout(n282),.clk(gclk));
	jand g197(.dina(w_dff_B_9AB076ns0_0),.dinb(n279),.dout(n283),.clk(gclk));
	jcb g198(.dina(n283),.dinb(w_dff_B_KYyTr8kZ9_1),.dout(G864gat));
	jxor g199(.dina(w_n239_0[2]),.dinb(w_G195gat_1[1]),.dout(n285),.clk(gclk));
	jand g200(.dina(w_n285_0[2]),.dinb(w_G228gat_2[1]),.dout(n286),.clk(gclk));
	jand g201(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n287),.clk(gclk));
	jand g202(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n288),.clk(gclk));
	jcb g203(.dina(n288),.dinb(w_G246gat_2[1]),.dout(n289));
	jand g204(.dina(w_dff_B_NElr3muP5_0),.dinb(w_n239_0[1]),.dout(n290),.clk(gclk));
	jcb g205(.dina(n290),.dinb(w_dff_B_oZ2mumHy2_1),.dout(n291));
	jand g206(.dina(w_n178_2[1]),.dinb(w_G195gat_0[2]),.dout(n292),.clk(gclk));
	jand g207(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n293),.clk(gclk));
	jcb g208(.dina(w_dff_B_cxlGlZI51_0),.dinb(n292),.dout(n294));
	jcb g209(.dina(w_dff_B_4bUShkSf5_0),.dinb(n291),.dout(n295));
	jcb g210(.dina(w_dff_B_0iPckTON6_0),.dinb(n286),.dout(n296));
	jcb g211(.dina(w_n285_0[1]),.dinb(w_n245_0[0]),.dout(n297));
	jnot g212(.din(w_n285_0[0]),.dout(n298),.clk(gclk));
	jcb g213(.dina(w_dff_B_oFKigCyb2_0),.dinb(w_n258_0[0]),.dout(n299));
	jand g214(.dina(n299),.dinb(w_G219gat_2[2]),.dout(n300),.clk(gclk));
	jand g215(.dina(w_dff_B_LWzEiq9O1_0),.dinb(n297),.dout(n301),.clk(gclk));
	jcb g216(.dina(n301),.dinb(w_dff_B_FX7SA9iW4_1),.dout(G865gat));
	jand g217(.dina(w_n168_0[0]),.dinb(w_G55gat_0[0]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n303_1[1]),.dinb(w_G143gat_0[0]),.dout(n304),.clk(gclk));
	jand g219(.dina(w_n146_0[0]),.dinb(w_G17gat_1[0]),.dout(n305),.clk(gclk));
	jand g220(.dina(n305),.dinb(w_n144_0[0]),.dout(n306),.clk(gclk));
	jcb g221(.dina(w_n306_1[1]),.dinb(w_dff_B_OZFlQu3P9_1),.dout(n307));
	jand g222(.dina(w_n164_2[0]),.dinb(w_G91gat_0[1]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n309),.clk(gclk));
	jcb g224(.dina(w_dff_B_aI0lAFX63_0),.dinb(n308),.dout(n310));
	jcb g225(.dina(n310),.dinb(n307),.dout(n311));
	jand g226(.dina(w_n311_1[2]),.dinb(w_G159gat_1[1]),.dout(n312),.clk(gclk));
	jcb g227(.dina(w_n311_1[1]),.dinb(w_G159gat_1[0]),.dout(n313));
	jand g228(.dina(w_n164_1[2]),.dinb(w_G96gat_0[1]),.dout(n314),.clk(gclk));
	jand g229(.dina(w_n303_1[0]),.dinb(w_G146gat_0[0]),.dout(n315),.clk(gclk));
	jand g230(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n316),.clk(gclk));
	jcb g231(.dina(w_dff_B_9JrxwEvH3_0),.dinb(n315),.dout(n317));
	jcb g232(.dina(w_dff_B_zVjBrFHL1_0),.dinb(n314),.dout(n318));
	jcb g233(.dina(n318),.dinb(w_n306_1[0]),.dout(n319));
	jand g234(.dina(w_n319_1[2]),.dinb(w_G165gat_1[1]),.dout(n320),.clk(gclk));
	jcb g235(.dina(w_n319_1[1]),.dinb(w_G165gat_1[0]),.dout(n321));
	jand g236(.dina(w_n164_1[1]),.dinb(w_G101gat_0[1]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n303_0[2]),.dinb(w_G149gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n324),.clk(gclk));
	jcb g239(.dina(w_dff_B_MSQsjCHr1_0),.dinb(n323),.dout(n325));
	jcb g240(.dina(w_dff_B_aSMCM9EO5_0),.dinb(n322),.dout(n326));
	jcb g241(.dina(n326),.dinb(w_n306_0[2]),.dout(n327));
	jand g242(.dina(w_n327_1[2]),.dinb(w_G171gat_1[1]),.dout(n328),.clk(gclk));
	jcb g243(.dina(w_n327_1[1]),.dinb(w_G171gat_1[0]),.dout(n329));
	jand g244(.dina(w_n164_1[0]),.dinb(w_G106gat_0[0]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n303_0[1]),.dinb(w_G153gat_0[0]),.dout(n331),.clk(gclk));
	jand g246(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n332),.clk(gclk));
	jcb g247(.dina(w_dff_B_xfwW9Hcw6_0),.dinb(n331),.dout(n333));
	jcb g248(.dina(w_dff_B_Fdm4RsM11_0),.dinb(n330),.dout(n334));
	jcb g249(.dina(n334),.dinb(w_n306_0[1]),.dout(n335));
	jand g250(.dina(w_n335_1[1]),.dinb(w_G177gat_1[1]),.dout(n336),.clk(gclk));
	jnot g251(.din(w_G177gat_1[0]),.dout(n337),.clk(gclk));
	jnot g252(.din(w_n335_1[0]),.dout(n338),.clk(gclk));
	jand g253(.dina(n338),.dinb(w_dff_B_6NKaHX122_1),.dout(n339),.clk(gclk));
	jnot g254(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jnot g255(.din(w_G183gat_0[1]),.dout(n341),.clk(gclk));
	jnot g256(.din(w_n218_0[1]),.dout(n342),.clk(gclk));
	jand g257(.dina(n342),.dinb(w_dff_B_HC1jVCeB8_1),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n343_0[1]),.dout(n344),.clk(gclk));
	jand g259(.dina(w_n249_0[0]),.dinb(w_dff_B_CFs5Y1xx7_1),.dout(n345),.clk(gclk));
	jcb g260(.dina(n345),.dinb(w_n222_0[1]),.dout(n346));
	jand g261(.dina(w_n346_0[1]),.dinb(w_dff_B_fnNvb5kg5_1),.dout(n347),.clk(gclk));
	jcb g262(.dina(n347),.dinb(w_n336_0[2]),.dout(n348));
	jand g263(.dina(w_n348_0[1]),.dinb(w_n329_0[1]),.dout(n349),.clk(gclk));
	jcb g264(.dina(n349),.dinb(w_n328_0[1]),.dout(n350));
	jand g265(.dina(w_n350_0[1]),.dinb(w_n321_0[1]),.dout(n351),.clk(gclk));
	jcb g266(.dina(n351),.dinb(w_n320_0[1]),.dout(n352));
	jand g267(.dina(w_n352_0[1]),.dinb(w_dff_B_TDFpNZwg1_1),.dout(n353),.clk(gclk));
	jcb g268(.dina(n353),.dinb(w_dff_B_q2WYnYNi0_1),.dout(G866gat));
	jxor g269(.dina(w_n335_0[2]),.dinb(w_G177gat_0[2]),.dout(n355),.clk(gclk));
	jnot g270(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n346_0[0]),.dinb(w_G219gat_2[1]),.dout(n357),.clk(gclk));
	jand g272(.dina(n357),.dinb(w_dff_B_4d6awUTU5_1),.dout(n358),.clk(gclk));
	jnot g273(.din(w_n222_0[0]),.dout(n359),.clk(gclk));
	jcb g274(.dina(w_n262_0[0]),.dinb(w_n343_0[0]),.dout(n360));
	jand g275(.dina(n360),.dinb(w_dff_B_iQF2qdDc8_1),.dout(n361),.clk(gclk));
	jand g276(.dina(w_n361_0[1]),.dinb(w_G219gat_2[0]),.dout(n362),.clk(gclk));
	jcb g277(.dina(n362),.dinb(w_G228gat_2[0]),.dout(n363));
	jand g278(.dina(n363),.dinb(w_n355_0[0]),.dout(n364),.clk(gclk));
	jand g279(.dina(w_n336_0[1]),.dinb(w_G237gat_2[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_n335_0[1]),.dinb(w_G246gat_2[0]),.dout(n366),.clk(gclk));
	jand g281(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n367),.clk(gclk));
	jand g282(.dina(w_n178_2[0]),.dinb(w_G177gat_0[1]),.dout(n368),.clk(gclk));
	jcb g283(.dina(n368),.dinb(w_dff_B_aeJyEo2r6_1),.dout(n369));
	jcb g284(.dina(w_dff_B_Q9e22nuI2_0),.dinb(n366),.dout(n370));
	jcb g285(.dina(w_dff_B_xJNQDe2B7_0),.dinb(n365),.dout(n371));
	jcb g286(.dina(w_dff_B_y7IukNiW4_0),.dinb(n364),.dout(n372));
	jcb g287(.dina(w_dff_B_FuP7dzmg7_0),.dinb(n358),.dout(G874gat));
	jand g288(.dina(w_n311_1[0]),.dinb(w_G237gat_1[2]),.dout(n374),.clk(gclk));
	jcb g289(.dina(n374),.dinb(w_n178_1[2]),.dout(n375));
	jand g290(.dina(n375),.dinb(w_G159gat_0[2]),.dout(n376),.clk(gclk));
	jxor g291(.dina(w_n311_0[2]),.dinb(w_G159gat_0[1]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_n377_0[2]),.dinb(w_G228gat_1[2]),.dout(n378),.clk(gclk));
	jand g293(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n379),.clk(gclk));
	jcb g294(.dina(w_dff_B_6wNC4TZh8_0),.dinb(n378),.dout(n380));
	jand g295(.dina(w_n311_0[1]),.dinb(w_G246gat_1[2]),.dout(n381),.clk(gclk));
	jcb g296(.dina(w_dff_B_tQydU9YP5_0),.dinb(n380),.dout(n382));
	jcb g297(.dina(n382),.dinb(n376),.dout(n383));
	jcb g298(.dina(w_n377_0[1]),.dinb(w_n352_0[0]),.dout(n384));
	jnot g299(.din(w_n320_0[0]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n321_0[0]),.dout(n386),.clk(gclk));
	jnot g301(.din(w_n328_0[0]),.dout(n387),.clk(gclk));
	jnot g302(.din(w_n329_0[0]),.dout(n388),.clk(gclk));
	jnot g303(.din(w_n336_0[0]),.dout(n389),.clk(gclk));
	jcb g304(.dina(w_n361_0[0]),.dinb(w_n339_0[0]),.dout(n390));
	jand g305(.dina(n390),.dinb(w_dff_B_CfTfS9m79_1),.dout(n391),.clk(gclk));
	jcb g306(.dina(w_n391_0[1]),.dinb(w_dff_B_03IvlBp05_1),.dout(n392));
	jand g307(.dina(n392),.dinb(w_dff_B_vHnDE2rC4_1),.dout(n393),.clk(gclk));
	jcb g308(.dina(w_n393_0[1]),.dinb(w_dff_B_kQCU9bhP1_1),.dout(n394));
	jand g309(.dina(n394),.dinb(w_dff_B_TReuXL9t2_1),.dout(n395),.clk(gclk));
	jnot g310(.din(w_n377_0[0]),.dout(n396),.clk(gclk));
	jcb g311(.dina(w_dff_B_l3ntDq6M2_0),.dinb(n395),.dout(n397));
	jand g312(.dina(n397),.dinb(w_G219gat_1[2]),.dout(n398),.clk(gclk));
	jand g313(.dina(w_dff_B_a7I7qVPu9_0),.dinb(n384),.dout(n399),.clk(gclk));
	jcb g314(.dina(n399),.dinb(w_dff_B_WIoMev244_1),.dout(G878gat));
	jand g315(.dina(w_n319_1[0]),.dinb(w_G237gat_1[1]),.dout(n401),.clk(gclk));
	jcb g316(.dina(n401),.dinb(w_n178_1[1]),.dout(n402));
	jand g317(.dina(n402),.dinb(w_G165gat_0[2]),.dout(n403),.clk(gclk));
	jxor g318(.dina(w_n319_0[2]),.dinb(w_G165gat_0[1]),.dout(n404),.clk(gclk));
	jand g319(.dina(w_n404_0[2]),.dinb(w_G228gat_1[1]),.dout(n405),.clk(gclk));
	jand g320(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n406),.clk(gclk));
	jcb g321(.dina(w_dff_B_AXPtbETS2_0),.dinb(n405),.dout(n407));
	jand g322(.dina(w_n319_0[1]),.dinb(w_G246gat_1[1]),.dout(n408),.clk(gclk));
	jcb g323(.dina(w_dff_B_vZpFLVwD0_0),.dinb(n407),.dout(n409));
	jcb g324(.dina(n409),.dinb(n403),.dout(n410));
	jcb g325(.dina(w_n404_0[1]),.dinb(w_n350_0[0]),.dout(n411));
	jnot g326(.din(w_n404_0[0]),.dout(n412),.clk(gclk));
	jcb g327(.dina(w_dff_B_cG3Xjw698_0),.dinb(w_n393_0[0]),.dout(n413));
	jand g328(.dina(n413),.dinb(w_G219gat_1[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(w_dff_B_E5KRjqAt4_0),.dinb(n411),.dout(n415),.clk(gclk));
	jcb g330(.dina(n415),.dinb(w_dff_B_5EfUWnzb2_1),.dout(G879gat));
	jand g331(.dina(w_n327_1[0]),.dinb(w_G237gat_1[0]),.dout(n417),.clk(gclk));
	jcb g332(.dina(n417),.dinb(w_n178_1[0]),.dout(n418));
	jand g333(.dina(n418),.dinb(w_G171gat_0[2]),.dout(n419),.clk(gclk));
	jxor g334(.dina(w_n327_0[2]),.dinb(w_G171gat_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n420_0[2]),.dinb(w_G228gat_1[0]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jcb g337(.dina(w_dff_B_sKQwZKGO0_0),.dinb(n421),.dout(n423));
	jand g338(.dina(w_n327_0[1]),.dinb(w_G246gat_1[0]),.dout(n424),.clk(gclk));
	jcb g339(.dina(w_dff_B_viTRVlxQ2_0),.dinb(n423),.dout(n425));
	jcb g340(.dina(n425),.dinb(n419),.dout(n426));
	jnot g341(.din(w_n420_0[1]),.dout(n427),.clk(gclk));
	jcb g342(.dina(w_dff_B_mYze1cyB0_0),.dinb(w_n391_0[0]),.dout(n428));
	jcb g343(.dina(w_n420_0[0]),.dinb(w_n348_0[0]),.dout(n429));
	jand g344(.dina(n429),.dinb(w_G219gat_1[0]),.dout(n430),.clk(gclk));
	jand g345(.dina(n430),.dinb(w_dff_B_74NRWyks0_1),.dout(n431),.clk(gclk));
	jcb g346(.dina(n431),.dinb(w_dff_B_Jmt0lTr00_1),.dout(G880gat));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_iCl7TOn50_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_dff_A_hw9j201Q8_1),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_kGD97uD18_0),.doutb(w_dff_A_R3mMVGf93_1),.doutc(w_G17gat_1[2]),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_dff_A_8o2GDxRU3_2),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_U5kbN1Si1_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_Okid8rW94_1),.doutc(w_dff_A_tuOdJaz41_2),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_dff_A_XDrhQoL33_0),.doutb(w_G42gat_1[1]),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_tZhBeJBZ3_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_YW6fEiix2_0),.doutb(w_dff_A_nmfxa6Js2_1),.doutc(w_G55gat_0[2]),.din(w_dff_B_i5JhTpjB3_3));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_dff_A_7uPyF1rD4_1),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_75Zmf9AN2_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_2b6CFqz22_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_tVvGk56O2_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_jJ3Agiua5_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_5QQC5bE49_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_7RxM1HFo4_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_wbINvpvQ9_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_bWkaAc2M5_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_KyQsSQ0E2_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl3 jspl3_w_G126gat_0(.douta(w_G126gat_0[0]),.doutb(w_dff_A_zkfDkXYw9_1),.doutc(w_G126gat_0[2]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_dff_A_cdbfX95G2_1),.din(G130gat));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_G143gat_0[1]),.din(w_dff_B_9ieTWPER3_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_G146gat_0[1]),.din(w_dff_B_NSpcUwYz7_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_G149gat_0[1]),.din(w_dff_B_yWvWJbNP7_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_xpiSFEr42_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_5PsbKJ721_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_dff_A_R3hqFTFh7_1),.doutc(w_dff_A_upcNwBLK1_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_dff_A_K3St2tcO9_0),.doutb(w_dff_A_ZUppNKUk6_1),.doutc(w_G159gat_1[2]),.din(w_G159gat_0[0]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_dff_A_Tm74dXJS5_1),.doutc(w_dff_A_yqRDbJJ93_2),.din(w_dff_B_jhSL01uD2_3));
	jspl3 jspl3_w_G165gat_1(.douta(w_dff_A_wJ0ToPjs9_0),.doutb(w_dff_A_565O5jmn6_1),.doutc(w_G165gat_1[2]),.din(w_G165gat_0[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_dff_A_pkWdKiuy2_1),.doutc(w_dff_A_4MhYOLGE7_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_dff_A_YmakPBz43_0),.doutb(w_dff_A_xrAKoSCS0_1),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_dff_A_HocxKQJ23_1),.doutc(w_dff_A_rKopKHok9_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_lUNGMeER4_1),.doutc(w_G177gat_1[2]),.din(w_G177gat_0[0]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_SOYVUpiV3_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_0kLhHTXP1_0),.doutb(w_dff_A_l1YZ2Gd11_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_Lb4784C42_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_3VLFMT3U3_1),.doutc(w_dff_A_8cuxrSrU0_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_otoplOJD7_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_hB4lQznq7_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_U1w57x487_1),.doutc(w_dff_A_SYPybmbJ0_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_nYxAQpCt9_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_dff_A_wB7S1cRe7_1),.doutc(w_G201gat_0[2]),.din(G201gat));
	jspl jspl_w_G201gat_1(.douta(w_dff_A_l2oQh35B4_0),.doutb(w_G201gat_1[1]),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_zS1JG0L90_0),.doutb(w_G219gat_0[1]),.doutc(w_dff_A_trNkA0at5_2),.din(w_dff_B_wDGhJLLo9_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_dff_A_Wf2H0hlY2_0),.doutb(w_G219gat_1[1]),.doutc(w_dff_A_ZjTjFceJ6_2),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_RcBFuB6l7_0),.doutb(w_dff_A_jOiGhT7j7_1),.doutc(w_G219gat_2[2]),.din(w_G219gat_0[1]));
	jspl3 jspl3_w_G219gat_3(.douta(w_G219gat_3[0]),.doutb(w_dff_A_wWjTsjEO8_1),.doutc(w_G219gat_3[2]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_G228gat_0[0]),.doutb(w_G228gat_0[1]),.doutc(w_G228gat_0[2]),.din(w_dff_B_PKDSliMz0_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_dff_A_SEYXpYpz4_0),.doutb(w_G228gat_2[1]),.doutc(w_G228gat_2[2]),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_dff_A_8YjeJZ702_1),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_dff_A_3StBpSnb5_0),.doutb(w_G237gat_0[1]),.doutc(w_dff_A_DwycHNr98_2),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_dff_A_JfoasXjw1_0),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_G237gat_3[1]),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_dff_A_XvYe7sEs4_0),.doutb(w_G246gat_0[1]),.doutc(w_dff_A_dio62ymb4_2),.din(w_dff_B_ML60B5756_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_dff_A_CGl3dEfJ4_0),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_G246gat_3[1]),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_7wpFEAVr2_0),.doutb(w_G261gat_0[1]),.doutc(w_dff_A_Xvcckb5q5_2),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_G390gat_0[1]),.doutc(G390gat),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_dff_A_GzPcAlQd1_2),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(G447gat),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_dff_A_8YW7iErV4_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.doutc(w_n95_0[2]),.din(n95));
	jspl jspl_w_n97_0(.douta(w_dff_A_AwLQZzfH2_0),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_dff_A_GrE8512v4_0),.doutb(w_n101_0[1]),.din(w_dff_B_Kxz2Dri24_2));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_CGqpf3Ic4_1),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.din(n113));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_dff_A_Cw9lnBBc6_1),.din(n122));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_nqtVZAax0_2));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_n148_1[0]),.doutb(w_n148_1[1]),.doutc(w_n148_1[2]),.din(w_n148_0[0]));
	jspl jspl_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.din(n149));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_EuLMJAVz8_1),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl3 jspl3_w_n164_1(.douta(w_n164_1[0]),.doutb(w_n164_1[1]),.doutc(w_n164_1[2]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n164_2(.douta(w_n164_2[0]),.doutb(w_n164_2[1]),.doutc(w_n164_2[2]),.din(w_n164_0[1]));
	jspl jspl_w_n164_3(.douta(w_n164_3[0]),.doutb(w_n164_3[1]),.din(w_n164_0[2]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_dOndz9hd4_1),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n170_1(.douta(w_n170_1[0]),.doutb(w_n170_1[1]),.din(w_n170_0[0]));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_xHTspfHT1_0),.doutb(w_n178_0[1]),.doutc(w_n178_0[2]),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n178_2(.douta(w_n178_2[0]),.doutb(w_n178_2[1]),.doutc(w_n178_2[2]),.din(w_n178_0[1]));
	jspl jspl_w_n178_3(.douta(w_n178_3[0]),.doutb(w_n178_3[1]),.din(w_n178_0[2]));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(w_dff_B_aeLYM4i55_3));
	jspl jspl_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.din(n185));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_ksjfY7GK7_1),.din(w_dff_B_tgNJEoev1_2));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl jspl_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_AkCmnQQX5_1),.doutc(w_n219_0[2]),.din(n219));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_dff_A_gnhZkBHY0_1),.doutc(w_n222_0[2]),.din(n222));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_dff_A_vVTloqkZ2_1),.din(n234));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_dff_A_LqsTnaKk6_1),.din(n235));
	jspl3 jspl3_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.doutc(w_n239_0[2]),.din(n239));
	jspl jspl_w_n239_1(.douta(w_n239_1[0]),.doutb(w_n239_1[1]),.din(w_n239_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_dff_A_gblR4WM46_1),.din(n240));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_dff_A_OPWn0AdZ8_1),.din(n241));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.din(n258));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_dff_A_R43HBhu72_1),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_dff_A_vSxnLJ9U6_1),.doutc(w_n285_0[2]),.din(n285));
	jspl3 jspl3_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.doutc(w_n303_0[2]),.din(n303));
	jspl jspl_w_n303_1(.douta(w_n303_1[0]),.doutb(w_n303_1[1]),.din(w_n303_0[0]));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.doutc(w_n306_0[2]),.din(n306));
	jspl jspl_w_n306_1(.douta(w_n306_1[0]),.doutb(w_n306_1[1]),.din(w_n306_0[0]));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.doutc(w_n311_0[2]),.din(n311));
	jspl3 jspl3_w_n311_1(.douta(w_n311_1[0]),.doutb(w_n311_1[1]),.doutc(w_n311_1[2]),.din(w_n311_0[0]));
	jspl3 jspl3_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.doutc(w_n319_0[2]),.din(n319));
	jspl3 jspl3_w_n319_1(.douta(w_n319_1[0]),.doutb(w_n319_1[1]),.doutc(w_n319_1[2]),.din(w_n319_0[0]));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_dff_A_tSEJwimh4_1),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_FEZopSkl9_1),.din(n321));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl3 jspl3_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.doutc(w_n327_1[2]),.din(w_n327_0[0]));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_dff_A_fQNP7HS99_1),.din(n328));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_dff_A_zqrSmoA51_1),.din(n329));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl jspl_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.din(w_n335_0[0]));
	jspl3 jspl3_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.doutc(w_dff_A_8pmlUdXC8_2),.din(n336));
	jspl jspl_w_n339_0(.douta(w_dff_A_6ChR3N6F0_0),.doutb(w_n339_0[1]),.din(n339));
	jspl jspl_w_n343_0(.douta(w_dff_A_Uex1Sy8D9_0),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.din(n352));
	jspl jspl_w_n355_0(.douta(w_dff_A_bDGdhnR76_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_J9C4nb5O7_1),.doutc(w_n377_0[2]),.din(n377));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_dff_A_QBszpqbZ2_1),.doutc(w_n404_0[2]),.din(n404));
	jspl3 jspl3_w_n420_0(.douta(w_dff_A_pXiBHGgW9_0),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jdff dff_A_CGqpf3Ic4_1(.dout(w_n103_0[1]),.din(w_dff_A_CGqpf3Ic4_1),.clk(gclk));
	jdff dff_A_GrE8512v4_0(.dout(w_n101_0[0]),.din(w_dff_A_GrE8512v4_0),.clk(gclk));
	jdff dff_B_Kxz2Dri24_2(.din(n101),.dout(w_dff_B_Kxz2Dri24_2),.clk(gclk));
	jdff dff_B_MUHJqlsa3_1(.din(G74gat),.dout(w_dff_B_MUHJqlsa3_1),.clk(gclk));
	jdff dff_B_D5KQVx4N8_1(.din(w_dff_B_MUHJqlsa3_1),.dout(w_dff_B_D5KQVx4N8_1),.clk(gclk));
	jdff dff_B_IMJTrLm56_1(.din(w_dff_B_D5KQVx4N8_1),.dout(w_dff_B_IMJTrLm56_1),.clk(gclk));
	jdff dff_B_kltv1uDD9_1(.din(n127),.dout(w_dff_B_kltv1uDD9_1),.clk(gclk));
	jdff dff_B_SWsBNjgP5_1(.din(G135gat),.dout(w_dff_B_SWsBNjgP5_1),.clk(gclk));
	jdff dff_B_SwAJvB7p8_1(.din(n136),.dout(w_dff_B_SwAJvB7p8_1),.clk(gclk));
	jdff dff_A_cdbfX95G2_1(.dout(w_G130gat_0[1]),.din(w_dff_A_cdbfX95G2_1),.clk(gclk));
	jdff dff_B_TPcV03838_1(.din(G207gat),.dout(w_dff_B_TPcV03838_1),.clk(gclk));
	jdff dff_B_8q5RoEtf6_1(.din(n207),.dout(w_dff_B_8q5RoEtf6_1),.clk(gclk));
	jdff dff_B_5ygL2A6b4_1(.din(w_dff_B_8q5RoEtf6_1),.dout(w_dff_B_5ygL2A6b4_1),.clk(gclk));
	jdff dff_B_atjGC3YD0_1(.din(n208),.dout(w_dff_B_atjGC3YD0_1),.clk(gclk));
	jdff dff_B_mOxQql009_1(.din(w_dff_B_atjGC3YD0_1),.dout(w_dff_B_mOxQql009_1),.clk(gclk));
	jdff dff_B_HNfNVR8z4_1(.din(n180),.dout(w_dff_B_HNfNVR8z4_1),.clk(gclk));
	jdff dff_B_sYsY2Xrd2_1(.din(w_dff_B_HNfNVR8z4_1),.dout(w_dff_B_sYsY2Xrd2_1),.clk(gclk));
	jdff dff_B_JNhqm3lS9_1(.din(w_dff_B_sYsY2Xrd2_1),.dout(w_dff_B_JNhqm3lS9_1),.clk(gclk));
	jdff dff_B_Tc3tWnSk6_0(.din(n205),.dout(w_dff_B_Tc3tWnSk6_0),.clk(gclk));
	jdff dff_B_9AOImXTe6_0(.din(w_dff_B_Tc3tWnSk6_0),.dout(w_dff_B_9AOImXTe6_0),.clk(gclk));
	jdff dff_B_18Whazdq0_0(.din(n204),.dout(w_dff_B_18Whazdq0_0),.clk(gclk));
	jdff dff_B_mmVXoTq22_0(.din(w_dff_B_18Whazdq0_0),.dout(w_dff_B_mmVXoTq22_0),.clk(gclk));
	jdff dff_B_9clIZ1G66_0(.din(w_dff_B_mmVXoTq22_0),.dout(w_dff_B_9clIZ1G66_0),.clk(gclk));
	jdff dff_B_i4hGdTD60_0(.din(w_dff_B_9clIZ1G66_0),.dout(w_dff_B_i4hGdTD60_0),.clk(gclk));
	jdff dff_B_x2sN5suX5_0(.din(w_dff_B_i4hGdTD60_0),.dout(w_dff_B_x2sN5suX5_0),.clk(gclk));
	jdff dff_B_mSd8cxZv9_0(.din(w_dff_B_x2sN5suX5_0),.dout(w_dff_B_mSd8cxZv9_0),.clk(gclk));
	jdff dff_B_JkHntt2U0_0(.din(w_dff_B_mSd8cxZv9_0),.dout(w_dff_B_JkHntt2U0_0),.clk(gclk));
	jdff dff_B_nzh4t6dO4_0(.din(n179),.dout(w_dff_B_nzh4t6dO4_0),.clk(gclk));
	jdff dff_B_KDBSoOv51_0(.din(w_dff_B_nzh4t6dO4_0),.dout(w_dff_B_KDBSoOv51_0),.clk(gclk));
	jdff dff_A_kcSaOgBj7_0(.dout(w_G201gat_1[0]),.din(w_dff_A_kcSaOgBj7_0),.clk(gclk));
	jdff dff_A_eOmbkkKK7_0(.dout(w_dff_A_kcSaOgBj7_0),.din(w_dff_A_eOmbkkKK7_0),.clk(gclk));
	jdff dff_A_ZJAKB7245_0(.dout(w_dff_A_eOmbkkKK7_0),.din(w_dff_A_ZJAKB7245_0),.clk(gclk));
	jdff dff_A_l2oQh35B4_0(.dout(w_dff_A_ZJAKB7245_0),.din(w_dff_A_l2oQh35B4_0),.clk(gclk));
	jdff dff_B_c76GNu681_1(.din(n229),.dout(w_dff_B_c76GNu681_1),.clk(gclk));
	jdff dff_B_VXEXTzTa3_1(.din(w_dff_B_c76GNu681_1),.dout(w_dff_B_VXEXTzTa3_1),.clk(gclk));
	jdff dff_B_twHoBtLm8_1(.din(w_dff_B_VXEXTzTa3_1),.dout(w_dff_B_twHoBtLm8_1),.clk(gclk));
	jdff dff_B_G23ZZq9F9_1(.din(w_dff_B_twHoBtLm8_1),.dout(w_dff_B_G23ZZq9F9_1),.clk(gclk));
	jdff dff_B_mPC2hAMR7_1(.din(w_dff_B_G23ZZq9F9_1),.dout(w_dff_B_mPC2hAMR7_1),.clk(gclk));
	jdff dff_B_swztmzOe3_1(.din(w_dff_B_mPC2hAMR7_1),.dout(w_dff_B_swztmzOe3_1),.clk(gclk));
	jdff dff_B_iVi9uWFn7_0(.din(n264),.dout(w_dff_B_iVi9uWFn7_0),.clk(gclk));
	jdff dff_B_vd8DefqJ3_1(.din(n251),.dout(w_dff_B_vd8DefqJ3_1),.clk(gclk));
	jdff dff_B_FEjPi52X4_1(.din(w_dff_B_vd8DefqJ3_1),.dout(w_dff_B_FEjPi52X4_1),.clk(gclk));
	jdff dff_B_kw8OM5yr9_1(.din(w_dff_B_FEjPi52X4_1),.dout(w_dff_B_kw8OM5yr9_1),.clk(gclk));
	jdff dff_B_mdY2YZjG4_1(.din(n221),.dout(w_dff_B_mdY2YZjG4_1),.clk(gclk));
	jdff dff_B_4sjJETFE3_1(.din(w_dff_B_mdY2YZjG4_1),.dout(w_dff_B_4sjJETFE3_1),.clk(gclk));
	jdff dff_B_FSdXD1d11_1(.din(w_dff_B_4sjJETFE3_1),.dout(w_dff_B_FSdXD1d11_1),.clk(gclk));
	jdff dff_B_abiyQRox7_0(.din(n226),.dout(w_dff_B_abiyQRox7_0),.clk(gclk));
	jdff dff_B_nUltx7Tg2_0(.din(n225),.dout(w_dff_B_nUltx7Tg2_0),.clk(gclk));
	jdff dff_B_sMTwHmq87_0(.din(w_dff_B_nUltx7Tg2_0),.dout(w_dff_B_sMTwHmq87_0),.clk(gclk));
	jdff dff_B_BM4PMVxL2_0(.din(w_dff_B_sMTwHmq87_0),.dout(w_dff_B_BM4PMVxL2_0),.clk(gclk));
	jdff dff_B_XYVWrlwg0_0(.din(w_dff_B_BM4PMVxL2_0),.dout(w_dff_B_XYVWrlwg0_0),.clk(gclk));
	jdff dff_B_peq3b0pW1_0(.din(w_dff_B_XYVWrlwg0_0),.dout(w_dff_B_peq3b0pW1_0),.clk(gclk));
	jdff dff_B_TciQSPIr2_0(.din(w_dff_B_peq3b0pW1_0),.dout(w_dff_B_TciQSPIr2_0),.clk(gclk));
	jdff dff_A_RTB5cNrH8_1(.dout(w_n219_0[1]),.din(w_dff_A_RTB5cNrH8_1),.clk(gclk));
	jdff dff_A_lT5BDjlx9_1(.dout(w_dff_A_RTB5cNrH8_1),.din(w_dff_A_lT5BDjlx9_1),.clk(gclk));
	jdff dff_A_7L9LTNAp1_1(.dout(w_dff_A_lT5BDjlx9_1),.din(w_dff_A_7L9LTNAp1_1),.clk(gclk));
	jdff dff_A_JhTgU0BS8_1(.dout(w_dff_A_7L9LTNAp1_1),.din(w_dff_A_JhTgU0BS8_1),.clk(gclk));
	jdff dff_A_ag8uLg3T9_1(.dout(w_dff_A_JhTgU0BS8_1),.din(w_dff_A_ag8uLg3T9_1),.clk(gclk));
	jdff dff_A_AkCmnQQX5_1(.dout(w_dff_A_ag8uLg3T9_1),.din(w_dff_A_AkCmnQQX5_1),.clk(gclk));
	jdff dff_A_TQi4cZKh2_0(.dout(w_G183gat_1[0]),.din(w_dff_A_TQi4cZKh2_0),.clk(gclk));
	jdff dff_A_dg5UlAL93_0(.dout(w_dff_A_TQi4cZKh2_0),.din(w_dff_A_dg5UlAL93_0),.clk(gclk));
	jdff dff_A_6qMOCYBK6_0(.dout(w_dff_A_dg5UlAL93_0),.din(w_dff_A_6qMOCYBK6_0),.clk(gclk));
	jdff dff_A_0kLhHTXP1_0(.dout(w_dff_A_6qMOCYBK6_0),.din(w_dff_A_0kLhHTXP1_0),.clk(gclk));
	jdff dff_A_cbz4fwcC7_1(.dout(w_G183gat_1[1]),.din(w_dff_A_cbz4fwcC7_1),.clk(gclk));
	jdff dff_A_YtPcYc5j3_1(.dout(w_dff_A_cbz4fwcC7_1),.din(w_dff_A_YtPcYc5j3_1),.clk(gclk));
	jdff dff_A_3EFehQgQ5_1(.dout(w_dff_A_YtPcYc5j3_1),.din(w_dff_A_3EFehQgQ5_1),.clk(gclk));
	jdff dff_A_QPAVvka71_1(.dout(w_dff_A_3EFehQgQ5_1),.din(w_dff_A_QPAVvka71_1),.clk(gclk));
	jdff dff_A_fHSpneZv5_1(.dout(w_dff_A_QPAVvka71_1),.din(w_dff_A_fHSpneZv5_1),.clk(gclk));
	jdff dff_A_l1YZ2Gd11_1(.dout(w_dff_A_fHSpneZv5_1),.din(w_dff_A_l1YZ2Gd11_1),.clk(gclk));
	jdff dff_A_GZUfWPL59_1(.dout(w_G228gat_3[1]),.din(w_dff_A_GZUfWPL59_1),.clk(gclk));
	jdff dff_A_8YjeJZ702_1(.dout(w_dff_A_GZUfWPL59_1),.din(w_dff_A_8YjeJZ702_1),.clk(gclk));
	jdff dff_B_vfrcgtj62_1(.din(n278),.dout(w_dff_B_vfrcgtj62_1),.clk(gclk));
	jdff dff_B_hpvNr7mY4_1(.din(w_dff_B_vfrcgtj62_1),.dout(w_dff_B_hpvNr7mY4_1),.clk(gclk));
	jdff dff_B_Qc5Ep4Et7_1(.din(w_dff_B_hpvNr7mY4_1),.dout(w_dff_B_Qc5Ep4Et7_1),.clk(gclk));
	jdff dff_B_mSYXw8eD5_1(.din(w_dff_B_Qc5Ep4Et7_1),.dout(w_dff_B_mSYXw8eD5_1),.clk(gclk));
	jdff dff_B_KYyTr8kZ9_1(.din(w_dff_B_mSYXw8eD5_1),.dout(w_dff_B_KYyTr8kZ9_1),.clk(gclk));
	jdff dff_B_9AB076ns0_0(.din(n282),.dout(w_dff_B_9AB076ns0_0),.clk(gclk));
	jdff dff_B_4IHM62Q08_0(.din(n280),.dout(w_dff_B_4IHM62Q08_0),.clk(gclk));
	jdff dff_B_eRAyobKB9_0(.din(w_dff_B_4IHM62Q08_0),.dout(w_dff_B_eRAyobKB9_0),.clk(gclk));
	jdff dff_A_wWjTsjEO8_1(.dout(w_G219gat_3[1]),.din(w_dff_A_wWjTsjEO8_1),.clk(gclk));
	jdff dff_B_w8J3QZD11_0(.din(n277),.dout(w_dff_B_w8J3QZD11_0),.clk(gclk));
	jdff dff_B_6pBXQl0J0_0(.din(n276),.dout(w_dff_B_6pBXQl0J0_0),.clk(gclk));
	jdff dff_B_i5rM6Lyh2_0(.din(w_dff_B_6pBXQl0J0_0),.dout(w_dff_B_i5rM6Lyh2_0),.clk(gclk));
	jdff dff_B_8bO6AFix8_1(.din(n274),.dout(w_dff_B_8bO6AFix8_1),.clk(gclk));
	jdff dff_B_Mhj4yigo2_1(.din(w_dff_B_8bO6AFix8_1),.dout(w_dff_B_Mhj4yigo2_1),.clk(gclk));
	jdff dff_B_5vQ5oGUA7_1(.din(w_dff_B_Mhj4yigo2_1),.dout(w_dff_B_5vQ5oGUA7_1),.clk(gclk));
	jdff dff_B_GPFA6cjJ3_1(.din(w_dff_B_5vQ5oGUA7_1),.dout(w_dff_B_GPFA6cjJ3_1),.clk(gclk));
	jdff dff_B_qcuLo3QQ8_1(.din(n269),.dout(w_dff_B_qcuLo3QQ8_1),.clk(gclk));
	jdff dff_B_7UHTb3y94_1(.din(w_dff_B_qcuLo3QQ8_1),.dout(w_dff_B_7UHTb3y94_1),.clk(gclk));
	jdff dff_B_z8ELfjDw5_1(.din(w_dff_B_7UHTb3y94_1),.dout(w_dff_B_z8ELfjDw5_1),.clk(gclk));
	jdff dff_B_OpAWbcsq9_1(.din(w_dff_B_z8ELfjDw5_1),.dout(w_dff_B_OpAWbcsq9_1),.clk(gclk));
	jdff dff_B_Fg1Gbfcy3_1(.din(w_dff_B_OpAWbcsq9_1),.dout(w_dff_B_Fg1Gbfcy3_1),.clk(gclk));
	jdff dff_B_cbzNglHz5_1(.din(w_dff_B_Fg1Gbfcy3_1),.dout(w_dff_B_cbzNglHz5_1),.clk(gclk));
	jdff dff_B_tLVV8sgM8_0(.din(n271),.dout(w_dff_B_tLVV8sgM8_0),.clk(gclk));
	jdff dff_B_ty9Yyy5w2_0(.din(w_dff_B_tLVV8sgM8_0),.dout(w_dff_B_ty9Yyy5w2_0),.clk(gclk));
	jdff dff_B_AOlezAnq9_0(.din(w_dff_B_ty9Yyy5w2_0),.dout(w_dff_B_AOlezAnq9_0),.clk(gclk));
	jdff dff_B_D1nOBTit1_0(.din(w_dff_B_AOlezAnq9_0),.dout(w_dff_B_D1nOBTit1_0),.clk(gclk));
	jdff dff_B_YtZGeX4D6_0(.din(w_dff_B_D1nOBTit1_0),.dout(w_dff_B_YtZGeX4D6_0),.clk(gclk));
	jdff dff_A_DzFSMGnM2_1(.dout(w_n267_0[1]),.din(w_dff_A_DzFSMGnM2_1),.clk(gclk));
	jdff dff_A_s39czw265_1(.dout(w_dff_A_DzFSMGnM2_1),.din(w_dff_A_s39czw265_1),.clk(gclk));
	jdff dff_A_7O3U6y6e2_1(.dout(w_dff_A_s39czw265_1),.din(w_dff_A_7O3U6y6e2_1),.clk(gclk));
	jdff dff_A_QFejvGR19_1(.dout(w_dff_A_7O3U6y6e2_1),.din(w_dff_A_QFejvGR19_1),.clk(gclk));
	jdff dff_A_R43HBhu72_1(.dout(w_dff_A_QFejvGR19_1),.din(w_dff_A_R43HBhu72_1),.clk(gclk));
	jdff dff_B_cAjIsP5b6_1(.din(n296),.dout(w_dff_B_cAjIsP5b6_1),.clk(gclk));
	jdff dff_B_Ger2NZoh9_1(.din(w_dff_B_cAjIsP5b6_1),.dout(w_dff_B_Ger2NZoh9_1),.clk(gclk));
	jdff dff_B_fGvbyBJA5_1(.din(w_dff_B_Ger2NZoh9_1),.dout(w_dff_B_fGvbyBJA5_1),.clk(gclk));
	jdff dff_B_FX7SA9iW4_1(.din(w_dff_B_fGvbyBJA5_1),.dout(w_dff_B_FX7SA9iW4_1),.clk(gclk));
	jdff dff_B_LWzEiq9O1_0(.din(n300),.dout(w_dff_B_LWzEiq9O1_0),.clk(gclk));
	jdff dff_B_oFKigCyb2_0(.din(n298),.dout(w_dff_B_oFKigCyb2_0),.clk(gclk));
	jdff dff_B_0iPckTON6_0(.din(n295),.dout(w_dff_B_0iPckTON6_0),.clk(gclk));
	jdff dff_B_5tk9Ng485_0(.din(n294),.dout(w_dff_B_5tk9Ng485_0),.clk(gclk));
	jdff dff_B_4bUShkSf5_0(.din(w_dff_B_5tk9Ng485_0),.dout(w_dff_B_4bUShkSf5_0),.clk(gclk));
	jdff dff_B_QeLuuleW6_0(.din(n293),.dout(w_dff_B_QeLuuleW6_0),.clk(gclk));
	jdff dff_B_ZfyCljN99_0(.din(w_dff_B_QeLuuleW6_0),.dout(w_dff_B_ZfyCljN99_0),.clk(gclk));
	jdff dff_B_jshBZBSI7_0(.din(w_dff_B_ZfyCljN99_0),.dout(w_dff_B_jshBZBSI7_0),.clk(gclk));
	jdff dff_B_cxlGlZI51_0(.din(w_dff_B_jshBZBSI7_0),.dout(w_dff_B_cxlGlZI51_0),.clk(gclk));
	jdff dff_B_qoyXegVq0_1(.din(n287),.dout(w_dff_B_qoyXegVq0_1),.clk(gclk));
	jdff dff_B_IVrEZG6f2_1(.din(w_dff_B_qoyXegVq0_1),.dout(w_dff_B_IVrEZG6f2_1),.clk(gclk));
	jdff dff_B_B3ass3li8_1(.din(w_dff_B_IVrEZG6f2_1),.dout(w_dff_B_B3ass3li8_1),.clk(gclk));
	jdff dff_B_pHz2bQjf1_1(.din(w_dff_B_B3ass3li8_1),.dout(w_dff_B_pHz2bQjf1_1),.clk(gclk));
	jdff dff_B_28Pg7Chg7_1(.din(w_dff_B_pHz2bQjf1_1),.dout(w_dff_B_28Pg7Chg7_1),.clk(gclk));
	jdff dff_B_oZ2mumHy2_1(.din(w_dff_B_28Pg7Chg7_1),.dout(w_dff_B_oZ2mumHy2_1),.clk(gclk));
	jdff dff_B_gLxFFouQ5_0(.din(n289),.dout(w_dff_B_gLxFFouQ5_0),.clk(gclk));
	jdff dff_B_KUqZWgip8_0(.din(w_dff_B_gLxFFouQ5_0),.dout(w_dff_B_KUqZWgip8_0),.clk(gclk));
	jdff dff_B_FssnNeB03_0(.din(w_dff_B_KUqZWgip8_0),.dout(w_dff_B_FssnNeB03_0),.clk(gclk));
	jdff dff_B_F7CSIpNA6_0(.din(w_dff_B_FssnNeB03_0),.dout(w_dff_B_F7CSIpNA6_0),.clk(gclk));
	jdff dff_B_NElr3muP5_0(.din(w_dff_B_F7CSIpNA6_0),.dout(w_dff_B_NElr3muP5_0),.clk(gclk));
	jdff dff_A_d7Xsperi1_1(.dout(w_n285_0[1]),.din(w_dff_A_d7Xsperi1_1),.clk(gclk));
	jdff dff_A_hjd6GLBh9_1(.dout(w_dff_A_d7Xsperi1_1),.din(w_dff_A_hjd6GLBh9_1),.clk(gclk));
	jdff dff_A_Bf1tSGQD0_1(.dout(w_dff_A_hjd6GLBh9_1),.din(w_dff_A_Bf1tSGQD0_1),.clk(gclk));
	jdff dff_A_vSxnLJ9U6_1(.dout(w_dff_A_Bf1tSGQD0_1),.din(w_dff_A_vSxnLJ9U6_1),.clk(gclk));
	jdff dff_B_9qzIs8wg5_1(.din(n312),.dout(w_dff_B_9qzIs8wg5_1),.clk(gclk));
	jdff dff_B_3a3WQmmx7_1(.din(w_dff_B_9qzIs8wg5_1),.dout(w_dff_B_3a3WQmmx7_1),.clk(gclk));
	jdff dff_B_q0XmMZTp5_1(.din(w_dff_B_3a3WQmmx7_1),.dout(w_dff_B_q0XmMZTp5_1),.clk(gclk));
	jdff dff_B_f4uRBHLF5_1(.din(w_dff_B_q0XmMZTp5_1),.dout(w_dff_B_f4uRBHLF5_1),.clk(gclk));
	jdff dff_B_ulRN76xC9_1(.din(w_dff_B_f4uRBHLF5_1),.dout(w_dff_B_ulRN76xC9_1),.clk(gclk));
	jdff dff_B_nduxFZnu9_1(.din(w_dff_B_ulRN76xC9_1),.dout(w_dff_B_nduxFZnu9_1),.clk(gclk));
	jdff dff_B_t3ezegcD5_1(.din(w_dff_B_nduxFZnu9_1),.dout(w_dff_B_t3ezegcD5_1),.clk(gclk));
	jdff dff_B_UNokS3si3_1(.din(w_dff_B_t3ezegcD5_1),.dout(w_dff_B_UNokS3si3_1),.clk(gclk));
	jdff dff_B_CBRBtQeq6_1(.din(w_dff_B_UNokS3si3_1),.dout(w_dff_B_CBRBtQeq6_1),.clk(gclk));
	jdff dff_B_WlG0mSKq4_1(.din(w_dff_B_CBRBtQeq6_1),.dout(w_dff_B_WlG0mSKq4_1),.clk(gclk));
	jdff dff_B_q2WYnYNi0_1(.din(w_dff_B_WlG0mSKq4_1),.dout(w_dff_B_q2WYnYNi0_1),.clk(gclk));
	jdff dff_B_FGgtUkCF1_1(.din(n313),.dout(w_dff_B_FGgtUkCF1_1),.clk(gclk));
	jdff dff_B_Dsin8gAB5_1(.din(w_dff_B_FGgtUkCF1_1),.dout(w_dff_B_Dsin8gAB5_1),.clk(gclk));
	jdff dff_B_0kJwRmP97_1(.din(w_dff_B_Dsin8gAB5_1),.dout(w_dff_B_0kJwRmP97_1),.clk(gclk));
	jdff dff_B_iGT7ybQT9_1(.din(w_dff_B_0kJwRmP97_1),.dout(w_dff_B_iGT7ybQT9_1),.clk(gclk));
	jdff dff_B_OcC37nY42_1(.din(w_dff_B_iGT7ybQT9_1),.dout(w_dff_B_OcC37nY42_1),.clk(gclk));
	jdff dff_B_dCPzLgYM7_1(.din(w_dff_B_OcC37nY42_1),.dout(w_dff_B_dCPzLgYM7_1),.clk(gclk));
	jdff dff_B_Aji7Bi1B0_1(.din(w_dff_B_dCPzLgYM7_1),.dout(w_dff_B_Aji7Bi1B0_1),.clk(gclk));
	jdff dff_B_iOYwoYdk4_1(.din(w_dff_B_Aji7Bi1B0_1),.dout(w_dff_B_iOYwoYdk4_1),.clk(gclk));
	jdff dff_B_dRqKBnj94_1(.din(w_dff_B_iOYwoYdk4_1),.dout(w_dff_B_dRqKBnj94_1),.clk(gclk));
	jdff dff_B_o1wsCmzP6_1(.din(w_dff_B_dRqKBnj94_1),.dout(w_dff_B_o1wsCmzP6_1),.clk(gclk));
	jdff dff_B_TDFpNZwg1_1(.din(w_dff_B_o1wsCmzP6_1),.dout(w_dff_B_TDFpNZwg1_1),.clk(gclk));
	jdff dff_A_dCMo2yu14_0(.dout(w_G159gat_1[0]),.din(w_dff_A_dCMo2yu14_0),.clk(gclk));
	jdff dff_A_HNKnGvbD6_0(.dout(w_dff_A_dCMo2yu14_0),.din(w_dff_A_HNKnGvbD6_0),.clk(gclk));
	jdff dff_A_w1A9S7e51_0(.dout(w_dff_A_HNKnGvbD6_0),.din(w_dff_A_w1A9S7e51_0),.clk(gclk));
	jdff dff_A_LwAixRhC6_0(.dout(w_dff_A_w1A9S7e51_0),.din(w_dff_A_LwAixRhC6_0),.clk(gclk));
	jdff dff_A_EuFvweOY7_0(.dout(w_dff_A_LwAixRhC6_0),.din(w_dff_A_EuFvweOY7_0),.clk(gclk));
	jdff dff_A_K3St2tcO9_0(.dout(w_dff_A_EuFvweOY7_0),.din(w_dff_A_K3St2tcO9_0),.clk(gclk));
	jdff dff_A_qIS9NgnR5_1(.dout(w_G159gat_1[1]),.din(w_dff_A_qIS9NgnR5_1),.clk(gclk));
	jdff dff_A_CDGiNcbs7_1(.dout(w_dff_A_qIS9NgnR5_1),.din(w_dff_A_CDGiNcbs7_1),.clk(gclk));
	jdff dff_A_0VuttSU13_1(.dout(w_dff_A_CDGiNcbs7_1),.din(w_dff_A_0VuttSU13_1),.clk(gclk));
	jdff dff_A_rCUEQCJY8_1(.dout(w_dff_A_0VuttSU13_1),.din(w_dff_A_rCUEQCJY8_1),.clk(gclk));
	jdff dff_A_Y0wwgnqY3_1(.dout(w_dff_A_rCUEQCJY8_1),.din(w_dff_A_Y0wwgnqY3_1),.clk(gclk));
	jdff dff_A_ZUppNKUk6_1(.dout(w_dff_A_Y0wwgnqY3_1),.din(w_dff_A_ZUppNKUk6_1),.clk(gclk));
	jdff dff_B_9LrSJ0Kr3_0(.din(n372),.dout(w_dff_B_9LrSJ0Kr3_0),.clk(gclk));
	jdff dff_B_FuP7dzmg7_0(.din(w_dff_B_9LrSJ0Kr3_0),.dout(w_dff_B_FuP7dzmg7_0),.clk(gclk));
	jdff dff_B_Mdi0xSTC6_0(.din(n371),.dout(w_dff_B_Mdi0xSTC6_0),.clk(gclk));
	jdff dff_B_FLIDAsOS3_0(.din(w_dff_B_Mdi0xSTC6_0),.dout(w_dff_B_FLIDAsOS3_0),.clk(gclk));
	jdff dff_B_mvBzfZ2u9_0(.din(w_dff_B_FLIDAsOS3_0),.dout(w_dff_B_mvBzfZ2u9_0),.clk(gclk));
	jdff dff_B_Nfcr0bzR3_0(.din(w_dff_B_mvBzfZ2u9_0),.dout(w_dff_B_Nfcr0bzR3_0),.clk(gclk));
	jdff dff_B_kSGpyvbW1_0(.din(w_dff_B_Nfcr0bzR3_0),.dout(w_dff_B_kSGpyvbW1_0),.clk(gclk));
	jdff dff_B_y7IukNiW4_0(.din(w_dff_B_kSGpyvbW1_0),.dout(w_dff_B_y7IukNiW4_0),.clk(gclk));
	jdff dff_B_xJNQDe2B7_0(.din(n370),.dout(w_dff_B_xJNQDe2B7_0),.clk(gclk));
	jdff dff_B_5e3LN8Mb1_0(.din(n369),.dout(w_dff_B_5e3LN8Mb1_0),.clk(gclk));
	jdff dff_B_Q9e22nuI2_0(.din(w_dff_B_5e3LN8Mb1_0),.dout(w_dff_B_Q9e22nuI2_0),.clk(gclk));
	jdff dff_B_W8HFDH5P9_1(.din(n367),.dout(w_dff_B_W8HFDH5P9_1),.clk(gclk));
	jdff dff_B_1JMh91Xp6_1(.din(w_dff_B_W8HFDH5P9_1),.dout(w_dff_B_1JMh91Xp6_1),.clk(gclk));
	jdff dff_B_jbJW216R2_1(.din(w_dff_B_1JMh91Xp6_1),.dout(w_dff_B_jbJW216R2_1),.clk(gclk));
	jdff dff_B_aeJyEo2r6_1(.din(w_dff_B_jbJW216R2_1),.dout(w_dff_B_aeJyEo2r6_1),.clk(gclk));
	jdff dff_A_982UkWgj0_0(.dout(w_G246gat_2[0]),.din(w_dff_A_982UkWgj0_0),.clk(gclk));
	jdff dff_A_0RAZQmfo6_0(.dout(w_dff_A_982UkWgj0_0),.din(w_dff_A_0RAZQmfo6_0),.clk(gclk));
	jdff dff_A_VcS46n8X2_0(.dout(w_dff_A_0RAZQmfo6_0),.din(w_dff_A_VcS46n8X2_0),.clk(gclk));
	jdff dff_A_7MmasVGu5_0(.dout(w_dff_A_VcS46n8X2_0),.din(w_dff_A_7MmasVGu5_0),.clk(gclk));
	jdff dff_A_CGl3dEfJ4_0(.dout(w_dff_A_7MmasVGu5_0),.din(w_dff_A_CGl3dEfJ4_0),.clk(gclk));
	jdff dff_A_LbkBKiXU0_0(.dout(w_G237gat_2[0]),.din(w_dff_A_LbkBKiXU0_0),.clk(gclk));
	jdff dff_A_SaVK1kLN8_0(.dout(w_dff_A_LbkBKiXU0_0),.din(w_dff_A_SaVK1kLN8_0),.clk(gclk));
	jdff dff_A_rNMfhchC8_0(.dout(w_dff_A_SaVK1kLN8_0),.din(w_dff_A_rNMfhchC8_0),.clk(gclk));
	jdff dff_A_S7Avvjfk1_0(.dout(w_dff_A_rNMfhchC8_0),.din(w_dff_A_S7Avvjfk1_0),.clk(gclk));
	jdff dff_A_dy2TlCbN1_0(.dout(w_dff_A_S7Avvjfk1_0),.din(w_dff_A_dy2TlCbN1_0),.clk(gclk));
	jdff dff_A_c1NVpzwA2_0(.dout(w_dff_A_dy2TlCbN1_0),.din(w_dff_A_c1NVpzwA2_0),.clk(gclk));
	jdff dff_A_JfoasXjw1_0(.dout(w_dff_A_c1NVpzwA2_0),.din(w_dff_A_JfoasXjw1_0),.clk(gclk));
	jdff dff_A_loYMBPnY5_0(.dout(w_G228gat_2[0]),.din(w_dff_A_loYMBPnY5_0),.clk(gclk));
	jdff dff_A_OQxJnndM3_0(.dout(w_dff_A_loYMBPnY5_0),.din(w_dff_A_OQxJnndM3_0),.clk(gclk));
	jdff dff_A_FMMyHLc56_0(.dout(w_dff_A_OQxJnndM3_0),.din(w_dff_A_FMMyHLc56_0),.clk(gclk));
	jdff dff_A_hLNHqSZs7_0(.dout(w_dff_A_FMMyHLc56_0),.din(w_dff_A_hLNHqSZs7_0),.clk(gclk));
	jdff dff_A_Z5EfJoiX1_0(.dout(w_dff_A_hLNHqSZs7_0),.din(w_dff_A_Z5EfJoiX1_0),.clk(gclk));
	jdff dff_A_SEYXpYpz4_0(.dout(w_dff_A_Z5EfJoiX1_0),.din(w_dff_A_SEYXpYpz4_0),.clk(gclk));
	jdff dff_B_Pgydenyu2_1(.din(n356),.dout(w_dff_B_Pgydenyu2_1),.clk(gclk));
	jdff dff_B_kigoaMPV8_1(.din(w_dff_B_Pgydenyu2_1),.dout(w_dff_B_kigoaMPV8_1),.clk(gclk));
	jdff dff_B_ua5mdZHW7_1(.din(w_dff_B_kigoaMPV8_1),.dout(w_dff_B_ua5mdZHW7_1),.clk(gclk));
	jdff dff_B_tIB9YUQI7_1(.din(w_dff_B_ua5mdZHW7_1),.dout(w_dff_B_tIB9YUQI7_1),.clk(gclk));
	jdff dff_B_Gryezse61_1(.din(w_dff_B_tIB9YUQI7_1),.dout(w_dff_B_Gryezse61_1),.clk(gclk));
	jdff dff_B_wHdF1m8M7_1(.din(w_dff_B_Gryezse61_1),.dout(w_dff_B_wHdF1m8M7_1),.clk(gclk));
	jdff dff_B_4d6awUTU5_1(.din(w_dff_B_wHdF1m8M7_1),.dout(w_dff_B_4d6awUTU5_1),.clk(gclk));
	jdff dff_A_NWvFy5Hw2_0(.dout(w_G219gat_2[0]),.din(w_dff_A_NWvFy5Hw2_0),.clk(gclk));
	jdff dff_A_Sdlj9REF0_0(.dout(w_dff_A_NWvFy5Hw2_0),.din(w_dff_A_Sdlj9REF0_0),.clk(gclk));
	jdff dff_A_RcBFuB6l7_0(.dout(w_dff_A_Sdlj9REF0_0),.din(w_dff_A_RcBFuB6l7_0),.clk(gclk));
	jdff dff_A_lFqBu8ff3_1(.dout(w_G219gat_2[1]),.din(w_dff_A_lFqBu8ff3_1),.clk(gclk));
	jdff dff_A_CIR6gLEO2_1(.dout(w_dff_A_lFqBu8ff3_1),.din(w_dff_A_CIR6gLEO2_1),.clk(gclk));
	jdff dff_A_yyLGguNy6_1(.dout(w_dff_A_CIR6gLEO2_1),.din(w_dff_A_yyLGguNy6_1),.clk(gclk));
	jdff dff_A_nKSADduP4_1(.dout(w_dff_A_yyLGguNy6_1),.din(w_dff_A_nKSADduP4_1),.clk(gclk));
	jdff dff_A_jOiGhT7j7_1(.dout(w_dff_A_nKSADduP4_1),.din(w_dff_A_jOiGhT7j7_1),.clk(gclk));
	jdff dff_A_dN2iwtJG6_0(.dout(w_n355_0[0]),.din(w_dff_A_dN2iwtJG6_0),.clk(gclk));
	jdff dff_A_tuWIrX232_0(.dout(w_dff_A_dN2iwtJG6_0),.din(w_dff_A_tuWIrX232_0),.clk(gclk));
	jdff dff_A_3nDModQ05_0(.dout(w_dff_A_tuWIrX232_0),.din(w_dff_A_3nDModQ05_0),.clk(gclk));
	jdff dff_A_6uVQRxkF7_0(.dout(w_dff_A_3nDModQ05_0),.din(w_dff_A_6uVQRxkF7_0),.clk(gclk));
	jdff dff_A_xCGh9Dik9_0(.dout(w_dff_A_6uVQRxkF7_0),.din(w_dff_A_xCGh9Dik9_0),.clk(gclk));
	jdff dff_A_bDGdhnR76_0(.dout(w_dff_A_xCGh9Dik9_0),.din(w_dff_A_bDGdhnR76_0),.clk(gclk));
	jdff dff_B_LdfayXuk2_1(.din(n383),.dout(w_dff_B_LdfayXuk2_1),.clk(gclk));
	jdff dff_B_0zEf7tRx3_1(.din(w_dff_B_LdfayXuk2_1),.dout(w_dff_B_0zEf7tRx3_1),.clk(gclk));
	jdff dff_B_idbxuYqm5_1(.din(w_dff_B_0zEf7tRx3_1),.dout(w_dff_B_idbxuYqm5_1),.clk(gclk));
	jdff dff_B_QB7OndPV7_1(.din(w_dff_B_idbxuYqm5_1),.dout(w_dff_B_QB7OndPV7_1),.clk(gclk));
	jdff dff_B_fZ38KBMZ0_1(.din(w_dff_B_QB7OndPV7_1),.dout(w_dff_B_fZ38KBMZ0_1),.clk(gclk));
	jdff dff_B_HFDlZuMX4_1(.din(w_dff_B_fZ38KBMZ0_1),.dout(w_dff_B_HFDlZuMX4_1),.clk(gclk));
	jdff dff_B_1JMPf21u8_1(.din(w_dff_B_HFDlZuMX4_1),.dout(w_dff_B_1JMPf21u8_1),.clk(gclk));
	jdff dff_B_r008HAdm7_1(.din(w_dff_B_1JMPf21u8_1),.dout(w_dff_B_r008HAdm7_1),.clk(gclk));
	jdff dff_B_qMihiaua6_1(.din(w_dff_B_r008HAdm7_1),.dout(w_dff_B_qMihiaua6_1),.clk(gclk));
	jdff dff_B_WIoMev244_1(.din(w_dff_B_qMihiaua6_1),.dout(w_dff_B_WIoMev244_1),.clk(gclk));
	jdff dff_B_a7I7qVPu9_0(.din(n398),.dout(w_dff_B_a7I7qVPu9_0),.clk(gclk));
	jdff dff_B_ADo2BB3P8_0(.din(n396),.dout(w_dff_B_ADo2BB3P8_0),.clk(gclk));
	jdff dff_B_hjgrIZ3j7_0(.din(w_dff_B_ADo2BB3P8_0),.dout(w_dff_B_hjgrIZ3j7_0),.clk(gclk));
	jdff dff_B_qjgcuFW77_0(.din(w_dff_B_hjgrIZ3j7_0),.dout(w_dff_B_qjgcuFW77_0),.clk(gclk));
	jdff dff_B_yiPhGhBJ3_0(.din(w_dff_B_qjgcuFW77_0),.dout(w_dff_B_yiPhGhBJ3_0),.clk(gclk));
	jdff dff_B_0h0mUdec1_0(.din(w_dff_B_yiPhGhBJ3_0),.dout(w_dff_B_0h0mUdec1_0),.clk(gclk));
	jdff dff_B_zTmpkxaA7_0(.din(w_dff_B_0h0mUdec1_0),.dout(w_dff_B_zTmpkxaA7_0),.clk(gclk));
	jdff dff_B_l3ntDq6M2_0(.din(w_dff_B_zTmpkxaA7_0),.dout(w_dff_B_l3ntDq6M2_0),.clk(gclk));
	jdff dff_B_WzdsCEQ61_1(.din(n385),.dout(w_dff_B_WzdsCEQ61_1),.clk(gclk));
	jdff dff_B_wOXiouiC2_1(.din(w_dff_B_WzdsCEQ61_1),.dout(w_dff_B_wOXiouiC2_1),.clk(gclk));
	jdff dff_B_1LLCSq9R4_1(.din(w_dff_B_wOXiouiC2_1),.dout(w_dff_B_1LLCSq9R4_1),.clk(gclk));
	jdff dff_B_rNEezTIS7_1(.din(w_dff_B_1LLCSq9R4_1),.dout(w_dff_B_rNEezTIS7_1),.clk(gclk));
	jdff dff_B_ZwnIq4qE3_1(.din(w_dff_B_rNEezTIS7_1),.dout(w_dff_B_ZwnIq4qE3_1),.clk(gclk));
	jdff dff_B_TReuXL9t2_1(.din(w_dff_B_ZwnIq4qE3_1),.dout(w_dff_B_TReuXL9t2_1),.clk(gclk));
	jdff dff_B_VAcRZKeS7_1(.din(n386),.dout(w_dff_B_VAcRZKeS7_1),.clk(gclk));
	jdff dff_B_WIKRwLFC7_1(.din(w_dff_B_VAcRZKeS7_1),.dout(w_dff_B_WIKRwLFC7_1),.clk(gclk));
	jdff dff_B_Fv3rBYbU3_1(.din(w_dff_B_WIKRwLFC7_1),.dout(w_dff_B_Fv3rBYbU3_1),.clk(gclk));
	jdff dff_B_tR9RhVxv1_1(.din(w_dff_B_Fv3rBYbU3_1),.dout(w_dff_B_tR9RhVxv1_1),.clk(gclk));
	jdff dff_B_oWFtll3n6_1(.din(w_dff_B_tR9RhVxv1_1),.dout(w_dff_B_oWFtll3n6_1),.clk(gclk));
	jdff dff_B_MQp7jTcs0_1(.din(w_dff_B_oWFtll3n6_1),.dout(w_dff_B_MQp7jTcs0_1),.clk(gclk));
	jdff dff_B_kQCU9bhP1_1(.din(w_dff_B_MQp7jTcs0_1),.dout(w_dff_B_kQCU9bhP1_1),.clk(gclk));
	jdff dff_A_Lw2nkXRA7_1(.dout(w_n321_0[1]),.din(w_dff_A_Lw2nkXRA7_1),.clk(gclk));
	jdff dff_A_2psb8fgB0_1(.dout(w_dff_A_Lw2nkXRA7_1),.din(w_dff_A_2psb8fgB0_1),.clk(gclk));
	jdff dff_A_ZW9u7zkC4_1(.dout(w_dff_A_2psb8fgB0_1),.din(w_dff_A_ZW9u7zkC4_1),.clk(gclk));
	jdff dff_A_VsPrxV389_1(.dout(w_dff_A_ZW9u7zkC4_1),.din(w_dff_A_VsPrxV389_1),.clk(gclk));
	jdff dff_A_ntaRptit4_1(.dout(w_dff_A_VsPrxV389_1),.din(w_dff_A_ntaRptit4_1),.clk(gclk));
	jdff dff_A_Ixj01O2b5_1(.dout(w_dff_A_ntaRptit4_1),.din(w_dff_A_Ixj01O2b5_1),.clk(gclk));
	jdff dff_A_1EgNIh4p0_1(.dout(w_dff_A_Ixj01O2b5_1),.din(w_dff_A_1EgNIh4p0_1),.clk(gclk));
	jdff dff_A_SHhAVmmh8_1(.dout(w_dff_A_1EgNIh4p0_1),.din(w_dff_A_SHhAVmmh8_1),.clk(gclk));
	jdff dff_A_T11TeQpQ0_1(.dout(w_dff_A_SHhAVmmh8_1),.din(w_dff_A_T11TeQpQ0_1),.clk(gclk));
	jdff dff_A_FEZopSkl9_1(.dout(w_dff_A_T11TeQpQ0_1),.din(w_dff_A_FEZopSkl9_1),.clk(gclk));
	jdff dff_A_Vfj7nTLU6_1(.dout(w_n320_0[1]),.din(w_dff_A_Vfj7nTLU6_1),.clk(gclk));
	jdff dff_A_uGUfn8pZ9_1(.dout(w_dff_A_Vfj7nTLU6_1),.din(w_dff_A_uGUfn8pZ9_1),.clk(gclk));
	jdff dff_A_OZAPhxzk8_1(.dout(w_dff_A_uGUfn8pZ9_1),.din(w_dff_A_OZAPhxzk8_1),.clk(gclk));
	jdff dff_A_xsg5iuCv3_1(.dout(w_dff_A_OZAPhxzk8_1),.din(w_dff_A_xsg5iuCv3_1),.clk(gclk));
	jdff dff_A_58KaghXt5_1(.dout(w_dff_A_xsg5iuCv3_1),.din(w_dff_A_58KaghXt5_1),.clk(gclk));
	jdff dff_A_QSLRiiCz1_1(.dout(w_dff_A_58KaghXt5_1),.din(w_dff_A_QSLRiiCz1_1),.clk(gclk));
	jdff dff_A_2iUk5Bju8_1(.dout(w_dff_A_QSLRiiCz1_1),.din(w_dff_A_2iUk5Bju8_1),.clk(gclk));
	jdff dff_A_Jc707j8k5_1(.dout(w_dff_A_2iUk5Bju8_1),.din(w_dff_A_Jc707j8k5_1),.clk(gclk));
	jdff dff_A_sopswqjr8_1(.dout(w_dff_A_Jc707j8k5_1),.din(w_dff_A_sopswqjr8_1),.clk(gclk));
	jdff dff_A_tSEJwimh4_1(.dout(w_dff_A_sopswqjr8_1),.din(w_dff_A_tSEJwimh4_1),.clk(gclk));
	jdff dff_A_WWdNkkQo7_0(.dout(w_G165gat_1[0]),.din(w_dff_A_WWdNkkQo7_0),.clk(gclk));
	jdff dff_A_6aj3ALzR6_0(.dout(w_dff_A_WWdNkkQo7_0),.din(w_dff_A_6aj3ALzR6_0),.clk(gclk));
	jdff dff_A_WKqgjHLf1_0(.dout(w_dff_A_6aj3ALzR6_0),.din(w_dff_A_WKqgjHLf1_0),.clk(gclk));
	jdff dff_A_mGkyNChX3_0(.dout(w_dff_A_WKqgjHLf1_0),.din(w_dff_A_mGkyNChX3_0),.clk(gclk));
	jdff dff_A_wJ0ToPjs9_0(.dout(w_dff_A_mGkyNChX3_0),.din(w_dff_A_wJ0ToPjs9_0),.clk(gclk));
	jdff dff_A_RIOFRY1c3_1(.dout(w_G165gat_1[1]),.din(w_dff_A_RIOFRY1c3_1),.clk(gclk));
	jdff dff_A_61SjS4mf6_1(.dout(w_dff_A_RIOFRY1c3_1),.din(w_dff_A_61SjS4mf6_1),.clk(gclk));
	jdff dff_A_UJ4GzRM53_1(.dout(w_dff_A_61SjS4mf6_1),.din(w_dff_A_UJ4GzRM53_1),.clk(gclk));
	jdff dff_A_VznsKQfu4_1(.dout(w_dff_A_UJ4GzRM53_1),.din(w_dff_A_VznsKQfu4_1),.clk(gclk));
	jdff dff_A_565O5jmn6_1(.dout(w_dff_A_VznsKQfu4_1),.din(w_dff_A_565O5jmn6_1),.clk(gclk));
	jdff dff_B_tQydU9YP5_0(.din(n381),.dout(w_dff_B_tQydU9YP5_0),.clk(gclk));
	jdff dff_B_Dkm7EISG0_0(.din(n379),.dout(w_dff_B_Dkm7EISG0_0),.clk(gclk));
	jdff dff_B_KD5l42ko3_0(.din(w_dff_B_Dkm7EISG0_0),.dout(w_dff_B_KD5l42ko3_0),.clk(gclk));
	jdff dff_B_f5EXtC6H9_0(.din(w_dff_B_KD5l42ko3_0),.dout(w_dff_B_f5EXtC6H9_0),.clk(gclk));
	jdff dff_B_Zb0KeNRc4_0(.din(w_dff_B_f5EXtC6H9_0),.dout(w_dff_B_Zb0KeNRc4_0),.clk(gclk));
	jdff dff_B_XlqSPRHB8_0(.din(w_dff_B_Zb0KeNRc4_0),.dout(w_dff_B_XlqSPRHB8_0),.clk(gclk));
	jdff dff_B_ykhVGkkf7_0(.din(w_dff_B_XlqSPRHB8_0),.dout(w_dff_B_ykhVGkkf7_0),.clk(gclk));
	jdff dff_B_6wNC4TZh8_0(.din(w_dff_B_ykhVGkkf7_0),.dout(w_dff_B_6wNC4TZh8_0),.clk(gclk));
	jdff dff_A_oDjmOo787_1(.dout(w_n377_0[1]),.din(w_dff_A_oDjmOo787_1),.clk(gclk));
	jdff dff_A_4YXFuWR95_1(.dout(w_dff_A_oDjmOo787_1),.din(w_dff_A_4YXFuWR95_1),.clk(gclk));
	jdff dff_A_Rtb4ygeS1_1(.dout(w_dff_A_4YXFuWR95_1),.din(w_dff_A_Rtb4ygeS1_1),.clk(gclk));
	jdff dff_A_5dzD6IV28_1(.dout(w_dff_A_Rtb4ygeS1_1),.din(w_dff_A_5dzD6IV28_1),.clk(gclk));
	jdff dff_A_Sti2pNHY4_1(.dout(w_dff_A_5dzD6IV28_1),.din(w_dff_A_Sti2pNHY4_1),.clk(gclk));
	jdff dff_A_0gJUaOWj9_1(.dout(w_dff_A_Sti2pNHY4_1),.din(w_dff_A_0gJUaOWj9_1),.clk(gclk));
	jdff dff_A_UpJRFN434_1(.dout(w_dff_A_0gJUaOWj9_1),.din(w_dff_A_UpJRFN434_1),.clk(gclk));
	jdff dff_A_LOMqImEe6_1(.dout(w_dff_A_UpJRFN434_1),.din(w_dff_A_LOMqImEe6_1),.clk(gclk));
	jdff dff_A_c1UHsm5x5_1(.dout(w_dff_A_LOMqImEe6_1),.din(w_dff_A_c1UHsm5x5_1),.clk(gclk));
	jdff dff_A_J9C4nb5O7_1(.dout(w_dff_A_c1UHsm5x5_1),.din(w_dff_A_J9C4nb5O7_1),.clk(gclk));
	jdff dff_B_yanJwCB44_0(.din(n309),.dout(w_dff_B_yanJwCB44_0),.clk(gclk));
	jdff dff_B_c6refnxp3_0(.din(w_dff_B_yanJwCB44_0),.dout(w_dff_B_c6refnxp3_0),.clk(gclk));
	jdff dff_B_LUQVtbp02_0(.din(w_dff_B_c6refnxp3_0),.dout(w_dff_B_LUQVtbp02_0),.clk(gclk));
	jdff dff_B_cI2qUmAb1_0(.din(w_dff_B_LUQVtbp02_0),.dout(w_dff_B_cI2qUmAb1_0),.clk(gclk));
	jdff dff_B_aI0lAFX63_0(.din(w_dff_B_cI2qUmAb1_0),.dout(w_dff_B_aI0lAFX63_0),.clk(gclk));
	jdff dff_B_OZFlQu3P9_1(.din(n304),.dout(w_dff_B_OZFlQu3P9_1),.clk(gclk));
	jdff dff_A_sF7pYkdu3_1(.dout(w_G159gat_0[1]),.din(w_dff_A_sF7pYkdu3_1),.clk(gclk));
	jdff dff_A_36UdQolH2_1(.dout(w_dff_A_sF7pYkdu3_1),.din(w_dff_A_36UdQolH2_1),.clk(gclk));
	jdff dff_A_ZSdgoZUi4_1(.dout(w_dff_A_36UdQolH2_1),.din(w_dff_A_ZSdgoZUi4_1),.clk(gclk));
	jdff dff_A_8WD9Ab1h0_1(.dout(w_dff_A_ZSdgoZUi4_1),.din(w_dff_A_8WD9Ab1h0_1),.clk(gclk));
	jdff dff_A_cXx4m2f19_1(.dout(w_dff_A_8WD9Ab1h0_1),.din(w_dff_A_cXx4m2f19_1),.clk(gclk));
	jdff dff_A_R3hqFTFh7_1(.dout(w_dff_A_cXx4m2f19_1),.din(w_dff_A_R3hqFTFh7_1),.clk(gclk));
	jdff dff_A_07ktnM4N1_2(.dout(w_G159gat_0[2]),.din(w_dff_A_07ktnM4N1_2),.clk(gclk));
	jdff dff_A_p7sELI7H8_2(.dout(w_dff_A_07ktnM4N1_2),.din(w_dff_A_p7sELI7H8_2),.clk(gclk));
	jdff dff_A_sKT9uFrm1_2(.dout(w_dff_A_p7sELI7H8_2),.din(w_dff_A_sKT9uFrm1_2),.clk(gclk));
	jdff dff_A_LYRp8ABC4_2(.dout(w_dff_A_sKT9uFrm1_2),.din(w_dff_A_LYRp8ABC4_2),.clk(gclk));
	jdff dff_A_MdwO1Gv75_2(.dout(w_dff_A_LYRp8ABC4_2),.din(w_dff_A_MdwO1Gv75_2),.clk(gclk));
	jdff dff_A_OYECsV1Y5_2(.dout(w_dff_A_MdwO1Gv75_2),.din(w_dff_A_OYECsV1Y5_2),.clk(gclk));
	jdff dff_A_upcNwBLK1_2(.dout(w_dff_A_OYECsV1Y5_2),.din(w_dff_A_upcNwBLK1_2),.clk(gclk));
	jdff dff_B_rW1EU6Te4_1(.din(n410),.dout(w_dff_B_rW1EU6Te4_1),.clk(gclk));
	jdff dff_B_EyTziCDF9_1(.din(w_dff_B_rW1EU6Te4_1),.dout(w_dff_B_EyTziCDF9_1),.clk(gclk));
	jdff dff_B_OBzCZk2W9_1(.din(w_dff_B_EyTziCDF9_1),.dout(w_dff_B_OBzCZk2W9_1),.clk(gclk));
	jdff dff_B_wEdu6AHF8_1(.din(w_dff_B_OBzCZk2W9_1),.dout(w_dff_B_wEdu6AHF8_1),.clk(gclk));
	jdff dff_B_MssoguAC5_1(.din(w_dff_B_wEdu6AHF8_1),.dout(w_dff_B_MssoguAC5_1),.clk(gclk));
	jdff dff_B_72sKcRBa7_1(.din(w_dff_B_MssoguAC5_1),.dout(w_dff_B_72sKcRBa7_1),.clk(gclk));
	jdff dff_B_BqekfUUL7_1(.din(w_dff_B_72sKcRBa7_1),.dout(w_dff_B_BqekfUUL7_1),.clk(gclk));
	jdff dff_B_woM3vRP19_1(.din(w_dff_B_BqekfUUL7_1),.dout(w_dff_B_woM3vRP19_1),.clk(gclk));
	jdff dff_B_5EfUWnzb2_1(.din(w_dff_B_woM3vRP19_1),.dout(w_dff_B_5EfUWnzb2_1),.clk(gclk));
	jdff dff_B_E5KRjqAt4_0(.din(n414),.dout(w_dff_B_E5KRjqAt4_0),.clk(gclk));
	jdff dff_B_PpYIByju5_0(.din(n412),.dout(w_dff_B_PpYIByju5_0),.clk(gclk));
	jdff dff_B_DjiXcTp32_0(.din(w_dff_B_PpYIByju5_0),.dout(w_dff_B_DjiXcTp32_0),.clk(gclk));
	jdff dff_B_qrNMyGa71_0(.din(w_dff_B_DjiXcTp32_0),.dout(w_dff_B_qrNMyGa71_0),.clk(gclk));
	jdff dff_B_bsbK8xZW9_0(.din(w_dff_B_qrNMyGa71_0),.dout(w_dff_B_bsbK8xZW9_0),.clk(gclk));
	jdff dff_B_Zbk6Cu6J0_0(.din(w_dff_B_bsbK8xZW9_0),.dout(w_dff_B_Zbk6Cu6J0_0),.clk(gclk));
	jdff dff_B_cG3Xjw698_0(.din(w_dff_B_Zbk6Cu6J0_0),.dout(w_dff_B_cG3Xjw698_0),.clk(gclk));
	jdff dff_B_mOUJgLFa0_1(.din(n387),.dout(w_dff_B_mOUJgLFa0_1),.clk(gclk));
	jdff dff_B_bNUevt1G2_1(.din(w_dff_B_mOUJgLFa0_1),.dout(w_dff_B_bNUevt1G2_1),.clk(gclk));
	jdff dff_B_dXgHK3Yp3_1(.din(w_dff_B_bNUevt1G2_1),.dout(w_dff_B_dXgHK3Yp3_1),.clk(gclk));
	jdff dff_B_cZMYYE268_1(.din(w_dff_B_dXgHK3Yp3_1),.dout(w_dff_B_cZMYYE268_1),.clk(gclk));
	jdff dff_B_vHnDE2rC4_1(.din(w_dff_B_cZMYYE268_1),.dout(w_dff_B_vHnDE2rC4_1),.clk(gclk));
	jdff dff_B_QkKGhZt22_1(.din(n388),.dout(w_dff_B_QkKGhZt22_1),.clk(gclk));
	jdff dff_B_rk1a4uK05_1(.din(w_dff_B_QkKGhZt22_1),.dout(w_dff_B_rk1a4uK05_1),.clk(gclk));
	jdff dff_B_h1z0VhRv5_1(.din(w_dff_B_rk1a4uK05_1),.dout(w_dff_B_h1z0VhRv5_1),.clk(gclk));
	jdff dff_B_7R8VIzpJ5_1(.din(w_dff_B_h1z0VhRv5_1),.dout(w_dff_B_7R8VIzpJ5_1),.clk(gclk));
	jdff dff_B_IfJ9V8Iv0_1(.din(w_dff_B_7R8VIzpJ5_1),.dout(w_dff_B_IfJ9V8Iv0_1),.clk(gclk));
	jdff dff_B_03IvlBp05_1(.din(w_dff_B_IfJ9V8Iv0_1),.dout(w_dff_B_03IvlBp05_1),.clk(gclk));
	jdff dff_A_SPHf5gbO2_1(.dout(w_n329_0[1]),.din(w_dff_A_SPHf5gbO2_1),.clk(gclk));
	jdff dff_A_mS5cLRA47_1(.dout(w_dff_A_SPHf5gbO2_1),.din(w_dff_A_mS5cLRA47_1),.clk(gclk));
	jdff dff_A_mGtiqhbr3_1(.dout(w_dff_A_mS5cLRA47_1),.din(w_dff_A_mGtiqhbr3_1),.clk(gclk));
	jdff dff_A_zbMvYBGP4_1(.dout(w_dff_A_mGtiqhbr3_1),.din(w_dff_A_zbMvYBGP4_1),.clk(gclk));
	jdff dff_A_hHCAGVJo6_1(.dout(w_dff_A_zbMvYBGP4_1),.din(w_dff_A_hHCAGVJo6_1),.clk(gclk));
	jdff dff_A_CTbhVQDo6_1(.dout(w_dff_A_hHCAGVJo6_1),.din(w_dff_A_CTbhVQDo6_1),.clk(gclk));
	jdff dff_A_9ObARDXq4_1(.dout(w_dff_A_CTbhVQDo6_1),.din(w_dff_A_9ObARDXq4_1),.clk(gclk));
	jdff dff_A_zJIgK1Bg2_1(.dout(w_dff_A_9ObARDXq4_1),.din(w_dff_A_zJIgK1Bg2_1),.clk(gclk));
	jdff dff_A_zqrSmoA51_1(.dout(w_dff_A_zJIgK1Bg2_1),.din(w_dff_A_zqrSmoA51_1),.clk(gclk));
	jdff dff_A_DedMGlCN7_1(.dout(w_n328_0[1]),.din(w_dff_A_DedMGlCN7_1),.clk(gclk));
	jdff dff_A_y6plcCYG4_1(.dout(w_dff_A_DedMGlCN7_1),.din(w_dff_A_y6plcCYG4_1),.clk(gclk));
	jdff dff_A_MkH3xeQL1_1(.dout(w_dff_A_y6plcCYG4_1),.din(w_dff_A_MkH3xeQL1_1),.clk(gclk));
	jdff dff_A_r0cTBsIR1_1(.dout(w_dff_A_MkH3xeQL1_1),.din(w_dff_A_r0cTBsIR1_1),.clk(gclk));
	jdff dff_A_IuZ5LARV5_1(.dout(w_dff_A_r0cTBsIR1_1),.din(w_dff_A_IuZ5LARV5_1),.clk(gclk));
	jdff dff_A_6HCHyGQQ9_1(.dout(w_dff_A_IuZ5LARV5_1),.din(w_dff_A_6HCHyGQQ9_1),.clk(gclk));
	jdff dff_A_TSZsjlpV1_1(.dout(w_dff_A_6HCHyGQQ9_1),.din(w_dff_A_TSZsjlpV1_1),.clk(gclk));
	jdff dff_A_DlXKxutM3_1(.dout(w_dff_A_TSZsjlpV1_1),.din(w_dff_A_DlXKxutM3_1),.clk(gclk));
	jdff dff_A_fQNP7HS99_1(.dout(w_dff_A_DlXKxutM3_1),.din(w_dff_A_fQNP7HS99_1),.clk(gclk));
	jdff dff_A_bD5zvcQ85_0(.dout(w_G171gat_1[0]),.din(w_dff_A_bD5zvcQ85_0),.clk(gclk));
	jdff dff_A_HYozMjNj5_0(.dout(w_dff_A_bD5zvcQ85_0),.din(w_dff_A_HYozMjNj5_0),.clk(gclk));
	jdff dff_A_o90QN0yh6_0(.dout(w_dff_A_HYozMjNj5_0),.din(w_dff_A_o90QN0yh6_0),.clk(gclk));
	jdff dff_A_ePc1xQin2_0(.dout(w_dff_A_o90QN0yh6_0),.din(w_dff_A_ePc1xQin2_0),.clk(gclk));
	jdff dff_A_7UQSFdWA5_0(.dout(w_dff_A_ePc1xQin2_0),.din(w_dff_A_7UQSFdWA5_0),.clk(gclk));
	jdff dff_A_YmakPBz43_0(.dout(w_dff_A_7UQSFdWA5_0),.din(w_dff_A_YmakPBz43_0),.clk(gclk));
	jdff dff_A_uSBCJs0L2_1(.dout(w_G171gat_1[1]),.din(w_dff_A_uSBCJs0L2_1),.clk(gclk));
	jdff dff_A_CJVIKroK9_1(.dout(w_dff_A_uSBCJs0L2_1),.din(w_dff_A_CJVIKroK9_1),.clk(gclk));
	jdff dff_A_jiVdyjUa6_1(.dout(w_dff_A_CJVIKroK9_1),.din(w_dff_A_jiVdyjUa6_1),.clk(gclk));
	jdff dff_A_dfbKhmrs3_1(.dout(w_dff_A_jiVdyjUa6_1),.din(w_dff_A_dfbKhmrs3_1),.clk(gclk));
	jdff dff_A_B16m9Pz97_1(.dout(w_dff_A_dfbKhmrs3_1),.din(w_dff_A_B16m9Pz97_1),.clk(gclk));
	jdff dff_A_xrAKoSCS0_1(.dout(w_dff_A_B16m9Pz97_1),.din(w_dff_A_xrAKoSCS0_1),.clk(gclk));
	jdff dff_B_vZpFLVwD0_0(.din(n408),.dout(w_dff_B_vZpFLVwD0_0),.clk(gclk));
	jdff dff_B_DrDOqf6g9_0(.din(n406),.dout(w_dff_B_DrDOqf6g9_0),.clk(gclk));
	jdff dff_B_ZLQlakEG2_0(.din(w_dff_B_DrDOqf6g9_0),.dout(w_dff_B_ZLQlakEG2_0),.clk(gclk));
	jdff dff_B_C0eZyB142_0(.din(w_dff_B_ZLQlakEG2_0),.dout(w_dff_B_C0eZyB142_0),.clk(gclk));
	jdff dff_B_JjyBe0Tl7_0(.din(w_dff_B_C0eZyB142_0),.dout(w_dff_B_JjyBe0Tl7_0),.clk(gclk));
	jdff dff_B_Rhue5dRa1_0(.din(w_dff_B_JjyBe0Tl7_0),.dout(w_dff_B_Rhue5dRa1_0),.clk(gclk));
	jdff dff_B_i3zowgiz9_0(.din(w_dff_B_Rhue5dRa1_0),.dout(w_dff_B_i3zowgiz9_0),.clk(gclk));
	jdff dff_B_AXPtbETS2_0(.din(w_dff_B_i3zowgiz9_0),.dout(w_dff_B_AXPtbETS2_0),.clk(gclk));
	jdff dff_A_0IQAcb3k1_1(.dout(w_G91gat_0[1]),.din(w_dff_A_0IQAcb3k1_1),.clk(gclk));
	jdff dff_A_SmWtqAwe8_1(.dout(w_dff_A_0IQAcb3k1_1),.din(w_dff_A_SmWtqAwe8_1),.clk(gclk));
	jdff dff_A_s16vtcMS6_1(.dout(w_dff_A_SmWtqAwe8_1),.din(w_dff_A_s16vtcMS6_1),.clk(gclk));
	jdff dff_A_uiFXOIqy7_1(.dout(w_dff_A_s16vtcMS6_1),.din(w_dff_A_uiFXOIqy7_1),.clk(gclk));
	jdff dff_A_tVvGk56O2_1(.dout(w_dff_A_uiFXOIqy7_1),.din(w_dff_A_tVvGk56O2_1),.clk(gclk));
	jdff dff_A_ehnFyZms5_1(.dout(w_n404_0[1]),.din(w_dff_A_ehnFyZms5_1),.clk(gclk));
	jdff dff_A_2H2vucLm3_1(.dout(w_dff_A_ehnFyZms5_1),.din(w_dff_A_2H2vucLm3_1),.clk(gclk));
	jdff dff_A_esZKSQfr0_1(.dout(w_dff_A_2H2vucLm3_1),.din(w_dff_A_esZKSQfr0_1),.clk(gclk));
	jdff dff_A_n2wj0pkY2_1(.dout(w_dff_A_esZKSQfr0_1),.din(w_dff_A_n2wj0pkY2_1),.clk(gclk));
	jdff dff_A_fKX7qDbX4_1(.dout(w_dff_A_n2wj0pkY2_1),.din(w_dff_A_fKX7qDbX4_1),.clk(gclk));
	jdff dff_A_AXBQXbDI0_1(.dout(w_dff_A_fKX7qDbX4_1),.din(w_dff_A_AXBQXbDI0_1),.clk(gclk));
	jdff dff_A_MKvadVPG1_1(.dout(w_dff_A_AXBQXbDI0_1),.din(w_dff_A_MKvadVPG1_1),.clk(gclk));
	jdff dff_A_SOubNi2I9_1(.dout(w_dff_A_MKvadVPG1_1),.din(w_dff_A_SOubNi2I9_1),.clk(gclk));
	jdff dff_A_QBszpqbZ2_1(.dout(w_dff_A_SOubNi2I9_1),.din(w_dff_A_QBszpqbZ2_1),.clk(gclk));
	jdff dff_B_zVjBrFHL1_0(.din(n317),.dout(w_dff_B_zVjBrFHL1_0),.clk(gclk));
	jdff dff_B_og1wBcb82_0(.din(n316),.dout(w_dff_B_og1wBcb82_0),.clk(gclk));
	jdff dff_B_ydvYg7mL0_0(.din(w_dff_B_og1wBcb82_0),.dout(w_dff_B_ydvYg7mL0_0),.clk(gclk));
	jdff dff_B_bQDqAH6q8_0(.din(w_dff_B_ydvYg7mL0_0),.dout(w_dff_B_bQDqAH6q8_0),.clk(gclk));
	jdff dff_B_9JrxwEvH3_0(.din(w_dff_B_bQDqAH6q8_0),.dout(w_dff_B_9JrxwEvH3_0),.clk(gclk));
	jdff dff_A_J3nc7o1c4_1(.dout(w_G165gat_0[1]),.din(w_dff_A_J3nc7o1c4_1),.clk(gclk));
	jdff dff_A_Qe7FKe0u8_1(.dout(w_dff_A_J3nc7o1c4_1),.din(w_dff_A_Qe7FKe0u8_1),.clk(gclk));
	jdff dff_A_cOvZmYvq4_1(.dout(w_dff_A_Qe7FKe0u8_1),.din(w_dff_A_cOvZmYvq4_1),.clk(gclk));
	jdff dff_A_ovxeSliI1_1(.dout(w_dff_A_cOvZmYvq4_1),.din(w_dff_A_ovxeSliI1_1),.clk(gclk));
	jdff dff_A_Tm74dXJS5_1(.dout(w_dff_A_ovxeSliI1_1),.din(w_dff_A_Tm74dXJS5_1),.clk(gclk));
	jdff dff_A_IqRzScHt9_2(.dout(w_G165gat_0[2]),.din(w_dff_A_IqRzScHt9_2),.clk(gclk));
	jdff dff_A_cUN7fqHM0_2(.dout(w_dff_A_IqRzScHt9_2),.din(w_dff_A_cUN7fqHM0_2),.clk(gclk));
	jdff dff_A_9DkCoM124_2(.dout(w_dff_A_cUN7fqHM0_2),.din(w_dff_A_9DkCoM124_2),.clk(gclk));
	jdff dff_A_eCraVxkm0_2(.dout(w_dff_A_9DkCoM124_2),.din(w_dff_A_eCraVxkm0_2),.clk(gclk));
	jdff dff_A_Vt9q6fv93_2(.dout(w_dff_A_eCraVxkm0_2),.din(w_dff_A_Vt9q6fv93_2),.clk(gclk));
	jdff dff_A_yqRDbJJ93_2(.dout(w_dff_A_Vt9q6fv93_2),.din(w_dff_A_yqRDbJJ93_2),.clk(gclk));
	jdff dff_B_jhSL01uD2_3(.din(G165gat),.dout(w_dff_B_jhSL01uD2_3),.clk(gclk));
	jdff dff_B_KJXC6WmS8_1(.din(n426),.dout(w_dff_B_KJXC6WmS8_1),.clk(gclk));
	jdff dff_B_dOaZpg373_1(.din(w_dff_B_KJXC6WmS8_1),.dout(w_dff_B_dOaZpg373_1),.clk(gclk));
	jdff dff_B_TlNcn5Pv4_1(.din(w_dff_B_dOaZpg373_1),.dout(w_dff_B_TlNcn5Pv4_1),.clk(gclk));
	jdff dff_B_uJlR2KdT4_1(.din(w_dff_B_TlNcn5Pv4_1),.dout(w_dff_B_uJlR2KdT4_1),.clk(gclk));
	jdff dff_B_aeYg415G4_1(.din(w_dff_B_uJlR2KdT4_1),.dout(w_dff_B_aeYg415G4_1),.clk(gclk));
	jdff dff_B_sMyLpKxq2_1(.din(w_dff_B_aeYg415G4_1),.dout(w_dff_B_sMyLpKxq2_1),.clk(gclk));
	jdff dff_B_3eVLZlkj4_1(.din(w_dff_B_sMyLpKxq2_1),.dout(w_dff_B_3eVLZlkj4_1),.clk(gclk));
	jdff dff_B_YSwBDnKS8_1(.din(w_dff_B_3eVLZlkj4_1),.dout(w_dff_B_YSwBDnKS8_1),.clk(gclk));
	jdff dff_B_Jmt0lTr00_1(.din(w_dff_B_YSwBDnKS8_1),.dout(w_dff_B_Jmt0lTr00_1),.clk(gclk));
	jdff dff_B_6FS7ywOQ1_1(.din(n428),.dout(w_dff_B_6FS7ywOQ1_1),.clk(gclk));
	jdff dff_B_aKQvAoRF6_1(.din(w_dff_B_6FS7ywOQ1_1),.dout(w_dff_B_aKQvAoRF6_1),.clk(gclk));
	jdff dff_B_74NRWyks0_1(.din(w_dff_B_aKQvAoRF6_1),.dout(w_dff_B_74NRWyks0_1),.clk(gclk));
	jdff dff_B_xuosGLmR3_1(.din(n340),.dout(w_dff_B_xuosGLmR3_1),.clk(gclk));
	jdff dff_B_SZO2vpfW5_1(.din(w_dff_B_xuosGLmR3_1),.dout(w_dff_B_SZO2vpfW5_1),.clk(gclk));
	jdff dff_B_vctFiGWx8_1(.din(w_dff_B_SZO2vpfW5_1),.dout(w_dff_B_vctFiGWx8_1),.clk(gclk));
	jdff dff_B_oWJGObSn8_1(.din(w_dff_B_vctFiGWx8_1),.dout(w_dff_B_oWJGObSn8_1),.clk(gclk));
	jdff dff_B_fnNvb5kg5_1(.din(w_dff_B_oWJGObSn8_1),.dout(w_dff_B_fnNvb5kg5_1),.clk(gclk));
	jdff dff_B_XXM4xDtG9_1(.din(n344),.dout(w_dff_B_XXM4xDtG9_1),.clk(gclk));
	jdff dff_B_NxF3yOF08_1(.din(w_dff_B_XXM4xDtG9_1),.dout(w_dff_B_NxF3yOF08_1),.clk(gclk));
	jdff dff_B_eyRduMUH2_1(.din(w_dff_B_NxF3yOF08_1),.dout(w_dff_B_eyRduMUH2_1),.clk(gclk));
	jdff dff_B_CFs5Y1xx7_1(.din(w_dff_B_eyRduMUH2_1),.dout(w_dff_B_CFs5Y1xx7_1),.clk(gclk));
	jdff dff_B_yMHv5IkB9_0(.din(n244),.dout(w_dff_B_yMHv5IkB9_0),.clk(gclk));
	jdff dff_B_zXYD6iSI0_0(.din(w_dff_B_yMHv5IkB9_0),.dout(w_dff_B_zXYD6iSI0_0),.clk(gclk));
	jdff dff_B_DWlw1QNO9_0(.din(w_dff_B_zXYD6iSI0_0),.dout(w_dff_B_DWlw1QNO9_0),.clk(gclk));
	jdff dff_B_S3sYJPcS1_0(.din(n171),.dout(w_dff_B_S3sYJPcS1_0),.clk(gclk));
	jdff dff_A_Wf2H0hlY2_0(.dout(w_G219gat_1[0]),.din(w_dff_A_Wf2H0hlY2_0),.clk(gclk));
	jdff dff_A_ZjTjFceJ6_2(.dout(w_G219gat_1[2]),.din(w_dff_A_ZjTjFceJ6_2),.clk(gclk));
	jdff dff_A_IAiiqf3i6_0(.dout(w_G219gat_0[0]),.din(w_dff_A_IAiiqf3i6_0),.clk(gclk));
	jdff dff_A_o97X8kgB7_0(.dout(w_dff_A_IAiiqf3i6_0),.din(w_dff_A_o97X8kgB7_0),.clk(gclk));
	jdff dff_A_Kbnq7u2O1_0(.dout(w_dff_A_o97X8kgB7_0),.din(w_dff_A_Kbnq7u2O1_0),.clk(gclk));
	jdff dff_A_Z46QNUuo2_0(.dout(w_dff_A_Kbnq7u2O1_0),.din(w_dff_A_Z46QNUuo2_0),.clk(gclk));
	jdff dff_A_zS1JG0L90_0(.dout(w_dff_A_Z46QNUuo2_0),.din(w_dff_A_zS1JG0L90_0),.clk(gclk));
	jdff dff_A_trNkA0at5_2(.dout(w_G219gat_0[2]),.din(w_dff_A_trNkA0at5_2),.clk(gclk));
	jdff dff_B_NFJP6KVg8_3(.din(G219gat),.dout(w_dff_B_NFJP6KVg8_3),.clk(gclk));
	jdff dff_B_zjjYFn9h6_3(.din(w_dff_B_NFJP6KVg8_3),.dout(w_dff_B_zjjYFn9h6_3),.clk(gclk));
	jdff dff_B_8A0IAFZs3_3(.din(w_dff_B_zjjYFn9h6_3),.dout(w_dff_B_8A0IAFZs3_3),.clk(gclk));
	jdff dff_B_TzjtyDDp6_3(.din(w_dff_B_8A0IAFZs3_3),.dout(w_dff_B_TzjtyDDp6_3),.clk(gclk));
	jdff dff_B_17y8TwHh1_3(.din(w_dff_B_TzjtyDDp6_3),.dout(w_dff_B_17y8TwHh1_3),.clk(gclk));
	jdff dff_B_1nGfh1w22_3(.din(w_dff_B_17y8TwHh1_3),.dout(w_dff_B_1nGfh1w22_3),.clk(gclk));
	jdff dff_B_qusmwgnb2_3(.din(w_dff_B_1nGfh1w22_3),.dout(w_dff_B_qusmwgnb2_3),.clk(gclk));
	jdff dff_B_lh7zMWQ93_3(.din(w_dff_B_qusmwgnb2_3),.dout(w_dff_B_lh7zMWQ93_3),.clk(gclk));
	jdff dff_B_wDGhJLLo9_3(.din(w_dff_B_lh7zMWQ93_3),.dout(w_dff_B_wDGhJLLo9_3),.clk(gclk));
	jdff dff_B_SWnVk3fM4_0(.din(n427),.dout(w_dff_B_SWnVk3fM4_0),.clk(gclk));
	jdff dff_B_faK5CgCR4_0(.din(w_dff_B_SWnVk3fM4_0),.dout(w_dff_B_faK5CgCR4_0),.clk(gclk));
	jdff dff_B_OpAQCHQY5_0(.din(w_dff_B_faK5CgCR4_0),.dout(w_dff_B_OpAQCHQY5_0),.clk(gclk));
	jdff dff_B_mVVOJtFA1_0(.din(w_dff_B_OpAQCHQY5_0),.dout(w_dff_B_mVVOJtFA1_0),.clk(gclk));
	jdff dff_B_mYze1cyB0_0(.din(w_dff_B_mVVOJtFA1_0),.dout(w_dff_B_mYze1cyB0_0),.clk(gclk));
	jdff dff_B_HgvTrgrE4_1(.din(n389),.dout(w_dff_B_HgvTrgrE4_1),.clk(gclk));
	jdff dff_B_9LoH4KPU1_1(.din(w_dff_B_HgvTrgrE4_1),.dout(w_dff_B_9LoH4KPU1_1),.clk(gclk));
	jdff dff_B_aTDe0dh08_1(.din(w_dff_B_9LoH4KPU1_1),.dout(w_dff_B_aTDe0dh08_1),.clk(gclk));
	jdff dff_B_CfTfS9m79_1(.din(w_dff_B_aTDe0dh08_1),.dout(w_dff_B_CfTfS9m79_1),.clk(gclk));
	jdff dff_B_odkAes6T3_1(.din(n359),.dout(w_dff_B_odkAes6T3_1),.clk(gclk));
	jdff dff_B_fFMHPjKW7_1(.din(w_dff_B_odkAes6T3_1),.dout(w_dff_B_fFMHPjKW7_1),.clk(gclk));
	jdff dff_B_iQF2qdDc8_1(.din(w_dff_B_fFMHPjKW7_1),.dout(w_dff_B_iQF2qdDc8_1),.clk(gclk));
	jdff dff_B_iAbdEwOF6_1(.din(n252),.dout(w_dff_B_iAbdEwOF6_1),.clk(gclk));
	jdff dff_B_174OM27a1_1(.din(w_dff_B_iAbdEwOF6_1),.dout(w_dff_B_174OM27a1_1),.clk(gclk));
	jdff dff_B_vhh45I5e9_1(.din(n253),.dout(w_dff_B_vhh45I5e9_1),.clk(gclk));
	jdff dff_B_TOWDjmT62_1(.din(w_dff_B_vhh45I5e9_1),.dout(w_dff_B_TOWDjmT62_1),.clk(gclk));
	jdff dff_B_qbt2vy6h2_1(.din(w_dff_B_TOWDjmT62_1),.dout(w_dff_B_qbt2vy6h2_1),.clk(gclk));
	jdff dff_B_mlaOqiYt2_1(.din(n254),.dout(w_dff_B_mlaOqiYt2_1),.clk(gclk));
	jdff dff_B_AEHREUcU6_1(.din(n255),.dout(w_dff_B_AEHREUcU6_1),.clk(gclk));
	jdff dff_B_KHqf8zhh8_1(.din(w_dff_B_AEHREUcU6_1),.dout(w_dff_B_KHqf8zhh8_1),.clk(gclk));
	jdff dff_A_dXaXVj1q0_1(.dout(w_n209_0[1]),.din(w_dff_A_dXaXVj1q0_1),.clk(gclk));
	jdff dff_A_ksjfY7GK7_1(.dout(w_dff_A_dXaXVj1q0_1),.din(w_dff_A_ksjfY7GK7_1),.clk(gclk));
	jdff dff_B_XdtsCMJR9_2(.din(n209),.dout(w_dff_B_XdtsCMJR9_2),.clk(gclk));
	jdff dff_B_SiCG6sbq2_2(.din(w_dff_B_XdtsCMJR9_2),.dout(w_dff_B_SiCG6sbq2_2),.clk(gclk));
	jdff dff_B_v0KGXehj0_2(.din(w_dff_B_SiCG6sbq2_2),.dout(w_dff_B_v0KGXehj0_2),.clk(gclk));
	jdff dff_B_JyUnwTMj7_2(.din(w_dff_B_v0KGXehj0_2),.dout(w_dff_B_JyUnwTMj7_2),.clk(gclk));
	jdff dff_B_8CLSBiVb8_2(.din(w_dff_B_JyUnwTMj7_2),.dout(w_dff_B_8CLSBiVb8_2),.clk(gclk));
	jdff dff_B_4SBoA1ic7_2(.din(w_dff_B_8CLSBiVb8_2),.dout(w_dff_B_4SBoA1ic7_2),.clk(gclk));
	jdff dff_B_tgNJEoev1_2(.din(w_dff_B_4SBoA1ic7_2),.dout(w_dff_B_tgNJEoev1_2),.clk(gclk));
	jdff dff_A_1IBYGsO18_0(.dout(w_G261gat_0[0]),.din(w_dff_A_1IBYGsO18_0),.clk(gclk));
	jdff dff_A_D4woEsY74_0(.dout(w_dff_A_1IBYGsO18_0),.din(w_dff_A_D4woEsY74_0),.clk(gclk));
	jdff dff_A_jB1P23PB0_0(.dout(w_dff_A_D4woEsY74_0),.din(w_dff_A_jB1P23PB0_0),.clk(gclk));
	jdff dff_A_SiiAtopi7_0(.dout(w_dff_A_jB1P23PB0_0),.din(w_dff_A_SiiAtopi7_0),.clk(gclk));
	jdff dff_A_gWlp2XUR5_0(.dout(w_dff_A_SiiAtopi7_0),.din(w_dff_A_gWlp2XUR5_0),.clk(gclk));
	jdff dff_A_CHDEXkLs0_0(.dout(w_dff_A_gWlp2XUR5_0),.din(w_dff_A_CHDEXkLs0_0),.clk(gclk));
	jdff dff_A_7wpFEAVr2_0(.dout(w_dff_A_CHDEXkLs0_0),.din(w_dff_A_7wpFEAVr2_0),.clk(gclk));
	jdff dff_A_6gRVB6vU5_2(.dout(w_G261gat_0[2]),.din(w_dff_A_6gRVB6vU5_2),.clk(gclk));
	jdff dff_A_oD1PAPfr0_2(.dout(w_dff_A_6gRVB6vU5_2),.din(w_dff_A_oD1PAPfr0_2),.clk(gclk));
	jdff dff_A_nnfEkIhN5_2(.dout(w_dff_A_oD1PAPfr0_2),.din(w_dff_A_nnfEkIhN5_2),.clk(gclk));
	jdff dff_A_UkosGhHV9_2(.dout(w_dff_A_nnfEkIhN5_2),.din(w_dff_A_UkosGhHV9_2),.clk(gclk));
	jdff dff_A_kLSexX1o4_2(.dout(w_dff_A_UkosGhHV9_2),.din(w_dff_A_kLSexX1o4_2),.clk(gclk));
	jdff dff_A_sL0toZFT4_2(.dout(w_dff_A_kLSexX1o4_2),.din(w_dff_A_sL0toZFT4_2),.clk(gclk));
	jdff dff_A_nqQkIykf5_2(.dout(w_dff_A_sL0toZFT4_2),.din(w_dff_A_nqQkIykf5_2),.clk(gclk));
	jdff dff_A_alRdQcG84_2(.dout(w_dff_A_nqQkIykf5_2),.din(w_dff_A_alRdQcG84_2),.clk(gclk));
	jdff dff_A_Xvcckb5q5_2(.dout(w_dff_A_alRdQcG84_2),.din(w_dff_A_Xvcckb5q5_2),.clk(gclk));
	jdff dff_B_EEo6iHmn8_0(.din(n196),.dout(w_dff_B_EEo6iHmn8_0),.clk(gclk));
	jdff dff_B_QHzuWFgV4_0(.din(w_dff_B_EEo6iHmn8_0),.dout(w_dff_B_QHzuWFgV4_0),.clk(gclk));
	jdff dff_B_yWnPKxVu2_0(.din(w_dff_B_QHzuWFgV4_0),.dout(w_dff_B_yWnPKxVu2_0),.clk(gclk));
	jdff dff_B_8rvGSJTv5_0(.din(n195),.dout(w_dff_B_8rvGSJTv5_0),.clk(gclk));
	jdff dff_B_LXHGXDS25_1(.din(n191),.dout(w_dff_B_LXHGXDS25_1),.clk(gclk));
	jdff dff_B_rjEnrd192_1(.din(n183),.dout(w_dff_B_rjEnrd192_1),.clk(gclk));
	jdff dff_B_VNrkrfuU0_1(.din(w_dff_B_rjEnrd192_1),.dout(w_dff_B_VNrkrfuU0_1),.clk(gclk));
	jdff dff_B_yzra5jcw6_0(.din(n187),.dout(w_dff_B_yzra5jcw6_0),.clk(gclk));
	jdff dff_A_UBalm7Lv3_1(.dout(w_G126gat_0[1]),.din(w_dff_A_UBalm7Lv3_1),.clk(gclk));
	jdff dff_A_pD37gmHI4_1(.dout(w_dff_A_UBalm7Lv3_1),.din(w_dff_A_pD37gmHI4_1),.clk(gclk));
	jdff dff_A_RBhIt13U0_1(.dout(w_dff_A_pD37gmHI4_1),.din(w_dff_A_RBhIt13U0_1),.clk(gclk));
	jdff dff_A_sOLrYTH73_1(.dout(w_dff_A_RBhIt13U0_1),.din(w_dff_A_sOLrYTH73_1),.clk(gclk));
	jdff dff_A_zkfDkXYw9_1(.dout(w_dff_A_sOLrYTH73_1),.din(w_dff_A_zkfDkXYw9_1),.clk(gclk));
	jdff dff_B_06ecEtg02_3(.din(n181),.dout(w_dff_B_06ecEtg02_3),.clk(gclk));
	jdff dff_B_oq7NxDPX3_3(.din(w_dff_B_06ecEtg02_3),.dout(w_dff_B_oq7NxDPX3_3),.clk(gclk));
	jdff dff_B_UEkLvT6m8_3(.din(w_dff_B_oq7NxDPX3_3),.dout(w_dff_B_UEkLvT6m8_3),.clk(gclk));
	jdff dff_B_yFgtCBhi9_3(.din(w_dff_B_UEkLvT6m8_3),.dout(w_dff_B_yFgtCBhi9_3),.clk(gclk));
	jdff dff_B_z5Smd1ad6_3(.din(w_dff_B_yFgtCBhi9_3),.dout(w_dff_B_z5Smd1ad6_3),.clk(gclk));
	jdff dff_B_rmc1moKw7_3(.din(w_dff_B_z5Smd1ad6_3),.dout(w_dff_B_rmc1moKw7_3),.clk(gclk));
	jdff dff_B_aeLYM4i55_3(.din(w_dff_B_rmc1moKw7_3),.dout(w_dff_B_aeLYM4i55_3),.clk(gclk));
	jdff dff_A_suOJKDa05_1(.dout(w_G201gat_0[1]),.din(w_dff_A_suOJKDa05_1),.clk(gclk));
	jdff dff_A_YZ83nlWG2_1(.dout(w_dff_A_suOJKDa05_1),.din(w_dff_A_YZ83nlWG2_1),.clk(gclk));
	jdff dff_A_IPvx8p3y3_1(.dout(w_dff_A_YZ83nlWG2_1),.din(w_dff_A_IPvx8p3y3_1),.clk(gclk));
	jdff dff_A_b2awXjOu8_1(.dout(w_dff_A_IPvx8p3y3_1),.din(w_dff_A_b2awXjOu8_1),.clk(gclk));
	jdff dff_A_H8RsPoNV2_1(.dout(w_dff_A_b2awXjOu8_1),.din(w_dff_A_H8RsPoNV2_1),.clk(gclk));
	jdff dff_A_wB7S1cRe7_1(.dout(w_dff_A_H8RsPoNV2_1),.din(w_dff_A_wB7S1cRe7_1),.clk(gclk));
	jdff dff_A_ULAE3HpL3_1(.dout(w_n241_0[1]),.din(w_dff_A_ULAE3HpL3_1),.clk(gclk));
	jdff dff_A_DpahGmAm1_1(.dout(w_dff_A_ULAE3HpL3_1),.din(w_dff_A_DpahGmAm1_1),.clk(gclk));
	jdff dff_A_d11fSYTr4_1(.dout(w_dff_A_DpahGmAm1_1),.din(w_dff_A_d11fSYTr4_1),.clk(gclk));
	jdff dff_A_ESlTA6IA9_1(.dout(w_dff_A_d11fSYTr4_1),.din(w_dff_A_ESlTA6IA9_1),.clk(gclk));
	jdff dff_A_OPWn0AdZ8_1(.dout(w_dff_A_ESlTA6IA9_1),.din(w_dff_A_OPWn0AdZ8_1),.clk(gclk));
	jdff dff_A_YSF8Dwbr8_1(.dout(w_G195gat_1[1]),.din(w_dff_A_YSF8Dwbr8_1),.clk(gclk));
	jdff dff_A_q5LsXBCT6_1(.dout(w_dff_A_YSF8Dwbr8_1),.din(w_dff_A_q5LsXBCT6_1),.clk(gclk));
	jdff dff_A_Zl6fLIM01_1(.dout(w_dff_A_q5LsXBCT6_1),.din(w_dff_A_Zl6fLIM01_1),.clk(gclk));
	jdff dff_A_5I7d8ltg5_1(.dout(w_dff_A_Zl6fLIM01_1),.din(w_dff_A_5I7d8ltg5_1),.clk(gclk));
	jdff dff_A_uvNG0BQX1_1(.dout(w_dff_A_5I7d8ltg5_1),.din(w_dff_A_uvNG0BQX1_1),.clk(gclk));
	jdff dff_A_U1w57x487_1(.dout(w_dff_A_uvNG0BQX1_1),.din(w_dff_A_U1w57x487_1),.clk(gclk));
	jdff dff_A_nEtWniCD5_2(.dout(w_G195gat_1[2]),.din(w_dff_A_nEtWniCD5_2),.clk(gclk));
	jdff dff_A_PZTH6ZlS0_2(.dout(w_dff_A_nEtWniCD5_2),.din(w_dff_A_PZTH6ZlS0_2),.clk(gclk));
	jdff dff_A_w7mMJzuS1_2(.dout(w_dff_A_PZTH6ZlS0_2),.din(w_dff_A_w7mMJzuS1_2),.clk(gclk));
	jdff dff_A_myQyaN844_2(.dout(w_dff_A_w7mMJzuS1_2),.din(w_dff_A_myQyaN844_2),.clk(gclk));
	jdff dff_A_oyiRnW668_2(.dout(w_dff_A_myQyaN844_2),.din(w_dff_A_oyiRnW668_2),.clk(gclk));
	jdff dff_A_SYPybmbJ0_2(.dout(w_dff_A_oyiRnW668_2),.din(w_dff_A_SYPybmbJ0_2),.clk(gclk));
	jdff dff_A_OQsddf6b0_1(.dout(w_n240_0[1]),.din(w_dff_A_OQsddf6b0_1),.clk(gclk));
	jdff dff_A_EQ06nY0c5_1(.dout(w_dff_A_OQsddf6b0_1),.din(w_dff_A_EQ06nY0c5_1),.clk(gclk));
	jdff dff_A_BONjA3LD0_1(.dout(w_dff_A_EQ06nY0c5_1),.din(w_dff_A_BONjA3LD0_1),.clk(gclk));
	jdff dff_A_JeGlmZaJ4_1(.dout(w_dff_A_BONjA3LD0_1),.din(w_dff_A_JeGlmZaJ4_1),.clk(gclk));
	jdff dff_A_gblR4WM46_1(.dout(w_dff_A_JeGlmZaJ4_1),.din(w_dff_A_gblR4WM46_1),.clk(gclk));
	jdff dff_B_GZeGIeJg7_0(.din(n237),.dout(w_dff_B_GZeGIeJg7_0),.clk(gclk));
	jdff dff_A_dCB7B7Mt5_0(.dout(w_G121gat_0[0]),.din(w_dff_A_dCB7B7Mt5_0),.clk(gclk));
	jdff dff_A_p8ekeHrl2_0(.dout(w_dff_A_dCB7B7Mt5_0),.din(w_dff_A_p8ekeHrl2_0),.clk(gclk));
	jdff dff_A_jyotcOTw4_0(.dout(w_dff_A_p8ekeHrl2_0),.din(w_dff_A_jyotcOTw4_0),.clk(gclk));
	jdff dff_A_XwizvcJe4_0(.dout(w_dff_A_jyotcOTw4_0),.din(w_dff_A_XwizvcJe4_0),.clk(gclk));
	jdff dff_A_KyQsSQ0E2_0(.dout(w_dff_A_XwizvcJe4_0),.din(w_dff_A_KyQsSQ0E2_0),.clk(gclk));
	jdff dff_A_r2rIaCPk6_0(.dout(w_G195gat_2[0]),.din(w_dff_A_r2rIaCPk6_0),.clk(gclk));
	jdff dff_A_8RPEXi2V4_0(.dout(w_dff_A_r2rIaCPk6_0),.din(w_dff_A_8RPEXi2V4_0),.clk(gclk));
	jdff dff_A_nWYoHk6q9_0(.dout(w_dff_A_8RPEXi2V4_0),.din(w_dff_A_nWYoHk6q9_0),.clk(gclk));
	jdff dff_A_CblQHe8Z2_0(.dout(w_dff_A_nWYoHk6q9_0),.din(w_dff_A_CblQHe8Z2_0),.clk(gclk));
	jdff dff_A_AugJmRfe2_0(.dout(w_dff_A_CblQHe8Z2_0),.din(w_dff_A_AugJmRfe2_0),.clk(gclk));
	jdff dff_A_nYxAQpCt9_0(.dout(w_dff_A_AugJmRfe2_0),.din(w_dff_A_nYxAQpCt9_0),.clk(gclk));
	jdff dff_A_mph99VEh3_2(.dout(w_G195gat_0[2]),.din(w_dff_A_mph99VEh3_2),.clk(gclk));
	jdff dff_A_E2JqAQvl6_2(.dout(w_dff_A_mph99VEh3_2),.din(w_dff_A_E2JqAQvl6_2),.clk(gclk));
	jdff dff_A_v8QyBFIZ8_2(.dout(w_dff_A_E2JqAQvl6_2),.din(w_dff_A_v8QyBFIZ8_2),.clk(gclk));
	jdff dff_A_hB4lQznq7_2(.dout(w_dff_A_v8QyBFIZ8_2),.din(w_dff_A_hB4lQznq7_2),.clk(gclk));
	jdff dff_A_nWno1Wal2_1(.dout(w_n235_0[1]),.din(w_dff_A_nWno1Wal2_1),.clk(gclk));
	jdff dff_A_re5dLjmD7_1(.dout(w_dff_A_nWno1Wal2_1),.din(w_dff_A_re5dLjmD7_1),.clk(gclk));
	jdff dff_A_sgBEVCZO9_1(.dout(w_dff_A_re5dLjmD7_1),.din(w_dff_A_sgBEVCZO9_1),.clk(gclk));
	jdff dff_A_fT2zX8mp0_1(.dout(w_dff_A_sgBEVCZO9_1),.din(w_dff_A_fT2zX8mp0_1),.clk(gclk));
	jdff dff_A_Cd0ItszR6_1(.dout(w_dff_A_fT2zX8mp0_1),.din(w_dff_A_Cd0ItszR6_1),.clk(gclk));
	jdff dff_A_LqsTnaKk6_1(.dout(w_dff_A_Cd0ItszR6_1),.din(w_dff_A_LqsTnaKk6_1),.clk(gclk));
	jdff dff_A_FObxGTHh5_1(.dout(w_G189gat_1[1]),.din(w_dff_A_FObxGTHh5_1),.clk(gclk));
	jdff dff_A_ktS4YwME7_1(.dout(w_dff_A_FObxGTHh5_1),.din(w_dff_A_ktS4YwME7_1),.clk(gclk));
	jdff dff_A_8u6x1zgP9_1(.dout(w_dff_A_ktS4YwME7_1),.din(w_dff_A_8u6x1zgP9_1),.clk(gclk));
	jdff dff_A_Y14E0BAy5_1(.dout(w_dff_A_8u6x1zgP9_1),.din(w_dff_A_Y14E0BAy5_1),.clk(gclk));
	jdff dff_A_CP88kakA0_1(.dout(w_dff_A_Y14E0BAy5_1),.din(w_dff_A_CP88kakA0_1),.clk(gclk));
	jdff dff_A_3VLFMT3U3_1(.dout(w_dff_A_CP88kakA0_1),.din(w_dff_A_3VLFMT3U3_1),.clk(gclk));
	jdff dff_A_Nhp5KMZX9_2(.dout(w_G189gat_1[2]),.din(w_dff_A_Nhp5KMZX9_2),.clk(gclk));
	jdff dff_A_MFyv88hl6_2(.dout(w_dff_A_Nhp5KMZX9_2),.din(w_dff_A_MFyv88hl6_2),.clk(gclk));
	jdff dff_A_d5bGZOk15_2(.dout(w_dff_A_MFyv88hl6_2),.din(w_dff_A_d5bGZOk15_2),.clk(gclk));
	jdff dff_A_vtQCxj908_2(.dout(w_dff_A_d5bGZOk15_2),.din(w_dff_A_vtQCxj908_2),.clk(gclk));
	jdff dff_A_87qMAd0C7_2(.dout(w_dff_A_vtQCxj908_2),.din(w_dff_A_87qMAd0C7_2),.clk(gclk));
	jdff dff_A_8cuxrSrU0_2(.dout(w_dff_A_87qMAd0C7_2),.din(w_dff_A_8cuxrSrU0_2),.clk(gclk));
	jdff dff_A_bXXcMXfy8_1(.dout(w_n234_0[1]),.din(w_dff_A_bXXcMXfy8_1),.clk(gclk));
	jdff dff_A_0lAv7VJc6_1(.dout(w_dff_A_bXXcMXfy8_1),.din(w_dff_A_0lAv7VJc6_1),.clk(gclk));
	jdff dff_A_2XhZqoQH4_1(.dout(w_dff_A_0lAv7VJc6_1),.din(w_dff_A_2XhZqoQH4_1),.clk(gclk));
	jdff dff_A_2iJHIspx2_1(.dout(w_dff_A_2XhZqoQH4_1),.din(w_dff_A_2iJHIspx2_1),.clk(gclk));
	jdff dff_A_2agpt3LK1_1(.dout(w_dff_A_2iJHIspx2_1),.din(w_dff_A_2agpt3LK1_1),.clk(gclk));
	jdff dff_A_vVTloqkZ2_1(.dout(w_dff_A_2agpt3LK1_1),.din(w_dff_A_vVTloqkZ2_1),.clk(gclk));
	jdff dff_B_FqU1p9qq9_0(.din(n231),.dout(w_dff_B_FqU1p9qq9_0),.clk(gclk));
	jdff dff_B_0ilOWy2G4_2(.din(G146gat),.dout(w_dff_B_0ilOWy2G4_2),.clk(gclk));
	jdff dff_B_MRjS1Njp8_2(.din(w_dff_B_0ilOWy2G4_2),.dout(w_dff_B_MRjS1Njp8_2),.clk(gclk));
	jdff dff_B_gRcPpe5u6_2(.din(w_dff_B_MRjS1Njp8_2),.dout(w_dff_B_gRcPpe5u6_2),.clk(gclk));
	jdff dff_B_NSpcUwYz7_2(.din(w_dff_B_gRcPpe5u6_2),.dout(w_dff_B_NSpcUwYz7_2),.clk(gclk));
	jdff dff_A_oZmKzSsl3_1(.dout(w_G116gat_0[1]),.din(w_dff_A_oZmKzSsl3_1),.clk(gclk));
	jdff dff_A_97LCpHz03_1(.dout(w_dff_A_oZmKzSsl3_1),.din(w_dff_A_97LCpHz03_1),.clk(gclk));
	jdff dff_A_crK0N7Vs8_1(.dout(w_dff_A_97LCpHz03_1),.din(w_dff_A_crK0N7Vs8_1),.clk(gclk));
	jdff dff_A_c1N16EQg6_1(.dout(w_dff_A_crK0N7Vs8_1),.din(w_dff_A_c1N16EQg6_1),.clk(gclk));
	jdff dff_A_bWkaAc2M5_1(.dout(w_dff_A_c1N16EQg6_1),.din(w_dff_A_bWkaAc2M5_1),.clk(gclk));
	jdff dff_A_tXEFaYxt1_0(.dout(w_G189gat_2[0]),.din(w_dff_A_tXEFaYxt1_0),.clk(gclk));
	jdff dff_A_tS9FdZ5z7_0(.dout(w_dff_A_tXEFaYxt1_0),.din(w_dff_A_tS9FdZ5z7_0),.clk(gclk));
	jdff dff_A_CwYXyIC57_0(.dout(w_dff_A_tS9FdZ5z7_0),.din(w_dff_A_CwYXyIC57_0),.clk(gclk));
	jdff dff_A_UzEpeajt9_0(.dout(w_dff_A_CwYXyIC57_0),.din(w_dff_A_UzEpeajt9_0),.clk(gclk));
	jdff dff_A_IHAUkHO70_0(.dout(w_dff_A_UzEpeajt9_0),.din(w_dff_A_IHAUkHO70_0),.clk(gclk));
	jdff dff_A_otoplOJD7_0(.dout(w_dff_A_IHAUkHO70_0),.din(w_dff_A_otoplOJD7_0),.clk(gclk));
	jdff dff_A_GI8UFyGU1_2(.dout(w_G189gat_0[2]),.din(w_dff_A_GI8UFyGU1_2),.clk(gclk));
	jdff dff_A_zDQ4ax1z6_2(.dout(w_dff_A_GI8UFyGU1_2),.din(w_dff_A_zDQ4ax1z6_2),.clk(gclk));
	jdff dff_A_MX0Zr1Yw4_2(.dout(w_dff_A_zDQ4ax1z6_2),.din(w_dff_A_MX0Zr1Yw4_2),.clk(gclk));
	jdff dff_A_Lb4784C42_2(.dout(w_dff_A_MX0Zr1Yw4_2),.din(w_dff_A_Lb4784C42_2),.clk(gclk));
	jdff dff_A_PotDqNv55_0(.dout(w_n343_0[0]),.din(w_dff_A_PotDqNv55_0),.clk(gclk));
	jdff dff_A_vcxIwZ0Q9_0(.dout(w_dff_A_PotDqNv55_0),.din(w_dff_A_vcxIwZ0Q9_0),.clk(gclk));
	jdff dff_A_Uex1Sy8D9_0(.dout(w_dff_A_vcxIwZ0Q9_0),.din(w_dff_A_Uex1Sy8D9_0),.clk(gclk));
	jdff dff_B_BFM5aiq04_1(.din(n341),.dout(w_dff_B_BFM5aiq04_1),.clk(gclk));
	jdff dff_B_aPH4xSno0_1(.din(w_dff_B_BFM5aiq04_1),.dout(w_dff_B_aPH4xSno0_1),.clk(gclk));
	jdff dff_B_LHtW3sfA3_1(.din(w_dff_B_aPH4xSno0_1),.dout(w_dff_B_LHtW3sfA3_1),.clk(gclk));
	jdff dff_B_1Wcb2P884_1(.din(w_dff_B_LHtW3sfA3_1),.dout(w_dff_B_1Wcb2P884_1),.clk(gclk));
	jdff dff_B_eiKI6U6S8_1(.din(w_dff_B_1Wcb2P884_1),.dout(w_dff_B_eiKI6U6S8_1),.clk(gclk));
	jdff dff_B_HC1jVCeB8_1(.din(w_dff_B_eiKI6U6S8_1),.dout(w_dff_B_HC1jVCeB8_1),.clk(gclk));
	jdff dff_A_5cxBnz5X5_1(.dout(w_n222_0[1]),.din(w_dff_A_5cxBnz5X5_1),.clk(gclk));
	jdff dff_A_fLnI7T5g4_1(.dout(w_dff_A_5cxBnz5X5_1),.din(w_dff_A_fLnI7T5g4_1),.clk(gclk));
	jdff dff_A_VOjLmj5e3_1(.dout(w_dff_A_fLnI7T5g4_1),.din(w_dff_A_VOjLmj5e3_1),.clk(gclk));
	jdff dff_A_YOt3qKd65_1(.dout(w_dff_A_VOjLmj5e3_1),.din(w_dff_A_YOt3qKd65_1),.clk(gclk));
	jdff dff_A_qjpVXUau6_1(.dout(w_dff_A_YOt3qKd65_1),.din(w_dff_A_qjpVXUau6_1),.clk(gclk));
	jdff dff_A_BVH0VYLg1_1(.dout(w_dff_A_qjpVXUau6_1),.din(w_dff_A_BVH0VYLg1_1),.clk(gclk));
	jdff dff_A_gnhZkBHY0_1(.dout(w_dff_A_BVH0VYLg1_1),.din(w_dff_A_gnhZkBHY0_1),.clk(gclk));
	jdff dff_B_tExV6k4Y7_0(.din(n216),.dout(w_dff_B_tExV6k4Y7_0),.clk(gclk));
	jdff dff_A_zQVbo4Md0_0(.dout(w_n97_0[0]),.din(w_dff_A_zQVbo4Md0_0),.clk(gclk));
	jdff dff_A_KthTLXre9_0(.dout(w_dff_A_zQVbo4Md0_0),.din(w_dff_A_KthTLXre9_0),.clk(gclk));
	jdff dff_A_AwLQZzfH2_0(.dout(w_dff_A_KthTLXre9_0),.din(w_dff_A_AwLQZzfH2_0),.clk(gclk));
	jdff dff_B_YcLKcsg87_2(.din(G143gat),.dout(w_dff_B_YcLKcsg87_2),.clk(gclk));
	jdff dff_B_MT7eeJA04_2(.din(w_dff_B_YcLKcsg87_2),.dout(w_dff_B_MT7eeJA04_2),.clk(gclk));
	jdff dff_B_DgHKgcrT3_2(.din(w_dff_B_MT7eeJA04_2),.dout(w_dff_B_DgHKgcrT3_2),.clk(gclk));
	jdff dff_B_9ieTWPER3_2(.din(w_dff_B_DgHKgcrT3_2),.dout(w_dff_B_9ieTWPER3_2),.clk(gclk));
	jdff dff_A_YkoPwWJI0_1(.dout(w_G111gat_0[1]),.din(w_dff_A_YkoPwWJI0_1),.clk(gclk));
	jdff dff_A_QhNNhfQG7_1(.dout(w_dff_A_YkoPwWJI0_1),.din(w_dff_A_QhNNhfQG7_1),.clk(gclk));
	jdff dff_A_zYDUrmcf6_1(.dout(w_dff_A_QhNNhfQG7_1),.din(w_dff_A_zYDUrmcf6_1),.clk(gclk));
	jdff dff_A_H8oosr1I6_1(.dout(w_dff_A_zYDUrmcf6_1),.din(w_dff_A_H8oosr1I6_1),.clk(gclk));
	jdff dff_A_wbINvpvQ9_1(.dout(w_dff_A_H8oosr1I6_1),.din(w_dff_A_wbINvpvQ9_1),.clk(gclk));
	jdff dff_A_ibJ16uri5_2(.dout(w_G183gat_0[2]),.din(w_dff_A_ibJ16uri5_2),.clk(gclk));
	jdff dff_A_USHhy8Zp4_2(.dout(w_dff_A_ibJ16uri5_2),.din(w_dff_A_USHhy8Zp4_2),.clk(gclk));
	jdff dff_A_pUoGMm6J3_2(.dout(w_dff_A_USHhy8Zp4_2),.din(w_dff_A_pUoGMm6J3_2),.clk(gclk));
	jdff dff_A_y0tuKOT93_2(.dout(w_dff_A_pUoGMm6J3_2),.din(w_dff_A_y0tuKOT93_2),.clk(gclk));
	jdff dff_A_EnOzxcB10_2(.dout(w_dff_A_y0tuKOT93_2),.din(w_dff_A_EnOzxcB10_2),.clk(gclk));
	jdff dff_A_SOYVUpiV3_2(.dout(w_dff_A_EnOzxcB10_2),.din(w_dff_A_SOYVUpiV3_2),.clk(gclk));
	jdff dff_A_ofK71HAU6_0(.dout(w_n339_0[0]),.din(w_dff_A_ofK71HAU6_0),.clk(gclk));
	jdff dff_A_oNxFUwe10_0(.dout(w_dff_A_ofK71HAU6_0),.din(w_dff_A_oNxFUwe10_0),.clk(gclk));
	jdff dff_A_xyIK1zVJ4_0(.dout(w_dff_A_oNxFUwe10_0),.din(w_dff_A_xyIK1zVJ4_0),.clk(gclk));
	jdff dff_A_6ChR3N6F0_0(.dout(w_dff_A_xyIK1zVJ4_0),.din(w_dff_A_6ChR3N6F0_0),.clk(gclk));
	jdff dff_B_PEHi7lLT7_1(.din(n337),.dout(w_dff_B_PEHi7lLT7_1),.clk(gclk));
	jdff dff_B_5pYlq4ee6_1(.din(w_dff_B_PEHi7lLT7_1),.dout(w_dff_B_5pYlq4ee6_1),.clk(gclk));
	jdff dff_B_OhZtvwu41_1(.din(w_dff_B_5pYlq4ee6_1),.dout(w_dff_B_OhZtvwu41_1),.clk(gclk));
	jdff dff_B_BuP4IWfi8_1(.din(w_dff_B_OhZtvwu41_1),.dout(w_dff_B_BuP4IWfi8_1),.clk(gclk));
	jdff dff_B_uT4SdLTS5_1(.din(w_dff_B_BuP4IWfi8_1),.dout(w_dff_B_uT4SdLTS5_1),.clk(gclk));
	jdff dff_B_6NKaHX122_1(.din(w_dff_B_uT4SdLTS5_1),.dout(w_dff_B_6NKaHX122_1),.clk(gclk));
	jdff dff_A_xSUtLzvB8_2(.dout(w_n336_0[2]),.din(w_dff_A_xSUtLzvB8_2),.clk(gclk));
	jdff dff_A_PkRi1psv1_2(.dout(w_dff_A_xSUtLzvB8_2),.din(w_dff_A_PkRi1psv1_2),.clk(gclk));
	jdff dff_A_QzUVvIL82_2(.dout(w_dff_A_PkRi1psv1_2),.din(w_dff_A_QzUVvIL82_2),.clk(gclk));
	jdff dff_A_a8LNnxp19_2(.dout(w_dff_A_QzUVvIL82_2),.din(w_dff_A_a8LNnxp19_2),.clk(gclk));
	jdff dff_A_4jYozLls1_2(.dout(w_dff_A_a8LNnxp19_2),.din(w_dff_A_4jYozLls1_2),.clk(gclk));
	jdff dff_A_svH6yMxW8_2(.dout(w_dff_A_4jYozLls1_2),.din(w_dff_A_svH6yMxW8_2),.clk(gclk));
	jdff dff_A_Rr19MyhV6_2(.dout(w_dff_A_svH6yMxW8_2),.din(w_dff_A_Rr19MyhV6_2),.clk(gclk));
	jdff dff_A_8pmlUdXC8_2(.dout(w_dff_A_Rr19MyhV6_2),.din(w_dff_A_8pmlUdXC8_2),.clk(gclk));
	jdff dff_B_Fdm4RsM11_0(.din(n333),.dout(w_dff_B_Fdm4RsM11_0),.clk(gclk));
	jdff dff_B_s1Db8RCQ1_0(.din(n332),.dout(w_dff_B_s1Db8RCQ1_0),.clk(gclk));
	jdff dff_B_EdJFt1En8_0(.din(w_dff_B_s1Db8RCQ1_0),.dout(w_dff_B_EdJFt1En8_0),.clk(gclk));
	jdff dff_B_jIabbdRv7_0(.din(w_dff_B_EdJFt1En8_0),.dout(w_dff_B_jIabbdRv7_0),.clk(gclk));
	jdff dff_B_xfwW9Hcw6_0(.din(w_dff_B_jIabbdRv7_0),.dout(w_dff_B_xfwW9Hcw6_0),.clk(gclk));
	jdff dff_A_fvIu41ZS9_0(.dout(w_G153gat_0[0]),.din(w_dff_A_fvIu41ZS9_0),.clk(gclk));
	jdff dff_A_My0mWd8l0_0(.dout(w_dff_A_fvIu41ZS9_0),.din(w_dff_A_My0mWd8l0_0),.clk(gclk));
	jdff dff_A_cac9qL9k1_0(.dout(w_dff_A_My0mWd8l0_0),.din(w_dff_A_cac9qL9k1_0),.clk(gclk));
	jdff dff_A_xpiSFEr42_0(.dout(w_dff_A_cac9qL9k1_0),.din(w_dff_A_xpiSFEr42_0),.clk(gclk));
	jdff dff_A_tVlgc52J8_2(.dout(w_G153gat_0[2]),.din(w_dff_A_tVlgc52J8_2),.clk(gclk));
	jdff dff_A_SoFnZV9s5_2(.dout(w_dff_A_tVlgc52J8_2),.din(w_dff_A_SoFnZV9s5_2),.clk(gclk));
	jdff dff_A_lFsG8WrJ4_2(.dout(w_dff_A_SoFnZV9s5_2),.din(w_dff_A_lFsG8WrJ4_2),.clk(gclk));
	jdff dff_A_5PsbKJ721_2(.dout(w_dff_A_lFsG8WrJ4_2),.din(w_dff_A_5PsbKJ721_2),.clk(gclk));
	jdff dff_A_TyLSCsX71_0(.dout(w_G106gat_0[0]),.din(w_dff_A_TyLSCsX71_0),.clk(gclk));
	jdff dff_A_jHSDHRod4_0(.dout(w_dff_A_TyLSCsX71_0),.din(w_dff_A_jHSDHRod4_0),.clk(gclk));
	jdff dff_A_29S4EfEs0_0(.dout(w_dff_A_jHSDHRod4_0),.din(w_dff_A_29S4EfEs0_0),.clk(gclk));
	jdff dff_A_tDyp7s3m2_0(.dout(w_dff_A_29S4EfEs0_0),.din(w_dff_A_tDyp7s3m2_0),.clk(gclk));
	jdff dff_A_7RxM1HFo4_0(.dout(w_dff_A_tDyp7s3m2_0),.din(w_dff_A_7RxM1HFo4_0),.clk(gclk));
	jdff dff_A_Q5tBt3Dt9_1(.dout(w_G177gat_1[1]),.din(w_dff_A_Q5tBt3Dt9_1),.clk(gclk));
	jdff dff_A_E1zMHKly0_1(.dout(w_dff_A_Q5tBt3Dt9_1),.din(w_dff_A_E1zMHKly0_1),.clk(gclk));
	jdff dff_A_giy5uNC20_1(.dout(w_dff_A_E1zMHKly0_1),.din(w_dff_A_giy5uNC20_1),.clk(gclk));
	jdff dff_A_VzVE7bFf2_1(.dout(w_dff_A_giy5uNC20_1),.din(w_dff_A_VzVE7bFf2_1),.clk(gclk));
	jdff dff_A_i1d2TrVF8_1(.dout(w_dff_A_VzVE7bFf2_1),.din(w_dff_A_i1d2TrVF8_1),.clk(gclk));
	jdff dff_A_lUNGMeER4_1(.dout(w_dff_A_i1d2TrVF8_1),.din(w_dff_A_lUNGMeER4_1),.clk(gclk));
	jdff dff_A_2tKN5lYi4_1(.dout(w_G177gat_0[1]),.din(w_dff_A_2tKN5lYi4_1),.clk(gclk));
	jdff dff_A_2rwWqu043_1(.dout(w_dff_A_2tKN5lYi4_1),.din(w_dff_A_2rwWqu043_1),.clk(gclk));
	jdff dff_A_hFupe5IP8_1(.dout(w_dff_A_2rwWqu043_1),.din(w_dff_A_hFupe5IP8_1),.clk(gclk));
	jdff dff_A_HocxKQJ23_1(.dout(w_dff_A_hFupe5IP8_1),.din(w_dff_A_HocxKQJ23_1),.clk(gclk));
	jdff dff_A_01X2N3y46_2(.dout(w_G177gat_0[2]),.din(w_dff_A_01X2N3y46_2),.clk(gclk));
	jdff dff_A_UGQgXXv72_2(.dout(w_dff_A_01X2N3y46_2),.din(w_dff_A_UGQgXXv72_2),.clk(gclk));
	jdff dff_A_eflLSDKj8_2(.dout(w_dff_A_UGQgXXv72_2),.din(w_dff_A_eflLSDKj8_2),.clk(gclk));
	jdff dff_A_VddeiRVt5_2(.dout(w_dff_A_eflLSDKj8_2),.din(w_dff_A_VddeiRVt5_2),.clk(gclk));
	jdff dff_A_9voGgNWk1_2(.dout(w_dff_A_VddeiRVt5_2),.din(w_dff_A_9voGgNWk1_2),.clk(gclk));
	jdff dff_A_rKopKHok9_2(.dout(w_dff_A_9voGgNWk1_2),.din(w_dff_A_rKopKHok9_2),.clk(gclk));
	jdff dff_B_viTRVlxQ2_0(.din(n424),.dout(w_dff_B_viTRVlxQ2_0),.clk(gclk));
	jdff dff_A_jBnBKk4m9_0(.dout(w_G246gat_0[0]),.din(w_dff_A_jBnBKk4m9_0),.clk(gclk));
	jdff dff_A_J4srjupc3_0(.dout(w_dff_A_jBnBKk4m9_0),.din(w_dff_A_J4srjupc3_0),.clk(gclk));
	jdff dff_A_me8cEVlX2_0(.dout(w_dff_A_J4srjupc3_0),.din(w_dff_A_me8cEVlX2_0),.clk(gclk));
	jdff dff_A_m2fWDuOw9_0(.dout(w_dff_A_me8cEVlX2_0),.din(w_dff_A_m2fWDuOw9_0),.clk(gclk));
	jdff dff_A_XvYe7sEs4_0(.dout(w_dff_A_m2fWDuOw9_0),.din(w_dff_A_XvYe7sEs4_0),.clk(gclk));
	jdff dff_A_hSenj8Fx6_2(.dout(w_G246gat_0[2]),.din(w_dff_A_hSenj8Fx6_2),.clk(gclk));
	jdff dff_A_pEiVFWVm5_2(.dout(w_dff_A_hSenj8Fx6_2),.din(w_dff_A_pEiVFWVm5_2),.clk(gclk));
	jdff dff_A_cWUMsuP71_2(.dout(w_dff_A_pEiVFWVm5_2),.din(w_dff_A_cWUMsuP71_2),.clk(gclk));
	jdff dff_A_XTSl5f3d1_2(.dout(w_dff_A_cWUMsuP71_2),.din(w_dff_A_XTSl5f3d1_2),.clk(gclk));
	jdff dff_A_dio62ymb4_2(.dout(w_dff_A_XTSl5f3d1_2),.din(w_dff_A_dio62ymb4_2),.clk(gclk));
	jdff dff_B_ML60B5756_3(.din(G246gat),.dout(w_dff_B_ML60B5756_3),.clk(gclk));
	jdff dff_B_Bgn1qL6f9_0(.din(n422),.dout(w_dff_B_Bgn1qL6f9_0),.clk(gclk));
	jdff dff_B_YSglphc89_0(.din(w_dff_B_Bgn1qL6f9_0),.dout(w_dff_B_YSglphc89_0),.clk(gclk));
	jdff dff_B_0gGQ4aty2_0(.din(w_dff_B_YSglphc89_0),.dout(w_dff_B_0gGQ4aty2_0),.clk(gclk));
	jdff dff_B_DowX2YEs5_0(.din(w_dff_B_0gGQ4aty2_0),.dout(w_dff_B_DowX2YEs5_0),.clk(gclk));
	jdff dff_B_dFK2gmNP0_0(.din(w_dff_B_DowX2YEs5_0),.dout(w_dff_B_dFK2gmNP0_0),.clk(gclk));
	jdff dff_B_UyXzk69G3_0(.din(w_dff_B_dFK2gmNP0_0),.dout(w_dff_B_UyXzk69G3_0),.clk(gclk));
	jdff dff_B_sKQwZKGO0_0(.din(w_dff_B_UyXzk69G3_0),.dout(w_dff_B_sKQwZKGO0_0),.clk(gclk));
	jdff dff_A_3S1ZAduI2_1(.dout(w_G96gat_0[1]),.din(w_dff_A_3S1ZAduI2_1),.clk(gclk));
	jdff dff_A_6NDJ6yQb2_1(.dout(w_dff_A_3S1ZAduI2_1),.din(w_dff_A_6NDJ6yQb2_1),.clk(gclk));
	jdff dff_A_eTmUPtl63_1(.dout(w_dff_A_6NDJ6yQb2_1),.din(w_dff_A_eTmUPtl63_1),.clk(gclk));
	jdff dff_A_aJpXrbLV9_1(.dout(w_dff_A_eTmUPtl63_1),.din(w_dff_A_aJpXrbLV9_1),.clk(gclk));
	jdff dff_A_jJ3Agiua5_1(.dout(w_dff_A_aJpXrbLV9_1),.din(w_dff_A_jJ3Agiua5_1),.clk(gclk));
	jdff dff_A_0cWndKis9_0(.dout(w_n420_0[0]),.din(w_dff_A_0cWndKis9_0),.clk(gclk));
	jdff dff_A_819gHp0h9_0(.dout(w_dff_A_0cWndKis9_0),.din(w_dff_A_819gHp0h9_0),.clk(gclk));
	jdff dff_A_Oac5nl3V1_0(.dout(w_dff_A_819gHp0h9_0),.din(w_dff_A_Oac5nl3V1_0),.clk(gclk));
	jdff dff_A_dfgJzSTR9_0(.dout(w_dff_A_Oac5nl3V1_0),.din(w_dff_A_dfgJzSTR9_0),.clk(gclk));
	jdff dff_A_oZNfvIV19_0(.dout(w_dff_A_dfgJzSTR9_0),.din(w_dff_A_oZNfvIV19_0),.clk(gclk));
	jdff dff_A_pv6Llxho5_0(.dout(w_dff_A_oZNfvIV19_0),.din(w_dff_A_pv6Llxho5_0),.clk(gclk));
	jdff dff_A_NZNGj85j5_0(.dout(w_dff_A_pv6Llxho5_0),.din(w_dff_A_NZNGj85j5_0),.clk(gclk));
	jdff dff_A_pXiBHGgW9_0(.dout(w_dff_A_NZNGj85j5_0),.din(w_dff_A_pXiBHGgW9_0),.clk(gclk));
	jdff dff_B_Zz8qS1RX9_3(.din(G228gat),.dout(w_dff_B_Zz8qS1RX9_3),.clk(gclk));
	jdff dff_B_zYXFjQ8f0_3(.din(w_dff_B_Zz8qS1RX9_3),.dout(w_dff_B_zYXFjQ8f0_3),.clk(gclk));
	jdff dff_B_FCpXZ9jE2_3(.din(w_dff_B_zYXFjQ8f0_3),.dout(w_dff_B_FCpXZ9jE2_3),.clk(gclk));
	jdff dff_B_yayIqxlm6_3(.din(w_dff_B_FCpXZ9jE2_3),.dout(w_dff_B_yayIqxlm6_3),.clk(gclk));
	jdff dff_B_6N5lYVNw8_3(.din(w_dff_B_yayIqxlm6_3),.dout(w_dff_B_6N5lYVNw8_3),.clk(gclk));
	jdff dff_B_AqJWYsQB9_3(.din(w_dff_B_6N5lYVNw8_3),.dout(w_dff_B_AqJWYsQB9_3),.clk(gclk));
	jdff dff_B_PKDSliMz0_3(.din(w_dff_B_AqJWYsQB9_3),.dout(w_dff_B_PKDSliMz0_3),.clk(gclk));
	jdff dff_B_aSMCM9EO5_0(.din(n325),.dout(w_dff_B_aSMCM9EO5_0),.clk(gclk));
	jdff dff_B_4QqzGzgF3_0(.din(n324),.dout(w_dff_B_4QqzGzgF3_0),.clk(gclk));
	jdff dff_B_O7heLr722_0(.din(w_dff_B_4QqzGzgF3_0),.dout(w_dff_B_O7heLr722_0),.clk(gclk));
	jdff dff_B_rR21cPeg6_0(.din(w_dff_B_O7heLr722_0),.dout(w_dff_B_rR21cPeg6_0),.clk(gclk));
	jdff dff_B_MSQsjCHr1_0(.din(w_dff_B_rR21cPeg6_0),.dout(w_dff_B_MSQsjCHr1_0),.clk(gclk));
	jdff dff_A_dOndz9hd4_1(.dout(w_n167_0[1]),.din(w_dff_A_dOndz9hd4_1),.clk(gclk));
	jdff dff_B_cxQVaFZO1_2(.din(G149gat),.dout(w_dff_B_cxQVaFZO1_2),.clk(gclk));
	jdff dff_B_Ts7w3xfM1_2(.din(w_dff_B_cxQVaFZO1_2),.dout(w_dff_B_Ts7w3xfM1_2),.clk(gclk));
	jdff dff_B_PZTWlNOE1_2(.din(w_dff_B_Ts7w3xfM1_2),.dout(w_dff_B_PZTWlNOE1_2),.clk(gclk));
	jdff dff_B_yWvWJbNP7_2(.din(w_dff_B_PZTWlNOE1_2),.dout(w_dff_B_yWvWJbNP7_2),.clk(gclk));
	jdff dff_B_S6JGZ4BK1_0(.din(n163),.dout(w_dff_B_S6JGZ4BK1_0),.clk(gclk));
	jdff dff_B_3Mit8GXY2_0(.din(w_dff_B_S6JGZ4BK1_0),.dout(w_dff_B_3Mit8GXY2_0),.clk(gclk));
	jdff dff_B_uBWyZ4wu8_1(.din(n150),.dout(w_dff_B_uBWyZ4wu8_1),.clk(gclk));
	jdff dff_A_EuLMJAVz8_1(.dout(w_n151_0[1]),.din(w_dff_A_EuLMJAVz8_1),.clk(gclk));
	jdff dff_A_XDrhQoL33_0(.dout(w_G42gat_1[0]),.din(w_dff_A_XDrhQoL33_0),.clk(gclk));
	jdff dff_A_svFjUYC56_2(.dout(w_G17gat_2[2]),.din(w_dff_A_svFjUYC56_2),.clk(gclk));
	jdff dff_A_8o2GDxRU3_2(.dout(w_dff_A_svFjUYC56_2),.din(w_dff_A_8o2GDxRU3_2),.clk(gclk));
	jdff dff_A_HBKRtCN28_1(.dout(w_G101gat_0[1]),.din(w_dff_A_HBKRtCN28_1),.clk(gclk));
	jdff dff_A_CGNMA64Z8_1(.dout(w_dff_A_HBKRtCN28_1),.din(w_dff_A_CGNMA64Z8_1),.clk(gclk));
	jdff dff_A_sojqwtga4_1(.dout(w_dff_A_CGNMA64Z8_1),.din(w_dff_A_sojqwtga4_1),.clk(gclk));
	jdff dff_A_kIJH5AZc0_1(.dout(w_dff_A_sojqwtga4_1),.din(w_dff_A_kIJH5AZc0_1),.clk(gclk));
	jdff dff_A_5QQC5bE49_1(.dout(w_dff_A_kIJH5AZc0_1),.din(w_dff_A_5QQC5bE49_1),.clk(gclk));
	jdff dff_A_GzPcAlQd1_2(.dout(w_G447gat_0[2]),.din(w_dff_A_GzPcAlQd1_2),.clk(gclk));
	jdff dff_A_tZhBeJBZ3_1(.dout(w_G51gat_1[1]),.din(w_dff_A_tZhBeJBZ3_1),.clk(gclk));
	jdff dff_A_rMq5VKvg8_0(.dout(w_G80gat_0[0]),.din(w_dff_A_rMq5VKvg8_0),.clk(gclk));
	jdff dff_A_75Zmf9AN2_0(.dout(w_dff_A_rMq5VKvg8_0),.din(w_dff_A_75Zmf9AN2_0),.clk(gclk));
	jdff dff_A_2b6CFqz22_2(.dout(w_G80gat_0[2]),.din(w_dff_A_2b6CFqz22_2),.clk(gclk));
	jdff dff_A_HumMNYpW3_0(.dout(w_n86_0[0]),.din(w_dff_A_HumMNYpW3_0),.clk(gclk));
	jdff dff_A_8YW7iErV4_0(.dout(w_dff_A_HumMNYpW3_0),.din(w_dff_A_8YW7iErV4_0),.clk(gclk));
	jdff dff_A_oWqVhi8U0_0(.dout(w_G29gat_0[0]),.din(w_dff_A_oWqVhi8U0_0),.clk(gclk));
	jdff dff_A_k2hAoUcH6_0(.dout(w_dff_A_oWqVhi8U0_0),.din(w_dff_A_k2hAoUcH6_0),.clk(gclk));
	jdff dff_A_U5kbN1Si1_0(.dout(w_dff_A_k2hAoUcH6_0),.din(w_dff_A_U5kbN1Si1_0),.clk(gclk));
	jdff dff_A_F5JMnWxN1_0(.dout(w_G17gat_1[0]),.din(w_dff_A_F5JMnWxN1_0),.clk(gclk));
	jdff dff_A_OYHwywK25_0(.dout(w_dff_A_F5JMnWxN1_0),.din(w_dff_A_OYHwywK25_0),.clk(gclk));
	jdff dff_A_ra75qUdI7_0(.dout(w_dff_A_OYHwywK25_0),.din(w_dff_A_ra75qUdI7_0),.clk(gclk));
	jdff dff_A_kGD97uD18_0(.dout(w_dff_A_ra75qUdI7_0),.din(w_dff_A_kGD97uD18_0),.clk(gclk));
	jdff dff_A_s4RucgmH5_1(.dout(w_G17gat_1[1]),.din(w_dff_A_s4RucgmH5_1),.clk(gclk));
	jdff dff_A_F6szztgT6_1(.dout(w_dff_A_s4RucgmH5_1),.din(w_dff_A_F6szztgT6_1),.clk(gclk));
	jdff dff_A_R3mMVGf93_1(.dout(w_dff_A_F6szztgT6_1),.din(w_dff_A_R3mMVGf93_1),.clk(gclk));
	jdff dff_B_6a7pafLu0_2(.din(n144),.dout(w_dff_B_6a7pafLu0_2),.clk(gclk));
	jdff dff_B_Z6YaJEQ33_2(.din(w_dff_B_6a7pafLu0_2),.dout(w_dff_B_Z6YaJEQ33_2),.clk(gclk));
	jdff dff_B_SNIlPIe11_2(.din(w_dff_B_Z6YaJEQ33_2),.dout(w_dff_B_SNIlPIe11_2),.clk(gclk));
	jdff dff_B_nqtVZAax0_2(.din(w_dff_B_SNIlPIe11_2),.dout(w_dff_B_nqtVZAax0_2),.clk(gclk));
	jdff dff_A_nKhPqxsF5_0(.dout(w_G237gat_0[0]),.din(w_dff_A_nKhPqxsF5_0),.clk(gclk));
	jdff dff_A_TfErT3cr0_0(.dout(w_dff_A_nKhPqxsF5_0),.din(w_dff_A_TfErT3cr0_0),.clk(gclk));
	jdff dff_A_7P5OOGI81_0(.dout(w_dff_A_TfErT3cr0_0),.din(w_dff_A_7P5OOGI81_0),.clk(gclk));
	jdff dff_A_wN3TuHHf4_0(.dout(w_dff_A_7P5OOGI81_0),.din(w_dff_A_wN3TuHHf4_0),.clk(gclk));
	jdff dff_A_eD2zl0ft8_0(.dout(w_dff_A_wN3TuHHf4_0),.din(w_dff_A_eD2zl0ft8_0),.clk(gclk));
	jdff dff_A_3StBpSnb5_0(.dout(w_dff_A_eD2zl0ft8_0),.din(w_dff_A_3StBpSnb5_0),.clk(gclk));
	jdff dff_A_Ms4I4KGx6_2(.dout(w_G237gat_0[2]),.din(w_dff_A_Ms4I4KGx6_2),.clk(gclk));
	jdff dff_A_j3KPQP6N1_2(.dout(w_dff_A_Ms4I4KGx6_2),.din(w_dff_A_j3KPQP6N1_2),.clk(gclk));
	jdff dff_A_QXsUzNsy5_2(.dout(w_dff_A_j3KPQP6N1_2),.din(w_dff_A_QXsUzNsy5_2),.clk(gclk));
	jdff dff_A_zz3gx5pR3_2(.dout(w_dff_A_QXsUzNsy5_2),.din(w_dff_A_zz3gx5pR3_2),.clk(gclk));
	jdff dff_A_aD3vSyb00_2(.dout(w_dff_A_zz3gx5pR3_2),.din(w_dff_A_aD3vSyb00_2),.clk(gclk));
	jdff dff_A_YjhNPzNL6_2(.dout(w_dff_A_aD3vSyb00_2),.din(w_dff_A_YjhNPzNL6_2),.clk(gclk));
	jdff dff_A_DwycHNr98_2(.dout(w_dff_A_YjhNPzNL6_2),.din(w_dff_A_DwycHNr98_2),.clk(gclk));
	jdff dff_A_JpqlyuDb6_0(.dout(w_n178_0[0]),.din(w_dff_A_JpqlyuDb6_0),.clk(gclk));
	jdff dff_A_LTmUMlhz6_0(.dout(w_dff_A_JpqlyuDb6_0),.din(w_dff_A_LTmUMlhz6_0),.clk(gclk));
	jdff dff_A_xHTspfHT1_0(.dout(w_dff_A_LTmUMlhz6_0),.din(w_dff_A_xHTspfHT1_0),.clk(gclk));
	jdff dff_B_MqzXXQpS0_0(.din(n176),.dout(w_dff_B_MqzXXQpS0_0),.clk(gclk));
	jdff dff_A_5mOXuFtE3_1(.dout(w_n122_0[1]),.din(w_dff_A_5mOXuFtE3_1),.clk(gclk));
	jdff dff_A_uX1ST8167_1(.dout(w_dff_A_5mOXuFtE3_1),.din(w_dff_A_uX1ST8167_1),.clk(gclk));
	jdff dff_A_Cw9lnBBc6_1(.dout(w_dff_A_uX1ST8167_1),.din(w_dff_A_Cw9lnBBc6_1),.clk(gclk));
	jdff dff_A_z6M065IR9_1(.dout(w_G68gat_0[1]),.din(w_dff_A_z6M065IR9_1),.clk(gclk));
	jdff dff_A_IxRrFqPx2_1(.dout(w_dff_A_z6M065IR9_1),.din(w_dff_A_IxRrFqPx2_1),.clk(gclk));
	jdff dff_A_uUTggaeS6_1(.dout(w_dff_A_IxRrFqPx2_1),.din(w_dff_A_uUTggaeS6_1),.clk(gclk));
	jdff dff_A_7uPyF1rD4_1(.dout(w_dff_A_uUTggaeS6_1),.din(w_dff_A_7uPyF1rD4_1),.clk(gclk));
	jdff dff_A_Okid8rW94_1(.dout(w_G42gat_0[1]),.din(w_dff_A_Okid8rW94_1),.clk(gclk));
	jdff dff_A_tuOdJaz41_2(.dout(w_G42gat_0[2]),.din(w_dff_A_tuOdJaz41_2),.clk(gclk));
	jdff dff_A_iCl7TOn50_1(.dout(w_G1gat_0[1]),.din(w_dff_A_iCl7TOn50_1),.clk(gclk));
	jdff dff_A_hw9j201Q8_1(.dout(w_G13gat_0[1]),.din(w_dff_A_hw9j201Q8_1),.clk(gclk));
	jdff dff_A_YW6fEiix2_0(.dout(w_G55gat_0[0]),.din(w_dff_A_YW6fEiix2_0),.clk(gclk));
	jdff dff_A_z1Q9CbA68_1(.dout(w_G55gat_0[1]),.din(w_dff_A_z1Q9CbA68_1),.clk(gclk));
	jdff dff_A_nmfxa6Js2_1(.dout(w_dff_A_z1Q9CbA68_1),.din(w_dff_A_nmfxa6Js2_1),.clk(gclk));
	jdff dff_B_mL6ahJM19_3(.din(G55gat),.dout(w_dff_B_mL6ahJM19_3),.clk(gclk));
	jdff dff_B_i5JhTpjB3_3(.din(w_dff_B_mL6ahJM19_3),.dout(w_dff_B_i5JhTpjB3_3),.clk(gclk));
	jdff dff_A_5NJTiXpF1_1(.dout(w_G171gat_0[1]),.din(w_dff_A_5NJTiXpF1_1),.clk(gclk));
	jdff dff_A_nKiX7A6H8_1(.dout(w_dff_A_5NJTiXpF1_1),.din(w_dff_A_nKiX7A6H8_1),.clk(gclk));
	jdff dff_A_sBEqGzWZ3_1(.dout(w_dff_A_nKiX7A6H8_1),.din(w_dff_A_sBEqGzWZ3_1),.clk(gclk));
	jdff dff_A_AWASG99i6_1(.dout(w_dff_A_sBEqGzWZ3_1),.din(w_dff_A_AWASG99i6_1),.clk(gclk));
	jdff dff_A_Q5vtmiXM1_1(.dout(w_dff_A_AWASG99i6_1),.din(w_dff_A_Q5vtmiXM1_1),.clk(gclk));
	jdff dff_A_pkWdKiuy2_1(.dout(w_dff_A_Q5vtmiXM1_1),.din(w_dff_A_pkWdKiuy2_1),.clk(gclk));
	jdff dff_A_qgJr1mYT1_2(.dout(w_G171gat_0[2]),.din(w_dff_A_qgJr1mYT1_2),.clk(gclk));
	jdff dff_A_UlNQ7CI57_2(.dout(w_dff_A_qgJr1mYT1_2),.din(w_dff_A_UlNQ7CI57_2),.clk(gclk));
	jdff dff_A_WoO4NXHP1_2(.dout(w_dff_A_UlNQ7CI57_2),.din(w_dff_A_WoO4NXHP1_2),.clk(gclk));
	jdff dff_A_ZSdoUlp44_2(.dout(w_dff_A_WoO4NXHP1_2),.din(w_dff_A_ZSdoUlp44_2),.clk(gclk));
	jdff dff_A_1aAZXfux4_2(.dout(w_dff_A_ZSdoUlp44_2),.din(w_dff_A_1aAZXfux4_2),.clk(gclk));
	jdff dff_A_iscgakJ79_2(.dout(w_dff_A_1aAZXfux4_2),.din(w_dff_A_iscgakJ79_2),.clk(gclk));
	jdff dff_A_4MhYOLGE7_2(.dout(w_dff_A_iscgakJ79_2),.din(w_dff_A_4MhYOLGE7_2),.clk(gclk));
endmodule

