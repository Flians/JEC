/*

c1908:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 1045
	jand: 128
	jor: 102

Summary:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 1045
	jand: 128
	jor: 102
*/

module c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n202;
	wire n204;
	wire n205;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n222;
	wire n224;
	wire n225;
	wire n226;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire [2:0] w_G101_0;
	wire [2:0] w_G104_0;
	wire [2:0] w_G107_0;
	wire [2:0] w_G110_0;
	wire [1:0] w_G110_1;
	wire [1:0] w_G113_0;
	wire [2:0] w_G116_0;
	wire [2:0] w_G119_0;
	wire [2:0] w_G122_0;
	wire [1:0] w_G122_1;
	wire [2:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [1:0] w_G128_1;
	wire [1:0] w_G131_0;
	wire [2:0] w_G134_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G140_0;
	wire [2:0] w_G143_0;
	wire [1:0] w_G143_1;
	wire [2:0] w_G146_0;
	wire [2:0] w_G210_0;
	wire [1:0] w_G214_0;
	wire [2:0] w_G217_0;
	wire [1:0] w_G221_0;
	wire [1:0] w_G224_0;
	wire [1:0] w_G227_0;
	wire [2:0] w_G234_0;
	wire [2:0] w_G237_0;
	wire [2:0] w_G469_0;
	wire [1:0] w_G472_0;
	wire [2:0] w_G475_0;
	wire [2:0] w_G478_0;
	wire [2:0] w_G902_0;
	wire [2:0] w_G902_1;
	wire [2:0] w_G902_2;
	wire [2:0] w_G902_3;
	wire [2:0] w_G952_0;
	wire [2:0] w_G953_0;
	wire [2:0] w_G953_1;
	wire [1:0] w_n59_0;
	wire [2:0] w_n60_0;
	wire [2:0] w_n61_0;
	wire [2:0] w_n61_1;
	wire [2:0] w_n61_2;
	wire [2:0] w_n61_3;
	wire [1:0] w_n62_0;
	wire [1:0] w_n67_0;
	wire [1:0] w_n68_0;
	wire [2:0] w_n70_0;
	wire [2:0] w_n70_1;
	wire [2:0] w_n70_2;
	wire [1:0] w_n70_3;
	wire [1:0] w_n71_0;
	wire [1:0] w_n73_0;
	wire [2:0] w_n74_0;
	wire [1:0] w_n74_1;
	wire [1:0] w_n77_0;
	wire [1:0] w_n79_0;
	wire [2:0] w_n81_0;
	wire [1:0] w_n82_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [2:0] w_n90_0;
	wire [2:0] w_n92_0;
	wire [2:0] w_n92_1;
	wire [2:0] w_n93_0;
	wire [1:0] w_n94_0;
	wire [2:0] w_n95_0;
	wire [2:0] w_n96_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [2:0] w_n107_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [2:0] w_n110_0;
	wire [2:0] w_n112_0;
	wire [1:0] w_n112_1;
	wire [2:0] w_n117_0;
	wire [1:0] w_n118_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [2:0] w_n121_0;
	wire [1:0] w_n121_1;
	wire [1:0] w_n122_0;
	wire [2:0] w_n130_0;
	wire [1:0] w_n131_0;
	wire [2:0] w_n132_0;
	wire [2:0] w_n141_0;
	wire [1:0] w_n142_0;
	wire [2:0] w_n143_0;
	wire [1:0] w_n143_1;
	wire [2:0] w_n144_0;
	wire [2:0] w_n144_1;
	wire [1:0] w_n145_0;
	wire [1:0] w_n146_0;
	wire [1:0] w_n147_0;
	wire [2:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n154_0;
	wire [1:0] w_n154_1;
	wire [2:0] w_n155_0;
	wire [1:0] w_n156_0;
	wire [2:0] w_n158_0;
	wire [1:0] w_n158_1;
	wire [2:0] w_n159_0;
	wire [1:0] w_n159_1;
	wire [1:0] w_n160_0;
	wire [2:0] w_n161_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n164_0;
	wire [2:0] w_n166_0;
	wire [1:0] w_n166_1;
	wire [1:0] w_n167_0;
	wire [2:0] w_n168_0;
	wire [1:0] w_n169_0;
	wire [1:0] w_n172_0;
	wire [2:0] w_n174_0;
	wire [1:0] w_n174_1;
	wire [1:0] w_n175_0;
	wire [1:0] w_n177_0;
	wire [2:0] w_n179_0;
	wire [1:0] w_n180_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n183_0;
	wire [2:0] w_n184_0;
	wire [1:0] w_n184_1;
	wire [2:0] w_n185_0;
	wire [1:0] w_n186_0;
	wire [2:0] w_n188_0;
	wire [1:0] w_n189_0;
	wire [1:0] w_n190_0;
	wire [2:0] w_n192_0;
	wire [1:0] w_n193_0;
	wire [2:0] w_n196_0;
	wire [2:0] w_n197_0;
	wire [1:0] w_n197_1;
	wire [2:0] w_n198_0;
	wire [1:0] w_n198_1;
	wire [1:0] w_n199_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n210_0;
	wire [1:0] w_n212_0;
	wire [1:0] w_n213_0;
	wire [2:0] w_n216_0;
	wire [2:0] w_n217_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [1:0] w_n219_0;
	wire [1:0] w_n220_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n226_0;
	wire [1:0] w_n228_0;
	wire [2:0] w_n244_0;
	wire [2:0] w_n244_1;
	wire [2:0] w_n244_2;
	wire [1:0] w_n252_0;
	wire [2:0] w_n253_0;
	wire [2:0] w_n254_0;
	wire [1:0] w_n254_1;
	wire [2:0] w_n273_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n275_0;
	wire [2:0] w_n276_0;
	wire [1:0] w_n276_1;
	wire [1:0] w_n277_0;
	wire [1:0] w_n278_0;
	wire [1:0] w_n280_0;
	wire [2:0] w_n281_0;
	wire [1:0] w_n282_0;
	wire [1:0] w_n286_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n289_0;
	wire [2:0] w_n290_0;
	wire [1:0] w_n291_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n309_0;
	wire [2:0] w_n311_0;
	wire [2:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n318_0;
	wire [1:0] w_n325_0;
	wire [1:0] w_n334_0;
	wire [2:0] w_n335_0;
	wire [2:0] w_n335_1;
	wire [1:0] w_n335_2;
	wire [1:0] w_n336_0;
	wire [2:0] w_n340_0;
	wire [2:0] w_n340_1;
	wire [1:0] w_n340_2;
	wire [1:0] w_n346_0;
	wire [1:0] w_n355_0;
	wire [1:0] w_n364_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n395_0;
	wire w_dff_B_6Tj43yLD7_0;
	wire w_dff_B_bkhnxK0n9_0;
	wire w_dff_B_mEmd24zc6_0;
	wire w_dff_B_aohSYRY50_0;
	wire w_dff_B_nGg3Q8VT6_0;
	wire w_dff_B_KYoJ6tCB8_0;
	wire w_dff_B_Lg0smOrj5_0;
	wire w_dff_B_ni4xBugN4_0;
	wire w_dff_B_Y771JsgA5_1;
	wire w_dff_B_UiVPnDn26_1;
	wire w_dff_B_8aigdvcU2_0;
	wire w_dff_B_mgpfL50U4_0;
	wire w_dff_A_XRjJXcUI0_1;
	wire w_dff_B_oMDeVr7b5_2;
	wire w_dff_B_f3bEe1Gh2_2;
	wire w_dff_B_piq5rTZj4_0;
	wire w_dff_B_vfSLBcRq1_0;
	wire w_dff_B_1psTim966_1;
	wire w_dff_B_fiJZxm4Z8_1;
	wire w_dff_B_keQD9Y6l7_1;
	wire w_dff_B_YCEUnVpZ7_1;
	wire w_dff_B_mD4x9hcs7_1;
	wire w_dff_B_dBMhKthn9_1;
	wire w_dff_B_GS8B36zJ7_1;
	wire w_dff_B_k1OSsfpz5_1;
	wire w_dff_B_c0cDSTjj5_1;
	wire w_dff_B_Wze0wzyd2_1;
	wire w_dff_B_rEFRVGKw1_1;
	wire w_dff_B_1ENNgSjZ1_1;
	wire w_dff_B_r8UYE5iT4_0;
	wire w_dff_B_5ETLHI0A6_0;
	wire w_dff_B_dUZCs7jr5_0;
	wire w_dff_B_AKSEso6s7_0;
	wire w_dff_B_DFzpmXxf4_0;
	wire w_dff_B_SsbS50495_0;
	wire w_dff_B_0NZxvEWX1_0;
	wire w_dff_B_2jxfQ34O3_0;
	wire w_dff_B_jEKe9zsj7_0;
	wire w_dff_B_deEBEmzQ3_0;
	wire w_dff_B_AR45nFuG8_0;
	wire w_dff_B_3E35odDm8_0;
	wire w_dff_B_JOhpdqEq1_0;
	wire w_dff_B_HuwMTHLf4_0;
	wire w_dff_A_xXznSd8I7_0;
	wire w_dff_A_6OrMfaJ90_0;
	wire w_dff_A_YmAvIMiq7_0;
	wire w_dff_A_t5Bh1HlL3_0;
	wire w_dff_A_PgDBrITs1_0;
	wire w_dff_A_Rzc3NOqW3_0;
	wire w_dff_A_c5pUAJpm7_0;
	wire w_dff_A_DhkEh3MU5_0;
	wire w_dff_A_hkU1notJ6_0;
	wire w_dff_A_KgHCMNRE3_0;
	wire w_dff_A_Bkj0KmFw3_0;
	wire w_dff_A_LJaleAfG1_0;
	wire w_dff_A_xV6AHXxs7_0;
	wire w_dff_A_TZZwCy5l3_0;
	wire w_dff_A_Z2vaiXFp1_0;
	wire w_dff_B_g2OF9prz8_1;
	wire w_dff_B_VEhLCr7G7_1;
	wire w_dff_B_XWBnabPj0_1;
	wire w_dff_B_SzE7DbvA0_1;
	wire w_dff_B_lrpHZXCg6_1;
	wire w_dff_B_idg45rYp0_1;
	wire w_dff_B_t6MrdRp72_1;
	wire w_dff_B_FaUJ5Y8Z3_1;
	wire w_dff_B_ZraIwppx8_1;
	wire w_dff_B_ELXaCA7H8_1;
	wire w_dff_B_6bEnps496_1;
	wire w_dff_B_9Nqzcnkn1_1;
	wire w_dff_B_H2CNrLJG0_0;
	wire w_dff_B_Y0JdRT1V6_0;
	wire w_dff_B_D6MFdtx69_0;
	wire w_dff_B_EfToIRyC9_0;
	wire w_dff_B_bg2glnvm3_0;
	wire w_dff_B_4tq0zEbH0_0;
	wire w_dff_B_EeBHlsE48_0;
	wire w_dff_B_aKeyEGGf3_0;
	wire w_dff_B_K5RX96Or7_0;
	wire w_dff_B_1qgJAdzW0_0;
	wire w_dff_B_ZwQVbcg82_0;
	wire w_dff_B_Ych6BOQm9_0;
	wire w_dff_B_RVrt5Roe8_0;
	wire w_dff_B_x8rUjeRO8_0;
	wire w_dff_A_a40ZrbBV0_0;
	wire w_dff_A_KS9CbfIl9_0;
	wire w_dff_A_x1JrpnHu2_0;
	wire w_dff_A_PjeSSwbs7_0;
	wire w_dff_A_pqi7Lsm11_0;
	wire w_dff_A_eDeewrIT1_0;
	wire w_dff_A_9jk7Iiux0_0;
	wire w_dff_A_1952PmuC5_0;
	wire w_dff_A_k4K5yYP36_0;
	wire w_dff_A_2j38ThGE6_0;
	wire w_dff_A_UcdqNdcy2_0;
	wire w_dff_A_cXUyKw9F2_0;
	wire w_dff_A_WX7shqmk3_0;
	wire w_dff_A_eBCgRtde7_0;
	wire w_dff_A_R35ciefN3_0;
	wire w_dff_B_2zSnQfFs1_1;
	wire w_dff_B_l8X87IZS8_1;
	wire w_dff_B_DfWMo8wB9_1;
	wire w_dff_B_3g5Nk9NH1_1;
	wire w_dff_B_MA4W0IWu2_1;
	wire w_dff_B_SH0MrZEv1_1;
	wire w_dff_B_9bOzUXyW0_1;
	wire w_dff_B_o1sQQcrB5_1;
	wire w_dff_B_sMMOgGKX7_1;
	wire w_dff_B_6INdmnwJ1_1;
	wire w_dff_B_kskOGiI54_1;
	wire w_dff_B_asEVOhQ28_1;
	wire w_dff_B_JUyNBap41_0;
	wire w_dff_B_rSUV66cp1_0;
	wire w_dff_B_QyQySQpP7_0;
	wire w_dff_B_G1D6aLzB0_0;
	wire w_dff_B_t4xgzVOG1_0;
	wire w_dff_B_3kqAcaaz4_0;
	wire w_dff_B_31AUgmxW9_0;
	wire w_dff_B_Bms54Ufo4_0;
	wire w_dff_B_cYH2h23q3_0;
	wire w_dff_B_eeIkLifw7_0;
	wire w_dff_B_hNMRWYNp3_0;
	wire w_dff_B_sPE2No0Z4_0;
	wire w_dff_B_3voJP80T0_0;
	wire w_dff_B_pgBGJOFz1_0;
	wire w_dff_A_xcYwUVsO8_0;
	wire w_dff_A_N6lIisni1_0;
	wire w_dff_A_7jPaRy5k4_0;
	wire w_dff_A_ak4shpa80_0;
	wire w_dff_A_NyE7DK9t8_0;
	wire w_dff_A_qjrtIxys2_0;
	wire w_dff_A_HcpEG8lA1_0;
	wire w_dff_A_1yBdBzXG3_0;
	wire w_dff_A_MneI7HUb6_0;
	wire w_dff_A_craBofKo4_0;
	wire w_dff_A_GIk3ME9r6_0;
	wire w_dff_A_xIxoSfj75_0;
	wire w_dff_A_rVfHl5V13_0;
	wire w_dff_A_3m4Gm8CY2_0;
	wire w_dff_A_LrjQo2z18_0;
	wire w_dff_B_wmO4A6qe3_1;
	wire w_dff_B_jmLswqoX8_1;
	wire w_dff_B_9h9Ky1mg4_1;
	wire w_dff_B_deW99Fmt3_1;
	wire w_dff_B_J9o3XUjZ7_1;
	wire w_dff_B_fUReB4hX0_1;
	wire w_dff_B_cqtGVioD4_1;
	wire w_dff_B_OajuNvdD9_1;
	wire w_dff_B_q63v1enh3_1;
	wire w_dff_B_9aVBX27z9_1;
	wire w_dff_B_PFtwNMs62_1;
	wire w_dff_B_7HXfiGRz1_1;
	wire w_dff_B_wYPCkrPE6_0;
	wire w_dff_B_yCtKu4ji2_0;
	wire w_dff_B_v0X3FtpK1_0;
	wire w_dff_B_MlQIv1ZU5_0;
	wire w_dff_B_6kqHQUWw3_0;
	wire w_dff_B_SOYqLUKg1_0;
	wire w_dff_B_xjELT74o9_0;
	wire w_dff_B_rYcgpTRV5_0;
	wire w_dff_B_WtvNf9XZ2_0;
	wire w_dff_B_HjZuLwPn8_0;
	wire w_dff_B_KurlW3CV9_0;
	wire w_dff_B_fBMT03aO5_0;
	wire w_dff_B_YPb2xc1Q6_0;
	wire w_dff_B_QxqH7i8L4_0;
	wire w_dff_A_iOWFAiQM5_0;
	wire w_dff_A_EYuRxxkG1_0;
	wire w_dff_A_4tEwtDPz3_0;
	wire w_dff_A_3akT1Pd26_0;
	wire w_dff_A_cbYSRxgy4_0;
	wire w_dff_A_4ykiYK3i2_0;
	wire w_dff_A_kCMJas7z6_0;
	wire w_dff_A_InaOq4ub2_0;
	wire w_dff_A_g4RHG3ie2_0;
	wire w_dff_A_9ovgboK87_0;
	wire w_dff_A_VbPYCV4X0_0;
	wire w_dff_A_lKUXeGMP7_0;
	wire w_dff_A_FtDOVRwm1_0;
	wire w_dff_A_U6VZd5uT4_0;
	wire w_dff_A_g4DgAnzk9_0;
	wire w_dff_B_Z1UoXxNG6_1;
	wire w_dff_B_TR4RPDZZ8_0;
	wire w_dff_B_O6hyf5kI2_0;
	wire w_dff_B_frALq1aB9_0;
	wire w_dff_B_2scBKyAd7_0;
	wire w_dff_B_Y8c7gJsy9_0;
	wire w_dff_B_1q9kFu5r6_0;
	wire w_dff_B_1vfvWWWA0_0;
	wire w_dff_B_4kM0jMEn1_0;
	wire w_dff_B_QgX8oHX47_0;
	wire w_dff_B_p43JBJuH3_0;
	wire w_dff_B_71GvA6f68_0;
	wire w_dff_B_af2l6ZNy0_0;
	wire w_dff_B_ybnAZrxV0_0;
	wire w_dff_B_oWeEm77E3_0;
	wire w_dff_A_Nv30eQLC1_1;
	wire w_dff_A_xmggtavh0_1;
	wire w_dff_A_95ILcNr92_1;
	wire w_dff_A_SMEdqSmF8_1;
	wire w_dff_A_b2oZaGwc0_1;
	wire w_dff_A_GcyNs0mk0_1;
	wire w_dff_A_YsLtPPyd4_1;
	wire w_dff_A_BJg2hu6n1_1;
	wire w_dff_A_nCy55j0m5_1;
	wire w_dff_A_94VjiY8l0_1;
	wire w_dff_A_5PIyMaYk5_1;
	wire w_dff_A_AHCK4zuY1_1;
	wire w_dff_A_5S1WgPzl9_1;
	wire w_dff_A_q94WGlpI1_1;
	wire w_dff_A_cfi4m6ds0_1;
	wire w_dff_B_auJy2zN15_1;
	wire w_dff_B_qsfCuBTl5_1;
	wire w_dff_B_KziesRIi4_1;
	wire w_dff_B_oytCqnNi5_1;
	wire w_dff_B_BOPJdd9c7_1;
	wire w_dff_B_Yc330sQ48_1;
	wire w_dff_B_c1neUtE09_1;
	wire w_dff_B_ZoSHi2uY1_1;
	wire w_dff_B_WR5UWy2s3_1;
	wire w_dff_B_kRtO0J5R1_1;
	wire w_dff_B_zdCjIH5i0_1;
	wire w_dff_B_hZt06uKP7_1;
	wire w_dff_B_4XIhDDXP0_1;
	wire w_dff_B_GTdvnyGC8_1;
	wire w_dff_B_TEb94CHB0_1;
	wire w_dff_B_6soSkoXO6_0;
	wire w_dff_B_Y3w9aD0W7_0;
	wire w_dff_B_yKKNmLjm2_0;
	wire w_dff_B_3h6HTqAb8_0;
	wire w_dff_B_40FnlNyZ3_0;
	wire w_dff_B_MMFoMroI5_0;
	wire w_dff_B_8RR9m6Ve9_0;
	wire w_dff_B_9D8b6rVG3_0;
	wire w_dff_B_wu922Bbp0_0;
	wire w_dff_B_btWV6d8S1_0;
	wire w_dff_B_SDE0ZuKW0_0;
	wire w_dff_B_VutXt6i25_0;
	wire w_dff_B_q8s1OkMF9_0;
	wire w_dff_B_GsXdjJPE0_0;
	wire w_dff_B_twuoMNpP3_0;
	wire w_dff_B_TKpuWm7I1_0;
	wire w_dff_B_vDz0SzSY1_0;
	wire w_dff_B_NUY7oWDt9_0;
	wire w_dff_B_Esqf7SVr8_0;
	wire w_dff_B_z3NEQ4bB6_0;
	wire w_dff_B_qvxlqp2j2_0;
	wire w_dff_B_WEKewzHa9_0;
	wire w_dff_B_bbuANj3p2_0;
	wire w_dff_B_4sBnFaE23_0;
	wire w_dff_B_3ezn6Tq90_0;
	wire w_dff_B_Hc6JuZM87_1;
	wire w_dff_B_6PMUkzqF5_1;
	wire w_dff_B_SllIQFCA4_0;
	wire w_dff_B_zFtMBBRt8_0;
	wire w_dff_B_AhKVwmre3_0;
	wire w_dff_B_kppAuLRK1_0;
	wire w_dff_B_f0LYQgLJ5_0;
	wire w_dff_B_ArSjcsta0_0;
	wire w_dff_B_3cKr2Jdv2_0;
	wire w_dff_B_kMhhQDeI1_0;
	wire w_dff_B_K6MMRE9n1_0;
	wire w_dff_B_4swiCMCz1_0;
	wire w_dff_B_PfseflL70_0;
	wire w_dff_B_sHmvpdd74_0;
	wire w_dff_B_PeeA8JVj0_0;
	wire w_dff_B_HjcMotW98_1;
	wire w_dff_B_h0UcXPex1_0;
	wire w_dff_A_9ps5Vm5Q7_0;
	wire w_dff_A_IHqyDOlI7_0;
	wire w_dff_A_JWHs09d71_2;
	wire w_dff_A_LORqUJdb7_2;
	wire w_dff_A_NQaIJkRP2_0;
	wire w_dff_A_8q8lNVYD4_2;
	wire w_dff_B_i6lhBmlg3_3;
	wire w_dff_B_mFbBRedQ8_0;
	wire w_dff_A_zDeAIA3f6_0;
	wire w_dff_A_mnwbm1S54_2;
	wire w_dff_A_HaA4EzaU8_2;
	wire w_dff_A_q3Bn0c1F6_0;
	wire w_dff_A_hiMHTam68_0;
	wire w_dff_A_tUnjq15O9_1;
	wire w_dff_A_H7gxCzUt6_1;
	wire w_dff_A_ppa3Ic6i2_0;
	wire w_dff_A_BItCi9uA1_2;
	wire w_dff_B_UBOMW93A9_3;
	wire w_dff_A_jmnqiUNg7_0;
	wire w_dff_A_4Gp49ERV3_0;
	wire w_dff_A_kmByPNTj0_1;
	wire w_dff_A_2KEevYyh8_1;
	wire w_dff_A_JLyGu4V98_2;
	wire w_dff_A_MLI46m0M2_2;
	wire w_dff_A_0CYnpiTc0_2;
	wire w_dff_B_Vs822WDe7_3;
	wire w_dff_A_ZeOdPqkX6_1;
	wire w_dff_A_VfQnigIX0_1;
	wire w_dff_A_95ZYmOEK6_1;
	wire w_dff_A_ArFhudP54_1;
	wire w_dff_A_BppLuG0Q2_2;
	wire w_dff_A_q0ph1p8R6_2;
	wire w_dff_A_jNgry8Oy4_2;
	wire w_dff_A_wq4tQ5FZ0_2;
	wire w_dff_B_l9DezJPm0_3;
	wire w_dff_B_WWkWQFP10_3;
	wire w_dff_B_KA9k3SP01_3;
	wire w_dff_B_wrDOKcW35_3;
	wire w_dff_B_5UkqvjVw4_3;
	wire w_dff_B_8DJu24hh8_3;
	wire w_dff_B_i4QGAl8O1_3;
	wire w_dff_B_DbVdrO6Q3_3;
	wire w_dff_B_VTHx8ntN8_3;
	wire w_dff_B_lmQytfA50_3;
	wire w_dff_B_xrTHEsuz2_3;
	wire w_dff_B_EjkoS64Q3_3;
	wire w_dff_B_Db3ZMv005_3;
	wire w_dff_B_dAipauU12_3;
	wire w_dff_B_xj0wtFRl3_3;
	wire w_dff_B_92ZUkadt7_3;
	wire w_dff_B_IbgITdg02_1;
	wire w_dff_B_ZGnttdhf7_1;
	wire w_dff_B_FTnw3Xg31_1;
	wire w_dff_B_LmGYBlcJ0_1;
	wire w_dff_B_hm38KX6z5_1;
	wire w_dff_B_GCOT9CSH3_1;
	wire w_dff_B_RLzrZUL35_1;
	wire w_dff_B_t14rLGUG9_1;
	wire w_dff_B_5ONNJ2aR7_1;
	wire w_dff_B_dFO8mxsd2_1;
	wire w_dff_B_w1bw6mgr0_1;
	wire w_dff_B_BudxxYAP4_0;
	wire w_dff_B_itO9ESq70_0;
	wire w_dff_B_uGzVBG4I4_0;
	wire w_dff_B_Eonx0fjG8_0;
	wire w_dff_B_z7ThNTPj4_0;
	wire w_dff_B_jJaHR3sF9_0;
	wire w_dff_B_87zgBDTl8_0;
	wire w_dff_B_PW4upquJ9_0;
	wire w_dff_B_kEp2i10w6_0;
	wire w_dff_B_cZCIEIF56_0;
	wire w_dff_B_tw1vjor82_0;
	wire w_dff_B_Ad4et2Xi9_0;
	wire w_dff_B_oS7eGAiL7_0;
	wire w_dff_B_CC303Aux6_0;
	wire w_dff_A_43sdw0E60_0;
	wire w_dff_A_b6tgVJP91_0;
	wire w_dff_A_9uWz4vrr6_0;
	wire w_dff_A_38kW0dit4_0;
	wire w_dff_A_VUERVbxm0_0;
	wire w_dff_A_1Xtr9VzC5_0;
	wire w_dff_A_L4eWfhTE0_0;
	wire w_dff_A_6u4U92tJ6_0;
	wire w_dff_A_Xtjrrr5O5_0;
	wire w_dff_A_AhSpaSA57_0;
	wire w_dff_A_cS1gB5A59_0;
	wire w_dff_A_IUbjxoHp6_0;
	wire w_dff_A_h3E7MLZb8_0;
	wire w_dff_A_whmcJS1k6_0;
	wire w_dff_A_hvRrNjYK1_0;
	wire w_dff_B_2X76qvum3_0;
	wire w_dff_B_C3EU4oge3_0;
	wire w_dff_A_Gsyd0ard9_1;
	wire w_dff_A_L6U6GY1b4_1;
	wire w_dff_B_JiY5AdFT7_2;
	wire w_dff_A_VjUM8A8S1_1;
	wire w_dff_A_BAYoBgXK4_1;
	wire w_dff_A_tczWpGTT9_2;
	wire w_dff_A_LGKbteRn7_2;
	wire w_dff_B_rWeVQahk1_3;
	wire w_dff_B_qYuHsMCP9_3;
	wire w_dff_A_JKWe0tgd8_0;
	wire w_dff_A_kPgkeHL59_1;
	wire w_dff_B_UkXvgx952_3;
	wire w_dff_A_9zwH7vGq2_1;
	wire w_dff_A_Y3bjhKXk0_2;
	wire w_dff_B_4fbkGuta1_3;
	wire w_dff_A_OwPFPiKc9_0;
	wire w_dff_A_D38mq5HD8_0;
	wire w_dff_A_lHFT4Hzt1_0;
	wire w_dff_A_IXDKr6J37_1;
	wire w_dff_A_twt0QH2O9_1;
	wire w_dff_A_eQpI6Izx1_1;
	wire w_dff_B_kw3WVZKl4_0;
	wire w_dff_B_dJvBFtKS2_1;
	wire w_dff_B_RWWx8zwf9_0;
	wire w_dff_A_cevCT52N3_1;
	wire w_dff_A_09aFEYq23_0;
	wire w_dff_B_tW00DcSv5_3;
	wire w_dff_A_fp2xXihd8_0;
	wire w_dff_A_35cPAWIb4_0;
	wire w_dff_B_Usf5N05v7_3;
	wire w_dff_A_G8WUL3kv2_0;
	wire w_dff_A_ZGKCYnYR1_0;
	wire w_dff_A_wYupysZH7_2;
	wire w_dff_A_rjUC9ARk0_2;
	wire w_dff_B_QNQfbk5n1_2;
	wire w_dff_A_77YZnQFx6_1;
	wire w_dff_A_EaD5zzkl9_1;
	wire w_dff_A_y4Ea0X3n9_2;
	wire w_dff_A_0mBEjIpT3_2;
	wire w_dff_B_n7nSzbcp3_1;
	wire w_dff_B_vdpK5TU17_1;
	wire w_dff_B_WZEIPPf01_1;
	wire w_dff_B_GZ9zm3sP0_1;
	wire w_dff_B_8YJPDxz80_1;
	wire w_dff_A_y3JAZ3pi5_0;
	wire w_dff_A_Ku2msB4J4_0;
	wire w_dff_A_TKKxVdUJ6_0;
	wire w_dff_A_RjJxRump3_0;
	wire w_dff_A_ntig2NOL4_0;
	wire w_dff_A_EQ0PWSxH9_0;
	wire w_dff_A_Yh7r2zhx9_0;
	wire w_dff_A_6DIvp8LB3_0;
	wire w_dff_A_ZK6n7x4R7_0;
	wire w_dff_A_TZpe6yX65_0;
	wire w_dff_A_tCNaVkta5_0;
	wire w_dff_A_tfIY17mv0_1;
	wire w_dff_B_4HOjDZJ16_3;
	wire w_dff_B_WJSuNHrv7_2;
	wire w_dff_A_cN8fX8Sm1_1;
	wire w_dff_A_uybc2Yyp3_1;
	wire w_dff_A_6VFVOl7i4_2;
	wire w_dff_A_OeuzmHsY5_2;
	wire w_dff_B_KIRixJ3S5_1;
	wire w_dff_B_32uTggt32_1;
	wire w_dff_B_mE7RG9PU7_1;
	wire w_dff_B_5LKhvowI7_1;
	wire w_dff_B_GPN843GF3_1;
	wire w_dff_A_12kEBCe27_0;
	wire w_dff_A_kUCrtOgj9_0;
	wire w_dff_A_fvXBlzga2_0;
	wire w_dff_A_ZxNX1Sgr7_0;
	wire w_dff_A_Y5zLzirL6_0;
	wire w_dff_A_sSbSow6S9_0;
	wire w_dff_A_WYtAyPVj2_0;
	wire w_dff_A_U4AwMOeS9_0;
	wire w_dff_A_iYSgMOEl1_0;
	wire w_dff_A_mpKgBLlT0_0;
	wire w_dff_A_lx7CktvA6_0;
	wire w_dff_A_r5bBon7e8_0;
	wire w_dff_B_10Srcflh0_1;
	wire w_dff_B_FqQKqgp44_1;
	wire w_dff_A_xJEj469K2_1;
	wire w_dff_A_3ZHx4Sfa5_1;
	wire w_dff_A_z3SmD95q2_1;
	wire w_dff_A_V1PZESwJ4_1;
	wire w_dff_A_cDqW9WV37_1;
	wire w_dff_A_Fen5hBPN4_1;
	wire w_dff_A_Dk9wjD6R1_0;
	wire w_dff_A_fb8SYfc44_0;
	wire w_dff_A_oovHH2GY4_0;
	wire w_dff_A_uqCwlZHn5_0;
	wire w_dff_A_bn6iy4Lk7_0;
	wire w_dff_A_s5dsEzNe8_0;
	wire w_dff_A_9LlXIY4a1_0;
	wire w_dff_A_4lE5uAY26_0;
	wire w_dff_A_4nBtkBNO7_0;
	wire w_dff_A_Bpjc5yAZ6_0;
	wire w_dff_A_mJFUkyte8_0;
	wire w_dff_A_7abemTm64_0;
	wire w_dff_B_RPK2d2Xf7_1;
	wire w_dff_B_SNUMfQmR4_1;
	wire w_dff_B_bnwWeJ3A0_1;
	wire w_dff_B_uMxwGq9V4_0;
	wire w_dff_A_2wfAFn5J6_1;
	wire w_dff_A_n8GTCpjy9_1;
	wire w_dff_A_yjmL5mQE3_1;
	wire w_dff_A_iHAj7Unf4_1;
	wire w_dff_A_q5UWtISA6_1;
	wire w_dff_A_P8vhbcLd3_1;
	wire w_dff_B_AsfZNo1y9_3;
	wire w_dff_B_F3v9r44p2_3;
	wire w_dff_A_Gijw0raT3_0;
	wire w_dff_A_AyTXD4nA2_0;
	wire w_dff_A_6OwQNu0J9_0;
	wire w_dff_A_pVs8Nnzn4_1;
	wire w_dff_A_04XLNkTB3_1;
	wire w_dff_A_Z17idjTY7_1;
	wire w_dff_B_gqqmwf5n4_1;
	wire w_dff_A_PkEGoEvi6_0;
	wire w_dff_A_uJhzAsOt0_1;
	wire w_dff_A_aYurxw2I2_1;
	wire w_dff_A_igt5OodG1_1;
	wire w_dff_A_rDsavkC15_1;
	wire w_dff_A_amWPkPxt1_1;
	wire w_dff_A_x3wg5B3h8_1;
	wire w_dff_A_PVbXV4xh1_1;
	wire w_dff_A_3FL4wCib1_1;
	wire w_dff_A_XJhtk5d93_1;
	wire w_dff_A_HgB1EC1h4_1;
	wire w_dff_A_rmgtX48U8_1;
	wire w_dff_A_skdxaJlv5_1;
	wire w_dff_A_sOYhJJgj6_1;
	wire w_dff_A_V62iRMJi4_1;
	wire w_dff_A_883NNCTR0_1;
	wire w_dff_A_8uRKuM9I3_1;
	wire w_dff_A_6XMG2iQb1_1;
	wire w_dff_A_Felw4Quu8_1;
	wire w_dff_A_2ZQnkBe39_1;
	wire w_dff_A_ioZ7jfd93_1;
	wire w_dff_A_OybXhudh7_1;
	wire w_dff_A_QS98rDnB1_1;
	wire w_dff_A_t1Ra9Q1I7_1;
	wire w_dff_A_401pkTmY4_1;
	wire w_dff_A_BdPtsxom3_1;
	wire w_dff_A_d75WGEe48_1;
	wire w_dff_A_GL5TIQ7d7_1;
	wire w_dff_B_aqHRAwgz1_3;
	wire w_dff_B_nVa2DG5s9_1;
	wire w_dff_A_ZalKv5WY2_2;
	wire w_dff_A_1P4uAqKF2_1;
	wire w_dff_A_WuJ6cgDg8_1;
	wire w_dff_A_jeN1wdfO5_2;
	wire w_dff_A_afyGrk4u3_2;
	wire w_dff_A_lWolemKd3_1;
	wire w_dff_A_zDWHIrcy1_1;
	wire w_dff_A_WQXVwCaB7_1;
	wire w_dff_A_syEcHXZs1_1;
	wire w_dff_A_MNtjag3F5_1;
	wire w_dff_A_hOgoEuEd3_1;
	wire w_dff_B_09PlH9TX2_2;
	wire w_dff_B_u4VfuVjA8_2;
	wire w_dff_B_mGhgz6K78_2;
	wire w_dff_B_WBIUpuZz2_2;
	wire w_dff_A_f1Cp3bG98_1;
	wire w_dff_A_tvjJs3Tl8_1;
	wire w_dff_A_4HiJw4826_2;
	wire w_dff_A_oGL2QCwY7_2;
	wire w_dff_A_QbcyzIER2_2;
	wire w_dff_A_KBqT75Wh0_0;
	wire w_dff_A_rAfPXC9K6_0;
	wire w_dff_A_NWX2EhTo2_0;
	wire w_dff_A_LsCdbSGK0_0;
	wire w_dff_A_e2ipIjke8_0;
	wire w_dff_A_yjeGonY34_0;
	wire w_dff_A_ooqiek5u7_0;
	wire w_dff_A_J9Kye0S65_0;
	wire w_dff_A_yWU1yxgg9_0;
	wire w_dff_A_tyPWgfYn3_0;
	wire w_dff_B_qVjn87qS0_1;
	wire w_dff_B_NQdxbq4y2_1;
	wire w_dff_B_9BtTOrGF3_1;
	wire w_dff_B_rV3lDE5L7_0;
	wire w_dff_B_CICOUOZh0_0;
	wire w_dff_B_XDCpQqw55_0;
	wire w_dff_A_rVz5rJYr1_2;
	wire w_dff_A_WkVPWE440_2;
	wire w_dff_A_sCpj0uGB3_2;
	wire w_dff_A_AWIT0A4U3_2;
	wire w_dff_A_D3arNb772_0;
	wire w_dff_A_0bAtBjHV7_0;
	wire w_dff_A_IBtRA15N5_0;
	wire w_dff_A_ooKg5vbG4_0;
	wire w_dff_A_Hcm2yFCB9_0;
	wire w_dff_A_Z03XvnuX8_0;
	wire w_dff_A_zP5OBylv6_0;
	wire w_dff_A_a6DH1R3z8_0;
	wire w_dff_A_QzUmoGbW1_0;
	wire w_dff_A_nXlO4NRF3_2;
	wire w_dff_A_6ggL88hA5_2;
	wire w_dff_A_0haDp6k33_2;
	wire w_dff_A_5pp87aYp3_2;
	wire w_dff_A_kIPf5GNX7_0;
	wire w_dff_B_kt5j7ogb8_3;
	wire w_dff_B_pUvsmUNx6_1;
	wire w_dff_B_hsa6jJmk4_1;
	wire w_dff_B_6090RKg83_1;
	wire w_dff_B_RdqqFmKd0_1;
	wire w_dff_B_vBQYwdZy1_1;
	wire w_dff_A_kn0O4zVs0_0;
	wire w_dff_A_R0blMJvl1_0;
	wire w_dff_A_0LejtOSm4_0;
	wire w_dff_A_3ddvpMdX2_0;
	wire w_dff_A_7zX1W30Z2_0;
	wire w_dff_A_iBWULkw02_0;
	wire w_dff_A_1BSELLl67_0;
	wire w_dff_A_bwzxMwcl3_0;
	wire w_dff_A_xRohhYjS0_0;
	wire w_dff_A_IwGUvFtv0_0;
	wire w_dff_A_XuFJb69N5_0;
	wire w_dff_A_GumpHgl86_0;
	wire w_dff_B_17TASBNk7_1;
	wire w_dff_B_t4FDx38c5_1;
	wire w_dff_B_ai20heMD3_2;
	wire w_dff_A_RCvN3C6T6_0;
	wire w_dff_A_LxU2gbhj5_0;
	wire w_dff_A_NZsG0kcp6_0;
	wire w_dff_A_wRSzDpwI1_0;
	wire w_dff_A_PEN5enCk8_0;
	wire w_dff_A_WcKIGJLU6_0;
	wire w_dff_A_JPnXOuYs9_0;
	wire w_dff_A_djOLakeL8_0;
	wire w_dff_A_zIy1Pbin5_0;
	wire w_dff_A_LqNjbebR4_0;
	wire w_dff_A_QJvkvlbc0_0;
	wire w_dff_A_d4WkHQ0Z2_0;
	wire w_dff_A_hnfjFiB41_2;
	wire w_dff_A_t9pIzLeU2_2;
	wire w_dff_A_VtLDsYHd1_2;
	wire w_dff_A_EKzrDLut8_2;
	wire w_dff_A_vE3DRFNW5_2;
	wire w_dff_A_cvbRW7X30_2;
	wire w_dff_B_qVbzvNhX4_2;
	wire w_dff_B_nFtuYOEF5_2;
	wire w_dff_B_mINt9NCA2_2;
	wire w_dff_A_zJEdtkcf1_0;
	wire w_dff_A_JJm11C8A9_0;
	wire w_dff_A_jeWGtTUG2_0;
	wire w_dff_A_TKvJNnJd2_0;
	wire w_dff_B_DLUqT1wF5_1;
	wire w_dff_A_FzWSr4BD6_0;
	wire w_dff_A_AHUzi0t56_0;
	wire w_dff_A_OUgUnslh1_0;
	wire w_dff_A_SuvM4uh57_0;
	wire w_dff_A_3s6b7g909_1;
	wire w_dff_A_tcZ97Uok8_2;
	wire w_dff_A_KBzpCBu49_1;
	wire w_dff_A_U8XN4OYU1_1;
	wire w_dff_A_GNKRvdAU7_1;
	wire w_dff_B_P7nnRRTv2_1;
	wire w_dff_B_1bk6M5GQ3_1;
	wire w_dff_B_4KWbCSTV9_1;
	wire w_dff_A_Mu8pssWn9_0;
	wire w_dff_A_Pb0nASbk4_0;
	wire w_dff_A_OqHcbhYV9_0;
	wire w_dff_A_5ziUDarr8_0;
	wire w_dff_A_FlESALGf8_0;
	wire w_dff_A_pBpvV1f40_0;
	wire w_dff_A_DFFuUNat0_0;
	wire w_dff_A_gFvpE0dd0_0;
	wire w_dff_A_vtIpbe572_0;
	wire w_dff_A_GUDFpytc8_0;
	wire w_dff_A_b5PWxoNR4_0;
	wire w_dff_A_L7Pb0JD02_0;
	wire w_dff_B_j7ORi5fJ4_1;
	wire w_dff_A_4wDg9vF33_0;
	wire w_dff_A_MXWL5hor6_0;
	wire w_dff_A_aqyJSxiM3_0;
	wire w_dff_A_jtM7ZKzT1_0;
	wire w_dff_A_dsDAIxOa7_0;
	wire w_dff_A_T2qMnk4w4_0;
	wire w_dff_A_TWFGBMQl6_0;
	wire w_dff_A_YZ9X46kS1_0;
	wire w_dff_A_66tUtsGc4_0;
	wire w_dff_A_hdQf4NJJ2_0;
	wire w_dff_A_z1J1XDfe3_0;
	wire w_dff_A_zgT0Dq8h2_0;
	wire w_dff_A_4QPWBgRY3_1;
	wire w_dff_A_CpdIIhVr7_1;
	wire w_dff_B_kmSRrjXT6_2;
	wire w_dff_A_hFLxOAdj0_0;
	wire w_dff_A_If4Cfjzg8_0;
	wire w_dff_A_6bajqFHh2_0;
	wire w_dff_A_hP0iS4SB2_0;
	wire w_dff_A_xluGOmX67_0;
	wire w_dff_A_VysrE9j18_0;
	wire w_dff_A_UwJ20bYM5_0;
	wire w_dff_A_7xs0rADG6_0;
	wire w_dff_A_gE4Z9ugN8_0;
	wire w_dff_A_7pHEecWW5_0;
	wire w_dff_A_ucgiOyXA1_0;
	wire w_dff_A_lzRQ1gWq6_0;
	wire w_dff_A_SKNglHc67_0;
	wire w_dff_B_5vl8XvmS1_1;
	wire w_dff_A_giLq9S0A9_0;
	wire w_dff_A_93JdGNrh0_0;
	wire w_dff_A_MvBygeNP4_0;
	wire w_dff_A_mLDWJFyI4_0;
	wire w_dff_A_VxnPZLMY8_0;
	wire w_dff_A_aivmkRLH2_0;
	wire w_dff_A_rMuGxJE06_0;
	wire w_dff_A_drDFIaqG9_0;
	wire w_dff_A_ZYdwwfIB7_0;
	wire w_dff_A_61NtS2Qr3_0;
	wire w_dff_A_B3U56SD00_0;
	wire w_dff_A_ZGo9KMbm9_0;
	wire w_dff_A_PpbxIOMY5_0;
	wire w_dff_A_giiRDZkl6_0;
	wire w_dff_A_gFO4fKnu8_0;
	wire w_dff_A_yUb77m495_0;
	wire w_dff_A_NoBqEcxZ5_0;
	wire w_dff_A_DKw5nSvP6_0;
	wire w_dff_A_ALrm9nvP8_0;
	wire w_dff_A_aTsbvFUy1_0;
	wire w_dff_A_7bcKgO1E1_0;
	wire w_dff_A_2HBKoYRK1_0;
	wire w_dff_A_dzbJfQrZ0_0;
	wire w_dff_A_VA4WSqGf3_0;
	wire w_dff_A_etYR0HCN8_1;
	wire w_dff_A_vdRpM4MQ1_1;
	wire w_dff_A_FhOJenYV3_1;
	wire w_dff_A_ydhDSGlf7_1;
	wire w_dff_A_sM50eAFw6_1;
	wire w_dff_A_ioKRfuF49_1;
	wire w_dff_A_VJEoO8Ns9_1;
	wire w_dff_A_zhEfnZEw1_1;
	wire w_dff_A_JEDRLKxa8_1;
	wire w_dff_A_AANOPBGj2_1;
	wire w_dff_A_UgnibWgb1_1;
	wire w_dff_A_IlKCEZte2_1;
	wire w_dff_A_wPeWIeJE3_1;
	wire w_dff_A_XM7YifRl2_1;
	wire w_dff_A_A11H96eB5_1;
	wire w_dff_A_CA6hxhaa2_2;
	wire w_dff_A_P1Y0U8u88_1;
	wire w_dff_A_kSXrRche8_1;
	wire w_dff_A_kkskv2WD1_1;
	wire w_dff_A_17WFrIPe7_1;
	wire w_dff_A_BlxwlLW53_1;
	wire w_dff_A_2YhUJvZh6_1;
	wire w_dff_A_IJnM518G8_1;
	wire w_dff_A_cT8yGlSW7_1;
	wire w_dff_A_7MjEoGRb8_1;
	wire w_dff_A_Q12is24H8_1;
	wire w_dff_A_tnAZyTG27_1;
	wire w_dff_A_3Ttm5HXl0_1;
	wire w_dff_A_3mxvC7sV4_1;
	wire w_dff_A_Ox3Ox4Mj2_1;
	wire w_dff_A_tvozGGvU1_1;
	wire w_dff_A_KWzCnMVZ9_1;
	wire w_dff_A_3jrU2D8Q1_1;
	wire w_dff_A_EtFij2pM5_1;
	wire w_dff_A_TqjaJjqP6_1;
	wire w_dff_A_GdEnrtP53_1;
	wire w_dff_A_1EvKxreK4_1;
	wire w_dff_A_sDiT8r3D9_1;
	wire w_dff_A_BiC8QFpX8_1;
	wire w_dff_A_qLKm3xvd3_1;
	wire w_dff_A_xyPaCXtD7_1;
	wire w_dff_A_Q9VlMNWd9_0;
	wire w_dff_A_0U42nwJQ0_0;
	wire w_dff_A_z9OCVGFs0_0;
	wire w_dff_A_3SNReyuh6_0;
	wire w_dff_A_CgzDlYLy2_0;
	wire w_dff_A_eccbc3R32_1;
	wire w_dff_A_XwczMQQv7_1;
	wire w_dff_A_25eBm0iU6_1;
	wire w_dff_A_GJx2WTsJ3_1;
	wire w_dff_A_F3e9q6nE5_1;
	wire w_dff_A_ljeLwGY25_2;
	wire w_dff_A_3HH2s7SH2_2;
	wire w_dff_A_YyFqHaP03_2;
	wire w_dff_A_lBjvXLsJ8_2;
	wire w_dff_A_MXJGJvzN2_2;
	wire w_dff_A_EzFCGtMC6_2;
	wire w_dff_A_1ct4tUVW5_2;
	wire w_dff_A_tDjuBF022_1;
	wire w_dff_A_TFlHmIqk2_0;
	wire w_dff_A_VoHE9fBq5_0;
	wire w_dff_A_e2jJr84u4_0;
	wire w_dff_A_vlfJkYt84_0;
	wire w_dff_A_psgFL68B2_0;
	wire w_dff_A_Y50veSqC4_0;
	wire w_dff_A_khJMROJi4_0;
	wire w_dff_A_7TayJBC28_0;
	wire w_dff_A_PgsX1UY79_0;
	wire w_dff_A_xwdIUY8b6_0;
	wire w_dff_A_wVPmatmG8_0;
	wire w_dff_A_ARU548hm1_0;
	wire w_dff_A_lu4iJZYK4_0;
	wire w_dff_A_C9fp8HEz8_0;
	wire w_dff_A_YPuRu8le4_0;
	wire w_dff_A_bB8PgO1H0_0;
	wire w_dff_A_6VQt6JLB0_0;
	wire w_dff_A_Ar2fbf4V7_0;
	wire w_dff_A_x0V1XLR20_0;
	wire w_dff_A_vGm6oouJ3_0;
	wire w_dff_A_zBiBCKun6_0;
	wire w_dff_A_pF8VoppL0_0;
	wire w_dff_A_AO545wsb5_0;
	wire w_dff_A_ReU8cIDJ8_0;
	wire w_dff_A_Tesifn7c3_1;
	wire w_dff_A_r5dHI0Mg5_1;
	wire w_dff_A_JaSSlB4U1_1;
	wire w_dff_A_01mEqRT91_1;
	wire w_dff_A_ep9tyags2_1;
	wire w_dff_A_c1QAZGLK1_1;
	wire w_dff_A_OsTznZ9H0_1;
	wire w_dff_A_GxhoUOcO6_1;
	wire w_dff_A_g1tDK9Uz9_1;
	wire w_dff_A_Lrt6JbTI1_1;
	wire w_dff_A_oXWUJnBQ8_1;
	wire w_dff_A_LvjoHDe40_1;
	wire w_dff_A_rP6NhMxu7_1;
	wire w_dff_A_nISm5J6t7_1;
	wire w_dff_A_4NxQWxMU5_1;
	wire w_dff_A_7YHlHYqo4_2;
	wire w_dff_A_c5zEmjNo8_2;
	wire w_dff_A_hxMpqtlg4_2;
	wire w_dff_A_E0DfOccd9_2;
	wire w_dff_A_BNiJlq0L4_2;
	wire w_dff_A_IOydEwTp7_2;
	wire w_dff_A_4wOHPwQ55_2;
	wire w_dff_A_V9BDueEv6_2;
	wire w_dff_A_4E1MKIdp5_2;
	wire w_dff_A_p6r6U7192_2;
	wire w_dff_A_YT0iPKEZ2_2;
	wire w_dff_A_uE5DdWu64_2;
	wire w_dff_A_lR96zMAH0_2;
	wire w_dff_A_2C4bJCot3_2;
	wire w_dff_A_aMzM9twT2_2;
	wire w_dff_A_hgRE24Ur4_1;
	wire w_dff_A_zDn1sl8B6_0;
	wire w_dff_A_Pl2UOARS7_0;
	wire w_dff_A_UcdiNOaL2_0;
	wire w_dff_A_L49YtfNm5_0;
	wire w_dff_A_YAKN5FWX1_0;
	wire w_dff_A_AIRXoOpO8_0;
	wire w_dff_A_BidEmMFn2_0;
	wire w_dff_A_NnIqgKkW5_0;
	wire w_dff_A_d0cJmlpv2_0;
	wire w_dff_A_AhXpHyez9_0;
	wire w_dff_A_t1gICSgz1_0;
	wire w_dff_A_MzGgJx775_2;
	wire w_dff_B_CNYfRje88_3;
	wire w_dff_A_dTNbfKqW2_1;
	wire w_dff_A_gySoFXbb7_0;
	wire w_dff_A_IzVn4X9S1_0;
	wire w_dff_A_a52UWG9N9_0;
	wire w_dff_A_ciRUgfln5_0;
	wire w_dff_A_0DQUmZFa0_0;
	wire w_dff_A_aL6OIHWs4_0;
	wire w_dff_A_cM89K7PN7_0;
	wire w_dff_A_bOgEq25R1_0;
	wire w_dff_A_QpA6hHJu8_0;
	wire w_dff_A_IyxPokaL6_0;
	wire w_dff_A_FWNJJz255_0;
	wire w_dff_A_JRMPtdzP8_0;
	wire w_dff_A_Jwv0xFl69_0;
	wire w_dff_A_Jrv4KkjY5_0;
	wire w_dff_A_hbsWC19E6_0;
	wire w_dff_A_nxKKuqmQ3_0;
	wire w_dff_A_5VAfND6l6_0;
	wire w_dff_A_PLCzIBgv4_0;
	wire w_dff_A_HnUe3F6y4_0;
	wire w_dff_A_nV6Otq3z1_0;
	wire w_dff_A_NqwXV67n3_0;
	wire w_dff_A_3wy2t2RS7_0;
	wire w_dff_A_vhvZQKxB3_0;
	wire w_dff_A_Q0lthbmY7_0;
	wire w_dff_A_W3bMojaO0_0;
	wire w_dff_A_xdonyWUW5_0;
	wire w_dff_A_5QXqa2PP2_0;
	wire w_dff_A_pLD4ERRR2_0;
	wire w_dff_A_g0l0pkBX9_0;
	wire w_dff_A_qpxDMKE01_0;
	wire w_dff_A_eYjeBoBV6_0;
	wire w_dff_A_I9y0xZiD0_0;
	wire w_dff_A_o0A0cI0X7_0;
	wire w_dff_A_xP5ed0Si7_0;
	wire w_dff_A_kpEjZ3k20_0;
	wire w_dff_A_qClEJX0E5_0;
	wire w_dff_B_0QcSUpE87_1;
	wire w_dff_A_OxbtqQiH3_0;
	wire w_dff_A_i5KrNt6T9_0;
	wire w_dff_A_yd3QNXME2_0;
	wire w_dff_A_acZ5Ytfb4_0;
	wire w_dff_A_cfTIUGSJ8_0;
	wire w_dff_A_JQrdEivi1_0;
	wire w_dff_A_QfZHXklO8_0;
	wire w_dff_A_o8Hxctjp1_0;
	wire w_dff_A_NH9undmQ0_0;
	wire w_dff_A_CNXFDjFT6_0;
	wire w_dff_A_UuCND0Wo4_0;
	wire w_dff_A_g4VM4Dvy0_0;
	wire w_dff_A_3DLO0SEv4_1;
	wire w_dff_A_KO2VCb6W2_1;
	wire w_dff_A_lUd35UYF5_1;
	wire w_dff_A_2ge8XyT67_1;
	wire w_dff_A_ZasxbszV9_1;
	wire w_dff_A_YL5btN9k8_1;
	wire w_dff_A_ausLFpKq4_1;
	wire w_dff_A_5KnuFEmd1_1;
	wire w_dff_A_xC3uKHfr6_1;
	wire w_dff_A_AKH3bdFV4_1;
	wire w_dff_A_sRTDwoK12_1;
	wire w_dff_A_ztNSLy4P5_1;
	wire w_dff_A_8uYIgGTS0_2;
	wire w_dff_A_UCIhReKV0_0;
	wire w_dff_A_pfVDzSTE0_1;
	wire w_dff_A_KgRkFrKY7_1;
	wire w_dff_A_kACUpb8O4_1;
	wire w_dff_A_AlS9pvZO9_1;
	wire w_dff_A_o6MO40ph5_1;
	wire w_dff_A_J2Q4ckKZ9_1;
	wire w_dff_A_UP4Oqxzk7_1;
	wire w_dff_A_MjJSgreQ2_1;
	wire w_dff_A_6UXBdWxc1_1;
	wire w_dff_A_zLLi7gXj2_1;
	wire w_dff_A_tfxBaH2f5_1;
	wire w_dff_A_NlFA4YzQ5_1;
	wire w_dff_A_RpMR2OxI7_1;
	wire w_dff_A_Aq2G3hRS3_0;
	wire w_dff_A_6sZriiSp8_0;
	wire w_dff_A_rBmApmgP5_0;
	wire w_dff_A_G4M8TZ2k6_0;
	wire w_dff_A_RFjz22497_0;
	wire w_dff_A_QCdRjKSu9_0;
	wire w_dff_A_5HrEIJzf6_0;
	wire w_dff_A_ZDdsL0xS4_0;
	wire w_dff_A_WLj5kph79_0;
	wire w_dff_A_DHFxyEwJ4_0;
	wire w_dff_A_cEYVCbYt4_0;
	wire w_dff_A_JyaBcpWa8_0;
	wire w_dff_A_Hcb55XUz0_0;
	wire w_dff_A_fq6alYdv7_0;
	wire w_dff_A_36Lp5GWA1_0;
	wire w_dff_A_RKopOPX02_0;
	wire w_dff_A_6PoYq1Wu0_0;
	wire w_dff_A_DVrloNLw8_0;
	wire w_dff_A_BwvDfDsI4_0;
	wire w_dff_A_qmWValbh4_0;
	wire w_dff_A_2H4Zhj1s8_0;
	wire w_dff_A_sbStELCV0_0;
	wire w_dff_A_YHUWyG7E9_0;
	wire w_dff_A_GtIiwpDE5_2;
	wire w_dff_A_W5ZQRB9x1_2;
	wire w_dff_B_GaHf3EBN6_3;
	wire w_dff_A_vGQfHwSI9_0;
	wire w_dff_A_xh7XY4I17_0;
	wire w_dff_A_VKKvjeLx6_0;
	wire w_dff_A_mjDFR3ZZ8_0;
	wire w_dff_A_cyVzZvfH3_0;
	wire w_dff_A_zvJDWPJX1_0;
	wire w_dff_A_rxR4Nddt3_0;
	wire w_dff_A_0nqpbG9k7_0;
	wire w_dff_A_7awu9U0n2_0;
	wire w_dff_A_dUMHazyn4_0;
	wire w_dff_A_j4u8WWwp4_0;
	wire w_dff_A_UfGRfBbx1_0;
	wire w_dff_A_YB2zu5zl1_2;
	wire w_dff_A_cdqCJLBY5_0;
	wire w_dff_A_PSCRMpSH3_0;
	wire w_dff_A_ZkCaUY862_0;
	wire w_dff_A_oBQTgxkS7_0;
	wire w_dff_A_BpVIvNa50_0;
	wire w_dff_A_mv8Apsd28_0;
	wire w_dff_A_pQ4XnbpO5_2;
	wire w_dff_A_S1ieWPyR5_0;
	wire w_dff_A_mOxFe7am8_0;
	wire w_dff_A_PvAxLKaP0_0;
	wire w_dff_A_uCKgvjuD2_0;
	wire w_dff_A_VsNLXOon8_0;
	wire w_dff_A_BeQV5WJi1_0;
	wire w_dff_A_ysQrHSkC2_2;
	wire w_dff_A_vN9CF0Gm8_0;
	wire w_dff_A_we0ql9Mr0_0;
	wire w_dff_A_Vwjcf8eh8_0;
	wire w_dff_A_1FVjeGYk7_0;
	wire w_dff_A_qYRMynfE0_0;
	wire w_dff_A_cZzKFklK0_0;
	wire w_dff_A_HmEPIFW31_2;
	wire w_dff_A_Yf84sPaq2_0;
	wire w_dff_A_xBjcXoJg3_0;
	wire w_dff_A_IUAawD926_0;
	wire w_dff_A_6ruDch8Q0_0;
	wire w_dff_A_fhOyMIsJ9_0;
	wire w_dff_A_IqqEoIAE2_0;
	wire w_dff_A_p6TGz3CQ7_2;
	wire w_dff_A_pcP2slpG1_0;
	wire w_dff_A_nLrVGHj24_0;
	wire w_dff_A_zDjIKNEK5_0;
	wire w_dff_A_ul1jI3C58_0;
	wire w_dff_A_4TF89CR94_0;
	wire w_dff_A_fZXszqZF7_0;
	wire w_dff_A_PXMQJc3d5_2;
	wire w_dff_A_2N3PY2Gp7_0;
	wire w_dff_A_MWnd850Z8_0;
	wire w_dff_A_q7w0t8Tn7_0;
	wire w_dff_A_4GBe8whH4_0;
	wire w_dff_A_9lS6el8A2_0;
	wire w_dff_A_rfva3CpZ6_0;
	wire w_dff_A_qNoSiuRR7_2;
	wire w_dff_A_v4RRjfoh9_0;
	wire w_dff_A_AoCrHRVr9_0;
	wire w_dff_A_1t0T9EDO3_0;
	wire w_dff_A_rT5XSn3U7_0;
	wire w_dff_A_2M8lKHt31_0;
	wire w_dff_A_Mtg6WqcU7_0;
	wire w_dff_A_39k7m2jl2_2;
	wire w_dff_A_7qsHetyr7_0;
	wire w_dff_A_Hwsv1vYt5_0;
	wire w_dff_A_hQTMbLAk3_0;
	wire w_dff_A_QBRE3wef0_0;
	wire w_dff_A_xgVmC8PK6_0;
	wire w_dff_A_bzv9FnAW3_0;
	wire w_dff_A_BLmIZlKE0_2;
	wire w_dff_A_i6juiczR6_0;
	wire w_dff_A_b8S6KonW0_0;
	wire w_dff_A_Ft2Yyr073_0;
	wire w_dff_A_mZTqoN8o6_0;
	wire w_dff_A_GXEhLkSL5_0;
	wire w_dff_A_FT3qtJPI0_0;
	wire w_dff_A_gNVWv1vW4_2;
	wire w_dff_A_sATPXdvY4_0;
	wire w_dff_A_F6qhPc3x8_0;
	wire w_dff_A_JQaKlUJk6_0;
	wire w_dff_A_uP6PnsRX4_0;
	wire w_dff_A_R4POdEhI4_0;
	wire w_dff_A_VJzf25z71_0;
	wire w_dff_A_2UJqkRKI1_2;
	wire w_dff_A_wfNajdZh6_0;
	wire w_dff_A_B7VUIsVW0_0;
	wire w_dff_A_wbhkfoiN6_0;
	wire w_dff_A_Ivbg4XuS0_0;
	wire w_dff_A_xYY1WJmk6_0;
	wire w_dff_A_4s4oRm1t2_0;
	wire w_dff_A_C3HB9a9M2_2;
	wire w_dff_A_W2j5GYVz1_0;
	wire w_dff_A_UoJPwRW47_0;
	wire w_dff_A_JEpQsdg96_0;
	wire w_dff_A_ixsuCzqR1_0;
	wire w_dff_A_pBSzkd7J0_0;
	wire w_dff_A_Kej9aHSI0_0;
	wire w_dff_A_m9hGZyC60_2;
	wire w_dff_A_ptNbcEFu4_0;
	wire w_dff_A_6mNYGtf30_0;
	wire w_dff_A_dQ51EN3j7_0;
	wire w_dff_A_q31Gen692_0;
	wire w_dff_A_VktOMNAv9_0;
	wire w_dff_A_P0wzao6F5_0;
	wire w_dff_A_l5uqOluA3_2;
	wire w_dff_A_f2h19v173_0;
	wire w_dff_A_z1MIvZhV2_0;
	wire w_dff_A_UKhPafOI0_0;
	wire w_dff_A_HGATsIzh4_0;
	wire w_dff_A_hZTYuz462_0;
	wire w_dff_A_wTV7cp5M7_0;
	wire w_dff_A_Q79VKY0V0_2;
	wire w_dff_A_zDAUhiBr7_0;
	wire w_dff_A_oOpvw8D26_0;
	wire w_dff_A_v0gXjNc76_0;
	wire w_dff_A_6VRRScJ37_0;
	wire w_dff_A_AxSq91kA5_0;
	wire w_dff_A_rRkmF9Gm9_0;
	wire w_dff_A_cx8NO26b9_2;
	wire w_dff_A_U1k4ksCe2_0;
	wire w_dff_A_AZVTyJzx7_0;
	wire w_dff_A_0HA9kgHt9_0;
	wire w_dff_A_VfTg2vxP4_0;
	wire w_dff_A_yEuuE7940_0;
	wire w_dff_A_lcECBcc08_0;
	wire w_dff_A_QcEcVxwy4_2;
	wire w_dff_A_hSV2AnXX1_2;
	wire w_dff_A_hZdDs68H3_2;
	wire w_dff_A_NAhYsgVu5_0;
	jnot g000(.din(w_G146_0[2]),.dout(n58),.clk(gclk));
	jxor g001(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n59),.clk(gclk));
	jxor g002(.dina(w_n59_0[1]),.dinb(n58),.dout(n60),.clk(gclk));
	jnot g003(.din(w_G953_1[2]),.dout(n61),.clk(gclk));
	jand g004(.dina(w_n61_3[2]),.dinb(w_G234_0[2]),.dout(n62),.clk(gclk));
	jand g005(.dina(w_n62_0[1]),.dinb(w_G221_0[1]),.dout(n63),.clk(gclk));
	jxor g006(.dina(n63),.dinb(w_G137_0[2]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_G128_1[1]),.dinb(w_G119_0[2]),.dout(n65),.clk(gclk));
	jxor g008(.dina(w_dff_B_XDCpQqw55_0),.dinb(n64),.dout(n66),.clk(gclk));
	jxor g009(.dina(n66),.dinb(w_G110_1[1]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_n67_0[1]),.dinb(w_n60_0[2]),.dout(n68),.clk(gclk));
	jor g011(.dina(w_n68_0[1]),.dinb(w_G902_3[2]),.dout(n69),.clk(gclk));
	jnot g012(.din(w_G902_3[1]),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_3[1]),.dinb(w_G234_0[1]),.dout(n71),.clk(gclk));
	jnot g014(.din(w_n71_0[1]),.dout(n72),.clk(gclk));
	jand g015(.dina(n72),.dinb(w_G217_0[2]),.dout(n73),.clk(gclk));
	jxor g016(.dina(w_n73_0[1]),.dinb(n69),.dout(n74),.clk(gclk));
	jnot g017(.din(w_G134_0[2]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_G137_0[1]),.dinb(n75),.dout(n76),.clk(gclk));
	jnot g019(.din(w_G131_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_G146_0[1]),.dinb(w_G143_1[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(n78),.dinb(w_G128_1[0]),.dout(n79),.clk(gclk));
	jxor g022(.dina(w_n79_0[1]),.dinb(w_n77_0[1]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_dff_B_0QcSUpE87_1),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[1]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(w_n82_0[1]),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_1[1]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[2]),.dinb(w_n70_3[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(n91),.dinb(w_G472_0[1]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[2]),.dinb(w_n74_1[1]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[0]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_0[2]),.dout(n96),.clk(gclk));
	jand g039(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n97),.clk(gclk));
	jnot g040(.din(w_G110_1[0]),.dout(n98),.clk(gclk));
	jxor g041(.dina(w_G122_1[1]),.dinb(n98),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n100),.clk(gclk));
	jxor g043(.dina(n100),.dinb(w_G101_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_n101_0[1]),.dinb(w_n84_0[0]),.dout(n102),.clk(gclk));
	jxor g045(.dina(n102),.dinb(w_dff_B_5vl8XvmS1_1),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n61_3[1]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n79_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(w_dff_B_j7ORi5fJ4_1),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n103_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[2]),.dinb(w_n70_2[2]),.dout(n108),.clk(gclk));
	jxor g051(.dina(w_n108_0[1]),.dinb(w_n97_0[1]),.dout(n109),.clk(gclk));
	jand g052(.dina(w_n109_0[1]),.dinb(w_n96_0[2]),.dout(n110),.clk(gclk));
	jnot g053(.din(w_G221_0[0]),.dout(n111),.clk(gclk));
	jor g054(.dina(w_n71_0[0]),.dinb(w_dff_B_DLUqT1wF5_1),.dout(n112),.clk(gclk));
	jxor g055(.dina(w_G140_0[1]),.dinb(w_G110_0[2]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n61_3[0]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(n114),.dinb(w_n101_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(w_dff_B_t4FDx38c5_1),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n81_0[1]),.dout(n117),.clk(gclk));
	jand g060(.dina(w_n117_0[2]),.dinb(w_n70_2[1]),.dout(n118),.clk(gclk));
	jxor g061(.dina(w_n118_0[1]),.dinb(w_G469_0[2]),.dout(n119),.clk(gclk));
	jand g062(.dina(w_n119_0[1]),.dinb(w_n112_1[1]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n110_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_1[1]),.dinb(w_n93_0[2]),.dout(n122),.clk(gclk));
	jnot g065(.din(w_G478_0[2]),.dout(n123),.clk(gclk));
	jxor g066(.dina(w_G143_1[0]),.dinb(w_G128_0[2]),.dout(n124),.clk(gclk));
	jand g067(.dina(w_n62_0[0]),.dinb(w_G217_0[1]),.dout(n125),.clk(gclk));
	jxor g068(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n126),.clk(gclk));
	jxor g069(.dina(w_G134_0[1]),.dinb(w_G107_0[1]),.dout(n127),.clk(gclk));
	jxor g070(.dina(n127),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g071(.dina(w_dff_B_uMxwGq9V4_0),.dinb(n125),.dout(n129),.clk(gclk));
	jxor g072(.dina(n129),.dinb(w_dff_B_bnwWeJ3A0_1),.dout(n130),.clk(gclk));
	jand g073(.dina(w_n130_0[2]),.dinb(w_n70_2[0]),.dout(n131),.clk(gclk));
	jxor g074(.dina(w_n131_0[1]),.dinb(w_dff_B_8YJPDxz80_1),.dout(n132),.clk(gclk));
	jnot g075(.din(w_G475_0[2]),.dout(n133),.clk(gclk));
	jxor g076(.dina(w_G143_0[2]),.dinb(w_n77_0[0]),.dout(n134),.clk(gclk));
	jxor g077(.dina(w_G122_0[2]),.dinb(w_n82_0[0]),.dout(n135),.clk(gclk));
	jxor g078(.dina(n135),.dinb(w_G104_0[1]),.dout(n136),.clk(gclk));
	jnot g079(.din(w_G214_0[0]),.dout(n137),.clk(gclk));
	jor g080(.dina(w_n86_0[0]),.dinb(n137),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(w_n60_0[1]),.dout(n139),.clk(gclk));
	jxor g082(.dina(n139),.dinb(n136),.dout(n140),.clk(gclk));
	jxor g083(.dina(n140),.dinb(w_dff_B_FqQKqgp44_1),.dout(n141),.clk(gclk));
	jand g084(.dina(w_n141_0[2]),.dinb(w_n70_1[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_n142_0[1]),.dinb(w_dff_B_GPN843GF3_1),.dout(n143),.clk(gclk));
	jand g086(.dina(w_n143_1[1]),.dinb(w_n132_0[2]),.dout(n144),.clk(gclk));
	jor g087(.dina(w_n61_2[2]),.dinb(w_dff_B_nVa2DG5s9_1),.dout(n145),.clk(gclk));
	jand g088(.dina(w_G237_0[0]),.dinb(w_G234_0[0]),.dout(n146),.clk(gclk));
	jor g089(.dina(w_n146_0[1]),.dinb(w_n70_1[1]),.dout(n147),.clk(gclk));
	jor g090(.dina(w_n147_0[1]),.dinb(w_n145_0[1]),.dout(n148),.clk(gclk));
	jnot g091(.din(w_n146_0[0]),.dout(n149),.clk(gclk));
	jand g092(.dina(w_n61_2[1]),.dinb(w_G952_0[2]),.dout(n150),.clk(gclk));
	jand g093(.dina(n150),.dinb(n149),.dout(n151),.clk(gclk));
	jnot g094(.din(w_n151_0[2]),.dout(n152),.clk(gclk));
	jand g095(.dina(w_n152_0[1]),.dinb(w_dff_B_gqqmwf5n4_1),.dout(n153),.clk(gclk));
	jnot g096(.din(w_n153_0[2]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n144_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[2]),.dinb(w_n122_0[1]),.dout(n156),.clk(gclk));
	jxor g099(.dina(w_n156_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_YB2zu5zl1_2),.clk(gclk));
	jnot g100(.din(w_n92_1[1]),.dout(n158),.clk(gclk));
	jand g101(.dina(w_n158_1[1]),.dinb(w_n74_1[0]),.dout(n159),.clk(gclk));
	jand g102(.dina(w_n159_1[1]),.dinb(w_n121_1[0]),.dout(n160),.clk(gclk));
	jxor g103(.dina(w_n142_0[0]),.dinb(w_G475_0[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_0[2]),.dinb(w_n132_0[1]),.dout(n162),.clk(gclk));
	jand g105(.dina(w_n162_0[1]),.dinb(w_n154_1[0]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_0[2]),.dinb(w_n160_0[1]),.dout(n164),.clk(gclk));
	jxor g107(.dina(w_n164_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_pQ4XnbpO5_2),.clk(gclk));
	jxor g108(.dina(w_n131_0[0]),.dinb(w_G478_0[1]),.dout(n166),.clk(gclk));
	jand g109(.dina(w_n143_1[0]),.dinb(w_n166_1[1]),.dout(n167),.clk(gclk));
	jand g110(.dina(w_n167_0[1]),.dinb(w_n154_0[2]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n168_0[2]),.dinb(w_n160_0[0]),.dout(n169),.clk(gclk));
	jxor g112(.dina(w_n169_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_ysQrHSkC2_2),.clk(gclk));
	jnot g113(.din(w_n60_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n67_0[0]),.dinb(w_dff_B_9BtTOrGF3_1),.dout(n172),.clk(gclk));
	jand g115(.dina(w_n172_0[1]),.dinb(w_n70_1[0]),.dout(n173),.clk(gclk));
	jxor g116(.dina(w_n73_0[0]),.dinb(n173),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n158_1[0]),.dinb(w_n174_1[1]),.dout(n175),.clk(gclk));
	jand g118(.dina(w_n175_0[1]),.dinb(w_n155_0[1]),.dout(n176),.clk(gclk));
	jand g119(.dina(n176),.dinb(w_n121_0[2]),.dout(n177),.clk(gclk));
	jxor g120(.dina(w_n177_0[1]),.dinb(w_G110_0[1]),.dout(w_dff_A_HmEPIFW31_2),.clk(gclk));
	jand g121(.dina(w_n92_1[0]),.dinb(w_n174_1[0]),.dout(n179),.clk(gclk));
	jand g122(.dina(w_n179_0[2]),.dinb(w_n121_0[1]),.dout(n180),.clk(gclk));
	jor g123(.dina(w_n61_2[0]),.dinb(w_dff_B_dJvBFtKS2_1),.dout(n181),.clk(gclk));
	jor g124(.dina(w_n181_0[2]),.dinb(w_n147_0[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(w_dff_B_kw3WVZKl4_0),.dinb(w_n152_0[0]),.dout(n183),.clk(gclk));
	jnot g126(.din(w_n183_0[2]),.dout(n184),.clk(gclk));
	jand g127(.dina(w_n184_1[1]),.dinb(w_n167_0[0]),.dout(n185),.clk(gclk));
	jand g128(.dina(w_n185_0[2]),.dinb(w_n180_0[1]),.dout(n186),.clk(gclk));
	jxor g129(.dina(w_n186_0[1]),.dinb(w_G128_0[1]),.dout(w_dff_A_p6TGz3CQ7_2),.clk(gclk));
	jand g130(.dina(w_n161_0[1]),.dinb(w_n166_1[0]),.dout(n188),.clk(gclk));
	jand g131(.dina(w_n188_0[2]),.dinb(w_n184_1[0]),.dout(n189),.clk(gclk));
	jand g132(.dina(w_n189_0[1]),.dinb(w_n122_0[0]),.dout(n190),.clk(gclk));
	jxor g133(.dina(w_n190_0[1]),.dinb(w_G143_0[1]),.dout(w_dff_A_PXMQJc3d5_2),.clk(gclk));
	jand g134(.dina(w_n184_0[2]),.dinb(w_n162_0[0]),.dout(n192),.clk(gclk));
	jand g135(.dina(w_n192_0[2]),.dinb(w_n180_0[0]),.dout(n193),.clk(gclk));
	jxor g136(.dina(w_n193_0[1]),.dinb(w_G146_0[0]),.dout(w_dff_A_qNoSiuRR7_2),.clk(gclk));
	jnot g137(.din(w_G469_0[1]),.dout(n195),.clk(gclk));
	jxor g138(.dina(w_n118_0[0]),.dinb(w_dff_B_vBQYwdZy1_1),.dout(n196),.clk(gclk));
	jand g139(.dina(w_n196_0[2]),.dinb(w_n112_1[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n110_0[1]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_1[1]),.dinb(w_n93_0[1]),.dout(n199),.clk(gclk));
	jand g142(.dina(w_n199_0[1]),.dinb(w_n163_0[1]),.dout(n200),.clk(gclk));
	jxor g143(.dina(w_n200_0[1]),.dinb(w_G113_0[0]),.dout(w_dff_A_39k7m2jl2_2),.clk(gclk));
	jand g144(.dina(w_n199_0[0]),.dinb(w_n168_0[1]),.dout(n202),.clk(gclk));
	jxor g145(.dina(w_n202_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_BLmIZlKE0_2),.clk(gclk));
	jand g146(.dina(w_n198_1[0]),.dinb(w_n179_0[1]),.dout(n204),.clk(gclk));
	jand g147(.dina(n204),.dinb(w_n155_0[0]),.dout(n205),.clk(gclk));
	jxor g148(.dina(w_n205_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_gNVWv1vW4_2),.clk(gclk));
	jand g149(.dina(w_n197_1[0]),.dinb(w_n159_1[0]),.dout(n207),.clk(gclk));
	jand g150(.dina(w_n154_0[1]),.dinb(w_n110_0[0]),.dout(n208),.clk(gclk));
	jand g151(.dina(n208),.dinb(w_n188_0[1]),.dout(n209),.clk(gclk));
	jand g152(.dina(w_dff_B_mFbBRedQ8_0),.dinb(w_n207_0[1]),.dout(n210),.clk(gclk));
	jxor g153(.dina(w_n210_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_2UJqkRKI1_2),.clk(gclk));
	jand g154(.dina(w_n192_0[1]),.dinb(w_n175_0[0]),.dout(n212),.clk(gclk));
	jand g155(.dina(w_n212_0[1]),.dinb(w_n198_0[2]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_n213_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_C3HB9a9M2_2),.clk(gclk));
	jnot g157(.din(w_n97_0[0]),.dout(n215),.clk(gclk));
	jxor g158(.dina(w_n108_0[0]),.dinb(w_dff_B_4KWbCSTV9_1),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_0[2]),.dinb(w_n96_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[2]),.dinb(w_n120_0[0]),.dout(n218),.clk(gclk));
	jand g161(.dina(w_n218_1[1]),.dinb(w_n93_0[0]),.dout(n219),.clk(gclk));
	jand g162(.dina(w_n219_0[1]),.dinb(w_n192_0[0]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_m9hGZyC60_2),.clk(gclk));
	jand g164(.dina(w_n219_0[0]),.dinb(w_n185_0[1]),.dout(n222),.clk(gclk));
	jxor g165(.dina(w_n222_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_l5uqOluA3_2),.clk(gclk));
	jand g166(.dina(w_n184_0[1]),.dinb(w_n144_1[1]),.dout(n224),.clk(gclk));
	jand g167(.dina(w_dff_B_h0UcXPex1_0),.dinb(w_n179_0[0]),.dout(n225),.clk(gclk));
	jand g168(.dina(n225),.dinb(w_n218_1[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_Q79VKY0V0_2),.clk(gclk));
	jand g170(.dina(w_n218_0[2]),.dinb(w_n212_0[0]),.dout(n228),.clk(gclk));
	jxor g171(.dina(w_n228_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_cx8NO26b9_2),.clk(gclk));
	jor g172(.dina(w_n177_0[0]),.dinb(w_n169_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n202_0[0]),.dinb(w_n164_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(n230),.dout(n232),.clk(gclk));
	jor g175(.dina(w_n205_0[0]),.dinb(w_n156_0[0]),.dout(n233),.clk(gclk));
	jor g176(.dina(w_n210_0[0]),.dinb(w_n200_0[0]),.dout(n234),.clk(gclk));
	jor g177(.dina(n234),.dinb(n233),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(n232),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n193_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n222_0[0]),.dinb(w_n186_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jor g182(.dina(w_n228_0[0]),.dinb(w_n190_0[0]),.dout(n240),.clk(gclk));
	jor g183(.dina(w_n226_0[0]),.dinb(w_n213_0[0]),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n240),.dout(n242),.clk(gclk));
	jor g185(.dina(n242),.dinb(n239),.dout(n243),.clk(gclk));
	jor g186(.dina(n243),.dinb(n236),.dout(n244),.clk(gclk));
	jor g187(.dina(w_n218_0[1]),.dinb(w_n198_0[1]),.dout(n245),.clk(gclk));
	jand g188(.dina(n245),.dinb(w_n144_1[0]),.dout(n246),.clk(gclk));
	jand g189(.dina(w_n217_0[1]),.dinb(w_n197_0[2]),.dout(n247),.clk(gclk));
	jxor g190(.dina(w_n143_0[2]),.dinb(w_n132_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(w_dff_B_vfSLBcRq1_0),.dinb(n247),.dout(n249),.clk(gclk));
	jor g192(.dina(w_dff_B_piq5rTZj4_0),.dinb(n246),.dout(n250),.clk(gclk));
	jand g193(.dina(n250),.dinb(w_n159_0[2]),.dout(n251),.clk(gclk));
	jand g194(.dina(w_n217_0[0]),.dinb(w_n144_0[2]),.dout(n252),.clk(gclk));
	jor g195(.dina(w_n92_0[2]),.dinb(w_n174_0[2]),.dout(n253),.clk(gclk));
	jor g196(.dina(w_n158_0[2]),.dinb(w_n74_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(w_n197_0[1]),.dinb(w_n254_1[1]),.dout(n255),.clk(gclk));
	jand g198(.dina(n255),.dinb(w_n253_0[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_n252_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(n257),.dinb(n251),.dout(n258),.clk(gclk));
	jand g201(.dina(n258),.dinb(w_n151_0[1]),.dout(n259),.clk(gclk));
	jxor g202(.dina(w_n112_0[2]),.dinb(w_n96_0[0]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n151_0[0]),.dout(n261),.clk(gclk));
	jand g204(.dina(w_dff_B_mgpfL50U4_0),.dinb(w_n196_0[1]),.dout(n262),.clk(gclk));
	jand g205(.dina(n262),.dinb(w_n216_0[1]),.dout(n263),.clk(gclk));
	jand g206(.dina(w_n159_0[1]),.dinb(w_n144_0[1]),.dout(n264),.clk(gclk));
	jand g207(.dina(n264),.dinb(w_dff_B_UiVPnDn26_1),.dout(n265),.clk(gclk));
	jor g208(.dina(w_dff_B_ni4xBugN4_0),.dinb(n259),.dout(n266),.clk(gclk));
	jor g209(.dina(n266),.dinb(w_n244_2[2]),.dout(n267),.clk(gclk));
	jand g210(.dina(n267),.dinb(w_G952_0[1]),.dout(n268),.clk(gclk));
	jand g211(.dina(w_n252_0[0]),.dinb(w_n207_0[0]),.dout(n269),.clk(gclk));
	jor g212(.dina(n269),.dinb(w_G953_1[0]),.dout(n270),.clk(gclk));
	jor g213(.dina(w_dff_B_nGg3Q8VT6_0),.dinb(n268),.dout(w_dff_A_QcEcVxwy4_2),.clk(gclk));
	jnot g214(.din(w_n107_0[1]),.dout(n272),.clk(gclk));
	jor g215(.dina(w_n216_0[0]),.dinb(w_n95_0[1]),.dout(n273),.clk(gclk));
	jnot g216(.din(w_n112_0[1]),.dout(n274),.clk(gclk));
	jor g217(.dina(w_n196_0[0]),.dinb(w_n274_0[1]),.dout(n275),.clk(gclk));
	jor g218(.dina(w_n275_0[1]),.dinb(w_n273_0[2]),.dout(n276),.clk(gclk));
	jor g219(.dina(w_n253_0[1]),.dinb(w_n276_1[1]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n168_0[0]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n278_0[1]),.dinb(w_n277_0[1]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n161_0[0]),.dinb(w_n166_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n153_0[1]),.dinb(w_n280_0[1]),.dout(n281),.clk(gclk));
	jor g224(.dina(w_n92_0[1]),.dinb(w_n74_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_0[1]),.dinb(w_n281_0[2]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n276_1[0]),.dout(n284),.clk(gclk));
	jand g227(.dina(n284),.dinb(n279),.dout(n285),.clk(gclk));
	jnot g228(.din(w_n163_0[0]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n277_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n158_0[1]),.dinb(w_n174_0[1]),.dout(n288),.clk(gclk));
	jor g231(.dina(w_n119_0[0]),.dinb(w_n274_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(w_n289_0[1]),.dinb(w_n273_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n290_0[2]),.dinb(w_n288_0[2]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n291_0[1]),.dinb(w_n278_0[0]),.dout(n292),.clk(gclk));
	jand g235(.dina(n292),.dinb(n287),.dout(n293),.clk(gclk));
	jand g236(.dina(n293),.dinb(n285),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n276_0[2]),.dinb(w_n288_0[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n281_0[1]),.dinb(w_n295_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(w_n290_0[1]),.dinb(w_n254_1[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(n297),.dinb(w_n281_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n296),.dout(n299),.clk(gclk));
	jor g242(.dina(w_n291_0[0]),.dinb(w_n286_0[0]),.dout(n300),.clk(gclk));
	jor g243(.dina(w_n289_0[0]),.dinb(w_n253_0[0]),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n188_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n153_0[0]),.dinb(w_n273_0[0]),.dout(n303),.clk(gclk));
	jor g246(.dina(n303),.dinb(n302),.dout(n304),.clk(gclk));
	jor g247(.dina(w_dff_B_RWWx8zwf9_0),.dinb(n301),.dout(n305),.clk(gclk));
	jand g248(.dina(n305),.dinb(n300),.dout(n306),.clk(gclk));
	jand g249(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jand g250(.dina(n307),.dinb(n294),.dout(n308),.clk(gclk));
	jor g251(.dina(w_n254_0[2]),.dinb(w_n276_0[1]),.dout(n309),.clk(gclk));
	jor g252(.dina(w_n143_0[1]),.dinb(w_n166_0[1]),.dout(n310),.clk(gclk));
	jor g253(.dina(w_n183_0[1]),.dinb(n310),.dout(n311),.clk(gclk));
	jor g254(.dina(w_n311_0[2]),.dinb(w_n309_0[1]),.dout(n312),.clk(gclk));
	jor g255(.dina(w_n109_0[0]),.dinb(w_n95_0[0]),.dout(n313),.clk(gclk));
	jor g256(.dina(n313),.dinb(w_n275_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n314_0[2]),.dinb(w_n288_0[0]),.dout(n315),.clk(gclk));
	jor g258(.dina(w_n315_0[1]),.dinb(w_n311_0[1]),.dout(n316),.clk(gclk));
	jand g259(.dina(n316),.dinb(n312),.dout(n317),.clk(gclk));
	jnot g260(.din(w_n185_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(w_n318_0[1]),.dinb(w_n309_0[0]),.dout(n319),.clk(gclk));
	jor g262(.dina(w_n315_0[0]),.dinb(w_n318_0[0]),.dout(n320),.clk(gclk));
	jand g263(.dina(n320),.dinb(n319),.dout(n321),.clk(gclk));
	jand g264(.dina(n321),.dinb(n317),.dout(n322),.clk(gclk));
	jnot g265(.din(w_n189_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(w_dff_B_C3EU4oge3_0),.dinb(w_n295_0[0]),.dout(n324),.clk(gclk));
	jor g267(.dina(w_n311_0[0]),.dinb(w_n282_0[0]),.dout(n325),.clk(gclk));
	jor g268(.dina(w_n314_0[1]),.dinb(w_n325_0[1]),.dout(n326),.clk(gclk));
	jand g269(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n325_0[0]),.dinb(w_n290_0[0]),.dout(n328),.clk(gclk));
	jor g271(.dina(w_n183_0[0]),.dinb(w_n280_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(w_dff_B_2X76qvum3_0),.dinb(w_n254_0[1]),.dout(n330),.clk(gclk));
	jor g273(.dina(n330),.dinb(w_n314_0[0]),.dout(n331),.clk(gclk));
	jand g274(.dina(n331),.dinb(n328),.dout(n332),.clk(gclk));
	jand g275(.dina(n332),.dinb(n327),.dout(n333),.clk(gclk));
	jand g276(.dina(n333),.dinb(n322),.dout(n334),.clk(gclk));
	jand g277(.dina(w_n334_0[1]),.dinb(w_n308_0[1]),.dout(n335),.clk(gclk));
	jand g278(.dina(w_G902_2[2]),.dinb(w_G210_0[0]),.dout(n336),.clk(gclk));
	jnot g279(.din(w_n336_0[1]),.dout(n337),.clk(gclk));
	jor g280(.dina(w_dff_B_HuwMTHLf4_0),.dinb(w_n335_2[1]),.dout(n338),.clk(gclk));
	jor g281(.dina(n338),.dinb(w_dff_B_1ENNgSjZ1_1),.dout(n339),.clk(gclk));
	jor g282(.dina(w_n61_1[2]),.dinb(w_G952_0[0]),.dout(n340),.clk(gclk));
	jand g283(.dina(w_n336_0[0]),.dinb(w_n244_2[1]),.dout(n341),.clk(gclk));
	jor g284(.dina(n341),.dinb(w_n107_0[0]),.dout(n342),.clk(gclk));
	jand g285(.dina(n342),.dinb(w_n340_2[1]),.dout(n343),.clk(gclk));
	jand g286(.dina(n343),.dinb(w_dff_B_1psTim966_1),.dout(G51),.clk(gclk));
	jnot g287(.din(w_n117_0[1]),.dout(n345),.clk(gclk));
	jand g288(.dina(w_G902_2[1]),.dinb(w_G469_0[0]),.dout(n346),.clk(gclk));
	jnot g289(.din(w_n346_0[1]),.dout(n347),.clk(gclk));
	jor g290(.dina(w_dff_B_x8rUjeRO8_0),.dinb(w_n335_2[0]),.dout(n348),.clk(gclk));
	jor g291(.dina(n348),.dinb(w_dff_B_9Nqzcnkn1_1),.dout(n349),.clk(gclk));
	jand g292(.dina(w_n346_0[0]),.dinb(w_n244_2[0]),.dout(n350),.clk(gclk));
	jor g293(.dina(n350),.dinb(w_n117_0[0]),.dout(n351),.clk(gclk));
	jand g294(.dina(n351),.dinb(w_n340_2[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_dff_B_g2OF9prz8_1),.dout(G54),.clk(gclk));
	jnot g296(.din(w_n141_0[1]),.dout(n354),.clk(gclk));
	jand g297(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n355),.clk(gclk));
	jnot g298(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jor g299(.dina(w_dff_B_pgBGJOFz1_0),.dinb(w_n335_1[2]),.dout(n357),.clk(gclk));
	jor g300(.dina(n357),.dinb(w_dff_B_asEVOhQ28_1),.dout(n358),.clk(gclk));
	jand g301(.dina(w_n355_0[0]),.dinb(w_n244_1[2]),.dout(n359),.clk(gclk));
	jor g302(.dina(n359),.dinb(w_n141_0[0]),.dout(n360),.clk(gclk));
	jand g303(.dina(n360),.dinb(w_n340_1[2]),.dout(n361),.clk(gclk));
	jand g304(.dina(n361),.dinb(w_dff_B_2zSnQfFs1_1),.dout(G60),.clk(gclk));
	jnot g305(.din(w_n130_0[1]),.dout(n363),.clk(gclk));
	jand g306(.dina(w_G902_1[2]),.dinb(w_G478_0[0]),.dout(n364),.clk(gclk));
	jnot g307(.din(w_n364_0[1]),.dout(n365),.clk(gclk));
	jor g308(.dina(w_dff_B_QxqH7i8L4_0),.dinb(w_n335_1[1]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(w_dff_B_7HXfiGRz1_1),.dout(n367),.clk(gclk));
	jand g310(.dina(w_n364_0[0]),.dinb(w_n244_1[1]),.dout(n368),.clk(gclk));
	jor g311(.dina(n368),.dinb(w_n130_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(n369),.dinb(w_n340_1[1]),.dout(n370),.clk(gclk));
	jand g313(.dina(n370),.dinb(w_dff_B_wmO4A6qe3_1),.dout(G63),.clk(gclk));
	jand g314(.dina(w_G902_1[1]),.dinb(w_G217_0[0]),.dout(n372),.clk(gclk));
	jand g315(.dina(w_n372_0[1]),.dinb(w_n244_1[0]),.dout(n373),.clk(gclk));
	jor g316(.dina(n373),.dinb(w_n172_0[0]),.dout(n374),.clk(gclk));
	jnot g317(.din(w_n372_0[0]),.dout(n375),.clk(gclk));
	jor g318(.dina(w_dff_B_oWeEm77E3_0),.dinb(w_n335_1[0]),.dout(n376),.clk(gclk));
	jor g319(.dina(n376),.dinb(w_n68_0[0]),.dout(n377),.clk(gclk));
	jand g320(.dina(n377),.dinb(w_n340_1[0]),.dout(n378),.clk(gclk));
	jand g321(.dina(n378),.dinb(w_dff_B_Z1UoXxNG6_1),.dout(G66),.clk(gclk));
	jnot g322(.din(w_n145_0[0]),.dout(n380),.clk(gclk));
	jor g323(.dina(w_n308_0[0]),.dinb(w_G953_0[2]),.dout(n381),.clk(gclk));
	jor g324(.dina(w_n61_1[1]),.dinb(w_G224_0[0]),.dout(n382),.clk(gclk));
	jand g325(.dina(w_dff_B_GsXdjJPE0_0),.dinb(n381),.dout(n383),.clk(gclk));
	jxor g326(.dina(n383),.dinb(w_n103_0[0]),.dout(n384),.clk(gclk));
	jor g327(.dina(n384),.dinb(w_dff_B_TEb94CHB0_1),.dout(w_dff_A_hSV2AnXX1_2),.clk(gclk));
	jor g328(.dina(w_n334_0[0]),.dinb(w_G953_0[1]),.dout(n386),.clk(gclk));
	jor g329(.dina(w_n61_1[0]),.dinb(w_G227_0[0]),.dout(n387),.clk(gclk));
	jand g330(.dina(n387),.dinb(w_n181_0[1]),.dout(n388),.clk(gclk));
	jand g331(.dina(w_dff_B_PeeA8JVj0_0),.dinb(n386),.dout(n389),.clk(gclk));
	jnot g332(.din(w_n181_0[0]),.dout(n390),.clk(gclk));
	jxor g333(.dina(w_n81_0[0]),.dinb(w_n59_0[0]),.dout(n391),.clk(gclk));
	jor g334(.dina(n391),.dinb(w_dff_B_6PMUkzqF5_1),.dout(n392),.clk(gclk));
	jxor g335(.dina(w_dff_B_3ezn6Tq90_0),.dinb(n389),.dout(w_dff_A_hZdDs68H3_2),.clk(gclk));
	jnot g336(.din(w_n90_0[1]),.dout(n394),.clk(gclk));
	jand g337(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n395),.clk(gclk));
	jnot g338(.din(w_n395_0[1]),.dout(n396),.clk(gclk));
	jor g339(.dina(w_dff_B_CC303Aux6_0),.dinb(w_n335_0[2]),.dout(n397),.clk(gclk));
	jor g340(.dina(n397),.dinb(w_dff_B_w1bw6mgr0_1),.dout(n398),.clk(gclk));
	jand g341(.dina(w_n395_0[0]),.dinb(w_n244_0[2]),.dout(n399),.clk(gclk));
	jor g342(.dina(n399),.dinb(w_n90_0[0]),.dout(n400),.clk(gclk));
	jand g343(.dina(n400),.dinb(w_n340_0[2]),.dout(n401),.clk(gclk));
	jand g344(.dina(n401),.dinb(w_dff_B_HjcMotW98_1),.dout(G57),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_t1gICSgz1_0),.doutb(w_G101_0[1]),.doutc(w_dff_A_MzGgJx775_2),.din(w_dff_B_CNYfRje88_3));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_VA4WSqGf3_0),.doutb(w_dff_A_vdRpM4MQ1_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_ZGo9KMbm9_0),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_G110_0[0]),.doutb(w_dff_A_3jrU2D8Q1_1),.doutc(w_G110_0[2]),.din(G110));
	jspl jspl_w_G110_1(.douta(w_G110_1[0]),.doutb(w_dff_A_BlxwlLW53_1),.din(w_G110_0[0]));
	jspl jspl_w_G113_0(.douta(w_dff_A_qClEJX0E5_0),.doutb(w_G113_0[1]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_Q0lthbmY7_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_JRMPtdzP8_0),.doutb(w_G119_0[1]),.doutc(w_G119_0[2]),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_A11H96eB5_1),.doutc(w_dff_A_CA6hxhaa2_2),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_dff_A_FhOJenYV3_1),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_zgT0Dq8h2_0),.doutb(w_dff_A_CpdIIhVr7_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_dff_A_NlFA4YzQ5_1),.doutc(w_G128_0[2]),.din(G128));
	jspl jspl_w_G128_1(.douta(w_dff_A_UCIhReKV0_0),.doutb(w_G128_1[1]),.din(w_G128_0[0]));
	jspl jspl_w_G131_0(.douta(w_dff_A_JyaBcpWa8_0),.doutb(w_G131_0[1]),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_UfGRfBbx1_0),.doutb(w_G134_0[1]),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_YHUWyG7E9_0),.doutb(w_G137_0[1]),.doutc(w_dff_A_W5ZQRB9x1_2),.din(w_dff_B_GaHf3EBN6_3));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_d4WkHQ0Z2_0),.doutb(w_G140_0[1]),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_dff_A_ztNSLy4P5_1),.doutc(w_dff_A_8uYIgGTS0_2),.din(G143));
	jspl jspl_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.din(w_G143_0[0]));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_g4VM4Dvy0_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(G146));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_dff_A_hgRE24Ur4_1),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_dff_A_tDjuBF022_1),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_G217_0[0]),.doutb(w_dff_A_tvjJs3Tl8_1),.doutc(w_dff_A_QbcyzIER2_2),.din(G217));
	jspl jspl_w_G221_0(.douta(w_G221_0[0]),.doutb(w_dff_A_U8XN4OYU1_1),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_G224_0[1]),.din(w_dff_B_kmSRrjXT6_2));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_G227_0[1]),.din(w_dff_B_ai20heMD3_2));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_dff_A_3s6b7g909_1),.doutc(w_dff_A_tcZ97Uok8_2),.din(G234));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_G469_0[0]),.doutb(w_G469_0[1]),.doutc(w_dff_A_cvbRW7X30_2),.din(G469));
	jspl jspl_w_G472_0(.douta(w_G472_0[0]),.doutb(w_dff_A_hOgoEuEd3_1),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_Fen5hBPN4_1),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_G478_0[0]),.doutb(w_dff_A_P8vhbcLd3_1),.doutc(w_G478_0[2]),.din(G478));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_G902_1[1]),.doutc(w_G902_1[2]),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_G902_2[1]),.doutc(w_G902_2[2]),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_G902_3[0]),.doutb(w_G902_3[1]),.doutc(w_dff_A_1ct4tUVW5_2),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_dff_A_GL5TIQ7d7_1),.doutc(w_G952_0[2]),.din(w_dff_B_aqHRAwgz1_3));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_dff_A_4NxQWxMU5_1),.doutc(w_dff_A_aMzM9twT2_2),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_ReU8cIDJ8_0),.doutb(w_G953_1[1]),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_n59_0(.douta(w_dff_A_IBtRA15N5_0),.doutb(w_n59_0[1]),.din(n59));
	jspl3 jspl3_w_n60_0(.douta(w_n60_0[0]),.doutb(w_n60_0[1]),.doutc(w_dff_A_AWIT0A4U3_2),.din(n60));
	jspl3 jspl3_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.doutc(w_n61_0[2]),.din(n61));
	jspl3 jspl3_w_n61_1(.douta(w_n61_1[0]),.doutb(w_n61_1[1]),.doutc(w_n61_1[2]),.din(w_n61_0[0]));
	jspl3 jspl3_w_n61_2(.douta(w_n61_2[0]),.doutb(w_n61_2[1]),.doutc(w_n61_2[2]),.din(w_n61_0[1]));
	jspl3 jspl3_w_n61_3(.douta(w_n61_3[0]),.doutb(w_n61_3[1]),.doutc(w_n61_3[2]),.din(w_n61_0[2]));
	jspl jspl_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n68_0(.douta(w_dff_A_TZpe6yX65_0),.doutb(w_n68_0[1]),.din(n68));
	jspl3 jspl3_w_n70_0(.douta(w_n70_0[0]),.doutb(w_dff_A_1EvKxreK4_1),.doutc(w_n70_0[2]),.din(n70));
	jspl3 jspl3_w_n70_1(.douta(w_dff_A_QzUmoGbW1_0),.doutb(w_n70_1[1]),.doutc(w_dff_A_5pp87aYp3_2),.din(w_n70_0[0]));
	jspl3 jspl3_w_n70_2(.douta(w_n70_2[0]),.doutb(w_n70_2[1]),.doutc(w_n70_2[2]),.din(w_n70_0[1]));
	jspl jspl_w_n70_3(.douta(w_dff_A_SuvM4uh57_0),.doutb(w_n70_3[1]),.din(w_n70_0[2]));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(w_dff_B_WBIUpuZz2_2));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_dff_A_RpMR2OxI7_1),.din(n77));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl jspl_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_dTNbfKqW2_1),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n90_0(.douta(w_dff_A_ARU548hm1_0),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_dff_A_WuJ6cgDg8_1),.doutc(w_dff_A_afyGrk4u3_2),.din(n92));
	jspl3 jspl3_w_n92_1(.douta(w_dff_A_ZGKCYnYR1_0),.doutb(w_n92_1[1]),.doutc(w_dff_A_rjUC9ARk0_2),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_dff_A_CgzDlYLy2_0),.doutb(w_dff_A_F3e9q6nE5_1),.doutc(w_n95_0[2]),.din(n95));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_ArFhudP54_1),.doutc(w_dff_A_wq4tQ5FZ0_2),.din(n96));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_dff_A_xyPaCXtD7_1),.din(n97));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_dff_A_SKNglHc67_0),.doutb(w_n103_0[1]),.din(n103));
	jspl3 jspl3_w_n107_0(.douta(w_dff_A_L7Pb0JD02_0),.doutb(w_n107_0[1]),.doutc(w_n107_0[2]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.doutc(w_n110_0[2]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_TKvJNnJd2_0),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_dff_A_GumpHgl86_0),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_dff_A_0CYnpiTc0_2),.din(w_dff_B_Vs822WDe7_3));
	jspl jspl_w_n121_1(.douta(w_n121_1[0]),.doutb(w_n121_1[1]),.din(w_n121_0[0]));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_7abemTm64_0),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n141_0(.douta(w_dff_A_r5bBon7e8_0),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl jspl_w_n143_1(.douta(w_n143_1[0]),.doutb(w_n143_1[1]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_dff_A_2KEevYyh8_1),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_dff_A_4Gp49ERV3_0),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl3 jspl3_w_n151_0(.douta(w_dff_A_PkEGoEvi6_0),.doutb(w_dff_A_rmgtX48U8_1),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_dff_A_6OwQNu0J9_0),.doutb(w_dff_A_Z17idjTY7_1),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(w_dff_B_F3v9r44p2_3));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_dff_A_ppa3Ic6i2_0),.doutb(w_n155_0[1]),.doutc(w_dff_A_BItCi9uA1_2),.din(w_dff_B_UBOMW93A9_3));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.doutc(w_n158_0[2]),.din(w_dff_B_Usf5N05v7_3));
	jspl jspl_w_n158_1(.douta(w_n158_1[0]),.doutb(w_n158_1[1]),.din(w_n158_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_dff_A_MLI46m0M2_2),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_dff_A_EaD5zzkl9_1),.doutc(w_dff_A_0mBEjIpT3_2),.din(n163));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl jspl_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.din(w_n166_0[0]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_dff_A_uybc2Yyp3_1),.doutc(w_dff_A_OeuzmHsY5_2),.din(n168));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n172_0(.douta(w_dff_A_tyPWgfYn3_0),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.doutc(w_n174_0[2]),.din(n174));
	jspl jspl_w_n174_1(.douta(w_n174_1[0]),.doutb(w_n174_1[1]),.din(w_n174_0[0]));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.doutc(w_n179_0[2]),.din(n179));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n183_0(.douta(w_dff_A_lHFT4Hzt1_0),.doutb(w_dff_A_eQpI6Izx1_1),.doutc(w_n183_0[2]),.din(n183));
	jspl3 jspl3_w_n184_0(.douta(w_n184_0[0]),.doutb(w_n184_0[1]),.doutc(w_n184_0[2]),.din(w_dff_B_qYuHsMCP9_3));
	jspl jspl_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_dff_A_BAYoBgXK4_1),.doutc(w_dff_A_LGKbteRn7_2),.din(n185));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl3 jspl3_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_cevCT52N3_1),.doutc(w_n188_0[2]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_dff_A_L6U6GY1b4_1),.din(n189));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_dff_A_NQaIJkRP2_0),.doutb(w_n192_0[1]),.doutc(w_dff_A_8q8lNVYD4_2),.din(w_dff_B_i6lhBmlg3_3));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl3 jspl3_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(n196));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_dff_A_H7gxCzUt6_1),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_dff_A_hiMHTam68_0),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_dff_A_zDeAIA3f6_0),.doutb(w_n198_0[1]),.doutc(w_dff_A_HaA4EzaU8_2),.din(n198));
	jspl jspl_w_n198_1(.douta(w_n198_1[0]),.doutb(w_n198_1[1]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_dff_A_GNKRvdAU7_1),.doutc(w_n216_0[2]),.din(n216));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl3 jspl3_w_n218_0(.douta(w_dff_A_IHqyDOlI7_0),.doutb(w_n218_0[1]),.doutc(w_dff_A_LORqUJdb7_2),.din(n218));
	jspl jspl_w_n218_1(.douta(w_dff_A_9ps5Vm5Q7_0),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl3 jspl3_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.doutc(w_n244_0[2]),.din(n244));
	jspl3 jspl3_w_n244_1(.douta(w_n244_1[0]),.doutb(w_n244_1[1]),.doutc(w_n244_1[2]),.din(w_n244_0[0]));
	jspl3 jspl3_w_n244_2(.douta(w_n244_2[0]),.doutb(w_n244_2[1]),.doutc(w_n244_2[2]),.din(w_n244_0[1]));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_XRjJXcUI0_1),.din(w_dff_B_f3bEe1Gh2_2));
	jspl3 jspl3_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.doutc(w_dff_A_ZalKv5WY2_2),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_mINt9NCA2_2));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_n276_0[2]),.din(w_dff_B_kt5j7ogb8_3));
	jspl jspl_w_n276_1(.douta(w_dff_A_kIPf5GNX7_0),.doutb(w_n276_1[1]),.din(w_n276_0[0]));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(w_dff_B_WJSuNHrv7_2));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n281_0(.douta(w_dff_A_tCNaVkta5_0),.doutb(w_dff_A_tfIY17mv0_1),.doutc(w_n281_0[2]),.din(w_dff_B_4HOjDZJ16_3));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(w_dff_B_QNQfbk5n1_2));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n289_0(.douta(w_dff_A_35cPAWIb4_0),.doutb(w_n289_0[1]),.din(n289));
	jspl3 jspl3_w_n290_0(.douta(w_dff_A_09aFEYq23_0),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(w_dff_B_tW00DcSv5_3));
	jspl jspl_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.din(n291));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_dff_A_9zwH7vGq2_1),.doutc(w_dff_A_Y3bjhKXk0_2),.din(w_dff_B_4fbkGuta1_3));
	jspl3 jspl3_w_n314_0(.douta(w_dff_A_JKWe0tgd8_0),.doutb(w_dff_A_kPgkeHL59_1),.doutc(w_n314_0[2]),.din(w_dff_B_UkXvgx952_3));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(w_dff_B_JiY5AdFT7_2));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.doutc(w_n335_1[2]),.din(w_n335_0[0]));
	jspl jspl_w_n335_2(.douta(w_n335_2[0]),.doutb(w_n335_2[1]),.din(w_n335_0[1]));
	jspl jspl_w_n336_0(.douta(w_dff_A_Z2vaiXFp1_0),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.doutc(w_n340_0[2]),.din(w_dff_B_92ZUkadt7_3));
	jspl3 jspl3_w_n340_1(.douta(w_n340_1[0]),.doutb(w_n340_1[1]),.doutc(w_n340_1[2]),.din(w_n340_0[0]));
	jspl jspl_w_n340_2(.douta(w_n340_2[0]),.doutb(w_n340_2[1]),.din(w_n340_0[1]));
	jspl jspl_w_n346_0(.douta(w_dff_A_R35ciefN3_0),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n355_0(.douta(w_dff_A_LrjQo2z18_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n364_0(.douta(w_dff_A_g4DgAnzk9_0),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_cfi4m6ds0_1),.din(n372));
	jspl jspl_w_n395_0(.douta(w_dff_A_hvRrNjYK1_0),.doutb(w_n395_0[1]),.din(n395));
	jdff dff_B_6Tj43yLD7_0(.din(n270),.dout(w_dff_B_6Tj43yLD7_0),.clk(gclk));
	jdff dff_B_bkhnxK0n9_0(.din(w_dff_B_6Tj43yLD7_0),.dout(w_dff_B_bkhnxK0n9_0),.clk(gclk));
	jdff dff_B_mEmd24zc6_0(.din(w_dff_B_bkhnxK0n9_0),.dout(w_dff_B_mEmd24zc6_0),.clk(gclk));
	jdff dff_B_aohSYRY50_0(.din(w_dff_B_mEmd24zc6_0),.dout(w_dff_B_aohSYRY50_0),.clk(gclk));
	jdff dff_B_nGg3Q8VT6_0(.din(w_dff_B_aohSYRY50_0),.dout(w_dff_B_nGg3Q8VT6_0),.clk(gclk));
	jdff dff_B_KYoJ6tCB8_0(.din(n265),.dout(w_dff_B_KYoJ6tCB8_0),.clk(gclk));
	jdff dff_B_Lg0smOrj5_0(.din(w_dff_B_KYoJ6tCB8_0),.dout(w_dff_B_Lg0smOrj5_0),.clk(gclk));
	jdff dff_B_ni4xBugN4_0(.din(w_dff_B_Lg0smOrj5_0),.dout(w_dff_B_ni4xBugN4_0),.clk(gclk));
	jdff dff_B_Y771JsgA5_1(.din(n263),.dout(w_dff_B_Y771JsgA5_1),.clk(gclk));
	jdff dff_B_UiVPnDn26_1(.din(w_dff_B_Y771JsgA5_1),.dout(w_dff_B_UiVPnDn26_1),.clk(gclk));
	jdff dff_B_8aigdvcU2_0(.din(n261),.dout(w_dff_B_8aigdvcU2_0),.clk(gclk));
	jdff dff_B_mgpfL50U4_0(.din(w_dff_B_8aigdvcU2_0),.dout(w_dff_B_mgpfL50U4_0),.clk(gclk));
	jdff dff_A_XRjJXcUI0_1(.dout(w_n252_0[1]),.din(w_dff_A_XRjJXcUI0_1),.clk(gclk));
	jdff dff_B_oMDeVr7b5_2(.din(n252),.dout(w_dff_B_oMDeVr7b5_2),.clk(gclk));
	jdff dff_B_f3bEe1Gh2_2(.din(w_dff_B_oMDeVr7b5_2),.dout(w_dff_B_f3bEe1Gh2_2),.clk(gclk));
	jdff dff_B_piq5rTZj4_0(.din(n249),.dout(w_dff_B_piq5rTZj4_0),.clk(gclk));
	jdff dff_B_vfSLBcRq1_0(.din(n248),.dout(w_dff_B_vfSLBcRq1_0),.clk(gclk));
	jdff dff_B_1psTim966_1(.din(n339),.dout(w_dff_B_1psTim966_1),.clk(gclk));
	jdff dff_B_fiJZxm4Z8_1(.din(n272),.dout(w_dff_B_fiJZxm4Z8_1),.clk(gclk));
	jdff dff_B_keQD9Y6l7_1(.din(w_dff_B_fiJZxm4Z8_1),.dout(w_dff_B_keQD9Y6l7_1),.clk(gclk));
	jdff dff_B_YCEUnVpZ7_1(.din(w_dff_B_keQD9Y6l7_1),.dout(w_dff_B_YCEUnVpZ7_1),.clk(gclk));
	jdff dff_B_mD4x9hcs7_1(.din(w_dff_B_YCEUnVpZ7_1),.dout(w_dff_B_mD4x9hcs7_1),.clk(gclk));
	jdff dff_B_dBMhKthn9_1(.din(w_dff_B_mD4x9hcs7_1),.dout(w_dff_B_dBMhKthn9_1),.clk(gclk));
	jdff dff_B_GS8B36zJ7_1(.din(w_dff_B_dBMhKthn9_1),.dout(w_dff_B_GS8B36zJ7_1),.clk(gclk));
	jdff dff_B_k1OSsfpz5_1(.din(w_dff_B_GS8B36zJ7_1),.dout(w_dff_B_k1OSsfpz5_1),.clk(gclk));
	jdff dff_B_c0cDSTjj5_1(.din(w_dff_B_k1OSsfpz5_1),.dout(w_dff_B_c0cDSTjj5_1),.clk(gclk));
	jdff dff_B_Wze0wzyd2_1(.din(w_dff_B_c0cDSTjj5_1),.dout(w_dff_B_Wze0wzyd2_1),.clk(gclk));
	jdff dff_B_rEFRVGKw1_1(.din(w_dff_B_Wze0wzyd2_1),.dout(w_dff_B_rEFRVGKw1_1),.clk(gclk));
	jdff dff_B_1ENNgSjZ1_1(.din(w_dff_B_rEFRVGKw1_1),.dout(w_dff_B_1ENNgSjZ1_1),.clk(gclk));
	jdff dff_B_r8UYE5iT4_0(.din(n337),.dout(w_dff_B_r8UYE5iT4_0),.clk(gclk));
	jdff dff_B_5ETLHI0A6_0(.din(w_dff_B_r8UYE5iT4_0),.dout(w_dff_B_5ETLHI0A6_0),.clk(gclk));
	jdff dff_B_dUZCs7jr5_0(.din(w_dff_B_5ETLHI0A6_0),.dout(w_dff_B_dUZCs7jr5_0),.clk(gclk));
	jdff dff_B_AKSEso6s7_0(.din(w_dff_B_dUZCs7jr5_0),.dout(w_dff_B_AKSEso6s7_0),.clk(gclk));
	jdff dff_B_DFzpmXxf4_0(.din(w_dff_B_AKSEso6s7_0),.dout(w_dff_B_DFzpmXxf4_0),.clk(gclk));
	jdff dff_B_SsbS50495_0(.din(w_dff_B_DFzpmXxf4_0),.dout(w_dff_B_SsbS50495_0),.clk(gclk));
	jdff dff_B_0NZxvEWX1_0(.din(w_dff_B_SsbS50495_0),.dout(w_dff_B_0NZxvEWX1_0),.clk(gclk));
	jdff dff_B_2jxfQ34O3_0(.din(w_dff_B_0NZxvEWX1_0),.dout(w_dff_B_2jxfQ34O3_0),.clk(gclk));
	jdff dff_B_jEKe9zsj7_0(.din(w_dff_B_2jxfQ34O3_0),.dout(w_dff_B_jEKe9zsj7_0),.clk(gclk));
	jdff dff_B_deEBEmzQ3_0(.din(w_dff_B_jEKe9zsj7_0),.dout(w_dff_B_deEBEmzQ3_0),.clk(gclk));
	jdff dff_B_AR45nFuG8_0(.din(w_dff_B_deEBEmzQ3_0),.dout(w_dff_B_AR45nFuG8_0),.clk(gclk));
	jdff dff_B_3E35odDm8_0(.din(w_dff_B_AR45nFuG8_0),.dout(w_dff_B_3E35odDm8_0),.clk(gclk));
	jdff dff_B_JOhpdqEq1_0(.din(w_dff_B_3E35odDm8_0),.dout(w_dff_B_JOhpdqEq1_0),.clk(gclk));
	jdff dff_B_HuwMTHLf4_0(.din(w_dff_B_JOhpdqEq1_0),.dout(w_dff_B_HuwMTHLf4_0),.clk(gclk));
	jdff dff_A_xXznSd8I7_0(.dout(w_n336_0[0]),.din(w_dff_A_xXznSd8I7_0),.clk(gclk));
	jdff dff_A_6OrMfaJ90_0(.dout(w_dff_A_xXznSd8I7_0),.din(w_dff_A_6OrMfaJ90_0),.clk(gclk));
	jdff dff_A_YmAvIMiq7_0(.dout(w_dff_A_6OrMfaJ90_0),.din(w_dff_A_YmAvIMiq7_0),.clk(gclk));
	jdff dff_A_t5Bh1HlL3_0(.dout(w_dff_A_YmAvIMiq7_0),.din(w_dff_A_t5Bh1HlL3_0),.clk(gclk));
	jdff dff_A_PgDBrITs1_0(.dout(w_dff_A_t5Bh1HlL3_0),.din(w_dff_A_PgDBrITs1_0),.clk(gclk));
	jdff dff_A_Rzc3NOqW3_0(.dout(w_dff_A_PgDBrITs1_0),.din(w_dff_A_Rzc3NOqW3_0),.clk(gclk));
	jdff dff_A_c5pUAJpm7_0(.dout(w_dff_A_Rzc3NOqW3_0),.din(w_dff_A_c5pUAJpm7_0),.clk(gclk));
	jdff dff_A_DhkEh3MU5_0(.dout(w_dff_A_c5pUAJpm7_0),.din(w_dff_A_DhkEh3MU5_0),.clk(gclk));
	jdff dff_A_hkU1notJ6_0(.dout(w_dff_A_DhkEh3MU5_0),.din(w_dff_A_hkU1notJ6_0),.clk(gclk));
	jdff dff_A_KgHCMNRE3_0(.dout(w_dff_A_hkU1notJ6_0),.din(w_dff_A_KgHCMNRE3_0),.clk(gclk));
	jdff dff_A_Bkj0KmFw3_0(.dout(w_dff_A_KgHCMNRE3_0),.din(w_dff_A_Bkj0KmFw3_0),.clk(gclk));
	jdff dff_A_LJaleAfG1_0(.dout(w_dff_A_Bkj0KmFw3_0),.din(w_dff_A_LJaleAfG1_0),.clk(gclk));
	jdff dff_A_xV6AHXxs7_0(.dout(w_dff_A_LJaleAfG1_0),.din(w_dff_A_xV6AHXxs7_0),.clk(gclk));
	jdff dff_A_TZZwCy5l3_0(.dout(w_dff_A_xV6AHXxs7_0),.din(w_dff_A_TZZwCy5l3_0),.clk(gclk));
	jdff dff_A_Z2vaiXFp1_0(.dout(w_dff_A_TZZwCy5l3_0),.din(w_dff_A_Z2vaiXFp1_0),.clk(gclk));
	jdff dff_B_g2OF9prz8_1(.din(n349),.dout(w_dff_B_g2OF9prz8_1),.clk(gclk));
	jdff dff_B_VEhLCr7G7_1(.din(n345),.dout(w_dff_B_VEhLCr7G7_1),.clk(gclk));
	jdff dff_B_XWBnabPj0_1(.din(w_dff_B_VEhLCr7G7_1),.dout(w_dff_B_XWBnabPj0_1),.clk(gclk));
	jdff dff_B_SzE7DbvA0_1(.din(w_dff_B_XWBnabPj0_1),.dout(w_dff_B_SzE7DbvA0_1),.clk(gclk));
	jdff dff_B_lrpHZXCg6_1(.din(w_dff_B_SzE7DbvA0_1),.dout(w_dff_B_lrpHZXCg6_1),.clk(gclk));
	jdff dff_B_idg45rYp0_1(.din(w_dff_B_lrpHZXCg6_1),.dout(w_dff_B_idg45rYp0_1),.clk(gclk));
	jdff dff_B_t6MrdRp72_1(.din(w_dff_B_idg45rYp0_1),.dout(w_dff_B_t6MrdRp72_1),.clk(gclk));
	jdff dff_B_FaUJ5Y8Z3_1(.din(w_dff_B_t6MrdRp72_1),.dout(w_dff_B_FaUJ5Y8Z3_1),.clk(gclk));
	jdff dff_B_ZraIwppx8_1(.din(w_dff_B_FaUJ5Y8Z3_1),.dout(w_dff_B_ZraIwppx8_1),.clk(gclk));
	jdff dff_B_ELXaCA7H8_1(.din(w_dff_B_ZraIwppx8_1),.dout(w_dff_B_ELXaCA7H8_1),.clk(gclk));
	jdff dff_B_6bEnps496_1(.din(w_dff_B_ELXaCA7H8_1),.dout(w_dff_B_6bEnps496_1),.clk(gclk));
	jdff dff_B_9Nqzcnkn1_1(.din(w_dff_B_6bEnps496_1),.dout(w_dff_B_9Nqzcnkn1_1),.clk(gclk));
	jdff dff_B_H2CNrLJG0_0(.din(n347),.dout(w_dff_B_H2CNrLJG0_0),.clk(gclk));
	jdff dff_B_Y0JdRT1V6_0(.din(w_dff_B_H2CNrLJG0_0),.dout(w_dff_B_Y0JdRT1V6_0),.clk(gclk));
	jdff dff_B_D6MFdtx69_0(.din(w_dff_B_Y0JdRT1V6_0),.dout(w_dff_B_D6MFdtx69_0),.clk(gclk));
	jdff dff_B_EfToIRyC9_0(.din(w_dff_B_D6MFdtx69_0),.dout(w_dff_B_EfToIRyC9_0),.clk(gclk));
	jdff dff_B_bg2glnvm3_0(.din(w_dff_B_EfToIRyC9_0),.dout(w_dff_B_bg2glnvm3_0),.clk(gclk));
	jdff dff_B_4tq0zEbH0_0(.din(w_dff_B_bg2glnvm3_0),.dout(w_dff_B_4tq0zEbH0_0),.clk(gclk));
	jdff dff_B_EeBHlsE48_0(.din(w_dff_B_4tq0zEbH0_0),.dout(w_dff_B_EeBHlsE48_0),.clk(gclk));
	jdff dff_B_aKeyEGGf3_0(.din(w_dff_B_EeBHlsE48_0),.dout(w_dff_B_aKeyEGGf3_0),.clk(gclk));
	jdff dff_B_K5RX96Or7_0(.din(w_dff_B_aKeyEGGf3_0),.dout(w_dff_B_K5RX96Or7_0),.clk(gclk));
	jdff dff_B_1qgJAdzW0_0(.din(w_dff_B_K5RX96Or7_0),.dout(w_dff_B_1qgJAdzW0_0),.clk(gclk));
	jdff dff_B_ZwQVbcg82_0(.din(w_dff_B_1qgJAdzW0_0),.dout(w_dff_B_ZwQVbcg82_0),.clk(gclk));
	jdff dff_B_Ych6BOQm9_0(.din(w_dff_B_ZwQVbcg82_0),.dout(w_dff_B_Ych6BOQm9_0),.clk(gclk));
	jdff dff_B_RVrt5Roe8_0(.din(w_dff_B_Ych6BOQm9_0),.dout(w_dff_B_RVrt5Roe8_0),.clk(gclk));
	jdff dff_B_x8rUjeRO8_0(.din(w_dff_B_RVrt5Roe8_0),.dout(w_dff_B_x8rUjeRO8_0),.clk(gclk));
	jdff dff_A_a40ZrbBV0_0(.dout(w_n346_0[0]),.din(w_dff_A_a40ZrbBV0_0),.clk(gclk));
	jdff dff_A_KS9CbfIl9_0(.dout(w_dff_A_a40ZrbBV0_0),.din(w_dff_A_KS9CbfIl9_0),.clk(gclk));
	jdff dff_A_x1JrpnHu2_0(.dout(w_dff_A_KS9CbfIl9_0),.din(w_dff_A_x1JrpnHu2_0),.clk(gclk));
	jdff dff_A_PjeSSwbs7_0(.dout(w_dff_A_x1JrpnHu2_0),.din(w_dff_A_PjeSSwbs7_0),.clk(gclk));
	jdff dff_A_pqi7Lsm11_0(.dout(w_dff_A_PjeSSwbs7_0),.din(w_dff_A_pqi7Lsm11_0),.clk(gclk));
	jdff dff_A_eDeewrIT1_0(.dout(w_dff_A_pqi7Lsm11_0),.din(w_dff_A_eDeewrIT1_0),.clk(gclk));
	jdff dff_A_9jk7Iiux0_0(.dout(w_dff_A_eDeewrIT1_0),.din(w_dff_A_9jk7Iiux0_0),.clk(gclk));
	jdff dff_A_1952PmuC5_0(.dout(w_dff_A_9jk7Iiux0_0),.din(w_dff_A_1952PmuC5_0),.clk(gclk));
	jdff dff_A_k4K5yYP36_0(.dout(w_dff_A_1952PmuC5_0),.din(w_dff_A_k4K5yYP36_0),.clk(gclk));
	jdff dff_A_2j38ThGE6_0(.dout(w_dff_A_k4K5yYP36_0),.din(w_dff_A_2j38ThGE6_0),.clk(gclk));
	jdff dff_A_UcdqNdcy2_0(.dout(w_dff_A_2j38ThGE6_0),.din(w_dff_A_UcdqNdcy2_0),.clk(gclk));
	jdff dff_A_cXUyKw9F2_0(.dout(w_dff_A_UcdqNdcy2_0),.din(w_dff_A_cXUyKw9F2_0),.clk(gclk));
	jdff dff_A_WX7shqmk3_0(.dout(w_dff_A_cXUyKw9F2_0),.din(w_dff_A_WX7shqmk3_0),.clk(gclk));
	jdff dff_A_eBCgRtde7_0(.dout(w_dff_A_WX7shqmk3_0),.din(w_dff_A_eBCgRtde7_0),.clk(gclk));
	jdff dff_A_R35ciefN3_0(.dout(w_dff_A_eBCgRtde7_0),.din(w_dff_A_R35ciefN3_0),.clk(gclk));
	jdff dff_B_2zSnQfFs1_1(.din(n358),.dout(w_dff_B_2zSnQfFs1_1),.clk(gclk));
	jdff dff_B_l8X87IZS8_1(.din(n354),.dout(w_dff_B_l8X87IZS8_1),.clk(gclk));
	jdff dff_B_DfWMo8wB9_1(.din(w_dff_B_l8X87IZS8_1),.dout(w_dff_B_DfWMo8wB9_1),.clk(gclk));
	jdff dff_B_3g5Nk9NH1_1(.din(w_dff_B_DfWMo8wB9_1),.dout(w_dff_B_3g5Nk9NH1_1),.clk(gclk));
	jdff dff_B_MA4W0IWu2_1(.din(w_dff_B_3g5Nk9NH1_1),.dout(w_dff_B_MA4W0IWu2_1),.clk(gclk));
	jdff dff_B_SH0MrZEv1_1(.din(w_dff_B_MA4W0IWu2_1),.dout(w_dff_B_SH0MrZEv1_1),.clk(gclk));
	jdff dff_B_9bOzUXyW0_1(.din(w_dff_B_SH0MrZEv1_1),.dout(w_dff_B_9bOzUXyW0_1),.clk(gclk));
	jdff dff_B_o1sQQcrB5_1(.din(w_dff_B_9bOzUXyW0_1),.dout(w_dff_B_o1sQQcrB5_1),.clk(gclk));
	jdff dff_B_sMMOgGKX7_1(.din(w_dff_B_o1sQQcrB5_1),.dout(w_dff_B_sMMOgGKX7_1),.clk(gclk));
	jdff dff_B_6INdmnwJ1_1(.din(w_dff_B_sMMOgGKX7_1),.dout(w_dff_B_6INdmnwJ1_1),.clk(gclk));
	jdff dff_B_kskOGiI54_1(.din(w_dff_B_6INdmnwJ1_1),.dout(w_dff_B_kskOGiI54_1),.clk(gclk));
	jdff dff_B_asEVOhQ28_1(.din(w_dff_B_kskOGiI54_1),.dout(w_dff_B_asEVOhQ28_1),.clk(gclk));
	jdff dff_B_JUyNBap41_0(.din(n356),.dout(w_dff_B_JUyNBap41_0),.clk(gclk));
	jdff dff_B_rSUV66cp1_0(.din(w_dff_B_JUyNBap41_0),.dout(w_dff_B_rSUV66cp1_0),.clk(gclk));
	jdff dff_B_QyQySQpP7_0(.din(w_dff_B_rSUV66cp1_0),.dout(w_dff_B_QyQySQpP7_0),.clk(gclk));
	jdff dff_B_G1D6aLzB0_0(.din(w_dff_B_QyQySQpP7_0),.dout(w_dff_B_G1D6aLzB0_0),.clk(gclk));
	jdff dff_B_t4xgzVOG1_0(.din(w_dff_B_G1D6aLzB0_0),.dout(w_dff_B_t4xgzVOG1_0),.clk(gclk));
	jdff dff_B_3kqAcaaz4_0(.din(w_dff_B_t4xgzVOG1_0),.dout(w_dff_B_3kqAcaaz4_0),.clk(gclk));
	jdff dff_B_31AUgmxW9_0(.din(w_dff_B_3kqAcaaz4_0),.dout(w_dff_B_31AUgmxW9_0),.clk(gclk));
	jdff dff_B_Bms54Ufo4_0(.din(w_dff_B_31AUgmxW9_0),.dout(w_dff_B_Bms54Ufo4_0),.clk(gclk));
	jdff dff_B_cYH2h23q3_0(.din(w_dff_B_Bms54Ufo4_0),.dout(w_dff_B_cYH2h23q3_0),.clk(gclk));
	jdff dff_B_eeIkLifw7_0(.din(w_dff_B_cYH2h23q3_0),.dout(w_dff_B_eeIkLifw7_0),.clk(gclk));
	jdff dff_B_hNMRWYNp3_0(.din(w_dff_B_eeIkLifw7_0),.dout(w_dff_B_hNMRWYNp3_0),.clk(gclk));
	jdff dff_B_sPE2No0Z4_0(.din(w_dff_B_hNMRWYNp3_0),.dout(w_dff_B_sPE2No0Z4_0),.clk(gclk));
	jdff dff_B_3voJP80T0_0(.din(w_dff_B_sPE2No0Z4_0),.dout(w_dff_B_3voJP80T0_0),.clk(gclk));
	jdff dff_B_pgBGJOFz1_0(.din(w_dff_B_3voJP80T0_0),.dout(w_dff_B_pgBGJOFz1_0),.clk(gclk));
	jdff dff_A_xcYwUVsO8_0(.dout(w_n355_0[0]),.din(w_dff_A_xcYwUVsO8_0),.clk(gclk));
	jdff dff_A_N6lIisni1_0(.dout(w_dff_A_xcYwUVsO8_0),.din(w_dff_A_N6lIisni1_0),.clk(gclk));
	jdff dff_A_7jPaRy5k4_0(.dout(w_dff_A_N6lIisni1_0),.din(w_dff_A_7jPaRy5k4_0),.clk(gclk));
	jdff dff_A_ak4shpa80_0(.dout(w_dff_A_7jPaRy5k4_0),.din(w_dff_A_ak4shpa80_0),.clk(gclk));
	jdff dff_A_NyE7DK9t8_0(.dout(w_dff_A_ak4shpa80_0),.din(w_dff_A_NyE7DK9t8_0),.clk(gclk));
	jdff dff_A_qjrtIxys2_0(.dout(w_dff_A_NyE7DK9t8_0),.din(w_dff_A_qjrtIxys2_0),.clk(gclk));
	jdff dff_A_HcpEG8lA1_0(.dout(w_dff_A_qjrtIxys2_0),.din(w_dff_A_HcpEG8lA1_0),.clk(gclk));
	jdff dff_A_1yBdBzXG3_0(.dout(w_dff_A_HcpEG8lA1_0),.din(w_dff_A_1yBdBzXG3_0),.clk(gclk));
	jdff dff_A_MneI7HUb6_0(.dout(w_dff_A_1yBdBzXG3_0),.din(w_dff_A_MneI7HUb6_0),.clk(gclk));
	jdff dff_A_craBofKo4_0(.dout(w_dff_A_MneI7HUb6_0),.din(w_dff_A_craBofKo4_0),.clk(gclk));
	jdff dff_A_GIk3ME9r6_0(.dout(w_dff_A_craBofKo4_0),.din(w_dff_A_GIk3ME9r6_0),.clk(gclk));
	jdff dff_A_xIxoSfj75_0(.dout(w_dff_A_GIk3ME9r6_0),.din(w_dff_A_xIxoSfj75_0),.clk(gclk));
	jdff dff_A_rVfHl5V13_0(.dout(w_dff_A_xIxoSfj75_0),.din(w_dff_A_rVfHl5V13_0),.clk(gclk));
	jdff dff_A_3m4Gm8CY2_0(.dout(w_dff_A_rVfHl5V13_0),.din(w_dff_A_3m4Gm8CY2_0),.clk(gclk));
	jdff dff_A_LrjQo2z18_0(.dout(w_dff_A_3m4Gm8CY2_0),.din(w_dff_A_LrjQo2z18_0),.clk(gclk));
	jdff dff_B_wmO4A6qe3_1(.din(n367),.dout(w_dff_B_wmO4A6qe3_1),.clk(gclk));
	jdff dff_B_jmLswqoX8_1(.din(n363),.dout(w_dff_B_jmLswqoX8_1),.clk(gclk));
	jdff dff_B_9h9Ky1mg4_1(.din(w_dff_B_jmLswqoX8_1),.dout(w_dff_B_9h9Ky1mg4_1),.clk(gclk));
	jdff dff_B_deW99Fmt3_1(.din(w_dff_B_9h9Ky1mg4_1),.dout(w_dff_B_deW99Fmt3_1),.clk(gclk));
	jdff dff_B_J9o3XUjZ7_1(.din(w_dff_B_deW99Fmt3_1),.dout(w_dff_B_J9o3XUjZ7_1),.clk(gclk));
	jdff dff_B_fUReB4hX0_1(.din(w_dff_B_J9o3XUjZ7_1),.dout(w_dff_B_fUReB4hX0_1),.clk(gclk));
	jdff dff_B_cqtGVioD4_1(.din(w_dff_B_fUReB4hX0_1),.dout(w_dff_B_cqtGVioD4_1),.clk(gclk));
	jdff dff_B_OajuNvdD9_1(.din(w_dff_B_cqtGVioD4_1),.dout(w_dff_B_OajuNvdD9_1),.clk(gclk));
	jdff dff_B_q63v1enh3_1(.din(w_dff_B_OajuNvdD9_1),.dout(w_dff_B_q63v1enh3_1),.clk(gclk));
	jdff dff_B_9aVBX27z9_1(.din(w_dff_B_q63v1enh3_1),.dout(w_dff_B_9aVBX27z9_1),.clk(gclk));
	jdff dff_B_PFtwNMs62_1(.din(w_dff_B_9aVBX27z9_1),.dout(w_dff_B_PFtwNMs62_1),.clk(gclk));
	jdff dff_B_7HXfiGRz1_1(.din(w_dff_B_PFtwNMs62_1),.dout(w_dff_B_7HXfiGRz1_1),.clk(gclk));
	jdff dff_B_wYPCkrPE6_0(.din(n365),.dout(w_dff_B_wYPCkrPE6_0),.clk(gclk));
	jdff dff_B_yCtKu4ji2_0(.din(w_dff_B_wYPCkrPE6_0),.dout(w_dff_B_yCtKu4ji2_0),.clk(gclk));
	jdff dff_B_v0X3FtpK1_0(.din(w_dff_B_yCtKu4ji2_0),.dout(w_dff_B_v0X3FtpK1_0),.clk(gclk));
	jdff dff_B_MlQIv1ZU5_0(.din(w_dff_B_v0X3FtpK1_0),.dout(w_dff_B_MlQIv1ZU5_0),.clk(gclk));
	jdff dff_B_6kqHQUWw3_0(.din(w_dff_B_MlQIv1ZU5_0),.dout(w_dff_B_6kqHQUWw3_0),.clk(gclk));
	jdff dff_B_SOYqLUKg1_0(.din(w_dff_B_6kqHQUWw3_0),.dout(w_dff_B_SOYqLUKg1_0),.clk(gclk));
	jdff dff_B_xjELT74o9_0(.din(w_dff_B_SOYqLUKg1_0),.dout(w_dff_B_xjELT74o9_0),.clk(gclk));
	jdff dff_B_rYcgpTRV5_0(.din(w_dff_B_xjELT74o9_0),.dout(w_dff_B_rYcgpTRV5_0),.clk(gclk));
	jdff dff_B_WtvNf9XZ2_0(.din(w_dff_B_rYcgpTRV5_0),.dout(w_dff_B_WtvNf9XZ2_0),.clk(gclk));
	jdff dff_B_HjZuLwPn8_0(.din(w_dff_B_WtvNf9XZ2_0),.dout(w_dff_B_HjZuLwPn8_0),.clk(gclk));
	jdff dff_B_KurlW3CV9_0(.din(w_dff_B_HjZuLwPn8_0),.dout(w_dff_B_KurlW3CV9_0),.clk(gclk));
	jdff dff_B_fBMT03aO5_0(.din(w_dff_B_KurlW3CV9_0),.dout(w_dff_B_fBMT03aO5_0),.clk(gclk));
	jdff dff_B_YPb2xc1Q6_0(.din(w_dff_B_fBMT03aO5_0),.dout(w_dff_B_YPb2xc1Q6_0),.clk(gclk));
	jdff dff_B_QxqH7i8L4_0(.din(w_dff_B_YPb2xc1Q6_0),.dout(w_dff_B_QxqH7i8L4_0),.clk(gclk));
	jdff dff_A_iOWFAiQM5_0(.dout(w_n364_0[0]),.din(w_dff_A_iOWFAiQM5_0),.clk(gclk));
	jdff dff_A_EYuRxxkG1_0(.dout(w_dff_A_iOWFAiQM5_0),.din(w_dff_A_EYuRxxkG1_0),.clk(gclk));
	jdff dff_A_4tEwtDPz3_0(.dout(w_dff_A_EYuRxxkG1_0),.din(w_dff_A_4tEwtDPz3_0),.clk(gclk));
	jdff dff_A_3akT1Pd26_0(.dout(w_dff_A_4tEwtDPz3_0),.din(w_dff_A_3akT1Pd26_0),.clk(gclk));
	jdff dff_A_cbYSRxgy4_0(.dout(w_dff_A_3akT1Pd26_0),.din(w_dff_A_cbYSRxgy4_0),.clk(gclk));
	jdff dff_A_4ykiYK3i2_0(.dout(w_dff_A_cbYSRxgy4_0),.din(w_dff_A_4ykiYK3i2_0),.clk(gclk));
	jdff dff_A_kCMJas7z6_0(.dout(w_dff_A_4ykiYK3i2_0),.din(w_dff_A_kCMJas7z6_0),.clk(gclk));
	jdff dff_A_InaOq4ub2_0(.dout(w_dff_A_kCMJas7z6_0),.din(w_dff_A_InaOq4ub2_0),.clk(gclk));
	jdff dff_A_g4RHG3ie2_0(.dout(w_dff_A_InaOq4ub2_0),.din(w_dff_A_g4RHG3ie2_0),.clk(gclk));
	jdff dff_A_9ovgboK87_0(.dout(w_dff_A_g4RHG3ie2_0),.din(w_dff_A_9ovgboK87_0),.clk(gclk));
	jdff dff_A_VbPYCV4X0_0(.dout(w_dff_A_9ovgboK87_0),.din(w_dff_A_VbPYCV4X0_0),.clk(gclk));
	jdff dff_A_lKUXeGMP7_0(.dout(w_dff_A_VbPYCV4X0_0),.din(w_dff_A_lKUXeGMP7_0),.clk(gclk));
	jdff dff_A_FtDOVRwm1_0(.dout(w_dff_A_lKUXeGMP7_0),.din(w_dff_A_FtDOVRwm1_0),.clk(gclk));
	jdff dff_A_U6VZd5uT4_0(.dout(w_dff_A_FtDOVRwm1_0),.din(w_dff_A_U6VZd5uT4_0),.clk(gclk));
	jdff dff_A_g4DgAnzk9_0(.dout(w_dff_A_U6VZd5uT4_0),.din(w_dff_A_g4DgAnzk9_0),.clk(gclk));
	jdff dff_B_Z1UoXxNG6_1(.din(n374),.dout(w_dff_B_Z1UoXxNG6_1),.clk(gclk));
	jdff dff_B_TR4RPDZZ8_0(.din(n375),.dout(w_dff_B_TR4RPDZZ8_0),.clk(gclk));
	jdff dff_B_O6hyf5kI2_0(.din(w_dff_B_TR4RPDZZ8_0),.dout(w_dff_B_O6hyf5kI2_0),.clk(gclk));
	jdff dff_B_frALq1aB9_0(.din(w_dff_B_O6hyf5kI2_0),.dout(w_dff_B_frALq1aB9_0),.clk(gclk));
	jdff dff_B_2scBKyAd7_0(.din(w_dff_B_frALq1aB9_0),.dout(w_dff_B_2scBKyAd7_0),.clk(gclk));
	jdff dff_B_Y8c7gJsy9_0(.din(w_dff_B_2scBKyAd7_0),.dout(w_dff_B_Y8c7gJsy9_0),.clk(gclk));
	jdff dff_B_1q9kFu5r6_0(.din(w_dff_B_Y8c7gJsy9_0),.dout(w_dff_B_1q9kFu5r6_0),.clk(gclk));
	jdff dff_B_1vfvWWWA0_0(.din(w_dff_B_1q9kFu5r6_0),.dout(w_dff_B_1vfvWWWA0_0),.clk(gclk));
	jdff dff_B_4kM0jMEn1_0(.din(w_dff_B_1vfvWWWA0_0),.dout(w_dff_B_4kM0jMEn1_0),.clk(gclk));
	jdff dff_B_QgX8oHX47_0(.din(w_dff_B_4kM0jMEn1_0),.dout(w_dff_B_QgX8oHX47_0),.clk(gclk));
	jdff dff_B_p43JBJuH3_0(.din(w_dff_B_QgX8oHX47_0),.dout(w_dff_B_p43JBJuH3_0),.clk(gclk));
	jdff dff_B_71GvA6f68_0(.din(w_dff_B_p43JBJuH3_0),.dout(w_dff_B_71GvA6f68_0),.clk(gclk));
	jdff dff_B_af2l6ZNy0_0(.din(w_dff_B_71GvA6f68_0),.dout(w_dff_B_af2l6ZNy0_0),.clk(gclk));
	jdff dff_B_ybnAZrxV0_0(.din(w_dff_B_af2l6ZNy0_0),.dout(w_dff_B_ybnAZrxV0_0),.clk(gclk));
	jdff dff_B_oWeEm77E3_0(.din(w_dff_B_ybnAZrxV0_0),.dout(w_dff_B_oWeEm77E3_0),.clk(gclk));
	jdff dff_A_Nv30eQLC1_1(.dout(w_n372_0[1]),.din(w_dff_A_Nv30eQLC1_1),.clk(gclk));
	jdff dff_A_xmggtavh0_1(.dout(w_dff_A_Nv30eQLC1_1),.din(w_dff_A_xmggtavh0_1),.clk(gclk));
	jdff dff_A_95ILcNr92_1(.dout(w_dff_A_xmggtavh0_1),.din(w_dff_A_95ILcNr92_1),.clk(gclk));
	jdff dff_A_SMEdqSmF8_1(.dout(w_dff_A_95ILcNr92_1),.din(w_dff_A_SMEdqSmF8_1),.clk(gclk));
	jdff dff_A_b2oZaGwc0_1(.dout(w_dff_A_SMEdqSmF8_1),.din(w_dff_A_b2oZaGwc0_1),.clk(gclk));
	jdff dff_A_GcyNs0mk0_1(.dout(w_dff_A_b2oZaGwc0_1),.din(w_dff_A_GcyNs0mk0_1),.clk(gclk));
	jdff dff_A_YsLtPPyd4_1(.dout(w_dff_A_GcyNs0mk0_1),.din(w_dff_A_YsLtPPyd4_1),.clk(gclk));
	jdff dff_A_BJg2hu6n1_1(.dout(w_dff_A_YsLtPPyd4_1),.din(w_dff_A_BJg2hu6n1_1),.clk(gclk));
	jdff dff_A_nCy55j0m5_1(.dout(w_dff_A_BJg2hu6n1_1),.din(w_dff_A_nCy55j0m5_1),.clk(gclk));
	jdff dff_A_94VjiY8l0_1(.dout(w_dff_A_nCy55j0m5_1),.din(w_dff_A_94VjiY8l0_1),.clk(gclk));
	jdff dff_A_5PIyMaYk5_1(.dout(w_dff_A_94VjiY8l0_1),.din(w_dff_A_5PIyMaYk5_1),.clk(gclk));
	jdff dff_A_AHCK4zuY1_1(.dout(w_dff_A_5PIyMaYk5_1),.din(w_dff_A_AHCK4zuY1_1),.clk(gclk));
	jdff dff_A_5S1WgPzl9_1(.dout(w_dff_A_AHCK4zuY1_1),.din(w_dff_A_5S1WgPzl9_1),.clk(gclk));
	jdff dff_A_q94WGlpI1_1(.dout(w_dff_A_5S1WgPzl9_1),.din(w_dff_A_q94WGlpI1_1),.clk(gclk));
	jdff dff_A_cfi4m6ds0_1(.dout(w_dff_A_q94WGlpI1_1),.din(w_dff_A_cfi4m6ds0_1),.clk(gclk));
	jdff dff_B_auJy2zN15_1(.din(n380),.dout(w_dff_B_auJy2zN15_1),.clk(gclk));
	jdff dff_B_qsfCuBTl5_1(.din(w_dff_B_auJy2zN15_1),.dout(w_dff_B_qsfCuBTl5_1),.clk(gclk));
	jdff dff_B_KziesRIi4_1(.din(w_dff_B_qsfCuBTl5_1),.dout(w_dff_B_KziesRIi4_1),.clk(gclk));
	jdff dff_B_oytCqnNi5_1(.din(w_dff_B_KziesRIi4_1),.dout(w_dff_B_oytCqnNi5_1),.clk(gclk));
	jdff dff_B_BOPJdd9c7_1(.din(w_dff_B_oytCqnNi5_1),.dout(w_dff_B_BOPJdd9c7_1),.clk(gclk));
	jdff dff_B_Yc330sQ48_1(.din(w_dff_B_BOPJdd9c7_1),.dout(w_dff_B_Yc330sQ48_1),.clk(gclk));
	jdff dff_B_c1neUtE09_1(.din(w_dff_B_Yc330sQ48_1),.dout(w_dff_B_c1neUtE09_1),.clk(gclk));
	jdff dff_B_ZoSHi2uY1_1(.din(w_dff_B_c1neUtE09_1),.dout(w_dff_B_ZoSHi2uY1_1),.clk(gclk));
	jdff dff_B_WR5UWy2s3_1(.din(w_dff_B_ZoSHi2uY1_1),.dout(w_dff_B_WR5UWy2s3_1),.clk(gclk));
	jdff dff_B_kRtO0J5R1_1(.din(w_dff_B_WR5UWy2s3_1),.dout(w_dff_B_kRtO0J5R1_1),.clk(gclk));
	jdff dff_B_zdCjIH5i0_1(.din(w_dff_B_kRtO0J5R1_1),.dout(w_dff_B_zdCjIH5i0_1),.clk(gclk));
	jdff dff_B_hZt06uKP7_1(.din(w_dff_B_zdCjIH5i0_1),.dout(w_dff_B_hZt06uKP7_1),.clk(gclk));
	jdff dff_B_4XIhDDXP0_1(.din(w_dff_B_hZt06uKP7_1),.dout(w_dff_B_4XIhDDXP0_1),.clk(gclk));
	jdff dff_B_GTdvnyGC8_1(.din(w_dff_B_4XIhDDXP0_1),.dout(w_dff_B_GTdvnyGC8_1),.clk(gclk));
	jdff dff_B_TEb94CHB0_1(.din(w_dff_B_GTdvnyGC8_1),.dout(w_dff_B_TEb94CHB0_1),.clk(gclk));
	jdff dff_B_6soSkoXO6_0(.din(n382),.dout(w_dff_B_6soSkoXO6_0),.clk(gclk));
	jdff dff_B_Y3w9aD0W7_0(.din(w_dff_B_6soSkoXO6_0),.dout(w_dff_B_Y3w9aD0W7_0),.clk(gclk));
	jdff dff_B_yKKNmLjm2_0(.din(w_dff_B_Y3w9aD0W7_0),.dout(w_dff_B_yKKNmLjm2_0),.clk(gclk));
	jdff dff_B_3h6HTqAb8_0(.din(w_dff_B_yKKNmLjm2_0),.dout(w_dff_B_3h6HTqAb8_0),.clk(gclk));
	jdff dff_B_40FnlNyZ3_0(.din(w_dff_B_3h6HTqAb8_0),.dout(w_dff_B_40FnlNyZ3_0),.clk(gclk));
	jdff dff_B_MMFoMroI5_0(.din(w_dff_B_40FnlNyZ3_0),.dout(w_dff_B_MMFoMroI5_0),.clk(gclk));
	jdff dff_B_8RR9m6Ve9_0(.din(w_dff_B_MMFoMroI5_0),.dout(w_dff_B_8RR9m6Ve9_0),.clk(gclk));
	jdff dff_B_9D8b6rVG3_0(.din(w_dff_B_8RR9m6Ve9_0),.dout(w_dff_B_9D8b6rVG3_0),.clk(gclk));
	jdff dff_B_wu922Bbp0_0(.din(w_dff_B_9D8b6rVG3_0),.dout(w_dff_B_wu922Bbp0_0),.clk(gclk));
	jdff dff_B_btWV6d8S1_0(.din(w_dff_B_wu922Bbp0_0),.dout(w_dff_B_btWV6d8S1_0),.clk(gclk));
	jdff dff_B_SDE0ZuKW0_0(.din(w_dff_B_btWV6d8S1_0),.dout(w_dff_B_SDE0ZuKW0_0),.clk(gclk));
	jdff dff_B_VutXt6i25_0(.din(w_dff_B_SDE0ZuKW0_0),.dout(w_dff_B_VutXt6i25_0),.clk(gclk));
	jdff dff_B_q8s1OkMF9_0(.din(w_dff_B_VutXt6i25_0),.dout(w_dff_B_q8s1OkMF9_0),.clk(gclk));
	jdff dff_B_GsXdjJPE0_0(.din(w_dff_B_q8s1OkMF9_0),.dout(w_dff_B_GsXdjJPE0_0),.clk(gclk));
	jdff dff_B_twuoMNpP3_0(.din(n392),.dout(w_dff_B_twuoMNpP3_0),.clk(gclk));
	jdff dff_B_TKpuWm7I1_0(.din(w_dff_B_twuoMNpP3_0),.dout(w_dff_B_TKpuWm7I1_0),.clk(gclk));
	jdff dff_B_vDz0SzSY1_0(.din(w_dff_B_TKpuWm7I1_0),.dout(w_dff_B_vDz0SzSY1_0),.clk(gclk));
	jdff dff_B_NUY7oWDt9_0(.din(w_dff_B_vDz0SzSY1_0),.dout(w_dff_B_NUY7oWDt9_0),.clk(gclk));
	jdff dff_B_Esqf7SVr8_0(.din(w_dff_B_NUY7oWDt9_0),.dout(w_dff_B_Esqf7SVr8_0),.clk(gclk));
	jdff dff_B_z3NEQ4bB6_0(.din(w_dff_B_Esqf7SVr8_0),.dout(w_dff_B_z3NEQ4bB6_0),.clk(gclk));
	jdff dff_B_qvxlqp2j2_0(.din(w_dff_B_z3NEQ4bB6_0),.dout(w_dff_B_qvxlqp2j2_0),.clk(gclk));
	jdff dff_B_WEKewzHa9_0(.din(w_dff_B_qvxlqp2j2_0),.dout(w_dff_B_WEKewzHa9_0),.clk(gclk));
	jdff dff_B_bbuANj3p2_0(.din(w_dff_B_WEKewzHa9_0),.dout(w_dff_B_bbuANj3p2_0),.clk(gclk));
	jdff dff_B_4sBnFaE23_0(.din(w_dff_B_bbuANj3p2_0),.dout(w_dff_B_4sBnFaE23_0),.clk(gclk));
	jdff dff_B_3ezn6Tq90_0(.din(w_dff_B_4sBnFaE23_0),.dout(w_dff_B_3ezn6Tq90_0),.clk(gclk));
	jdff dff_B_Hc6JuZM87_1(.din(n390),.dout(w_dff_B_Hc6JuZM87_1),.clk(gclk));
	jdff dff_B_6PMUkzqF5_1(.din(w_dff_B_Hc6JuZM87_1),.dout(w_dff_B_6PMUkzqF5_1),.clk(gclk));
	jdff dff_B_SllIQFCA4_0(.din(n388),.dout(w_dff_B_SllIQFCA4_0),.clk(gclk));
	jdff dff_B_zFtMBBRt8_0(.din(w_dff_B_SllIQFCA4_0),.dout(w_dff_B_zFtMBBRt8_0),.clk(gclk));
	jdff dff_B_AhKVwmre3_0(.din(w_dff_B_zFtMBBRt8_0),.dout(w_dff_B_AhKVwmre3_0),.clk(gclk));
	jdff dff_B_kppAuLRK1_0(.din(w_dff_B_AhKVwmre3_0),.dout(w_dff_B_kppAuLRK1_0),.clk(gclk));
	jdff dff_B_f0LYQgLJ5_0(.din(w_dff_B_kppAuLRK1_0),.dout(w_dff_B_f0LYQgLJ5_0),.clk(gclk));
	jdff dff_B_ArSjcsta0_0(.din(w_dff_B_f0LYQgLJ5_0),.dout(w_dff_B_ArSjcsta0_0),.clk(gclk));
	jdff dff_B_3cKr2Jdv2_0(.din(w_dff_B_ArSjcsta0_0),.dout(w_dff_B_3cKr2Jdv2_0),.clk(gclk));
	jdff dff_B_kMhhQDeI1_0(.din(w_dff_B_3cKr2Jdv2_0),.dout(w_dff_B_kMhhQDeI1_0),.clk(gclk));
	jdff dff_B_K6MMRE9n1_0(.din(w_dff_B_kMhhQDeI1_0),.dout(w_dff_B_K6MMRE9n1_0),.clk(gclk));
	jdff dff_B_4swiCMCz1_0(.din(w_dff_B_K6MMRE9n1_0),.dout(w_dff_B_4swiCMCz1_0),.clk(gclk));
	jdff dff_B_PfseflL70_0(.din(w_dff_B_4swiCMCz1_0),.dout(w_dff_B_PfseflL70_0),.clk(gclk));
	jdff dff_B_sHmvpdd74_0(.din(w_dff_B_PfseflL70_0),.dout(w_dff_B_sHmvpdd74_0),.clk(gclk));
	jdff dff_B_PeeA8JVj0_0(.din(w_dff_B_sHmvpdd74_0),.dout(w_dff_B_PeeA8JVj0_0),.clk(gclk));
	jdff dff_B_HjcMotW98_1(.din(n398),.dout(w_dff_B_HjcMotW98_1),.clk(gclk));
	jdff dff_B_h0UcXPex1_0(.din(n224),.dout(w_dff_B_h0UcXPex1_0),.clk(gclk));
	jdff dff_A_9ps5Vm5Q7_0(.dout(w_n218_1[0]),.din(w_dff_A_9ps5Vm5Q7_0),.clk(gclk));
	jdff dff_A_IHqyDOlI7_0(.dout(w_n218_0[0]),.din(w_dff_A_IHqyDOlI7_0),.clk(gclk));
	jdff dff_A_JWHs09d71_2(.dout(w_n218_0[2]),.din(w_dff_A_JWHs09d71_2),.clk(gclk));
	jdff dff_A_LORqUJdb7_2(.dout(w_dff_A_JWHs09d71_2),.din(w_dff_A_LORqUJdb7_2),.clk(gclk));
	jdff dff_A_NQaIJkRP2_0(.dout(w_n192_0[0]),.din(w_dff_A_NQaIJkRP2_0),.clk(gclk));
	jdff dff_A_8q8lNVYD4_2(.dout(w_n192_0[2]),.din(w_dff_A_8q8lNVYD4_2),.clk(gclk));
	jdff dff_B_i6lhBmlg3_3(.din(n192),.dout(w_dff_B_i6lhBmlg3_3),.clk(gclk));
	jdff dff_B_mFbBRedQ8_0(.din(n209),.dout(w_dff_B_mFbBRedQ8_0),.clk(gclk));
	jdff dff_A_zDeAIA3f6_0(.dout(w_n198_0[0]),.din(w_dff_A_zDeAIA3f6_0),.clk(gclk));
	jdff dff_A_mnwbm1S54_2(.dout(w_n198_0[2]),.din(w_dff_A_mnwbm1S54_2),.clk(gclk));
	jdff dff_A_HaA4EzaU8_2(.dout(w_dff_A_mnwbm1S54_2),.din(w_dff_A_HaA4EzaU8_2),.clk(gclk));
	jdff dff_A_q3Bn0c1F6_0(.dout(w_n197_1[0]),.din(w_dff_A_q3Bn0c1F6_0),.clk(gclk));
	jdff dff_A_hiMHTam68_0(.dout(w_dff_A_q3Bn0c1F6_0),.din(w_dff_A_hiMHTam68_0),.clk(gclk));
	jdff dff_A_tUnjq15O9_1(.dout(w_n197_0[1]),.din(w_dff_A_tUnjq15O9_1),.clk(gclk));
	jdff dff_A_H7gxCzUt6_1(.dout(w_dff_A_tUnjq15O9_1),.din(w_dff_A_H7gxCzUt6_1),.clk(gclk));
	jdff dff_A_ppa3Ic6i2_0(.dout(w_n155_0[0]),.din(w_dff_A_ppa3Ic6i2_0),.clk(gclk));
	jdff dff_A_BItCi9uA1_2(.dout(w_n155_0[2]),.din(w_dff_A_BItCi9uA1_2),.clk(gclk));
	jdff dff_B_UBOMW93A9_3(.din(n155),.dout(w_dff_B_UBOMW93A9_3),.clk(gclk));
	jdff dff_A_jmnqiUNg7_0(.dout(w_n144_1[0]),.din(w_dff_A_jmnqiUNg7_0),.clk(gclk));
	jdff dff_A_4Gp49ERV3_0(.dout(w_dff_A_jmnqiUNg7_0),.din(w_dff_A_4Gp49ERV3_0),.clk(gclk));
	jdff dff_A_kmByPNTj0_1(.dout(w_n144_0[1]),.din(w_dff_A_kmByPNTj0_1),.clk(gclk));
	jdff dff_A_2KEevYyh8_1(.dout(w_dff_A_kmByPNTj0_1),.din(w_dff_A_2KEevYyh8_1),.clk(gclk));
	jdff dff_A_JLyGu4V98_2(.dout(w_n159_0[2]),.din(w_dff_A_JLyGu4V98_2),.clk(gclk));
	jdff dff_A_MLI46m0M2_2(.dout(w_dff_A_JLyGu4V98_2),.din(w_dff_A_MLI46m0M2_2),.clk(gclk));
	jdff dff_A_0CYnpiTc0_2(.dout(w_n121_0[2]),.din(w_dff_A_0CYnpiTc0_2),.clk(gclk));
	jdff dff_B_Vs822WDe7_3(.din(n121),.dout(w_dff_B_Vs822WDe7_3),.clk(gclk));
	jdff dff_A_ZeOdPqkX6_1(.dout(w_n96_0[1]),.din(w_dff_A_ZeOdPqkX6_1),.clk(gclk));
	jdff dff_A_VfQnigIX0_1(.dout(w_dff_A_ZeOdPqkX6_1),.din(w_dff_A_VfQnigIX0_1),.clk(gclk));
	jdff dff_A_95ZYmOEK6_1(.dout(w_dff_A_VfQnigIX0_1),.din(w_dff_A_95ZYmOEK6_1),.clk(gclk));
	jdff dff_A_ArFhudP54_1(.dout(w_dff_A_95ZYmOEK6_1),.din(w_dff_A_ArFhudP54_1),.clk(gclk));
	jdff dff_A_BppLuG0Q2_2(.dout(w_n96_0[2]),.din(w_dff_A_BppLuG0Q2_2),.clk(gclk));
	jdff dff_A_q0ph1p8R6_2(.dout(w_dff_A_BppLuG0Q2_2),.din(w_dff_A_q0ph1p8R6_2),.clk(gclk));
	jdff dff_A_jNgry8Oy4_2(.dout(w_dff_A_q0ph1p8R6_2),.din(w_dff_A_jNgry8Oy4_2),.clk(gclk));
	jdff dff_A_wq4tQ5FZ0_2(.dout(w_dff_A_jNgry8Oy4_2),.din(w_dff_A_wq4tQ5FZ0_2),.clk(gclk));
	jdff dff_B_l9DezJPm0_3(.din(n340),.dout(w_dff_B_l9DezJPm0_3),.clk(gclk));
	jdff dff_B_WWkWQFP10_3(.din(w_dff_B_l9DezJPm0_3),.dout(w_dff_B_WWkWQFP10_3),.clk(gclk));
	jdff dff_B_KA9k3SP01_3(.din(w_dff_B_WWkWQFP10_3),.dout(w_dff_B_KA9k3SP01_3),.clk(gclk));
	jdff dff_B_wrDOKcW35_3(.din(w_dff_B_KA9k3SP01_3),.dout(w_dff_B_wrDOKcW35_3),.clk(gclk));
	jdff dff_B_5UkqvjVw4_3(.din(w_dff_B_wrDOKcW35_3),.dout(w_dff_B_5UkqvjVw4_3),.clk(gclk));
	jdff dff_B_8DJu24hh8_3(.din(w_dff_B_5UkqvjVw4_3),.dout(w_dff_B_8DJu24hh8_3),.clk(gclk));
	jdff dff_B_i4QGAl8O1_3(.din(w_dff_B_8DJu24hh8_3),.dout(w_dff_B_i4QGAl8O1_3),.clk(gclk));
	jdff dff_B_DbVdrO6Q3_3(.din(w_dff_B_i4QGAl8O1_3),.dout(w_dff_B_DbVdrO6Q3_3),.clk(gclk));
	jdff dff_B_VTHx8ntN8_3(.din(w_dff_B_DbVdrO6Q3_3),.dout(w_dff_B_VTHx8ntN8_3),.clk(gclk));
	jdff dff_B_lmQytfA50_3(.din(w_dff_B_VTHx8ntN8_3),.dout(w_dff_B_lmQytfA50_3),.clk(gclk));
	jdff dff_B_xrTHEsuz2_3(.din(w_dff_B_lmQytfA50_3),.dout(w_dff_B_xrTHEsuz2_3),.clk(gclk));
	jdff dff_B_EjkoS64Q3_3(.din(w_dff_B_xrTHEsuz2_3),.dout(w_dff_B_EjkoS64Q3_3),.clk(gclk));
	jdff dff_B_Db3ZMv005_3(.din(w_dff_B_EjkoS64Q3_3),.dout(w_dff_B_Db3ZMv005_3),.clk(gclk));
	jdff dff_B_dAipauU12_3(.din(w_dff_B_Db3ZMv005_3),.dout(w_dff_B_dAipauU12_3),.clk(gclk));
	jdff dff_B_xj0wtFRl3_3(.din(w_dff_B_dAipauU12_3),.dout(w_dff_B_xj0wtFRl3_3),.clk(gclk));
	jdff dff_B_92ZUkadt7_3(.din(w_dff_B_xj0wtFRl3_3),.dout(w_dff_B_92ZUkadt7_3),.clk(gclk));
	jdff dff_B_IbgITdg02_1(.din(n394),.dout(w_dff_B_IbgITdg02_1),.clk(gclk));
	jdff dff_B_ZGnttdhf7_1(.din(w_dff_B_IbgITdg02_1),.dout(w_dff_B_ZGnttdhf7_1),.clk(gclk));
	jdff dff_B_FTnw3Xg31_1(.din(w_dff_B_ZGnttdhf7_1),.dout(w_dff_B_FTnw3Xg31_1),.clk(gclk));
	jdff dff_B_LmGYBlcJ0_1(.din(w_dff_B_FTnw3Xg31_1),.dout(w_dff_B_LmGYBlcJ0_1),.clk(gclk));
	jdff dff_B_hm38KX6z5_1(.din(w_dff_B_LmGYBlcJ0_1),.dout(w_dff_B_hm38KX6z5_1),.clk(gclk));
	jdff dff_B_GCOT9CSH3_1(.din(w_dff_B_hm38KX6z5_1),.dout(w_dff_B_GCOT9CSH3_1),.clk(gclk));
	jdff dff_B_RLzrZUL35_1(.din(w_dff_B_GCOT9CSH3_1),.dout(w_dff_B_RLzrZUL35_1),.clk(gclk));
	jdff dff_B_t14rLGUG9_1(.din(w_dff_B_RLzrZUL35_1),.dout(w_dff_B_t14rLGUG9_1),.clk(gclk));
	jdff dff_B_5ONNJ2aR7_1(.din(w_dff_B_t14rLGUG9_1),.dout(w_dff_B_5ONNJ2aR7_1),.clk(gclk));
	jdff dff_B_dFO8mxsd2_1(.din(w_dff_B_5ONNJ2aR7_1),.dout(w_dff_B_dFO8mxsd2_1),.clk(gclk));
	jdff dff_B_w1bw6mgr0_1(.din(w_dff_B_dFO8mxsd2_1),.dout(w_dff_B_w1bw6mgr0_1),.clk(gclk));
	jdff dff_B_BudxxYAP4_0(.din(n396),.dout(w_dff_B_BudxxYAP4_0),.clk(gclk));
	jdff dff_B_itO9ESq70_0(.din(w_dff_B_BudxxYAP4_0),.dout(w_dff_B_itO9ESq70_0),.clk(gclk));
	jdff dff_B_uGzVBG4I4_0(.din(w_dff_B_itO9ESq70_0),.dout(w_dff_B_uGzVBG4I4_0),.clk(gclk));
	jdff dff_B_Eonx0fjG8_0(.din(w_dff_B_uGzVBG4I4_0),.dout(w_dff_B_Eonx0fjG8_0),.clk(gclk));
	jdff dff_B_z7ThNTPj4_0(.din(w_dff_B_Eonx0fjG8_0),.dout(w_dff_B_z7ThNTPj4_0),.clk(gclk));
	jdff dff_B_jJaHR3sF9_0(.din(w_dff_B_z7ThNTPj4_0),.dout(w_dff_B_jJaHR3sF9_0),.clk(gclk));
	jdff dff_B_87zgBDTl8_0(.din(w_dff_B_jJaHR3sF9_0),.dout(w_dff_B_87zgBDTl8_0),.clk(gclk));
	jdff dff_B_PW4upquJ9_0(.din(w_dff_B_87zgBDTl8_0),.dout(w_dff_B_PW4upquJ9_0),.clk(gclk));
	jdff dff_B_kEp2i10w6_0(.din(w_dff_B_PW4upquJ9_0),.dout(w_dff_B_kEp2i10w6_0),.clk(gclk));
	jdff dff_B_cZCIEIF56_0(.din(w_dff_B_kEp2i10w6_0),.dout(w_dff_B_cZCIEIF56_0),.clk(gclk));
	jdff dff_B_tw1vjor82_0(.din(w_dff_B_cZCIEIF56_0),.dout(w_dff_B_tw1vjor82_0),.clk(gclk));
	jdff dff_B_Ad4et2Xi9_0(.din(w_dff_B_tw1vjor82_0),.dout(w_dff_B_Ad4et2Xi9_0),.clk(gclk));
	jdff dff_B_oS7eGAiL7_0(.din(w_dff_B_Ad4et2Xi9_0),.dout(w_dff_B_oS7eGAiL7_0),.clk(gclk));
	jdff dff_B_CC303Aux6_0(.din(w_dff_B_oS7eGAiL7_0),.dout(w_dff_B_CC303Aux6_0),.clk(gclk));
	jdff dff_A_43sdw0E60_0(.dout(w_n395_0[0]),.din(w_dff_A_43sdw0E60_0),.clk(gclk));
	jdff dff_A_b6tgVJP91_0(.dout(w_dff_A_43sdw0E60_0),.din(w_dff_A_b6tgVJP91_0),.clk(gclk));
	jdff dff_A_9uWz4vrr6_0(.dout(w_dff_A_b6tgVJP91_0),.din(w_dff_A_9uWz4vrr6_0),.clk(gclk));
	jdff dff_A_38kW0dit4_0(.dout(w_dff_A_9uWz4vrr6_0),.din(w_dff_A_38kW0dit4_0),.clk(gclk));
	jdff dff_A_VUERVbxm0_0(.dout(w_dff_A_38kW0dit4_0),.din(w_dff_A_VUERVbxm0_0),.clk(gclk));
	jdff dff_A_1Xtr9VzC5_0(.dout(w_dff_A_VUERVbxm0_0),.din(w_dff_A_1Xtr9VzC5_0),.clk(gclk));
	jdff dff_A_L4eWfhTE0_0(.dout(w_dff_A_1Xtr9VzC5_0),.din(w_dff_A_L4eWfhTE0_0),.clk(gclk));
	jdff dff_A_6u4U92tJ6_0(.dout(w_dff_A_L4eWfhTE0_0),.din(w_dff_A_6u4U92tJ6_0),.clk(gclk));
	jdff dff_A_Xtjrrr5O5_0(.dout(w_dff_A_6u4U92tJ6_0),.din(w_dff_A_Xtjrrr5O5_0),.clk(gclk));
	jdff dff_A_AhSpaSA57_0(.dout(w_dff_A_Xtjrrr5O5_0),.din(w_dff_A_AhSpaSA57_0),.clk(gclk));
	jdff dff_A_cS1gB5A59_0(.dout(w_dff_A_AhSpaSA57_0),.din(w_dff_A_cS1gB5A59_0),.clk(gclk));
	jdff dff_A_IUbjxoHp6_0(.dout(w_dff_A_cS1gB5A59_0),.din(w_dff_A_IUbjxoHp6_0),.clk(gclk));
	jdff dff_A_h3E7MLZb8_0(.dout(w_dff_A_IUbjxoHp6_0),.din(w_dff_A_h3E7MLZb8_0),.clk(gclk));
	jdff dff_A_whmcJS1k6_0(.dout(w_dff_A_h3E7MLZb8_0),.din(w_dff_A_whmcJS1k6_0),.clk(gclk));
	jdff dff_A_hvRrNjYK1_0(.dout(w_dff_A_whmcJS1k6_0),.din(w_dff_A_hvRrNjYK1_0),.clk(gclk));
	jdff dff_B_2X76qvum3_0(.din(n329),.dout(w_dff_B_2X76qvum3_0),.clk(gclk));
	jdff dff_B_C3EU4oge3_0(.din(n323),.dout(w_dff_B_C3EU4oge3_0),.clk(gclk));
	jdff dff_A_Gsyd0ard9_1(.dout(w_n189_0[1]),.din(w_dff_A_Gsyd0ard9_1),.clk(gclk));
	jdff dff_A_L6U6GY1b4_1(.dout(w_dff_A_Gsyd0ard9_1),.din(w_dff_A_L6U6GY1b4_1),.clk(gclk));
	jdff dff_B_JiY5AdFT7_2(.din(n318),.dout(w_dff_B_JiY5AdFT7_2),.clk(gclk));
	jdff dff_A_VjUM8A8S1_1(.dout(w_n185_0[1]),.din(w_dff_A_VjUM8A8S1_1),.clk(gclk));
	jdff dff_A_BAYoBgXK4_1(.dout(w_dff_A_VjUM8A8S1_1),.din(w_dff_A_BAYoBgXK4_1),.clk(gclk));
	jdff dff_A_tczWpGTT9_2(.dout(w_n185_0[2]),.din(w_dff_A_tczWpGTT9_2),.clk(gclk));
	jdff dff_A_LGKbteRn7_2(.dout(w_dff_A_tczWpGTT9_2),.din(w_dff_A_LGKbteRn7_2),.clk(gclk));
	jdff dff_B_rWeVQahk1_3(.din(n184),.dout(w_dff_B_rWeVQahk1_3),.clk(gclk));
	jdff dff_B_qYuHsMCP9_3(.din(w_dff_B_rWeVQahk1_3),.dout(w_dff_B_qYuHsMCP9_3),.clk(gclk));
	jdff dff_A_JKWe0tgd8_0(.dout(w_n314_0[0]),.din(w_dff_A_JKWe0tgd8_0),.clk(gclk));
	jdff dff_A_kPgkeHL59_1(.dout(w_n314_0[1]),.din(w_dff_A_kPgkeHL59_1),.clk(gclk));
	jdff dff_B_UkXvgx952_3(.din(n314),.dout(w_dff_B_UkXvgx952_3),.clk(gclk));
	jdff dff_A_9zwH7vGq2_1(.dout(w_n311_0[1]),.din(w_dff_A_9zwH7vGq2_1),.clk(gclk));
	jdff dff_A_Y3bjhKXk0_2(.dout(w_n311_0[2]),.din(w_dff_A_Y3bjhKXk0_2),.clk(gclk));
	jdff dff_B_4fbkGuta1_3(.din(n311),.dout(w_dff_B_4fbkGuta1_3),.clk(gclk));
	jdff dff_A_OwPFPiKc9_0(.dout(w_n183_0[0]),.din(w_dff_A_OwPFPiKc9_0),.clk(gclk));
	jdff dff_A_D38mq5HD8_0(.dout(w_dff_A_OwPFPiKc9_0),.din(w_dff_A_D38mq5HD8_0),.clk(gclk));
	jdff dff_A_lHFT4Hzt1_0(.dout(w_dff_A_D38mq5HD8_0),.din(w_dff_A_lHFT4Hzt1_0),.clk(gclk));
	jdff dff_A_IXDKr6J37_1(.dout(w_n183_0[1]),.din(w_dff_A_IXDKr6J37_1),.clk(gclk));
	jdff dff_A_twt0QH2O9_1(.dout(w_dff_A_IXDKr6J37_1),.din(w_dff_A_twt0QH2O9_1),.clk(gclk));
	jdff dff_A_eQpI6Izx1_1(.dout(w_dff_A_twt0QH2O9_1),.din(w_dff_A_eQpI6Izx1_1),.clk(gclk));
	jdff dff_B_kw3WVZKl4_0(.din(n182),.dout(w_dff_B_kw3WVZKl4_0),.clk(gclk));
	jdff dff_B_dJvBFtKS2_1(.din(G900),.dout(w_dff_B_dJvBFtKS2_1),.clk(gclk));
	jdff dff_B_RWWx8zwf9_0(.din(n304),.dout(w_dff_B_RWWx8zwf9_0),.clk(gclk));
	jdff dff_A_cevCT52N3_1(.dout(w_n188_0[1]),.din(w_dff_A_cevCT52N3_1),.clk(gclk));
	jdff dff_A_09aFEYq23_0(.dout(w_n290_0[0]),.din(w_dff_A_09aFEYq23_0),.clk(gclk));
	jdff dff_B_tW00DcSv5_3(.din(n290),.dout(w_dff_B_tW00DcSv5_3),.clk(gclk));
	jdff dff_A_fp2xXihd8_0(.dout(w_n289_0[0]),.din(w_dff_A_fp2xXihd8_0),.clk(gclk));
	jdff dff_A_35cPAWIb4_0(.dout(w_dff_A_fp2xXihd8_0),.din(w_dff_A_35cPAWIb4_0),.clk(gclk));
	jdff dff_B_Usf5N05v7_3(.din(n158),.dout(w_dff_B_Usf5N05v7_3),.clk(gclk));
	jdff dff_A_G8WUL3kv2_0(.dout(w_n92_1[0]),.din(w_dff_A_G8WUL3kv2_0),.clk(gclk));
	jdff dff_A_ZGKCYnYR1_0(.dout(w_dff_A_G8WUL3kv2_0),.din(w_dff_A_ZGKCYnYR1_0),.clk(gclk));
	jdff dff_A_wYupysZH7_2(.dout(w_n92_1[2]),.din(w_dff_A_wYupysZH7_2),.clk(gclk));
	jdff dff_A_rjUC9ARk0_2(.dout(w_dff_A_wYupysZH7_2),.din(w_dff_A_rjUC9ARk0_2),.clk(gclk));
	jdff dff_B_QNQfbk5n1_2(.din(n286),.dout(w_dff_B_QNQfbk5n1_2),.clk(gclk));
	jdff dff_A_77YZnQFx6_1(.dout(w_n163_0[1]),.din(w_dff_A_77YZnQFx6_1),.clk(gclk));
	jdff dff_A_EaD5zzkl9_1(.dout(w_dff_A_77YZnQFx6_1),.din(w_dff_A_EaD5zzkl9_1),.clk(gclk));
	jdff dff_A_y4Ea0X3n9_2(.dout(w_n163_0[2]),.din(w_dff_A_y4Ea0X3n9_2),.clk(gclk));
	jdff dff_A_0mBEjIpT3_2(.dout(w_dff_A_y4Ea0X3n9_2),.din(w_dff_A_0mBEjIpT3_2),.clk(gclk));
	jdff dff_B_n7nSzbcp3_1(.din(n123),.dout(w_dff_B_n7nSzbcp3_1),.clk(gclk));
	jdff dff_B_vdpK5TU17_1(.din(w_dff_B_n7nSzbcp3_1),.dout(w_dff_B_vdpK5TU17_1),.clk(gclk));
	jdff dff_B_WZEIPPf01_1(.din(w_dff_B_vdpK5TU17_1),.dout(w_dff_B_WZEIPPf01_1),.clk(gclk));
	jdff dff_B_GZ9zm3sP0_1(.din(w_dff_B_WZEIPPf01_1),.dout(w_dff_B_GZ9zm3sP0_1),.clk(gclk));
	jdff dff_B_8YJPDxz80_1(.din(w_dff_B_GZ9zm3sP0_1),.dout(w_dff_B_8YJPDxz80_1),.clk(gclk));
	jdff dff_A_y3JAZ3pi5_0(.dout(w_n68_0[0]),.din(w_dff_A_y3JAZ3pi5_0),.clk(gclk));
	jdff dff_A_Ku2msB4J4_0(.dout(w_dff_A_y3JAZ3pi5_0),.din(w_dff_A_Ku2msB4J4_0),.clk(gclk));
	jdff dff_A_TKKxVdUJ6_0(.dout(w_dff_A_Ku2msB4J4_0),.din(w_dff_A_TKKxVdUJ6_0),.clk(gclk));
	jdff dff_A_RjJxRump3_0(.dout(w_dff_A_TKKxVdUJ6_0),.din(w_dff_A_RjJxRump3_0),.clk(gclk));
	jdff dff_A_ntig2NOL4_0(.dout(w_dff_A_RjJxRump3_0),.din(w_dff_A_ntig2NOL4_0),.clk(gclk));
	jdff dff_A_EQ0PWSxH9_0(.dout(w_dff_A_ntig2NOL4_0),.din(w_dff_A_EQ0PWSxH9_0),.clk(gclk));
	jdff dff_A_Yh7r2zhx9_0(.dout(w_dff_A_EQ0PWSxH9_0),.din(w_dff_A_Yh7r2zhx9_0),.clk(gclk));
	jdff dff_A_6DIvp8LB3_0(.dout(w_dff_A_Yh7r2zhx9_0),.din(w_dff_A_6DIvp8LB3_0),.clk(gclk));
	jdff dff_A_ZK6n7x4R7_0(.dout(w_dff_A_6DIvp8LB3_0),.din(w_dff_A_ZK6n7x4R7_0),.clk(gclk));
	jdff dff_A_TZpe6yX65_0(.dout(w_dff_A_ZK6n7x4R7_0),.din(w_dff_A_TZpe6yX65_0),.clk(gclk));
	jdff dff_A_tCNaVkta5_0(.dout(w_n281_0[0]),.din(w_dff_A_tCNaVkta5_0),.clk(gclk));
	jdff dff_A_tfIY17mv0_1(.dout(w_n281_0[1]),.din(w_dff_A_tfIY17mv0_1),.clk(gclk));
	jdff dff_B_4HOjDZJ16_3(.din(n281),.dout(w_dff_B_4HOjDZJ16_3),.clk(gclk));
	jdff dff_B_WJSuNHrv7_2(.din(n278),.dout(w_dff_B_WJSuNHrv7_2),.clk(gclk));
	jdff dff_A_cN8fX8Sm1_1(.dout(w_n168_0[1]),.din(w_dff_A_cN8fX8Sm1_1),.clk(gclk));
	jdff dff_A_uybc2Yyp3_1(.dout(w_dff_A_cN8fX8Sm1_1),.din(w_dff_A_uybc2Yyp3_1),.clk(gclk));
	jdff dff_A_6VFVOl7i4_2(.dout(w_n168_0[2]),.din(w_dff_A_6VFVOl7i4_2),.clk(gclk));
	jdff dff_A_OeuzmHsY5_2(.dout(w_dff_A_6VFVOl7i4_2),.din(w_dff_A_OeuzmHsY5_2),.clk(gclk));
	jdff dff_B_KIRixJ3S5_1(.din(n133),.dout(w_dff_B_KIRixJ3S5_1),.clk(gclk));
	jdff dff_B_32uTggt32_1(.din(w_dff_B_KIRixJ3S5_1),.dout(w_dff_B_32uTggt32_1),.clk(gclk));
	jdff dff_B_mE7RG9PU7_1(.din(w_dff_B_32uTggt32_1),.dout(w_dff_B_mE7RG9PU7_1),.clk(gclk));
	jdff dff_B_5LKhvowI7_1(.din(w_dff_B_mE7RG9PU7_1),.dout(w_dff_B_5LKhvowI7_1),.clk(gclk));
	jdff dff_B_GPN843GF3_1(.din(w_dff_B_5LKhvowI7_1),.dout(w_dff_B_GPN843GF3_1),.clk(gclk));
	jdff dff_A_12kEBCe27_0(.dout(w_n141_0[0]),.din(w_dff_A_12kEBCe27_0),.clk(gclk));
	jdff dff_A_kUCrtOgj9_0(.dout(w_dff_A_12kEBCe27_0),.din(w_dff_A_kUCrtOgj9_0),.clk(gclk));
	jdff dff_A_fvXBlzga2_0(.dout(w_dff_A_kUCrtOgj9_0),.din(w_dff_A_fvXBlzga2_0),.clk(gclk));
	jdff dff_A_ZxNX1Sgr7_0(.dout(w_dff_A_fvXBlzga2_0),.din(w_dff_A_ZxNX1Sgr7_0),.clk(gclk));
	jdff dff_A_Y5zLzirL6_0(.dout(w_dff_A_ZxNX1Sgr7_0),.din(w_dff_A_Y5zLzirL6_0),.clk(gclk));
	jdff dff_A_sSbSow6S9_0(.dout(w_dff_A_Y5zLzirL6_0),.din(w_dff_A_sSbSow6S9_0),.clk(gclk));
	jdff dff_A_WYtAyPVj2_0(.dout(w_dff_A_sSbSow6S9_0),.din(w_dff_A_WYtAyPVj2_0),.clk(gclk));
	jdff dff_A_U4AwMOeS9_0(.dout(w_dff_A_WYtAyPVj2_0),.din(w_dff_A_U4AwMOeS9_0),.clk(gclk));
	jdff dff_A_iYSgMOEl1_0(.dout(w_dff_A_U4AwMOeS9_0),.din(w_dff_A_iYSgMOEl1_0),.clk(gclk));
	jdff dff_A_mpKgBLlT0_0(.dout(w_dff_A_iYSgMOEl1_0),.din(w_dff_A_mpKgBLlT0_0),.clk(gclk));
	jdff dff_A_lx7CktvA6_0(.dout(w_dff_A_mpKgBLlT0_0),.din(w_dff_A_lx7CktvA6_0),.clk(gclk));
	jdff dff_A_r5bBon7e8_0(.dout(w_dff_A_lx7CktvA6_0),.din(w_dff_A_r5bBon7e8_0),.clk(gclk));
	jdff dff_B_10Srcflh0_1(.din(n134),.dout(w_dff_B_10Srcflh0_1),.clk(gclk));
	jdff dff_B_FqQKqgp44_1(.din(w_dff_B_10Srcflh0_1),.dout(w_dff_B_FqQKqgp44_1),.clk(gclk));
	jdff dff_A_xJEj469K2_1(.dout(w_G475_0[1]),.din(w_dff_A_xJEj469K2_1),.clk(gclk));
	jdff dff_A_3ZHx4Sfa5_1(.dout(w_dff_A_xJEj469K2_1),.din(w_dff_A_3ZHx4Sfa5_1),.clk(gclk));
	jdff dff_A_z3SmD95q2_1(.dout(w_dff_A_3ZHx4Sfa5_1),.din(w_dff_A_z3SmD95q2_1),.clk(gclk));
	jdff dff_A_V1PZESwJ4_1(.dout(w_dff_A_z3SmD95q2_1),.din(w_dff_A_V1PZESwJ4_1),.clk(gclk));
	jdff dff_A_cDqW9WV37_1(.dout(w_dff_A_V1PZESwJ4_1),.din(w_dff_A_cDqW9WV37_1),.clk(gclk));
	jdff dff_A_Fen5hBPN4_1(.dout(w_dff_A_cDqW9WV37_1),.din(w_dff_A_Fen5hBPN4_1),.clk(gclk));
	jdff dff_A_Dk9wjD6R1_0(.dout(w_n130_0[0]),.din(w_dff_A_Dk9wjD6R1_0),.clk(gclk));
	jdff dff_A_fb8SYfc44_0(.dout(w_dff_A_Dk9wjD6R1_0),.din(w_dff_A_fb8SYfc44_0),.clk(gclk));
	jdff dff_A_oovHH2GY4_0(.dout(w_dff_A_fb8SYfc44_0),.din(w_dff_A_oovHH2GY4_0),.clk(gclk));
	jdff dff_A_uqCwlZHn5_0(.dout(w_dff_A_oovHH2GY4_0),.din(w_dff_A_uqCwlZHn5_0),.clk(gclk));
	jdff dff_A_bn6iy4Lk7_0(.dout(w_dff_A_uqCwlZHn5_0),.din(w_dff_A_bn6iy4Lk7_0),.clk(gclk));
	jdff dff_A_s5dsEzNe8_0(.dout(w_dff_A_bn6iy4Lk7_0),.din(w_dff_A_s5dsEzNe8_0),.clk(gclk));
	jdff dff_A_9LlXIY4a1_0(.dout(w_dff_A_s5dsEzNe8_0),.din(w_dff_A_9LlXIY4a1_0),.clk(gclk));
	jdff dff_A_4lE5uAY26_0(.dout(w_dff_A_9LlXIY4a1_0),.din(w_dff_A_4lE5uAY26_0),.clk(gclk));
	jdff dff_A_4nBtkBNO7_0(.dout(w_dff_A_4lE5uAY26_0),.din(w_dff_A_4nBtkBNO7_0),.clk(gclk));
	jdff dff_A_Bpjc5yAZ6_0(.dout(w_dff_A_4nBtkBNO7_0),.din(w_dff_A_Bpjc5yAZ6_0),.clk(gclk));
	jdff dff_A_mJFUkyte8_0(.dout(w_dff_A_Bpjc5yAZ6_0),.din(w_dff_A_mJFUkyte8_0),.clk(gclk));
	jdff dff_A_7abemTm64_0(.dout(w_dff_A_mJFUkyte8_0),.din(w_dff_A_7abemTm64_0),.clk(gclk));
	jdff dff_B_RPK2d2Xf7_1(.din(n124),.dout(w_dff_B_RPK2d2Xf7_1),.clk(gclk));
	jdff dff_B_SNUMfQmR4_1(.din(w_dff_B_RPK2d2Xf7_1),.dout(w_dff_B_SNUMfQmR4_1),.clk(gclk));
	jdff dff_B_bnwWeJ3A0_1(.din(w_dff_B_SNUMfQmR4_1),.dout(w_dff_B_bnwWeJ3A0_1),.clk(gclk));
	jdff dff_B_uMxwGq9V4_0(.din(n128),.dout(w_dff_B_uMxwGq9V4_0),.clk(gclk));
	jdff dff_A_2wfAFn5J6_1(.dout(w_G478_0[1]),.din(w_dff_A_2wfAFn5J6_1),.clk(gclk));
	jdff dff_A_n8GTCpjy9_1(.dout(w_dff_A_2wfAFn5J6_1),.din(w_dff_A_n8GTCpjy9_1),.clk(gclk));
	jdff dff_A_yjmL5mQE3_1(.dout(w_dff_A_n8GTCpjy9_1),.din(w_dff_A_yjmL5mQE3_1),.clk(gclk));
	jdff dff_A_iHAj7Unf4_1(.dout(w_dff_A_yjmL5mQE3_1),.din(w_dff_A_iHAj7Unf4_1),.clk(gclk));
	jdff dff_A_q5UWtISA6_1(.dout(w_dff_A_iHAj7Unf4_1),.din(w_dff_A_q5UWtISA6_1),.clk(gclk));
	jdff dff_A_P8vhbcLd3_1(.dout(w_dff_A_q5UWtISA6_1),.din(w_dff_A_P8vhbcLd3_1),.clk(gclk));
	jdff dff_B_AsfZNo1y9_3(.din(n154),.dout(w_dff_B_AsfZNo1y9_3),.clk(gclk));
	jdff dff_B_F3v9r44p2_3(.din(w_dff_B_AsfZNo1y9_3),.dout(w_dff_B_F3v9r44p2_3),.clk(gclk));
	jdff dff_A_Gijw0raT3_0(.dout(w_n153_0[0]),.din(w_dff_A_Gijw0raT3_0),.clk(gclk));
	jdff dff_A_AyTXD4nA2_0(.dout(w_dff_A_Gijw0raT3_0),.din(w_dff_A_AyTXD4nA2_0),.clk(gclk));
	jdff dff_A_6OwQNu0J9_0(.dout(w_dff_A_AyTXD4nA2_0),.din(w_dff_A_6OwQNu0J9_0),.clk(gclk));
	jdff dff_A_pVs8Nnzn4_1(.dout(w_n153_0[1]),.din(w_dff_A_pVs8Nnzn4_1),.clk(gclk));
	jdff dff_A_04XLNkTB3_1(.dout(w_dff_A_pVs8Nnzn4_1),.din(w_dff_A_04XLNkTB3_1),.clk(gclk));
	jdff dff_A_Z17idjTY7_1(.dout(w_dff_A_04XLNkTB3_1),.din(w_dff_A_Z17idjTY7_1),.clk(gclk));
	jdff dff_B_gqqmwf5n4_1(.din(n148),.dout(w_dff_B_gqqmwf5n4_1),.clk(gclk));
	jdff dff_A_PkEGoEvi6_0(.dout(w_n151_0[0]),.din(w_dff_A_PkEGoEvi6_0),.clk(gclk));
	jdff dff_A_uJhzAsOt0_1(.dout(w_n151_0[1]),.din(w_dff_A_uJhzAsOt0_1),.clk(gclk));
	jdff dff_A_aYurxw2I2_1(.dout(w_dff_A_uJhzAsOt0_1),.din(w_dff_A_aYurxw2I2_1),.clk(gclk));
	jdff dff_A_igt5OodG1_1(.dout(w_dff_A_aYurxw2I2_1),.din(w_dff_A_igt5OodG1_1),.clk(gclk));
	jdff dff_A_rDsavkC15_1(.dout(w_dff_A_igt5OodG1_1),.din(w_dff_A_rDsavkC15_1),.clk(gclk));
	jdff dff_A_amWPkPxt1_1(.dout(w_dff_A_rDsavkC15_1),.din(w_dff_A_amWPkPxt1_1),.clk(gclk));
	jdff dff_A_x3wg5B3h8_1(.dout(w_dff_A_amWPkPxt1_1),.din(w_dff_A_x3wg5B3h8_1),.clk(gclk));
	jdff dff_A_PVbXV4xh1_1(.dout(w_dff_A_x3wg5B3h8_1),.din(w_dff_A_PVbXV4xh1_1),.clk(gclk));
	jdff dff_A_3FL4wCib1_1(.dout(w_dff_A_PVbXV4xh1_1),.din(w_dff_A_3FL4wCib1_1),.clk(gclk));
	jdff dff_A_XJhtk5d93_1(.dout(w_dff_A_3FL4wCib1_1),.din(w_dff_A_XJhtk5d93_1),.clk(gclk));
	jdff dff_A_HgB1EC1h4_1(.dout(w_dff_A_XJhtk5d93_1),.din(w_dff_A_HgB1EC1h4_1),.clk(gclk));
	jdff dff_A_rmgtX48U8_1(.dout(w_dff_A_HgB1EC1h4_1),.din(w_dff_A_rmgtX48U8_1),.clk(gclk));
	jdff dff_A_skdxaJlv5_1(.dout(w_G952_0[1]),.din(w_dff_A_skdxaJlv5_1),.clk(gclk));
	jdff dff_A_sOYhJJgj6_1(.dout(w_dff_A_skdxaJlv5_1),.din(w_dff_A_sOYhJJgj6_1),.clk(gclk));
	jdff dff_A_V62iRMJi4_1(.dout(w_dff_A_sOYhJJgj6_1),.din(w_dff_A_V62iRMJi4_1),.clk(gclk));
	jdff dff_A_883NNCTR0_1(.dout(w_dff_A_V62iRMJi4_1),.din(w_dff_A_883NNCTR0_1),.clk(gclk));
	jdff dff_A_8uRKuM9I3_1(.dout(w_dff_A_883NNCTR0_1),.din(w_dff_A_8uRKuM9I3_1),.clk(gclk));
	jdff dff_A_6XMG2iQb1_1(.dout(w_dff_A_8uRKuM9I3_1),.din(w_dff_A_6XMG2iQb1_1),.clk(gclk));
	jdff dff_A_Felw4Quu8_1(.dout(w_dff_A_6XMG2iQb1_1),.din(w_dff_A_Felw4Quu8_1),.clk(gclk));
	jdff dff_A_2ZQnkBe39_1(.dout(w_dff_A_Felw4Quu8_1),.din(w_dff_A_2ZQnkBe39_1),.clk(gclk));
	jdff dff_A_ioZ7jfd93_1(.dout(w_dff_A_2ZQnkBe39_1),.din(w_dff_A_ioZ7jfd93_1),.clk(gclk));
	jdff dff_A_OybXhudh7_1(.dout(w_dff_A_ioZ7jfd93_1),.din(w_dff_A_OybXhudh7_1),.clk(gclk));
	jdff dff_A_QS98rDnB1_1(.dout(w_dff_A_OybXhudh7_1),.din(w_dff_A_QS98rDnB1_1),.clk(gclk));
	jdff dff_A_t1Ra9Q1I7_1(.dout(w_dff_A_QS98rDnB1_1),.din(w_dff_A_t1Ra9Q1I7_1),.clk(gclk));
	jdff dff_A_401pkTmY4_1(.dout(w_dff_A_t1Ra9Q1I7_1),.din(w_dff_A_401pkTmY4_1),.clk(gclk));
	jdff dff_A_BdPtsxom3_1(.dout(w_dff_A_401pkTmY4_1),.din(w_dff_A_BdPtsxom3_1),.clk(gclk));
	jdff dff_A_d75WGEe48_1(.dout(w_dff_A_BdPtsxom3_1),.din(w_dff_A_d75WGEe48_1),.clk(gclk));
	jdff dff_A_GL5TIQ7d7_1(.dout(w_dff_A_d75WGEe48_1),.din(w_dff_A_GL5TIQ7d7_1),.clk(gclk));
	jdff dff_B_aqHRAwgz1_3(.din(G952),.dout(w_dff_B_aqHRAwgz1_3),.clk(gclk));
	jdff dff_B_nVa2DG5s9_1(.din(G898),.dout(w_dff_B_nVa2DG5s9_1),.clk(gclk));
	jdff dff_A_ZalKv5WY2_2(.dout(w_n253_0[2]),.din(w_dff_A_ZalKv5WY2_2),.clk(gclk));
	jdff dff_A_1P4uAqKF2_1(.dout(w_n92_0[1]),.din(w_dff_A_1P4uAqKF2_1),.clk(gclk));
	jdff dff_A_WuJ6cgDg8_1(.dout(w_dff_A_1P4uAqKF2_1),.din(w_dff_A_WuJ6cgDg8_1),.clk(gclk));
	jdff dff_A_jeN1wdfO5_2(.dout(w_n92_0[2]),.din(w_dff_A_jeN1wdfO5_2),.clk(gclk));
	jdff dff_A_afyGrk4u3_2(.dout(w_dff_A_jeN1wdfO5_2),.din(w_dff_A_afyGrk4u3_2),.clk(gclk));
	jdff dff_A_lWolemKd3_1(.dout(w_G472_0[1]),.din(w_dff_A_lWolemKd3_1),.clk(gclk));
	jdff dff_A_zDWHIrcy1_1(.dout(w_dff_A_lWolemKd3_1),.din(w_dff_A_zDWHIrcy1_1),.clk(gclk));
	jdff dff_A_WQXVwCaB7_1(.dout(w_dff_A_zDWHIrcy1_1),.din(w_dff_A_WQXVwCaB7_1),.clk(gclk));
	jdff dff_A_syEcHXZs1_1(.dout(w_dff_A_WQXVwCaB7_1),.din(w_dff_A_syEcHXZs1_1),.clk(gclk));
	jdff dff_A_MNtjag3F5_1(.dout(w_dff_A_syEcHXZs1_1),.din(w_dff_A_MNtjag3F5_1),.clk(gclk));
	jdff dff_A_hOgoEuEd3_1(.dout(w_dff_A_MNtjag3F5_1),.din(w_dff_A_hOgoEuEd3_1),.clk(gclk));
	jdff dff_B_09PlH9TX2_2(.din(n73),.dout(w_dff_B_09PlH9TX2_2),.clk(gclk));
	jdff dff_B_u4VfuVjA8_2(.din(w_dff_B_09PlH9TX2_2),.dout(w_dff_B_u4VfuVjA8_2),.clk(gclk));
	jdff dff_B_mGhgz6K78_2(.din(w_dff_B_u4VfuVjA8_2),.dout(w_dff_B_mGhgz6K78_2),.clk(gclk));
	jdff dff_B_WBIUpuZz2_2(.din(w_dff_B_mGhgz6K78_2),.dout(w_dff_B_WBIUpuZz2_2),.clk(gclk));
	jdff dff_A_f1Cp3bG98_1(.dout(w_G217_0[1]),.din(w_dff_A_f1Cp3bG98_1),.clk(gclk));
	jdff dff_A_tvjJs3Tl8_1(.dout(w_dff_A_f1Cp3bG98_1),.din(w_dff_A_tvjJs3Tl8_1),.clk(gclk));
	jdff dff_A_4HiJw4826_2(.dout(w_G217_0[2]),.din(w_dff_A_4HiJw4826_2),.clk(gclk));
	jdff dff_A_oGL2QCwY7_2(.dout(w_dff_A_4HiJw4826_2),.din(w_dff_A_oGL2QCwY7_2),.clk(gclk));
	jdff dff_A_QbcyzIER2_2(.dout(w_dff_A_oGL2QCwY7_2),.din(w_dff_A_QbcyzIER2_2),.clk(gclk));
	jdff dff_A_KBqT75Wh0_0(.dout(w_n172_0[0]),.din(w_dff_A_KBqT75Wh0_0),.clk(gclk));
	jdff dff_A_rAfPXC9K6_0(.dout(w_dff_A_KBqT75Wh0_0),.din(w_dff_A_rAfPXC9K6_0),.clk(gclk));
	jdff dff_A_NWX2EhTo2_0(.dout(w_dff_A_rAfPXC9K6_0),.din(w_dff_A_NWX2EhTo2_0),.clk(gclk));
	jdff dff_A_LsCdbSGK0_0(.dout(w_dff_A_NWX2EhTo2_0),.din(w_dff_A_LsCdbSGK0_0),.clk(gclk));
	jdff dff_A_e2ipIjke8_0(.dout(w_dff_A_LsCdbSGK0_0),.din(w_dff_A_e2ipIjke8_0),.clk(gclk));
	jdff dff_A_yjeGonY34_0(.dout(w_dff_A_e2ipIjke8_0),.din(w_dff_A_yjeGonY34_0),.clk(gclk));
	jdff dff_A_ooqiek5u7_0(.dout(w_dff_A_yjeGonY34_0),.din(w_dff_A_ooqiek5u7_0),.clk(gclk));
	jdff dff_A_J9Kye0S65_0(.dout(w_dff_A_ooqiek5u7_0),.din(w_dff_A_J9Kye0S65_0),.clk(gclk));
	jdff dff_A_yWU1yxgg9_0(.dout(w_dff_A_J9Kye0S65_0),.din(w_dff_A_yWU1yxgg9_0),.clk(gclk));
	jdff dff_A_tyPWgfYn3_0(.dout(w_dff_A_yWU1yxgg9_0),.din(w_dff_A_tyPWgfYn3_0),.clk(gclk));
	jdff dff_B_qVjn87qS0_1(.din(n171),.dout(w_dff_B_qVjn87qS0_1),.clk(gclk));
	jdff dff_B_NQdxbq4y2_1(.din(w_dff_B_qVjn87qS0_1),.dout(w_dff_B_NQdxbq4y2_1),.clk(gclk));
	jdff dff_B_9BtTOrGF3_1(.din(w_dff_B_NQdxbq4y2_1),.dout(w_dff_B_9BtTOrGF3_1),.clk(gclk));
	jdff dff_B_rV3lDE5L7_0(.din(n65),.dout(w_dff_B_rV3lDE5L7_0),.clk(gclk));
	jdff dff_B_CICOUOZh0_0(.din(w_dff_B_rV3lDE5L7_0),.dout(w_dff_B_CICOUOZh0_0),.clk(gclk));
	jdff dff_B_XDCpQqw55_0(.din(w_dff_B_CICOUOZh0_0),.dout(w_dff_B_XDCpQqw55_0),.clk(gclk));
	jdff dff_A_rVz5rJYr1_2(.dout(w_n60_0[2]),.din(w_dff_A_rVz5rJYr1_2),.clk(gclk));
	jdff dff_A_WkVPWE440_2(.dout(w_dff_A_rVz5rJYr1_2),.din(w_dff_A_WkVPWE440_2),.clk(gclk));
	jdff dff_A_sCpj0uGB3_2(.dout(w_dff_A_WkVPWE440_2),.din(w_dff_A_sCpj0uGB3_2),.clk(gclk));
	jdff dff_A_AWIT0A4U3_2(.dout(w_dff_A_sCpj0uGB3_2),.din(w_dff_A_AWIT0A4U3_2),.clk(gclk));
	jdff dff_A_D3arNb772_0(.dout(w_n59_0[0]),.din(w_dff_A_D3arNb772_0),.clk(gclk));
	jdff dff_A_0bAtBjHV7_0(.dout(w_dff_A_D3arNb772_0),.din(w_dff_A_0bAtBjHV7_0),.clk(gclk));
	jdff dff_A_IBtRA15N5_0(.dout(w_dff_A_0bAtBjHV7_0),.din(w_dff_A_IBtRA15N5_0),.clk(gclk));
	jdff dff_A_ooKg5vbG4_0(.dout(w_n70_1[0]),.din(w_dff_A_ooKg5vbG4_0),.clk(gclk));
	jdff dff_A_Hcm2yFCB9_0(.dout(w_dff_A_ooKg5vbG4_0),.din(w_dff_A_Hcm2yFCB9_0),.clk(gclk));
	jdff dff_A_Z03XvnuX8_0(.dout(w_dff_A_Hcm2yFCB9_0),.din(w_dff_A_Z03XvnuX8_0),.clk(gclk));
	jdff dff_A_zP5OBylv6_0(.dout(w_dff_A_Z03XvnuX8_0),.din(w_dff_A_zP5OBylv6_0),.clk(gclk));
	jdff dff_A_a6DH1R3z8_0(.dout(w_dff_A_zP5OBylv6_0),.din(w_dff_A_a6DH1R3z8_0),.clk(gclk));
	jdff dff_A_QzUmoGbW1_0(.dout(w_dff_A_a6DH1R3z8_0),.din(w_dff_A_QzUmoGbW1_0),.clk(gclk));
	jdff dff_A_nXlO4NRF3_2(.dout(w_n70_1[2]),.din(w_dff_A_nXlO4NRF3_2),.clk(gclk));
	jdff dff_A_6ggL88hA5_2(.dout(w_dff_A_nXlO4NRF3_2),.din(w_dff_A_6ggL88hA5_2),.clk(gclk));
	jdff dff_A_0haDp6k33_2(.dout(w_dff_A_6ggL88hA5_2),.din(w_dff_A_0haDp6k33_2),.clk(gclk));
	jdff dff_A_5pp87aYp3_2(.dout(w_dff_A_0haDp6k33_2),.din(w_dff_A_5pp87aYp3_2),.clk(gclk));
	jdff dff_A_kIPf5GNX7_0(.dout(w_n276_1[0]),.din(w_dff_A_kIPf5GNX7_0),.clk(gclk));
	jdff dff_B_kt5j7ogb8_3(.din(n276),.dout(w_dff_B_kt5j7ogb8_3),.clk(gclk));
	jdff dff_B_pUvsmUNx6_1(.din(n195),.dout(w_dff_B_pUvsmUNx6_1),.clk(gclk));
	jdff dff_B_hsa6jJmk4_1(.din(w_dff_B_pUvsmUNx6_1),.dout(w_dff_B_hsa6jJmk4_1),.clk(gclk));
	jdff dff_B_6090RKg83_1(.din(w_dff_B_hsa6jJmk4_1),.dout(w_dff_B_6090RKg83_1),.clk(gclk));
	jdff dff_B_RdqqFmKd0_1(.din(w_dff_B_6090RKg83_1),.dout(w_dff_B_RdqqFmKd0_1),.clk(gclk));
	jdff dff_B_vBQYwdZy1_1(.din(w_dff_B_RdqqFmKd0_1),.dout(w_dff_B_vBQYwdZy1_1),.clk(gclk));
	jdff dff_A_kn0O4zVs0_0(.dout(w_n117_0[0]),.din(w_dff_A_kn0O4zVs0_0),.clk(gclk));
	jdff dff_A_R0blMJvl1_0(.dout(w_dff_A_kn0O4zVs0_0),.din(w_dff_A_R0blMJvl1_0),.clk(gclk));
	jdff dff_A_0LejtOSm4_0(.dout(w_dff_A_R0blMJvl1_0),.din(w_dff_A_0LejtOSm4_0),.clk(gclk));
	jdff dff_A_3ddvpMdX2_0(.dout(w_dff_A_0LejtOSm4_0),.din(w_dff_A_3ddvpMdX2_0),.clk(gclk));
	jdff dff_A_7zX1W30Z2_0(.dout(w_dff_A_3ddvpMdX2_0),.din(w_dff_A_7zX1W30Z2_0),.clk(gclk));
	jdff dff_A_iBWULkw02_0(.dout(w_dff_A_7zX1W30Z2_0),.din(w_dff_A_iBWULkw02_0),.clk(gclk));
	jdff dff_A_1BSELLl67_0(.dout(w_dff_A_iBWULkw02_0),.din(w_dff_A_1BSELLl67_0),.clk(gclk));
	jdff dff_A_bwzxMwcl3_0(.dout(w_dff_A_1BSELLl67_0),.din(w_dff_A_bwzxMwcl3_0),.clk(gclk));
	jdff dff_A_xRohhYjS0_0(.dout(w_dff_A_bwzxMwcl3_0),.din(w_dff_A_xRohhYjS0_0),.clk(gclk));
	jdff dff_A_IwGUvFtv0_0(.dout(w_dff_A_xRohhYjS0_0),.din(w_dff_A_IwGUvFtv0_0),.clk(gclk));
	jdff dff_A_XuFJb69N5_0(.dout(w_dff_A_IwGUvFtv0_0),.din(w_dff_A_XuFJb69N5_0),.clk(gclk));
	jdff dff_A_GumpHgl86_0(.dout(w_dff_A_XuFJb69N5_0),.din(w_dff_A_GumpHgl86_0),.clk(gclk));
	jdff dff_B_17TASBNk7_1(.din(n113),.dout(w_dff_B_17TASBNk7_1),.clk(gclk));
	jdff dff_B_t4FDx38c5_1(.din(w_dff_B_17TASBNk7_1),.dout(w_dff_B_t4FDx38c5_1),.clk(gclk));
	jdff dff_B_ai20heMD3_2(.din(G227),.dout(w_dff_B_ai20heMD3_2),.clk(gclk));
	jdff dff_A_RCvN3C6T6_0(.dout(w_G140_0[0]),.din(w_dff_A_RCvN3C6T6_0),.clk(gclk));
	jdff dff_A_LxU2gbhj5_0(.dout(w_dff_A_RCvN3C6T6_0),.din(w_dff_A_LxU2gbhj5_0),.clk(gclk));
	jdff dff_A_NZsG0kcp6_0(.dout(w_dff_A_LxU2gbhj5_0),.din(w_dff_A_NZsG0kcp6_0),.clk(gclk));
	jdff dff_A_wRSzDpwI1_0(.dout(w_dff_A_NZsG0kcp6_0),.din(w_dff_A_wRSzDpwI1_0),.clk(gclk));
	jdff dff_A_PEN5enCk8_0(.dout(w_dff_A_wRSzDpwI1_0),.din(w_dff_A_PEN5enCk8_0),.clk(gclk));
	jdff dff_A_WcKIGJLU6_0(.dout(w_dff_A_PEN5enCk8_0),.din(w_dff_A_WcKIGJLU6_0),.clk(gclk));
	jdff dff_A_JPnXOuYs9_0(.dout(w_dff_A_WcKIGJLU6_0),.din(w_dff_A_JPnXOuYs9_0),.clk(gclk));
	jdff dff_A_djOLakeL8_0(.dout(w_dff_A_JPnXOuYs9_0),.din(w_dff_A_djOLakeL8_0),.clk(gclk));
	jdff dff_A_zIy1Pbin5_0(.dout(w_dff_A_djOLakeL8_0),.din(w_dff_A_zIy1Pbin5_0),.clk(gclk));
	jdff dff_A_LqNjbebR4_0(.dout(w_dff_A_zIy1Pbin5_0),.din(w_dff_A_LqNjbebR4_0),.clk(gclk));
	jdff dff_A_QJvkvlbc0_0(.dout(w_dff_A_LqNjbebR4_0),.din(w_dff_A_QJvkvlbc0_0),.clk(gclk));
	jdff dff_A_d4WkHQ0Z2_0(.dout(w_dff_A_QJvkvlbc0_0),.din(w_dff_A_d4WkHQ0Z2_0),.clk(gclk));
	jdff dff_A_hnfjFiB41_2(.dout(w_G469_0[2]),.din(w_dff_A_hnfjFiB41_2),.clk(gclk));
	jdff dff_A_t9pIzLeU2_2(.dout(w_dff_A_hnfjFiB41_2),.din(w_dff_A_t9pIzLeU2_2),.clk(gclk));
	jdff dff_A_VtLDsYHd1_2(.dout(w_dff_A_t9pIzLeU2_2),.din(w_dff_A_VtLDsYHd1_2),.clk(gclk));
	jdff dff_A_EKzrDLut8_2(.dout(w_dff_A_VtLDsYHd1_2),.din(w_dff_A_EKzrDLut8_2),.clk(gclk));
	jdff dff_A_vE3DRFNW5_2(.dout(w_dff_A_EKzrDLut8_2),.din(w_dff_A_vE3DRFNW5_2),.clk(gclk));
	jdff dff_A_cvbRW7X30_2(.dout(w_dff_A_vE3DRFNW5_2),.din(w_dff_A_cvbRW7X30_2),.clk(gclk));
	jdff dff_B_qVbzvNhX4_2(.din(n274),.dout(w_dff_B_qVbzvNhX4_2),.clk(gclk));
	jdff dff_B_nFtuYOEF5_2(.din(w_dff_B_qVbzvNhX4_2),.dout(w_dff_B_nFtuYOEF5_2),.clk(gclk));
	jdff dff_B_mINt9NCA2_2(.din(w_dff_B_nFtuYOEF5_2),.dout(w_dff_B_mINt9NCA2_2),.clk(gclk));
	jdff dff_A_zJEdtkcf1_0(.dout(w_n112_0[0]),.din(w_dff_A_zJEdtkcf1_0),.clk(gclk));
	jdff dff_A_JJm11C8A9_0(.dout(w_dff_A_zJEdtkcf1_0),.din(w_dff_A_JJm11C8A9_0),.clk(gclk));
	jdff dff_A_jeWGtTUG2_0(.dout(w_dff_A_JJm11C8A9_0),.din(w_dff_A_jeWGtTUG2_0),.clk(gclk));
	jdff dff_A_TKvJNnJd2_0(.dout(w_dff_A_jeWGtTUG2_0),.din(w_dff_A_TKvJNnJd2_0),.clk(gclk));
	jdff dff_B_DLUqT1wF5_1(.din(n111),.dout(w_dff_B_DLUqT1wF5_1),.clk(gclk));
	jdff dff_A_FzWSr4BD6_0(.dout(w_n70_3[0]),.din(w_dff_A_FzWSr4BD6_0),.clk(gclk));
	jdff dff_A_AHUzi0t56_0(.dout(w_dff_A_FzWSr4BD6_0),.din(w_dff_A_AHUzi0t56_0),.clk(gclk));
	jdff dff_A_OUgUnslh1_0(.dout(w_dff_A_AHUzi0t56_0),.din(w_dff_A_OUgUnslh1_0),.clk(gclk));
	jdff dff_A_SuvM4uh57_0(.dout(w_dff_A_OUgUnslh1_0),.din(w_dff_A_SuvM4uh57_0),.clk(gclk));
	jdff dff_A_3s6b7g909_1(.dout(w_G234_0[1]),.din(w_dff_A_3s6b7g909_1),.clk(gclk));
	jdff dff_A_tcZ97Uok8_2(.dout(w_G234_0[2]),.din(w_dff_A_tcZ97Uok8_2),.clk(gclk));
	jdff dff_A_KBzpCBu49_1(.dout(w_G221_0[1]),.din(w_dff_A_KBzpCBu49_1),.clk(gclk));
	jdff dff_A_U8XN4OYU1_1(.dout(w_dff_A_KBzpCBu49_1),.din(w_dff_A_U8XN4OYU1_1),.clk(gclk));
	jdff dff_A_GNKRvdAU7_1(.dout(w_n216_0[1]),.din(w_dff_A_GNKRvdAU7_1),.clk(gclk));
	jdff dff_B_P7nnRRTv2_1(.din(n215),.dout(w_dff_B_P7nnRRTv2_1),.clk(gclk));
	jdff dff_B_1bk6M5GQ3_1(.din(w_dff_B_P7nnRRTv2_1),.dout(w_dff_B_1bk6M5GQ3_1),.clk(gclk));
	jdff dff_B_4KWbCSTV9_1(.din(w_dff_B_1bk6M5GQ3_1),.dout(w_dff_B_4KWbCSTV9_1),.clk(gclk));
	jdff dff_A_Mu8pssWn9_0(.dout(w_n107_0[0]),.din(w_dff_A_Mu8pssWn9_0),.clk(gclk));
	jdff dff_A_Pb0nASbk4_0(.dout(w_dff_A_Mu8pssWn9_0),.din(w_dff_A_Pb0nASbk4_0),.clk(gclk));
	jdff dff_A_OqHcbhYV9_0(.dout(w_dff_A_Pb0nASbk4_0),.din(w_dff_A_OqHcbhYV9_0),.clk(gclk));
	jdff dff_A_5ziUDarr8_0(.dout(w_dff_A_OqHcbhYV9_0),.din(w_dff_A_5ziUDarr8_0),.clk(gclk));
	jdff dff_A_FlESALGf8_0(.dout(w_dff_A_5ziUDarr8_0),.din(w_dff_A_FlESALGf8_0),.clk(gclk));
	jdff dff_A_pBpvV1f40_0(.dout(w_dff_A_FlESALGf8_0),.din(w_dff_A_pBpvV1f40_0),.clk(gclk));
	jdff dff_A_DFFuUNat0_0(.dout(w_dff_A_pBpvV1f40_0),.din(w_dff_A_DFFuUNat0_0),.clk(gclk));
	jdff dff_A_gFvpE0dd0_0(.dout(w_dff_A_DFFuUNat0_0),.din(w_dff_A_gFvpE0dd0_0),.clk(gclk));
	jdff dff_A_vtIpbe572_0(.dout(w_dff_A_gFvpE0dd0_0),.din(w_dff_A_vtIpbe572_0),.clk(gclk));
	jdff dff_A_GUDFpytc8_0(.dout(w_dff_A_vtIpbe572_0),.din(w_dff_A_GUDFpytc8_0),.clk(gclk));
	jdff dff_A_b5PWxoNR4_0(.dout(w_dff_A_GUDFpytc8_0),.din(w_dff_A_b5PWxoNR4_0),.clk(gclk));
	jdff dff_A_L7Pb0JD02_0(.dout(w_dff_A_b5PWxoNR4_0),.din(w_dff_A_L7Pb0JD02_0),.clk(gclk));
	jdff dff_B_j7ORi5fJ4_1(.din(n104),.dout(w_dff_B_j7ORi5fJ4_1),.clk(gclk));
	jdff dff_A_4wDg9vF33_0(.dout(w_G125_0[0]),.din(w_dff_A_4wDg9vF33_0),.clk(gclk));
	jdff dff_A_MXWL5hor6_0(.dout(w_dff_A_4wDg9vF33_0),.din(w_dff_A_MXWL5hor6_0),.clk(gclk));
	jdff dff_A_aqyJSxiM3_0(.dout(w_dff_A_MXWL5hor6_0),.din(w_dff_A_aqyJSxiM3_0),.clk(gclk));
	jdff dff_A_jtM7ZKzT1_0(.dout(w_dff_A_aqyJSxiM3_0),.din(w_dff_A_jtM7ZKzT1_0),.clk(gclk));
	jdff dff_A_dsDAIxOa7_0(.dout(w_dff_A_jtM7ZKzT1_0),.din(w_dff_A_dsDAIxOa7_0),.clk(gclk));
	jdff dff_A_T2qMnk4w4_0(.dout(w_dff_A_dsDAIxOa7_0),.din(w_dff_A_T2qMnk4w4_0),.clk(gclk));
	jdff dff_A_TWFGBMQl6_0(.dout(w_dff_A_T2qMnk4w4_0),.din(w_dff_A_TWFGBMQl6_0),.clk(gclk));
	jdff dff_A_YZ9X46kS1_0(.dout(w_dff_A_TWFGBMQl6_0),.din(w_dff_A_YZ9X46kS1_0),.clk(gclk));
	jdff dff_A_66tUtsGc4_0(.dout(w_dff_A_YZ9X46kS1_0),.din(w_dff_A_66tUtsGc4_0),.clk(gclk));
	jdff dff_A_hdQf4NJJ2_0(.dout(w_dff_A_66tUtsGc4_0),.din(w_dff_A_hdQf4NJJ2_0),.clk(gclk));
	jdff dff_A_z1J1XDfe3_0(.dout(w_dff_A_hdQf4NJJ2_0),.din(w_dff_A_z1J1XDfe3_0),.clk(gclk));
	jdff dff_A_zgT0Dq8h2_0(.dout(w_dff_A_z1J1XDfe3_0),.din(w_dff_A_zgT0Dq8h2_0),.clk(gclk));
	jdff dff_A_4QPWBgRY3_1(.dout(w_G125_0[1]),.din(w_dff_A_4QPWBgRY3_1),.clk(gclk));
	jdff dff_A_CpdIIhVr7_1(.dout(w_dff_A_4QPWBgRY3_1),.din(w_dff_A_CpdIIhVr7_1),.clk(gclk));
	jdff dff_B_kmSRrjXT6_2(.din(G224),.dout(w_dff_B_kmSRrjXT6_2),.clk(gclk));
	jdff dff_A_hFLxOAdj0_0(.dout(w_n103_0[0]),.din(w_dff_A_hFLxOAdj0_0),.clk(gclk));
	jdff dff_A_If4Cfjzg8_0(.dout(w_dff_A_hFLxOAdj0_0),.din(w_dff_A_If4Cfjzg8_0),.clk(gclk));
	jdff dff_A_6bajqFHh2_0(.dout(w_dff_A_If4Cfjzg8_0),.din(w_dff_A_6bajqFHh2_0),.clk(gclk));
	jdff dff_A_hP0iS4SB2_0(.dout(w_dff_A_6bajqFHh2_0),.din(w_dff_A_hP0iS4SB2_0),.clk(gclk));
	jdff dff_A_xluGOmX67_0(.dout(w_dff_A_hP0iS4SB2_0),.din(w_dff_A_xluGOmX67_0),.clk(gclk));
	jdff dff_A_VysrE9j18_0(.dout(w_dff_A_xluGOmX67_0),.din(w_dff_A_VysrE9j18_0),.clk(gclk));
	jdff dff_A_UwJ20bYM5_0(.dout(w_dff_A_VysrE9j18_0),.din(w_dff_A_UwJ20bYM5_0),.clk(gclk));
	jdff dff_A_7xs0rADG6_0(.dout(w_dff_A_UwJ20bYM5_0),.din(w_dff_A_7xs0rADG6_0),.clk(gclk));
	jdff dff_A_gE4Z9ugN8_0(.dout(w_dff_A_7xs0rADG6_0),.din(w_dff_A_gE4Z9ugN8_0),.clk(gclk));
	jdff dff_A_7pHEecWW5_0(.dout(w_dff_A_gE4Z9ugN8_0),.din(w_dff_A_7pHEecWW5_0),.clk(gclk));
	jdff dff_A_ucgiOyXA1_0(.dout(w_dff_A_7pHEecWW5_0),.din(w_dff_A_ucgiOyXA1_0),.clk(gclk));
	jdff dff_A_lzRQ1gWq6_0(.dout(w_dff_A_ucgiOyXA1_0),.din(w_dff_A_lzRQ1gWq6_0),.clk(gclk));
	jdff dff_A_SKNglHc67_0(.dout(w_dff_A_lzRQ1gWq6_0),.din(w_dff_A_SKNglHc67_0),.clk(gclk));
	jdff dff_B_5vl8XvmS1_1(.din(n99),.dout(w_dff_B_5vl8XvmS1_1),.clk(gclk));
	jdff dff_A_giLq9S0A9_0(.dout(w_G107_0[0]),.din(w_dff_A_giLq9S0A9_0),.clk(gclk));
	jdff dff_A_93JdGNrh0_0(.dout(w_dff_A_giLq9S0A9_0),.din(w_dff_A_93JdGNrh0_0),.clk(gclk));
	jdff dff_A_MvBygeNP4_0(.dout(w_dff_A_93JdGNrh0_0),.din(w_dff_A_MvBygeNP4_0),.clk(gclk));
	jdff dff_A_mLDWJFyI4_0(.dout(w_dff_A_MvBygeNP4_0),.din(w_dff_A_mLDWJFyI4_0),.clk(gclk));
	jdff dff_A_VxnPZLMY8_0(.dout(w_dff_A_mLDWJFyI4_0),.din(w_dff_A_VxnPZLMY8_0),.clk(gclk));
	jdff dff_A_aivmkRLH2_0(.dout(w_dff_A_VxnPZLMY8_0),.din(w_dff_A_aivmkRLH2_0),.clk(gclk));
	jdff dff_A_rMuGxJE06_0(.dout(w_dff_A_aivmkRLH2_0),.din(w_dff_A_rMuGxJE06_0),.clk(gclk));
	jdff dff_A_drDFIaqG9_0(.dout(w_dff_A_rMuGxJE06_0),.din(w_dff_A_drDFIaqG9_0),.clk(gclk));
	jdff dff_A_ZYdwwfIB7_0(.dout(w_dff_A_drDFIaqG9_0),.din(w_dff_A_ZYdwwfIB7_0),.clk(gclk));
	jdff dff_A_61NtS2Qr3_0(.dout(w_dff_A_ZYdwwfIB7_0),.din(w_dff_A_61NtS2Qr3_0),.clk(gclk));
	jdff dff_A_B3U56SD00_0(.dout(w_dff_A_61NtS2Qr3_0),.din(w_dff_A_B3U56SD00_0),.clk(gclk));
	jdff dff_A_ZGo9KMbm9_0(.dout(w_dff_A_B3U56SD00_0),.din(w_dff_A_ZGo9KMbm9_0),.clk(gclk));
	jdff dff_A_PpbxIOMY5_0(.dout(w_G104_0[0]),.din(w_dff_A_PpbxIOMY5_0),.clk(gclk));
	jdff dff_A_giiRDZkl6_0(.dout(w_dff_A_PpbxIOMY5_0),.din(w_dff_A_giiRDZkl6_0),.clk(gclk));
	jdff dff_A_gFO4fKnu8_0(.dout(w_dff_A_giiRDZkl6_0),.din(w_dff_A_gFO4fKnu8_0),.clk(gclk));
	jdff dff_A_yUb77m495_0(.dout(w_dff_A_gFO4fKnu8_0),.din(w_dff_A_yUb77m495_0),.clk(gclk));
	jdff dff_A_NoBqEcxZ5_0(.dout(w_dff_A_yUb77m495_0),.din(w_dff_A_NoBqEcxZ5_0),.clk(gclk));
	jdff dff_A_DKw5nSvP6_0(.dout(w_dff_A_NoBqEcxZ5_0),.din(w_dff_A_DKw5nSvP6_0),.clk(gclk));
	jdff dff_A_ALrm9nvP8_0(.dout(w_dff_A_DKw5nSvP6_0),.din(w_dff_A_ALrm9nvP8_0),.clk(gclk));
	jdff dff_A_aTsbvFUy1_0(.dout(w_dff_A_ALrm9nvP8_0),.din(w_dff_A_aTsbvFUy1_0),.clk(gclk));
	jdff dff_A_7bcKgO1E1_0(.dout(w_dff_A_aTsbvFUy1_0),.din(w_dff_A_7bcKgO1E1_0),.clk(gclk));
	jdff dff_A_2HBKoYRK1_0(.dout(w_dff_A_7bcKgO1E1_0),.din(w_dff_A_2HBKoYRK1_0),.clk(gclk));
	jdff dff_A_dzbJfQrZ0_0(.dout(w_dff_A_2HBKoYRK1_0),.din(w_dff_A_dzbJfQrZ0_0),.clk(gclk));
	jdff dff_A_VA4WSqGf3_0(.dout(w_dff_A_dzbJfQrZ0_0),.din(w_dff_A_VA4WSqGf3_0),.clk(gclk));
	jdff dff_A_etYR0HCN8_1(.dout(w_G104_0[1]),.din(w_dff_A_etYR0HCN8_1),.clk(gclk));
	jdff dff_A_vdRpM4MQ1_1(.dout(w_dff_A_etYR0HCN8_1),.din(w_dff_A_vdRpM4MQ1_1),.clk(gclk));
	jdff dff_A_FhOJenYV3_1(.dout(w_G122_1[1]),.din(w_dff_A_FhOJenYV3_1),.clk(gclk));
	jdff dff_A_ydhDSGlf7_1(.dout(w_G122_0[1]),.din(w_dff_A_ydhDSGlf7_1),.clk(gclk));
	jdff dff_A_sM50eAFw6_1(.dout(w_dff_A_ydhDSGlf7_1),.din(w_dff_A_sM50eAFw6_1),.clk(gclk));
	jdff dff_A_ioKRfuF49_1(.dout(w_dff_A_sM50eAFw6_1),.din(w_dff_A_ioKRfuF49_1),.clk(gclk));
	jdff dff_A_VJEoO8Ns9_1(.dout(w_dff_A_ioKRfuF49_1),.din(w_dff_A_VJEoO8Ns9_1),.clk(gclk));
	jdff dff_A_zhEfnZEw1_1(.dout(w_dff_A_VJEoO8Ns9_1),.din(w_dff_A_zhEfnZEw1_1),.clk(gclk));
	jdff dff_A_JEDRLKxa8_1(.dout(w_dff_A_zhEfnZEw1_1),.din(w_dff_A_JEDRLKxa8_1),.clk(gclk));
	jdff dff_A_AANOPBGj2_1(.dout(w_dff_A_JEDRLKxa8_1),.din(w_dff_A_AANOPBGj2_1),.clk(gclk));
	jdff dff_A_UgnibWgb1_1(.dout(w_dff_A_AANOPBGj2_1),.din(w_dff_A_UgnibWgb1_1),.clk(gclk));
	jdff dff_A_IlKCEZte2_1(.dout(w_dff_A_UgnibWgb1_1),.din(w_dff_A_IlKCEZte2_1),.clk(gclk));
	jdff dff_A_wPeWIeJE3_1(.dout(w_dff_A_IlKCEZte2_1),.din(w_dff_A_wPeWIeJE3_1),.clk(gclk));
	jdff dff_A_XM7YifRl2_1(.dout(w_dff_A_wPeWIeJE3_1),.din(w_dff_A_XM7YifRl2_1),.clk(gclk));
	jdff dff_A_A11H96eB5_1(.dout(w_dff_A_XM7YifRl2_1),.din(w_dff_A_A11H96eB5_1),.clk(gclk));
	jdff dff_A_CA6hxhaa2_2(.dout(w_G122_0[2]),.din(w_dff_A_CA6hxhaa2_2),.clk(gclk));
	jdff dff_A_P1Y0U8u88_1(.dout(w_G110_1[1]),.din(w_dff_A_P1Y0U8u88_1),.clk(gclk));
	jdff dff_A_kSXrRche8_1(.dout(w_dff_A_P1Y0U8u88_1),.din(w_dff_A_kSXrRche8_1),.clk(gclk));
	jdff dff_A_kkskv2WD1_1(.dout(w_dff_A_kSXrRche8_1),.din(w_dff_A_kkskv2WD1_1),.clk(gclk));
	jdff dff_A_17WFrIPe7_1(.dout(w_dff_A_kkskv2WD1_1),.din(w_dff_A_17WFrIPe7_1),.clk(gclk));
	jdff dff_A_BlxwlLW53_1(.dout(w_dff_A_17WFrIPe7_1),.din(w_dff_A_BlxwlLW53_1),.clk(gclk));
	jdff dff_A_2YhUJvZh6_1(.dout(w_G110_0[1]),.din(w_dff_A_2YhUJvZh6_1),.clk(gclk));
	jdff dff_A_IJnM518G8_1(.dout(w_dff_A_2YhUJvZh6_1),.din(w_dff_A_IJnM518G8_1),.clk(gclk));
	jdff dff_A_cT8yGlSW7_1(.dout(w_dff_A_IJnM518G8_1),.din(w_dff_A_cT8yGlSW7_1),.clk(gclk));
	jdff dff_A_7MjEoGRb8_1(.dout(w_dff_A_cT8yGlSW7_1),.din(w_dff_A_7MjEoGRb8_1),.clk(gclk));
	jdff dff_A_Q12is24H8_1(.dout(w_dff_A_7MjEoGRb8_1),.din(w_dff_A_Q12is24H8_1),.clk(gclk));
	jdff dff_A_tnAZyTG27_1(.dout(w_dff_A_Q12is24H8_1),.din(w_dff_A_tnAZyTG27_1),.clk(gclk));
	jdff dff_A_3Ttm5HXl0_1(.dout(w_dff_A_tnAZyTG27_1),.din(w_dff_A_3Ttm5HXl0_1),.clk(gclk));
	jdff dff_A_3mxvC7sV4_1(.dout(w_dff_A_3Ttm5HXl0_1),.din(w_dff_A_3mxvC7sV4_1),.clk(gclk));
	jdff dff_A_Ox3Ox4Mj2_1(.dout(w_dff_A_3mxvC7sV4_1),.din(w_dff_A_Ox3Ox4Mj2_1),.clk(gclk));
	jdff dff_A_tvozGGvU1_1(.dout(w_dff_A_Ox3Ox4Mj2_1),.din(w_dff_A_tvozGGvU1_1),.clk(gclk));
	jdff dff_A_KWzCnMVZ9_1(.dout(w_dff_A_tvozGGvU1_1),.din(w_dff_A_KWzCnMVZ9_1),.clk(gclk));
	jdff dff_A_3jrU2D8Q1_1(.dout(w_dff_A_KWzCnMVZ9_1),.din(w_dff_A_3jrU2D8Q1_1),.clk(gclk));
	jdff dff_A_EtFij2pM5_1(.dout(w_n70_0[1]),.din(w_dff_A_EtFij2pM5_1),.clk(gclk));
	jdff dff_A_TqjaJjqP6_1(.dout(w_dff_A_EtFij2pM5_1),.din(w_dff_A_TqjaJjqP6_1),.clk(gclk));
	jdff dff_A_GdEnrtP53_1(.dout(w_dff_A_TqjaJjqP6_1),.din(w_dff_A_GdEnrtP53_1),.clk(gclk));
	jdff dff_A_1EvKxreK4_1(.dout(w_dff_A_GdEnrtP53_1),.din(w_dff_A_1EvKxreK4_1),.clk(gclk));
	jdff dff_A_sDiT8r3D9_1(.dout(w_n97_0[1]),.din(w_dff_A_sDiT8r3D9_1),.clk(gclk));
	jdff dff_A_BiC8QFpX8_1(.dout(w_dff_A_sDiT8r3D9_1),.din(w_dff_A_BiC8QFpX8_1),.clk(gclk));
	jdff dff_A_qLKm3xvd3_1(.dout(w_dff_A_BiC8QFpX8_1),.din(w_dff_A_qLKm3xvd3_1),.clk(gclk));
	jdff dff_A_xyPaCXtD7_1(.dout(w_dff_A_qLKm3xvd3_1),.din(w_dff_A_xyPaCXtD7_1),.clk(gclk));
	jdff dff_A_Q9VlMNWd9_0(.dout(w_n95_0[0]),.din(w_dff_A_Q9VlMNWd9_0),.clk(gclk));
	jdff dff_A_0U42nwJQ0_0(.dout(w_dff_A_Q9VlMNWd9_0),.din(w_dff_A_0U42nwJQ0_0),.clk(gclk));
	jdff dff_A_z9OCVGFs0_0(.dout(w_dff_A_0U42nwJQ0_0),.din(w_dff_A_z9OCVGFs0_0),.clk(gclk));
	jdff dff_A_3SNReyuh6_0(.dout(w_dff_A_z9OCVGFs0_0),.din(w_dff_A_3SNReyuh6_0),.clk(gclk));
	jdff dff_A_CgzDlYLy2_0(.dout(w_dff_A_3SNReyuh6_0),.din(w_dff_A_CgzDlYLy2_0),.clk(gclk));
	jdff dff_A_eccbc3R32_1(.dout(w_n95_0[1]),.din(w_dff_A_eccbc3R32_1),.clk(gclk));
	jdff dff_A_XwczMQQv7_1(.dout(w_dff_A_eccbc3R32_1),.din(w_dff_A_XwczMQQv7_1),.clk(gclk));
	jdff dff_A_25eBm0iU6_1(.dout(w_dff_A_XwczMQQv7_1),.din(w_dff_A_25eBm0iU6_1),.clk(gclk));
	jdff dff_A_GJx2WTsJ3_1(.dout(w_dff_A_25eBm0iU6_1),.din(w_dff_A_GJx2WTsJ3_1),.clk(gclk));
	jdff dff_A_F3e9q6nE5_1(.dout(w_dff_A_GJx2WTsJ3_1),.din(w_dff_A_F3e9q6nE5_1),.clk(gclk));
	jdff dff_A_ljeLwGY25_2(.dout(w_G902_3[2]),.din(w_dff_A_ljeLwGY25_2),.clk(gclk));
	jdff dff_A_3HH2s7SH2_2(.dout(w_dff_A_ljeLwGY25_2),.din(w_dff_A_3HH2s7SH2_2),.clk(gclk));
	jdff dff_A_YyFqHaP03_2(.dout(w_dff_A_3HH2s7SH2_2),.din(w_dff_A_YyFqHaP03_2),.clk(gclk));
	jdff dff_A_lBjvXLsJ8_2(.dout(w_dff_A_YyFqHaP03_2),.din(w_dff_A_lBjvXLsJ8_2),.clk(gclk));
	jdff dff_A_MXJGJvzN2_2(.dout(w_dff_A_lBjvXLsJ8_2),.din(w_dff_A_MXJGJvzN2_2),.clk(gclk));
	jdff dff_A_EzFCGtMC6_2(.dout(w_dff_A_MXJGJvzN2_2),.din(w_dff_A_EzFCGtMC6_2),.clk(gclk));
	jdff dff_A_1ct4tUVW5_2(.dout(w_dff_A_EzFCGtMC6_2),.din(w_dff_A_1ct4tUVW5_2),.clk(gclk));
	jdff dff_A_tDjuBF022_1(.dout(w_G214_0[1]),.din(w_dff_A_tDjuBF022_1),.clk(gclk));
	jdff dff_A_TFlHmIqk2_0(.dout(w_n90_0[0]),.din(w_dff_A_TFlHmIqk2_0),.clk(gclk));
	jdff dff_A_VoHE9fBq5_0(.dout(w_dff_A_TFlHmIqk2_0),.din(w_dff_A_VoHE9fBq5_0),.clk(gclk));
	jdff dff_A_e2jJr84u4_0(.dout(w_dff_A_VoHE9fBq5_0),.din(w_dff_A_e2jJr84u4_0),.clk(gclk));
	jdff dff_A_vlfJkYt84_0(.dout(w_dff_A_e2jJr84u4_0),.din(w_dff_A_vlfJkYt84_0),.clk(gclk));
	jdff dff_A_psgFL68B2_0(.dout(w_dff_A_vlfJkYt84_0),.din(w_dff_A_psgFL68B2_0),.clk(gclk));
	jdff dff_A_Y50veSqC4_0(.dout(w_dff_A_psgFL68B2_0),.din(w_dff_A_Y50veSqC4_0),.clk(gclk));
	jdff dff_A_khJMROJi4_0(.dout(w_dff_A_Y50veSqC4_0),.din(w_dff_A_khJMROJi4_0),.clk(gclk));
	jdff dff_A_7TayJBC28_0(.dout(w_dff_A_khJMROJi4_0),.din(w_dff_A_7TayJBC28_0),.clk(gclk));
	jdff dff_A_PgsX1UY79_0(.dout(w_dff_A_7TayJBC28_0),.din(w_dff_A_PgsX1UY79_0),.clk(gclk));
	jdff dff_A_xwdIUY8b6_0(.dout(w_dff_A_PgsX1UY79_0),.din(w_dff_A_xwdIUY8b6_0),.clk(gclk));
	jdff dff_A_wVPmatmG8_0(.dout(w_dff_A_xwdIUY8b6_0),.din(w_dff_A_wVPmatmG8_0),.clk(gclk));
	jdff dff_A_ARU548hm1_0(.dout(w_dff_A_wVPmatmG8_0),.din(w_dff_A_ARU548hm1_0),.clk(gclk));
	jdff dff_A_lu4iJZYK4_0(.dout(w_G953_1[0]),.din(w_dff_A_lu4iJZYK4_0),.clk(gclk));
	jdff dff_A_C9fp8HEz8_0(.dout(w_dff_A_lu4iJZYK4_0),.din(w_dff_A_C9fp8HEz8_0),.clk(gclk));
	jdff dff_A_YPuRu8le4_0(.dout(w_dff_A_C9fp8HEz8_0),.din(w_dff_A_YPuRu8le4_0),.clk(gclk));
	jdff dff_A_bB8PgO1H0_0(.dout(w_dff_A_YPuRu8le4_0),.din(w_dff_A_bB8PgO1H0_0),.clk(gclk));
	jdff dff_A_6VQt6JLB0_0(.dout(w_dff_A_bB8PgO1H0_0),.din(w_dff_A_6VQt6JLB0_0),.clk(gclk));
	jdff dff_A_Ar2fbf4V7_0(.dout(w_dff_A_6VQt6JLB0_0),.din(w_dff_A_Ar2fbf4V7_0),.clk(gclk));
	jdff dff_A_x0V1XLR20_0(.dout(w_dff_A_Ar2fbf4V7_0),.din(w_dff_A_x0V1XLR20_0),.clk(gclk));
	jdff dff_A_vGm6oouJ3_0(.dout(w_dff_A_x0V1XLR20_0),.din(w_dff_A_vGm6oouJ3_0),.clk(gclk));
	jdff dff_A_zBiBCKun6_0(.dout(w_dff_A_vGm6oouJ3_0),.din(w_dff_A_zBiBCKun6_0),.clk(gclk));
	jdff dff_A_pF8VoppL0_0(.dout(w_dff_A_zBiBCKun6_0),.din(w_dff_A_pF8VoppL0_0),.clk(gclk));
	jdff dff_A_AO545wsb5_0(.dout(w_dff_A_pF8VoppL0_0),.din(w_dff_A_AO545wsb5_0),.clk(gclk));
	jdff dff_A_ReU8cIDJ8_0(.dout(w_dff_A_AO545wsb5_0),.din(w_dff_A_ReU8cIDJ8_0),.clk(gclk));
	jdff dff_A_Tesifn7c3_1(.dout(w_G953_0[1]),.din(w_dff_A_Tesifn7c3_1),.clk(gclk));
	jdff dff_A_r5dHI0Mg5_1(.dout(w_dff_A_Tesifn7c3_1),.din(w_dff_A_r5dHI0Mg5_1),.clk(gclk));
	jdff dff_A_JaSSlB4U1_1(.dout(w_dff_A_r5dHI0Mg5_1),.din(w_dff_A_JaSSlB4U1_1),.clk(gclk));
	jdff dff_A_01mEqRT91_1(.dout(w_dff_A_JaSSlB4U1_1),.din(w_dff_A_01mEqRT91_1),.clk(gclk));
	jdff dff_A_ep9tyags2_1(.dout(w_dff_A_01mEqRT91_1),.din(w_dff_A_ep9tyags2_1),.clk(gclk));
	jdff dff_A_c1QAZGLK1_1(.dout(w_dff_A_ep9tyags2_1),.din(w_dff_A_c1QAZGLK1_1),.clk(gclk));
	jdff dff_A_OsTznZ9H0_1(.dout(w_dff_A_c1QAZGLK1_1),.din(w_dff_A_OsTznZ9H0_1),.clk(gclk));
	jdff dff_A_GxhoUOcO6_1(.dout(w_dff_A_OsTznZ9H0_1),.din(w_dff_A_GxhoUOcO6_1),.clk(gclk));
	jdff dff_A_g1tDK9Uz9_1(.dout(w_dff_A_GxhoUOcO6_1),.din(w_dff_A_g1tDK9Uz9_1),.clk(gclk));
	jdff dff_A_Lrt6JbTI1_1(.dout(w_dff_A_g1tDK9Uz9_1),.din(w_dff_A_Lrt6JbTI1_1),.clk(gclk));
	jdff dff_A_oXWUJnBQ8_1(.dout(w_dff_A_Lrt6JbTI1_1),.din(w_dff_A_oXWUJnBQ8_1),.clk(gclk));
	jdff dff_A_LvjoHDe40_1(.dout(w_dff_A_oXWUJnBQ8_1),.din(w_dff_A_LvjoHDe40_1),.clk(gclk));
	jdff dff_A_rP6NhMxu7_1(.dout(w_dff_A_LvjoHDe40_1),.din(w_dff_A_rP6NhMxu7_1),.clk(gclk));
	jdff dff_A_nISm5J6t7_1(.dout(w_dff_A_rP6NhMxu7_1),.din(w_dff_A_nISm5J6t7_1),.clk(gclk));
	jdff dff_A_4NxQWxMU5_1(.dout(w_dff_A_nISm5J6t7_1),.din(w_dff_A_4NxQWxMU5_1),.clk(gclk));
	jdff dff_A_7YHlHYqo4_2(.dout(w_G953_0[2]),.din(w_dff_A_7YHlHYqo4_2),.clk(gclk));
	jdff dff_A_c5zEmjNo8_2(.dout(w_dff_A_7YHlHYqo4_2),.din(w_dff_A_c5zEmjNo8_2),.clk(gclk));
	jdff dff_A_hxMpqtlg4_2(.dout(w_dff_A_c5zEmjNo8_2),.din(w_dff_A_hxMpqtlg4_2),.clk(gclk));
	jdff dff_A_E0DfOccd9_2(.dout(w_dff_A_hxMpqtlg4_2),.din(w_dff_A_E0DfOccd9_2),.clk(gclk));
	jdff dff_A_BNiJlq0L4_2(.dout(w_dff_A_E0DfOccd9_2),.din(w_dff_A_BNiJlq0L4_2),.clk(gclk));
	jdff dff_A_IOydEwTp7_2(.dout(w_dff_A_BNiJlq0L4_2),.din(w_dff_A_IOydEwTp7_2),.clk(gclk));
	jdff dff_A_4wOHPwQ55_2(.dout(w_dff_A_IOydEwTp7_2),.din(w_dff_A_4wOHPwQ55_2),.clk(gclk));
	jdff dff_A_V9BDueEv6_2(.dout(w_dff_A_4wOHPwQ55_2),.din(w_dff_A_V9BDueEv6_2),.clk(gclk));
	jdff dff_A_4E1MKIdp5_2(.dout(w_dff_A_V9BDueEv6_2),.din(w_dff_A_4E1MKIdp5_2),.clk(gclk));
	jdff dff_A_p6r6U7192_2(.dout(w_dff_A_4E1MKIdp5_2),.din(w_dff_A_p6r6U7192_2),.clk(gclk));
	jdff dff_A_YT0iPKEZ2_2(.dout(w_dff_A_p6r6U7192_2),.din(w_dff_A_YT0iPKEZ2_2),.clk(gclk));
	jdff dff_A_uE5DdWu64_2(.dout(w_dff_A_YT0iPKEZ2_2),.din(w_dff_A_uE5DdWu64_2),.clk(gclk));
	jdff dff_A_lR96zMAH0_2(.dout(w_dff_A_uE5DdWu64_2),.din(w_dff_A_lR96zMAH0_2),.clk(gclk));
	jdff dff_A_2C4bJCot3_2(.dout(w_dff_A_lR96zMAH0_2),.din(w_dff_A_2C4bJCot3_2),.clk(gclk));
	jdff dff_A_aMzM9twT2_2(.dout(w_dff_A_2C4bJCot3_2),.din(w_dff_A_aMzM9twT2_2),.clk(gclk));
	jdff dff_A_hgRE24Ur4_1(.dout(w_G210_0[1]),.din(w_dff_A_hgRE24Ur4_1),.clk(gclk));
	jdff dff_A_zDn1sl8B6_0(.dout(w_G101_0[0]),.din(w_dff_A_zDn1sl8B6_0),.clk(gclk));
	jdff dff_A_Pl2UOARS7_0(.dout(w_dff_A_zDn1sl8B6_0),.din(w_dff_A_Pl2UOARS7_0),.clk(gclk));
	jdff dff_A_UcdiNOaL2_0(.dout(w_dff_A_Pl2UOARS7_0),.din(w_dff_A_UcdiNOaL2_0),.clk(gclk));
	jdff dff_A_L49YtfNm5_0(.dout(w_dff_A_UcdiNOaL2_0),.din(w_dff_A_L49YtfNm5_0),.clk(gclk));
	jdff dff_A_YAKN5FWX1_0(.dout(w_dff_A_L49YtfNm5_0),.din(w_dff_A_YAKN5FWX1_0),.clk(gclk));
	jdff dff_A_AIRXoOpO8_0(.dout(w_dff_A_YAKN5FWX1_0),.din(w_dff_A_AIRXoOpO8_0),.clk(gclk));
	jdff dff_A_BidEmMFn2_0(.dout(w_dff_A_AIRXoOpO8_0),.din(w_dff_A_BidEmMFn2_0),.clk(gclk));
	jdff dff_A_NnIqgKkW5_0(.dout(w_dff_A_BidEmMFn2_0),.din(w_dff_A_NnIqgKkW5_0),.clk(gclk));
	jdff dff_A_d0cJmlpv2_0(.dout(w_dff_A_NnIqgKkW5_0),.din(w_dff_A_d0cJmlpv2_0),.clk(gclk));
	jdff dff_A_AhXpHyez9_0(.dout(w_dff_A_d0cJmlpv2_0),.din(w_dff_A_AhXpHyez9_0),.clk(gclk));
	jdff dff_A_t1gICSgz1_0(.dout(w_dff_A_AhXpHyez9_0),.din(w_dff_A_t1gICSgz1_0),.clk(gclk));
	jdff dff_A_MzGgJx775_2(.dout(w_G101_0[2]),.din(w_dff_A_MzGgJx775_2),.clk(gclk));
	jdff dff_B_CNYfRje88_3(.din(G101),.dout(w_dff_B_CNYfRje88_3),.clk(gclk));
	jdff dff_A_dTNbfKqW2_1(.dout(w_n84_0[1]),.din(w_dff_A_dTNbfKqW2_1),.clk(gclk));
	jdff dff_A_gySoFXbb7_0(.dout(w_G119_0[0]),.din(w_dff_A_gySoFXbb7_0),.clk(gclk));
	jdff dff_A_IzVn4X9S1_0(.dout(w_dff_A_gySoFXbb7_0),.din(w_dff_A_IzVn4X9S1_0),.clk(gclk));
	jdff dff_A_a52UWG9N9_0(.dout(w_dff_A_IzVn4X9S1_0),.din(w_dff_A_a52UWG9N9_0),.clk(gclk));
	jdff dff_A_ciRUgfln5_0(.dout(w_dff_A_a52UWG9N9_0),.din(w_dff_A_ciRUgfln5_0),.clk(gclk));
	jdff dff_A_0DQUmZFa0_0(.dout(w_dff_A_ciRUgfln5_0),.din(w_dff_A_0DQUmZFa0_0),.clk(gclk));
	jdff dff_A_aL6OIHWs4_0(.dout(w_dff_A_0DQUmZFa0_0),.din(w_dff_A_aL6OIHWs4_0),.clk(gclk));
	jdff dff_A_cM89K7PN7_0(.dout(w_dff_A_aL6OIHWs4_0),.din(w_dff_A_cM89K7PN7_0),.clk(gclk));
	jdff dff_A_bOgEq25R1_0(.dout(w_dff_A_cM89K7PN7_0),.din(w_dff_A_bOgEq25R1_0),.clk(gclk));
	jdff dff_A_QpA6hHJu8_0(.dout(w_dff_A_bOgEq25R1_0),.din(w_dff_A_QpA6hHJu8_0),.clk(gclk));
	jdff dff_A_IyxPokaL6_0(.dout(w_dff_A_QpA6hHJu8_0),.din(w_dff_A_IyxPokaL6_0),.clk(gclk));
	jdff dff_A_FWNJJz255_0(.dout(w_dff_A_IyxPokaL6_0),.din(w_dff_A_FWNJJz255_0),.clk(gclk));
	jdff dff_A_JRMPtdzP8_0(.dout(w_dff_A_FWNJJz255_0),.din(w_dff_A_JRMPtdzP8_0),.clk(gclk));
	jdff dff_A_Jwv0xFl69_0(.dout(w_G116_0[0]),.din(w_dff_A_Jwv0xFl69_0),.clk(gclk));
	jdff dff_A_Jrv4KkjY5_0(.dout(w_dff_A_Jwv0xFl69_0),.din(w_dff_A_Jrv4KkjY5_0),.clk(gclk));
	jdff dff_A_hbsWC19E6_0(.dout(w_dff_A_Jrv4KkjY5_0),.din(w_dff_A_hbsWC19E6_0),.clk(gclk));
	jdff dff_A_nxKKuqmQ3_0(.dout(w_dff_A_hbsWC19E6_0),.din(w_dff_A_nxKKuqmQ3_0),.clk(gclk));
	jdff dff_A_5VAfND6l6_0(.dout(w_dff_A_nxKKuqmQ3_0),.din(w_dff_A_5VAfND6l6_0),.clk(gclk));
	jdff dff_A_PLCzIBgv4_0(.dout(w_dff_A_5VAfND6l6_0),.din(w_dff_A_PLCzIBgv4_0),.clk(gclk));
	jdff dff_A_HnUe3F6y4_0(.dout(w_dff_A_PLCzIBgv4_0),.din(w_dff_A_HnUe3F6y4_0),.clk(gclk));
	jdff dff_A_nV6Otq3z1_0(.dout(w_dff_A_HnUe3F6y4_0),.din(w_dff_A_nV6Otq3z1_0),.clk(gclk));
	jdff dff_A_NqwXV67n3_0(.dout(w_dff_A_nV6Otq3z1_0),.din(w_dff_A_NqwXV67n3_0),.clk(gclk));
	jdff dff_A_3wy2t2RS7_0(.dout(w_dff_A_NqwXV67n3_0),.din(w_dff_A_3wy2t2RS7_0),.clk(gclk));
	jdff dff_A_vhvZQKxB3_0(.dout(w_dff_A_3wy2t2RS7_0),.din(w_dff_A_vhvZQKxB3_0),.clk(gclk));
	jdff dff_A_Q0lthbmY7_0(.dout(w_dff_A_vhvZQKxB3_0),.din(w_dff_A_Q0lthbmY7_0),.clk(gclk));
	jdff dff_A_W3bMojaO0_0(.dout(w_G113_0[0]),.din(w_dff_A_W3bMojaO0_0),.clk(gclk));
	jdff dff_A_xdonyWUW5_0(.dout(w_dff_A_W3bMojaO0_0),.din(w_dff_A_xdonyWUW5_0),.clk(gclk));
	jdff dff_A_5QXqa2PP2_0(.dout(w_dff_A_xdonyWUW5_0),.din(w_dff_A_5QXqa2PP2_0),.clk(gclk));
	jdff dff_A_pLD4ERRR2_0(.dout(w_dff_A_5QXqa2PP2_0),.din(w_dff_A_pLD4ERRR2_0),.clk(gclk));
	jdff dff_A_g0l0pkBX9_0(.dout(w_dff_A_pLD4ERRR2_0),.din(w_dff_A_g0l0pkBX9_0),.clk(gclk));
	jdff dff_A_qpxDMKE01_0(.dout(w_dff_A_g0l0pkBX9_0),.din(w_dff_A_qpxDMKE01_0),.clk(gclk));
	jdff dff_A_eYjeBoBV6_0(.dout(w_dff_A_qpxDMKE01_0),.din(w_dff_A_eYjeBoBV6_0),.clk(gclk));
	jdff dff_A_I9y0xZiD0_0(.dout(w_dff_A_eYjeBoBV6_0),.din(w_dff_A_I9y0xZiD0_0),.clk(gclk));
	jdff dff_A_o0A0cI0X7_0(.dout(w_dff_A_I9y0xZiD0_0),.din(w_dff_A_o0A0cI0X7_0),.clk(gclk));
	jdff dff_A_xP5ed0Si7_0(.dout(w_dff_A_o0A0cI0X7_0),.din(w_dff_A_xP5ed0Si7_0),.clk(gclk));
	jdff dff_A_kpEjZ3k20_0(.dout(w_dff_A_xP5ed0Si7_0),.din(w_dff_A_kpEjZ3k20_0),.clk(gclk));
	jdff dff_A_qClEJX0E5_0(.dout(w_dff_A_kpEjZ3k20_0),.din(w_dff_A_qClEJX0E5_0),.clk(gclk));
	jdff dff_B_0QcSUpE87_1(.din(n76),.dout(w_dff_B_0QcSUpE87_1),.clk(gclk));
	jdff dff_A_OxbtqQiH3_0(.dout(w_G146_0[0]),.din(w_dff_A_OxbtqQiH3_0),.clk(gclk));
	jdff dff_A_i5KrNt6T9_0(.dout(w_dff_A_OxbtqQiH3_0),.din(w_dff_A_i5KrNt6T9_0),.clk(gclk));
	jdff dff_A_yd3QNXME2_0(.dout(w_dff_A_i5KrNt6T9_0),.din(w_dff_A_yd3QNXME2_0),.clk(gclk));
	jdff dff_A_acZ5Ytfb4_0(.dout(w_dff_A_yd3QNXME2_0),.din(w_dff_A_acZ5Ytfb4_0),.clk(gclk));
	jdff dff_A_cfTIUGSJ8_0(.dout(w_dff_A_acZ5Ytfb4_0),.din(w_dff_A_cfTIUGSJ8_0),.clk(gclk));
	jdff dff_A_JQrdEivi1_0(.dout(w_dff_A_cfTIUGSJ8_0),.din(w_dff_A_JQrdEivi1_0),.clk(gclk));
	jdff dff_A_QfZHXklO8_0(.dout(w_dff_A_JQrdEivi1_0),.din(w_dff_A_QfZHXklO8_0),.clk(gclk));
	jdff dff_A_o8Hxctjp1_0(.dout(w_dff_A_QfZHXklO8_0),.din(w_dff_A_o8Hxctjp1_0),.clk(gclk));
	jdff dff_A_NH9undmQ0_0(.dout(w_dff_A_o8Hxctjp1_0),.din(w_dff_A_NH9undmQ0_0),.clk(gclk));
	jdff dff_A_CNXFDjFT6_0(.dout(w_dff_A_NH9undmQ0_0),.din(w_dff_A_CNXFDjFT6_0),.clk(gclk));
	jdff dff_A_UuCND0Wo4_0(.dout(w_dff_A_CNXFDjFT6_0),.din(w_dff_A_UuCND0Wo4_0),.clk(gclk));
	jdff dff_A_g4VM4Dvy0_0(.dout(w_dff_A_UuCND0Wo4_0),.din(w_dff_A_g4VM4Dvy0_0),.clk(gclk));
	jdff dff_A_3DLO0SEv4_1(.dout(w_G143_0[1]),.din(w_dff_A_3DLO0SEv4_1),.clk(gclk));
	jdff dff_A_KO2VCb6W2_1(.dout(w_dff_A_3DLO0SEv4_1),.din(w_dff_A_KO2VCb6W2_1),.clk(gclk));
	jdff dff_A_lUd35UYF5_1(.dout(w_dff_A_KO2VCb6W2_1),.din(w_dff_A_lUd35UYF5_1),.clk(gclk));
	jdff dff_A_2ge8XyT67_1(.dout(w_dff_A_lUd35UYF5_1),.din(w_dff_A_2ge8XyT67_1),.clk(gclk));
	jdff dff_A_ZasxbszV9_1(.dout(w_dff_A_2ge8XyT67_1),.din(w_dff_A_ZasxbszV9_1),.clk(gclk));
	jdff dff_A_YL5btN9k8_1(.dout(w_dff_A_ZasxbszV9_1),.din(w_dff_A_YL5btN9k8_1),.clk(gclk));
	jdff dff_A_ausLFpKq4_1(.dout(w_dff_A_YL5btN9k8_1),.din(w_dff_A_ausLFpKq4_1),.clk(gclk));
	jdff dff_A_5KnuFEmd1_1(.dout(w_dff_A_ausLFpKq4_1),.din(w_dff_A_5KnuFEmd1_1),.clk(gclk));
	jdff dff_A_xC3uKHfr6_1(.dout(w_dff_A_5KnuFEmd1_1),.din(w_dff_A_xC3uKHfr6_1),.clk(gclk));
	jdff dff_A_AKH3bdFV4_1(.dout(w_dff_A_xC3uKHfr6_1),.din(w_dff_A_AKH3bdFV4_1),.clk(gclk));
	jdff dff_A_sRTDwoK12_1(.dout(w_dff_A_AKH3bdFV4_1),.din(w_dff_A_sRTDwoK12_1),.clk(gclk));
	jdff dff_A_ztNSLy4P5_1(.dout(w_dff_A_sRTDwoK12_1),.din(w_dff_A_ztNSLy4P5_1),.clk(gclk));
	jdff dff_A_8uYIgGTS0_2(.dout(w_G143_0[2]),.din(w_dff_A_8uYIgGTS0_2),.clk(gclk));
	jdff dff_A_UCIhReKV0_0(.dout(w_G128_1[0]),.din(w_dff_A_UCIhReKV0_0),.clk(gclk));
	jdff dff_A_pfVDzSTE0_1(.dout(w_G128_0[1]),.din(w_dff_A_pfVDzSTE0_1),.clk(gclk));
	jdff dff_A_KgRkFrKY7_1(.dout(w_dff_A_pfVDzSTE0_1),.din(w_dff_A_KgRkFrKY7_1),.clk(gclk));
	jdff dff_A_kACUpb8O4_1(.dout(w_dff_A_KgRkFrKY7_1),.din(w_dff_A_kACUpb8O4_1),.clk(gclk));
	jdff dff_A_AlS9pvZO9_1(.dout(w_dff_A_kACUpb8O4_1),.din(w_dff_A_AlS9pvZO9_1),.clk(gclk));
	jdff dff_A_o6MO40ph5_1(.dout(w_dff_A_AlS9pvZO9_1),.din(w_dff_A_o6MO40ph5_1),.clk(gclk));
	jdff dff_A_J2Q4ckKZ9_1(.dout(w_dff_A_o6MO40ph5_1),.din(w_dff_A_J2Q4ckKZ9_1),.clk(gclk));
	jdff dff_A_UP4Oqxzk7_1(.dout(w_dff_A_J2Q4ckKZ9_1),.din(w_dff_A_UP4Oqxzk7_1),.clk(gclk));
	jdff dff_A_MjJSgreQ2_1(.dout(w_dff_A_UP4Oqxzk7_1),.din(w_dff_A_MjJSgreQ2_1),.clk(gclk));
	jdff dff_A_6UXBdWxc1_1(.dout(w_dff_A_MjJSgreQ2_1),.din(w_dff_A_6UXBdWxc1_1),.clk(gclk));
	jdff dff_A_zLLi7gXj2_1(.dout(w_dff_A_6UXBdWxc1_1),.din(w_dff_A_zLLi7gXj2_1),.clk(gclk));
	jdff dff_A_tfxBaH2f5_1(.dout(w_dff_A_zLLi7gXj2_1),.din(w_dff_A_tfxBaH2f5_1),.clk(gclk));
	jdff dff_A_NlFA4YzQ5_1(.dout(w_dff_A_tfxBaH2f5_1),.din(w_dff_A_NlFA4YzQ5_1),.clk(gclk));
	jdff dff_A_RpMR2OxI7_1(.dout(w_n77_0[1]),.din(w_dff_A_RpMR2OxI7_1),.clk(gclk));
	jdff dff_A_Aq2G3hRS3_0(.dout(w_G131_0[0]),.din(w_dff_A_Aq2G3hRS3_0),.clk(gclk));
	jdff dff_A_6sZriiSp8_0(.dout(w_dff_A_Aq2G3hRS3_0),.din(w_dff_A_6sZriiSp8_0),.clk(gclk));
	jdff dff_A_rBmApmgP5_0(.dout(w_dff_A_6sZriiSp8_0),.din(w_dff_A_rBmApmgP5_0),.clk(gclk));
	jdff dff_A_G4M8TZ2k6_0(.dout(w_dff_A_rBmApmgP5_0),.din(w_dff_A_G4M8TZ2k6_0),.clk(gclk));
	jdff dff_A_RFjz22497_0(.dout(w_dff_A_G4M8TZ2k6_0),.din(w_dff_A_RFjz22497_0),.clk(gclk));
	jdff dff_A_QCdRjKSu9_0(.dout(w_dff_A_RFjz22497_0),.din(w_dff_A_QCdRjKSu9_0),.clk(gclk));
	jdff dff_A_5HrEIJzf6_0(.dout(w_dff_A_QCdRjKSu9_0),.din(w_dff_A_5HrEIJzf6_0),.clk(gclk));
	jdff dff_A_ZDdsL0xS4_0(.dout(w_dff_A_5HrEIJzf6_0),.din(w_dff_A_ZDdsL0xS4_0),.clk(gclk));
	jdff dff_A_WLj5kph79_0(.dout(w_dff_A_ZDdsL0xS4_0),.din(w_dff_A_WLj5kph79_0),.clk(gclk));
	jdff dff_A_DHFxyEwJ4_0(.dout(w_dff_A_WLj5kph79_0),.din(w_dff_A_DHFxyEwJ4_0),.clk(gclk));
	jdff dff_A_cEYVCbYt4_0(.dout(w_dff_A_DHFxyEwJ4_0),.din(w_dff_A_cEYVCbYt4_0),.clk(gclk));
	jdff dff_A_JyaBcpWa8_0(.dout(w_dff_A_cEYVCbYt4_0),.din(w_dff_A_JyaBcpWa8_0),.clk(gclk));
	jdff dff_A_Hcb55XUz0_0(.dout(w_G137_0[0]),.din(w_dff_A_Hcb55XUz0_0),.clk(gclk));
	jdff dff_A_fq6alYdv7_0(.dout(w_dff_A_Hcb55XUz0_0),.din(w_dff_A_fq6alYdv7_0),.clk(gclk));
	jdff dff_A_36Lp5GWA1_0(.dout(w_dff_A_fq6alYdv7_0),.din(w_dff_A_36Lp5GWA1_0),.clk(gclk));
	jdff dff_A_RKopOPX02_0(.dout(w_dff_A_36Lp5GWA1_0),.din(w_dff_A_RKopOPX02_0),.clk(gclk));
	jdff dff_A_6PoYq1Wu0_0(.dout(w_dff_A_RKopOPX02_0),.din(w_dff_A_6PoYq1Wu0_0),.clk(gclk));
	jdff dff_A_DVrloNLw8_0(.dout(w_dff_A_6PoYq1Wu0_0),.din(w_dff_A_DVrloNLw8_0),.clk(gclk));
	jdff dff_A_BwvDfDsI4_0(.dout(w_dff_A_DVrloNLw8_0),.din(w_dff_A_BwvDfDsI4_0),.clk(gclk));
	jdff dff_A_qmWValbh4_0(.dout(w_dff_A_BwvDfDsI4_0),.din(w_dff_A_qmWValbh4_0),.clk(gclk));
	jdff dff_A_2H4Zhj1s8_0(.dout(w_dff_A_qmWValbh4_0),.din(w_dff_A_2H4Zhj1s8_0),.clk(gclk));
	jdff dff_A_sbStELCV0_0(.dout(w_dff_A_2H4Zhj1s8_0),.din(w_dff_A_sbStELCV0_0),.clk(gclk));
	jdff dff_A_YHUWyG7E9_0(.dout(w_dff_A_sbStELCV0_0),.din(w_dff_A_YHUWyG7E9_0),.clk(gclk));
	jdff dff_A_GtIiwpDE5_2(.dout(w_G137_0[2]),.din(w_dff_A_GtIiwpDE5_2),.clk(gclk));
	jdff dff_A_W5ZQRB9x1_2(.dout(w_dff_A_GtIiwpDE5_2),.din(w_dff_A_W5ZQRB9x1_2),.clk(gclk));
	jdff dff_B_GaHf3EBN6_3(.din(G137),.dout(w_dff_B_GaHf3EBN6_3),.clk(gclk));
	jdff dff_A_vGQfHwSI9_0(.dout(w_G134_0[0]),.din(w_dff_A_vGQfHwSI9_0),.clk(gclk));
	jdff dff_A_xh7XY4I17_0(.dout(w_dff_A_vGQfHwSI9_0),.din(w_dff_A_xh7XY4I17_0),.clk(gclk));
	jdff dff_A_VKKvjeLx6_0(.dout(w_dff_A_xh7XY4I17_0),.din(w_dff_A_VKKvjeLx6_0),.clk(gclk));
	jdff dff_A_mjDFR3ZZ8_0(.dout(w_dff_A_VKKvjeLx6_0),.din(w_dff_A_mjDFR3ZZ8_0),.clk(gclk));
	jdff dff_A_cyVzZvfH3_0(.dout(w_dff_A_mjDFR3ZZ8_0),.din(w_dff_A_cyVzZvfH3_0),.clk(gclk));
	jdff dff_A_zvJDWPJX1_0(.dout(w_dff_A_cyVzZvfH3_0),.din(w_dff_A_zvJDWPJX1_0),.clk(gclk));
	jdff dff_A_rxR4Nddt3_0(.dout(w_dff_A_zvJDWPJX1_0),.din(w_dff_A_rxR4Nddt3_0),.clk(gclk));
	jdff dff_A_0nqpbG9k7_0(.dout(w_dff_A_rxR4Nddt3_0),.din(w_dff_A_0nqpbG9k7_0),.clk(gclk));
	jdff dff_A_7awu9U0n2_0(.dout(w_dff_A_0nqpbG9k7_0),.din(w_dff_A_7awu9U0n2_0),.clk(gclk));
	jdff dff_A_dUMHazyn4_0(.dout(w_dff_A_7awu9U0n2_0),.din(w_dff_A_dUMHazyn4_0),.clk(gclk));
	jdff dff_A_j4u8WWwp4_0(.dout(w_dff_A_dUMHazyn4_0),.din(w_dff_A_j4u8WWwp4_0),.clk(gclk));
	jdff dff_A_UfGRfBbx1_0(.dout(w_dff_A_j4u8WWwp4_0),.din(w_dff_A_UfGRfBbx1_0),.clk(gclk));
	jdff dff_A_YB2zu5zl1_2(.dout(w_dff_A_cdqCJLBY5_0),.din(w_dff_A_YB2zu5zl1_2),.clk(gclk));
	jdff dff_A_cdqCJLBY5_0(.dout(w_dff_A_PSCRMpSH3_0),.din(w_dff_A_cdqCJLBY5_0),.clk(gclk));
	jdff dff_A_PSCRMpSH3_0(.dout(w_dff_A_ZkCaUY862_0),.din(w_dff_A_PSCRMpSH3_0),.clk(gclk));
	jdff dff_A_ZkCaUY862_0(.dout(w_dff_A_oBQTgxkS7_0),.din(w_dff_A_ZkCaUY862_0),.clk(gclk));
	jdff dff_A_oBQTgxkS7_0(.dout(w_dff_A_BpVIvNa50_0),.din(w_dff_A_oBQTgxkS7_0),.clk(gclk));
	jdff dff_A_BpVIvNa50_0(.dout(w_dff_A_mv8Apsd28_0),.din(w_dff_A_BpVIvNa50_0),.clk(gclk));
	jdff dff_A_mv8Apsd28_0(.dout(G3),.din(w_dff_A_mv8Apsd28_0),.clk(gclk));
	jdff dff_A_pQ4XnbpO5_2(.dout(w_dff_A_S1ieWPyR5_0),.din(w_dff_A_pQ4XnbpO5_2),.clk(gclk));
	jdff dff_A_S1ieWPyR5_0(.dout(w_dff_A_mOxFe7am8_0),.din(w_dff_A_S1ieWPyR5_0),.clk(gclk));
	jdff dff_A_mOxFe7am8_0(.dout(w_dff_A_PvAxLKaP0_0),.din(w_dff_A_mOxFe7am8_0),.clk(gclk));
	jdff dff_A_PvAxLKaP0_0(.dout(w_dff_A_uCKgvjuD2_0),.din(w_dff_A_PvAxLKaP0_0),.clk(gclk));
	jdff dff_A_uCKgvjuD2_0(.dout(w_dff_A_VsNLXOon8_0),.din(w_dff_A_uCKgvjuD2_0),.clk(gclk));
	jdff dff_A_VsNLXOon8_0(.dout(w_dff_A_BeQV5WJi1_0),.din(w_dff_A_VsNLXOon8_0),.clk(gclk));
	jdff dff_A_BeQV5WJi1_0(.dout(G6),.din(w_dff_A_BeQV5WJi1_0),.clk(gclk));
	jdff dff_A_ysQrHSkC2_2(.dout(w_dff_A_vN9CF0Gm8_0),.din(w_dff_A_ysQrHSkC2_2),.clk(gclk));
	jdff dff_A_vN9CF0Gm8_0(.dout(w_dff_A_we0ql9Mr0_0),.din(w_dff_A_vN9CF0Gm8_0),.clk(gclk));
	jdff dff_A_we0ql9Mr0_0(.dout(w_dff_A_Vwjcf8eh8_0),.din(w_dff_A_we0ql9Mr0_0),.clk(gclk));
	jdff dff_A_Vwjcf8eh8_0(.dout(w_dff_A_1FVjeGYk7_0),.din(w_dff_A_Vwjcf8eh8_0),.clk(gclk));
	jdff dff_A_1FVjeGYk7_0(.dout(w_dff_A_qYRMynfE0_0),.din(w_dff_A_1FVjeGYk7_0),.clk(gclk));
	jdff dff_A_qYRMynfE0_0(.dout(w_dff_A_cZzKFklK0_0),.din(w_dff_A_qYRMynfE0_0),.clk(gclk));
	jdff dff_A_cZzKFklK0_0(.dout(G9),.din(w_dff_A_cZzKFklK0_0),.clk(gclk));
	jdff dff_A_HmEPIFW31_2(.dout(w_dff_A_Yf84sPaq2_0),.din(w_dff_A_HmEPIFW31_2),.clk(gclk));
	jdff dff_A_Yf84sPaq2_0(.dout(w_dff_A_xBjcXoJg3_0),.din(w_dff_A_Yf84sPaq2_0),.clk(gclk));
	jdff dff_A_xBjcXoJg3_0(.dout(w_dff_A_IUAawD926_0),.din(w_dff_A_xBjcXoJg3_0),.clk(gclk));
	jdff dff_A_IUAawD926_0(.dout(w_dff_A_6ruDch8Q0_0),.din(w_dff_A_IUAawD926_0),.clk(gclk));
	jdff dff_A_6ruDch8Q0_0(.dout(w_dff_A_fhOyMIsJ9_0),.din(w_dff_A_6ruDch8Q0_0),.clk(gclk));
	jdff dff_A_fhOyMIsJ9_0(.dout(w_dff_A_IqqEoIAE2_0),.din(w_dff_A_fhOyMIsJ9_0),.clk(gclk));
	jdff dff_A_IqqEoIAE2_0(.dout(G12),.din(w_dff_A_IqqEoIAE2_0),.clk(gclk));
	jdff dff_A_p6TGz3CQ7_2(.dout(w_dff_A_pcP2slpG1_0),.din(w_dff_A_p6TGz3CQ7_2),.clk(gclk));
	jdff dff_A_pcP2slpG1_0(.dout(w_dff_A_nLrVGHj24_0),.din(w_dff_A_pcP2slpG1_0),.clk(gclk));
	jdff dff_A_nLrVGHj24_0(.dout(w_dff_A_zDjIKNEK5_0),.din(w_dff_A_nLrVGHj24_0),.clk(gclk));
	jdff dff_A_zDjIKNEK5_0(.dout(w_dff_A_ul1jI3C58_0),.din(w_dff_A_zDjIKNEK5_0),.clk(gclk));
	jdff dff_A_ul1jI3C58_0(.dout(w_dff_A_4TF89CR94_0),.din(w_dff_A_ul1jI3C58_0),.clk(gclk));
	jdff dff_A_4TF89CR94_0(.dout(w_dff_A_fZXszqZF7_0),.din(w_dff_A_4TF89CR94_0),.clk(gclk));
	jdff dff_A_fZXszqZF7_0(.dout(G30),.din(w_dff_A_fZXszqZF7_0),.clk(gclk));
	jdff dff_A_PXMQJc3d5_2(.dout(w_dff_A_2N3PY2Gp7_0),.din(w_dff_A_PXMQJc3d5_2),.clk(gclk));
	jdff dff_A_2N3PY2Gp7_0(.dout(w_dff_A_MWnd850Z8_0),.din(w_dff_A_2N3PY2Gp7_0),.clk(gclk));
	jdff dff_A_MWnd850Z8_0(.dout(w_dff_A_q7w0t8Tn7_0),.din(w_dff_A_MWnd850Z8_0),.clk(gclk));
	jdff dff_A_q7w0t8Tn7_0(.dout(w_dff_A_4GBe8whH4_0),.din(w_dff_A_q7w0t8Tn7_0),.clk(gclk));
	jdff dff_A_4GBe8whH4_0(.dout(w_dff_A_9lS6el8A2_0),.din(w_dff_A_4GBe8whH4_0),.clk(gclk));
	jdff dff_A_9lS6el8A2_0(.dout(w_dff_A_rfva3CpZ6_0),.din(w_dff_A_9lS6el8A2_0),.clk(gclk));
	jdff dff_A_rfva3CpZ6_0(.dout(G45),.din(w_dff_A_rfva3CpZ6_0),.clk(gclk));
	jdff dff_A_qNoSiuRR7_2(.dout(w_dff_A_v4RRjfoh9_0),.din(w_dff_A_qNoSiuRR7_2),.clk(gclk));
	jdff dff_A_v4RRjfoh9_0(.dout(w_dff_A_AoCrHRVr9_0),.din(w_dff_A_v4RRjfoh9_0),.clk(gclk));
	jdff dff_A_AoCrHRVr9_0(.dout(w_dff_A_1t0T9EDO3_0),.din(w_dff_A_AoCrHRVr9_0),.clk(gclk));
	jdff dff_A_1t0T9EDO3_0(.dout(w_dff_A_rT5XSn3U7_0),.din(w_dff_A_1t0T9EDO3_0),.clk(gclk));
	jdff dff_A_rT5XSn3U7_0(.dout(w_dff_A_2M8lKHt31_0),.din(w_dff_A_rT5XSn3U7_0),.clk(gclk));
	jdff dff_A_2M8lKHt31_0(.dout(w_dff_A_Mtg6WqcU7_0),.din(w_dff_A_2M8lKHt31_0),.clk(gclk));
	jdff dff_A_Mtg6WqcU7_0(.dout(G48),.din(w_dff_A_Mtg6WqcU7_0),.clk(gclk));
	jdff dff_A_39k7m2jl2_2(.dout(w_dff_A_7qsHetyr7_0),.din(w_dff_A_39k7m2jl2_2),.clk(gclk));
	jdff dff_A_7qsHetyr7_0(.dout(w_dff_A_Hwsv1vYt5_0),.din(w_dff_A_7qsHetyr7_0),.clk(gclk));
	jdff dff_A_Hwsv1vYt5_0(.dout(w_dff_A_hQTMbLAk3_0),.din(w_dff_A_Hwsv1vYt5_0),.clk(gclk));
	jdff dff_A_hQTMbLAk3_0(.dout(w_dff_A_QBRE3wef0_0),.din(w_dff_A_hQTMbLAk3_0),.clk(gclk));
	jdff dff_A_QBRE3wef0_0(.dout(w_dff_A_xgVmC8PK6_0),.din(w_dff_A_QBRE3wef0_0),.clk(gclk));
	jdff dff_A_xgVmC8PK6_0(.dout(w_dff_A_bzv9FnAW3_0),.din(w_dff_A_xgVmC8PK6_0),.clk(gclk));
	jdff dff_A_bzv9FnAW3_0(.dout(G15),.din(w_dff_A_bzv9FnAW3_0),.clk(gclk));
	jdff dff_A_BLmIZlKE0_2(.dout(w_dff_A_i6juiczR6_0),.din(w_dff_A_BLmIZlKE0_2),.clk(gclk));
	jdff dff_A_i6juiczR6_0(.dout(w_dff_A_b8S6KonW0_0),.din(w_dff_A_i6juiczR6_0),.clk(gclk));
	jdff dff_A_b8S6KonW0_0(.dout(w_dff_A_Ft2Yyr073_0),.din(w_dff_A_b8S6KonW0_0),.clk(gclk));
	jdff dff_A_Ft2Yyr073_0(.dout(w_dff_A_mZTqoN8o6_0),.din(w_dff_A_Ft2Yyr073_0),.clk(gclk));
	jdff dff_A_mZTqoN8o6_0(.dout(w_dff_A_GXEhLkSL5_0),.din(w_dff_A_mZTqoN8o6_0),.clk(gclk));
	jdff dff_A_GXEhLkSL5_0(.dout(w_dff_A_FT3qtJPI0_0),.din(w_dff_A_GXEhLkSL5_0),.clk(gclk));
	jdff dff_A_FT3qtJPI0_0(.dout(G18),.din(w_dff_A_FT3qtJPI0_0),.clk(gclk));
	jdff dff_A_gNVWv1vW4_2(.dout(w_dff_A_sATPXdvY4_0),.din(w_dff_A_gNVWv1vW4_2),.clk(gclk));
	jdff dff_A_sATPXdvY4_0(.dout(w_dff_A_F6qhPc3x8_0),.din(w_dff_A_sATPXdvY4_0),.clk(gclk));
	jdff dff_A_F6qhPc3x8_0(.dout(w_dff_A_JQaKlUJk6_0),.din(w_dff_A_F6qhPc3x8_0),.clk(gclk));
	jdff dff_A_JQaKlUJk6_0(.dout(w_dff_A_uP6PnsRX4_0),.din(w_dff_A_JQaKlUJk6_0),.clk(gclk));
	jdff dff_A_uP6PnsRX4_0(.dout(w_dff_A_R4POdEhI4_0),.din(w_dff_A_uP6PnsRX4_0),.clk(gclk));
	jdff dff_A_R4POdEhI4_0(.dout(w_dff_A_VJzf25z71_0),.din(w_dff_A_R4POdEhI4_0),.clk(gclk));
	jdff dff_A_VJzf25z71_0(.dout(G21),.din(w_dff_A_VJzf25z71_0),.clk(gclk));
	jdff dff_A_2UJqkRKI1_2(.dout(w_dff_A_wfNajdZh6_0),.din(w_dff_A_2UJqkRKI1_2),.clk(gclk));
	jdff dff_A_wfNajdZh6_0(.dout(w_dff_A_B7VUIsVW0_0),.din(w_dff_A_wfNajdZh6_0),.clk(gclk));
	jdff dff_A_B7VUIsVW0_0(.dout(w_dff_A_wbhkfoiN6_0),.din(w_dff_A_B7VUIsVW0_0),.clk(gclk));
	jdff dff_A_wbhkfoiN6_0(.dout(w_dff_A_Ivbg4XuS0_0),.din(w_dff_A_wbhkfoiN6_0),.clk(gclk));
	jdff dff_A_Ivbg4XuS0_0(.dout(w_dff_A_xYY1WJmk6_0),.din(w_dff_A_Ivbg4XuS0_0),.clk(gclk));
	jdff dff_A_xYY1WJmk6_0(.dout(w_dff_A_4s4oRm1t2_0),.din(w_dff_A_xYY1WJmk6_0),.clk(gclk));
	jdff dff_A_4s4oRm1t2_0(.dout(G24),.din(w_dff_A_4s4oRm1t2_0),.clk(gclk));
	jdff dff_A_C3HB9a9M2_2(.dout(w_dff_A_W2j5GYVz1_0),.din(w_dff_A_C3HB9a9M2_2),.clk(gclk));
	jdff dff_A_W2j5GYVz1_0(.dout(w_dff_A_UoJPwRW47_0),.din(w_dff_A_W2j5GYVz1_0),.clk(gclk));
	jdff dff_A_UoJPwRW47_0(.dout(w_dff_A_JEpQsdg96_0),.din(w_dff_A_UoJPwRW47_0),.clk(gclk));
	jdff dff_A_JEpQsdg96_0(.dout(w_dff_A_ixsuCzqR1_0),.din(w_dff_A_JEpQsdg96_0),.clk(gclk));
	jdff dff_A_ixsuCzqR1_0(.dout(w_dff_A_pBSzkd7J0_0),.din(w_dff_A_ixsuCzqR1_0),.clk(gclk));
	jdff dff_A_pBSzkd7J0_0(.dout(w_dff_A_Kej9aHSI0_0),.din(w_dff_A_pBSzkd7J0_0),.clk(gclk));
	jdff dff_A_Kej9aHSI0_0(.dout(G27),.din(w_dff_A_Kej9aHSI0_0),.clk(gclk));
	jdff dff_A_m9hGZyC60_2(.dout(w_dff_A_ptNbcEFu4_0),.din(w_dff_A_m9hGZyC60_2),.clk(gclk));
	jdff dff_A_ptNbcEFu4_0(.dout(w_dff_A_6mNYGtf30_0),.din(w_dff_A_ptNbcEFu4_0),.clk(gclk));
	jdff dff_A_6mNYGtf30_0(.dout(w_dff_A_dQ51EN3j7_0),.din(w_dff_A_6mNYGtf30_0),.clk(gclk));
	jdff dff_A_dQ51EN3j7_0(.dout(w_dff_A_q31Gen692_0),.din(w_dff_A_dQ51EN3j7_0),.clk(gclk));
	jdff dff_A_q31Gen692_0(.dout(w_dff_A_VktOMNAv9_0),.din(w_dff_A_q31Gen692_0),.clk(gclk));
	jdff dff_A_VktOMNAv9_0(.dout(w_dff_A_P0wzao6F5_0),.din(w_dff_A_VktOMNAv9_0),.clk(gclk));
	jdff dff_A_P0wzao6F5_0(.dout(G33),.din(w_dff_A_P0wzao6F5_0),.clk(gclk));
	jdff dff_A_l5uqOluA3_2(.dout(w_dff_A_f2h19v173_0),.din(w_dff_A_l5uqOluA3_2),.clk(gclk));
	jdff dff_A_f2h19v173_0(.dout(w_dff_A_z1MIvZhV2_0),.din(w_dff_A_f2h19v173_0),.clk(gclk));
	jdff dff_A_z1MIvZhV2_0(.dout(w_dff_A_UKhPafOI0_0),.din(w_dff_A_z1MIvZhV2_0),.clk(gclk));
	jdff dff_A_UKhPafOI0_0(.dout(w_dff_A_HGATsIzh4_0),.din(w_dff_A_UKhPafOI0_0),.clk(gclk));
	jdff dff_A_HGATsIzh4_0(.dout(w_dff_A_hZTYuz462_0),.din(w_dff_A_HGATsIzh4_0),.clk(gclk));
	jdff dff_A_hZTYuz462_0(.dout(w_dff_A_wTV7cp5M7_0),.din(w_dff_A_hZTYuz462_0),.clk(gclk));
	jdff dff_A_wTV7cp5M7_0(.dout(G36),.din(w_dff_A_wTV7cp5M7_0),.clk(gclk));
	jdff dff_A_Q79VKY0V0_2(.dout(w_dff_A_zDAUhiBr7_0),.din(w_dff_A_Q79VKY0V0_2),.clk(gclk));
	jdff dff_A_zDAUhiBr7_0(.dout(w_dff_A_oOpvw8D26_0),.din(w_dff_A_zDAUhiBr7_0),.clk(gclk));
	jdff dff_A_oOpvw8D26_0(.dout(w_dff_A_v0gXjNc76_0),.din(w_dff_A_oOpvw8D26_0),.clk(gclk));
	jdff dff_A_v0gXjNc76_0(.dout(w_dff_A_6VRRScJ37_0),.din(w_dff_A_v0gXjNc76_0),.clk(gclk));
	jdff dff_A_6VRRScJ37_0(.dout(w_dff_A_AxSq91kA5_0),.din(w_dff_A_6VRRScJ37_0),.clk(gclk));
	jdff dff_A_AxSq91kA5_0(.dout(w_dff_A_rRkmF9Gm9_0),.din(w_dff_A_AxSq91kA5_0),.clk(gclk));
	jdff dff_A_rRkmF9Gm9_0(.dout(G39),.din(w_dff_A_rRkmF9Gm9_0),.clk(gclk));
	jdff dff_A_cx8NO26b9_2(.dout(w_dff_A_U1k4ksCe2_0),.din(w_dff_A_cx8NO26b9_2),.clk(gclk));
	jdff dff_A_U1k4ksCe2_0(.dout(w_dff_A_AZVTyJzx7_0),.din(w_dff_A_U1k4ksCe2_0),.clk(gclk));
	jdff dff_A_AZVTyJzx7_0(.dout(w_dff_A_0HA9kgHt9_0),.din(w_dff_A_AZVTyJzx7_0),.clk(gclk));
	jdff dff_A_0HA9kgHt9_0(.dout(w_dff_A_VfTg2vxP4_0),.din(w_dff_A_0HA9kgHt9_0),.clk(gclk));
	jdff dff_A_VfTg2vxP4_0(.dout(w_dff_A_yEuuE7940_0),.din(w_dff_A_VfTg2vxP4_0),.clk(gclk));
	jdff dff_A_yEuuE7940_0(.dout(w_dff_A_lcECBcc08_0),.din(w_dff_A_yEuuE7940_0),.clk(gclk));
	jdff dff_A_lcECBcc08_0(.dout(G42),.din(w_dff_A_lcECBcc08_0),.clk(gclk));
	jdff dff_A_QcEcVxwy4_2(.dout(G75),.din(w_dff_A_QcEcVxwy4_2),.clk(gclk));
	jdff dff_A_hSV2AnXX1_2(.dout(G69),.din(w_dff_A_hSV2AnXX1_2),.clk(gclk));
	jdff dff_A_hZdDs68H3_2(.dout(w_dff_A_NAhYsgVu5_0),.din(w_dff_A_hZdDs68H3_2),.clk(gclk));
	jdff dff_A_NAhYsgVu5_0(.dout(G72),.din(w_dff_A_NAhYsgVu5_0),.clk(gclk));
endmodule

