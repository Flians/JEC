/*
gf_c6288:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 8046
	jand: 664
	jor: 312

Summary:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 8046
	jand: 664
	jor: 312

The maximum logic level gap of any gate:
	gf_c6288: 57
*/

module gf_c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G1gat_1;
	wire [2:0] w_G1gat_2;
	wire [2:0] w_G1gat_3;
	wire [2:0] w_G1gat_4;
	wire [2:0] w_G1gat_5;
	wire [2:0] w_G1gat_6;
	wire [1:0] w_G1gat_7;
	wire [2:0] w_G18gat_0;
	wire [2:0] w_G18gat_1;
	wire [2:0] w_G18gat_2;
	wire [2:0] w_G18gat_3;
	wire [2:0] w_G18gat_4;
	wire [2:0] w_G18gat_5;
	wire [2:0] w_G18gat_6;
	wire [1:0] w_G18gat_7;
	wire [2:0] w_G35gat_0;
	wire [2:0] w_G35gat_1;
	wire [2:0] w_G35gat_2;
	wire [2:0] w_G35gat_3;
	wire [2:0] w_G35gat_4;
	wire [2:0] w_G35gat_5;
	wire [2:0] w_G35gat_6;
	wire [2:0] w_G35gat_7;
	wire [2:0] w_G52gat_0;
	wire [2:0] w_G52gat_1;
	wire [2:0] w_G52gat_2;
	wire [2:0] w_G52gat_3;
	wire [2:0] w_G52gat_4;
	wire [2:0] w_G52gat_5;
	wire [2:0] w_G52gat_6;
	wire [2:0] w_G52gat_7;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G69gat_1;
	wire [2:0] w_G69gat_2;
	wire [2:0] w_G69gat_3;
	wire [2:0] w_G69gat_4;
	wire [2:0] w_G69gat_5;
	wire [2:0] w_G69gat_6;
	wire [1:0] w_G69gat_7;
	wire [2:0] w_G86gat_0;
	wire [2:0] w_G86gat_1;
	wire [2:0] w_G86gat_2;
	wire [2:0] w_G86gat_3;
	wire [2:0] w_G86gat_4;
	wire [2:0] w_G86gat_5;
	wire [2:0] w_G86gat_6;
	wire [1:0] w_G86gat_7;
	wire [2:0] w_G103gat_0;
	wire [2:0] w_G103gat_1;
	wire [2:0] w_G103gat_2;
	wire [2:0] w_G103gat_3;
	wire [2:0] w_G103gat_4;
	wire [2:0] w_G103gat_5;
	wire [2:0] w_G103gat_6;
	wire [1:0] w_G103gat_7;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G120gat_1;
	wire [2:0] w_G120gat_2;
	wire [2:0] w_G120gat_3;
	wire [2:0] w_G120gat_4;
	wire [2:0] w_G120gat_5;
	wire [2:0] w_G120gat_6;
	wire [1:0] w_G120gat_7;
	wire [2:0] w_G137gat_0;
	wire [2:0] w_G137gat_1;
	wire [2:0] w_G137gat_2;
	wire [2:0] w_G137gat_3;
	wire [2:0] w_G137gat_4;
	wire [2:0] w_G137gat_5;
	wire [2:0] w_G137gat_6;
	wire [1:0] w_G137gat_7;
	wire [2:0] w_G154gat_0;
	wire [2:0] w_G154gat_1;
	wire [2:0] w_G154gat_2;
	wire [2:0] w_G154gat_3;
	wire [2:0] w_G154gat_4;
	wire [2:0] w_G154gat_5;
	wire [2:0] w_G154gat_6;
	wire [1:0] w_G154gat_7;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G171gat_2;
	wire [2:0] w_G171gat_3;
	wire [2:0] w_G171gat_4;
	wire [2:0] w_G171gat_5;
	wire [2:0] w_G171gat_6;
	wire [1:0] w_G171gat_7;
	wire [2:0] w_G188gat_0;
	wire [2:0] w_G188gat_1;
	wire [2:0] w_G188gat_2;
	wire [2:0] w_G188gat_3;
	wire [2:0] w_G188gat_4;
	wire [2:0] w_G188gat_5;
	wire [2:0] w_G188gat_6;
	wire [1:0] w_G188gat_7;
	wire [2:0] w_G205gat_0;
	wire [2:0] w_G205gat_1;
	wire [2:0] w_G205gat_2;
	wire [2:0] w_G205gat_3;
	wire [2:0] w_G205gat_4;
	wire [2:0] w_G205gat_5;
	wire [2:0] w_G205gat_6;
	wire [1:0] w_G205gat_7;
	wire [2:0] w_G222gat_0;
	wire [2:0] w_G222gat_1;
	wire [2:0] w_G222gat_2;
	wire [2:0] w_G222gat_3;
	wire [2:0] w_G222gat_4;
	wire [2:0] w_G222gat_5;
	wire [2:0] w_G222gat_6;
	wire [1:0] w_G222gat_7;
	wire [2:0] w_G239gat_0;
	wire [2:0] w_G239gat_1;
	wire [2:0] w_G239gat_2;
	wire [2:0] w_G239gat_3;
	wire [2:0] w_G239gat_4;
	wire [2:0] w_G239gat_5;
	wire [2:0] w_G239gat_6;
	wire [1:0] w_G239gat_7;
	wire [2:0] w_G256gat_0;
	wire [2:0] w_G256gat_1;
	wire [2:0] w_G256gat_2;
	wire [2:0] w_G256gat_3;
	wire [2:0] w_G256gat_4;
	wire [2:0] w_G256gat_5;
	wire [2:0] w_G256gat_6;
	wire [1:0] w_G256gat_7;
	wire [2:0] w_G273gat_0;
	wire [2:0] w_G273gat_1;
	wire [2:0] w_G273gat_2;
	wire [2:0] w_G273gat_3;
	wire [2:0] w_G273gat_4;
	wire [2:0] w_G273gat_5;
	wire [2:0] w_G273gat_6;
	wire [1:0] w_G273gat_7;
	wire [2:0] w_G290gat_0;
	wire [2:0] w_G290gat_1;
	wire [2:0] w_G290gat_2;
	wire [2:0] w_G290gat_3;
	wire [2:0] w_G290gat_4;
	wire [2:0] w_G290gat_5;
	wire [2:0] w_G290gat_6;
	wire [2:0] w_G290gat_7;
	wire [2:0] w_G307gat_0;
	wire [2:0] w_G307gat_1;
	wire [2:0] w_G307gat_2;
	wire [2:0] w_G307gat_3;
	wire [2:0] w_G307gat_4;
	wire [2:0] w_G307gat_5;
	wire [2:0] w_G307gat_6;
	wire [1:0] w_G307gat_7;
	wire [2:0] w_G324gat_0;
	wire [2:0] w_G324gat_1;
	wire [2:0] w_G324gat_2;
	wire [2:0] w_G324gat_3;
	wire [2:0] w_G324gat_4;
	wire [2:0] w_G324gat_5;
	wire [2:0] w_G324gat_6;
	wire [1:0] w_G324gat_7;
	wire [2:0] w_G341gat_0;
	wire [2:0] w_G341gat_1;
	wire [2:0] w_G341gat_2;
	wire [2:0] w_G341gat_3;
	wire [2:0] w_G341gat_4;
	wire [2:0] w_G341gat_5;
	wire [2:0] w_G341gat_6;
	wire [1:0] w_G341gat_7;
	wire [2:0] w_G358gat_0;
	wire [2:0] w_G358gat_1;
	wire [2:0] w_G358gat_2;
	wire [2:0] w_G358gat_3;
	wire [2:0] w_G358gat_4;
	wire [2:0] w_G358gat_5;
	wire [2:0] w_G358gat_6;
	wire [1:0] w_G358gat_7;
	wire [2:0] w_G375gat_0;
	wire [2:0] w_G375gat_1;
	wire [2:0] w_G375gat_2;
	wire [2:0] w_G375gat_3;
	wire [2:0] w_G375gat_4;
	wire [2:0] w_G375gat_5;
	wire [2:0] w_G375gat_6;
	wire [1:0] w_G375gat_7;
	wire [2:0] w_G392gat_0;
	wire [2:0] w_G392gat_1;
	wire [2:0] w_G392gat_2;
	wire [2:0] w_G392gat_3;
	wire [2:0] w_G392gat_4;
	wire [2:0] w_G392gat_5;
	wire [2:0] w_G392gat_6;
	wire [1:0] w_G392gat_7;
	wire [2:0] w_G409gat_0;
	wire [2:0] w_G409gat_1;
	wire [2:0] w_G409gat_2;
	wire [2:0] w_G409gat_3;
	wire [2:0] w_G409gat_4;
	wire [2:0] w_G409gat_5;
	wire [2:0] w_G409gat_6;
	wire [1:0] w_G409gat_7;
	wire [2:0] w_G426gat_0;
	wire [2:0] w_G426gat_1;
	wire [2:0] w_G426gat_2;
	wire [2:0] w_G426gat_3;
	wire [2:0] w_G426gat_4;
	wire [2:0] w_G426gat_5;
	wire [2:0] w_G426gat_6;
	wire [1:0] w_G426gat_7;
	wire [2:0] w_G443gat_0;
	wire [2:0] w_G443gat_1;
	wire [2:0] w_G443gat_2;
	wire [2:0] w_G443gat_3;
	wire [2:0] w_G443gat_4;
	wire [2:0] w_G443gat_5;
	wire [2:0] w_G443gat_6;
	wire [1:0] w_G443gat_7;
	wire [2:0] w_G460gat_0;
	wire [2:0] w_G460gat_1;
	wire [2:0] w_G460gat_2;
	wire [2:0] w_G460gat_3;
	wire [2:0] w_G460gat_4;
	wire [2:0] w_G460gat_5;
	wire [2:0] w_G460gat_6;
	wire [1:0] w_G460gat_7;
	wire [2:0] w_G477gat_0;
	wire [2:0] w_G477gat_1;
	wire [2:0] w_G477gat_2;
	wire [2:0] w_G477gat_3;
	wire [2:0] w_G477gat_4;
	wire [2:0] w_G477gat_5;
	wire [2:0] w_G477gat_6;
	wire [1:0] w_G477gat_7;
	wire [2:0] w_G494gat_0;
	wire [2:0] w_G494gat_1;
	wire [2:0] w_G494gat_2;
	wire [2:0] w_G494gat_3;
	wire [2:0] w_G494gat_4;
	wire [2:0] w_G494gat_5;
	wire [2:0] w_G494gat_6;
	wire [1:0] w_G494gat_7;
	wire [2:0] w_G511gat_0;
	wire [2:0] w_G511gat_1;
	wire [2:0] w_G511gat_2;
	wire [2:0] w_G511gat_3;
	wire [2:0] w_G511gat_4;
	wire [2:0] w_G511gat_5;
	wire [2:0] w_G511gat_6;
	wire [1:0] w_G511gat_7;
	wire [2:0] w_G528gat_0;
	wire [2:0] w_G528gat_1;
	wire [2:0] w_G528gat_2;
	wire [2:0] w_G528gat_3;
	wire [2:0] w_G528gat_4;
	wire [2:0] w_G528gat_5;
	wire [2:0] w_G528gat_6;
	wire [1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire [1:0] w_n65_0;
	wire [1:0] w_n66_0;
	wire [1:0] w_n67_0;
	wire [1:0] w_n69_0;
	wire [1:0] w_n70_0;
	wire [1:0] w_n75_0;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [2:0] w_n80_0;
	wire [1:0] w_n83_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [1:0] w_n90_0;
	wire [1:0] w_n91_0;
	wire [1:0] w_n93_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n99_0;
	wire [2:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n106_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n112_0;
	wire [2:0] w_n117_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n122_0;
	wire [1:0] w_n123_0;
	wire [1:0] w_n125_0;
	wire [1:0] w_n127_0;
	wire [1:0] w_n128_0;
	wire [1:0] w_n129_0;
	wire [1:0] w_n130_0;
	wire [1:0] w_n132_0;
	wire [1:0] w_n133_0;
	wire [1:0] w_n135_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n141_0;
	wire [2:0] w_n146_0;
	wire [1:0] w_n148_0;
	wire [1:0] w_n152_0;
	wire [1:0] w_n154_0;
	wire [1:0] w_n155_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n157_0;
	wire [1:0] w_n158_0;
	wire [1:0] w_n160_0;
	wire [1:0] w_n161_0;
	wire [1:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [1:0] w_n164_0;
	wire [1:0] w_n165_0;
	wire [1:0] w_n167_0;
	wire [1:0] w_n168_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n175_0;
	wire [1:0] w_n176_0;
	wire [2:0] w_n181_0;
	wire [1:0] w_n183_0;
	wire [1:0] w_n186_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n192_0;
	wire [1:0] w_n194_0;
	wire [1:0] w_n195_0;
	wire [2:0] w_n196_0;
	wire [1:0] w_n198_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n203_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n206_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n209_0;
	wire [1:0] w_n210_0;
	wire [1:0] w_n212_0;
	wire [1:0] w_n217_0;
	wire [1:0] w_n218_0;
	wire [2:0] w_n223_0;
	wire [1:0] w_n225_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n230_0;
	wire [1:0] w_n233_0;
	wire [1:0] w_n235_0;
	wire [1:0] w_n239_0;
	wire [1:0] w_n241_0;
	wire [1:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [1:0] w_n245_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n248_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n250_0;
	wire [1:0] w_n251_0;
	wire [1:0] w_n252_0;
	wire [1:0] w_n253_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n255_0;
	wire [1:0] w_n256_0;
	wire [1:0] w_n258_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n266_0;
	wire [1:0] w_n267_0;
	wire [2:0] w_n272_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n277_0;
	wire [1:0] w_n279_0;
	wire [1:0] w_n282_0;
	wire [1:0] w_n284_0;
	wire [1:0] w_n287_0;
	wire [1:0] w_n289_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n296_0;
	wire [2:0] w_n297_0;
	wire [1:0] w_n299_0;
	wire [1:0] w_n301_0;
	wire [1:0] w_n302_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n304_0;
	wire [1:0] w_n305_0;
	wire [1:0] w_n306_0;
	wire [1:0] w_n307_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n309_0;
	wire [1:0] w_n310_0;
	wire [1:0] w_n311_0;
	wire [1:0] w_n312_0;
	wire [1:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n317_0;
	wire [1:0] w_n322_0;
	wire [1:0] w_n323_0;
	wire [2:0] w_n328_0;
	wire [1:0] w_n330_0;
	wire [1:0] w_n333_0;
	wire [1:0] w_n335_0;
	wire [1:0] w_n338_0;
	wire [1:0] w_n340_0;
	wire [1:0] w_n343_0;
	wire [1:0] w_n345_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n354_0;
	wire [1:0] w_n356_0;
	wire [1:0] w_n357_0;
	wire [2:0] w_n358_0;
	wire [1:0] w_n360_0;
	wire [1:0] w_n362_0;
	wire [1:0] w_n363_0;
	wire [1:0] w_n364_0;
	wire [1:0] w_n365_0;
	wire [1:0] w_n366_0;
	wire [1:0] w_n367_0;
	wire [1:0] w_n368_0;
	wire [1:0] w_n369_0;
	wire [1:0] w_n370_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n373_0;
	wire [1:0] w_n374_0;
	wire [1:0] w_n375_0;
	wire [1:0] w_n377_0;
	wire [1:0] w_n378_0;
	wire [1:0] w_n380_0;
	wire [1:0] w_n385_0;
	wire [1:0] w_n386_0;
	wire [2:0] w_n391_0;
	wire [1:0] w_n393_0;
	wire [1:0] w_n396_0;
	wire [1:0] w_n398_0;
	wire [1:0] w_n401_0;
	wire [1:0] w_n403_0;
	wire [1:0] w_n406_0;
	wire [1:0] w_n408_0;
	wire [1:0] w_n411_0;
	wire [1:0] w_n413_0;
	wire [1:0] w_n416_0;
	wire [1:0] w_n418_0;
	wire [1:0] w_n423_0;
	wire [1:0] w_n425_0;
	wire [1:0] w_n426_0;
	wire [2:0] w_n427_0;
	wire [1:0] w_n429_0;
	wire [1:0] w_n431_0;
	wire [1:0] w_n432_0;
	wire [1:0] w_n433_0;
	wire [1:0] w_n434_0;
	wire [1:0] w_n435_0;
	wire [1:0] w_n436_0;
	wire [1:0] w_n437_0;
	wire [1:0] w_n438_0;
	wire [1:0] w_n439_0;
	wire [1:0] w_n440_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n442_0;
	wire [1:0] w_n443_0;
	wire [1:0] w_n444_0;
	wire [1:0] w_n445_0;
	wire [1:0] w_n446_0;
	wire [1:0] w_n448_0;
	wire [1:0] w_n449_0;
	wire [1:0] w_n451_0;
	wire [1:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [2:0] w_n462_0;
	wire [1:0] w_n464_0;
	wire [1:0] w_n467_0;
	wire [1:0] w_n469_0;
	wire [1:0] w_n472_0;
	wire [1:0] w_n474_0;
	wire [1:0] w_n477_0;
	wire [1:0] w_n479_0;
	wire [1:0] w_n482_0;
	wire [1:0] w_n484_0;
	wire [1:0] w_n487_0;
	wire [1:0] w_n489_0;
	wire [1:0] w_n492_0;
	wire [1:0] w_n494_0;
	wire [1:0] w_n499_0;
	wire [1:0] w_n501_0;
	wire [1:0] w_n502_0;
	wire [2:0] w_n503_0;
	wire [1:0] w_n505_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n508_0;
	wire [1:0] w_n509_0;
	wire [1:0] w_n510_0;
	wire [1:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n513_0;
	wire [1:0] w_n514_0;
	wire [1:0] w_n515_0;
	wire [1:0] w_n516_0;
	wire [1:0] w_n517_0;
	wire [1:0] w_n518_0;
	wire [1:0] w_n519_0;
	wire [1:0] w_n520_0;
	wire [1:0] w_n521_0;
	wire [1:0] w_n522_0;
	wire [1:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [1:0] w_n526_0;
	wire [1:0] w_n527_0;
	wire [1:0] w_n529_0;
	wire [1:0] w_n534_0;
	wire [1:0] w_n535_0;
	wire [2:0] w_n540_0;
	wire [1:0] w_n542_0;
	wire [1:0] w_n545_0;
	wire [1:0] w_n547_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n552_0;
	wire [1:0] w_n555_0;
	wire [1:0] w_n557_0;
	wire [1:0] w_n560_0;
	wire [1:0] w_n562_0;
	wire [1:0] w_n565_0;
	wire [1:0] w_n567_0;
	wire [1:0] w_n570_0;
	wire [1:0] w_n572_0;
	wire [1:0] w_n575_0;
	wire [1:0] w_n577_0;
	wire [1:0] w_n582_0;
	wire [1:0] w_n584_0;
	wire [1:0] w_n585_0;
	wire [2:0] w_n586_0;
	wire [1:0] w_n588_0;
	wire [1:0] w_n590_0;
	wire [1:0] w_n591_0;
	wire [1:0] w_n592_0;
	wire [1:0] w_n593_0;
	wire [1:0] w_n594_0;
	wire [1:0] w_n595_0;
	wire [1:0] w_n596_0;
	wire [1:0] w_n597_0;
	wire [1:0] w_n598_0;
	wire [1:0] w_n599_0;
	wire [1:0] w_n600_0;
	wire [1:0] w_n601_0;
	wire [1:0] w_n602_0;
	wire [1:0] w_n603_0;
	wire [1:0] w_n604_0;
	wire [1:0] w_n605_0;
	wire [1:0] w_n606_0;
	wire [1:0] w_n607_0;
	wire [1:0] w_n608_0;
	wire [1:0] w_n609_0;
	wire [1:0] w_n611_0;
	wire [1:0] w_n612_0;
	wire [1:0] w_n614_0;
	wire [1:0] w_n619_0;
	wire [1:0] w_n620_0;
	wire [2:0] w_n625_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n630_0;
	wire [1:0] w_n632_0;
	wire [1:0] w_n635_0;
	wire [1:0] w_n637_0;
	wire [1:0] w_n640_0;
	wire [1:0] w_n642_0;
	wire [1:0] w_n645_0;
	wire [1:0] w_n647_0;
	wire [1:0] w_n650_0;
	wire [1:0] w_n652_0;
	wire [1:0] w_n655_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n660_0;
	wire [1:0] w_n662_0;
	wire [1:0] w_n665_0;
	wire [1:0] w_n667_0;
	wire [1:0] w_n672_0;
	wire [1:0] w_n674_0;
	wire [1:0] w_n675_0;
	wire [2:0] w_n676_0;
	wire [1:0] w_n678_0;
	wire [1:0] w_n680_0;
	wire [1:0] w_n681_0;
	wire [1:0] w_n682_0;
	wire [1:0] w_n683_0;
	wire [1:0] w_n684_0;
	wire [1:0] w_n685_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n688_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n690_0;
	wire [1:0] w_n691_0;
	wire [1:0] w_n692_0;
	wire [1:0] w_n693_0;
	wire [1:0] w_n694_0;
	wire [1:0] w_n695_0;
	wire [1:0] w_n696_0;
	wire [1:0] w_n697_0;
	wire [1:0] w_n698_0;
	wire [1:0] w_n699_0;
	wire [1:0] w_n700_0;
	wire [1:0] w_n701_0;
	wire [1:0] w_n703_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n706_0;
	wire [1:0] w_n711_0;
	wire [1:0] w_n712_0;
	wire [2:0] w_n717_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n722_0;
	wire [1:0] w_n724_0;
	wire [1:0] w_n727_0;
	wire [1:0] w_n729_0;
	wire [1:0] w_n732_0;
	wire [1:0] w_n734_0;
	wire [1:0] w_n737_0;
	wire [1:0] w_n739_0;
	wire [1:0] w_n742_0;
	wire [1:0] w_n744_0;
	wire [1:0] w_n747_0;
	wire [1:0] w_n749_0;
	wire [1:0] w_n752_0;
	wire [1:0] w_n754_0;
	wire [1:0] w_n757_0;
	wire [1:0] w_n759_0;
	wire [1:0] w_n762_0;
	wire [1:0] w_n764_0;
	wire [1:0] w_n769_0;
	wire [1:0] w_n771_0;
	wire [1:0] w_n772_0;
	wire [1:0] w_n773_0;
	wire [1:0] w_n774_0;
	wire [1:0] w_n775_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n778_0;
	wire [1:0] w_n779_0;
	wire [1:0] w_n780_0;
	wire [1:0] w_n781_0;
	wire [1:0] w_n782_0;
	wire [1:0] w_n783_0;
	wire [1:0] w_n784_0;
	wire [1:0] w_n785_0;
	wire [1:0] w_n786_0;
	wire [1:0] w_n787_0;
	wire [1:0] w_n788_0;
	wire [1:0] w_n789_0;
	wire [1:0] w_n790_0;
	wire [1:0] w_n791_0;
	wire [1:0] w_n792_0;
	wire [1:0] w_n793_0;
	wire [1:0] w_n794_0;
	wire [1:0] w_n795_0;
	wire [1:0] w_n796_0;
	wire [1:0] w_n797_0;
	wire [1:0] w_n798_0;
	wire [1:0] w_n799_0;
	wire [1:0] w_n800_0;
	wire [1:0] w_n802_0;
	wire [1:0] w_n803_0;
	wire [1:0] w_n805_0;
	wire [1:0] w_n810_0;
	wire [1:0] w_n811_0;
	wire [1:0] w_n815_0;
	wire [1:0] w_n816_0;
	wire [2:0] w_n820_0;
	wire [1:0] w_n822_0;
	wire [1:0] w_n825_0;
	wire [1:0] w_n827_0;
	wire [1:0] w_n830_0;
	wire [1:0] w_n832_0;
	wire [1:0] w_n835_0;
	wire [1:0] w_n837_0;
	wire [1:0] w_n840_0;
	wire [1:0] w_n842_0;
	wire [1:0] w_n845_0;
	wire [1:0] w_n847_0;
	wire [1:0] w_n850_0;
	wire [1:0] w_n852_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n857_0;
	wire [1:0] w_n860_0;
	wire [1:0] w_n862_0;
	wire [1:0] w_n865_0;
	wire [1:0] w_n867_0;
	wire [1:0] w_n872_0;
	wire [1:0] w_n874_0;
	wire [1:0] w_n875_0;
	wire [1:0] w_n877_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n880_0;
	wire [1:0] w_n881_0;
	wire [1:0] w_n882_0;
	wire [1:0] w_n883_0;
	wire [1:0] w_n884_0;
	wire [1:0] w_n885_0;
	wire [1:0] w_n886_0;
	wire [1:0] w_n887_0;
	wire [1:0] w_n888_0;
	wire [1:0] w_n889_0;
	wire [1:0] w_n890_0;
	wire [1:0] w_n891_0;
	wire [1:0] w_n892_0;
	wire [1:0] w_n893_0;
	wire [1:0] w_n894_0;
	wire [1:0] w_n895_0;
	wire [1:0] w_n896_0;
	wire [1:0] w_n897_0;
	wire [1:0] w_n898_0;
	wire [1:0] w_n899_0;
	wire [2:0] w_n900_0;
	wire [1:0] w_n902_0;
	wire [1:0] w_n903_0;
	wire [1:0] w_n904_0;
	wire [1:0] w_n905_0;
	wire [1:0] w_n910_0;
	wire [1:0] w_n911_0;
	wire [2:0] w_n915_0;
	wire [1:0] w_n916_0;
	wire [1:0] w_n922_0;
	wire [1:0] w_n924_0;
	wire [1:0] w_n927_0;
	wire [1:0] w_n929_0;
	wire [1:0] w_n932_0;
	wire [1:0] w_n934_0;
	wire [1:0] w_n937_0;
	wire [1:0] w_n939_0;
	wire [1:0] w_n942_0;
	wire [1:0] w_n944_0;
	wire [1:0] w_n947_0;
	wire [1:0] w_n949_0;
	wire [1:0] w_n952_0;
	wire [1:0] w_n954_0;
	wire [1:0] w_n957_0;
	wire [1:0] w_n959_0;
	wire [1:0] w_n962_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n967_0;
	wire [1:0] w_n969_0;
	wire [1:0] w_n972_0;
	wire [1:0] w_n974_0;
	wire [1:0] w_n978_0;
	wire [1:0] w_n980_0;
	wire [1:0] w_n982_0;
	wire [1:0] w_n983_0;
	wire [1:0] w_n984_0;
	wire [1:0] w_n985_0;
	wire [1:0] w_n986_0;
	wire [1:0] w_n987_0;
	wire [1:0] w_n988_0;
	wire [1:0] w_n989_0;
	wire [1:0] w_n990_0;
	wire [1:0] w_n991_0;
	wire [1:0] w_n992_0;
	wire [1:0] w_n993_0;
	wire [1:0] w_n994_0;
	wire [1:0] w_n995_0;
	wire [1:0] w_n996_0;
	wire [1:0] w_n997_0;
	wire [1:0] w_n998_0;
	wire [1:0] w_n999_0;
	wire [1:0] w_n1000_0;
	wire [1:0] w_n1001_0;
	wire [1:0] w_n1002_0;
	wire [1:0] w_n1003_0;
	wire [1:0] w_n1004_0;
	wire [1:0] w_n1005_0;
	wire [1:0] w_n1006_0;
	wire [1:0] w_n1007_0;
	wire [1:0] w_n1008_0;
	wire [1:0] w_n1009_0;
	wire [1:0] w_n1011_0;
	wire [1:0] w_n1013_0;
	wire [1:0] w_n1017_0;
	wire [1:0] w_n1018_0;
	wire [1:0] w_n1022_0;
	wire [1:0] w_n1023_0;
	wire [1:0] w_n1026_0;
	wire [1:0] w_n1028_0;
	wire [1:0] w_n1031_0;
	wire [1:0] w_n1033_0;
	wire [1:0] w_n1036_0;
	wire [1:0] w_n1038_0;
	wire [1:0] w_n1041_0;
	wire [1:0] w_n1043_0;
	wire [1:0] w_n1046_0;
	wire [1:0] w_n1048_0;
	wire [1:0] w_n1051_0;
	wire [1:0] w_n1053_0;
	wire [1:0] w_n1056_0;
	wire [1:0] w_n1058_0;
	wire [1:0] w_n1061_0;
	wire [1:0] w_n1063_0;
	wire [1:0] w_n1066_0;
	wire [1:0] w_n1068_0;
	wire [1:0] w_n1071_0;
	wire [1:0] w_n1073_0;
	wire [1:0] w_n1076_0;
	wire [1:0] w_n1077_0;
	wire [1:0] w_n1078_0;
	wire [1:0] w_n1080_0;
	wire [1:0] w_n1082_0;
	wire [1:0] w_n1083_0;
	wire [1:0] w_n1084_0;
	wire [1:0] w_n1085_0;
	wire [1:0] w_n1086_0;
	wire [1:0] w_n1087_0;
	wire [1:0] w_n1088_0;
	wire [1:0] w_n1089_0;
	wire [1:0] w_n1090_0;
	wire [1:0] w_n1091_0;
	wire [1:0] w_n1092_0;
	wire [1:0] w_n1093_0;
	wire [1:0] w_n1094_0;
	wire [1:0] w_n1095_0;
	wire [1:0] w_n1096_0;
	wire [1:0] w_n1097_0;
	wire [1:0] w_n1098_0;
	wire [1:0] w_n1099_0;
	wire [1:0] w_n1100_0;
	wire [1:0] w_n1101_0;
	wire [1:0] w_n1102_0;
	wire [1:0] w_n1103_0;
	wire [1:0] w_n1105_0;
	wire [1:0] w_n1106_0;
	wire [1:0] w_n1107_0;
	wire [1:0] w_n1108_0;
	wire [1:0] w_n1109_0;
	wire [1:0] w_n1115_0;
	wire [1:0] w_n1119_0;
	wire [1:0] w_n1120_0;
	wire [1:0] w_n1124_0;
	wire [1:0] w_n1126_0;
	wire [1:0] w_n1129_0;
	wire [1:0] w_n1131_0;
	wire [1:0] w_n1134_0;
	wire [1:0] w_n1136_0;
	wire [1:0] w_n1139_0;
	wire [1:0] w_n1141_0;
	wire [1:0] w_n1144_0;
	wire [1:0] w_n1146_0;
	wire [1:0] w_n1149_0;
	wire [1:0] w_n1151_0;
	wire [1:0] w_n1154_0;
	wire [1:0] w_n1156_0;
	wire [1:0] w_n1159_0;
	wire [1:0] w_n1161_0;
	wire [1:0] w_n1164_0;
	wire [1:0] w_n1166_0;
	wire [1:0] w_n1169_0;
	wire [1:0] w_n1171_0;
	wire [1:0] w_n1174_0;
	wire [1:0] w_n1175_0;
	wire [1:0] w_n1176_0;
	wire [1:0] w_n1179_0;
	wire [1:0] w_n1181_0;
	wire [1:0] w_n1182_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1184_0;
	wire [1:0] w_n1185_0;
	wire [1:0] w_n1186_0;
	wire [1:0] w_n1187_0;
	wire [1:0] w_n1188_0;
	wire [1:0] w_n1189_0;
	wire [1:0] w_n1190_0;
	wire [1:0] w_n1191_0;
	wire [1:0] w_n1192_0;
	wire [1:0] w_n1193_0;
	wire [1:0] w_n1194_0;
	wire [1:0] w_n1195_0;
	wire [1:0] w_n1196_0;
	wire [1:0] w_n1197_0;
	wire [1:0] w_n1198_0;
	wire [1:0] w_n1199_0;
	wire [1:0] w_n1200_0;
	wire [1:0] w_n1201_0;
	wire [1:0] w_n1203_0;
	wire [1:0] w_n1205_0;
	wire [1:0] w_n1206_0;
	wire [1:0] w_n1207_0;
	wire [1:0] w_n1213_0;
	wire [1:0] w_n1216_0;
	wire [1:0] w_n1217_0;
	wire [1:0] w_n1220_0;
	wire [1:0] w_n1222_0;
	wire [1:0] w_n1225_0;
	wire [1:0] w_n1227_0;
	wire [1:0] w_n1230_0;
	wire [1:0] w_n1232_0;
	wire [1:0] w_n1235_0;
	wire [1:0] w_n1237_0;
	wire [1:0] w_n1240_0;
	wire [1:0] w_n1242_0;
	wire [1:0] w_n1245_0;
	wire [1:0] w_n1247_0;
	wire [1:0] w_n1250_0;
	wire [1:0] w_n1252_0;
	wire [1:0] w_n1255_0;
	wire [1:0] w_n1257_0;
	wire [1:0] w_n1260_0;
	wire [1:0] w_n1262_0;
	wire [1:0] w_n1265_0;
	wire [1:0] w_n1266_0;
	wire [1:0] w_n1267_0;
	wire [1:0] w_n1270_0;
	wire [1:0] w_n1272_0;
	wire [1:0] w_n1273_0;
	wire [1:0] w_n1274_0;
	wire [1:0] w_n1275_0;
	wire [1:0] w_n1276_0;
	wire [1:0] w_n1277_0;
	wire [1:0] w_n1278_0;
	wire [1:0] w_n1279_0;
	wire [1:0] w_n1280_0;
	wire [1:0] w_n1281_0;
	wire [1:0] w_n1282_0;
	wire [1:0] w_n1283_0;
	wire [1:0] w_n1284_0;
	wire [1:0] w_n1285_0;
	wire [1:0] w_n1286_0;
	wire [1:0] w_n1287_0;
	wire [1:0] w_n1288_0;
	wire [1:0] w_n1289_0;
	wire [1:0] w_n1290_0;
	wire [1:0] w_n1291_0;
	wire [1:0] w_n1293_0;
	wire [1:0] w_n1294_0;
	wire [1:0] w_n1295_0;
	wire [1:0] w_n1301_0;
	wire [1:0] w_n1306_0;
	wire [1:0] w_n1307_0;
	wire [1:0] w_n1310_0;
	wire [1:0] w_n1312_0;
	wire [1:0] w_n1315_0;
	wire [1:0] w_n1317_0;
	wire [1:0] w_n1320_0;
	wire [1:0] w_n1322_0;
	wire [1:0] w_n1325_0;
	wire [1:0] w_n1327_0;
	wire [1:0] w_n1330_0;
	wire [1:0] w_n1332_0;
	wire [1:0] w_n1335_0;
	wire [1:0] w_n1337_0;
	wire [1:0] w_n1340_0;
	wire [1:0] w_n1342_0;
	wire [1:0] w_n1345_0;
	wire [1:0] w_n1347_0;
	wire [1:0] w_n1350_0;
	wire [1:0] w_n1351_0;
	wire [1:0] w_n1352_0;
	wire [1:0] w_n1355_0;
	wire [1:0] w_n1357_0;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1359_0;
	wire [1:0] w_n1360_0;
	wire [1:0] w_n1361_0;
	wire [1:0] w_n1362_0;
	wire [1:0] w_n1363_0;
	wire [1:0] w_n1364_0;
	wire [1:0] w_n1365_0;
	wire [1:0] w_n1366_0;
	wire [1:0] w_n1367_0;
	wire [1:0] w_n1368_0;
	wire [1:0] w_n1369_0;
	wire [1:0] w_n1370_0;
	wire [1:0] w_n1371_0;
	wire [1:0] w_n1372_0;
	wire [1:0] w_n1373_0;
	wire [1:0] w_n1374_0;
	wire [1:0] w_n1376_0;
	wire [1:0] w_n1378_0;
	wire [1:0] w_n1379_0;
	wire [1:0] w_n1384_0;
	wire [1:0] w_n1389_0;
	wire [1:0] w_n1390_0;
	wire [1:0] w_n1393_0;
	wire [1:0] w_n1395_0;
	wire [1:0] w_n1398_0;
	wire [1:0] w_n1400_0;
	wire [1:0] w_n1403_0;
	wire [1:0] w_n1405_0;
	wire [1:0] w_n1408_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1413_0;
	wire [1:0] w_n1415_0;
	wire [1:0] w_n1418_0;
	wire [1:0] w_n1420_0;
	wire [1:0] w_n1423_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1428_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1430_0;
	wire [1:0] w_n1433_0;
	wire [1:0] w_n1435_0;
	wire [1:0] w_n1436_0;
	wire [1:0] w_n1437_0;
	wire [1:0] w_n1438_0;
	wire [1:0] w_n1439_0;
	wire [1:0] w_n1440_0;
	wire [1:0] w_n1441_0;
	wire [1:0] w_n1442_0;
	wire [1:0] w_n1443_0;
	wire [1:0] w_n1444_0;
	wire [1:0] w_n1445_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1447_0;
	wire [1:0] w_n1448_0;
	wire [1:0] w_n1449_0;
	wire [1:0] w_n1450_0;
	wire [1:0] w_n1452_0;
	wire [1:0] w_n1454_0;
	wire [1:0] w_n1455_0;
	wire [1:0] w_n1460_0;
	wire [1:0] w_n1465_0;
	wire [1:0] w_n1466_0;
	wire [1:0] w_n1469_0;
	wire [1:0] w_n1471_0;
	wire [1:0] w_n1474_0;
	wire [1:0] w_n1476_0;
	wire [1:0] w_n1479_0;
	wire [1:0] w_n1481_0;
	wire [1:0] w_n1484_0;
	wire [1:0] w_n1486_0;
	wire [1:0] w_n1489_0;
	wire [1:0] w_n1491_0;
	wire [1:0] w_n1494_0;
	wire [1:0] w_n1496_0;
	wire [1:0] w_n1499_0;
	wire [1:0] w_n1500_0;
	wire [1:0] w_n1501_0;
	wire [1:0] w_n1504_0;
	wire [1:0] w_n1506_0;
	wire [1:0] w_n1507_0;
	wire [1:0] w_n1508_0;
	wire [1:0] w_n1509_0;
	wire [1:0] w_n1510_0;
	wire [1:0] w_n1511_0;
	wire [1:0] w_n1512_0;
	wire [1:0] w_n1513_0;
	wire [1:0] w_n1514_0;
	wire [1:0] w_n1515_0;
	wire [1:0] w_n1516_0;
	wire [1:0] w_n1517_0;
	wire [1:0] w_n1518_0;
	wire [1:0] w_n1519_0;
	wire [1:0] w_n1521_0;
	wire [1:0] w_n1523_0;
	wire [1:0] w_n1524_0;
	wire [1:0] w_n1529_0;
	wire [1:0] w_n1534_0;
	wire [1:0] w_n1535_0;
	wire [1:0] w_n1538_0;
	wire [1:0] w_n1540_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1548_0;
	wire [1:0] w_n1550_0;
	wire [1:0] w_n1553_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1558_0;
	wire [1:0] w_n1560_0;
	wire [1:0] w_n1563_0;
	wire [1:0] w_n1564_0;
	wire [1:0] w_n1565_0;
	wire [1:0] w_n1568_0;
	wire [1:0] w_n1570_0;
	wire [1:0] w_n1571_0;
	wire [1:0] w_n1572_0;
	wire [1:0] w_n1573_0;
	wire [1:0] w_n1574_0;
	wire [1:0] w_n1575_0;
	wire [1:0] w_n1576_0;
	wire [1:0] w_n1577_0;
	wire [1:0] w_n1578_0;
	wire [1:0] w_n1579_0;
	wire [1:0] w_n1580_0;
	wire [1:0] w_n1581_0;
	wire [1:0] w_n1583_0;
	wire [1:0] w_n1585_0;
	wire [1:0] w_n1586_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1597_0;
	wire [1:0] w_n1600_0;
	wire [1:0] w_n1602_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1607_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1612_0;
	wire [1:0] w_n1615_0;
	wire [1:0] w_n1617_0;
	wire [1:0] w_n1620_0;
	wire [1:0] w_n1621_0;
	wire [1:0] w_n1622_0;
	wire [1:0] w_n1625_0;
	wire [1:0] w_n1627_0;
	wire [1:0] w_n1628_0;
	wire [1:0] w_n1629_0;
	wire [1:0] w_n1630_0;
	wire [1:0] w_n1631_0;
	wire [1:0] w_n1632_0;
	wire [1:0] w_n1633_0;
	wire [1:0] w_n1634_0;
	wire [1:0] w_n1635_0;
	wire [1:0] w_n1636_0;
	wire [1:0] w_n1638_0;
	wire [1:0] w_n1640_0;
	wire [1:0] w_n1641_0;
	wire [1:0] w_n1646_0;
	wire [1:0] w_n1651_0;
	wire [1:0] w_n1653_0;
	wire [1:0] w_n1656_0;
	wire [1:0] w_n1658_0;
	wire [1:0] w_n1661_0;
	wire [1:0] w_n1663_0;
	wire [1:0] w_n1666_0;
	wire [1:0] w_n1668_0;
	wire [1:0] w_n1671_0;
	wire [1:0] w_n1672_0;
	wire [1:0] w_n1673_0;
	wire [1:0] w_n1676_0;
	wire [1:0] w_n1678_0;
	wire [1:0] w_n1679_0;
	wire [1:0] w_n1680_0;
	wire [1:0] w_n1681_0;
	wire [1:0] w_n1682_0;
	wire [1:0] w_n1683_0;
	wire [1:0] w_n1684_0;
	wire [1:0] w_n1685_0;
	wire [1:0] w_n1686_0;
	wire [1:0] w_n1688_0;
	wire [1:0] w_n1689_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1697_0;
	wire [1:0] w_n1699_0;
	wire [1:0] w_n1702_0;
	wire [1:0] w_n1704_0;
	wire [1:0] w_n1707_0;
	wire [1:0] w_n1709_0;
	wire [1:0] w_n1712_0;
	wire [1:0] w_n1713_0;
	wire [1:0] w_n1714_0;
	wire [1:0] w_n1717_0;
	wire [1:0] w_n1719_0;
	wire [1:0] w_n1720_0;
	wire [1:0] w_n1721_0;
	wire [1:0] w_n1722_0;
	wire [1:0] w_n1723_0;
	wire [1:0] w_n1724_0;
	wire [1:0] w_n1725_0;
	wire [1:0] w_n1726_0;
	wire [1:0] w_n1727_0;
	wire [1:0] w_n1734_0;
	wire [1:0] w_n1737_0;
	wire [1:0] w_n1739_0;
	wire [1:0] w_n1742_0;
	wire [1:0] w_n1744_0;
	wire [1:0] w_n1747_0;
	wire [1:0] w_n1748_0;
	wire [1:0] w_n1749_0;
	wire [1:0] w_n1752_0;
	wire [1:0] w_n1754_0;
	wire [1:0] w_n1755_0;
	wire [1:0] w_n1756_0;
	wire [1:0] w_n1757_0;
	wire [1:0] w_n1758_0;
	wire [1:0] w_n1759_0;
	wire [1:0] w_n1760_0;
	wire [1:0] w_n1767_0;
	wire [1:0] w_n1770_0;
	wire [1:0] w_n1772_0;
	wire [1:0] w_n1775_0;
	wire [1:0] w_n1776_0;
	wire [1:0] w_n1777_0;
	wire [1:0] w_n1780_0;
	wire [1:0] w_n1782_0;
	wire [1:0] w_n1783_0;
	wire [1:0] w_n1784_0;
	wire [1:0] w_n1785_0;
	wire [1:0] w_n1786_0;
	wire [1:0] w_n1793_0;
	wire [1:0] w_n1796_0;
	wire [1:0] w_n1797_0;
	wire [1:0] w_n1798_0;
	wire [1:0] w_n1801_0;
	wire [1:0] w_n1803_0;
	wire [1:0] w_n1804_0;
	wire [1:0] w_n1805_0;
	wire [1:0] w_n1807_0;
	wire [1:0] w_n1810_0;
	wire [1:0] w_n1817_0;
	wire [1:0] w_n1818_0;
	wire w_dff_B_CQzbtU104_0;
	wire w_dff_B_lEuxbv5F0_0;
	wire w_dff_B_m2YFsOFD9_1;
	wire w_dff_B_b2YnYtSV1_1;
	wire w_dff_B_5LuDeCfj3_1;
	wire w_dff_B_WFVxcR7l8_1;
	wire w_dff_B_A4lZUm4M2_1;
	wire w_dff_B_6FQXuesw2_1;
	wire w_dff_B_0gcEPcrz3_1;
	wire w_dff_B_KvMrhP0T4_1;
	wire w_dff_B_HfeP3lcw0_1;
	wire w_dff_B_i8xu0OGh6_1;
	wire w_dff_B_OQQcgr6h1_1;
	wire w_dff_B_q9eLr02q1_1;
	wire w_dff_B_I3Ru0P1g5_1;
	wire w_dff_B_7YBUKEnd7_1;
	wire w_dff_B_Zkre0t9S8_1;
	wire w_dff_B_QCM5rOcm5_1;
	wire w_dff_B_vmjV8cet6_1;
	wire w_dff_B_k71p4s1n3_1;
	wire w_dff_B_HH8HPvVI0_1;
	wire w_dff_B_QqQK8s0U3_1;
	wire w_dff_B_kCeu8XBG1_1;
	wire w_dff_B_dxQzISG90_1;
	wire w_dff_B_FGCQnwCp5_1;
	wire w_dff_B_1CSPJc2a0_1;
	wire w_dff_B_uPvNFZ5c1_1;
	wire w_dff_B_BNbxdmAq4_1;
	wire w_dff_B_tBwCKQwe8_1;
	wire w_dff_B_DPQZ5tvD5_1;
	wire w_dff_B_fqpEbCij6_1;
	wire w_dff_B_PcDM2u6M1_1;
	wire w_dff_B_yAJYlebs5_1;
	wire w_dff_B_L9zoaLbS3_1;
	wire w_dff_B_ZF4KR1sm0_1;
	wire w_dff_B_IUAIBhO16_1;
	wire w_dff_B_zZlEm5fz8_1;
	wire w_dff_B_vjaNgyfC6_1;
	wire w_dff_B_U7jcckH96_1;
	wire w_dff_B_kWtxciCH1_1;
	wire w_dff_B_cL18KVjY0_1;
	wire w_dff_B_5OBCqHq93_1;
	wire w_dff_B_SFJx1Xso7_1;
	wire w_dff_B_Kja5SFmP6_1;
	wire w_dff_B_tYDsVwD79_1;
	wire w_dff_B_r7koO1Cd2_1;
	wire w_dff_B_5lzuWr6g6_1;
	wire w_dff_B_rvQUMrX54_1;
	wire w_dff_B_lXCG7Vdi4_1;
	wire w_dff_B_QcjPscN71_1;
	wire w_dff_B_8Z8mEQet0_1;
	wire w_dff_B_vqGt22TA8_1;
	wire w_dff_B_buYVPwG02_1;
	wire w_dff_B_axfIYrza8_1;
	wire w_dff_B_GcG9iY9w2_1;
	wire w_dff_B_bOkHvbh19_1;
	wire w_dff_B_DVNXvqNt3_1;
	wire w_dff_B_HqbXxAvh1_1;
	wire w_dff_B_OAhj6Tw48_1;
	wire w_dff_B_aRs7Cx5P3_1;
	wire w_dff_B_wZ0tyaKd6_1;
	wire w_dff_B_ZY3QDktq1_1;
	wire w_dff_B_9qnEvK782_1;
	wire w_dff_B_gPfvKI8H1_1;
	wire w_dff_B_so7U7eC87_1;
	wire w_dff_B_BUyvwPbb1_1;
	wire w_dff_B_elVOzZ7q4_1;
	wire w_dff_B_Vh7Y9NNi4_1;
	wire w_dff_B_JULEhToh9_1;
	wire w_dff_B_ZH3oGxlj7_1;
	wire w_dff_B_xsy6icMC9_1;
	wire w_dff_B_WTuFu6Cv4_1;
	wire w_dff_B_cRFxGYkK1_1;
	wire w_dff_B_AgMqf6K30_1;
	wire w_dff_B_XYW3L56N0_1;
	wire w_dff_B_lQf1FyrY4_1;
	wire w_dff_B_CLGPZbuj3_1;
	wire w_dff_B_4CV3vP6I7_1;
	wire w_dff_B_RUUqzdH85_1;
	wire w_dff_B_A4zxo8ba5_1;
	wire w_dff_B_PkSuJ1jH0_1;
	wire w_dff_B_IwnpOftq1_1;
	wire w_dff_B_rgS15Ok66_1;
	wire w_dff_B_EpuBHSCh7_1;
	wire w_dff_B_0esQzCRK8_1;
	wire w_dff_B_m3PEL1Gm3_1;
	wire w_dff_B_om5yi6oo6_1;
	wire w_dff_B_RNaMrRvH6_1;
	wire w_dff_B_SENSpIqz4_1;
	wire w_dff_B_P9Uq7ySz0_1;
	wire w_dff_B_gGLWvwHE0_1;
	wire w_dff_B_5xawmo587_1;
	wire w_dff_B_HF85Sorq0_1;
	wire w_dff_B_McV18ixf3_1;
	wire w_dff_B_tspBcsNe5_1;
	wire w_dff_B_8KvmIXAE4_1;
	wire w_dff_B_1PlvDrQ21_1;
	wire w_dff_B_RRqtvSfw5_1;
	wire w_dff_B_nSHEtc8K3_1;
	wire w_dff_B_p4kuG29k6_1;
	wire w_dff_B_dd5qWz7c1_1;
	wire w_dff_B_G8juxv5v1_1;
	wire w_dff_B_s2YN9vxX1_1;
	wire w_dff_B_5YcMWnSx7_1;
	wire w_dff_B_GfcNu1Pm8_1;
	wire w_dff_B_Q0U8vNiJ5_1;
	wire w_dff_B_RTNinQqY8_1;
	wire w_dff_B_xgb81Vz88_1;
	wire w_dff_B_RoA3tBvL4_1;
	wire w_dff_B_vGQOMZBB4_1;
	wire w_dff_B_1thrLE4J6_1;
	wire w_dff_B_d6xtxwtY7_1;
	wire w_dff_B_pBJyrQGT0_1;
	wire w_dff_B_zfMrTPdX8_1;
	wire w_dff_B_rqsZCN590_1;
	wire w_dff_B_RgPVaUv77_1;
	wire w_dff_B_2YqoXrLH1_1;
	wire w_dff_B_oRoaPbra3_1;
	wire w_dff_B_xaVLPsu49_1;
	wire w_dff_B_wQlgNhLa9_1;
	wire w_dff_B_WrfQEx1C9_1;
	wire w_dff_B_Sd5vFueX7_1;
	wire w_dff_B_SN7GOMXW4_1;
	wire w_dff_B_fK4bgWEk7_1;
	wire w_dff_B_fW7d0Ilt6_1;
	wire w_dff_B_Uq6KDSWv2_1;
	wire w_dff_B_JW9BKxOH9_1;
	wire w_dff_B_JV781Cy01_1;
	wire w_dff_B_bY10uaJ73_1;
	wire w_dff_B_sgIQiEtB3_1;
	wire w_dff_B_C2SNLFqJ7_1;
	wire w_dff_B_ahZNrPcM3_1;
	wire w_dff_B_PRVmNAZi2_1;
	wire w_dff_B_JoZcubzt1_1;
	wire w_dff_B_n3g5oXJa5_1;
	wire w_dff_B_BznF3FIb6_1;
	wire w_dff_B_0X766xLg1_1;
	wire w_dff_B_Ohaxnjpv1_1;
	wire w_dff_B_Wv2zYr603_1;
	wire w_dff_B_qCibCRSU7_1;
	wire w_dff_B_esUgqMcf7_1;
	wire w_dff_B_g5YFE9H99_1;
	wire w_dff_B_QQv9vc7A3_1;
	wire w_dff_B_QcL6UJab8_1;
	wire w_dff_B_TSTDwVwp3_1;
	wire w_dff_B_Uf0UaQSc9_1;
	wire w_dff_B_xKDbCvj80_1;
	wire w_dff_B_a9NgOcio2_1;
	wire w_dff_B_HcrrAszy4_1;
	wire w_dff_B_BX3Q1osR8_1;
	wire w_dff_B_b7YPd1iR0_1;
	wire w_dff_B_mKgddXPJ7_1;
	wire w_dff_B_Ul9xBQiK3_1;
	wire w_dff_B_TpvobFwx6_1;
	wire w_dff_B_lpnll1dX3_1;
	wire w_dff_B_RYRal4Ol3_1;
	wire w_dff_B_hHpZTndD7_1;
	wire w_dff_B_3B7n4IN74_1;
	wire w_dff_B_x8QwSilg4_1;
	wire w_dff_B_apnd5IDr9_1;
	wire w_dff_B_IHiiTo3O6_1;
	wire w_dff_B_sIpOpXkx0_1;
	wire w_dff_B_s83mAJLg8_1;
	wire w_dff_B_yeVQDdmo1_1;
	wire w_dff_B_zfGdRU5l7_1;
	wire w_dff_B_67DesMrR9_1;
	wire w_dff_B_1Aoe1Zp02_1;
	wire w_dff_B_KJ8ERTgx0_1;
	wire w_dff_B_t6pgtpSN5_1;
	wire w_dff_B_0wvmjINJ5_1;
	wire w_dff_B_c1bT9x5k3_1;
	wire w_dff_B_4LN2QOOh6_1;
	wire w_dff_B_OfhxVnc54_1;
	wire w_dff_B_tiIEoovw4_1;
	wire w_dff_B_b53M9FKu8_1;
	wire w_dff_B_XxgO3fsy4_1;
	wire w_dff_B_Xlc5vSBR1_1;
	wire w_dff_B_aoAsfADC9_1;
	wire w_dff_B_2Mb77foR9_1;
	wire w_dff_B_5WwukQxC4_1;
	wire w_dff_B_RQ5xwhgu3_1;
	wire w_dff_B_bYMdPLlh5_1;
	wire w_dff_B_iwxCcSjO6_1;
	wire w_dff_B_fQfxNQOK0_1;
	wire w_dff_B_s8kfIGKo6_1;
	wire w_dff_B_tyYRCZIO8_1;
	wire w_dff_B_OEb6m1KX0_1;
	wire w_dff_B_Vo9cFIp64_1;
	wire w_dff_B_8y9R6sCY2_1;
	wire w_dff_B_tmAYfzY61_1;
	wire w_dff_B_LL1POgVB0_1;
	wire w_dff_B_1ywzHM0E6_1;
	wire w_dff_B_G2YRkX784_1;
	wire w_dff_B_euuIZCO06_1;
	wire w_dff_B_AOLl8XXU4_1;
	wire w_dff_B_3tJ6Ru2z1_1;
	wire w_dff_B_1xWW39aW4_1;
	wire w_dff_B_igPDpLnN4_1;
	wire w_dff_B_BQUck8pw6_1;
	wire w_dff_B_EMXdE2Dp7_1;
	wire w_dff_B_o5KyN9Av8_1;
	wire w_dff_B_iRKRjkPD3_1;
	wire w_dff_B_bNiXRNEt7_1;
	wire w_dff_B_VEZuYu6E5_1;
	wire w_dff_B_b0yhfW5y1_1;
	wire w_dff_B_XmdeWYy09_1;
	wire w_dff_B_RvcMJutV0_1;
	wire w_dff_B_q54efvMt6_1;
	wire w_dff_B_LZfvazFs7_1;
	wire w_dff_B_zkdoqCH55_1;
	wire w_dff_B_ldcZC9kl6_1;
	wire w_dff_B_zyZGnLg48_1;
	wire w_dff_B_6PCwuYHb9_1;
	wire w_dff_B_KO4JF4GX2_1;
	wire w_dff_B_xlK0L1Ug7_1;
	wire w_dff_B_wJjdlrfB6_1;
	wire w_dff_B_3Ji2gMQm7_1;
	wire w_dff_B_PfB9bUjh7_1;
	wire w_dff_B_dC8IHqIJ1_1;
	wire w_dff_B_HBS5AwK51_1;
	wire w_dff_B_EouPxaki8_1;
	wire w_dff_B_RrulAtdA1_1;
	wire w_dff_B_pF2aKIxn5_1;
	wire w_dff_B_MU30OuBi8_1;
	wire w_dff_B_2OfEKHBX4_1;
	wire w_dff_B_LS0Nnnbe9_1;
	wire w_dff_B_UI1ALbJ59_1;
	wire w_dff_B_i2YItJvF0_1;
	wire w_dff_B_u8OfvAuj2_1;
	wire w_dff_B_46lwCQV27_1;
	wire w_dff_B_ieZy9wnn7_1;
	wire w_dff_B_UM2IZ2TQ9_1;
	wire w_dff_B_G7fpRx6n5_1;
	wire w_dff_B_lWOX5vnu7_1;
	wire w_dff_B_w8mdgQxL8_1;
	wire w_dff_B_g0rjQRyU7_1;
	wire w_dff_B_mSkAwcO57_1;
	wire w_dff_B_8aKZDA7T4_1;
	wire w_dff_B_qiYe6hHG4_1;
	wire w_dff_B_p2oC7vdN4_1;
	wire w_dff_B_JbZNPpgs7_1;
	wire w_dff_B_HaaH6aMG8_1;
	wire w_dff_B_J7folQdM4_1;
	wire w_dff_B_yizmqqar9_1;
	wire w_dff_B_35aKkuzV0_1;
	wire w_dff_B_EHn5wVSy5_1;
	wire w_dff_B_JFgDmkrW3_1;
	wire w_dff_B_uXi9tDhs3_1;
	wire w_dff_B_vdqwhCzo3_1;
	wire w_dff_B_FqzXHXep2_1;
	wire w_dff_B_5UKeuiYK9_1;
	wire w_dff_B_qvxQFtuE9_1;
	wire w_dff_B_bXpVsNP53_1;
	wire w_dff_B_0fmmWaq16_1;
	wire w_dff_B_OeStJnji3_1;
	wire w_dff_B_LDuQEcWd1_1;
	wire w_dff_B_xifPqPjM2_1;
	wire w_dff_B_tXSItKuV4_1;
	wire w_dff_B_i0Qc3n010_1;
	wire w_dff_B_4Qc3BT602_1;
	wire w_dff_B_oKhZ9Px72_1;
	wire w_dff_B_r7Cgy82A9_1;
	wire w_dff_B_azoRYASO7_1;
	wire w_dff_B_5LPQTviR3_1;
	wire w_dff_B_oalh4PKc8_1;
	wire w_dff_B_VSJ31bKI6_1;
	wire w_dff_B_ERF1bee34_1;
	wire w_dff_B_GjShUze15_1;
	wire w_dff_B_xBN9sYd73_1;
	wire w_dff_B_TrtEvN463_1;
	wire w_dff_B_Dto28vYA0_1;
	wire w_dff_B_Wd6tI4do1_1;
	wire w_dff_B_nrI87EEZ2_1;
	wire w_dff_B_WuR5d0mp4_1;
	wire w_dff_B_R5ONn5iw7_1;
	wire w_dff_B_PP0smkJr0_1;
	wire w_dff_B_Z6uSNpOy7_1;
	wire w_dff_B_FkH7Nsub6_1;
	wire w_dff_B_bMddaBju1_1;
	wire w_dff_B_aNQnMqfL8_1;
	wire w_dff_B_cfoY5vZH4_1;
	wire w_dff_B_D1TEAkdy4_1;
	wire w_dff_B_nYixf4ck7_1;
	wire w_dff_B_E7GihjsA6_1;
	wire w_dff_B_OsmL041d6_1;
	wire w_dff_B_H0AYqXlV5_1;
	wire w_dff_B_AqCS8Wmr0_1;
	wire w_dff_B_5E5N8fbG7_1;
	wire w_dff_B_mbyGOUyK7_1;
	wire w_dff_B_NE2Esbso4_1;
	wire w_dff_B_hKZQVC1B9_1;
	wire w_dff_B_OaZI88vZ2_1;
	wire w_dff_B_QS0AaBq25_1;
	wire w_dff_B_nR662HS23_1;
	wire w_dff_B_fCejSuMv7_1;
	wire w_dff_B_fAWzTRaQ1_1;
	wire w_dff_B_yOrbzuPC5_1;
	wire w_dff_B_pzsHEBWb6_1;
	wire w_dff_B_Zn469Bwc7_1;
	wire w_dff_B_VLtRZy4v3_1;
	wire w_dff_B_ptQ25fex8_1;
	wire w_dff_B_jVX8F6Xl3_1;
	wire w_dff_B_CawEFLW32_1;
	wire w_dff_B_6Uk0kY1J5_1;
	wire w_dff_B_bbrhRmbf2_1;
	wire w_dff_B_Z3OEavTf6_1;
	wire w_dff_B_igpowbij3_1;
	wire w_dff_B_olWfDcaN6_1;
	wire w_dff_B_YXhLdMks0_1;
	wire w_dff_B_NQAj0qbZ9_1;
	wire w_dff_B_ngqDtuqD7_1;
	wire w_dff_B_kNPbp8J69_1;
	wire w_dff_B_8VV8Qc1M7_1;
	wire w_dff_B_ttafBy0w3_1;
	wire w_dff_B_bHVB0p1Z3_1;
	wire w_dff_B_AiGyld9I4_1;
	wire w_dff_B_6y3Mt8UG5_1;
	wire w_dff_B_z8w0zcKB8_0;
	wire w_dff_B_hV2wI3hE3_1;
	wire w_dff_B_tPuf6rMo7_1;
	wire w_dff_B_NK12tZbp3_1;
	wire w_dff_B_SKk71p9z7_1;
	wire w_dff_B_GiwqYT4t5_1;
	wire w_dff_B_gzxu1Q299_1;
	wire w_dff_B_7eVcSRTQ8_1;
	wire w_dff_B_DQvoTz455_1;
	wire w_dff_B_6cc3BkZ72_1;
	wire w_dff_B_IkXUt7xC5_1;
	wire w_dff_B_B10s512I5_1;
	wire w_dff_B_US89lrvl8_1;
	wire w_dff_B_hSmZqu2u0_1;
	wire w_dff_B_bJ7asy1c2_1;
	wire w_dff_B_huyM6Sbm7_1;
	wire w_dff_B_Zzjqdy094_0;
	wire w_dff_B_Lx8y4Qgd1_0;
	wire w_dff_B_n1DYH6Eu0_0;
	wire w_dff_B_BbkwgzEX7_0;
	wire w_dff_B_AnWxIQvn7_0;
	wire w_dff_B_Cu2zUTVv4_0;
	wire w_dff_B_fCzsxwc23_0;
	wire w_dff_B_hC0stYPe2_0;
	wire w_dff_B_xDjbwjZR5_0;
	wire w_dff_B_22CDTs6g3_0;
	wire w_dff_B_y0h7Pa8r2_0;
	wire w_dff_B_nUH4L31U6_0;
	wire w_dff_B_sQArDvcX8_0;
	wire w_dff_A_zNSE46Vu5_0;
	wire w_dff_A_V2Fsx7BU9_0;
	wire w_dff_A_bvULOijl7_0;
	wire w_dff_A_YY2plMGm3_0;
	wire w_dff_A_ccwjmVMm4_0;
	wire w_dff_A_AmWwTINm2_0;
	wire w_dff_A_jj2KitXd6_0;
	wire w_dff_A_0QE3QVJE9_0;
	wire w_dff_A_rZ7ONRVB7_0;
	wire w_dff_A_WEIV3QYS9_0;
	wire w_dff_A_rErx2SLH9_0;
	wire w_dff_A_gxGqzSXs2_0;
	wire w_dff_A_pgjsqp0w8_0;
	wire w_dff_A_L8ueDPvO2_0;
	wire w_dff_B_CwRSeIak2_1;
	wire w_dff_B_JdEVAEq01_1;
	wire w_dff_B_9c9ST8518_2;
	wire w_dff_B_MdcDDMGE5_2;
	wire w_dff_B_oGKanOkl0_2;
	wire w_dff_B_NgeIEH9P2_2;
	wire w_dff_B_DzNTginG5_2;
	wire w_dff_B_eKoW9Bcr7_2;
	wire w_dff_B_xKfx4z0l9_2;
	wire w_dff_B_47pJCbFJ9_2;
	wire w_dff_B_md9S7CLo4_2;
	wire w_dff_B_Wug8SRLh9_2;
	wire w_dff_B_c5thFNV69_2;
	wire w_dff_B_avL0NWVT2_2;
	wire w_dff_B_yldM4uHr4_2;
	wire w_dff_B_yyCtVycQ4_2;
	wire w_dff_B_Fb5PdAwy2_2;
	wire w_dff_B_4XwPFce52_2;
	wire w_dff_B_SPLC5CPS6_2;
	wire w_dff_B_HaKW4JTM6_2;
	wire w_dff_B_88C9hQyN6_2;
	wire w_dff_B_gda2oCd96_2;
	wire w_dff_B_QoPMMl6n7_2;
	wire w_dff_B_1DjAqkbo8_2;
	wire w_dff_B_EaUyJfyk4_2;
	wire w_dff_B_4p0V0LEh8_2;
	wire w_dff_B_GwtcKxKR3_2;
	wire w_dff_B_8dBBk3Rk7_2;
	wire w_dff_B_PMIi69VZ4_2;
	wire w_dff_B_GMkvc1yV0_2;
	wire w_dff_B_jO2yocm39_2;
	wire w_dff_B_Tv2aRw1p4_2;
	wire w_dff_B_6g1LHoz31_2;
	wire w_dff_B_dEqZoGSd7_2;
	wire w_dff_B_hQI3iIFS4_2;
	wire w_dff_B_WO3SNvig4_2;
	wire w_dff_B_p620AGEX3_2;
	wire w_dff_B_UDwP52Ud7_2;
	wire w_dff_B_wsO7XN0l8_2;
	wire w_dff_B_TSTtLijB6_2;
	wire w_dff_B_ijDm1qaW2_2;
	wire w_dff_B_0EXD4U4H2_2;
	wire w_dff_B_ia58TNRU7_2;
	wire w_dff_B_xNE0itga9_2;
	wire w_dff_B_KIGMbyhU2_2;
	wire w_dff_B_TrggROkz2_2;
	wire w_dff_B_mPZEw0Sx3_2;
	wire w_dff_B_2wUTUvBm1_2;
	wire w_dff_B_Zbsd94kw5_2;
	wire w_dff_B_qUOymOHe4_2;
	wire w_dff_B_bPgX9GmS9_2;
	wire w_dff_B_9eiVS16e5_2;
	wire w_dff_B_gdKuuyar9_2;
	wire w_dff_B_iT1HOUD15_2;
	wire w_dff_B_pls9ok3V1_2;
	wire w_dff_B_Ao8U18wJ8_2;
	wire w_dff_B_vA60CrKa1_2;
	wire w_dff_B_ulT9deez7_2;
	wire w_dff_B_TnNJYkFP3_2;
	wire w_dff_B_7cLve7654_1;
	wire w_dff_B_B7AqmFwC0_1;
	wire w_dff_B_ZBDtyjBf7_1;
	wire w_dff_B_nfKhVY6U7_1;
	wire w_dff_B_s2zwTIMK9_1;
	wire w_dff_B_fH90MPwb5_1;
	wire w_dff_B_yYdbQXdC5_1;
	wire w_dff_B_kcXlAPcu8_1;
	wire w_dff_B_hl3AyHsE8_1;
	wire w_dff_B_lViDSS2w3_1;
	wire w_dff_B_TIDP2gBH7_1;
	wire w_dff_B_Jif6Ryib0_1;
	wire w_dff_B_rKvz3qNj9_1;
	wire w_dff_B_NTsVBm794_0;
	wire w_dff_B_X3m0Mhqr1_0;
	wire w_dff_B_JJsjNdCn2_0;
	wire w_dff_B_xpjB9u8B6_0;
	wire w_dff_B_fMFD8vZA7_0;
	wire w_dff_B_XbszIEMB1_0;
	wire w_dff_B_pdpPE8Ce2_0;
	wire w_dff_B_uFpunoN25_0;
	wire w_dff_B_Bz1ltoA82_0;
	wire w_dff_B_1vNNiMQ23_0;
	wire w_dff_B_oT7xWidf7_0;
	wire w_dff_B_uG0G052K0_0;
	wire w_dff_A_WPGvsqm03_1;
	wire w_dff_A_hETNtujh0_1;
	wire w_dff_A_78BxAME50_1;
	wire w_dff_A_KFoJGfPx5_1;
	wire w_dff_A_TzyQriov7_1;
	wire w_dff_A_SczVSiE31_1;
	wire w_dff_A_DqlTu6MF6_1;
	wire w_dff_A_MSz7eijY0_1;
	wire w_dff_A_yQFGxJ9h3_1;
	wire w_dff_A_Mgt8YJNu3_1;
	wire w_dff_A_hP7rHZ7F3_1;
	wire w_dff_A_rstKqXmV5_1;
	wire w_dff_A_bKLg2vTL0_1;
	wire w_dff_B_YmazJ7807_1;
	wire w_dff_B_bGUZDYX04_1;
	wire w_dff_B_LjhZY2LC8_1;
	wire w_dff_B_LrYV5Ntu7_1;
	wire w_dff_B_oawRA7Kw5_1;
	wire w_dff_B_8vfzK27C1_1;
	wire w_dff_B_aKUpKm3y4_1;
	wire w_dff_B_RFLUSRNx9_1;
	wire w_dff_B_iDbRK6Ty8_1;
	wire w_dff_B_ix4VJOmh3_1;
	wire w_dff_B_JpgOkr6L9_1;
	wire w_dff_B_mwwiw5lE1_1;
	wire w_dff_B_yRWuqKkw5_1;
	wire w_dff_B_GnbcdT6s3_0;
	wire w_dff_B_PQTROi1O5_0;
	wire w_dff_B_fXrwwZH15_0;
	wire w_dff_B_2Mux3wgO2_0;
	wire w_dff_B_pwpySj0Q4_0;
	wire w_dff_B_Ys9Lr5Gk2_0;
	wire w_dff_B_YKptjCab5_0;
	wire w_dff_B_8sy3xX1L0_0;
	wire w_dff_B_7XPHU3ij2_0;
	wire w_dff_B_6MQAk3Jk8_0;
	wire w_dff_B_Ue28N7Wt2_0;
	wire w_dff_B_ZeYPt54T0_0;
	wire w_dff_A_DRe20etP5_1;
	wire w_dff_A_Payo0NRM4_1;
	wire w_dff_A_NCnB7HKx1_1;
	wire w_dff_A_xtky17vQ9_1;
	wire w_dff_A_76v08Zms2_1;
	wire w_dff_A_GHVd2Zyw9_1;
	wire w_dff_A_J7RdBkdz0_1;
	wire w_dff_A_r3anLi1b9_1;
	wire w_dff_A_1l4xKHte9_1;
	wire w_dff_A_BzNfuLlh3_1;
	wire w_dff_A_9SNYp1wM0_1;
	wire w_dff_A_Rjsuyn4I3_1;
	wire w_dff_A_7qFQCJai5_1;
	wire w_dff_B_eNlUkgVG5_1;
	wire w_dff_B_YWAHMO8q9_1;
	wire w_dff_B_dtiGdofG0_1;
	wire w_dff_B_4duU7BmE7_1;
	wire w_dff_B_Z8govWyO5_1;
	wire w_dff_B_HzdqHQ8b1_1;
	wire w_dff_B_49hZUSiv5_1;
	wire w_dff_B_yBNeNkrt9_1;
	wire w_dff_B_NV8Mmotu3_1;
	wire w_dff_B_UfNvOxqL0_1;
	wire w_dff_B_DuRBjKw84_1;
	wire w_dff_B_JQXNLPIO4_1;
	wire w_dff_B_7RvKsDtP2_1;
	wire w_dff_B_amPhIF7z0_0;
	wire w_dff_B_0jufnKom3_0;
	wire w_dff_B_FhmQjCn73_0;
	wire w_dff_B_HT2msORh7_0;
	wire w_dff_B_RkqyehRP2_0;
	wire w_dff_B_NSVuilWk4_0;
	wire w_dff_B_RNWkcmDE6_0;
	wire w_dff_B_mRCXoC721_0;
	wire w_dff_B_P1j5d9o49_0;
	wire w_dff_B_gmYC9GAI3_0;
	wire w_dff_B_DpBUIqX74_0;
	wire w_dff_B_uwUQSseo9_0;
	wire w_dff_A_tVT1kRa81_1;
	wire w_dff_A_m27y9gzO1_1;
	wire w_dff_A_xd4Zz27l4_1;
	wire w_dff_A_Kc73B2Dy1_1;
	wire w_dff_A_Imk16Ha12_1;
	wire w_dff_A_rcnkaNm23_1;
	wire w_dff_A_iChtqyvu4_1;
	wire w_dff_A_ThzbdRSI1_1;
	wire w_dff_A_jm8Lkqrz0_1;
	wire w_dff_A_e6Ndbnko0_1;
	wire w_dff_A_kMsrLRUe9_1;
	wire w_dff_A_oPgmPD5s8_1;
	wire w_dff_A_RXQQeR0j4_1;
	wire w_dff_B_Nxv2lKfY3_1;
	wire w_dff_B_Svgiq7dL8_1;
	wire w_dff_B_90TNmHwt5_1;
	wire w_dff_B_FrOJXGS59_1;
	wire w_dff_B_sxy5MF9o5_1;
	wire w_dff_B_Nq6ZbYhD8_1;
	wire w_dff_B_hj7KsYkM8_1;
	wire w_dff_B_EuXoRDHk3_1;
	wire w_dff_B_SD6C0Zyb9_1;
	wire w_dff_B_N8NeO2o61_1;
	wire w_dff_B_GRBTspeu4_1;
	wire w_dff_B_mLqofTnu3_1;
	wire w_dff_B_gEpp6YSE9_1;
	wire w_dff_B_5xmx5qGV8_0;
	wire w_dff_B_eLSVE3a04_0;
	wire w_dff_B_gncrlQUf1_0;
	wire w_dff_B_uOqhqrZZ5_0;
	wire w_dff_B_Uh3br8OP1_0;
	wire w_dff_B_sNHTtnzO9_0;
	wire w_dff_B_BzJNnD1D7_0;
	wire w_dff_B_BH4Of6eP9_0;
	wire w_dff_B_aVgAbiVL2_0;
	wire w_dff_B_A9IBnHUG1_0;
	wire w_dff_B_CZSJDSlp4_0;
	wire w_dff_B_CZ6KcnlD1_0;
	wire w_dff_A_Xqu6oyos0_1;
	wire w_dff_A_FZsRS98w9_1;
	wire w_dff_A_c2ocHHsM0_1;
	wire w_dff_A_4hJbz2qi8_1;
	wire w_dff_A_UMsmR2nH5_1;
	wire w_dff_A_XA7goTYL7_1;
	wire w_dff_A_zak9b8nx1_1;
	wire w_dff_A_6AwDm7zx1_1;
	wire w_dff_A_ZVsb9R9N5_1;
	wire w_dff_A_3MqrD0346_1;
	wire w_dff_A_y6QKNNti8_1;
	wire w_dff_A_9f82srkK4_1;
	wire w_dff_A_5HE7nm6i7_1;
	wire w_dff_B_NiDVM0IL5_1;
	wire w_dff_B_THVXFYeH5_1;
	wire w_dff_B_7I4s2tqs1_1;
	wire w_dff_B_RMbF241J6_1;
	wire w_dff_B_BmFgoTeU9_1;
	wire w_dff_B_DTPtxRqV5_1;
	wire w_dff_B_U4l6Lo1O8_1;
	wire w_dff_B_opdsPIUC0_1;
	wire w_dff_B_R2IaWWdf9_1;
	wire w_dff_B_CfiCXOBP8_1;
	wire w_dff_B_d17h1mHL1_1;
	wire w_dff_B_mKcOYGMj2_1;
	wire w_dff_B_BJyvovda8_1;
	wire w_dff_B_PHS5PLeG6_0;
	wire w_dff_B_JIpurjGO8_0;
	wire w_dff_B_sG6rwZFY1_0;
	wire w_dff_B_oBhBHtF84_0;
	wire w_dff_B_OdtYtcLg4_0;
	wire w_dff_B_xsNTFTtr1_0;
	wire w_dff_B_WNGqTnbW3_0;
	wire w_dff_B_FKsoa0ir1_0;
	wire w_dff_B_RQHNHvPB1_0;
	wire w_dff_B_hxzfebwW3_0;
	wire w_dff_B_OfOjkk3r2_0;
	wire w_dff_A_vpGPPpDK3_1;
	wire w_dff_A_pSKzezHl3_1;
	wire w_dff_A_Rusjejt27_1;
	wire w_dff_A_M9euufRg3_1;
	wire w_dff_A_eRHyMjoD2_1;
	wire w_dff_A_PVXk5nwi7_1;
	wire w_dff_A_MfpC0Ifo4_1;
	wire w_dff_A_hMwGH2CM1_1;
	wire w_dff_A_Ybb0AtZm0_1;
	wire w_dff_A_aXTdrMCm9_1;
	wire w_dff_A_S3s5DZjn4_1;
	wire w_dff_A_tcFSoMZz5_1;
	wire w_dff_B_e3ghwwLt7_1;
	wire w_dff_B_L9j5KGTg7_1;
	wire w_dff_B_2GY2a0XT6_1;
	wire w_dff_B_HVPxgTXN8_1;
	wire w_dff_B_mJSyy9Rn2_1;
	wire w_dff_B_Aigm1sfF2_1;
	wire w_dff_B_s606KOLh5_1;
	wire w_dff_B_OF9NdZiU4_1;
	wire w_dff_B_xoSSOig16_1;
	wire w_dff_B_m1bmlMH42_1;
	wire w_dff_B_s8cq0cag8_1;
	wire w_dff_B_Dr5rfgtG5_1;
	wire w_dff_B_D1a7pTL46_0;
	wire w_dff_B_OyFgyPyf2_0;
	wire w_dff_B_3Ws6aF4L7_0;
	wire w_dff_B_ymzlpt8I1_0;
	wire w_dff_B_OnHE1AtY9_0;
	wire w_dff_B_1oA95bXm2_0;
	wire w_dff_B_dgtYZbqV3_0;
	wire w_dff_B_Jo74UEam3_0;
	wire w_dff_B_0nBRYLJG4_0;
	wire w_dff_B_Dmfo7PaF5_0;
	wire w_dff_A_4gYtos4m5_1;
	wire w_dff_A_FV8rHZS99_1;
	wire w_dff_A_ydxLPViJ9_1;
	wire w_dff_A_dhhiH5bd2_1;
	wire w_dff_A_Vcc0JimF0_1;
	wire w_dff_A_V8eDVjaH6_1;
	wire w_dff_A_GwGo1QBI6_1;
	wire w_dff_A_njHiTBld0_1;
	wire w_dff_A_S8IsL0Ib0_1;
	wire w_dff_A_DhK7EMWn8_1;
	wire w_dff_A_0iecNvAh2_1;
	wire w_dff_B_LJJlWnk41_1;
	wire w_dff_B_3piuALWv7_1;
	wire w_dff_B_oTDNCRoU0_1;
	wire w_dff_B_9Cz1FamL9_1;
	wire w_dff_B_Ag025cPL1_1;
	wire w_dff_B_lk0hO8Yq2_1;
	wire w_dff_B_Z6oXm97H1_1;
	wire w_dff_B_WQEF9ekj2_1;
	wire w_dff_B_hmfNt6b79_1;
	wire w_dff_B_fPT3ph2e2_1;
	wire w_dff_B_lxy4xvBU3_0;
	wire w_dff_B_zpgqweIC2_0;
	wire w_dff_B_PrMF6BJ27_0;
	wire w_dff_B_dNHn36ia0_0;
	wire w_dff_B_dMpuQB7g0_0;
	wire w_dff_B_vyKnG3id5_0;
	wire w_dff_B_FU2qZ6LP7_0;
	wire w_dff_B_7MkU68A62_0;
	wire w_dff_A_MRcvc1uA4_1;
	wire w_dff_A_yu7UUQFT7_1;
	wire w_dff_A_OthvHi1X1_1;
	wire w_dff_A_bF84zSeK2_1;
	wire w_dff_A_ENBa59xu0_1;
	wire w_dff_A_1h5GEteT0_1;
	wire w_dff_A_Usz5I9JG5_1;
	wire w_dff_A_2sHKpfZJ6_1;
	wire w_dff_A_xuraak5w1_1;
	wire w_dff_B_ufxgNgqS8_1;
	wire w_dff_B_ztb9utD51_1;
	wire w_dff_B_kKiGYkkF8_1;
	wire w_dff_B_FLJ4YpMp7_1;
	wire w_dff_B_sDoBt1Vb4_1;
	wire w_dff_B_pgsVoisl2_1;
	wire w_dff_B_wJdjq6UD9_1;
	wire w_dff_B_la4C7ecR3_1;
	wire w_dff_B_dWAYz2Rc7_0;
	wire w_dff_B_1epMpAng0_0;
	wire w_dff_B_Bz65Kcuo5_0;
	wire w_dff_B_98FrXcK27_0;
	wire w_dff_B_5zVSnA2z6_0;
	wire w_dff_B_NW2B2g9Z9_0;
	wire w_dff_A_XFDpb1RG5_1;
	wire w_dff_A_3JmpqIru4_1;
	wire w_dff_A_xbN7cE4m9_1;
	wire w_dff_A_AGCUTb3e5_1;
	wire w_dff_A_o1mjaOtS0_1;
	wire w_dff_A_CzaZjN317_1;
	wire w_dff_A_G45fXfk25_1;
	wire w_dff_B_99jEtv879_1;
	wire w_dff_B_RwJTWK5E1_1;
	wire w_dff_B_D62o8hER1_1;
	wire w_dff_B_JohTtuWZ5_1;
	wire w_dff_B_zctOC7Yx2_1;
	wire w_dff_B_u2wEuWIl8_1;
	wire w_dff_B_6M8TUMrb7_1;
	wire w_dff_B_uzcjNXjC1_0;
	wire w_dff_B_zq4uOzPE2_0;
	wire w_dff_B_7hI0vCHj9_0;
	wire w_dff_B_HrYEjpWa5_0;
	wire w_dff_B_HRfc0iEy8_0;
	wire w_dff_A_Lrjqb8Q71_1;
	wire w_dff_A_ggzCto9m0_1;
	wire w_dff_A_VVPVeflc3_1;
	wire w_dff_A_6UoLyPy62_1;
	wire w_dff_A_ajr6RC2b0_1;
	wire w_dff_A_vTJCgUqr5_1;
	wire w_dff_B_DtWOtbt48_1;
	wire w_dff_B_x6YGrWCP2_1;
	wire w_dff_B_cgKo1uKb5_1;
	wire w_dff_B_sNmOolNm6_1;
	wire w_dff_B_Ly4X3evK3_1;
	wire w_dff_B_5Qqva24S8_1;
	wire w_dff_B_0BX5uYEF9_0;
	wire w_dff_B_b6oP3IBR6_0;
	wire w_dff_B_2pCn1TmJ8_0;
	wire w_dff_B_ZlZ6Nbus7_0;
	wire w_dff_A_4ONEt3wy6_1;
	wire w_dff_A_2j2h0TO31_1;
	wire w_dff_A_LPtiH6V44_1;
	wire w_dff_A_ytACUHtR0_1;
	wire w_dff_A_eCoR4Xyq0_1;
	wire w_dff_B_ciEhE5oa1_1;
	wire w_dff_B_CwNbjt9l7_1;
	wire w_dff_B_kUkGjYFU6_1;
	wire w_dff_A_LFIfuljK0_0;
	wire w_dff_A_HSElSoIF5_0;
	wire w_dff_B_4lbaaL8i8_1;
	wire w_dff_A_PYphhLrQ4_0;
	wire w_dff_B_RwNnqVnb6_1;
	wire w_dff_A_0ILHXRq21_1;
	wire w_dff_B_T4lBY7sl2_2;
	wire w_dff_B_4xi7J29C7_1;
	wire w_dff_A_7wZHuWQL2_0;
	wire w_dff_A_6cJ0fW5k2_0;
	wire w_dff_A_uhSwwA6H0_0;
	wire w_dff_A_f0TEMAuq8_0;
	wire w_dff_A_h7EAVs6D4_0;
	wire w_dff_A_rq093ssw9_0;
	wire w_dff_A_tdctkbOV7_0;
	wire w_dff_A_IRIJoYKg8_0;
	wire w_dff_A_x3REjARl0_0;
	wire w_dff_A_BnG97WkD2_0;
	wire w_dff_A_519OxtWA7_0;
	wire w_dff_A_GUR3HTEq2_0;
	wire w_dff_A_Ol7f7Yt26_0;
	wire w_dff_A_qEkqeOYb4_0;
	wire w_dff_A_p7tFtE577_0;
	wire w_dff_A_ZBV2MSCJ5_0;
	wire w_dff_A_Ye1uCfar5_0;
	wire w_dff_A_U3V8u78H4_0;
	wire w_dff_A_pvdl4QGc7_0;
	wire w_dff_A_hJ8zBZk38_0;
	wire w_dff_A_UAq6hRJH3_0;
	wire w_dff_A_NGo2YtPo8_0;
	wire w_dff_A_2sVv8gC40_0;
	wire w_dff_A_G5Ho0abw3_0;
	wire w_dff_A_zQaSjH4w4_0;
	wire w_dff_A_6vw6P3qt7_0;
	wire w_dff_A_fSUzXhIk9_0;
	wire w_dff_A_5ulZx8a16_0;
	wire w_dff_A_VItp2do45_0;
	wire w_dff_A_xLxnb5Pd4_0;
	wire w_dff_A_mADrcsg95_0;
	wire w_dff_A_gL54cPH75_0;
	wire w_dff_A_IORHVl6G9_0;
	wire w_dff_A_TyhxclkV9_0;
	wire w_dff_A_3vCRfo9D2_0;
	wire w_dff_A_DWvgFadZ6_0;
	wire w_dff_A_yC5md7O78_0;
	wire w_dff_A_Pamahlte9_0;
	wire w_dff_A_SlVhe1Ga5_0;
	wire w_dff_A_ozVsdxvV6_0;
	wire w_dff_A_2j9truBF6_0;
	wire w_dff_A_nCOFFhXa2_0;
	wire w_dff_A_fOMSH2Sk7_0;
	wire w_dff_A_ra8b89sL4_1;
	wire w_dff_B_fUgsaO6R2_1;
	wire w_dff_A_9MiIiI5w5_0;
	wire w_dff_A_waEKkhjf6_0;
	wire w_dff_A_69ytUQ3A2_0;
	wire w_dff_A_cricFCtc1_0;
	wire w_dff_A_FqntZ5Tl4_0;
	wire w_dff_A_BDf71oEe9_0;
	wire w_dff_A_VV4S4COs5_0;
	wire w_dff_A_iEuW9GLf4_0;
	wire w_dff_A_wGF92iH39_0;
	wire w_dff_A_0cM9jCbq7_0;
	wire w_dff_A_1RFis5Qd1_0;
	wire w_dff_A_M7FYKQnL0_0;
	wire w_dff_A_ZuQNXriM2_0;
	wire w_dff_A_A8vXEfk04_0;
	wire w_dff_A_fHoQzASn9_0;
	wire w_dff_A_q3L2bRJV4_0;
	wire w_dff_A_BHblP0pF8_0;
	wire w_dff_A_80Ax4HiU1_0;
	wire w_dff_A_a7bQXuza9_0;
	wire w_dff_A_d3Gl7lLy4_0;
	wire w_dff_A_meFxOqsl9_0;
	wire w_dff_A_S2lwdrPZ8_0;
	wire w_dff_A_y5gs4Hco1_0;
	wire w_dff_A_2QmPDKaM1_0;
	wire w_dff_A_82jbZI446_0;
	wire w_dff_A_rK3tfZIg7_0;
	wire w_dff_A_UAWSx7hy1_0;
	wire w_dff_A_Ko96IlfN0_0;
	wire w_dff_A_j9RYdZ2H2_0;
	wire w_dff_A_Q0cTpnbQ8_0;
	wire w_dff_A_wNsxdpsx3_0;
	wire w_dff_A_avqQY4bb2_0;
	wire w_dff_A_infK8D7j8_0;
	wire w_dff_A_pbCOyc8h0_0;
	wire w_dff_A_DtMsdpwU6_0;
	wire w_dff_A_A5FpTrrD7_0;
	wire w_dff_A_CVFsShbn7_0;
	wire w_dff_A_75sGKR2N7_0;
	wire w_dff_A_juJ0YWCi8_0;
	wire w_dff_A_Evzuf2IR8_0;
	wire w_dff_A_8ocpneNJ7_1;
	wire w_dff_B_f2s8ll5S7_1;
	wire w_dff_B_7zUKubWB6_1;
	wire w_dff_B_g3NAIaP19_1;
	wire w_dff_B_zKyZ22v46_1;
	wire w_dff_B_mpMOliPw9_1;
	wire w_dff_B_bcE9CSpy9_1;
	wire w_dff_B_dlzDynoQ1_1;
	wire w_dff_B_j0tIeTl78_1;
	wire w_dff_B_pLlDu1QI6_1;
	wire w_dff_B_IPAGpyNa0_1;
	wire w_dff_B_u30lyc8x6_1;
	wire w_dff_B_g9Bj4mR33_1;
	wire w_dff_B_nKzF8pWz9_1;
	wire w_dff_B_TEq6th2s5_1;
	wire w_dff_B_nKuV32Vx8_1;
	wire w_dff_B_h6kLfVcb0_1;
	wire w_dff_B_RiyIr1VH1_1;
	wire w_dff_B_Gympt39G8_1;
	wire w_dff_B_auS0WcJ65_1;
	wire w_dff_B_uHsCIQpA1_1;
	wire w_dff_B_pOAFj4aZ1_1;
	wire w_dff_B_aYxePEI51_1;
	wire w_dff_B_KW18rf0u3_1;
	wire w_dff_B_hygbpTQG2_1;
	wire w_dff_B_l2DXJUKw7_1;
	wire w_dff_B_bpVekJAE0_1;
	wire w_dff_B_P0Vt5Ayd2_1;
	wire w_dff_B_whaAqAAA6_1;
	wire w_dff_B_CGGRfG9D1_1;
	wire w_dff_B_jqOp89Qm7_1;
	wire w_dff_B_cPDyFdle6_1;
	wire w_dff_B_vWgwoJ0C9_1;
	wire w_dff_B_WcWjvEIU6_1;
	wire w_dff_B_gumcnGAx1_1;
	wire w_dff_B_nBj5gObl3_1;
	wire w_dff_B_BYWga9r30_1;
	wire w_dff_B_fCo7Mjhw4_1;
	wire w_dff_A_ZJqsWTE38_0;
	wire w_dff_A_DCweRg5G9_0;
	wire w_dff_A_hX73WQSW0_0;
	wire w_dff_A_USYjXc4M0_0;
	wire w_dff_A_ixLA7BGJ6_0;
	wire w_dff_A_wxoBXF8s7_0;
	wire w_dff_A_qEHhoYL80_0;
	wire w_dff_A_cX3KY70c8_0;
	wire w_dff_A_ijblW0et0_0;
	wire w_dff_A_O56tFSYs1_0;
	wire w_dff_A_0qlK8UcB2_0;
	wire w_dff_A_0ai6Xu861_0;
	wire w_dff_A_c7qtzy478_0;
	wire w_dff_A_WcqWStd04_0;
	wire w_dff_A_fdY2wFf83_0;
	wire w_dff_A_iYs6F8116_0;
	wire w_dff_A_T5gWcaLG1_0;
	wire w_dff_A_JudO6DsY1_0;
	wire w_dff_A_poqCqyYs2_0;
	wire w_dff_A_su1z9E7p4_0;
	wire w_dff_A_fSXXNJlq9_0;
	wire w_dff_A_wEsTfLSH6_0;
	wire w_dff_A_xCLZBxnn9_0;
	wire w_dff_A_ZGgbvMH67_0;
	wire w_dff_A_Sej4oIN88_0;
	wire w_dff_A_oyV8gBJ34_0;
	wire w_dff_A_l7rrKOUt6_0;
	wire w_dff_A_IM9QaROx9_0;
	wire w_dff_A_g2VpbbBh7_0;
	wire w_dff_A_cx1u4WQ89_0;
	wire w_dff_A_e7tTKAds4_0;
	wire w_dff_A_XqkBEqQ31_0;
	wire w_dff_A_PWjDeHci6_0;
	wire w_dff_A_dY0r4lcd6_0;
	wire w_dff_A_5BRhJD7N1_0;
	wire w_dff_A_vAxDeasC0_0;
	wire w_dff_A_QDiMJm2D6_0;
	wire w_dff_A_iUY45Q7M8_1;
	wire w_dff_B_A9VAm78q2_1;
	wire w_dff_B_LzmwLakx0_1;
	wire w_dff_B_ZSyUTwRc7_1;
	wire w_dff_B_42Ahjxve6_1;
	wire w_dff_B_WlzyMSi54_1;
	wire w_dff_B_2rCRDrJq6_1;
	wire w_dff_B_L977e37d9_1;
	wire w_dff_B_6CTHGhie9_1;
	wire w_dff_B_cZeONxXS9_1;
	wire w_dff_B_JNLUcxS15_1;
	wire w_dff_B_LogmgIUp3_1;
	wire w_dff_B_mgBfWcrG7_1;
	wire w_dff_B_EumMpXXp3_1;
	wire w_dff_B_7qv4UN6Y2_1;
	wire w_dff_B_gnVaiatE6_1;
	wire w_dff_B_mECXKtel3_1;
	wire w_dff_B_MIaqtrIC0_1;
	wire w_dff_B_3oUq2jOq1_1;
	wire w_dff_B_zgz4uphr2_1;
	wire w_dff_B_rd9DjhPC2_1;
	wire w_dff_B_7AHnIwJO3_1;
	wire w_dff_B_V2fvPVmd2_1;
	wire w_dff_B_vCZDwaJ74_1;
	wire w_dff_B_qLM4d4355_1;
	wire w_dff_B_DwxN9Yr58_1;
	wire w_dff_B_00rLh3e55_1;
	wire w_dff_B_fYR1K5me0_1;
	wire w_dff_B_KKRx64nL9_1;
	wire w_dff_B_eEHalRt61_1;
	wire w_dff_B_vuomH4Em3_1;
	wire w_dff_B_m0uvBwCu9_1;
	wire w_dff_B_SoQs1uK54_1;
	wire w_dff_B_0W0p7jUR3_1;
	wire w_dff_B_ZVITaAWb1_1;
	wire w_dff_A_nhDvlxFe4_0;
	wire w_dff_A_hEzlDyid1_0;
	wire w_dff_A_LMN6QWFi3_0;
	wire w_dff_A_zdwR896X3_0;
	wire w_dff_A_Cmglstuh2_0;
	wire w_dff_A_Nl0zI5LZ5_0;
	wire w_dff_A_RSNCOae38_0;
	wire w_dff_A_N1FfJhoA5_0;
	wire w_dff_A_HYh079cz5_0;
	wire w_dff_A_tZljyAks7_0;
	wire w_dff_A_8X8Jhouy3_0;
	wire w_dff_A_Gie4ZqOK9_0;
	wire w_dff_A_xgNC3I4N5_0;
	wire w_dff_A_iSccoqyV6_0;
	wire w_dff_A_boqlekLb4_0;
	wire w_dff_A_nOoTvesv8_0;
	wire w_dff_A_OuPDWl9o5_0;
	wire w_dff_A_IFEyOzj68_0;
	wire w_dff_A_hu77U5f90_0;
	wire w_dff_A_lIkyySYt0_0;
	wire w_dff_A_atsADPc67_0;
	wire w_dff_A_6ZuKJLlt6_0;
	wire w_dff_A_w7li6z5p6_0;
	wire w_dff_A_DmifbVad4_0;
	wire w_dff_A_PCxv85Wy7_0;
	wire w_dff_A_31BEGkBD1_0;
	wire w_dff_A_CFjU7RDm6_0;
	wire w_dff_A_2drIfCX83_0;
	wire w_dff_A_ek3ulER84_0;
	wire w_dff_A_IItxrOUx2_0;
	wire w_dff_A_AMAesH8T0_0;
	wire w_dff_A_vIpGoxcf1_0;
	wire w_dff_A_qHCW8PGe7_0;
	wire w_dff_A_bu9jZuxo2_0;
	wire w_dff_A_tWZbizCL0_1;
	wire w_dff_B_kCHBFrzY0_1;
	wire w_dff_B_Rd8TzzGj5_1;
	wire w_dff_B_tENXyBbO8_1;
	wire w_dff_B_g6xqOmz25_1;
	wire w_dff_B_hrUXolzj6_1;
	wire w_dff_B_ugocssaZ4_1;
	wire w_dff_B_CSr6RIpv1_1;
	wire w_dff_B_iBwWptcJ3_1;
	wire w_dff_B_Fj0Pwj9V7_1;
	wire w_dff_B_ER53Vsgq1_1;
	wire w_dff_B_uXHMzpMj3_1;
	wire w_dff_B_i2aGU7eZ7_1;
	wire w_dff_B_Ko8H580d3_1;
	wire w_dff_B_qqmrnoyj5_1;
	wire w_dff_B_M5TtD4UT8_1;
	wire w_dff_B_gEHEpSTY6_1;
	wire w_dff_B_p8LGoybh8_1;
	wire w_dff_B_V5hUxEtK1_1;
	wire w_dff_B_25lRxmGI1_1;
	wire w_dff_B_IyNrAS8v8_1;
	wire w_dff_B_y8CD5oan6_1;
	wire w_dff_B_748Wehi27_1;
	wire w_dff_B_kh3cpPPq2_1;
	wire w_dff_B_yOohTYGP9_1;
	wire w_dff_B_FEgnCTD95_1;
	wire w_dff_B_AnnayLHC9_1;
	wire w_dff_B_Uyh8CFlP1_1;
	wire w_dff_B_fq7cDSzQ7_1;
	wire w_dff_B_9mT4DgtD6_1;
	wire w_dff_B_vR0plZ4L4_1;
	wire w_dff_B_VXK70yMo3_1;
	wire w_dff_A_OTZF4ZFo9_0;
	wire w_dff_A_Cb8ck3cf5_0;
	wire w_dff_A_N3kcUESC7_0;
	wire w_dff_A_fBeDrGu99_0;
	wire w_dff_A_hHwR3u782_0;
	wire w_dff_A_AUvVvqXm5_0;
	wire w_dff_A_OSAg4mRU4_0;
	wire w_dff_A_hSXfgab13_0;
	wire w_dff_A_aVSZUbVy0_0;
	wire w_dff_A_tZZZ0Cgd1_0;
	wire w_dff_A_a4zs17Eo1_0;
	wire w_dff_A_GcPPHrYn8_0;
	wire w_dff_A_vJB0qnwq9_0;
	wire w_dff_A_pfhOpkfR0_0;
	wire w_dff_A_2QKP8nLj5_0;
	wire w_dff_A_lhi8bUCk6_0;
	wire w_dff_A_n9iK2LAY2_0;
	wire w_dff_A_pCPGAd0k0_0;
	wire w_dff_A_AdIacxm98_0;
	wire w_dff_A_wi5K90kP1_0;
	wire w_dff_A_OzyeiJQp1_0;
	wire w_dff_A_IzGg7SBo5_0;
	wire w_dff_A_1tXWoT3N0_0;
	wire w_dff_A_Yhmi73pX0_0;
	wire w_dff_A_HW5x8sja4_0;
	wire w_dff_A_JCaxpzaX2_0;
	wire w_dff_A_79MTMddy7_0;
	wire w_dff_A_bvmvRzxa6_0;
	wire w_dff_A_56tZM1Q22_0;
	wire w_dff_A_90ofgxfk4_0;
	wire w_dff_A_ERRIE9kX2_0;
	wire w_dff_A_kiwmOoXQ4_1;
	wire w_dff_B_zBMuKWgD3_1;
	wire w_dff_B_DnZAdYla3_1;
	wire w_dff_B_R4Ar9KN49_1;
	wire w_dff_B_KcFTeE4h5_1;
	wire w_dff_B_RXR5pRJ54_1;
	wire w_dff_B_G6ai8QNX2_1;
	wire w_dff_B_LTqYmLE73_1;
	wire w_dff_B_c7cHTrDQ1_1;
	wire w_dff_B_vwTbbMfu9_1;
	wire w_dff_B_qzxyu0aN4_1;
	wire w_dff_B_HIYPKxAn3_1;
	wire w_dff_B_jU9d4w7i2_1;
	wire w_dff_B_4z6oZ8he6_1;
	wire w_dff_B_XvF1Glm41_1;
	wire w_dff_B_zXNSOptH7_1;
	wire w_dff_B_otfm0FSw6_1;
	wire w_dff_B_8O76r0r17_1;
	wire w_dff_B_UUJVWsuS2_1;
	wire w_dff_B_FF4VzAs23_1;
	wire w_dff_B_WsWMziBW5_1;
	wire w_dff_B_Hwa1W5oB3_1;
	wire w_dff_B_uyrPcFlQ2_1;
	wire w_dff_B_ODTl2ZlX6_1;
	wire w_dff_B_Ak0VIRh19_1;
	wire w_dff_B_YezfJTEd4_1;
	wire w_dff_B_YrzUY8kt2_1;
	wire w_dff_B_YUvxqxm79_1;
	wire w_dff_B_LJWEIvt20_1;
	wire w_dff_A_xFbdq81z3_0;
	wire w_dff_A_FCQ7mtkf0_0;
	wire w_dff_A_FEfsb2Wf5_0;
	wire w_dff_A_Ri2JnhyP2_0;
	wire w_dff_A_RVueaT9M4_0;
	wire w_dff_A_6peDFwnx9_0;
	wire w_dff_A_4aofisUd7_0;
	wire w_dff_A_7GCzgXLn8_0;
	wire w_dff_A_SRM2ThGz5_0;
	wire w_dff_A_Gqg9NpGL7_0;
	wire w_dff_A_TpbmBRl95_0;
	wire w_dff_A_Nmm34HsN3_0;
	wire w_dff_A_qz0O7cJg1_0;
	wire w_dff_A_t4KNzypt8_0;
	wire w_dff_A_HYwUUR276_0;
	wire w_dff_A_UADPqvIj5_0;
	wire w_dff_A_RzRk2Cvz2_0;
	wire w_dff_A_TulId1XP1_0;
	wire w_dff_A_z1uLUdZy3_0;
	wire w_dff_A_kiJJroz33_0;
	wire w_dff_A_niUUt0470_0;
	wire w_dff_A_G00qHLd81_0;
	wire w_dff_A_X0F482pz5_0;
	wire w_dff_A_MCwLeiD24_0;
	wire w_dff_A_7H8fdpvx4_0;
	wire w_dff_A_QCgajTaP8_0;
	wire w_dff_A_Cffrl4qT1_0;
	wire w_dff_A_mhHgcLc15_0;
	wire w_dff_A_RSzIhc3H1_1;
	wire w_dff_B_8IzsM0oD3_1;
	wire w_dff_B_jL7slHTw7_1;
	wire w_dff_B_MxMOhbsl4_1;
	wire w_dff_B_kYRKIEJe8_1;
	wire w_dff_B_AzhsXSAm8_1;
	wire w_dff_B_l27U4c4U9_1;
	wire w_dff_B_Y2BR2rwX8_1;
	wire w_dff_B_dQ7RhL0j2_1;
	wire w_dff_B_M3EBURiR6_1;
	wire w_dff_B_wBDy8Uej1_1;
	wire w_dff_B_DVoJ7zCR3_1;
	wire w_dff_B_S9ZaIGoN3_1;
	wire w_dff_B_mc7YIRdA1_1;
	wire w_dff_B_ci266ybB5_1;
	wire w_dff_B_UWT8ro7g5_1;
	wire w_dff_B_QskdNfw20_1;
	wire w_dff_B_75B13Y7W2_1;
	wire w_dff_B_Ag1D4aU29_1;
	wire w_dff_B_15cdKQOx4_1;
	wire w_dff_B_5Sw6A1Cq3_1;
	wire w_dff_B_7SAOGW3R3_1;
	wire w_dff_B_vMg1hHGn4_1;
	wire w_dff_B_BGqwVxJj0_1;
	wire w_dff_B_o39bPTKi1_1;
	wire w_dff_B_qUFUEihJ6_1;
	wire w_dff_A_6OLEzaXf3_0;
	wire w_dff_A_eY119YXw3_0;
	wire w_dff_A_n9av7IQb4_0;
	wire w_dff_A_auMVzTH99_0;
	wire w_dff_A_XrQEAPYG6_0;
	wire w_dff_A_0nzDlDOa0_0;
	wire w_dff_A_eSBgJxCX8_0;
	wire w_dff_A_Ila1lE2m4_0;
	wire w_dff_A_WKUXKNJR6_0;
	wire w_dff_A_8xVbUGRS1_0;
	wire w_dff_A_MJZC7UVW9_0;
	wire w_dff_A_P7rHvVYo6_0;
	wire w_dff_A_c9UHDsyl7_0;
	wire w_dff_A_ERqEylzL4_0;
	wire w_dff_A_MJGTWWdj1_0;
	wire w_dff_A_U95dLSqh6_0;
	wire w_dff_A_G2zgbwfV5_0;
	wire w_dff_A_o2RSMPzA4_0;
	wire w_dff_A_RXOCSMT92_0;
	wire w_dff_A_WtEesyWf0_0;
	wire w_dff_A_vDLIzGEw7_0;
	wire w_dff_A_WCsDVMnX1_0;
	wire w_dff_A_6vSefmfV5_0;
	wire w_dff_A_7HWt21FX3_0;
	wire w_dff_A_k1BBpuyE8_0;
	wire w_dff_A_Bovu7nZx1_1;
	wire w_dff_B_e8GjJcCW9_1;
	wire w_dff_B_BuGj6LmC7_1;
	wire w_dff_B_RqGqG74g8_1;
	wire w_dff_B_WImsQgUi5_1;
	wire w_dff_B_vF7Lls0q3_1;
	wire w_dff_B_Gy6lrtYG3_1;
	wire w_dff_B_eKfU6hzp1_1;
	wire w_dff_B_yndFDEJi3_1;
	wire w_dff_B_sbJdPLQ23_1;
	wire w_dff_B_ibPIAYSx6_1;
	wire w_dff_B_feS9UsVx4_1;
	wire w_dff_B_FurDQtN38_1;
	wire w_dff_B_5HMl790y2_1;
	wire w_dff_B_jyvY51ll4_1;
	wire w_dff_B_td2FHD193_1;
	wire w_dff_B_KbefJUfY2_1;
	wire w_dff_B_eBGwZBbY3_1;
	wire w_dff_B_WzNbvo4m5_1;
	wire w_dff_B_1d3JgBps1_1;
	wire w_dff_B_oEH0J9py3_1;
	wire w_dff_B_Y7eTPMcT7_1;
	wire w_dff_B_P7NpbNA11_1;
	wire w_dff_A_D0Qidzpm9_0;
	wire w_dff_A_yMczb0lx9_0;
	wire w_dff_A_DMy0DIpY8_0;
	wire w_dff_A_oiy70Ye71_0;
	wire w_dff_A_V1h4Rjwg7_0;
	wire w_dff_A_CWeX05oF3_0;
	wire w_dff_A_5qC8yfzW7_0;
	wire w_dff_A_13OJlsHp3_0;
	wire w_dff_A_h5S33M530_0;
	wire w_dff_A_poXiEqOV4_0;
	wire w_dff_A_5kNhbh6y7_0;
	wire w_dff_A_e8JIFoMd9_0;
	wire w_dff_A_9EEJxgeo5_0;
	wire w_dff_A_ZOgyuoVn7_0;
	wire w_dff_A_Cf2f3QFx5_0;
	wire w_dff_A_zvRImTZy9_0;
	wire w_dff_A_D6LMTFrW8_0;
	wire w_dff_A_k7yBVQ1b5_0;
	wire w_dff_A_r7j8Heqh9_0;
	wire w_dff_A_Hn8yPNAj3_0;
	wire w_dff_A_HRlk4xJI7_0;
	wire w_dff_A_MScdtDYV3_0;
	wire w_dff_A_z1v3IO1U1_1;
	wire w_dff_B_OatZHRhl5_1;
	wire w_dff_B_E2m2I4tc4_1;
	wire w_dff_B_chenxPSq4_1;
	wire w_dff_B_J1Ave9H68_1;
	wire w_dff_B_AnLyatS00_1;
	wire w_dff_B_FhbxRMqo2_1;
	wire w_dff_B_Nns16vPM0_1;
	wire w_dff_B_XjGdVqET9_1;
	wire w_dff_B_GfNLBomx2_1;
	wire w_dff_B_EwLD71nM2_1;
	wire w_dff_B_zMiVHBW53_1;
	wire w_dff_B_6Z095BjI0_1;
	wire w_dff_B_DZPrepAl3_1;
	wire w_dff_B_xkW8tMkH8_1;
	wire w_dff_B_ZkP7TBDr9_1;
	wire w_dff_B_LQ6f3UFc1_1;
	wire w_dff_B_odZ837622_1;
	wire w_dff_B_vzXoSk9X4_1;
	wire w_dff_B_adsMT2n22_1;
	wire w_dff_A_k4xenT4h7_0;
	wire w_dff_A_a7we9Gva3_0;
	wire w_dff_A_I0ImGIF14_0;
	wire w_dff_A_13YisptX2_0;
	wire w_dff_A_I9Lt9Vzd6_0;
	wire w_dff_A_BTmGs1Yk9_0;
	wire w_dff_A_tPINrfYB9_0;
	wire w_dff_A_BPjLgJLX3_0;
	wire w_dff_A_ucfuI76z7_0;
	wire w_dff_A_dkBXmf8y8_0;
	wire w_dff_A_5HtJrMS99_0;
	wire w_dff_A_5zkDC9HT5_0;
	wire w_dff_A_YOSbSJAe4_0;
	wire w_dff_A_Aw2O2uyB6_0;
	wire w_dff_A_2eztFaSA8_0;
	wire w_dff_A_6D4g2EIK1_0;
	wire w_dff_A_wbKw1Hd12_0;
	wire w_dff_A_Z720XUCY7_0;
	wire w_dff_A_mzsbKJ0A0_0;
	wire w_dff_A_mMzflZNv3_1;
	wire w_dff_B_AdKknkAd7_1;
	wire w_dff_B_Ym6Vbl3d6_1;
	wire w_dff_B_ATfipyHE7_1;
	wire w_dff_B_psPElH7X9_1;
	wire w_dff_B_o9LOOIpQ2_1;
	wire w_dff_B_57Rkjt1g2_1;
	wire w_dff_B_oYqScWT52_1;
	wire w_dff_B_lV0f9tA09_1;
	wire w_dff_B_hVxklnD74_1;
	wire w_dff_B_5jGr5oyl7_1;
	wire w_dff_B_Dcg3VGSg8_1;
	wire w_dff_B_ptQJVMAC3_1;
	wire w_dff_B_b6MtkQpX9_1;
	wire w_dff_B_rKwLbcEY2_1;
	wire w_dff_B_aBcORKe87_1;
	wire w_dff_B_e2lxoe595_1;
	wire w_dff_A_0pDleJ5R5_0;
	wire w_dff_A_mHUCRWvC3_0;
	wire w_dff_A_KvTRu6M32_0;
	wire w_dff_A_NMlXlc5E6_0;
	wire w_dff_A_6Vq3yUtu1_0;
	wire w_dff_A_EnQjXoip4_0;
	wire w_dff_A_Lr4elQOt6_0;
	wire w_dff_A_8UBRyQ647_0;
	wire w_dff_A_JYv7GULW8_0;
	wire w_dff_A_GscKWzc12_0;
	wire w_dff_A_guE4PUy30_0;
	wire w_dff_A_Ju6eZYVy8_0;
	wire w_dff_A_R1jzM2gi9_0;
	wire w_dff_A_MElvZuSi2_0;
	wire w_dff_A_8MtG78A65_0;
	wire w_dff_A_O45etuQo1_0;
	wire w_dff_A_w1J36y282_1;
	wire w_dff_B_kMJdIi8X0_1;
	wire w_dff_B_acniKS1l7_1;
	wire w_dff_B_sKMPpX0Y6_1;
	wire w_dff_B_lkREedsx8_1;
	wire w_dff_B_LuK1vCnM8_1;
	wire w_dff_B_7iCANmHr3_1;
	wire w_dff_B_5R1v7BSg4_1;
	wire w_dff_B_lIklxeFu5_1;
	wire w_dff_B_EMIjIBl47_1;
	wire w_dff_B_pRj0KyJu7_1;
	wire w_dff_B_Zyuwm4wT3_1;
	wire w_dff_B_223yyBnc1_1;
	wire w_dff_B_mivY9yYO3_1;
	wire w_dff_A_YghuRqzn2_0;
	wire w_dff_A_mCe75unF2_0;
	wire w_dff_A_LLBwnret3_0;
	wire w_dff_A_A2uk5kT93_0;
	wire w_dff_A_GRq9yJjw4_0;
	wire w_dff_A_IbVR6JTN4_0;
	wire w_dff_A_Kcu7LNBs7_0;
	wire w_dff_A_rGT5YZ3j4_0;
	wire w_dff_A_ApxXQGR94_0;
	wire w_dff_A_V76GR7Iw8_0;
	wire w_dff_A_2TC2PRkm0_0;
	wire w_dff_A_ItZ3DfJD9_0;
	wire w_dff_A_vEHJDhK88_0;
	wire w_dff_A_RjMD47tF9_1;
	wire w_dff_B_uW5YyeLi5_1;
	wire w_dff_B_F8HT6iDB7_1;
	wire w_dff_B_spgkFarl1_1;
	wire w_dff_B_Cl3PKAn14_1;
	wire w_dff_B_H0hHKyTQ3_1;
	wire w_dff_B_3NaMh7mf2_1;
	wire w_dff_B_8u50gTNV8_1;
	wire w_dff_B_U8ykEoTV5_1;
	wire w_dff_B_kHBgj2ct0_1;
	wire w_dff_B_gf04LRoR5_1;
	wire w_dff_A_KFtXeObF6_0;
	wire w_dff_A_gDAG2uvu0_0;
	wire w_dff_A_l3fN9AQo9_0;
	wire w_dff_A_zmhu8g9k0_0;
	wire w_dff_A_DlyKsRMP4_0;
	wire w_dff_A_4nmWnb527_0;
	wire w_dff_A_valVlmqL2_0;
	wire w_dff_A_gF5BJC1H4_0;
	wire w_dff_A_CxuUWjyH7_0;
	wire w_dff_A_mRes1rl40_0;
	wire w_dff_A_WxYnSB6O0_1;
	wire w_dff_B_IuinFrhh4_1;
	wire w_dff_B_BQSZpY1a8_1;
	wire w_dff_B_PdmuyN320_1;
	wire w_dff_B_W36D3cMK6_1;
	wire w_dff_B_NGmeOSA00_1;
	wire w_dff_B_Su360Bny1_1;
	wire w_dff_B_wzAgij7Z4_1;
	wire w_dff_A_9U95j5xh3_0;
	wire w_dff_A_ZP3HyAxE7_0;
	wire w_dff_A_uiWKBazU3_0;
	wire w_dff_A_kFeW8RfP9_0;
	wire w_dff_A_KoVx2Kan5_0;
	wire w_dff_A_Ylz2tDqD9_0;
	wire w_dff_A_GHg8aXye0_0;
	wire w_dff_A_GQBtAAG96_1;
	wire w_dff_B_Uv9ReWOd9_1;
	wire w_dff_B_NMrMQwpv2_1;
	wire w_dff_B_cXBzVoJC3_1;
	wire w_dff_B_bRNIW5P95_1;
	wire w_dff_B_9Vf5Icva4_2;
	wire w_dff_A_CH6f1AEo0_0;
	wire w_dff_A_BfS0jTiv1_0;
	wire w_dff_A_HwO8AQJo2_0;
	wire w_dff_A_eQtCUR2S4_0;
	wire w_dff_B_QKLZD07U2_0;
	wire w_dff_A_HWHyE6Iw3_0;
	wire w_dff_A_eAFIM9nI2_0;
	wire w_dff_A_ezmFXke16_1;
	wire w_dff_B_ha1f2K3W5_1;
	wire w_dff_B_SVlH4JPV1_2;
	wire w_dff_B_1dCmcIVs7_2;
	wire w_dff_B_HXwN8Lw13_2;
	wire w_dff_B_z04SlnyX3_2;
	wire w_dff_B_Yq8ukHI04_2;
	wire w_dff_B_NmQc9hKf4_2;
	wire w_dff_B_XuNwJZp97_2;
	wire w_dff_B_fKhPNZ3o0_2;
	wire w_dff_B_13MhYITO2_2;
	wire w_dff_B_XFPRGYNU8_2;
	wire w_dff_B_buTV6WBg6_2;
	wire w_dff_B_UjuXZ5CJ3_2;
	wire w_dff_B_05ly3pzf6_2;
	wire w_dff_B_1BVgJJ1u8_2;
	wire w_dff_B_XLESq5Yo7_2;
	wire w_dff_B_bvomDQYL5_2;
	wire w_dff_B_q9w15ckF9_2;
	wire w_dff_B_hD4v8Ou89_2;
	wire w_dff_B_X7ecC6Wd5_2;
	wire w_dff_B_QafV0eiG5_2;
	wire w_dff_B_RrjQB6hy1_2;
	wire w_dff_B_NGJoTSCz3_2;
	wire w_dff_B_ayq64um91_2;
	wire w_dff_B_19hUALFP2_2;
	wire w_dff_B_MGeJWS6N6_2;
	wire w_dff_B_S4elgKpK0_2;
	wire w_dff_B_NUkd8ZMM3_2;
	wire w_dff_B_Pdm31MgI0_2;
	wire w_dff_B_ST9919Fo5_2;
	wire w_dff_B_rykJtCo34_2;
	wire w_dff_B_v9OHv9Jy7_2;
	wire w_dff_B_9UDA5jTH7_2;
	wire w_dff_B_o96nVqcz0_2;
	wire w_dff_B_dsntBdmM9_2;
	wire w_dff_B_PGcsK3oM3_2;
	wire w_dff_B_DW5CnjLJ6_2;
	wire w_dff_B_kPbPoVDA1_2;
	wire w_dff_B_U2tUafzD3_2;
	wire w_dff_B_eWjOhlCz6_2;
	wire w_dff_B_n3CbNZ7m1_2;
	wire w_dff_B_h19lBGnf6_2;
	wire w_dff_B_YmRQM7ho6_2;
	wire w_dff_B_5PjTactY9_2;
	wire w_dff_A_2JoOJDSK2_0;
	wire w_dff_B_dHhXXkpS5_1;
	wire w_dff_B_J4iVVmD45_2;
	wire w_dff_B_kRUpxviw3_2;
	wire w_dff_B_00tmrzpk5_2;
	wire w_dff_B_sX4AHlqn2_2;
	wire w_dff_B_XiFH1nWY4_2;
	wire w_dff_B_JjgOmFdZ7_2;
	wire w_dff_B_xCXM2NdE3_2;
	wire w_dff_B_tXtJZLsf3_2;
	wire w_dff_B_C68lsUKi6_2;
	wire w_dff_B_o8ytgLja9_2;
	wire w_dff_B_5maTWP3Q7_2;
	wire w_dff_B_EOLkSml62_2;
	wire w_dff_B_5J2p2Z6a5_2;
	wire w_dff_B_wiSXpisI5_2;
	wire w_dff_B_T20hXRdQ5_2;
	wire w_dff_B_hyFsdzvO5_2;
	wire w_dff_B_ZHpLUpvA3_2;
	wire w_dff_B_C6MODavM5_2;
	wire w_dff_B_Q4GKMZ6Q8_2;
	wire w_dff_B_yBBfHVMM8_2;
	wire w_dff_B_6rFDfqKX0_2;
	wire w_dff_B_rYoQMKwM4_2;
	wire w_dff_B_mC83W5Rc5_2;
	wire w_dff_B_uJtnMJem2_2;
	wire w_dff_B_QKsNVTjd3_2;
	wire w_dff_B_oqvn98nS2_2;
	wire w_dff_B_7BcMa4337_2;
	wire w_dff_B_8hs0nVhs3_2;
	wire w_dff_B_Vc8OozMm0_2;
	wire w_dff_B_PYBsMJ9P9_2;
	wire w_dff_B_xMXPbBb82_2;
	wire w_dff_B_p2nWBI8F7_2;
	wire w_dff_B_ddwJvNLP0_2;
	wire w_dff_B_KjfHu9ii9_2;
	wire w_dff_B_0AxgoCU34_2;
	wire w_dff_B_FGlZw0UB6_2;
	wire w_dff_B_apCgWL839_2;
	wire w_dff_B_AgWRX1l88_2;
	wire w_dff_B_WQwPjHer9_2;
	wire w_dff_B_hfAiVJWe3_2;
	wire w_dff_A_5cOfMQR71_1;
	wire w_dff_B_RNAk0Tkx4_1;
	wire w_dff_B_PhiVPLAi5_1;
	wire w_dff_B_InFZxYzN7_1;
	wire w_dff_B_oBaMsv0G5_1;
	wire w_dff_B_jMryvljm0_1;
	wire w_dff_B_jMceVpjg0_1;
	wire w_dff_B_heRGCE8B9_1;
	wire w_dff_B_GaBfpLVx4_1;
	wire w_dff_B_9uO6NMfn0_1;
	wire w_dff_B_x3ieAqcX2_1;
	wire w_dff_B_7IiFwS3P8_1;
	wire w_dff_B_MMbV8bfs2_1;
	wire w_dff_B_EwlDGIH42_1;
	wire w_dff_B_cdFzpImB1_1;
	wire w_dff_B_dl5NeYNR9_1;
	wire w_dff_B_5vqpXoGX5_1;
	wire w_dff_B_ZjGfVioi1_1;
	wire w_dff_B_0q1L5jKI0_1;
	wire w_dff_B_G80Po5kR9_1;
	wire w_dff_B_huyKn8U95_1;
	wire w_dff_B_VSsqfEtz9_1;
	wire w_dff_B_fHp5JBK31_1;
	wire w_dff_B_Y50gPpK19_1;
	wire w_dff_B_3ivmdiVg8_1;
	wire w_dff_B_iX1uKm0m5_1;
	wire w_dff_B_SyEwpmjE0_1;
	wire w_dff_B_lZFbIdAi7_1;
	wire w_dff_B_p6NBbtwH1_1;
	wire w_dff_B_yEzUR16l3_1;
	wire w_dff_B_BVIuilGA2_1;
	wire w_dff_B_9Dp1CswD9_1;
	wire w_dff_B_0UZTnRyO1_1;
	wire w_dff_B_mGM3q0Vz8_1;
	wire w_dff_B_KUOq6v4B6_1;
	wire w_dff_B_Ga6U3ZaT1_1;
	wire w_dff_B_i87Plare9_1;
	wire w_dff_B_Z8LzQloI7_1;
	wire w_dff_A_nvzMUPSq9_0;
	wire w_dff_A_mFVKxGu34_0;
	wire w_dff_A_irLXAV5G9_0;
	wire w_dff_A_RyDPdlYE3_0;
	wire w_dff_A_cE9ToscC4_0;
	wire w_dff_A_E4D3sfKA6_0;
	wire w_dff_A_Jk9NLDmv1_0;
	wire w_dff_A_MX7Ewhas0_0;
	wire w_dff_A_B8nYgEY25_0;
	wire w_dff_A_eZzfNJOH7_0;
	wire w_dff_A_UsNuXq1X7_0;
	wire w_dff_A_MXIAfFn31_0;
	wire w_dff_A_yO15gPJr5_0;
	wire w_dff_A_vP0gkV1y6_0;
	wire w_dff_A_kdFHnUVh3_0;
	wire w_dff_A_Lm5Gs0yh8_0;
	wire w_dff_A_TOM3HrQ90_0;
	wire w_dff_A_dViOtFSk2_0;
	wire w_dff_A_AZWB3P7r5_0;
	wire w_dff_A_60ukqH3e5_0;
	wire w_dff_A_k9uGuW0y1_0;
	wire w_dff_A_aJjaHec75_0;
	wire w_dff_A_DnOZtxGb6_0;
	wire w_dff_A_KYdOX3r87_0;
	wire w_dff_A_h8Kp11Vq8_0;
	wire w_dff_A_Bt6sxac45_0;
	wire w_dff_A_BPXW0qTw3_0;
	wire w_dff_A_t55fvk2X7_0;
	wire w_dff_A_MaHfv1FW1_0;
	wire w_dff_A_Y7GbduvZ9_0;
	wire w_dff_A_14xhSJk46_0;
	wire w_dff_A_ImEE9lU15_0;
	wire w_dff_A_iLKi4kvh6_0;
	wire w_dff_A_9KENl70F9_0;
	wire w_dff_A_4Rx08WPt0_0;
	wire w_dff_A_RF7ZFcvi5_0;
	wire w_dff_A_4Ww2YHwk1_0;
	wire w_dff_A_CozEEMQj4_0;
	wire w_dff_B_BOjcivN93_1;
	wire w_dff_A_BxerMc0E2_0;
	wire w_dff_A_cimKIYuX4_0;
	wire w_dff_A_WayADUjb1_0;
	wire w_dff_A_KuDZC9I02_0;
	wire w_dff_A_08M9oir51_0;
	wire w_dff_A_tL04Z9ZC3_0;
	wire w_dff_A_lQBRQG533_0;
	wire w_dff_A_yc2Ulbxy7_0;
	wire w_dff_A_WALWMKSr5_0;
	wire w_dff_A_kTz6nelh8_0;
	wire w_dff_A_CBnURHp55_0;
	wire w_dff_A_FbDy6Hqa8_0;
	wire w_dff_A_wE4lDe5G2_0;
	wire w_dff_A_6gPJGe730_0;
	wire w_dff_A_VhV8I7eJ5_0;
	wire w_dff_A_gzDa1RYH1_0;
	wire w_dff_A_nwetkaC47_0;
	wire w_dff_A_9EQNKs7y2_0;
	wire w_dff_A_0n1Cb1087_0;
	wire w_dff_A_0CZJAKpG5_0;
	wire w_dff_A_X2SkhwMt9_0;
	wire w_dff_A_F5OZ1ssi3_0;
	wire w_dff_A_f3oK9d4V5_0;
	wire w_dff_A_lOdRId168_0;
	wire w_dff_A_SyaBC5oX3_0;
	wire w_dff_A_PNUyjw2S6_0;
	wire w_dff_A_VHH0K7Fk1_0;
	wire w_dff_A_I0vO1TjO2_0;
	wire w_dff_A_QcxV2Gco2_0;
	wire w_dff_A_Uz29G7AQ7_0;
	wire w_dff_A_AALeN3uJ1_0;
	wire w_dff_A_VUxJTziZ8_0;
	wire w_dff_A_8AzY1BgI9_0;
	wire w_dff_A_z3WtrQqV4_0;
	wire w_dff_A_UaJP31Zr4_0;
	wire w_dff_B_L54OtKa01_1;
	wire w_dff_A_j5LpYyAI9_0;
	wire w_dff_A_4GuMcs7N8_0;
	wire w_dff_A_p0kP9c4r6_0;
	wire w_dff_A_za4cIv037_0;
	wire w_dff_A_wAJFscVw8_0;
	wire w_dff_A_b7g7ZcYN2_0;
	wire w_dff_A_z2ZGlGEA4_0;
	wire w_dff_A_umsH6zCL8_0;
	wire w_dff_A_JLlDFbRd2_0;
	wire w_dff_A_x5KzGJFz5_0;
	wire w_dff_A_NdGpRJNo7_0;
	wire w_dff_A_MvVhzOVP0_0;
	wire w_dff_A_mh6JhjAo7_0;
	wire w_dff_A_7hFL9iPU2_0;
	wire w_dff_A_zEVAQUr66_0;
	wire w_dff_A_SnifY13u4_0;
	wire w_dff_A_k3fn1NIj1_0;
	wire w_dff_A_6zqEzYZu6_0;
	wire w_dff_A_7XWCDsIC5_0;
	wire w_dff_A_fNutgw799_0;
	wire w_dff_A_rUtuXh2z2_0;
	wire w_dff_A_X6Mg3W7K6_0;
	wire w_dff_A_WuETERNJ9_0;
	wire w_dff_A_m8Rt0BIM9_0;
	wire w_dff_A_ZhwonHSi7_0;
	wire w_dff_A_CULjJBlH4_0;
	wire w_dff_A_TdxwIVvD1_0;
	wire w_dff_A_HfS7QI0y6_0;
	wire w_dff_A_bim36IMe0_0;
	wire w_dff_A_PDCWZ8WG3_0;
	wire w_dff_A_fuaXEbQU2_0;
	wire w_dff_A_tK0LOVYt9_0;
	wire w_dff_B_25LyZmhv8_1;
	wire w_dff_A_1DTD4n8o4_0;
	wire w_dff_A_27Vjn8E55_0;
	wire w_dff_A_BliCZHBw1_0;
	wire w_dff_A_fXjxcnL24_0;
	wire w_dff_A_HOjB8P6M0_0;
	wire w_dff_A_1EmnySFl3_0;
	wire w_dff_A_FuMXZAhx2_0;
	wire w_dff_A_UxwMdAWx5_0;
	wire w_dff_A_pWCk4pl57_0;
	wire w_dff_A_VAfjNRrt7_0;
	wire w_dff_A_fOvk9cU14_0;
	wire w_dff_A_wAk2BdGn2_0;
	wire w_dff_A_Zz4QNO8u9_0;
	wire w_dff_A_kqjg2sC43_0;
	wire w_dff_A_bHnznFdG8_0;
	wire w_dff_A_aVJMZtkD3_0;
	wire w_dff_A_TliCd5nd7_0;
	wire w_dff_A_vgzIR9E05_0;
	wire w_dff_A_86JmCiBZ5_0;
	wire w_dff_A_z9Z0vJC13_0;
	wire w_dff_A_bVLbzTMZ9_0;
	wire w_dff_A_OanEgcdL1_0;
	wire w_dff_A_ZQtBZvJU8_0;
	wire w_dff_A_qfSXjFBA6_0;
	wire w_dff_A_L6IHRjm13_0;
	wire w_dff_A_4Wo6oDnA2_0;
	wire w_dff_A_CqY9cvf81_0;
	wire w_dff_A_ufPHR4DL3_0;
	wire w_dff_A_ZUZuYvs31_0;
	wire w_dff_B_n8ulN2hL2_1;
	wire w_dff_A_xjivaEHV1_0;
	wire w_dff_A_ZvFdidse1_0;
	wire w_dff_A_xFCNRFwu0_0;
	wire w_dff_A_Kua27kwP5_0;
	wire w_dff_A_1FeNvmBt3_0;
	wire w_dff_A_IxzFZAqA6_0;
	wire w_dff_A_2qGJEOFE4_0;
	wire w_dff_A_kaogT0kH7_0;
	wire w_dff_A_bKpgsxEn1_0;
	wire w_dff_A_NZwXKZmx8_0;
	wire w_dff_A_KHPVtjxh0_0;
	wire w_dff_A_xrEJUqYf1_0;
	wire w_dff_A_jY8NaeET5_0;
	wire w_dff_A_POqxp1OC9_0;
	wire w_dff_A_cgWZzR0d5_0;
	wire w_dff_A_e5NLw3368_0;
	wire w_dff_A_L0BiFdBL6_0;
	wire w_dff_A_iW3Ri9iE7_0;
	wire w_dff_A_xoUAkCg02_0;
	wire w_dff_A_K3HezAHJ7_0;
	wire w_dff_A_HGeg1hHW6_0;
	wire w_dff_A_gL9w6xVe1_0;
	wire w_dff_A_w2bfYK5X3_0;
	wire w_dff_A_rkplaC5G5_0;
	wire w_dff_A_9rwQQ0ko5_0;
	wire w_dff_A_WZktrhNT6_0;
	wire w_dff_B_XzZDx8md5_1;
	wire w_dff_A_S8SNoUsr9_0;
	wire w_dff_A_wpuGUwG39_0;
	wire w_dff_A_FvzflmIP5_0;
	wire w_dff_A_X1Fed3WN2_0;
	wire w_dff_A_4EEzFBoY1_0;
	wire w_dff_A_4guQfGBD0_0;
	wire w_dff_A_wS0E1z5y9_0;
	wire w_dff_A_YrXEYsNd4_0;
	wire w_dff_A_OjWPk9ni2_0;
	wire w_dff_A_YignJEAz3_0;
	wire w_dff_A_UPRj53l43_0;
	wire w_dff_A_RHGOpSsd7_0;
	wire w_dff_A_4aoOijak7_0;
	wire w_dff_A_6Ja7ZXuS3_0;
	wire w_dff_A_pWKTwEMx6_0;
	wire w_dff_A_7gdt2f474_0;
	wire w_dff_A_4U1aKAbU6_0;
	wire w_dff_A_28mJBR7X3_0;
	wire w_dff_A_0vlo5Euv3_0;
	wire w_dff_A_b3Uh1PC65_0;
	wire w_dff_A_GzMRwxlk0_0;
	wire w_dff_A_Y1PZdxHC4_0;
	wire w_dff_A_pUfXEeqD8_0;
	wire w_dff_B_qxEaHlTH9_1;
	wire w_dff_A_TgP2QZxM9_0;
	wire w_dff_A_0OEhDnkf8_0;
	wire w_dff_A_OZmavzp60_0;
	wire w_dff_A_dUy6AJW28_0;
	wire w_dff_A_eGm3zfLS4_0;
	wire w_dff_A_Z04TkIfy3_0;
	wire w_dff_A_we4WEDFt3_0;
	wire w_dff_A_KjXsNrp10_0;
	wire w_dff_A_rjJE9DLc2_0;
	wire w_dff_A_glNc0pJw3_0;
	wire w_dff_A_BEOL1gef2_0;
	wire w_dff_A_617rBd9v6_0;
	wire w_dff_A_gUGhPz4P7_0;
	wire w_dff_A_SIE3Puh01_0;
	wire w_dff_A_DuFthvhz9_0;
	wire w_dff_A_byQnZsMu2_0;
	wire w_dff_A_ggmsijOl8_0;
	wire w_dff_A_HEERYzqX3_0;
	wire w_dff_A_07ryFYOn6_0;
	wire w_dff_A_9FZh6byn6_0;
	wire w_dff_B_r4hNDjzn8_1;
	wire w_dff_A_I8DUMGoX0_0;
	wire w_dff_A_Lq53wyEv9_0;
	wire w_dff_A_ZDDJNgU28_0;
	wire w_dff_A_lIx0bLKJ0_0;
	wire w_dff_A_MfRrB5g66_0;
	wire w_dff_A_Y63wSNTp3_0;
	wire w_dff_A_iwE2BmLL0_0;
	wire w_dff_A_I1qV6Jaa1_0;
	wire w_dff_A_yRNag3fp1_0;
	wire w_dff_A_RlUYuPSY5_0;
	wire w_dff_A_rAoiwxM79_0;
	wire w_dff_A_k0fiZLEa3_0;
	wire w_dff_A_aFVBh2xO5_0;
	wire w_dff_A_9jfXyD3y3_0;
	wire w_dff_A_U1tuxpQ13_0;
	wire w_dff_A_ZGD17F2e9_0;
	wire w_dff_A_nhN25l222_0;
	wire w_dff_B_3vhxBByS6_1;
	wire w_dff_A_Ps0Tcvho8_0;
	wire w_dff_A_25z5P6Bh1_0;
	wire w_dff_A_WkQvTt551_0;
	wire w_dff_A_npWI4njK8_0;
	wire w_dff_A_YRLimjjR8_0;
	wire w_dff_A_jBdQNVfI9_0;
	wire w_dff_A_7PdzuaE90_0;
	wire w_dff_A_nA7dc5BY9_0;
	wire w_dff_A_jhRbLA6Q7_0;
	wire w_dff_A_4EuBYuut9_0;
	wire w_dff_A_yhwUhhM33_0;
	wire w_dff_A_m062pSjM0_0;
	wire w_dff_A_Usx6TU591_0;
	wire w_dff_A_xTHqHmzl2_0;
	wire w_dff_B_HfKmuf415_1;
	wire w_dff_A_0qNLck1J0_0;
	wire w_dff_A_17ZMACWF0_0;
	wire w_dff_A_Gc39vKPx9_0;
	wire w_dff_A_RtNC1uB15_0;
	wire w_dff_A_PV9EYaJr3_0;
	wire w_dff_A_OMyJ6xQq8_0;
	wire w_dff_A_UFZvJpGt8_0;
	wire w_dff_A_E2NoMfwW0_0;
	wire w_dff_A_jALWbNxy6_0;
	wire w_dff_A_Ub9v0iXs2_0;
	wire w_dff_A_uGHgRN7S4_0;
	wire w_dff_B_BZ4iv02w0_1;
	wire w_dff_A_DMVcyFUf3_0;
	wire w_dff_A_mIiBCANF5_0;
	wire w_dff_A_oJ5GVM8I1_0;
	wire w_dff_A_lfYOIB5d5_0;
	wire w_dff_A_3gPfbbnv4_0;
	wire w_dff_A_kYqYKoxr2_0;
	wire w_dff_A_yz2g5o3T1_0;
	wire w_dff_A_OcGInJTO8_0;
	wire w_dff_B_lka824er8_1;
	wire w_dff_A_ZdyDGYRF6_0;
	wire w_dff_A_7RScKASn6_0;
	wire w_dff_A_G0LNzcrn8_0;
	wire w_dff_A_wyHhALjm2_0;
	wire w_dff_B_AsRBWcbj0_0;
	wire w_dff_A_iGsqUyTS8_0;
	wire w_dff_A_kHDRHVTJ0_0;
	wire w_dff_B_cMjIhJEV7_2;
	wire w_dff_B_sWP56mRH1_2;
	wire w_dff_B_z2gJh9B52_2;
	wire w_dff_B_s9MKeXFT0_2;
	wire w_dff_B_BlJtStrS9_2;
	wire w_dff_B_4ZrApfOc7_2;
	wire w_dff_B_8WTIScRC8_2;
	wire w_dff_B_aaE8ibXH6_2;
	wire w_dff_B_p8XQ9mHl2_2;
	wire w_dff_B_rsoZITgZ2_2;
	wire w_dff_B_jskZ009W2_2;
	wire w_dff_B_xaX5NC4Z6_2;
	wire w_dff_B_zVOHL91y4_2;
	wire w_dff_B_AoneoiBe9_2;
	wire w_dff_B_oa4YAf3i9_2;
	wire w_dff_B_JsRxpWHk4_2;
	wire w_dff_B_V75BtALJ3_2;
	wire w_dff_B_wMJb6RMj2_2;
	wire w_dff_B_C2abLtti9_2;
	wire w_dff_B_aiyDfmbh1_2;
	wire w_dff_B_kFzdtis48_2;
	wire w_dff_B_9puinoJx4_2;
	wire w_dff_B_PJWfu2Pf8_2;
	wire w_dff_B_DYGmZ1rB0_2;
	wire w_dff_B_9ImUXCEc7_2;
	wire w_dff_B_AqnN7G0m1_2;
	wire w_dff_B_AGVbdhUS4_2;
	wire w_dff_B_ItjhBvyb7_2;
	wire w_dff_B_q11eEC790_2;
	wire w_dff_B_GlJLWQMp1_2;
	wire w_dff_B_w76aUxrT4_2;
	wire w_dff_B_0gDijboI2_2;
	wire w_dff_B_jGYKGauk4_2;
	wire w_dff_B_rLjNOMb91_2;
	wire w_dff_B_zAdSHiSq5_2;
	wire w_dff_B_2emaucSo3_2;
	wire w_dff_B_Eevua5uk6_2;
	wire w_dff_B_shMmYz582_2;
	wire w_dff_B_NZ4Gurnf1_2;
	wire w_dff_B_htANaIDt2_2;
	wire w_dff_B_lJ5FMkbB7_2;
	wire w_dff_B_F9pzeo6i8_2;
	wire w_dff_B_eu71PbNQ2_2;
	wire w_dff_B_SYqhYXJy0_2;
	wire w_dff_A_pjjutMCB9_0;
	wire w_dff_B_YGBk4d6B0_1;
	wire w_dff_B_DNzvvfS67_2;
	wire w_dff_B_9PEsjT5o3_2;
	wire w_dff_B_F9IZMHeN6_2;
	wire w_dff_B_n4xbpcwy0_2;
	wire w_dff_B_TX0PA1M27_2;
	wire w_dff_B_s0ldgvR69_2;
	wire w_dff_B_ufuef6bT3_2;
	wire w_dff_B_AWDttdoo6_2;
	wire w_dff_B_46xmwMo04_2;
	wire w_dff_B_DdNHP23u2_2;
	wire w_dff_B_3si6Bylu5_2;
	wire w_dff_B_6md3Pfvk6_2;
	wire w_dff_B_zMoJKukp6_2;
	wire w_dff_B_T7pmnkJE6_2;
	wire w_dff_B_pJFDvR551_2;
	wire w_dff_B_XdTbbgsw2_2;
	wire w_dff_B_3GcBCU8N6_2;
	wire w_dff_B_ONcR3NhH2_2;
	wire w_dff_B_mKjN1i3f4_2;
	wire w_dff_B_bLNxqumJ4_2;
	wire w_dff_B_bBPrEfQk3_2;
	wire w_dff_B_dfR48Bq79_2;
	wire w_dff_B_tkF1pB0Z6_2;
	wire w_dff_B_4DlmKAeM9_2;
	wire w_dff_B_6oKVEMCU6_2;
	wire w_dff_B_EnQPCE8p7_2;
	wire w_dff_B_cHf5ylHZ9_2;
	wire w_dff_B_BAK4Yd0c4_2;
	wire w_dff_B_SlQVWnTe7_2;
	wire w_dff_B_S8kf8kxz5_2;
	wire w_dff_B_fsWyEvLm5_2;
	wire w_dff_B_kvg1jy7G3_2;
	wire w_dff_B_zxP7er6f1_2;
	wire w_dff_B_lYmcxQpE6_2;
	wire w_dff_B_dDExMTO48_2;
	wire w_dff_B_vl2mcgNi2_2;
	wire w_dff_B_TgsGOfhP3_2;
	wire w_dff_B_DyxWsHIf6_2;
	wire w_dff_B_aPoveLqF9_2;
	wire w_dff_B_h1Ll7FdX5_2;
	wire w_dff_A_hK4FPsXJ4_1;
	wire w_dff_A_IkfscCdt0_0;
	wire w_dff_A_o7mAy3Ez9_0;
	wire w_dff_A_0GxAqjJG5_0;
	wire w_dff_A_5SACCQAh5_0;
	wire w_dff_A_Ik0Oth9e5_0;
	wire w_dff_A_nsYC6Hbg7_0;
	wire w_dff_A_An1SyVrE2_0;
	wire w_dff_A_M7gSdpXs0_0;
	wire w_dff_A_5rpS1fqF4_0;
	wire w_dff_A_pSdRuKNy8_0;
	wire w_dff_A_XKVGVf5W9_0;
	wire w_dff_A_VWHnLsL63_0;
	wire w_dff_A_WEnicOu88_0;
	wire w_dff_A_1zrSoqdJ3_0;
	wire w_dff_A_yVQzp8SB4_0;
	wire w_dff_A_xslBY8zI0_0;
	wire w_dff_A_35C7cfdF6_0;
	wire w_dff_A_8cBoGORk7_0;
	wire w_dff_A_egw93r2D5_0;
	wire w_dff_A_WZxTySWC9_0;
	wire w_dff_A_DZBG9ZFJ8_0;
	wire w_dff_A_R99VK25B9_0;
	wire w_dff_A_wHvWHxvY7_0;
	wire w_dff_A_Q1y6kjRc2_0;
	wire w_dff_A_JRrZcsmk8_0;
	wire w_dff_A_LYjliNrx4_0;
	wire w_dff_A_vGqp6JRk5_0;
	wire w_dff_A_mR8NV3dy0_0;
	wire w_dff_A_lBdYvBH87_0;
	wire w_dff_A_RC3CelW55_0;
	wire w_dff_A_YHXS3FzX4_0;
	wire w_dff_A_WlHj1mDf7_0;
	wire w_dff_A_eaK2RJ0m7_0;
	wire w_dff_A_uca9syKp0_0;
	wire w_dff_A_lio901276_0;
	wire w_dff_A_1EnTW8GZ1_0;
	wire w_dff_A_4lszyFn33_0;
	wire w_dff_A_PaeTrKK39_1;
	wire w_dff_A_1ezDC40J1_2;
	wire w_dff_B_S4ORdUCC3_1;
	wire w_dff_B_OKyzk8Am3_2;
	wire w_dff_B_QrOMOxpq3_2;
	wire w_dff_B_HQ5mZaLc5_2;
	wire w_dff_B_mWzklsGZ8_2;
	wire w_dff_B_sPbXZwBI1_2;
	wire w_dff_B_Hy6mtHDx0_2;
	wire w_dff_B_x3l5EV4w5_2;
	wire w_dff_B_4cEYmsvB1_2;
	wire w_dff_B_8MIdHzbJ5_2;
	wire w_dff_B_kdifOqQd7_2;
	wire w_dff_B_vrR4YgeA2_2;
	wire w_dff_B_lJIkTdyN4_2;
	wire w_dff_B_jDm2Xwa08_2;
	wire w_dff_B_RYTP8VTC3_2;
	wire w_dff_B_HFKsYVuF3_2;
	wire w_dff_B_I4ktasz51_2;
	wire w_dff_B_nw3p254o3_2;
	wire w_dff_B_QimNdpqH1_2;
	wire w_dff_B_mbMrcQet5_2;
	wire w_dff_B_dy8Lzjex8_2;
	wire w_dff_B_30BLDKRy9_2;
	wire w_dff_B_1NGgOigZ9_2;
	wire w_dff_B_FN4SjH7s3_2;
	wire w_dff_B_Ppqrb9gF4_2;
	wire w_dff_B_ikvOKAlh6_2;
	wire w_dff_B_3TVZMWGu1_2;
	wire w_dff_B_KW8k5q2W6_2;
	wire w_dff_B_JAMLgE5S9_2;
	wire w_dff_B_xLQ3FboZ2_2;
	wire w_dff_B_SuUU2NdK7_2;
	wire w_dff_B_6GiWr4pP6_2;
	wire w_dff_B_iI2UZcQj6_2;
	wire w_dff_B_48MqtL2S3_2;
	wire w_dff_B_Ch8v8ZGe5_2;
	wire w_dff_B_HgCApr8i9_1;
	wire w_dff_B_7rpKxDZC5_2;
	wire w_dff_B_PA0FYVIU6_2;
	wire w_dff_B_udIlobvs4_2;
	wire w_dff_B_4RYQuMem5_2;
	wire w_dff_B_CrwMvU7m9_2;
	wire w_dff_B_tNMH12mS0_2;
	wire w_dff_B_l5jHD8MR4_2;
	wire w_dff_B_qePmiZwV4_2;
	wire w_dff_B_OLuMQmi39_2;
	wire w_dff_B_8KIr8lb44_2;
	wire w_dff_B_czveACIn4_2;
	wire w_dff_B_hAZy3l651_2;
	wire w_dff_B_NQ8nkmsP1_2;
	wire w_dff_B_fk6Cz92y8_2;
	wire w_dff_B_ZqHVFzJZ2_2;
	wire w_dff_B_mTFfpFVL5_2;
	wire w_dff_B_GDRo23Pv9_2;
	wire w_dff_B_QiA1G6pS1_2;
	wire w_dff_B_niBFkt3b7_2;
	wire w_dff_B_QKoQBLWg2_2;
	wire w_dff_B_HEmFGvd54_2;
	wire w_dff_B_mKI4ZSl27_2;
	wire w_dff_B_jULFZCLS9_2;
	wire w_dff_B_KtQEJS3O6_2;
	wire w_dff_B_IYezIVQ78_2;
	wire w_dff_B_foWNZZ9p7_2;
	wire w_dff_B_UZL6lfpx4_2;
	wire w_dff_B_ZPYN26713_2;
	wire w_dff_B_ellVHP0T5_2;
	wire w_dff_B_QaEcDSuD5_2;
	wire w_dff_B_TJA2DPQ43_2;
	wire w_dff_B_AAk7rBFR0_1;
	wire w_dff_B_ZWLLn9iO4_2;
	wire w_dff_B_B5DJdmPx2_2;
	wire w_dff_B_B0ltlHbD7_2;
	wire w_dff_B_rtksfZyz1_2;
	wire w_dff_B_IZqBLimd3_2;
	wire w_dff_B_L5uThb3m5_2;
	wire w_dff_B_edTWyWv18_2;
	wire w_dff_B_oXxetAOU7_2;
	wire w_dff_B_buIo5cxD3_2;
	wire w_dff_B_OzSw6qXi9_2;
	wire w_dff_B_TiI6N7T87_2;
	wire w_dff_B_RCrHm3Xz7_2;
	wire w_dff_B_it2SQyoQ9_2;
	wire w_dff_B_QMs1OM2m9_2;
	wire w_dff_B_ybz9E4168_2;
	wire w_dff_B_zgUtsPIU0_2;
	wire w_dff_B_95oHT9fe1_2;
	wire w_dff_B_eRILAvIh6_2;
	wire w_dff_B_Md6ppQSk7_2;
	wire w_dff_B_etzLcrmj9_2;
	wire w_dff_B_SinFgzVt4_2;
	wire w_dff_B_SvLkIe8e0_2;
	wire w_dff_B_1q12hnRw7_2;
	wire w_dff_B_xBntAbYr8_2;
	wire w_dff_B_An2QI8fG8_2;
	wire w_dff_B_ehX91O2y4_2;
	wire w_dff_B_SabJs8jz7_2;
	wire w_dff_B_hR5poCbV0_2;
	wire w_dff_B_E0zn4wyP8_1;
	wire w_dff_B_ZZyPhveW8_2;
	wire w_dff_B_MIqa1AyF2_2;
	wire w_dff_B_qBmtmQtj2_2;
	wire w_dff_B_rd3rvPc38_2;
	wire w_dff_B_usGTkVpu1_2;
	wire w_dff_B_825KKHae9_2;
	wire w_dff_B_N8ROcOzd9_2;
	wire w_dff_B_xYtmxULo3_2;
	wire w_dff_B_nrQD752S8_2;
	wire w_dff_B_EMqMMHyE5_2;
	wire w_dff_B_Q106ELUE1_2;
	wire w_dff_B_uaLusQio5_2;
	wire w_dff_B_q8welTEc0_2;
	wire w_dff_B_oDDvjCoj2_2;
	wire w_dff_B_8HwWkaG32_2;
	wire w_dff_B_MIVvcWb63_2;
	wire w_dff_B_B0z1MmyT0_2;
	wire w_dff_B_9EBzyWvx7_2;
	wire w_dff_B_5monQgmX4_2;
	wire w_dff_B_rmr0cjqc3_2;
	wire w_dff_B_ULDb7L4G2_2;
	wire w_dff_B_TtEmYi327_2;
	wire w_dff_B_w0Tkh8XO5_2;
	wire w_dff_B_q57hWTjr9_2;
	wire w_dff_B_0xyfVBWM7_2;
	wire w_dff_B_Jh6lq4521_1;
	wire w_dff_B_lANTmmel5_2;
	wire w_dff_B_0ZG2LOSb2_2;
	wire w_dff_B_c7ztxUz32_2;
	wire w_dff_B_sXmtubWl5_2;
	wire w_dff_B_yb5GS2Gt2_2;
	wire w_dff_B_mtJ3BfXa4_2;
	wire w_dff_B_KDc0nzDV6_2;
	wire w_dff_B_k8XBaHQ05_2;
	wire w_dff_B_lJSoHneo5_2;
	wire w_dff_B_NSEFXBjI0_2;
	wire w_dff_B_rMwsg27l6_2;
	wire w_dff_B_BgW5oD0n5_2;
	wire w_dff_B_KZPQY57t3_2;
	wire w_dff_B_B70Eamoi1_2;
	wire w_dff_B_Jl3RscIH9_2;
	wire w_dff_B_LcQSTCgc3_2;
	wire w_dff_B_UduQqCAt0_2;
	wire w_dff_B_mzj2trgd0_2;
	wire w_dff_B_uUV632eO3_2;
	wire w_dff_B_KPaKpPg85_2;
	wire w_dff_B_TLAx6knM4_2;
	wire w_dff_B_1M3mdTob1_2;
	wire w_dff_B_ZPrv69rY1_1;
	wire w_dff_B_lLyytNMO4_2;
	wire w_dff_B_q9Gu2eiS7_2;
	wire w_dff_B_Qnk4Z3XI8_2;
	wire w_dff_B_JDG4hyvH6_2;
	wire w_dff_B_YibEVKDh6_2;
	wire w_dff_B_mbI4Fcqw5_2;
	wire w_dff_B_TYspeDOi8_2;
	wire w_dff_B_I7HuwlUW0_2;
	wire w_dff_B_ZJeV8KQq0_2;
	wire w_dff_B_UyzBVT2o6_2;
	wire w_dff_B_D39Jdf8i9_2;
	wire w_dff_B_0ErRhg7G6_2;
	wire w_dff_B_V8zmzqOd3_2;
	wire w_dff_B_vlvm1FA74_2;
	wire w_dff_B_Odve1Lhe6_2;
	wire w_dff_B_delXOXpE8_2;
	wire w_dff_B_bvDYa1ZN5_2;
	wire w_dff_B_ciueZflC7_2;
	wire w_dff_B_sqKLcQOC4_2;
	wire w_dff_B_TLyREf666_1;
	wire w_dff_B_IrrZjGgS5_2;
	wire w_dff_B_cGe2yHM70_2;
	wire w_dff_B_1wgzXjHn1_2;
	wire w_dff_B_1jjrzbDi0_2;
	wire w_dff_B_heFUKkxg4_2;
	wire w_dff_B_1VszxwXr2_2;
	wire w_dff_B_csLb90T36_2;
	wire w_dff_B_R6PbYK4y9_2;
	wire w_dff_B_T7akaYFz9_2;
	wire w_dff_B_4HVlGHnt6_2;
	wire w_dff_B_IfJ7XFg28_2;
	wire w_dff_B_YFvkUf2B4_2;
	wire w_dff_B_vQSkTbsO0_2;
	wire w_dff_B_gOonVgmw2_2;
	wire w_dff_B_DlfQu4jH3_2;
	wire w_dff_B_jQbxvzmW2_2;
	wire w_dff_B_genMed2k6_1;
	wire w_dff_B_euvDCGwU1_2;
	wire w_dff_B_jm1HdqEf7_2;
	wire w_dff_B_PvityzRU3_2;
	wire w_dff_B_fbqMY5Fy7_2;
	wire w_dff_B_XlrAH4nN9_2;
	wire w_dff_B_VDOgafZk5_2;
	wire w_dff_B_yIxQC1JB1_2;
	wire w_dff_B_R9KdxMF81_2;
	wire w_dff_B_PFtbiEVC2_2;
	wire w_dff_B_qmSAHCoo1_2;
	wire w_dff_B_YeWPrfTF1_2;
	wire w_dff_B_4w5HXiWm6_2;
	wire w_dff_B_tnSzTt9L3_2;
	wire w_dff_B_wrVJX94M6_1;
	wire w_dff_B_895YVFTo0_2;
	wire w_dff_B_4s2w8K9Y7_2;
	wire w_dff_B_ZI8ipCT06_2;
	wire w_dff_B_bX9VQi0l8_2;
	wire w_dff_B_3eTLC9ts9_2;
	wire w_dff_B_042cQft63_2;
	wire w_dff_B_Acj0Q3uf9_2;
	wire w_dff_B_Hotdf22T6_2;
	wire w_dff_B_e4Sw9TXZ8_2;
	wire w_dff_B_ezZqCDx86_2;
	wire w_dff_B_APnmgULd0_1;
	wire w_dff_B_4chyMujv4_2;
	wire w_dff_B_OyqFo2pv3_2;
	wire w_dff_B_YlC1PFSL0_2;
	wire w_dff_B_hgHBTYbN4_2;
	wire w_dff_B_RwhEWNGK6_2;
	wire w_dff_B_NaR232Rg3_2;
	wire w_dff_B_Z5Otzmzb1_2;
	wire w_dff_B_577uiCVg7_2;
	wire w_dff_B_sx2C9rLO4_2;
	wire w_dff_B_O43b9nPM6_2;
	wire w_dff_B_dzB81Hgh7_0;
	wire w_dff_B_LoIPBci80_0;
	wire w_dff_A_qpxHJBxk7_1;
	wire w_dff_A_2JNqYLSr2_1;
	wire w_dff_B_1fupoCDN4_1;
	wire w_dff_B_bDw6z2Oz2_1;
	wire w_dff_B_agULwE7d2_2;
	wire w_dff_B_9G69aGdd5_2;
	wire w_dff_B_tKOA0cNV7_2;
	wire w_dff_B_I8NQoZMb0_2;
	wire w_dff_B_3d7BK34F9_2;
	wire w_dff_B_Z7r1eV5q3_2;
	wire w_dff_B_0Lb0Z4XO1_2;
	wire w_dff_B_nQFnVsln3_2;
	wire w_dff_B_Kb7Zeb3Y6_2;
	wire w_dff_B_2X3IdqpE8_2;
	wire w_dff_B_AM3Gsmgg2_2;
	wire w_dff_B_js2o9Z0f2_2;
	wire w_dff_B_jABkcMLU9_2;
	wire w_dff_B_GEq0rs3t1_2;
	wire w_dff_B_z3jHJwCv0_2;
	wire w_dff_B_OsDbvXug6_2;
	wire w_dff_B_yCyNaL3H4_2;
	wire w_dff_B_qc7t4wag4_2;
	wire w_dff_B_zNShhUgA5_2;
	wire w_dff_B_ZfHSKcpl7_2;
	wire w_dff_B_4nWPXNbs0_2;
	wire w_dff_B_p2gXxWfN5_2;
	wire w_dff_B_zJyTFgA67_2;
	wire w_dff_B_rz3cbqO80_2;
	wire w_dff_B_6zMnba1y1_2;
	wire w_dff_B_79eag0Im4_2;
	wire w_dff_B_s7YJnI191_2;
	wire w_dff_B_QQAIagTG4_2;
	wire w_dff_B_1lIRuHz28_2;
	wire w_dff_B_IidVnOHl6_2;
	wire w_dff_B_Tp1iF3st0_2;
	wire w_dff_B_WkK6Jg3g3_2;
	wire w_dff_B_lH4z1VnS0_2;
	wire w_dff_B_rEbARcMs4_2;
	wire w_dff_B_g7WqY3Vk1_2;
	wire w_dff_B_NUMWLlKW5_2;
	wire w_dff_B_JrUy5QGY1_2;
	wire w_dff_B_aPPa0fvm0_2;
	wire w_dff_B_7H0YXTN93_2;
	wire w_dff_B_1nH08Sja8_2;
	wire w_dff_B_XG3sNIfl3_2;
	wire w_dff_B_yXpJVcTT4_2;
	wire w_dff_B_R2JGXC7W8_2;
	wire w_dff_B_Yl0vInWa3_2;
	wire w_dff_B_wGGF3adj5_2;
	wire w_dff_B_cdwtbpXo2_2;
	wire w_dff_B_DqGxwHbC1_1;
	wire w_dff_B_VV78izEa9_2;
	wire w_dff_B_JMfHh7yQ0_2;
	wire w_dff_B_ZYCJzGjH1_2;
	wire w_dff_B_wf8qKgqo5_2;
	wire w_dff_B_Ob14SXDA6_2;
	wire w_dff_B_H8wrZPF16_2;
	wire w_dff_B_t6MrAjES9_2;
	wire w_dff_B_XnWuqa858_2;
	wire w_dff_B_kZDBTZal0_2;
	wire w_dff_B_6yvoHXFB8_2;
	wire w_dff_B_kmO6vQG50_2;
	wire w_dff_B_4k5jc4My3_2;
	wire w_dff_B_vr977IGf2_2;
	wire w_dff_B_nSYaRnhO1_2;
	wire w_dff_B_vJ78mm8x6_2;
	wire w_dff_B_RyP6E7gn7_2;
	wire w_dff_B_Myshnbe47_2;
	wire w_dff_B_qKkLw8Kc0_2;
	wire w_dff_B_IisZFHk28_2;
	wire w_dff_B_173zE3wI9_2;
	wire w_dff_B_iRmfp9v25_2;
	wire w_dff_B_Q9WrxAtQ0_2;
	wire w_dff_B_IneNu71y8_2;
	wire w_dff_B_u2K4lrpV7_2;
	wire w_dff_B_gfMryNpa4_2;
	wire w_dff_B_fRjP8YWz6_2;
	wire w_dff_B_D5pOJyV48_2;
	wire w_dff_B_lrRpCMSJ2_2;
	wire w_dff_B_Xvy2Y6VW9_2;
	wire w_dff_B_kapuTbQO3_2;
	wire w_dff_B_XGW6OSEY6_2;
	wire w_dff_B_vCc9X8W45_2;
	wire w_dff_B_it0Mh74z4_2;
	wire w_dff_B_hFTNOiXp8_2;
	wire w_dff_B_r37wjaCq0_2;
	wire w_dff_B_xdNBrZCi3_2;
	wire w_dff_B_hbOlwcAs2_2;
	wire w_dff_B_czKOHofc8_2;
	wire w_dff_B_ygtjzrFC1_2;
	wire w_dff_B_QYiA9Km83_2;
	wire w_dff_B_73M7BQO13_2;
	wire w_dff_B_falzzeP72_2;
	wire w_dff_B_hUWPJ5Ia0_1;
	wire w_dff_B_38pXlEXW0_2;
	wire w_dff_B_Crpe4JDv4_2;
	wire w_dff_B_97xQvbry6_2;
	wire w_dff_B_mrqPKc1Z9_2;
	wire w_dff_B_jt0FEUrP4_2;
	wire w_dff_B_mGJMO9eB6_2;
	wire w_dff_B_RT6MvAg04_2;
	wire w_dff_B_1LtO1l2e5_2;
	wire w_dff_B_Q2eDYiTU0_2;
	wire w_dff_B_ezHkWKvm5_2;
	wire w_dff_B_M6PcMdri6_2;
	wire w_dff_B_P3VgKcs09_2;
	wire w_dff_B_yBk1mHDO0_2;
	wire w_dff_B_BlxQOUZS7_2;
	wire w_dff_B_ltFOv6Vo1_2;
	wire w_dff_B_4J8Yf2W26_2;
	wire w_dff_B_BYr64GK65_2;
	wire w_dff_B_8rB9nKcx1_2;
	wire w_dff_B_wqUHvkBj8_2;
	wire w_dff_B_ywuXpUg47_2;
	wire w_dff_B_8gURS7ci2_2;
	wire w_dff_B_7jpLkQnA1_2;
	wire w_dff_B_ZxD3NAAN4_2;
	wire w_dff_B_V06AWYwM1_2;
	wire w_dff_B_9SUaudRb2_2;
	wire w_dff_B_VrWv7SJo9_2;
	wire w_dff_B_Apnxg2Su3_2;
	wire w_dff_B_a4hT12As6_2;
	wire w_dff_B_iJMMg6Ci0_2;
	wire w_dff_B_udsFMJq63_2;
	wire w_dff_B_nh31iq2e9_2;
	wire w_dff_B_3OVzZOA39_2;
	wire w_dff_B_HTKKiomk7_2;
	wire w_dff_B_35qTgeS53_2;
	wire w_dff_B_Zn1pUUIV4_2;
	wire w_dff_B_TERMiXSN4_2;
	wire w_dff_B_0s0TzxQu7_2;
	wire w_dff_B_kcbxlRjy9_1;
	wire w_dff_B_sXUB0K114_2;
	wire w_dff_B_YYgudbEX2_2;
	wire w_dff_B_vJXMOotG0_2;
	wire w_dff_B_NTZ2dVIL2_2;
	wire w_dff_B_X4nHCl4w9_2;
	wire w_dff_B_gAE62IgG1_2;
	wire w_dff_B_aQZGDkUz8_2;
	wire w_dff_B_onVMGKRj3_2;
	wire w_dff_B_FgjOxEOF1_2;
	wire w_dff_B_bfyIWMSJ1_2;
	wire w_dff_B_xDZnBuEW5_2;
	wire w_dff_B_GErPVUKH1_2;
	wire w_dff_B_Gd7Hg6vj8_2;
	wire w_dff_B_pMVFnvOx5_2;
	wire w_dff_B_AehMOhl39_2;
	wire w_dff_B_TpH9i84D8_2;
	wire w_dff_B_AQPdMPZB4_2;
	wire w_dff_B_GU4ROdY50_2;
	wire w_dff_B_hoyULrMt1_2;
	wire w_dff_B_REC2RIuZ3_2;
	wire w_dff_B_3WRI4TEW0_2;
	wire w_dff_B_AOovrG2I8_2;
	wire w_dff_B_iVdF1zSj9_2;
	wire w_dff_B_CSJejrr00_2;
	wire w_dff_B_TmgQY7aq7_2;
	wire w_dff_B_h0FRUO3j1_2;
	wire w_dff_B_cxljlFJk5_2;
	wire w_dff_B_YT0MdckA4_2;
	wire w_dff_B_G4X87IfJ0_2;
	wire w_dff_B_CXA7bD8E7_2;
	wire w_dff_B_Kr04a6zH7_2;
	wire w_dff_B_wiemeGC85_2;
	wire w_dff_B_6PAvUIMV1_2;
	wire w_dff_B_2oTC1IeI8_2;
	wire w_dff_B_ga3xMME42_1;
	wire w_dff_B_vTMbvAtu7_2;
	wire w_dff_B_G4nAPH1o3_2;
	wire w_dff_B_NnmeNfwY3_2;
	wire w_dff_B_rfwclIUl9_2;
	wire w_dff_B_2qcbZqSG7_2;
	wire w_dff_B_Jv9X6WHL8_2;
	wire w_dff_B_7tMLKjnG5_2;
	wire w_dff_B_7001iSvU5_2;
	wire w_dff_B_i7ycTdzN4_2;
	wire w_dff_B_IIDlM1ND3_2;
	wire w_dff_B_9dRHixW77_2;
	wire w_dff_B_PYVcYUhh0_2;
	wire w_dff_B_6uRsDfVo0_2;
	wire w_dff_B_bIISXcli7_2;
	wire w_dff_B_Et2FDZtn3_2;
	wire w_dff_B_8qZZ8Nt57_2;
	wire w_dff_B_AERnxkmb3_2;
	wire w_dff_B_dpix5o353_2;
	wire w_dff_B_XSC01LDr4_2;
	wire w_dff_B_VzC8j6nj0_2;
	wire w_dff_B_rXnnaJ8p2_2;
	wire w_dff_B_99nxWuam3_2;
	wire w_dff_B_7xjFRmPL5_2;
	wire w_dff_B_mRuCOBGJ1_2;
	wire w_dff_B_oXeNmgWz7_2;
	wire w_dff_B_ycWV6Zts4_2;
	wire w_dff_B_fZhepIFF1_2;
	wire w_dff_B_5V2BFPIT7_2;
	wire w_dff_B_MY9aCvZg6_2;
	wire w_dff_B_dn6khCWy1_2;
	wire w_dff_B_kQ3pLChE1_2;
	wire w_dff_B_72vJHDRm4_1;
	wire w_dff_B_WNXECbNp2_2;
	wire w_dff_B_6yy8D0MW7_2;
	wire w_dff_B_095mUswf9_2;
	wire w_dff_B_ra6e7fzJ3_2;
	wire w_dff_B_bnGmFO3i5_2;
	wire w_dff_B_dIlXzTbE6_2;
	wire w_dff_B_ke0Ex4BD3_2;
	wire w_dff_B_KAHiQ5MD5_2;
	wire w_dff_B_bQJjeAAb6_2;
	wire w_dff_B_S8pShqH10_2;
	wire w_dff_B_MxzhyBte1_2;
	wire w_dff_B_jbY18xuA5_2;
	wire w_dff_B_GjZpbovM5_2;
	wire w_dff_B_NsfHKnrZ2_2;
	wire w_dff_B_WaTfX6FN6_2;
	wire w_dff_B_arKz1MVK2_2;
	wire w_dff_B_Ud9JqVjp2_2;
	wire w_dff_B_wf0MDSsA7_2;
	wire w_dff_B_GvL24ZfN1_2;
	wire w_dff_B_M83a0Eab1_2;
	wire w_dff_B_ME0FJdGH6_2;
	wire w_dff_B_mQ5KoUqM3_2;
	wire w_dff_B_87p6jvvS3_2;
	wire w_dff_B_0HG02Vwh6_2;
	wire w_dff_B_UfNS9ONN4_2;
	wire w_dff_B_Toz374d67_2;
	wire w_dff_B_SVn0Kq5S2_2;
	wire w_dff_B_QMXPycXa7_2;
	wire w_dff_B_pzUmcCNM8_1;
	wire w_dff_B_C42Mg9dF7_2;
	wire w_dff_B_pVjvpTb82_2;
	wire w_dff_B_QZ5Ergr54_2;
	wire w_dff_B_0F1z5oQc6_2;
	wire w_dff_B_UeUDiyVH4_2;
	wire w_dff_B_LanzuH9v9_2;
	wire w_dff_B_z233RMrP0_2;
	wire w_dff_B_NqmiiqCc0_2;
	wire w_dff_B_FkWLYgRS5_2;
	wire w_dff_B_cGomwskl3_2;
	wire w_dff_B_hqs1QI3m7_2;
	wire w_dff_B_SMA1iwBW7_2;
	wire w_dff_B_8CGju51P5_2;
	wire w_dff_B_4P63Sk099_2;
	wire w_dff_B_8RovYKMb4_2;
	wire w_dff_B_fmaC9uC59_2;
	wire w_dff_B_lF1rxL5v7_2;
	wire w_dff_B_Cwkc5HQG3_2;
	wire w_dff_B_aKonAQ029_2;
	wire w_dff_B_qCDbyKzR8_2;
	wire w_dff_B_tmX8AwQQ1_2;
	wire w_dff_B_0YCRTGia0_2;
	wire w_dff_B_dLSiwg0c4_2;
	wire w_dff_B_uGOp2fnT2_2;
	wire w_dff_B_m8OWrTci8_2;
	wire w_dff_B_TF5vSIb98_1;
	wire w_dff_B_tQ4qXZ1x6_2;
	wire w_dff_B_mClwyOzS8_2;
	wire w_dff_B_Kxlplazs1_2;
	wire w_dff_B_N5a60De67_2;
	wire w_dff_B_ektGJC4b7_2;
	wire w_dff_B_kUC2MXDG0_2;
	wire w_dff_B_BWCi4y7u3_2;
	wire w_dff_B_yKfef8Pu0_2;
	wire w_dff_B_Fp8V6JlI0_2;
	wire w_dff_B_DnZORb424_2;
	wire w_dff_B_7p2Mnrod6_2;
	wire w_dff_B_NzmfXrmJ6_2;
	wire w_dff_B_CkSWZqT83_2;
	wire w_dff_B_Gb3iBuFG9_2;
	wire w_dff_B_mOkqK3Gg9_2;
	wire w_dff_B_JWUZTMPr4_2;
	wire w_dff_B_AyP0BeJS5_2;
	wire w_dff_B_2AWjIdOv7_2;
	wire w_dff_B_oh0qzwZ21_2;
	wire w_dff_B_2gms4NKT4_2;
	wire w_dff_B_1obje77m9_2;
	wire w_dff_B_yR9CiLXM5_2;
	wire w_dff_B_dbiXsX4n4_1;
	wire w_dff_B_S6ClhJNw1_2;
	wire w_dff_B_WSKv8KBR4_2;
	wire w_dff_B_xbLX4O0F3_2;
	wire w_dff_B_S23IViRA3_2;
	wire w_dff_B_W2KmOD0e8_2;
	wire w_dff_B_8F2KyJNg0_2;
	wire w_dff_B_cCmCpYAe2_2;
	wire w_dff_B_4ViM8jpT8_2;
	wire w_dff_B_iqCsRr4K0_2;
	wire w_dff_B_b3U0LBdv4_2;
	wire w_dff_B_GxMsT4im8_2;
	wire w_dff_B_esmiuX8b5_2;
	wire w_dff_B_3HHKbp6f0_2;
	wire w_dff_B_PLmQuOCZ8_2;
	wire w_dff_B_mkCIRXr34_2;
	wire w_dff_B_iOstxyim7_2;
	wire w_dff_B_IV2nnOEA5_2;
	wire w_dff_B_0vg8Nkm94_2;
	wire w_dff_B_a3vhh17j0_2;
	wire w_dff_B_8KXdKmmc6_1;
	wire w_dff_B_81DpVl7v2_2;
	wire w_dff_B_kAjE0D7I4_2;
	wire w_dff_B_RAeSevz53_2;
	wire w_dff_B_IuAArMSN9_2;
	wire w_dff_B_DgacSUbd6_2;
	wire w_dff_B_N6zbtjUG2_2;
	wire w_dff_B_87EYA9Y24_2;
	wire w_dff_B_j7nDCuoL8_2;
	wire w_dff_B_7EixtPTM1_2;
	wire w_dff_B_eJVg4sHJ5_2;
	wire w_dff_B_VMoPedRs6_2;
	wire w_dff_B_01JQ4hfl9_2;
	wire w_dff_B_DjleBzKY8_2;
	wire w_dff_B_c9L2D4CH9_2;
	wire w_dff_B_4GGfpT8Z2_2;
	wire w_dff_B_hUuxM9Cj6_2;
	wire w_dff_B_npBmo3FI2_1;
	wire w_dff_B_RhK0niGN5_2;
	wire w_dff_B_OEwf7hP66_2;
	wire w_dff_B_MtaKCeQ73_2;
	wire w_dff_B_cqrkvAVp5_2;
	wire w_dff_B_NgYT9d8Q1_2;
	wire w_dff_B_K1oAFODJ0_2;
	wire w_dff_B_7lGNjVI75_2;
	wire w_dff_B_kWvFYJsq6_2;
	wire w_dff_B_1vqvDT3b4_2;
	wire w_dff_B_4jZlZdKo0_2;
	wire w_dff_B_eHDaJjSf8_2;
	wire w_dff_B_YuxiLJVP8_2;
	wire w_dff_B_FPWiNprk3_2;
	wire w_dff_B_Y4Mwki8N8_1;
	wire w_dff_B_buPbW46o2_2;
	wire w_dff_B_SDqNf5448_2;
	wire w_dff_B_jdejU4C27_2;
	wire w_dff_B_0AFkGHTD9_2;
	wire w_dff_B_NAGmiFYT7_2;
	wire w_dff_B_taqlKBRo7_2;
	wire w_dff_B_brYJ81LH6_2;
	wire w_dff_B_lNswk0dg6_2;
	wire w_dff_B_NoOfWuhP6_2;
	wire w_dff_B_uVj7vMka2_2;
	wire w_dff_B_FHDfKqcc2_1;
	wire w_dff_B_fUk4hqjq2_2;
	wire w_dff_B_NMJW5qQQ6_2;
	wire w_dff_B_p0VVpxOD7_2;
	wire w_dff_B_fcmW6xwU6_2;
	wire w_dff_B_guLnpw2S4_2;
	wire w_dff_B_Z7m1PGz53_2;
	wire w_dff_B_9pL1rP5c5_2;
	wire w_dff_B_2iH3l9Ps9_2;
	wire w_dff_B_rcPjiLWS1_2;
	wire w_dff_B_qFMZlzBN6_2;
	wire w_dff_B_p96wqOZf1_0;
	wire w_dff_A_hn2ihA4X7_0;
	wire w_dff_A_uRE18QYz7_0;
	wire w_dff_A_9DHjInrX5_0;
	wire w_dff_A_VnVkTe6E1_0;
	wire w_dff_B_QzRqY8Wk5_1;
	wire w_dff_B_EkBsbp5C6_2;
	wire w_dff_B_V9gy66MR8_2;
	wire w_dff_B_yvxOb0tX3_2;
	wire w_dff_B_0htVR8JQ3_2;
	wire w_dff_B_kgx9rspv3_2;
	wire w_dff_B_wW5J3Qoh9_2;
	wire w_dff_B_soxLtRFc3_2;
	wire w_dff_B_FWVnXE4p0_2;
	wire w_dff_B_WzvgQYNR4_2;
	wire w_dff_B_mAyzAEGv6_2;
	wire w_dff_B_5kND4eji3_2;
	wire w_dff_B_DbAaB1HS5_2;
	wire w_dff_B_e4KXCDof2_2;
	wire w_dff_B_49mKgtxF0_2;
	wire w_dff_B_9CdU1SOe2_2;
	wire w_dff_B_5hYqEvx10_2;
	wire w_dff_B_pvutrAiR3_2;
	wire w_dff_B_AqLBlfe52_2;
	wire w_dff_B_2GA041mq3_2;
	wire w_dff_B_C2zU20Io9_2;
	wire w_dff_B_rU33edgr0_2;
	wire w_dff_B_OjLXyaVm5_2;
	wire w_dff_B_81I1jSqI7_2;
	wire w_dff_B_U93Whbfi2_2;
	wire w_dff_B_OyWiSILw4_2;
	wire w_dff_B_4PLsqf2P9_2;
	wire w_dff_B_YFt1gIIa4_2;
	wire w_dff_B_v7PNWjxa0_2;
	wire w_dff_B_z7Ry1QkT6_2;
	wire w_dff_B_cDt5Zpe71_2;
	wire w_dff_B_OoEpJWQ75_2;
	wire w_dff_B_qZ5tv5vY1_2;
	wire w_dff_B_kwTMnRty0_2;
	wire w_dff_B_1Xdjdf6N3_2;
	wire w_dff_B_Pmgh6Obo0_2;
	wire w_dff_B_AnrDfWcl1_2;
	wire w_dff_B_cROquOB40_2;
	wire w_dff_B_8iPXoG4N2_2;
	wire w_dff_B_dFmAg3GA4_2;
	wire w_dff_B_MBQbCFaM1_2;
	wire w_dff_B_r03NUlUN3_2;
	wire w_dff_B_XQyldepu8_2;
	wire w_dff_B_ihKtn3974_2;
	wire w_dff_B_lMmJApGb6_2;
	wire w_dff_B_qZbCVfzj9_0;
	wire w_dff_A_KSJU7kjs1_1;
	wire w_dff_B_PIGqr8be1_1;
	wire w_dff_B_Ty8a6ple1_2;
	wire w_dff_B_TgjVLXRI8_2;
	wire w_dff_B_iX1SIyCK9_2;
	wire w_dff_B_Bpbbljzn2_2;
	wire w_dff_B_BWbAjSqr9_2;
	wire w_dff_B_QiCnsXfR8_2;
	wire w_dff_B_ndOyVV2j6_2;
	wire w_dff_B_61lASTgb5_2;
	wire w_dff_B_5DdOldDp4_2;
	wire w_dff_B_MW2rohRv5_2;
	wire w_dff_B_vw7WS6Vh2_2;
	wire w_dff_B_O72Qgpf74_2;
	wire w_dff_B_y1TaDchZ3_2;
	wire w_dff_B_tUTWzf819_2;
	wire w_dff_B_YFiYT1dE0_2;
	wire w_dff_B_zvHLBJFV5_2;
	wire w_dff_B_2Mx7iK5f4_2;
	wire w_dff_B_bRBWLhek8_2;
	wire w_dff_B_otkSlVI13_2;
	wire w_dff_B_ENapcN2Q7_2;
	wire w_dff_B_wznB5eDK4_2;
	wire w_dff_B_3GKlaIZe6_2;
	wire w_dff_B_uoHfKMwe3_2;
	wire w_dff_B_QUFRqTmT9_2;
	wire w_dff_B_DtG11sPz5_2;
	wire w_dff_B_XgtGxpl03_2;
	wire w_dff_B_1vmPD2DE7_2;
	wire w_dff_B_YZQ42WSY0_2;
	wire w_dff_B_KYsVBEqh2_2;
	wire w_dff_B_sQAQDt9x0_2;
	wire w_dff_B_oyWSxQ8s7_2;
	wire w_dff_B_VVkazXL08_2;
	wire w_dff_B_p14iwy2s5_2;
	wire w_dff_B_nWvH51cH1_2;
	wire w_dff_B_mXrTqje64_2;
	wire w_dff_B_mMzPzBnB3_2;
	wire w_dff_B_pDd7DsGf2_2;
	wire w_dff_B_7UA23h9k2_2;
	wire w_dff_B_b70qJSYz4_2;
	wire w_dff_B_5iKIACOp3_2;
	wire w_dff_B_sd11iQz02_1;
	wire w_dff_B_hEbWQPmX7_2;
	wire w_dff_B_iSAHyJDU1_2;
	wire w_dff_B_fWquE1lm3_2;
	wire w_dff_B_IXoj6phy2_2;
	wire w_dff_B_F6nurJeV8_2;
	wire w_dff_B_6BhQ51V03_2;
	wire w_dff_B_bCwoT1087_2;
	wire w_dff_B_63redlre2_2;
	wire w_dff_B_KhVip9yp2_2;
	wire w_dff_B_9eFEpYFy0_2;
	wire w_dff_B_IiLtqin01_2;
	wire w_dff_B_p2cgsK5s6_2;
	wire w_dff_B_of7gZplG1_2;
	wire w_dff_B_bs3hwhOS7_2;
	wire w_dff_B_eduZAaEZ4_2;
	wire w_dff_B_S0g0nGY06_2;
	wire w_dff_B_3MpBENIv7_2;
	wire w_dff_B_wtFYxcyM4_2;
	wire w_dff_B_AV4j1lCr9_2;
	wire w_dff_B_ppbbj4CA7_2;
	wire w_dff_B_CgPF2nQd7_2;
	wire w_dff_B_zHiCCIu05_2;
	wire w_dff_B_LfNVZFHD4_2;
	wire w_dff_B_3PL62WaT2_2;
	wire w_dff_B_ZSbUGnJW2_2;
	wire w_dff_B_pWWTM2Y27_2;
	wire w_dff_B_Al4mrGMr3_2;
	wire w_dff_B_6nyFcD707_2;
	wire w_dff_B_hcK1CvGR3_2;
	wire w_dff_B_EzUzla1W5_2;
	wire w_dff_B_FmlE7YQ12_2;
	wire w_dff_B_zAg5CuoL4_2;
	wire w_dff_B_cHCEvE6K0_2;
	wire w_dff_B_hiXhoUJe8_2;
	wire w_dff_B_GAIlJRWL5_2;
	wire w_dff_B_yxORPfpV4_2;
	wire w_dff_B_kFtO13Jo8_2;
	wire w_dff_B_h5RKjoXL7_1;
	wire w_dff_B_NnjAGsoU7_2;
	wire w_dff_B_LYVkxd7D5_2;
	wire w_dff_B_VmWTAZtv4_2;
	wire w_dff_B_tnMALOZq3_2;
	wire w_dff_B_d7bR3JMp8_2;
	wire w_dff_B_ruUHm3AQ6_2;
	wire w_dff_B_TC4EuuNo9_2;
	wire w_dff_B_yM2L6Mdt9_2;
	wire w_dff_B_0IPI0RnW8_2;
	wire w_dff_B_Q3q1zVDc1_2;
	wire w_dff_B_bI9xB2bZ9_2;
	wire w_dff_B_TjPZ7ovH1_2;
	wire w_dff_B_Lm9FGTjR5_2;
	wire w_dff_B_tZNQvoH75_2;
	wire w_dff_B_4pJm1sHH8_2;
	wire w_dff_B_H4pbYAZF2_2;
	wire w_dff_B_sVdGHBeJ4_2;
	wire w_dff_B_so5KxBVc1_2;
	wire w_dff_B_OLx5nN6y6_2;
	wire w_dff_B_A6cRI4CC0_2;
	wire w_dff_B_H5aKrbt48_2;
	wire w_dff_B_tQKB44Qv3_2;
	wire w_dff_B_cFMP2liM2_2;
	wire w_dff_B_mAIyepEz8_2;
	wire w_dff_B_kTr9xOqP9_2;
	wire w_dff_B_vCH8Yl6s0_2;
	wire w_dff_B_zXluw1Pn2_2;
	wire w_dff_B_9colIbKg8_2;
	wire w_dff_B_ZAZGKhV92_2;
	wire w_dff_B_cPn2rPyx0_2;
	wire w_dff_B_cn1O666u4_2;
	wire w_dff_B_41p4QyuJ8_2;
	wire w_dff_B_uKmEUj662_2;
	wire w_dff_B_ZU10pe9H4_2;
	wire w_dff_B_btAzBAx92_1;
	wire w_dff_B_VfH5eDLA1_2;
	wire w_dff_B_oaqYiaht3_2;
	wire w_dff_B_0yXjSoOC4_2;
	wire w_dff_B_0M9xiurG3_2;
	wire w_dff_B_NHpPM4v32_2;
	wire w_dff_B_tOnSlKTU0_2;
	wire w_dff_B_2ODDkCKI1_2;
	wire w_dff_B_joaL3qXE0_2;
	wire w_dff_B_CLQvEiQE2_2;
	wire w_dff_B_jDHRomNs2_2;
	wire w_dff_B_gUogtGF26_2;
	wire w_dff_B_OQVanudn7_2;
	wire w_dff_B_6SX5KmRQ8_2;
	wire w_dff_B_yzV2Or5e4_2;
	wire w_dff_B_tvV6kvBu0_2;
	wire w_dff_B_5K8zSqgW8_2;
	wire w_dff_B_kxCncmAs0_2;
	wire w_dff_B_Ag3YV6zH0_2;
	wire w_dff_B_PlsJUzfM3_2;
	wire w_dff_B_l2dIo4kx2_2;
	wire w_dff_B_U0akR9E61_2;
	wire w_dff_B_NNCM58xX8_2;
	wire w_dff_B_oixyRztc2_2;
	wire w_dff_B_OXM9SkIO4_2;
	wire w_dff_B_oC5ZLoHu2_2;
	wire w_dff_B_mOPvEqd12_2;
	wire w_dff_B_zUZlpJFU2_2;
	wire w_dff_B_5ICvawnu0_2;
	wire w_dff_B_aBYRBPMW7_2;
	wire w_dff_B_l0x3636S9_2;
	wire w_dff_B_8D3wYtpI7_2;
	wire w_dff_B_njc17Ywt8_1;
	wire w_dff_B_6cC8yWm12_2;
	wire w_dff_B_plZlpx0s6_2;
	wire w_dff_B_xb8gVmEt6_2;
	wire w_dff_B_w5Xido9G2_2;
	wire w_dff_B_HOPuzNZf5_2;
	wire w_dff_B_Qvz7TyA18_2;
	wire w_dff_B_wuIZJW1W9_2;
	wire w_dff_B_bvELdRvx3_2;
	wire w_dff_B_ceOTJzh47_2;
	wire w_dff_B_TKpfZjDq6_2;
	wire w_dff_B_WuACwFQS9_2;
	wire w_dff_B_tx0XA0783_2;
	wire w_dff_B_NWz40CIk0_2;
	wire w_dff_B_vIFXtAW55_2;
	wire w_dff_B_bzFWu4ny1_2;
	wire w_dff_B_75wCUuzk0_2;
	wire w_dff_B_tfdl6AfL5_2;
	wire w_dff_B_YZpG7Fea5_2;
	wire w_dff_B_LaH0a9xn0_2;
	wire w_dff_B_UJ4MCAKo1_2;
	wire w_dff_B_fOYjXp3i4_2;
	wire w_dff_B_vJoXqYFp8_2;
	wire w_dff_B_g2y8LwN22_2;
	wire w_dff_B_i2MIQDRW4_2;
	wire w_dff_B_NIJGMWC59_2;
	wire w_dff_B_51UgwMD87_2;
	wire w_dff_B_uISdzOLI9_2;
	wire w_dff_B_xUzkRPVC2_2;
	wire w_dff_B_xlYWbEmV9_1;
	wire w_dff_B_pt8vCAy86_2;
	wire w_dff_B_s5txgLny6_2;
	wire w_dff_B_t4oyNgGK6_2;
	wire w_dff_B_yTAOYG8R6_2;
	wire w_dff_B_qt64Ig8W3_2;
	wire w_dff_B_2Eme1FDV3_2;
	wire w_dff_B_6tjTP7AH4_2;
	wire w_dff_B_9RCxY58A2_2;
	wire w_dff_B_aTQZ94k94_2;
	wire w_dff_B_sJyoePeo2_2;
	wire w_dff_B_ImeqOoTv9_2;
	wire w_dff_B_1Itl3AOh3_2;
	wire w_dff_B_mZbG4vqC8_2;
	wire w_dff_B_rSfylnvx7_2;
	wire w_dff_B_m61EIGg49_2;
	wire w_dff_B_MqoDtEPs3_2;
	wire w_dff_B_2MiqQLhx2_2;
	wire w_dff_B_1Gyz0rPC4_2;
	wire w_dff_B_FiWusDru0_2;
	wire w_dff_B_slO8bQ4h7_2;
	wire w_dff_B_7A5LtFVb7_2;
	wire w_dff_B_rKjJMvQ06_2;
	wire w_dff_B_hZEEUm4Y3_2;
	wire w_dff_B_5DMS3Dqa4_2;
	wire w_dff_B_cHYOWHXB5_2;
	wire w_dff_B_zA1fVh209_1;
	wire w_dff_B_1TX4ygRy1_2;
	wire w_dff_B_2Ap0Oqjh9_2;
	wire w_dff_B_fy72smUI6_2;
	wire w_dff_B_v6yxoG7W3_2;
	wire w_dff_B_9xjHvdEt9_2;
	wire w_dff_B_Pcfv2wn50_2;
	wire w_dff_B_XPrzWFuJ1_2;
	wire w_dff_B_jWl5kXsp0_2;
	wire w_dff_B_dgaqfbzw1_2;
	wire w_dff_B_moLpdjUd3_2;
	wire w_dff_B_yKpLB11R7_2;
	wire w_dff_B_Lcg9y8Rs8_2;
	wire w_dff_B_dYU88pkw3_2;
	wire w_dff_B_jAOlGQVv3_2;
	wire w_dff_B_anPlZ8127_2;
	wire w_dff_B_GHpfCaqR4_2;
	wire w_dff_B_RLwUrAon2_2;
	wire w_dff_B_stLmgViI4_2;
	wire w_dff_B_N3kdYXo48_2;
	wire w_dff_B_MgyIN9sG8_2;
	wire w_dff_B_EPOCiutL4_2;
	wire w_dff_B_EnMmaieR2_2;
	wire w_dff_B_5tQ7JrXv8_1;
	wire w_dff_B_unxCXfma1_2;
	wire w_dff_B_DP6qr3E65_2;
	wire w_dff_B_8WCx9P2a0_2;
	wire w_dff_B_s9KaS7nA7_2;
	wire w_dff_B_Qk2RJZfU0_2;
	wire w_dff_B_HucCc95M5_2;
	wire w_dff_B_aEXFm0rz2_2;
	wire w_dff_B_8bl8lquq5_2;
	wire w_dff_B_Yhzy4Ndu3_2;
	wire w_dff_B_njnJNp6A2_2;
	wire w_dff_B_cS8zJBEm8_2;
	wire w_dff_B_5CUOBbrJ7_2;
	wire w_dff_B_HqXxARjb4_2;
	wire w_dff_B_xOSps5fC8_2;
	wire w_dff_B_iZ8ykPvT0_2;
	wire w_dff_B_2ZKYKSsb9_2;
	wire w_dff_B_tsuREzKB2_2;
	wire w_dff_B_4CxapzYz1_2;
	wire w_dff_B_4qBsAPLP7_2;
	wire w_dff_B_OJBqW99N0_1;
	wire w_dff_B_8TiqfJm83_2;
	wire w_dff_B_spq7FsAY6_2;
	wire w_dff_B_iU8hxj5e1_2;
	wire w_dff_B_PoU6hK8L2_2;
	wire w_dff_B_YEs4TTuI8_2;
	wire w_dff_B_aKduiEst8_2;
	wire w_dff_B_4qvfDN7q2_2;
	wire w_dff_B_8hgihRAU9_2;
	wire w_dff_B_1GD3gS9O6_2;
	wire w_dff_B_EOP7VZoZ8_2;
	wire w_dff_B_lovxccja4_2;
	wire w_dff_B_itFyY2Vu1_2;
	wire w_dff_B_gQntoKex1_2;
	wire w_dff_B_9hBpI5fz1_2;
	wire w_dff_B_BS4fxE5g2_2;
	wire w_dff_B_r0V17XPo8_2;
	wire w_dff_B_SU23IKnx1_1;
	wire w_dff_B_Qg4SlNPd6_2;
	wire w_dff_B_mZfea7FP3_2;
	wire w_dff_B_Cq93G2qv7_2;
	wire w_dff_B_kpgUEfDk0_2;
	wire w_dff_B_Kfx9Yzom1_2;
	wire w_dff_B_FE3Gv6zn0_2;
	wire w_dff_B_zx2YoD5R1_2;
	wire w_dff_B_DxyAWonr9_2;
	wire w_dff_B_elgOHi1A7_2;
	wire w_dff_B_Hm7V5PC60_2;
	wire w_dff_B_cbYwfaWm6_2;
	wire w_dff_B_aXqrKbzR6_2;
	wire w_dff_B_wdsUzH4j4_2;
	wire w_dff_B_7jaHZNBo7_1;
	wire w_dff_B_7DToSdmf9_2;
	wire w_dff_B_M4yhwTvW1_2;
	wire w_dff_B_lcqc8b7C2_2;
	wire w_dff_B_epfj3P5X7_2;
	wire w_dff_B_MansYrIu4_2;
	wire w_dff_B_EQiZtGhV6_2;
	wire w_dff_B_AdXqyWo67_2;
	wire w_dff_B_JKAZmDuY8_2;
	wire w_dff_B_vjmx9RdH1_2;
	wire w_dff_B_waBKwR1N6_2;
	wire w_dff_B_bwQLdsF85_1;
	wire w_dff_B_rWS67cWL3_2;
	wire w_dff_B_eJtv3WUt9_2;
	wire w_dff_B_cYqClYIx4_2;
	wire w_dff_B_CV3Uu8y61_2;
	wire w_dff_B_atcqW1Xi4_2;
	wire w_dff_B_MLy6fGzE4_2;
	wire w_dff_B_NTfgZDis7_2;
	wire w_dff_B_pD4IhY2h2_2;
	wire w_dff_B_vgbS1Rp80_2;
	wire w_dff_B_cj34X8qx6_2;
	wire w_dff_B_Bo96JeWH4_0;
	wire w_dff_A_9FnJfSj86_0;
	wire w_dff_A_0Gfv49f07_0;
	wire w_dff_A_bfPU2Rw02_0;
	wire w_dff_A_NFpSeRGc1_0;
	wire w_dff_B_82kEDmpO3_2;
	wire w_dff_B_p8CFYD8r0_1;
	wire w_dff_B_HI0qfoCK6_2;
	wire w_dff_B_w73QtY3Q9_2;
	wire w_dff_B_LNYBxVAH7_2;
	wire w_dff_B_lPzsAtnl1_2;
	wire w_dff_B_i6rbg7Gh2_2;
	wire w_dff_B_H2vf3QHQ9_2;
	wire w_dff_B_644zwNW39_2;
	wire w_dff_B_AUHmEi0s6_2;
	wire w_dff_B_0XDnDoZu7_2;
	wire w_dff_B_GWh1cxgr8_2;
	wire w_dff_B_Mc1DBr5L5_2;
	wire w_dff_B_OaBZf7ZE6_2;
	wire w_dff_B_58AJcBXl5_2;
	wire w_dff_B_5tmlsUO70_2;
	wire w_dff_B_Tmk9yV9w1_2;
	wire w_dff_B_WdOXA5mO3_2;
	wire w_dff_B_Zs0lAgYe5_2;
	wire w_dff_B_ZBSGuona0_2;
	wire w_dff_B_DSnE9pEi0_2;
	wire w_dff_B_N3MGM5NK5_2;
	wire w_dff_B_0QJHOML52_2;
	wire w_dff_B_DAQtcvhJ1_2;
	wire w_dff_B_JhCNHU203_2;
	wire w_dff_B_iPkvAayr1_2;
	wire w_dff_B_yIxlhDMw1_2;
	wire w_dff_B_ANWPsLnT1_2;
	wire w_dff_B_8OEexEgb5_2;
	wire w_dff_B_PX4UNlqr5_2;
	wire w_dff_B_oa0pRPl03_2;
	wire w_dff_B_FibqFtvc0_2;
	wire w_dff_B_zzVScD3D7_2;
	wire w_dff_B_luxOHkko4_2;
	wire w_dff_B_yfR7hewW4_2;
	wire w_dff_B_jRtBBDC25_2;
	wire w_dff_B_WxJYm7pB9_2;
	wire w_dff_B_uMKWbvTc7_2;
	wire w_dff_B_CvaJ2SY51_2;
	wire w_dff_B_FmLZ3YRa6_2;
	wire w_dff_B_obwItojH0_2;
	wire w_dff_B_bC6drbKZ5_2;
	wire w_dff_B_2xx4hGKK8_2;
	wire w_dff_B_78y7PVT11_2;
	wire w_dff_B_SmH6ODnO9_2;
	wire w_dff_B_RRUhEdFG0_2;
	wire w_dff_B_8gNLrgrL5_1;
	wire w_dff_B_EGvTs1xQ9_2;
	wire w_dff_B_vmsMTtn00_2;
	wire w_dff_B_Zzdhxzqe1_2;
	wire w_dff_B_r0mzhX8g9_2;
	wire w_dff_B_ABwxiugB5_2;
	wire w_dff_B_QmTSpFZp3_2;
	wire w_dff_B_FWRpa9tG3_2;
	wire w_dff_B_CuoKJ7Sx5_2;
	wire w_dff_B_WowdH8jj9_2;
	wire w_dff_B_fSLnroM98_2;
	wire w_dff_B_SDYmAZBe9_2;
	wire w_dff_B_CnjXIl4S1_2;
	wire w_dff_B_RTL4yCjC8_2;
	wire w_dff_B_YEiyUClY1_2;
	wire w_dff_B_M6m0kAGz4_2;
	wire w_dff_B_RNWrOxw22_2;
	wire w_dff_B_VZj7Jbbp9_2;
	wire w_dff_B_gL287Ds75_2;
	wire w_dff_B_noyylPMX4_2;
	wire w_dff_B_GUT3ncYz4_2;
	wire w_dff_B_Qye8awiK7_2;
	wire w_dff_B_O7kn2KFC2_2;
	wire w_dff_B_xaYz8JMU4_2;
	wire w_dff_B_QzuES2Gt2_2;
	wire w_dff_B_frUWt0if3_2;
	wire w_dff_B_gPjMMraJ6_2;
	wire w_dff_B_rQAbOnRM8_2;
	wire w_dff_B_iTUhyJ955_2;
	wire w_dff_B_gO1OiREC7_2;
	wire w_dff_B_GI2S4c4N1_2;
	wire w_dff_B_PbHefd6e7_2;
	wire w_dff_B_20oLcZmG6_2;
	wire w_dff_B_xMYI3rRT2_2;
	wire w_dff_B_CSBp4CcL0_2;
	wire w_dff_B_k0b7nD5x0_2;
	wire w_dff_B_odrsetPv7_2;
	wire w_dff_B_CWleIVRD5_2;
	wire w_dff_B_ZrBCp82e3_2;
	wire w_dff_B_kISjt9Nd0_2;
	wire w_dff_B_6d1qojQz1_1;
	wire w_dff_B_arPmkPW94_2;
	wire w_dff_B_eYb4nYSB6_2;
	wire w_dff_B_UA0qZu8p6_2;
	wire w_dff_B_ycShQNNf1_2;
	wire w_dff_B_vwywIjc38_2;
	wire w_dff_B_at1gFTkX8_2;
	wire w_dff_B_cmhlqIXG9_2;
	wire w_dff_B_pISZsA3N8_2;
	wire w_dff_B_mMikUdx37_2;
	wire w_dff_B_QLYrlFXX6_2;
	wire w_dff_B_jHcBvwUM4_2;
	wire w_dff_B_1QeLrvrj9_2;
	wire w_dff_B_y537y5px3_2;
	wire w_dff_B_7EOGJAyi0_2;
	wire w_dff_B_SRZiTzNW4_2;
	wire w_dff_B_BBsEUafp8_2;
	wire w_dff_B_SuLWa2X11_2;
	wire w_dff_B_N1fq99Ep3_2;
	wire w_dff_B_LbBO6qaN2_2;
	wire w_dff_B_TyOotS5b3_2;
	wire w_dff_B_sG5fA6rP3_2;
	wire w_dff_B_9Mr5x8V88_2;
	wire w_dff_B_5rC9Sz629_2;
	wire w_dff_B_2XOD3RCs5_2;
	wire w_dff_B_iUV9ddRP3_2;
	wire w_dff_B_lmhbLABn6_2;
	wire w_dff_B_gd9OMT3T3_2;
	wire w_dff_B_LDYzMncT7_2;
	wire w_dff_B_kP9rWVYB7_2;
	wire w_dff_B_0lC176QA7_2;
	wire w_dff_B_hQAH83qA2_2;
	wire w_dff_B_kq3TksPn3_2;
	wire w_dff_B_9RGTEren2_2;
	wire w_dff_B_eo8HzTsY9_2;
	wire w_dff_B_vCCULbSY1_2;
	wire w_dff_B_K4Sn2Y1Z6_2;
	wire w_dff_B_LiVhcqFl1_1;
	wire w_dff_B_5T1BUQmj0_2;
	wire w_dff_B_6hDLsMDT8_2;
	wire w_dff_B_sA8hbA520_2;
	wire w_dff_B_THETvd4u5_2;
	wire w_dff_B_VxDt8xz84_2;
	wire w_dff_B_xFbP1kHF3_2;
	wire w_dff_B_silobUlP7_2;
	wire w_dff_B_0jBhBDnc6_2;
	wire w_dff_B_04O1bZi03_2;
	wire w_dff_B_t02yxgQk1_2;
	wire w_dff_B_MewjG7D89_2;
	wire w_dff_B_dFCn7i5V6_2;
	wire w_dff_B_aVcUdzfJ1_2;
	wire w_dff_B_5CNxMRfU1_2;
	wire w_dff_B_cFdAtfq98_2;
	wire w_dff_B_CqDelUtY8_2;
	wire w_dff_B_HN26A4Ni0_2;
	wire w_dff_B_ESmp7wAC2_2;
	wire w_dff_B_6SQQFuWk0_2;
	wire w_dff_B_ZdHZhSpi1_2;
	wire w_dff_B_ydtLEszk5_2;
	wire w_dff_B_yJlNFCTq1_2;
	wire w_dff_B_T9STk5IL3_2;
	wire w_dff_B_jr5fRvJ45_2;
	wire w_dff_B_EdQo7zSe0_2;
	wire w_dff_B_GCfu9r2u5_2;
	wire w_dff_B_GbPeGblU3_2;
	wire w_dff_B_ETSuWgpd3_2;
	wire w_dff_B_BBvFPJw66_2;
	wire w_dff_B_ZkoKZYV51_2;
	wire w_dff_B_Tv3gA1nG5_2;
	wire w_dff_B_ExnYwyxT1_2;
	wire w_dff_B_bJ48C7vN1_2;
	wire w_dff_B_TOvxfCyx5_1;
	wire w_dff_B_OOBUTOR80_2;
	wire w_dff_B_D8hCKFkA6_2;
	wire w_dff_B_b1EnRnaB3_2;
	wire w_dff_B_BXIPDdgF9_2;
	wire w_dff_B_v2VkihFM1_2;
	wire w_dff_B_AVv2Zxrm7_2;
	wire w_dff_B_MH4fLmfQ2_2;
	wire w_dff_B_fPbrqTmk8_2;
	wire w_dff_B_jT1SUDCg2_2;
	wire w_dff_B_WKMyKDQw5_2;
	wire w_dff_B_mJQtkapL5_2;
	wire w_dff_B_1MfXvMZP2_2;
	wire w_dff_B_9DHT5X8f3_2;
	wire w_dff_B_351IfMQB1_2;
	wire w_dff_B_y4NHOxFn7_2;
	wire w_dff_B_YPCthopJ1_2;
	wire w_dff_B_4awknyCS9_2;
	wire w_dff_B_DWLC9RBZ3_2;
	wire w_dff_B_OqWSA1Nw7_2;
	wire w_dff_B_gCtn49xw4_2;
	wire w_dff_B_Pi0nXxgR0_2;
	wire w_dff_B_8AZnS9pP3_2;
	wire w_dff_B_Xxba8x8E1_2;
	wire w_dff_B_Ehs56RKh6_2;
	wire w_dff_B_HD4A2ZOK1_2;
	wire w_dff_B_tGNUhpZH2_2;
	wire w_dff_B_pfjyruZ24_2;
	wire w_dff_B_JbvP0yVV6_2;
	wire w_dff_B_Ob6Fd71d9_2;
	wire w_dff_B_pOWat9C22_2;
	wire w_dff_B_3pE5dkfD9_1;
	wire w_dff_B_Sdv33Ges1_2;
	wire w_dff_B_aGtrsy8H2_2;
	wire w_dff_B_gwpL6CsZ7_2;
	wire w_dff_B_JJvg7gsc7_2;
	wire w_dff_B_gFquDKE14_2;
	wire w_dff_B_IHxtHSjZ1_2;
	wire w_dff_B_SP6uV0Fr4_2;
	wire w_dff_B_EUc7JVss8_2;
	wire w_dff_B_Gq3OZvl68_2;
	wire w_dff_B_OlSijAxY2_2;
	wire w_dff_B_mvxnN1Jh5_2;
	wire w_dff_B_7WigKAb76_2;
	wire w_dff_B_mOah6vMx6_2;
	wire w_dff_B_bv47knXu4_2;
	wire w_dff_B_tujRlVA13_2;
	wire w_dff_B_ZTTkuLQJ6_2;
	wire w_dff_B_EJc5b1yF0_2;
	wire w_dff_B_ksKWp9c14_2;
	wire w_dff_B_SERcjpHn4_2;
	wire w_dff_B_tvqRN6p74_2;
	wire w_dff_B_QfL4rNG06_2;
	wire w_dff_B_CZvNo3Yr6_2;
	wire w_dff_B_ucpVJGBH3_2;
	wire w_dff_B_toF0Zfpz7_2;
	wire w_dff_B_28ZkR1Dl2_2;
	wire w_dff_B_nS4ZgaTO2_2;
	wire w_dff_B_oweQ0Jal5_2;
	wire w_dff_B_R0z19Jep3_1;
	wire w_dff_B_QXRnl56v5_2;
	wire w_dff_B_v8ZdHMr87_2;
	wire w_dff_B_V1zqU0I55_2;
	wire w_dff_B_CisTQMR80_2;
	wire w_dff_B_fe4cb1eZ6_2;
	wire w_dff_B_ijIuYNse6_2;
	wire w_dff_B_566cVKcr4_2;
	wire w_dff_B_WqcfleWR4_2;
	wire w_dff_B_S3eKu4XR9_2;
	wire w_dff_B_pQ4tXXlM0_2;
	wire w_dff_B_VWJBY6Ak9_2;
	wire w_dff_B_144ktcIl9_2;
	wire w_dff_B_rTcU2Qbc6_2;
	wire w_dff_B_5txrRGBZ7_2;
	wire w_dff_B_ceTNVhgU7_2;
	wire w_dff_B_oM1CwD9C8_2;
	wire w_dff_B_FCiStozC3_2;
	wire w_dff_B_uCabLax15_2;
	wire w_dff_B_MMFxZGqu2_2;
	wire w_dff_B_ptfX8f457_2;
	wire w_dff_B_Cnn5jTTL5_2;
	wire w_dff_B_2ydK2cuO5_2;
	wire w_dff_B_ZUEycug21_2;
	wire w_dff_B_QgQgfMTD9_2;
	wire w_dff_B_y8GhzqHs6_1;
	wire w_dff_B_wKUwr2961_2;
	wire w_dff_B_cAHx3hjm3_2;
	wire w_dff_B_hZNCI5Hf4_2;
	wire w_dff_B_sP1w03i44_2;
	wire w_dff_B_9iWZnr7B6_2;
	wire w_dff_B_knllvzOm7_2;
	wire w_dff_B_8Ck0rVff5_2;
	wire w_dff_B_9gBWMI4B5_2;
	wire w_dff_B_rgx9td3J4_2;
	wire w_dff_B_WQ171XwV0_2;
	wire w_dff_B_dwY2m9UF3_2;
	wire w_dff_B_JUxIufPX6_2;
	wire w_dff_B_PV8T9nrb8_2;
	wire w_dff_B_5h6mvSNl8_2;
	wire w_dff_B_Ojy9qFaM2_2;
	wire w_dff_B_dol2pIu93_2;
	wire w_dff_B_FRJtNm0V9_2;
	wire w_dff_B_YOq2of3r1_2;
	wire w_dff_B_IyBLy1eD9_2;
	wire w_dff_B_jQaiMMzj2_2;
	wire w_dff_B_N8U5UmxG3_2;
	wire w_dff_B_tzp9z56e2_1;
	wire w_dff_B_jPNCXNaj2_2;
	wire w_dff_B_Cpi0dReh1_2;
	wire w_dff_B_OWU55v149_2;
	wire w_dff_B_wvPkt51q9_2;
	wire w_dff_B_3juSFDU49_2;
	wire w_dff_B_Lrkf98dy0_2;
	wire w_dff_B_yl3iKIQG4_2;
	wire w_dff_B_yZdKaMai2_2;
	wire w_dff_B_DLeQDyfQ9_2;
	wire w_dff_B_2bPKmKWU6_2;
	wire w_dff_B_GcPNPhsu4_2;
	wire w_dff_B_rndqwl6u4_2;
	wire w_dff_B_DknIx0LD7_2;
	wire w_dff_B_t4DhqEG94_2;
	wire w_dff_B_Td7YVL914_2;
	wire w_dff_B_mlVKHcth2_2;
	wire w_dff_B_GZaXYlnM9_2;
	wire w_dff_B_ImxTX2uV5_2;
	wire w_dff_B_yLerp6T52_1;
	wire w_dff_B_xh23TJQr8_2;
	wire w_dff_B_09jGHuYQ8_2;
	wire w_dff_B_6ejMo3wB8_2;
	wire w_dff_B_c5X5DqdK8_2;
	wire w_dff_B_HGtgy4R34_2;
	wire w_dff_B_yCSnzhs16_2;
	wire w_dff_B_SFvSsLEM0_2;
	wire w_dff_B_1jqv8wRl7_2;
	wire w_dff_B_dBRo2nOc2_2;
	wire w_dff_B_ZzuDrKUA1_2;
	wire w_dff_B_fd8RLpn81_2;
	wire w_dff_B_HZl9l0B42_2;
	wire w_dff_B_TcTb2V1f6_2;
	wire w_dff_B_8kyQZQZ51_2;
	wire w_dff_B_JfRbc5xr0_2;
	wire w_dff_B_AwApN28D3_1;
	wire w_dff_B_ui3Vok8d8_2;
	wire w_dff_B_rycLXFoe9_2;
	wire w_dff_B_BAIFFObf8_2;
	wire w_dff_B_i6dKyt5G1_2;
	wire w_dff_B_zAncI7QG6_2;
	wire w_dff_B_duj50ZVH5_2;
	wire w_dff_B_5QHiVTBT2_2;
	wire w_dff_B_Eli7zVJp5_2;
	wire w_dff_B_HuYzGv3G8_2;
	wire w_dff_B_vM8hH5fA0_2;
	wire w_dff_B_2wEY9y9G1_2;
	wire w_dff_B_4Ews6Nh30_2;
	wire w_dff_B_NBaNDCuu2_1;
	wire w_dff_B_em16gT3f0_2;
	wire w_dff_B_UhREfVy77_2;
	wire w_dff_B_ZGV8XdVu4_2;
	wire w_dff_B_FiMxoM3v3_2;
	wire w_dff_B_NhkCPPxv1_2;
	wire w_dff_B_oWJ8I7fA0_2;
	wire w_dff_B_U5HSUCU58_2;
	wire w_dff_B_RIt4nk6Q7_2;
	wire w_dff_B_bhrnvtsu1_2;
	wire w_dff_B_AZjjbSdA3_2;
	wire w_dff_B_vTLeOGiF5_1;
	wire w_dff_B_96ZCAOpF3_2;
	wire w_dff_B_yrshsnC17_2;
	wire w_dff_B_9AaqN74H3_2;
	wire w_dff_B_Tn8aBqFA4_2;
	wire w_dff_B_w4EXgv7l6_2;
	wire w_dff_B_uIrpoRSt3_2;
	wire w_dff_B_008ENNDH2_2;
	wire w_dff_B_9mLinlEm2_2;
	wire w_dff_B_lGbCP0C67_2;
	wire w_dff_B_lTV9VUfa5_2;
	wire w_dff_B_GV8eUhdT1_0;
	wire w_dff_A_GLXUj7kV6_0;
	wire w_dff_A_PJAIXXDw9_0;
	wire w_dff_A_yrorCRtU1_1;
	wire w_dff_A_q9M9gnBA4_1;
	wire w_dff_B_w8ZEJdi97_2;
	wire w_dff_B_3QFD0j615_1;
	wire w_dff_B_k2wqKZQZ9_2;
	wire w_dff_B_SQ3Agozi2_2;
	wire w_dff_B_Ub5cjh3i8_2;
	wire w_dff_B_5c4vqkeX8_2;
	wire w_dff_B_3Nuek61q6_2;
	wire w_dff_B_sfNeiznr8_2;
	wire w_dff_B_Mp7ndH4q8_2;
	wire w_dff_B_ArSjtfMa1_2;
	wire w_dff_B_wnb6lGO95_2;
	wire w_dff_B_x3L7vdKr0_2;
	wire w_dff_B_3pbMwHA09_2;
	wire w_dff_B_CnP5aY734_2;
	wire w_dff_B_StkDG3hZ3_2;
	wire w_dff_B_eybkSGqS9_2;
	wire w_dff_B_AqZy4FWR8_2;
	wire w_dff_B_3fuGERfV3_2;
	wire w_dff_B_xO7fNMXW9_2;
	wire w_dff_B_MPmlsFHX5_2;
	wire w_dff_B_QflfAzRo9_2;
	wire w_dff_B_IPHjuRXg6_2;
	wire w_dff_B_iNBJO3Iw4_2;
	wire w_dff_B_p1UJ8gvY2_2;
	wire w_dff_B_A70XKMX65_2;
	wire w_dff_B_xVATjQpv2_2;
	wire w_dff_B_FfQGHvcz9_2;
	wire w_dff_B_tpDpCILF9_2;
	wire w_dff_B_y7UBxaVe9_2;
	wire w_dff_B_t3zvDPvW5_2;
	wire w_dff_B_sdIisz9O7_2;
	wire w_dff_B_j20DL4N69_2;
	wire w_dff_B_8ay992s14_2;
	wire w_dff_B_0a14F5911_2;
	wire w_dff_B_ljbBY7Lj5_2;
	wire w_dff_B_vAfuBllz1_2;
	wire w_dff_B_9R6hN7230_2;
	wire w_dff_B_6eoxZfhQ4_2;
	wire w_dff_B_6LRWDamo4_2;
	wire w_dff_B_8fNPFrdf1_2;
	wire w_dff_B_aapST4Cv0_2;
	wire w_dff_B_UJh4Cvpm5_2;
	wire w_dff_B_3Rj94cVZ0_2;
	wire w_dff_B_xrHz6jpY7_2;
	wire w_dff_B_UUKJBab72_2;
	wire w_dff_B_bWkcc7Z69_2;
	wire w_dff_B_Jayjf1Sp4_2;
	wire w_dff_B_okZPYfUy4_1;
	wire w_dff_B_2FHgVOBY5_2;
	wire w_dff_B_AiUKz9DE9_2;
	wire w_dff_B_GxH1MmvG7_2;
	wire w_dff_B_m4tnjpuY3_2;
	wire w_dff_B_cfai8G0e3_2;
	wire w_dff_B_KKUPwmjX8_2;
	wire w_dff_B_aDOm0Xx91_2;
	wire w_dff_B_Rj9sCT1D3_2;
	wire w_dff_B_CPqFrG2y8_2;
	wire w_dff_B_3tQuH77c7_2;
	wire w_dff_B_0e7vG31u5_2;
	wire w_dff_B_TdBal9S57_2;
	wire w_dff_B_ft8Dn88k7_2;
	wire w_dff_B_e01OjxXX3_2;
	wire w_dff_B_AW0MOot52_2;
	wire w_dff_B_jl81WEhp0_2;
	wire w_dff_B_rBITXdHJ1_2;
	wire w_dff_B_RMp93ep76_2;
	wire w_dff_B_Pq315Gmc5_2;
	wire w_dff_B_GjW8idSO6_2;
	wire w_dff_B_PcNx6c0N0_2;
	wire w_dff_B_7AyP6H7O7_2;
	wire w_dff_B_rY2At0qi5_2;
	wire w_dff_B_uQXcYRnD8_2;
	wire w_dff_B_3HOUjZ767_2;
	wire w_dff_B_Q8KQnlZG4_2;
	wire w_dff_B_BfZmWP7T6_2;
	wire w_dff_B_TsQO7Wvf1_2;
	wire w_dff_B_zzPrbLCm3_2;
	wire w_dff_B_Te1i66hV5_2;
	wire w_dff_B_htUOUhmr2_2;
	wire w_dff_B_SvxBL2CX5_2;
	wire w_dff_B_XFH8kGgb9_2;
	wire w_dff_B_Eat20wwF4_2;
	wire w_dff_B_p53BAToJ1_2;
	wire w_dff_B_1If2QCPg3_2;
	wire w_dff_B_QzXJUNAG0_2;
	wire w_dff_B_Yt2BTntV6_2;
	wire w_dff_B_5Tscc3mU5_2;
	wire w_dff_B_46wlq6IK4_2;
	wire w_dff_B_GkOsAjCA5_1;
	wire w_dff_B_qCfy96cX7_2;
	wire w_dff_B_qWFkwedW8_2;
	wire w_dff_B_ETqTeCqg5_2;
	wire w_dff_B_mrs8oaK01_2;
	wire w_dff_B_Ym8bGeRl2_2;
	wire w_dff_B_DsylCa3W7_2;
	wire w_dff_B_ij8RsBNT2_2;
	wire w_dff_B_s822BQXD2_2;
	wire w_dff_B_4LJR26Zz4_2;
	wire w_dff_B_I8FsOP383_2;
	wire w_dff_B_4TyCm9ea4_2;
	wire w_dff_B_jNm1oBz20_2;
	wire w_dff_B_yDvWNEvw1_2;
	wire w_dff_B_jQSi0nhl7_2;
	wire w_dff_B_zYfO4QD10_2;
	wire w_dff_B_npo0KMU07_2;
	wire w_dff_B_zNGsRY8g2_2;
	wire w_dff_B_rm5N9AZt7_2;
	wire w_dff_B_wgWjRY6A8_2;
	wire w_dff_B_BOFFIOU05_2;
	wire w_dff_B_Gxmvnb5R5_2;
	wire w_dff_B_XvF3he9e9_2;
	wire w_dff_B_3LlcdKAo3_2;
	wire w_dff_B_a6VJsaRx5_2;
	wire w_dff_B_fj0iVqtX8_2;
	wire w_dff_B_fhlgibW17_2;
	wire w_dff_B_Cp7XneBh6_2;
	wire w_dff_B_5IhKFno72_2;
	wire w_dff_B_SDTPaPew4_2;
	wire w_dff_B_LosGJHyD2_2;
	wire w_dff_B_olGrOOJb1_2;
	wire w_dff_B_2MIsppXc9_2;
	wire w_dff_B_t4jWqFVG6_2;
	wire w_dff_B_OZ6qpPTy4_2;
	wire w_dff_B_wnkFhy2N6_2;
	wire w_dff_B_XlSilwFu7_2;
	wire w_dff_B_yriLKFxM6_2;
	wire w_dff_B_eWRukfmw4_1;
	wire w_dff_B_ydnRlVpB3_2;
	wire w_dff_B_w7fsqj4P0_2;
	wire w_dff_B_ObquUWuS3_2;
	wire w_dff_B_HB8JQfSM1_2;
	wire w_dff_B_F02MSOvL3_2;
	wire w_dff_B_FGbvqy2Q7_2;
	wire w_dff_B_QQupTRmD1_2;
	wire w_dff_B_71fpE7MR4_2;
	wire w_dff_B_NauiZ4Fy0_2;
	wire w_dff_B_RX9WqM9h0_2;
	wire w_dff_B_XI0Fftw28_2;
	wire w_dff_B_JPYRxwGb9_2;
	wire w_dff_B_5PY4syl25_2;
	wire w_dff_B_rM1B12IR7_2;
	wire w_dff_B_kzbweZEn4_2;
	wire w_dff_B_hPe3EIBr9_2;
	wire w_dff_B_jlKiSpEy3_2;
	wire w_dff_B_SvRxmqY43_2;
	wire w_dff_B_sVpnHyj48_2;
	wire w_dff_B_ZtETKS3z6_2;
	wire w_dff_B_moEckjPF2_2;
	wire w_dff_B_go3ZHA9c7_2;
	wire w_dff_B_nbiclrTt7_2;
	wire w_dff_B_ZGsriYPt7_2;
	wire w_dff_B_H2jBMIvq9_2;
	wire w_dff_B_RGsD2Ahi9_2;
	wire w_dff_B_3h3hCPL00_2;
	wire w_dff_B_MAN844QY8_2;
	wire w_dff_B_iHtcMqOh4_2;
	wire w_dff_B_KCXcFZxf4_2;
	wire w_dff_B_Ba1c2bqR6_2;
	wire w_dff_B_nAh4pjQW7_2;
	wire w_dff_B_L0ho2uIT0_2;
	wire w_dff_B_2vJ0ECc04_2;
	wire w_dff_B_FmIUrn9u6_1;
	wire w_dff_B_YhOheFMg0_2;
	wire w_dff_B_5cIrRVT33_2;
	wire w_dff_B_kOYBXiHE9_2;
	wire w_dff_B_M6Wwa9E80_2;
	wire w_dff_B_IbJm1Q2G1_2;
	wire w_dff_B_o65yV4W44_2;
	wire w_dff_B_oq3h95fv5_2;
	wire w_dff_B_YPRjFFTg2_2;
	wire w_dff_B_9jWxiIwf0_2;
	wire w_dff_B_9oihohtO2_2;
	wire w_dff_B_3L40jCqf7_2;
	wire w_dff_B_zL8YWxPk1_2;
	wire w_dff_B_5xWILhr79_2;
	wire w_dff_B_gRWqRPTD8_2;
	wire w_dff_B_Xvrm9jtV6_2;
	wire w_dff_B_M2GUvrHP8_2;
	wire w_dff_B_ezwzdqy06_2;
	wire w_dff_B_UTwgntyC9_2;
	wire w_dff_B_SyqnNlG53_2;
	wire w_dff_B_dXG8MYI47_2;
	wire w_dff_B_bivUJdQg9_2;
	wire w_dff_B_0hyWc2yJ5_2;
	wire w_dff_B_YkUMhdsQ6_2;
	wire w_dff_B_ALrXiQfO9_2;
	wire w_dff_B_3o62TwvU7_2;
	wire w_dff_B_hv9kSpGt7_2;
	wire w_dff_B_Cl89ITno8_2;
	wire w_dff_B_bvYFSfcm1_2;
	wire w_dff_B_4xLBcRnD9_2;
	wire w_dff_B_pMWVECVB6_2;
	wire w_dff_B_UImGPrEg1_2;
	wire w_dff_B_X9x5eONG1_1;
	wire w_dff_B_lfBrzUrz6_2;
	wire w_dff_B_I4gDPI392_2;
	wire w_dff_B_BYaGUQBu7_2;
	wire w_dff_B_4SEIkHOT4_2;
	wire w_dff_B_FoWaM2DB1_2;
	wire w_dff_B_vtqDLHrl3_2;
	wire w_dff_B_qlO9WPcz7_2;
	wire w_dff_B_Gv3WRA0O5_2;
	wire w_dff_B_Hym1lT2v2_2;
	wire w_dff_B_QnELvtVC3_2;
	wire w_dff_B_z5fmOBeh4_2;
	wire w_dff_B_xfTH8nsm5_2;
	wire w_dff_B_PwRJ4YaM8_2;
	wire w_dff_B_VIYUXkdD6_2;
	wire w_dff_B_c2ygEIGp6_2;
	wire w_dff_B_8K4SJKp38_2;
	wire w_dff_B_8WTgtnfC7_2;
	wire w_dff_B_URCHDs8v9_2;
	wire w_dff_B_y35Sv2AP7_2;
	wire w_dff_B_Oyr3oh2T5_2;
	wire w_dff_B_kj4TQQJI6_2;
	wire w_dff_B_U5nNO81N0_2;
	wire w_dff_B_W06xmaZP0_2;
	wire w_dff_B_gq6YKjlZ3_2;
	wire w_dff_B_bm1ZlNgl4_2;
	wire w_dff_B_HD6R4fCa1_2;
	wire w_dff_B_GZNE8dma7_2;
	wire w_dff_B_VDExURbU0_2;
	wire w_dff_B_70voapNf1_1;
	wire w_dff_B_TnajQOjF5_2;
	wire w_dff_B_nX7Vn4xJ0_2;
	wire w_dff_B_T0Uzh5Y36_2;
	wire w_dff_B_x0u8nhnw7_2;
	wire w_dff_B_jaIlhc4N4_2;
	wire w_dff_B_e4TP2vWq7_2;
	wire w_dff_B_nxV8kibe6_2;
	wire w_dff_B_c0u3t53e8_2;
	wire w_dff_B_PIbZcqUT2_2;
	wire w_dff_B_91UUNVtU3_2;
	wire w_dff_B_wFMIMidM1_2;
	wire w_dff_B_8t7O4wBV8_2;
	wire w_dff_B_tRlUm20j6_2;
	wire w_dff_B_QyVkVUSp4_2;
	wire w_dff_B_YymKICMc9_2;
	wire w_dff_B_aCMHH9qC4_2;
	wire w_dff_B_hwY2v7cA7_2;
	wire w_dff_B_vVhDKRVx4_2;
	wire w_dff_B_6WwIKGxL4_2;
	wire w_dff_B_TRxvA4oM1_2;
	wire w_dff_B_QFo2R29W7_2;
	wire w_dff_B_lWDsRKFF7_2;
	wire w_dff_B_Wa67a40Z2_2;
	wire w_dff_B_2mA5JmjA2_2;
	wire w_dff_B_5ffPzOR82_2;
	wire w_dff_B_AojH413d8_1;
	wire w_dff_B_bojL8AXu1_2;
	wire w_dff_B_SFc7Rnd68_2;
	wire w_dff_B_UEQUFxnz8_2;
	wire w_dff_B_5pgdEYHc1_2;
	wire w_dff_B_Ek4SrkcL4_2;
	wire w_dff_B_Ykuj1MrY5_2;
	wire w_dff_B_Z8op9tpd0_2;
	wire w_dff_B_5E3MbnFt2_2;
	wire w_dff_B_WVyxDF8I4_2;
	wire w_dff_B_b1NwTAOJ4_2;
	wire w_dff_B_lNHeQRKb6_2;
	wire w_dff_B_VAyTxHL41_2;
	wire w_dff_B_fTBCHUgh1_2;
	wire w_dff_B_DQMvKJ7t2_2;
	wire w_dff_B_g8yulbvU8_2;
	wire w_dff_B_H6I1go5J2_2;
	wire w_dff_B_DWQ0Z7NF1_2;
	wire w_dff_B_3naLMSS43_2;
	wire w_dff_B_LKYOLMbw2_2;
	wire w_dff_B_Xe8hfpQ35_2;
	wire w_dff_B_djo0VUY31_2;
	wire w_dff_B_IUpPIGVx7_2;
	wire w_dff_B_fmHAL9ae8_1;
	wire w_dff_B_p0tE444d6_2;
	wire w_dff_B_K7UTe42L6_2;
	wire w_dff_B_usZ9fHwx7_2;
	wire w_dff_B_CbklaxfM4_2;
	wire w_dff_B_nYoSMv0S4_2;
	wire w_dff_B_Y01bI1t40_2;
	wire w_dff_B_lyYWGvSQ6_2;
	wire w_dff_B_SpMFarON3_2;
	wire w_dff_B_wHlfpW2R6_2;
	wire w_dff_B_2SCrIjwV1_2;
	wire w_dff_B_DAxOj5kw2_2;
	wire w_dff_B_F5LGktB03_2;
	wire w_dff_B_dL8pwDjZ5_2;
	wire w_dff_B_4125E9pF6_2;
	wire w_dff_B_ouX0EVPl2_2;
	wire w_dff_B_cMnm8UwX8_2;
	wire w_dff_B_YZicZTeH6_2;
	wire w_dff_B_JOVUyAjR9_2;
	wire w_dff_B_XIqTUG0R2_2;
	wire w_dff_B_C3gKgd3D9_1;
	wire w_dff_B_UIQ4Tq8K0_2;
	wire w_dff_B_xZKQC6Z66_2;
	wire w_dff_B_lNb5zbNw0_2;
	wire w_dff_B_ga64F56D5_2;
	wire w_dff_B_d7xdTB787_2;
	wire w_dff_B_2feWtac50_2;
	wire w_dff_B_WQK4Y9oX0_2;
	wire w_dff_B_Yk8M5kI21_2;
	wire w_dff_B_f4xQt3x57_2;
	wire w_dff_B_eYPa24kv9_2;
	wire w_dff_B_5xrQ4LJY0_2;
	wire w_dff_B_fErRU8Wa4_2;
	wire w_dff_B_Bd6Lq7wK7_2;
	wire w_dff_B_x36fGRs87_2;
	wire w_dff_B_D8eIa9Ef0_2;
	wire w_dff_B_uF078E1D9_2;
	wire w_dff_B_sw5cd2Qe4_1;
	wire w_dff_B_FGIlsyaX8_2;
	wire w_dff_B_n0mfdLxC7_2;
	wire w_dff_B_62jIwzj55_2;
	wire w_dff_B_XhVzmfEv7_2;
	wire w_dff_B_5eJCXF1s5_2;
	wire w_dff_B_NOQRRBaB4_2;
	wire w_dff_B_kHeG3J936_2;
	wire w_dff_B_YZ9xqlzj5_2;
	wire w_dff_B_iHiiKhso8_2;
	wire w_dff_B_1lthIbJN1_2;
	wire w_dff_B_ZEY1crJr7_2;
	wire w_dff_B_54IVPH8S9_2;
	wire w_dff_B_jEXVVydu5_2;
	wire w_dff_B_w72PYw6U1_1;
	wire w_dff_B_GVirOKkz8_2;
	wire w_dff_B_8VwgNTfV6_2;
	wire w_dff_B_LGWtgeBN4_2;
	wire w_dff_B_p1Qsan2p5_2;
	wire w_dff_B_KAxhzIm75_2;
	wire w_dff_B_FNNwejJq3_2;
	wire w_dff_B_BMlDPU3H2_2;
	wire w_dff_B_j38HnXvi8_2;
	wire w_dff_B_LmNVtie13_2;
	wire w_dff_B_LCG7Dk6n8_2;
	wire w_dff_B_JyHIx9uu1_2;
	wire w_dff_B_thuy0MMT4_1;
	wire w_dff_B_ljJHdLN36_2;
	wire w_dff_B_h6o6Ds5F7_2;
	wire w_dff_B_YtVsayaB5_2;
	wire w_dff_B_cjpEUtrF4_2;
	wire w_dff_B_5WzQe57n6_2;
	wire w_dff_B_sUOIGnBS8_2;
	wire w_dff_B_6texNomC5_2;
	wire w_dff_B_q5ZAGjY43_2;
	wire w_dff_B_ZYfDr3Pu6_2;
	wire w_dff_B_rXwee7iy7_2;
	wire w_dff_B_z4cPPlU19_0;
	wire w_dff_A_UHb6hdmf2_0;
	wire w_dff_A_OoN2Prmy8_0;
	wire w_dff_A_xqfz72US4_1;
	wire w_dff_A_U7KNUsVf3_1;
	wire w_dff_B_QvWK9LdJ4_1;
	wire w_dff_B_ppWMHWH82_2;
	wire w_dff_B_Du9yRvuv4_2;
	wire w_dff_B_rfOzPZWh0_2;
	wire w_dff_B_YRD4GLRA9_2;
	wire w_dff_B_qtVBLd7Y9_2;
	wire w_dff_B_xXxxeo2k8_2;
	wire w_dff_B_d8ZyoDXL4_2;
	wire w_dff_B_ZSyl96Lv8_2;
	wire w_dff_B_ty4Ue4Zf2_2;
	wire w_dff_B_QUKVixNC3_2;
	wire w_dff_B_EAF4somy5_2;
	wire w_dff_B_C9a3ZSxp0_2;
	wire w_dff_B_tNmU4ROw3_2;
	wire w_dff_B_8gGogAKO4_2;
	wire w_dff_B_iHw0yWVS2_2;
	wire w_dff_B_BfLDeT4F0_2;
	wire w_dff_B_HHnTZyAA9_2;
	wire w_dff_B_6myBpVsI6_2;
	wire w_dff_B_RKm6MBC72_2;
	wire w_dff_B_CYVv1W5i4_2;
	wire w_dff_B_l3al1kNK2_2;
	wire w_dff_B_6DiyvSLa4_2;
	wire w_dff_B_coAxeVZi2_2;
	wire w_dff_B_Bm9ZbwX94_2;
	wire w_dff_B_DSTJ5NN37_2;
	wire w_dff_B_bvZFtliG9_2;
	wire w_dff_B_U2I4LaUO3_2;
	wire w_dff_B_3EmoHhCN9_2;
	wire w_dff_B_vpWzQMEl9_2;
	wire w_dff_B_RaFgWQMW8_2;
	wire w_dff_B_85e4b9YS0_2;
	wire w_dff_B_TwqKLTjI6_2;
	wire w_dff_B_IJpz2FlE4_2;
	wire w_dff_B_RXGS2Cq57_2;
	wire w_dff_B_NqeVhiCF4_2;
	wire w_dff_B_KE23DJSF1_2;
	wire w_dff_B_27oEDSQy4_2;
	wire w_dff_B_WcwpsT4j7_2;
	wire w_dff_B_OhiqQqoW1_2;
	wire w_dff_B_e4TzaCi25_2;
	wire w_dff_B_zgaLzjm17_2;
	wire w_dff_B_ufmkUT7W0_2;
	wire w_dff_B_OfDykzgp6_2;
	wire w_dff_B_769FflUu8_2;
	wire w_dff_B_cWIKRbme5_2;
	wire w_dff_B_bG14cOkU1_2;
	wire w_dff_B_xTRmInr30_0;
	wire w_dff_A_Z1NK3AwW0_1;
	wire w_dff_B_JumOCHSu3_1;
	wire w_dff_B_djXDBNZ67_2;
	wire w_dff_B_rgShl3M96_2;
	wire w_dff_B_MbQSwguy8_2;
	wire w_dff_B_rTXAzY9u6_2;
	wire w_dff_B_TAxIsREk8_2;
	wire w_dff_B_SWI5FPZO2_2;
	wire w_dff_B_nES1lzeJ1_2;
	wire w_dff_B_6yVykT7u9_2;
	wire w_dff_B_X9DvH45u2_2;
	wire w_dff_B_TOFT54Yp0_2;
	wire w_dff_B_OdCsBtY38_2;
	wire w_dff_B_g10y2h3c7_2;
	wire w_dff_B_f3DeNnlr7_2;
	wire w_dff_B_SxCiQWFo4_2;
	wire w_dff_B_v9SIsnLb9_2;
	wire w_dff_B_ZNzTCBjo3_2;
	wire w_dff_B_egjYoBMq4_2;
	wire w_dff_B_k4CU2HWw1_2;
	wire w_dff_B_faOXZq9f7_2;
	wire w_dff_B_Ztrfcz5F5_2;
	wire w_dff_B_an9KytBv9_2;
	wire w_dff_B_LTd2AH0n9_2;
	wire w_dff_B_vd0NwYDS0_2;
	wire w_dff_B_jpAy5BiJ6_2;
	wire w_dff_B_Jx3w7Wv96_2;
	wire w_dff_B_mx0KoNRe1_2;
	wire w_dff_B_Lrim48jw3_2;
	wire w_dff_B_Gywrwyt91_2;
	wire w_dff_B_4stycAfw9_2;
	wire w_dff_B_5v1tJlmS4_2;
	wire w_dff_B_o9DQ50o20_2;
	wire w_dff_B_EMoVDda25_2;
	wire w_dff_B_480Yo4J14_2;
	wire w_dff_B_KftfVnJe9_2;
	wire w_dff_B_6Q6U5BxS6_2;
	wire w_dff_B_lgHEpE4d0_2;
	wire w_dff_B_KgXNBHXA8_2;
	wire w_dff_B_0qqmCVOu2_2;
	wire w_dff_B_cyDokG0S9_2;
	wire w_dff_B_GRujP2cX2_2;
	wire w_dff_B_sDfgSwXx5_2;
	wire w_dff_B_OeZSAjlN6_2;
	wire w_dff_B_48fLUiLC1_1;
	wire w_dff_B_Ze3kLx3K1_2;
	wire w_dff_B_D0RzeeaR9_2;
	wire w_dff_B_uvEPI7238_2;
	wire w_dff_B_1GtuQFdD7_2;
	wire w_dff_B_6I9bN3aj2_2;
	wire w_dff_B_pDkBuq3W4_2;
	wire w_dff_B_l6egQqTq1_2;
	wire w_dff_B_EeIx6lWu5_2;
	wire w_dff_B_ZKzze1G45_2;
	wire w_dff_B_5EIQBByw2_2;
	wire w_dff_B_WnUd9fAB9_2;
	wire w_dff_B_XJ7ye8VP4_2;
	wire w_dff_B_iATijlvg3_2;
	wire w_dff_B_WJsVMLVr2_2;
	wire w_dff_B_SoQN8u6O6_2;
	wire w_dff_B_WMpKEzfw9_2;
	wire w_dff_B_VyaUp4V64_2;
	wire w_dff_B_eOWDQZM86_2;
	wire w_dff_B_9fiXV1DK3_2;
	wire w_dff_B_cVKcOvl73_2;
	wire w_dff_B_2cCtsE6g0_2;
	wire w_dff_B_QFeoGzuf5_2;
	wire w_dff_B_MpVpW8QW2_2;
	wire w_dff_B_9I3MpTzM1_2;
	wire w_dff_B_FsC1pxoD0_2;
	wire w_dff_B_npHzAUx52_2;
	wire w_dff_B_lmkokJKy3_2;
	wire w_dff_B_Nla71nIv1_2;
	wire w_dff_B_rBTTfBLi3_2;
	wire w_dff_B_OsS6zM8y5_2;
	wire w_dff_B_j7TGoQOg7_2;
	wire w_dff_B_1xncBhks8_2;
	wire w_dff_B_aauT4CO23_2;
	wire w_dff_B_hK8ZzDrd1_2;
	wire w_dff_B_OzuIHOuw2_2;
	wire w_dff_B_SyOUUt9X8_2;
	wire w_dff_B_yX9rmHxl6_2;
	wire w_dff_B_tUH2K1Kj7_2;
	wire w_dff_B_lcTOel7j3_2;
	wire w_dff_B_uDtCWuTI2_1;
	wire w_dff_B_6Yaw6uqx5_2;
	wire w_dff_B_LKpBOd4S8_2;
	wire w_dff_B_yJLB6yw02_2;
	wire w_dff_B_GsbWfNwj8_2;
	wire w_dff_B_z9ITqEVW7_2;
	wire w_dff_B_p9IB5jVJ4_2;
	wire w_dff_B_EDkMg6i13_2;
	wire w_dff_B_lP6sjAII6_2;
	wire w_dff_B_8h7NaPld4_2;
	wire w_dff_B_J6f9wVXD2_2;
	wire w_dff_B_KD3qxIVs4_2;
	wire w_dff_B_txNDtw8o4_2;
	wire w_dff_B_GpM0pypo0_2;
	wire w_dff_B_iCeFsNNo9_2;
	wire w_dff_B_CUFHkhrZ5_2;
	wire w_dff_B_GIlZr1Dv9_2;
	wire w_dff_B_DEd7KeBy8_2;
	wire w_dff_B_NrOlrH518_2;
	wire w_dff_B_Lth8MXWF7_2;
	wire w_dff_B_GH5mXvln3_2;
	wire w_dff_B_nWFoS2jl6_2;
	wire w_dff_B_xiXCikwH9_2;
	wire w_dff_B_jQFxVyoR7_2;
	wire w_dff_B_i0DgvZ6z9_2;
	wire w_dff_B_psaKYNCg1_2;
	wire w_dff_B_zO67d4XR7_2;
	wire w_dff_B_PchzTo831_2;
	wire w_dff_B_FhYYglJE0_2;
	wire w_dff_B_0Z8dxuCq2_2;
	wire w_dff_B_raInsWt43_2;
	wire w_dff_B_xjhE7TFx1_2;
	wire w_dff_B_wtkhyI6N7_2;
	wire w_dff_B_MB2L94Ng8_2;
	wire w_dff_B_Jhi8veVz7_2;
	wire w_dff_B_1dOlMKis6_2;
	wire w_dff_B_Jne99qpP9_2;
	wire w_dff_B_wqdKiwbS9_1;
	wire w_dff_B_CHpjLhuk3_2;
	wire w_dff_B_LpyoHiG38_2;
	wire w_dff_B_oT9evhYB1_2;
	wire w_dff_B_YfPu9CoH1_2;
	wire w_dff_B_58QxJlSM5_2;
	wire w_dff_B_zteXz2tj4_2;
	wire w_dff_B_tzSbd6xs9_2;
	wire w_dff_B_QoKpxNwm7_2;
	wire w_dff_B_1HGe7cXS1_2;
	wire w_dff_B_btzooBeW8_2;
	wire w_dff_B_pWBrxOSL1_2;
	wire w_dff_B_DPu6pGJB2_2;
	wire w_dff_B_AzLLaukc4_2;
	wire w_dff_B_9VsHYNVU5_2;
	wire w_dff_B_R2wqIfy29_2;
	wire w_dff_B_61Mi9vDS6_2;
	wire w_dff_B_m9xDWTid6_2;
	wire w_dff_B_CcgNIaTM2_2;
	wire w_dff_B_h5OAkxsp3_2;
	wire w_dff_B_HEGYzhwY5_2;
	wire w_dff_B_kfbk9PY04_2;
	wire w_dff_B_jmaO7NWx0_2;
	wire w_dff_B_TShXzsna3_2;
	wire w_dff_B_pNS8rVN69_2;
	wire w_dff_B_hFPCJFyh2_2;
	wire w_dff_B_A0tafV0w9_2;
	wire w_dff_B_AEbfou5c6_2;
	wire w_dff_B_K75tx89b6_2;
	wire w_dff_B_wzPUwsfF3_2;
	wire w_dff_B_ZZcJZLBn4_2;
	wire w_dff_B_4VF6pijT7_2;
	wire w_dff_B_4HCmCGDr6_2;
	wire w_dff_B_xjUxkvVQ5_2;
	wire w_dff_B_Ks3Cgzof9_1;
	wire w_dff_B_LotTPgHT2_2;
	wire w_dff_B_eiVwXRlF0_2;
	wire w_dff_B_GApNkSkT3_2;
	wire w_dff_B_0UPiT9ic9_2;
	wire w_dff_B_Il2GKSpk7_2;
	wire w_dff_B_lUTGmdDb2_2;
	wire w_dff_B_xuW5NKz55_2;
	wire w_dff_B_w1R3Xp8i3_2;
	wire w_dff_B_DQw6JW6I5_2;
	wire w_dff_B_ThdgcyjF7_2;
	wire w_dff_B_Fm0jZ2AS0_2;
	wire w_dff_B_9hfurshI2_2;
	wire w_dff_B_fFRCeOFU6_2;
	wire w_dff_B_sL9yCUtx2_2;
	wire w_dff_B_zBNIm5ku7_2;
	wire w_dff_B_35zlfNO25_2;
	wire w_dff_B_ozIz7hsk9_2;
	wire w_dff_B_iBDx4kTa8_2;
	wire w_dff_B_FRqwOUtL0_2;
	wire w_dff_B_5SioB8bi0_2;
	wire w_dff_B_dRfhkIXO6_2;
	wire w_dff_B_meGfJ4Ml7_2;
	wire w_dff_B_THRXSfUE3_2;
	wire w_dff_B_djv53PIm9_2;
	wire w_dff_B_EQBEhJzu3_2;
	wire w_dff_B_SbD6dXDL5_2;
	wire w_dff_B_PZcz0VKj4_2;
	wire w_dff_B_Vv5vw15y6_2;
	wire w_dff_B_wqQfrI6j6_2;
	wire w_dff_B_xho3upNn0_2;
	wire w_dff_B_fiFeTNe63_1;
	wire w_dff_B_9HwILk8E8_2;
	wire w_dff_B_BmLP96EL6_2;
	wire w_dff_B_95OsEaqm3_2;
	wire w_dff_B_u1vD9SdR2_2;
	wire w_dff_B_iyhTj8nm2_2;
	wire w_dff_B_M4IeJZNd0_2;
	wire w_dff_B_ZEyAsnHN7_2;
	wire w_dff_B_4WlfT4Mr9_2;
	wire w_dff_B_tbs6DpMD0_2;
	wire w_dff_B_L8MrorfR3_2;
	wire w_dff_B_u8g5p00Q1_2;
	wire w_dff_B_5dMGJnKw8_2;
	wire w_dff_B_auTy16xV2_2;
	wire w_dff_B_jzl2WbeF3_2;
	wire w_dff_B_VAok8B1c7_2;
	wire w_dff_B_UYzEA5X27_2;
	wire w_dff_B_d2Gkv2e39_2;
	wire w_dff_B_0eXg0p0U9_2;
	wire w_dff_B_xiRj92M16_2;
	wire w_dff_B_u6oZYj6j5_2;
	wire w_dff_B_TnozkIyp2_2;
	wire w_dff_B_qnhEsylH2_2;
	wire w_dff_B_qkhO7al72_2;
	wire w_dff_B_y6kwC2sf6_2;
	wire w_dff_B_vV0bDt1L1_2;
	wire w_dff_B_lZ5Qjorr3_2;
	wire w_dff_B_bcP0E7Hi5_2;
	wire w_dff_B_PDENw4BN8_1;
	wire w_dff_B_hNgHePwe0_2;
	wire w_dff_B_LygJ5N0O7_2;
	wire w_dff_B_vLA6d5pQ6_2;
	wire w_dff_B_Cgfh33L38_2;
	wire w_dff_B_SlTnutle6_2;
	wire w_dff_B_piViiJcf3_2;
	wire w_dff_B_o90DMMD02_2;
	wire w_dff_B_4XRK2MfO1_2;
	wire w_dff_B_Umx2e0Ti1_2;
	wire w_dff_B_V9ZXbxxY2_2;
	wire w_dff_B_ptmoT6kf6_2;
	wire w_dff_B_uyGMp8xf6_2;
	wire w_dff_B_0aqzSceQ4_2;
	wire w_dff_B_WfaHkpyi8_2;
	wire w_dff_B_FQgo4IeQ5_2;
	wire w_dff_B_aHhwdnR76_2;
	wire w_dff_B_EZTUX7EG6_2;
	wire w_dff_B_11je3hXV5_2;
	wire w_dff_B_dNzfvh2j6_2;
	wire w_dff_B_ii4FWdKs3_2;
	wire w_dff_B_PMTWwnZD2_2;
	wire w_dff_B_2R7uQTqB7_2;
	wire w_dff_B_Jyz2QApv5_2;
	wire w_dff_B_JBIaOyn81_2;
	wire w_dff_B_yT5jobxk4_1;
	wire w_dff_B_7JAqNfso5_2;
	wire w_dff_B_retg5sal1_2;
	wire w_dff_B_A4vrtnSH3_2;
	wire w_dff_B_qlYry9lt8_2;
	wire w_dff_B_r1y2DTad6_2;
	wire w_dff_B_IpJS6Yjr3_2;
	wire w_dff_B_aSytTE3v5_2;
	wire w_dff_B_eA3eVsOS5_2;
	wire w_dff_B_NmyyoUbH7_2;
	wire w_dff_B_N30qgxtY5_2;
	wire w_dff_B_sBD5fOAS7_2;
	wire w_dff_B_ROiWYELl3_2;
	wire w_dff_B_JwGCPUiN1_2;
	wire w_dff_B_QP6oDmvm3_2;
	wire w_dff_B_IrJyoUG20_2;
	wire w_dff_B_Vh5xl8JH8_2;
	wire w_dff_B_uhyn0yt57_2;
	wire w_dff_B_8vJAl03n1_2;
	wire w_dff_B_3r6Rjrm44_2;
	wire w_dff_B_QJ1fA5oe5_2;
	wire w_dff_B_OBfPOlGw5_2;
	wire w_dff_B_Y00TVUep1_1;
	wire w_dff_B_GBVQ5kQi4_2;
	wire w_dff_B_emarn5hR8_2;
	wire w_dff_B_xo7lOydL0_2;
	wire w_dff_B_1y3bl1DT5_2;
	wire w_dff_B_S8pJRnZ08_2;
	wire w_dff_B_zyBgXcK69_2;
	wire w_dff_B_2l6JgLO20_2;
	wire w_dff_B_vvGstb3u6_2;
	wire w_dff_B_Ojxe2w5V1_2;
	wire w_dff_B_NJQC5RLN1_2;
	wire w_dff_B_xkyLc5QC5_2;
	wire w_dff_B_g4Xk05fy1_2;
	wire w_dff_B_LojWqOlZ3_2;
	wire w_dff_B_B9DS5n4x2_2;
	wire w_dff_B_UzAZefYP7_2;
	wire w_dff_B_zRtuluKM3_2;
	wire w_dff_B_uqRp0sXY8_2;
	wire w_dff_B_dnBmfhxP0_2;
	wire w_dff_B_3HGlLHHK0_1;
	wire w_dff_B_YfSYz0J25_2;
	wire w_dff_B_zRZmOvmZ9_2;
	wire w_dff_B_vHLmVdCp7_2;
	wire w_dff_B_WeDC8Aqf4_2;
	wire w_dff_B_pCDmsHui1_2;
	wire w_dff_B_A5EVWbOE0_2;
	wire w_dff_B_ygM08s7E1_2;
	wire w_dff_B_IIZZ6ubz3_2;
	wire w_dff_B_rCEn5z0B8_2;
	wire w_dff_B_Xo7uSpIc3_2;
	wire w_dff_B_AUIvz5kU7_2;
	wire w_dff_B_6J6Zapwv8_2;
	wire w_dff_B_Qds8q9tS3_2;
	wire w_dff_B_3uAKOUMy2_2;
	wire w_dff_B_aW03qvsr3_2;
	wire w_dff_B_5W1HNHhA0_1;
	wire w_dff_B_zeqJF3l42_2;
	wire w_dff_B_EX0KBTux0_2;
	wire w_dff_B_40DQ05gC1_2;
	wire w_dff_B_ispNmflQ4_2;
	wire w_dff_B_SUYk7Gpm9_2;
	wire w_dff_B_0wiadfvI9_2;
	wire w_dff_B_wCwrZ7sT0_2;
	wire w_dff_B_Ez6ZSNkI5_2;
	wire w_dff_B_9qG03qPU5_2;
	wire w_dff_B_lFuhzVqH5_2;
	wire w_dff_B_YFOUAA3M5_2;
	wire w_dff_B_H0YJAthz5_2;
	wire w_dff_B_TG7ggu479_1;
	wire w_dff_B_gICaoszp8_2;
	wire w_dff_B_AQ3BNbBd1_2;
	wire w_dff_B_LpODIpdX2_2;
	wire w_dff_B_qCK0mbns7_2;
	wire w_dff_B_yM5iZlxK9_2;
	wire w_dff_B_dE0RJCMY2_2;
	wire w_dff_B_BnSvBPJn0_2;
	wire w_dff_B_a5JaWE737_2;
	wire w_dff_B_StYRvpWz0_2;
	wire w_dff_B_xBcKVmxU9_2;
	wire w_dff_B_Baav93bQ4_2;
	wire w_dff_B_Cecb2C139_1;
	wire w_dff_B_LhXZKNt04_1;
	wire w_dff_B_GQQ7GrVa6_2;
	wire w_dff_B_tssskMr49_2;
	wire w_dff_B_XzIhFrPZ0_2;
	wire w_dff_B_wHOweIil2_0;
	wire w_dff_A_kPRBdduK3_0;
	wire w_dff_A_hmDCpiYY5_0;
	wire w_dff_A_ONStMVIT2_1;
	wire w_dff_A_Cqil93OE8_1;
	wire w_dff_B_tH64gZ2p2_1;
	wire w_dff_B_vsBkSVvQ9_2;
	wire w_dff_B_YDKIcx736_2;
	wire w_dff_B_wiQ12gCq0_2;
	wire w_dff_B_bc7mP5u12_2;
	wire w_dff_B_pJwiY3L16_2;
	wire w_dff_B_CfVTyzbr7_2;
	wire w_dff_B_3nC7AJco0_2;
	wire w_dff_B_z5Zy6f9Q3_2;
	wire w_dff_B_JiiRaLyT6_2;
	wire w_dff_B_dWWWBkCr0_2;
	wire w_dff_B_hVJNX2qw9_2;
	wire w_dff_B_8JGAj5iT2_2;
	wire w_dff_B_b6KKmoqP2_2;
	wire w_dff_B_p2xCU6m46_2;
	wire w_dff_B_uJrcZC8F0_2;
	wire w_dff_B_g1fcwlwt0_2;
	wire w_dff_B_gBggXZDR0_2;
	wire w_dff_B_qYAFNbPN4_2;
	wire w_dff_B_LXBC5JLy0_2;
	wire w_dff_B_BEpY2dra0_2;
	wire w_dff_B_oNRq0rgT5_2;
	wire w_dff_B_FUrM4H2e0_2;
	wire w_dff_B_hE4UHJNO5_2;
	wire w_dff_B_XpKPpW862_2;
	wire w_dff_B_Pukwssw95_2;
	wire w_dff_B_iDh9LQAv8_2;
	wire w_dff_B_zZ0kqyn91_2;
	wire w_dff_B_91ISSEBv4_2;
	wire w_dff_B_qPa29pS04_2;
	wire w_dff_B_kfwyd9nP9_2;
	wire w_dff_B_yrxVOoOE8_2;
	wire w_dff_B_AY7lYIUV9_2;
	wire w_dff_B_mrrtY6pt7_2;
	wire w_dff_B_LKQUuxjj8_2;
	wire w_dff_B_1kTDukAs5_2;
	wire w_dff_B_hUXzn7KH6_2;
	wire w_dff_B_njlmG7O59_2;
	wire w_dff_B_POyDQKv68_2;
	wire w_dff_B_4EvScwfw9_2;
	wire w_dff_B_Th3njhLC2_2;
	wire w_dff_B_w1gSjeAf4_2;
	wire w_dff_B_OsKlf9aE8_2;
	wire w_dff_B_2lysxwuL8_2;
	wire w_dff_B_NUZsT6f97_2;
	wire w_dff_B_ulbJp4165_2;
	wire w_dff_B_ERHUrecI3_2;
	wire w_dff_B_gnw9YzMm7_0;
	wire w_dff_A_0VYyg8st6_1;
	wire w_dff_B_mEub8Cht3_1;
	wire w_dff_B_04aaA9Pj2_2;
	wire w_dff_B_uGPEyDWy3_2;
	wire w_dff_B_Jw4gCK698_2;
	wire w_dff_B_4MHLehCB7_2;
	wire w_dff_B_mho9pv3N5_2;
	wire w_dff_B_9cKZPClz3_2;
	wire w_dff_B_aL7DujUi5_2;
	wire w_dff_B_WNed0ixx4_2;
	wire w_dff_B_RlHJfAZj3_2;
	wire w_dff_B_OXey3Q4g5_2;
	wire w_dff_B_Fb4TIpvM9_2;
	wire w_dff_B_hvDhxpSV8_2;
	wire w_dff_B_IlmlciXJ9_2;
	wire w_dff_B_NU3PDFub9_2;
	wire w_dff_B_kjDWGwKC5_2;
	wire w_dff_B_5EXv2p1d4_2;
	wire w_dff_B_f1JfoURg7_2;
	wire w_dff_B_VRDgX8f18_2;
	wire w_dff_B_GZkdl9En5_2;
	wire w_dff_B_I8KzF8wc2_2;
	wire w_dff_B_gaRqe6bL1_2;
	wire w_dff_B_kkHFDaT97_2;
	wire w_dff_B_SLCXx6yq3_2;
	wire w_dff_B_CIHttLD85_2;
	wire w_dff_B_LAMs7jrJ3_2;
	wire w_dff_B_Qp8Tv7Y91_2;
	wire w_dff_B_oeu70c2d3_2;
	wire w_dff_B_QyTblDHL5_2;
	wire w_dff_B_YqwMphmv2_2;
	wire w_dff_B_pC1cg0cG3_2;
	wire w_dff_B_D3KQpFdg0_2;
	wire w_dff_B_gDvfvCPO2_2;
	wire w_dff_B_zJAf4Cmw7_2;
	wire w_dff_B_IpZCzPRt6_2;
	wire w_dff_B_en0pEEKL1_2;
	wire w_dff_B_wsaxXHHs7_2;
	wire w_dff_B_IUhOhLE62_2;
	wire w_dff_B_jTOsY1Br4_2;
	wire w_dff_B_t6m14mr58_2;
	wire w_dff_B_7I4L68L81_2;
	wire w_dff_B_q3UgyzgI7_2;
	wire w_dff_B_LidCqk3d7_2;
	wire w_dff_B_0Um9Rg9s4_1;
	wire w_dff_B_FYeqss1r8_2;
	wire w_dff_B_0W5GxR8j8_2;
	wire w_dff_B_NEVodtvL7_2;
	wire w_dff_B_dS7nhfoN4_2;
	wire w_dff_B_DxMaCaeA6_2;
	wire w_dff_B_4DuoXHBK1_2;
	wire w_dff_B_xnHIWkkX9_2;
	wire w_dff_B_OguhmY5w5_2;
	wire w_dff_B_lrRq2WNd1_2;
	wire w_dff_B_LUS16xPf8_2;
	wire w_dff_B_0c9zDrv27_2;
	wire w_dff_B_2lR4bZBX6_2;
	wire w_dff_B_KgCCofJ52_2;
	wire w_dff_B_VJZliVqm8_2;
	wire w_dff_B_pbKSCjGs5_2;
	wire w_dff_B_XnRPovyT7_2;
	wire w_dff_B_u0kxdFDU7_2;
	wire w_dff_B_MNcbHyEE3_2;
	wire w_dff_B_Q4OwdjlL3_2;
	wire w_dff_B_o4bAO1UA8_2;
	wire w_dff_B_bBxnxwqF7_2;
	wire w_dff_B_nCngdcef7_2;
	wire w_dff_B_b1sbFnIp3_2;
	wire w_dff_B_Z51BpY3j1_2;
	wire w_dff_B_g0EJDHDJ5_2;
	wire w_dff_B_4gtwUJOe7_2;
	wire w_dff_B_XGXJ9S162_2;
	wire w_dff_B_lqSVTLqO9_2;
	wire w_dff_B_1ccNLfBt2_2;
	wire w_dff_B_ySeAm6lW3_2;
	wire w_dff_B_Tma7Mkyr4_2;
	wire w_dff_B_ry4mptlp7_2;
	wire w_dff_B_Y7zLzYTy3_2;
	wire w_dff_B_20eYAsih1_2;
	wire w_dff_B_WyUNR5Ew3_2;
	wire w_dff_B_P6uXQ72v4_2;
	wire w_dff_B_oSg6BDzv9_2;
	wire w_dff_B_i3Ve0M2d3_2;
	wire w_dff_B_389B8GSI6_2;
	wire w_dff_B_EEFDNy893_1;
	wire w_dff_B_9McnlYsm1_2;
	wire w_dff_B_pKf1HR1x4_2;
	wire w_dff_B_ZzQzMXrZ2_2;
	wire w_dff_B_rFb84YWB2_2;
	wire w_dff_B_7nHviEfH9_2;
	wire w_dff_B_81ooFWeb5_2;
	wire w_dff_B_YoHzIqbB8_2;
	wire w_dff_B_1ydIIUHn3_2;
	wire w_dff_B_s5ig4Y2j8_2;
	wire w_dff_B_rNt2kuqR7_2;
	wire w_dff_B_CgeR1ohU2_2;
	wire w_dff_B_0kXB4qhL2_2;
	wire w_dff_B_KB8LWmM05_2;
	wire w_dff_B_WiRQ99eB1_2;
	wire w_dff_B_suPLVpzt2_2;
	wire w_dff_B_XNBJe3SD3_2;
	wire w_dff_B_2Jcdb9cm1_2;
	wire w_dff_B_SxIBpEx52_2;
	wire w_dff_B_xp7BD0NP4_2;
	wire w_dff_B_fKc2By9A8_2;
	wire w_dff_B_x1gpd9tU7_2;
	wire w_dff_B_KWAnneZX5_2;
	wire w_dff_B_pK1bjzOe0_2;
	wire w_dff_B_qKvLM4Iq3_2;
	wire w_dff_B_nhlIYQLz9_2;
	wire w_dff_B_JB3bG6Ez7_2;
	wire w_dff_B_rE2btYBL6_2;
	wire w_dff_B_jamFC7LZ3_2;
	wire w_dff_B_4FG32wZ97_2;
	wire w_dff_B_sh2kcuiY3_2;
	wire w_dff_B_Cwv5OEyC3_2;
	wire w_dff_B_E6RTjQmc2_2;
	wire w_dff_B_b5uOftRa7_2;
	wire w_dff_B_m4B0bsaM0_2;
	wire w_dff_B_sJDrkbVR3_2;
	wire w_dff_B_IP2xz7gk6_2;
	wire w_dff_B_8fyuWS3C8_1;
	wire w_dff_B_CZ4lnBnU4_2;
	wire w_dff_B_uJTWmKKg9_2;
	wire w_dff_B_W8kdiqNn7_2;
	wire w_dff_B_DMpF30di2_2;
	wire w_dff_B_jObhIa4m8_2;
	wire w_dff_B_DkXtiUhh5_2;
	wire w_dff_B_3AZzWK5K9_2;
	wire w_dff_B_RB8EGyzc3_2;
	wire w_dff_B_2Rkc27738_2;
	wire w_dff_B_8bct5HR39_2;
	wire w_dff_B_TTeqG0FQ9_2;
	wire w_dff_B_blGsaODc0_2;
	wire w_dff_B_dC8F7YR52_2;
	wire w_dff_B_0CWn7SjJ2_2;
	wire w_dff_B_nwh0I2Wz3_2;
	wire w_dff_B_RUdayj0h1_2;
	wire w_dff_B_0taMoH0W1_2;
	wire w_dff_B_N06HOcfl0_2;
	wire w_dff_B_S6kSeQDQ7_2;
	wire w_dff_B_TnDkHids0_2;
	wire w_dff_B_QcMnnVQb5_2;
	wire w_dff_B_LZyd5xTg3_2;
	wire w_dff_B_jpyCYVHf7_2;
	wire w_dff_B_clxmQnR12_2;
	wire w_dff_B_tSSBfNa53_2;
	wire w_dff_B_EMA8cHjx2_2;
	wire w_dff_B_vPuxReyu7_2;
	wire w_dff_B_WpTXQUJm7_2;
	wire w_dff_B_ZwD6HCR57_2;
	wire w_dff_B_ywKQgdwa4_2;
	wire w_dff_B_j0Buq58s5_2;
	wire w_dff_B_yeqhcbgU8_2;
	wire w_dff_B_rRpQxRXk6_2;
	wire w_dff_B_CsyphyLd6_1;
	wire w_dff_B_hwIpHyGz5_2;
	wire w_dff_B_JaLNPF1R5_2;
	wire w_dff_B_Zoz5qMIX0_2;
	wire w_dff_B_3WYuB6Xe5_2;
	wire w_dff_B_O26byoBL3_2;
	wire w_dff_B_Wq22OHV66_2;
	wire w_dff_B_OMek1LYa7_2;
	wire w_dff_B_umbRiCSr6_2;
	wire w_dff_B_rLrmj8R86_2;
	wire w_dff_B_TGZvNaf38_2;
	wire w_dff_B_L6VddQaT1_2;
	wire w_dff_B_IeuTQqpa0_2;
	wire w_dff_B_bMmCb6Ng6_2;
	wire w_dff_B_3ObcaEG11_2;
	wire w_dff_B_1Nz5Iy0p0_2;
	wire w_dff_B_I8eRL6Ot3_2;
	wire w_dff_B_tlWbOF6S3_2;
	wire w_dff_B_JkJ5zbY76_2;
	wire w_dff_B_vJoA67bg3_2;
	wire w_dff_B_8zk7mE1u7_2;
	wire w_dff_B_4XKKqanO3_2;
	wire w_dff_B_4rGBuJul6_2;
	wire w_dff_B_bEemoxrx1_2;
	wire w_dff_B_xrQzQvAZ3_2;
	wire w_dff_B_gtHlNTOL7_2;
	wire w_dff_B_mwnWALYY4_2;
	wire w_dff_B_6rzBcZzE7_2;
	wire w_dff_B_eGjzVzzH4_2;
	wire w_dff_B_95Ba9HeD1_2;
	wire w_dff_B_Hv6YVCsr6_2;
	wire w_dff_B_LQq7XSgV1_1;
	wire w_dff_B_vcJIzG6e5_2;
	wire w_dff_B_KyAy0u7z2_2;
	wire w_dff_B_bwFVgsCd8_2;
	wire w_dff_B_ryv10emY7_2;
	wire w_dff_B_QLutS9cy4_2;
	wire w_dff_B_v9840jYK1_2;
	wire w_dff_B_BrCgUxQT1_2;
	wire w_dff_B_93aRqduI4_2;
	wire w_dff_B_PNnW47wB3_2;
	wire w_dff_B_rbEFlcNa3_2;
	wire w_dff_B_wvnIlnOQ6_2;
	wire w_dff_B_Dr87KwPU9_2;
	wire w_dff_B_iVVXmieo7_2;
	wire w_dff_B_XlvhNH716_2;
	wire w_dff_B_AgCiMPqe9_2;
	wire w_dff_B_7texvTvg8_2;
	wire w_dff_B_hYW46rO79_2;
	wire w_dff_B_tfZRLX5F1_2;
	wire w_dff_B_fdfRDlZi0_2;
	wire w_dff_B_KkekWbYD4_2;
	wire w_dff_B_DA453B0D7_2;
	wire w_dff_B_Tsr0aNow7_2;
	wire w_dff_B_bbOFfDPy5_2;
	wire w_dff_B_XGlQejHS2_2;
	wire w_dff_B_tpqpxOud6_2;
	wire w_dff_B_NgZUA2VO6_2;
	wire w_dff_B_a8DfgMyJ2_2;
	wire w_dff_B_VQ99M6Cp9_1;
	wire w_dff_B_fLOEm6OU5_2;
	wire w_dff_B_b7EgqpGf5_2;
	wire w_dff_B_IsKYsYA35_2;
	wire w_dff_B_mmaiWdOm9_2;
	wire w_dff_B_uifbmBo90_2;
	wire w_dff_B_VPp2sZDf3_2;
	wire w_dff_B_qSggmim50_2;
	wire w_dff_B_mvAoWqJI4_2;
	wire w_dff_B_QYgGxJNT9_2;
	wire w_dff_B_OjC2kcUA2_2;
	wire w_dff_B_ihnlVSrx3_2;
	wire w_dff_B_MMmXR79t3_2;
	wire w_dff_B_YZu4mbko4_2;
	wire w_dff_B_R2YHob0V1_2;
	wire w_dff_B_HGKn9FQW3_2;
	wire w_dff_B_KHbhU1An3_2;
	wire w_dff_B_dfrDS8QZ4_2;
	wire w_dff_B_VpsGrLNj7_2;
	wire w_dff_B_1iysCM1M1_2;
	wire w_dff_B_dbbJhbRE7_2;
	wire w_dff_B_m9jNYSza4_2;
	wire w_dff_B_fYo9iQxr0_2;
	wire w_dff_B_AJ278F735_2;
	wire w_dff_B_6UGA7hQZ1_2;
	wire w_dff_B_0oMYSq0L6_1;
	wire w_dff_B_loGNozgi9_2;
	wire w_dff_B_WwYCtl412_2;
	wire w_dff_B_0n1Jadz66_2;
	wire w_dff_B_PVehoIcG1_2;
	wire w_dff_B_vgegI7jV3_2;
	wire w_dff_B_1Pkxkatc6_2;
	wire w_dff_B_8YPRvzTG9_2;
	wire w_dff_B_5BL8usaY8_2;
	wire w_dff_B_5Wt5ibDr7_2;
	wire w_dff_B_HGp057y16_2;
	wire w_dff_B_N3HA4PbK2_2;
	wire w_dff_B_YP7WalGR7_2;
	wire w_dff_B_xXCczbKI4_2;
	wire w_dff_B_GG2LoV179_2;
	wire w_dff_B_7rTj1hxk0_2;
	wire w_dff_B_CU0GAnsS0_2;
	wire w_dff_B_lOPgQupd8_2;
	wire w_dff_B_r7yNn4561_2;
	wire w_dff_B_U5REUEV02_2;
	wire w_dff_B_nKiBMnI58_2;
	wire w_dff_B_OuUO3ksH5_2;
	wire w_dff_B_ze7CwRxD5_1;
	wire w_dff_B_t2qiqlq82_2;
	wire w_dff_B_hO8a1Kat6_2;
	wire w_dff_B_vIvEHoZA5_2;
	wire w_dff_B_M4VIBpVI8_2;
	wire w_dff_B_rie1OaCW6_2;
	wire w_dff_B_Q64ShAcO6_2;
	wire w_dff_B_0aDQFoDM4_2;
	wire w_dff_B_LU8Dum5u8_2;
	wire w_dff_B_cM3drlQI4_2;
	wire w_dff_B_Vl92Qsgo9_2;
	wire w_dff_B_uEBfFmQA5_2;
	wire w_dff_B_1JArMmMc1_2;
	wire w_dff_B_i5U1hvRO7_2;
	wire w_dff_B_SGnsI4oE7_2;
	wire w_dff_B_zEE62LWO5_2;
	wire w_dff_B_Y9rOaHPJ9_2;
	wire w_dff_B_XlNQGqbr8_2;
	wire w_dff_B_5kYk2Ixa5_2;
	wire w_dff_B_yZ1ZLZMX3_1;
	wire w_dff_B_9aoLueLy1_2;
	wire w_dff_B_NKCKydGn2_2;
	wire w_dff_B_EnS2MZHq4_2;
	wire w_dff_B_H4nkGOZq9_2;
	wire w_dff_B_I65d36uz4_2;
	wire w_dff_B_ODDEud1P6_2;
	wire w_dff_B_YOraFkZV4_2;
	wire w_dff_B_Do3QMKhj3_2;
	wire w_dff_B_5ngNZ9rE4_2;
	wire w_dff_B_MMv7rcA25_2;
	wire w_dff_B_PfO4DHBQ4_2;
	wire w_dff_B_LksThUh49_2;
	wire w_dff_B_o4GO084i3_2;
	wire w_dff_B_ZD8FogMh6_2;
	wire w_dff_B_YZpFnkvY4_2;
	wire w_dff_B_2TtZjgDR4_1;
	wire w_dff_B_Fjt8NB8M0_2;
	wire w_dff_B_u3Ye1c305_2;
	wire w_dff_B_gUTxaUXY9_2;
	wire w_dff_B_oevza0wB1_2;
	wire w_dff_B_a5k7dsn76_2;
	wire w_dff_B_jd9iXizh0_2;
	wire w_dff_B_Gg90a2hp3_2;
	wire w_dff_B_3CvsAI2d8_2;
	wire w_dff_B_yuFhykAK8_2;
	wire w_dff_B_7cHnDViy2_2;
	wire w_dff_B_hpCVcopu1_2;
	wire w_dff_B_N8xVdQVc1_2;
	wire w_dff_B_xDE2wZ4o5_1;
	wire w_dff_B_RVTKO89N5_2;
	wire w_dff_B_A9ghjFdp7_2;
	wire w_dff_B_WMQLPQZL3_2;
	wire w_dff_B_aFF7X2kQ6_2;
	wire w_dff_B_XU1FHgmb0_2;
	wire w_dff_B_DxLwwvlN7_2;
	wire w_dff_B_T9Gfyxhh1_2;
	wire w_dff_B_enx57Ify0_2;
	wire w_dff_B_NtmhkJ5H6_2;
	wire w_dff_B_s5WQ3C6t1_2;
	wire w_dff_B_HmdH1K3B2_2;
	wire w_dff_B_9yuZU2o59_1;
	wire w_dff_B_UTv53eIV5_1;
	wire w_dff_B_tWtgbXPF4_2;
	wire w_dff_B_ac57eWrJ6_2;
	wire w_dff_B_qT2GWI6i5_2;
	wire w_dff_B_tFhInTpS8_0;
	wire w_dff_A_Nr7FDlQy8_0;
	wire w_dff_A_ld5XHP2q6_0;
	wire w_dff_A_eYh6xHTD4_1;
	wire w_dff_A_iGOTVGdz2_1;
	wire w_dff_B_H4YrT5Qg7_2;
	wire w_dff_B_8u82OTEk1_1;
	wire w_dff_B_FGBf8jTf5_2;
	wire w_dff_B_U6B4oF6j0_2;
	wire w_dff_B_3fEIf1bE7_2;
	wire w_dff_B_yMlOjoPT8_2;
	wire w_dff_B_kCyg5rZc0_2;
	wire w_dff_B_ss9DrP9Y1_2;
	wire w_dff_B_dvk5yyze7_2;
	wire w_dff_B_4ywqs0yT2_2;
	wire w_dff_B_Gh7a08yD4_2;
	wire w_dff_B_JdaNaoCJ2_2;
	wire w_dff_B_pectrKqf5_2;
	wire w_dff_B_3R9HEZGO0_2;
	wire w_dff_B_9ygUsPbc1_2;
	wire w_dff_B_bOpPDq8M7_2;
	wire w_dff_B_Yj0muCWl6_2;
	wire w_dff_B_se3wxhWY6_2;
	wire w_dff_B_F3XBj8p07_2;
	wire w_dff_B_VVdkneR19_2;
	wire w_dff_B_LpBLNGRS6_2;
	wire w_dff_B_2VuZlde11_2;
	wire w_dff_B_nFCJ8jKP4_2;
	wire w_dff_B_KJT6IcWt6_2;
	wire w_dff_B_yRnuStW29_2;
	wire w_dff_B_f7ZKQCdD4_2;
	wire w_dff_B_cXNZhmIG1_2;
	wire w_dff_B_crvvGL4B9_2;
	wire w_dff_B_UhOpIEwD0_2;
	wire w_dff_B_ORNnKSAZ3_2;
	wire w_dff_B_O8kLOrDs2_2;
	wire w_dff_B_uDZeASMP8_2;
	wire w_dff_B_7PCcJPzQ8_2;
	wire w_dff_B_Wr61stAb9_2;
	wire w_dff_B_QiQR7aMu3_2;
	wire w_dff_B_i18PVtYj0_2;
	wire w_dff_B_CaZbuqti0_2;
	wire w_dff_B_KjIXxOAI4_2;
	wire w_dff_B_yNlJaCvY2_2;
	wire w_dff_B_0vT1vTWF3_2;
	wire w_dff_B_txootfBz2_2;
	wire w_dff_B_kNuXWdfu9_2;
	wire w_dff_B_detvEDeQ7_2;
	wire w_dff_B_sWByKdUo7_2;
	wire w_dff_B_2AclVfkZ8_2;
	wire w_dff_B_q3Jkis7o0_2;
	wire w_dff_B_Atz20Po82_2;
	wire w_dff_B_r2TRi9Mw7_2;
	wire w_dff_B_5fqpPpqw5_1;
	wire w_dff_B_QrfLMSFN7_2;
	wire w_dff_B_SwO2J2EG7_2;
	wire w_dff_B_Dhp19eWZ8_2;
	wire w_dff_B_oEFFDRTh8_2;
	wire w_dff_B_n4yAV2wC8_2;
	wire w_dff_B_3SGtO3pG8_2;
	wire w_dff_B_WPmYJb8g0_2;
	wire w_dff_B_vamdq46V0_2;
	wire w_dff_B_2c0lb1Bf7_2;
	wire w_dff_B_Sm94U7RC0_2;
	wire w_dff_B_tovPr3Gj6_2;
	wire w_dff_B_zPC9L6st9_2;
	wire w_dff_B_sTXdIzQA2_2;
	wire w_dff_B_x1NngZmO0_2;
	wire w_dff_B_azJUgKoO7_2;
	wire w_dff_B_u3P2LWv37_2;
	wire w_dff_B_cdPaMq575_2;
	wire w_dff_B_Zq5If9UR2_2;
	wire w_dff_B_w6kQEEtk9_2;
	wire w_dff_B_fbeGPNnm0_2;
	wire w_dff_B_BkEWtN9y7_2;
	wire w_dff_B_lvhUxNJ98_2;
	wire w_dff_B_ecqrKTUu2_2;
	wire w_dff_B_Y5dEumy19_2;
	wire w_dff_B_s2o6rmh26_2;
	wire w_dff_B_NMEG0RSD1_2;
	wire w_dff_B_JC3shGiu0_2;
	wire w_dff_B_pXr7CSBT4_2;
	wire w_dff_B_8w5qjcmb8_2;
	wire w_dff_B_z0CxYak16_2;
	wire w_dff_B_n8slCP0C6_2;
	wire w_dff_B_VT0uZWCC8_2;
	wire w_dff_B_bADfbBni1_2;
	wire w_dff_B_4BIGkTLY9_2;
	wire w_dff_B_4emyKrqa6_2;
	wire w_dff_B_m5RFnYi50_2;
	wire w_dff_B_HUgFLPur3_2;
	wire w_dff_B_a4usGJD99_2;
	wire w_dff_B_74qhYA3S4_2;
	wire w_dff_B_K35Yb9Sz9_2;
	wire w_dff_B_KK9cnNdY5_2;
	wire w_dff_B_qGDh7Zs29_2;
	wire w_dff_B_nhG2MuVO0_1;
	wire w_dff_B_a1J0J8zG7_2;
	wire w_dff_B_sLsiD19P3_2;
	wire w_dff_B_kZurIMWo1_2;
	wire w_dff_B_v1clK4ii3_2;
	wire w_dff_B_kbrYLWt37_2;
	wire w_dff_B_C1Pb4Yuh2_2;
	wire w_dff_B_Dut4g0gZ1_2;
	wire w_dff_B_MpKWRWAR2_2;
	wire w_dff_B_Fql4Qd7Y3_2;
	wire w_dff_B_HHxpagHl6_2;
	wire w_dff_B_PZ1KQNwm2_2;
	wire w_dff_B_nKl0y47p4_2;
	wire w_dff_B_OYBpVMMG4_2;
	wire w_dff_B_DhW66jAU8_2;
	wire w_dff_B_PKuxjvw20_2;
	wire w_dff_B_XO8h7PGg5_2;
	wire w_dff_B_6upL2GWj7_2;
	wire w_dff_B_GFhoQmhn0_2;
	wire w_dff_B_SY94yo6c3_2;
	wire w_dff_B_usDLdEv52_2;
	wire w_dff_B_sQZJRW9M8_2;
	wire w_dff_B_RS1zbws18_2;
	wire w_dff_B_oizmTqgH0_2;
	wire w_dff_B_7PiZW7l29_2;
	wire w_dff_B_A6TJtnUN1_2;
	wire w_dff_B_ohZEdczW6_2;
	wire w_dff_B_qy9MKSzC9_2;
	wire w_dff_B_iIQ3jMah6_2;
	wire w_dff_B_R38DuS625_2;
	wire w_dff_B_vIsaCBPL2_2;
	wire w_dff_B_cUbWS54X7_2;
	wire w_dff_B_eOyqHQmx1_2;
	wire w_dff_B_i0NGRoIy4_2;
	wire w_dff_B_QUAW3t0y8_2;
	wire w_dff_B_fLeIxoKr1_2;
	wire w_dff_B_hKsMYOUV6_2;
	wire w_dff_B_9uGbm21M2_2;
	wire w_dff_B_azQbmOOL5_2;
	wire w_dff_B_BHERS2qa9_2;
	wire w_dff_B_zf6t6t9G7_1;
	wire w_dff_B_dHAvEPUM8_2;
	wire w_dff_B_9vA585IV4_2;
	wire w_dff_B_5Ot79jrZ1_2;
	wire w_dff_B_bQt6pq1O5_2;
	wire w_dff_B_aCRvs3vO8_2;
	wire w_dff_B_OuMRJDx00_2;
	wire w_dff_B_7rnNunb37_2;
	wire w_dff_B_UNyA0LNQ6_2;
	wire w_dff_B_NkuPCib06_2;
	wire w_dff_B_HrWAqTVg2_2;
	wire w_dff_B_jr0H6M1h2_2;
	wire w_dff_B_SWrWulLa4_2;
	wire w_dff_B_Jct4dJkK5_2;
	wire w_dff_B_gvxPh2zu3_2;
	wire w_dff_B_irv6qS638_2;
	wire w_dff_B_77RqiY8q1_2;
	wire w_dff_B_4vLrbhgG4_2;
	wire w_dff_B_oshIgT4C9_2;
	wire w_dff_B_m3SBlrPt7_2;
	wire w_dff_B_tfumFg1C3_2;
	wire w_dff_B_wLCrObGZ6_2;
	wire w_dff_B_VVLKQ5Q39_2;
	wire w_dff_B_ezfXU9GF3_2;
	wire w_dff_B_cdb9Mvoj9_2;
	wire w_dff_B_lLLZcuUT7_2;
	wire w_dff_B_6O5EvuP08_2;
	wire w_dff_B_Ooj3M8kE1_2;
	wire w_dff_B_MKSnQWk41_2;
	wire w_dff_B_oLOudchR1_2;
	wire w_dff_B_zLTCYzRl5_2;
	wire w_dff_B_16exLBNQ7_2;
	wire w_dff_B_EdcHSJMl5_2;
	wire w_dff_B_shG9GEvp3_2;
	wire w_dff_B_27VPICdG5_2;
	wire w_dff_B_S6AkPJPj3_2;
	wire w_dff_B_YJTAuJ945_2;
	wire w_dff_B_vokYGC0b9_1;
	wire w_dff_B_Rs2hwzpB6_2;
	wire w_dff_B_aasmsvVd2_2;
	wire w_dff_B_4LFEAv2j1_2;
	wire w_dff_B_eaDDy6O16_2;
	wire w_dff_B_OcaGUfCW3_2;
	wire w_dff_B_PNv8s8b13_2;
	wire w_dff_B_vBZLomtJ0_2;
	wire w_dff_B_pFNvnAe62_2;
	wire w_dff_B_JH47gPyU9_2;
	wire w_dff_B_rV3xResR9_2;
	wire w_dff_B_63Ip9KMa2_2;
	wire w_dff_B_6M2EC8Sh4_2;
	wire w_dff_B_bcnpDTA37_2;
	wire w_dff_B_CZEdGSg04_2;
	wire w_dff_B_mm5R5TOt7_2;
	wire w_dff_B_60Pm7ex72_2;
	wire w_dff_B_PblsyD8d8_2;
	wire w_dff_B_RwT1Wr1B0_2;
	wire w_dff_B_vzNWISLk7_2;
	wire w_dff_B_3Kovejb60_2;
	wire w_dff_B_fYZ8xuDg6_2;
	wire w_dff_B_chM9taEi2_2;
	wire w_dff_B_74WmtdW34_2;
	wire w_dff_B_j07Wur1H8_2;
	wire w_dff_B_oqLzKfjo0_2;
	wire w_dff_B_AcLahKgS3_2;
	wire w_dff_B_t5uMJZv03_2;
	wire w_dff_B_3hXUBDKd9_2;
	wire w_dff_B_V6ganN2S2_2;
	wire w_dff_B_ZnWklMm30_2;
	wire w_dff_B_HPrd3aYp5_2;
	wire w_dff_B_FQxKZDL89_2;
	wire w_dff_B_Iax4cSnN7_2;
	wire w_dff_B_UmQpK0rO6_1;
	wire w_dff_B_FsbPAJqs4_2;
	wire w_dff_B_hr2bwteo6_2;
	wire w_dff_B_SPLLnP7V4_2;
	wire w_dff_B_ZQK7VYsx0_2;
	wire w_dff_B_eP6flCHu8_2;
	wire w_dff_B_brZIFypa5_2;
	wire w_dff_B_pqV4ZWSR7_2;
	wire w_dff_B_UYsBVN7x8_2;
	wire w_dff_B_tBOkJJb40_2;
	wire w_dff_B_nsVhCZI74_2;
	wire w_dff_B_cuijBt0D2_2;
	wire w_dff_B_9wj8SFYG0_2;
	wire w_dff_B_tsTS65vP0_2;
	wire w_dff_B_9Kcyb6XJ9_2;
	wire w_dff_B_9PupgfsD7_2;
	wire w_dff_B_6XqStstz9_2;
	wire w_dff_B_6eOq1zfV8_2;
	wire w_dff_B_ILwT88TU8_2;
	wire w_dff_B_BUWLskyo8_2;
	wire w_dff_B_N4sZZfxb6_2;
	wire w_dff_B_eqDd9iGy1_2;
	wire w_dff_B_wpPzMh8I8_2;
	wire w_dff_B_c7gFdwpw1_2;
	wire w_dff_B_cIlPVjOn5_2;
	wire w_dff_B_NqV9IsLF5_2;
	wire w_dff_B_Rb0pOu6w7_2;
	wire w_dff_B_662tQZJI7_2;
	wire w_dff_B_kSVCW75S1_2;
	wire w_dff_B_BJnENFj11_2;
	wire w_dff_B_iPNammup2_2;
	wire w_dff_B_kV5BDMjF1_1;
	wire w_dff_B_XhDtq3AJ2_2;
	wire w_dff_B_OtLSsN8s5_2;
	wire w_dff_B_bnGijKmp3_2;
	wire w_dff_B_hG63Xueq7_2;
	wire w_dff_B_n7O1Vi9l0_2;
	wire w_dff_B_EFcVe6XA3_2;
	wire w_dff_B_gUOyplqD7_2;
	wire w_dff_B_fOUSJ79E6_2;
	wire w_dff_B_C8o3RLos2_2;
	wire w_dff_B_pFQjw1tg7_2;
	wire w_dff_B_FI3zd4kB1_2;
	wire w_dff_B_2OInZIqZ2_2;
	wire w_dff_B_UZfuMZFs9_2;
	wire w_dff_B_7JcPBHQe5_2;
	wire w_dff_B_ndH0dVsQ9_2;
	wire w_dff_B_pkbBsHLO6_2;
	wire w_dff_B_NnntY5257_2;
	wire w_dff_B_iOERsrR15_2;
	wire w_dff_B_XxpYyPVq8_2;
	wire w_dff_B_Q5tekKKe3_2;
	wire w_dff_B_vLguwKsV5_2;
	wire w_dff_B_0dbO5Wv47_2;
	wire w_dff_B_OtmVuPkN3_2;
	wire w_dff_B_zByO5G0a4_2;
	wire w_dff_B_7Pig3tyK4_2;
	wire w_dff_B_JryGpri68_2;
	wire w_dff_B_Plxwei5y9_2;
	wire w_dff_B_OjcRlY2h2_1;
	wire w_dff_B_HPLnmYZ77_2;
	wire w_dff_B_LbOgLdUB8_2;
	wire w_dff_B_8NvYTmhn2_2;
	wire w_dff_B_MEBeBxjM5_2;
	wire w_dff_B_IGindAYx2_2;
	wire w_dff_B_ZQPs9dvB0_2;
	wire w_dff_B_ZCpSSidV1_2;
	wire w_dff_B_jXxu9ANi9_2;
	wire w_dff_B_tu67hxLv5_2;
	wire w_dff_B_0blAYzrs3_2;
	wire w_dff_B_TbBUV0R14_2;
	wire w_dff_B_JDREr97s5_2;
	wire w_dff_B_yb7PB9Q66_2;
	wire w_dff_B_nb3SKiOT1_2;
	wire w_dff_B_WWQgLknE4_2;
	wire w_dff_B_3O4752CT8_2;
	wire w_dff_B_vQ44mGwc6_2;
	wire w_dff_B_raAU1QSt2_2;
	wire w_dff_B_mvcsrnVc6_2;
	wire w_dff_B_TNAedXlp4_2;
	wire w_dff_B_UNstYPRl4_2;
	wire w_dff_B_86jlqXc21_2;
	wire w_dff_B_tSTxillR3_2;
	wire w_dff_B_hTlA5sbm7_2;
	wire w_dff_B_4uKjXcCu3_1;
	wire w_dff_B_fQlxMl3S2_2;
	wire w_dff_B_vOfmXFxe6_2;
	wire w_dff_B_Dnm3OYAp9_2;
	wire w_dff_B_6BoHQNdw7_2;
	wire w_dff_B_8skwEj4r5_2;
	wire w_dff_B_SDPVJy5z0_2;
	wire w_dff_B_1eEa4Tww7_2;
	wire w_dff_B_5oxYSuVg4_2;
	wire w_dff_B_qVWTOqfh8_2;
	wire w_dff_B_ebnHM4xV7_2;
	wire w_dff_B_NnQfzU9z1_2;
	wire w_dff_B_IozRSbbz6_2;
	wire w_dff_B_vM7YJ0Xz1_2;
	wire w_dff_B_qD9Fs3SU4_2;
	wire w_dff_B_xmQi2xox5_2;
	wire w_dff_B_jBhYpXq06_2;
	wire w_dff_B_CAA55B1Q4_2;
	wire w_dff_B_abYapm3v1_2;
	wire w_dff_B_x7NgL6XT6_2;
	wire w_dff_B_f5N2DkNH4_2;
	wire w_dff_B_D286X2Hh9_2;
	wire w_dff_B_UxsF3NTc2_1;
	wire w_dff_B_hX83ipm33_2;
	wire w_dff_B_zHvMk9Xz7_2;
	wire w_dff_B_HWcn8jjT1_2;
	wire w_dff_B_mGgKSy1w6_2;
	wire w_dff_B_LkwT9Bz25_2;
	wire w_dff_B_UygJsp3C1_2;
	wire w_dff_B_Fj9SQ95y6_2;
	wire w_dff_B_OOIce2499_2;
	wire w_dff_B_fCJYw80P6_2;
	wire w_dff_B_3bHjyah09_2;
	wire w_dff_B_Bz4Qlem84_2;
	wire w_dff_B_5G53VeFP1_2;
	wire w_dff_B_ydf0zOwQ6_2;
	wire w_dff_B_Mr9PeNBM7_2;
	wire w_dff_B_mijPNv5Q7_2;
	wire w_dff_B_EfAza7EV0_2;
	wire w_dff_B_QFBFxzKh3_2;
	wire w_dff_B_FYrpa1pl8_2;
	wire w_dff_B_0SQLVANx9_1;
	wire w_dff_B_JMyW1ypF9_2;
	wire w_dff_B_ZabHqtev9_2;
	wire w_dff_B_IgmttBZF3_2;
	wire w_dff_B_kxWji1ZO6_2;
	wire w_dff_B_d0AN3yjj9_2;
	wire w_dff_B_Yyo1N9A11_2;
	wire w_dff_B_vNMxwU1F8_2;
	wire w_dff_B_WhY8Jqys4_2;
	wire w_dff_B_E0b8Qx8l9_2;
	wire w_dff_B_FGUSWCTU2_2;
	wire w_dff_B_wZjoefnz4_2;
	wire w_dff_B_DLMpgKeL7_2;
	wire w_dff_B_KgWTyaJP3_2;
	wire w_dff_B_VRnjLZMF3_2;
	wire w_dff_B_1GKvZS0y0_2;
	wire w_dff_B_L9dAiNeY6_1;
	wire w_dff_B_2hQyrjfp5_2;
	wire w_dff_B_BOZk9Qht4_2;
	wire w_dff_B_r1xfYZN53_2;
	wire w_dff_B_EPQRGGMb7_2;
	wire w_dff_B_iIKiHArP0_2;
	wire w_dff_B_Eu9Ud1cb9_2;
	wire w_dff_B_kH1awpSJ2_2;
	wire w_dff_B_epbDVz3U0_2;
	wire w_dff_B_KZTDu68j0_2;
	wire w_dff_B_v20WeeIt3_2;
	wire w_dff_B_RmOrkIc96_2;
	wire w_dff_B_6vOacekQ0_2;
	wire w_dff_B_fhsB5pI32_1;
	wire w_dff_B_j6r1Pr0z6_2;
	wire w_dff_B_RyfUBfVm0_2;
	wire w_dff_B_ZW9y5cSy0_2;
	wire w_dff_B_zvjJeL4G4_2;
	wire w_dff_B_oPHvr82C4_2;
	wire w_dff_B_Gng1ttnp6_2;
	wire w_dff_B_IDqVQHuX0_2;
	wire w_dff_B_SF8nTlbT9_2;
	wire w_dff_B_1peuGQj02_2;
	wire w_dff_B_ioxh8fVC2_2;
	wire w_dff_B_7qNLUpmv4_2;
	wire w_dff_B_4LAuJUSU0_1;
	wire w_dff_B_Zdg8hQQA3_1;
	wire w_dff_B_ESJgNDMp1_2;
	wire w_dff_B_L6eWh6e09_2;
	wire w_dff_B_7ZZLxOsm6_2;
	wire w_dff_B_pZTOoJE89_0;
	wire w_dff_A_5Se624DU4_0;
	wire w_dff_A_tI7GeNyK3_0;
	wire w_dff_A_ZWzEZO8B7_1;
	wire w_dff_A_4MM8phz66_1;
	wire w_dff_B_GwYof2122_1;
	wire w_dff_A_SwQ6ri8m3_1;
	wire w_dff_B_2BO5H3Fh3_1;
	wire w_dff_B_RcXJoA6M0_2;
	wire w_dff_B_Y2oKoKr14_2;
	wire w_dff_B_AqPVFHW88_2;
	wire w_dff_B_LXSgQJGn9_2;
	wire w_dff_B_tnyuM3JP5_2;
	wire w_dff_B_EsATly1H6_2;
	wire w_dff_B_drNmJrFC1_2;
	wire w_dff_B_IZfbzlGw3_2;
	wire w_dff_B_kwFoYC738_2;
	wire w_dff_B_48rGiQOT0_2;
	wire w_dff_B_SJPeioDR3_2;
	wire w_dff_B_lFPka0Mg0_2;
	wire w_dff_B_q4jIGpo08_2;
	wire w_dff_B_6I0723fN9_2;
	wire w_dff_B_4Rmj2au51_2;
	wire w_dff_B_QsbgupvY5_2;
	wire w_dff_B_gR31hLuU8_2;
	wire w_dff_B_ayIruosr3_2;
	wire w_dff_B_FR4NXnEc2_2;
	wire w_dff_B_U8P0ZI8H6_2;
	wire w_dff_B_3uuSu37e9_2;
	wire w_dff_B_pJgnBA9L0_2;
	wire w_dff_B_oMVFEaJZ8_2;
	wire w_dff_B_SNcH6jEJ1_2;
	wire w_dff_B_Y9glgvmM9_2;
	wire w_dff_B_FSEjjpyd0_2;
	wire w_dff_B_1crG85sG9_2;
	wire w_dff_B_vTiA19Pk2_2;
	wire w_dff_B_Lyc5LJAo0_2;
	wire w_dff_B_bGXVEpuy0_2;
	wire w_dff_B_mSs1jPUu0_2;
	wire w_dff_B_Pku4wRHZ5_2;
	wire w_dff_B_B7nL4GdN8_2;
	wire w_dff_B_KGXfH1jC9_2;
	wire w_dff_B_J2KmmILp8_2;
	wire w_dff_B_OJ7Z7NdO4_2;
	wire w_dff_B_4gXtPzDy4_2;
	wire w_dff_B_JGdoBNXQ8_2;
	wire w_dff_B_VD9mQd8f7_2;
	wire w_dff_B_Ch4NS9AK4_2;
	wire w_dff_B_J1tycnE23_2;
	wire w_dff_B_aVyGAD361_2;
	wire w_dff_B_7v498nzy0_2;
	wire w_dff_B_JaHyIaEv7_2;
	wire w_dff_B_0Z2jdXNz8_2;
	wire w_dff_B_nBxfy3Zo3_2;
	wire w_dff_B_toABSUla3_2;
	wire w_dff_B_fL374ioq5_1;
	wire w_dff_B_srz84Pgv4_2;
	wire w_dff_B_sUGcgf2X2_2;
	wire w_dff_B_RUO0MwKQ6_2;
	wire w_dff_B_5CxXe5pG9_2;
	wire w_dff_B_50FqWL0Y6_2;
	wire w_dff_B_ArT0Qvck4_2;
	wire w_dff_B_QYaoqqG31_2;
	wire w_dff_B_bRblvbew7_2;
	wire w_dff_B_WLVMwxOw3_2;
	wire w_dff_B_vqFZ7Nlo6_2;
	wire w_dff_B_azEYAeet3_2;
	wire w_dff_B_6GDNLp3L0_2;
	wire w_dff_B_GR1mAU6h5_2;
	wire w_dff_B_iG84c0cQ4_2;
	wire w_dff_B_c0IoGkQP4_2;
	wire w_dff_B_gmBvsdYM9_2;
	wire w_dff_B_NrddrdD48_2;
	wire w_dff_B_qbGeRZxD1_2;
	wire w_dff_B_2ser7ZdF1_2;
	wire w_dff_B_47goirtf3_2;
	wire w_dff_B_D7XGDyVJ9_2;
	wire w_dff_B_sHbW1fKC7_2;
	wire w_dff_B_0Vhg79P96_2;
	wire w_dff_B_hvuTvXpA6_2;
	wire w_dff_B_5xX9sl2J5_2;
	wire w_dff_B_NQN0w1Pi1_2;
	wire w_dff_B_Ch0jz0Lk7_2;
	wire w_dff_B_6RVLTVQF5_2;
	wire w_dff_B_VKIDSFkq0_2;
	wire w_dff_B_6WOtqA6l9_2;
	wire w_dff_B_EUwzOq7b3_2;
	wire w_dff_B_YLDpHNXV0_2;
	wire w_dff_B_36NqWeYd2_2;
	wire w_dff_B_2brQbtMX9_2;
	wire w_dff_B_DqxQL4XO5_2;
	wire w_dff_B_NniZN1Ep7_2;
	wire w_dff_B_mgg01KfN9_2;
	wire w_dff_B_O9TiFwU31_2;
	wire w_dff_B_KzSalANb9_2;
	wire w_dff_B_Z8fkM5Ii2_2;
	wire w_dff_B_IPbenLDB9_2;
	wire w_dff_B_7sCSoUGO2_2;
	wire w_dff_B_JeVevLGF2_2;
	wire w_dff_B_72FCd2WI3_1;
	wire w_dff_B_0Vkd3RTi3_2;
	wire w_dff_B_viszoCbb1_2;
	wire w_dff_B_HKpayDrq0_2;
	wire w_dff_B_E9oVdWO76_2;
	wire w_dff_B_jhOmsjKU5_2;
	wire w_dff_B_xtnw1jPq3_2;
	wire w_dff_B_vMVUCDk53_2;
	wire w_dff_B_LLlFAXGO4_2;
	wire w_dff_B_WSTci83g3_2;
	wire w_dff_B_Sy19B0WV3_2;
	wire w_dff_B_hSeXNY4M3_2;
	wire w_dff_B_knrWhgjB0_2;
	wire w_dff_B_AlE2HCrZ7_2;
	wire w_dff_B_pUKBjtUL4_2;
	wire w_dff_B_x9Vc4eVj3_2;
	wire w_dff_B_YlLyWT2v8_2;
	wire w_dff_B_hE1A2bxz0_2;
	wire w_dff_B_RViGyZXN7_2;
	wire w_dff_B_js2biHo04_2;
	wire w_dff_B_WXYXMVMO7_2;
	wire w_dff_B_P71syNyq0_2;
	wire w_dff_B_3ubAaHD18_2;
	wire w_dff_B_ZKTx0qP55_2;
	wire w_dff_B_NRRn0mRd2_2;
	wire w_dff_B_qGaMJt2o9_2;
	wire w_dff_B_UOKfX48y1_2;
	wire w_dff_B_UAhTtrPE9_2;
	wire w_dff_B_qp6leGgL9_2;
	wire w_dff_B_Fun1EjNk6_2;
	wire w_dff_B_9F7rfMuK1_2;
	wire w_dff_B_N588Bo4B8_2;
	wire w_dff_B_jIJU7zvh7_2;
	wire w_dff_B_ywrMII1O9_2;
	wire w_dff_B_HHFWSoPB6_2;
	wire w_dff_B_FCpTu1Oa8_2;
	wire w_dff_B_Xjo0NHRN6_2;
	wire w_dff_B_6gaVyu1c2_2;
	wire w_dff_B_T9xSZq4u2_2;
	wire w_dff_B_rtoEWXzK4_1;
	wire w_dff_B_gnbereKi1_2;
	wire w_dff_B_4sCXKAMt1_2;
	wire w_dff_B_6isl9lQp4_2;
	wire w_dff_B_Hdl40UF99_2;
	wire w_dff_B_k3FqWsEE3_2;
	wire w_dff_B_iWKtQyWh8_2;
	wire w_dff_B_nvr54PpG3_2;
	wire w_dff_B_AK8tEOvm0_2;
	wire w_dff_B_1R9eaqrL3_2;
	wire w_dff_B_AtGAz6sJ3_2;
	wire w_dff_B_bxWflXCE9_2;
	wire w_dff_B_SIXSQ67O1_2;
	wire w_dff_B_7fkhM7wJ7_2;
	wire w_dff_B_zYeiN5JJ3_2;
	wire w_dff_B_JMkfEVJD1_2;
	wire w_dff_B_Tzx18ChG4_2;
	wire w_dff_B_yVYF2ret0_2;
	wire w_dff_B_VbsMSVfW1_2;
	wire w_dff_B_GRIBojrQ9_2;
	wire w_dff_B_ufNGh5Nz9_2;
	wire w_dff_B_DDVDSGGr2_2;
	wire w_dff_B_mNTMWGwj0_2;
	wire w_dff_B_VTye8jUV5_2;
	wire w_dff_B_UOQW4Sx61_2;
	wire w_dff_B_AXAewekX7_2;
	wire w_dff_B_I64BCFFe1_2;
	wire w_dff_B_GV3oyR2n5_2;
	wire w_dff_B_mjDJMCsb6_2;
	wire w_dff_B_8bAUqhY71_2;
	wire w_dff_B_WnYZ6jln3_2;
	wire w_dff_B_5mHy322U6_2;
	wire w_dff_B_w2IKrN7g5_2;
	wire w_dff_B_Qx7mxZdT6_2;
	wire w_dff_B_V8sIV8sd4_2;
	wire w_dff_B_YklFauZj3_2;
	wire w_dff_B_p7AWjSaB0_2;
	wire w_dff_B_ISJUd31I5_1;
	wire w_dff_B_ojx5wQ788_2;
	wire w_dff_B_QrGb6vKY1_2;
	wire w_dff_B_XmWNjiDD2_2;
	wire w_dff_B_U0fFuZLV2_2;
	wire w_dff_B_OcXYIF8E9_2;
	wire w_dff_B_gsfkJpD56_2;
	wire w_dff_B_lX7IsoW62_2;
	wire w_dff_B_R6nnz4UU4_2;
	wire w_dff_B_iseOWATe5_2;
	wire w_dff_B_ekQc6uMI0_2;
	wire w_dff_B_Tg2ton5F5_2;
	wire w_dff_B_NC6bMZWi2_2;
	wire w_dff_B_OV4Ev9ke2_2;
	wire w_dff_B_is4k58l98_2;
	wire w_dff_B_lyz9BWDG1_2;
	wire w_dff_B_guYPLWXn1_2;
	wire w_dff_B_mCemIItI9_2;
	wire w_dff_B_TqwFgypW8_2;
	wire w_dff_B_xYAQw4AV9_2;
	wire w_dff_B_EdqLmb3R3_2;
	wire w_dff_B_wCYtV0fA5_2;
	wire w_dff_B_C2u7cuHN4_2;
	wire w_dff_B_57zDsbaF2_2;
	wire w_dff_B_jHyEaw602_2;
	wire w_dff_B_EGWOWf9O9_2;
	wire w_dff_B_3Q829Jkz3_2;
	wire w_dff_B_sJTrjs2W8_2;
	wire w_dff_B_tCRWd8Nn7_2;
	wire w_dff_B_lgAIjsaz4_2;
	wire w_dff_B_gFPDvHSl5_2;
	wire w_dff_B_XWMtnGVA1_2;
	wire w_dff_B_b6jgOv2c9_2;
	wire w_dff_B_OMXvXjla2_2;
	wire w_dff_B_Np1v8xsj0_1;
	wire w_dff_B_r9gpkzOX2_2;
	wire w_dff_B_Q5FUyK8T8_2;
	wire w_dff_B_WR9kmS2X1_2;
	wire w_dff_B_1DoWVFXC1_2;
	wire w_dff_B_ZAbB7ElF1_2;
	wire w_dff_B_DPWgG65B2_2;
	wire w_dff_B_d4tDt8xY2_2;
	wire w_dff_B_SE9M4N407_2;
	wire w_dff_B_4KpCWajW6_2;
	wire w_dff_B_7rAnPWkD7_2;
	wire w_dff_B_OAgzgMeN7_2;
	wire w_dff_B_f3bO6ym16_2;
	wire w_dff_B_HesHG1wa0_2;
	wire w_dff_B_n536rLtD1_2;
	wire w_dff_B_6lxU23xG7_2;
	wire w_dff_B_oK34vapg7_2;
	wire w_dff_B_RIE4rCTD5_2;
	wire w_dff_B_tP5Jx9bR0_2;
	wire w_dff_B_jY14pEFG1_2;
	wire w_dff_B_MnnwXFB70_2;
	wire w_dff_B_3EnhQxlt8_2;
	wire w_dff_B_exRvzMEK2_2;
	wire w_dff_B_yAKnvj3u6_2;
	wire w_dff_B_j4vFqJ064_2;
	wire w_dff_B_yJX6VZx83_2;
	wire w_dff_B_GWUwXBzq6_2;
	wire w_dff_B_YFRCnf3a8_2;
	wire w_dff_B_8IqsvRsL8_2;
	wire w_dff_B_FIqkKil95_2;
	wire w_dff_B_QCqWFUuj5_2;
	wire w_dff_B_sVmjXq6O1_1;
	wire w_dff_B_EEabGscb2_2;
	wire w_dff_B_C5w2kazg8_2;
	wire w_dff_B_r9Sv5kHl7_2;
	wire w_dff_B_uGOE5r0T1_2;
	wire w_dff_B_9TwJOURK2_2;
	wire w_dff_B_TfOF2y5w2_2;
	wire w_dff_B_6IR98p932_2;
	wire w_dff_B_btSoseQP4_2;
	wire w_dff_B_fS0yraMI8_2;
	wire w_dff_B_scyRMOS63_2;
	wire w_dff_B_pVniVI5P7_2;
	wire w_dff_B_9uNclzfI9_2;
	wire w_dff_B_c3VBUoBz3_2;
	wire w_dff_B_4ifoD7h11_2;
	wire w_dff_B_hlolFbYN3_2;
	wire w_dff_B_GcVyUEG90_2;
	wire w_dff_B_IVrARRAJ7_2;
	wire w_dff_B_7JJpx3z64_2;
	wire w_dff_B_Jewm9tFG1_2;
	wire w_dff_B_p9A0L6m08_2;
	wire w_dff_B_lHK1nEr31_2;
	wire w_dff_B_xgDKfvmL6_2;
	wire w_dff_B_9SBAGRw60_2;
	wire w_dff_B_77LkU9Lp6_2;
	wire w_dff_B_oo3hJmBa6_2;
	wire w_dff_B_lI9bCXDS3_2;
	wire w_dff_B_vcCq38sD8_2;
	wire w_dff_B_D0MLO62s7_1;
	wire w_dff_B_lDD5EwiP7_2;
	wire w_dff_B_Hdwz1ovf6_2;
	wire w_dff_B_jqabLlTY0_2;
	wire w_dff_B_uKePzSI57_2;
	wire w_dff_B_gaOYESsH8_2;
	wire w_dff_B_CniT0wFX8_2;
	wire w_dff_B_dHg9dOE06_2;
	wire w_dff_B_NIVvBHeG0_2;
	wire w_dff_B_VzNCio8K6_2;
	wire w_dff_B_8w6j5v7y6_2;
	wire w_dff_B_pcyUuP953_2;
	wire w_dff_B_0Hiugs2T1_2;
	wire w_dff_B_BAdALqCA6_2;
	wire w_dff_B_mSwIxkXj7_2;
	wire w_dff_B_T0QRnaFX5_2;
	wire w_dff_B_GNuTaNYm0_2;
	wire w_dff_B_Dy29BoGg8_2;
	wire w_dff_B_tSwhzLp33_2;
	wire w_dff_B_gGSt85UG0_2;
	wire w_dff_B_YYxGgZYu9_2;
	wire w_dff_B_d5I3Ey5t8_2;
	wire w_dff_B_QuqzS3fK1_2;
	wire w_dff_B_mNza9tcW4_2;
	wire w_dff_B_WUYVu1hl2_2;
	wire w_dff_B_QMF8uRl06_1;
	wire w_dff_B_GWeOCnPO4_2;
	wire w_dff_B_dp9fFCs86_2;
	wire w_dff_B_VCj82tDn3_2;
	wire w_dff_B_vR181oxi7_2;
	wire w_dff_B_IxfaIcaT8_2;
	wire w_dff_B_IztkZPXG7_2;
	wire w_dff_B_hrt4Mc5x8_2;
	wire w_dff_B_8G0zxng01_2;
	wire w_dff_B_iSS9SgOM1_2;
	wire w_dff_B_61yb0ejX0_2;
	wire w_dff_B_DyhUzHgK1_2;
	wire w_dff_B_Q1Z70QoM6_2;
	wire w_dff_B_rKgbTX9Z3_2;
	wire w_dff_B_ZyRBvNaZ5_2;
	wire w_dff_B_JiEXtOrC9_2;
	wire w_dff_B_Ac5JdQf82_2;
	wire w_dff_B_QPIfgRm07_2;
	wire w_dff_B_dvVVJkmv8_2;
	wire w_dff_B_9c7T0okH9_2;
	wire w_dff_B_652yf0Nx1_2;
	wire w_dff_B_NeEOwLOI0_2;
	wire w_dff_B_Fipv8Gnp4_1;
	wire w_dff_B_D7jdRNo73_2;
	wire w_dff_B_BtA0HKAD4_2;
	wire w_dff_B_AhycjzWL7_2;
	wire w_dff_B_3xKiqqXz9_2;
	wire w_dff_B_T7FWyf9u6_2;
	wire w_dff_B_OU22KPS90_2;
	wire w_dff_B_RjM9ejhg4_2;
	wire w_dff_B_gab97HyR4_2;
	wire w_dff_B_rMKqRuTO1_2;
	wire w_dff_B_dSkZkfJE4_2;
	wire w_dff_B_sN3aDqCS2_2;
	wire w_dff_B_ncNNF4w89_2;
	wire w_dff_B_mNnMG2Nw2_2;
	wire w_dff_B_Nu24rtER5_2;
	wire w_dff_B_EH87Q9Ja2_2;
	wire w_dff_B_v7n9ZdN78_2;
	wire w_dff_B_vel3G9qh4_2;
	wire w_dff_B_BygthE7M4_2;
	wire w_dff_B_8eTRNjEg9_1;
	wire w_dff_B_dSdzBKzL6_2;
	wire w_dff_B_kRD1cGHm0_2;
	wire w_dff_B_XSB0ImkT2_2;
	wire w_dff_B_XFmF0o247_2;
	wire w_dff_B_PD1NDFcd8_2;
	wire w_dff_B_NB5zcMHp8_2;
	wire w_dff_B_LoTM9iGp8_2;
	wire w_dff_B_vh1z7EQf4_2;
	wire w_dff_B_zQxCkmZz4_2;
	wire w_dff_B_f8lY0Vet6_2;
	wire w_dff_B_dx4pguYu7_2;
	wire w_dff_B_QmuKa4eK6_2;
	wire w_dff_B_7X7O8SjT0_2;
	wire w_dff_B_y521lsx49_2;
	wire w_dff_B_nNHk4TPi9_2;
	wire w_dff_B_ls7eEVDF7_1;
	wire w_dff_B_zKkPmLf05_2;
	wire w_dff_B_TqMtYgbm1_2;
	wire w_dff_B_jE18dZpw0_2;
	wire w_dff_B_DJpvfd7x3_2;
	wire w_dff_B_RhTWUUQC2_2;
	wire w_dff_B_lUQaqNA31_2;
	wire w_dff_B_jhO1V4YD3_2;
	wire w_dff_B_OmTWrffi8_2;
	wire w_dff_B_6XF6CHzP5_2;
	wire w_dff_B_AZbtr5c57_2;
	wire w_dff_B_L4nzzlCr2_2;
	wire w_dff_B_t4bNrN1L3_2;
	wire w_dff_B_MeaEWRaU7_1;
	wire w_dff_B_BHp6WDKG1_2;
	wire w_dff_B_DSmInTRM0_2;
	wire w_dff_B_3QYMA24v9_2;
	wire w_dff_B_SFGCOXC16_2;
	wire w_dff_B_PjFtCOgg4_2;
	wire w_dff_B_gWzcO45F1_2;
	wire w_dff_B_e3dMIBCj6_2;
	wire w_dff_B_KiS2yLUk1_2;
	wire w_dff_B_5fbQ0Tdx8_2;
	wire w_dff_B_FXkMh77Y8_2;
	wire w_dff_B_BJLQn1AZ7_2;
	wire w_dff_B_HdovCmk45_1;
	wire w_dff_B_Q8Jhx20V3_1;
	wire w_dff_B_uImFXF9W3_2;
	wire w_dff_B_Mzhg2ssD0_2;
	wire w_dff_B_ts3WuSzZ2_2;
	wire w_dff_B_vPj7a03l5_0;
	wire w_dff_A_KX7Rd5572_0;
	wire w_dff_A_rWc83jMO0_0;
	wire w_dff_A_gy46G8l43_1;
	wire w_dff_A_mOLit72c0_1;
	wire w_dff_B_s9lPq6nu2_1;
	wire w_dff_A_xWpozIyr6_1;
	wire w_dff_B_iOR8SBie2_1;
	wire w_dff_B_xvidG6BS0_2;
	wire w_dff_B_H2JOajln6_2;
	wire w_dff_B_Ycn68z6x2_2;
	wire w_dff_B_Qkicp0Nj0_2;
	wire w_dff_B_zlxqnU5T9_2;
	wire w_dff_B_mSDuYZpA9_2;
	wire w_dff_B_vmDLUHHK1_2;
	wire w_dff_B_eHd2FTqC3_2;
	wire w_dff_B_uBOGlqrS6_2;
	wire w_dff_B_gyLmnItY4_2;
	wire w_dff_B_A0NbFXRA3_2;
	wire w_dff_B_KZ3Pl0a95_2;
	wire w_dff_B_68pFLTaF9_2;
	wire w_dff_B_Nblkd6oV4_2;
	wire w_dff_B_msA6pmMP5_2;
	wire w_dff_B_OTPIfpTj9_2;
	wire w_dff_B_ThheJh362_2;
	wire w_dff_B_78wLyOoW3_2;
	wire w_dff_B_K1WphjVx7_2;
	wire w_dff_B_y3jsG4hi1_2;
	wire w_dff_B_wBCu0QuX0_2;
	wire w_dff_B_k9OXH5N45_2;
	wire w_dff_B_mcAs9FME2_2;
	wire w_dff_B_xzlCFREP8_2;
	wire w_dff_B_EFUzlIud0_2;
	wire w_dff_B_0yo6G0Im4_2;
	wire w_dff_B_KIwlVoas2_2;
	wire w_dff_B_usAQ4Qhc7_2;
	wire w_dff_B_QKoOKo823_2;
	wire w_dff_B_D7HvH2q07_2;
	wire w_dff_B_iZ8Cg2jB2_2;
	wire w_dff_B_XrxrqQa70_2;
	wire w_dff_B_AimAZ4rY5_2;
	wire w_dff_B_0mGKjRwK7_2;
	wire w_dff_B_SLqgLeUz6_2;
	wire w_dff_B_0Notq8cF1_2;
	wire w_dff_B_cmmxr5wm9_2;
	wire w_dff_B_HsDwihJM1_2;
	wire w_dff_B_kU29M0Bi9_2;
	wire w_dff_B_OO6lC5Ma8_2;
	wire w_dff_B_u8os5wxt0_2;
	wire w_dff_B_9aw1YUF01_2;
	wire w_dff_B_H41Oumqr2_2;
	wire w_dff_B_MLozTtSE3_2;
	wire w_dff_B_u2iNC7Yd9_2;
	wire w_dff_B_lFhYoAov1_2;
	wire w_dff_B_FFxwMcAg2_2;
	wire w_dff_B_4Kjf9Xzu5_2;
	wire w_dff_B_AUJVVuZs7_2;
	wire w_dff_B_rhnCP9QY2_1;
	wire w_dff_B_C7LHpqBI3_2;
	wire w_dff_B_UeWfbcrz7_2;
	wire w_dff_B_n4tpqdkJ5_2;
	wire w_dff_B_G7YogIVE9_2;
	wire w_dff_B_J8LjVr9Z2_2;
	wire w_dff_B_Y0KJbX4N0_2;
	wire w_dff_B_4qNiEXOt8_2;
	wire w_dff_B_9kFeaxVf5_2;
	wire w_dff_B_HsptdJyG0_2;
	wire w_dff_B_TKzAi6Gl3_2;
	wire w_dff_B_6ynsMQ2l0_2;
	wire w_dff_B_bhnIZjwp3_2;
	wire w_dff_B_tXVk6FcT9_2;
	wire w_dff_B_58LdgK666_2;
	wire w_dff_B_gzIk7S020_2;
	wire w_dff_B_szxKorJG7_2;
	wire w_dff_B_f5OiTOd96_2;
	wire w_dff_B_e6WLPQm50_2;
	wire w_dff_B_2F000M8A6_2;
	wire w_dff_B_IFocsjVe8_2;
	wire w_dff_B_1Y0NbcHw4_2;
	wire w_dff_B_8w1rBpYa0_2;
	wire w_dff_B_eGCw48JR6_2;
	wire w_dff_B_Ym96BF5n5_2;
	wire w_dff_B_7GNR9CiQ1_2;
	wire w_dff_B_jydhBZkv3_2;
	wire w_dff_B_XwbwARax8_2;
	wire w_dff_B_XUXLl9PZ6_2;
	wire w_dff_B_9s5BgiKq1_2;
	wire w_dff_B_cbhmIanl0_2;
	wire w_dff_B_53C2nhS84_2;
	wire w_dff_B_UbLtddzG5_2;
	wire w_dff_B_KsXZ429F1_2;
	wire w_dff_B_rrGJcutx6_2;
	wire w_dff_B_mdjShcxc7_2;
	wire w_dff_B_6MPxDqRq9_2;
	wire w_dff_B_Uj77CKxn5_2;
	wire w_dff_B_VDZ8DIOG4_2;
	wire w_dff_B_lS3yPT7e4_2;
	wire w_dff_B_8uBAOWGH5_2;
	wire w_dff_B_26cPxGU03_2;
	wire w_dff_B_LrqcIO5M8_2;
	wire w_dff_B_aE2A8Mk01_2;
	wire w_dff_B_x0b2LiBp2_2;
	wire w_dff_B_oh5mULbq1_2;
	wire w_dff_B_eWtrvpIs8_1;
	wire w_dff_B_SEXWdAiT6_2;
	wire w_dff_B_mNob9bnb3_2;
	wire w_dff_B_Rq2NlqbI9_2;
	wire w_dff_B_Mx0VVGVZ5_2;
	wire w_dff_B_dViLjMkg3_2;
	wire w_dff_B_2ZNy9ijD6_2;
	wire w_dff_B_zYGaFDGy4_2;
	wire w_dff_B_tEeN3z9T5_2;
	wire w_dff_B_AxSFZzne9_2;
	wire w_dff_B_tWQnD0L75_2;
	wire w_dff_B_sDYprePW0_2;
	wire w_dff_B_WQqs7YsP8_2;
	wire w_dff_B_OG5ng1w95_2;
	wire w_dff_B_MiR8bfbQ0_2;
	wire w_dff_B_YZLiTGSk0_2;
	wire w_dff_B_EnkYOP629_2;
	wire w_dff_B_Mr0QJ2Rl2_2;
	wire w_dff_B_7Sbwzsal4_2;
	wire w_dff_B_ZBxEJg4i8_2;
	wire w_dff_B_D6LTuJuE5_2;
	wire w_dff_B_saW3zqss9_2;
	wire w_dff_B_KcjWQJfm3_2;
	wire w_dff_B_i9E5E1I67_2;
	wire w_dff_B_JW1bkQxN0_2;
	wire w_dff_B_e2OkxWGi5_2;
	wire w_dff_B_xJhJw2nF1_2;
	wire w_dff_B_wXwwq99M3_2;
	wire w_dff_B_GbvRjd4Z4_2;
	wire w_dff_B_wEKKARbf3_2;
	wire w_dff_B_Apw4MyEK7_2;
	wire w_dff_B_vVS5O0Tl3_2;
	wire w_dff_B_bhfZ3va88_2;
	wire w_dff_B_P4om3MHF6_2;
	wire w_dff_B_ulKX7iad3_2;
	wire w_dff_B_7qJFgdvK6_2;
	wire w_dff_B_1c96IQu83_2;
	wire w_dff_B_9Dh0EJpF6_2;
	wire w_dff_B_wYij6kNY8_2;
	wire w_dff_B_4GVMkThx5_2;
	wire w_dff_B_KFTi04Gr6_2;
	wire w_dff_B_lTDcgB0E7_2;
	wire w_dff_B_EBXg5wWk4_1;
	wire w_dff_B_CS0Eygq89_2;
	wire w_dff_B_tZDpSqCR3_2;
	wire w_dff_B_KbDKyaV90_2;
	wire w_dff_B_aNfeVkdx7_2;
	wire w_dff_B_HjDldspW8_2;
	wire w_dff_B_vsXKsXhd8_2;
	wire w_dff_B_mworufgv5_2;
	wire w_dff_B_EAgftY1d4_2;
	wire w_dff_B_5mH1526m9_2;
	wire w_dff_B_MGMWnnIC6_2;
	wire w_dff_B_gsLYPoQi5_2;
	wire w_dff_B_EznCGRIn1_2;
	wire w_dff_B_CHsZoZUY8_2;
	wire w_dff_B_JsWHldx16_2;
	wire w_dff_B_LYm6CVXr4_2;
	wire w_dff_B_jWypSJo20_2;
	wire w_dff_B_Sqw4sEgo6_2;
	wire w_dff_B_kVl59ngq4_2;
	wire w_dff_B_k48YUVn62_2;
	wire w_dff_B_JXehVPJs1_2;
	wire w_dff_B_d9IGH2WH9_2;
	wire w_dff_B_EFMcX0Bi4_2;
	wire w_dff_B_pBk6d6VG7_2;
	wire w_dff_B_B7dy0SCz9_2;
	wire w_dff_B_wV1OtUmf9_2;
	wire w_dff_B_0fkp3bTY3_2;
	wire w_dff_B_Jug4uxFi6_2;
	wire w_dff_B_dHAEEWK13_2;
	wire w_dff_B_fQPqUJfB7_2;
	wire w_dff_B_dsG3ScMA0_2;
	wire w_dff_B_xXtdYtIG7_2;
	wire w_dff_B_MJMUtV6s6_2;
	wire w_dff_B_JAChyVXO1_2;
	wire w_dff_B_cC53jNmb5_2;
	wire w_dff_B_Ypjycl5A1_2;
	wire w_dff_B_Qs83rpz59_2;
	wire w_dff_B_g95BrBah1_2;
	wire w_dff_B_kTo0wJwr9_1;
	wire w_dff_B_xXfvTIEd0_2;
	wire w_dff_B_ctNTb8Vz8_2;
	wire w_dff_B_OYTBoBDN5_2;
	wire w_dff_B_sxvJC70M6_2;
	wire w_dff_B_x7kPA3hh2_2;
	wire w_dff_B_A0qOBcfU0_2;
	wire w_dff_B_dNMv3fYf8_2;
	wire w_dff_B_MLygmdTh6_2;
	wire w_dff_B_qHf0FhW84_2;
	wire w_dff_B_hG1YzoXd2_2;
	wire w_dff_B_EyEr9Flw2_2;
	wire w_dff_B_Yq8VIdSQ8_2;
	wire w_dff_B_Gku1QtqH0_2;
	wire w_dff_B_RNxEJiZe6_2;
	wire w_dff_B_m2PhG3Yg5_2;
	wire w_dff_B_LxhWNwgI0_2;
	wire w_dff_B_l56bxpkC6_2;
	wire w_dff_B_YpCP5Imj6_2;
	wire w_dff_B_Bf7M6seD1_2;
	wire w_dff_B_MmXmCIyY0_2;
	wire w_dff_B_Spc6bhKa1_2;
	wire w_dff_B_r5cNsBke1_2;
	wire w_dff_B_nHrTzs1x6_2;
	wire w_dff_B_z8BuF0Ov7_2;
	wire w_dff_B_Qy6Ze7tF0_2;
	wire w_dff_B_g8XNXJmE1_2;
	wire w_dff_B_YcrhXcAJ0_2;
	wire w_dff_B_DyvprqCN1_2;
	wire w_dff_B_iVPqHczQ2_2;
	wire w_dff_B_Ui4cwZhr5_2;
	wire w_dff_B_ugUEf2eZ9_2;
	wire w_dff_B_6ZFVxRWY6_2;
	wire w_dff_B_IFTw00kJ0_1;
	wire w_dff_B_RdtKvNYk3_2;
	wire w_dff_B_PYP44jYz2_2;
	wire w_dff_B_VC9rdrPe5_2;
	wire w_dff_B_683VvSZM6_2;
	wire w_dff_B_HDIY0YNw2_2;
	wire w_dff_B_alUXG5IP2_2;
	wire w_dff_B_SH10VcSh0_2;
	wire w_dff_B_7aTyqGo02_2;
	wire w_dff_B_plSKXuKT6_2;
	wire w_dff_B_EPFTNTCF3_2;
	wire w_dff_B_Aqhfj5nR5_2;
	wire w_dff_B_YfFf0rx90_2;
	wire w_dff_B_59uJ2E770_2;
	wire w_dff_B_NU8mHIPF2_2;
	wire w_dff_B_Nh5cQURV0_2;
	wire w_dff_B_Qwg1tJgI4_2;
	wire w_dff_B_oBTCs1Ic9_2;
	wire w_dff_B_XklLRYk78_2;
	wire w_dff_B_GPxNX4dw3_2;
	wire w_dff_B_jDbtH2FR7_2;
	wire w_dff_B_7ezMDUGa6_2;
	wire w_dff_B_ieCxqmrM1_2;
	wire w_dff_B_58kcIXwr5_2;
	wire w_dff_B_jgVScGte7_2;
	wire w_dff_B_kVei2QwS4_2;
	wire w_dff_B_G6KMSaKk6_2;
	wire w_dff_B_0MYWOVCF2_2;
	wire w_dff_B_RqFGWpq18_2;
	wire w_dff_B_SaWBszGf8_2;
	wire w_dff_B_DMjZiILv3_2;
	wire w_dff_B_P7pV3xtN2_1;
	wire w_dff_B_cAv5JQXD4_2;
	wire w_dff_B_Ci97n3TX3_2;
	wire w_dff_B_QUZc3E899_2;
	wire w_dff_B_OXQttdKS8_2;
	wire w_dff_B_MrVLvbVi6_2;
	wire w_dff_B_2r5jHqnC5_2;
	wire w_dff_B_yNIcBTNp0_2;
	wire w_dff_B_uLGDsaIN0_2;
	wire w_dff_B_y1WSSNpM2_2;
	wire w_dff_B_YtGwdiAQ3_2;
	wire w_dff_B_qe8iiywU7_2;
	wire w_dff_B_6l0Wpm4N9_2;
	wire w_dff_B_VZVm6zFy0_2;
	wire w_dff_B_q2C1g8q56_2;
	wire w_dff_B_boap64Cn4_2;
	wire w_dff_B_oxSfq6k95_2;
	wire w_dff_B_WVnCnoJi5_2;
	wire w_dff_B_Q0dkQHni8_2;
	wire w_dff_B_xlSSTIkI9_2;
	wire w_dff_B_rUa4M8Eg4_2;
	wire w_dff_B_OTarkhj05_2;
	wire w_dff_B_Xh3xVpyD0_2;
	wire w_dff_B_7AhYg2xx1_2;
	wire w_dff_B_IDndbqFh3_2;
	wire w_dff_B_MbvSBqjA3_2;
	wire w_dff_B_59Rap77Z8_2;
	wire w_dff_B_8SaeRHr09_2;
	wire w_dff_B_fvBuavZm2_1;
	wire w_dff_B_rikRDUoQ1_2;
	wire w_dff_B_ODqYfBd60_2;
	wire w_dff_B_stjmCUix9_2;
	wire w_dff_B_W1CnToUL2_2;
	wire w_dff_B_nQibsh9b1_2;
	wire w_dff_B_kKp3HgM66_2;
	wire w_dff_B_umLtDdPn9_2;
	wire w_dff_B_BPR8izXS1_2;
	wire w_dff_B_qkOfTQAf0_2;
	wire w_dff_B_WLXmD37M5_2;
	wire w_dff_B_1jGcuY3J0_2;
	wire w_dff_B_MssQaZhz4_2;
	wire w_dff_B_4Y6TmLK67_2;
	wire w_dff_B_aI1Fc56f5_2;
	wire w_dff_B_3pmW3EdN4_2;
	wire w_dff_B_72SL8DNq3_2;
	wire w_dff_B_LGk9zbWS5_2;
	wire w_dff_B_O5NBdmpQ8_2;
	wire w_dff_B_2AiuQ0aa5_2;
	wire w_dff_B_R4gBO1sg1_2;
	wire w_dff_B_6S7DUVKu4_2;
	wire w_dff_B_s3V2nT0A2_2;
	wire w_dff_B_mIQobraJ3_2;
	wire w_dff_B_FU4KmCfZ3_2;
	wire w_dff_B_8eTcrcM07_1;
	wire w_dff_B_BpDJCnWy6_2;
	wire w_dff_B_c4Ac7gBD1_2;
	wire w_dff_B_q5sa0PWj0_2;
	wire w_dff_B_embPnHVU0_2;
	wire w_dff_B_VdXsQq5V5_2;
	wire w_dff_B_ClWm7J4h1_2;
	wire w_dff_B_96uQTumw9_2;
	wire w_dff_B_ZlA23hll0_2;
	wire w_dff_B_8DPtsfbq1_2;
	wire w_dff_B_1qKzQJJP8_2;
	wire w_dff_B_M0w7T2lc0_2;
	wire w_dff_B_mBifnvAS7_2;
	wire w_dff_B_8JcM7pM71_2;
	wire w_dff_B_EwOgen9I2_2;
	wire w_dff_B_Vcf7JBKS5_2;
	wire w_dff_B_e7VYbVbi1_2;
	wire w_dff_B_9pHvuOoV7_2;
	wire w_dff_B_83EA3s7T5_2;
	wire w_dff_B_V6q3kUu22_2;
	wire w_dff_B_sx23HeQZ2_2;
	wire w_dff_B_aZm2xLBW4_2;
	wire w_dff_B_S4B5uJt66_1;
	wire w_dff_B_WJNUuhNB8_2;
	wire w_dff_B_ErLCSPMA9_2;
	wire w_dff_B_3U4Xjlvm5_2;
	wire w_dff_B_7nm19qju8_2;
	wire w_dff_B_3fJvhWbh9_2;
	wire w_dff_B_oSfWurtQ4_2;
	wire w_dff_B_f4WRCaVE0_2;
	wire w_dff_B_2Mtrg2IV3_2;
	wire w_dff_B_1F4gxY6Q7_2;
	wire w_dff_B_NuWwU2qs6_2;
	wire w_dff_B_MIncjyIH1_2;
	wire w_dff_B_ZgAoVJIJ3_2;
	wire w_dff_B_efVkfXK28_2;
	wire w_dff_B_kFYl820U7_2;
	wire w_dff_B_M8n77AtN2_2;
	wire w_dff_B_qFN8LtCW0_2;
	wire w_dff_B_7weLBBiR8_2;
	wire w_dff_B_3TVnsZem2_2;
	wire w_dff_B_tEIsuwSY6_1;
	wire w_dff_B_7D12UUX70_2;
	wire w_dff_B_eHnnMSzG1_2;
	wire w_dff_B_S24SvMsw7_2;
	wire w_dff_B_345aMDvI1_2;
	wire w_dff_B_oLj4Ws795_2;
	wire w_dff_B_bq8Tivif7_2;
	wire w_dff_B_PKtjp3DY0_2;
	wire w_dff_B_D8Aa3MQq6_2;
	wire w_dff_B_kwYhMsJa9_2;
	wire w_dff_B_ShhZK4Dh8_2;
	wire w_dff_B_BrJCwibb1_2;
	wire w_dff_B_R3ndHCbo9_2;
	wire w_dff_B_YR6wcwMd9_2;
	wire w_dff_B_0qnDpiRu7_2;
	wire w_dff_B_8aMSco662_2;
	wire w_dff_B_dvYDu3121_1;
	wire w_dff_B_sGKYpW7A1_2;
	wire w_dff_B_bfIW92sH1_2;
	wire w_dff_B_Fsgw87Dp9_2;
	wire w_dff_B_9T1ypWOQ6_2;
	wire w_dff_B_OcvriUyv4_2;
	wire w_dff_B_1L2foCBo2_2;
	wire w_dff_B_dbicMcUa1_2;
	wire w_dff_B_2INhwtRo7_2;
	wire w_dff_B_WjTeDR5t1_2;
	wire w_dff_B_lhZez3Wi3_2;
	wire w_dff_B_lEt3Fjqo3_2;
	wire w_dff_B_Vd6fMmaD0_2;
	wire w_dff_B_rX2M1cWh8_1;
	wire w_dff_B_c50el4ku7_2;
	wire w_dff_B_c98Z24RB0_2;
	wire w_dff_B_h0AshvrR1_2;
	wire w_dff_B_Cl50itll5_2;
	wire w_dff_B_lq4ZSHCx9_2;
	wire w_dff_B_I93lvMkg4_2;
	wire w_dff_B_oe9DYwCn9_2;
	wire w_dff_B_GURg5o5w9_2;
	wire w_dff_B_VI1NDn6o2_2;
	wire w_dff_B_ifZxfT5A3_2;
	wire w_dff_B_9WGQxfkY6_2;
	wire w_dff_B_kuP3yNXd4_1;
	wire w_dff_B_6JvFeimc6_1;
	wire w_dff_B_j4e8ueRL0_2;
	wire w_dff_B_bJXOhhWn9_2;
	wire w_dff_B_3QPnI6HQ7_2;
	wire w_dff_B_P53qelmo0_0;
	wire w_dff_A_46UlZCZ00_0;
	wire w_dff_A_Y85roqRL0_0;
	wire w_dff_A_c6VNpxpW0_1;
	wire w_dff_A_as2XVWPH6_1;
	wire w_dff_B_IuxRMeHR7_1;
	wire w_dff_A_XICyd0S42_1;
	wire w_dff_B_cNIx8qef4_1;
	wire w_dff_B_5VH3S5KC4_2;
	wire w_dff_B_eonfFV8u8_2;
	wire w_dff_B_56vQnV2A8_2;
	wire w_dff_B_eO0lWiz65_2;
	wire w_dff_B_oC8nM5Yi5_2;
	wire w_dff_B_vwgx5DcS3_2;
	wire w_dff_B_fFVJZIG67_2;
	wire w_dff_B_d4FGOjfo9_2;
	wire w_dff_B_UILQIAy54_2;
	wire w_dff_B_KoF4gMht1_2;
	wire w_dff_B_Wn5ugI7L7_2;
	wire w_dff_B_rjqHnoJX9_2;
	wire w_dff_B_n6GBJcvL2_2;
	wire w_dff_B_Dt4sJqKx5_2;
	wire w_dff_B_BJI9yP0M9_2;
	wire w_dff_B_vrLlW9cl6_2;
	wire w_dff_B_3LRHKtQS9_2;
	wire w_dff_B_aCKGDVyq4_2;
	wire w_dff_B_ORugJqgg6_2;
	wire w_dff_B_5efZ3p6X7_2;
	wire w_dff_B_UwK4YVAB1_2;
	wire w_dff_B_euxLNvD36_2;
	wire w_dff_B_Dd2Sk7f24_2;
	wire w_dff_B_LVENd3dJ2_2;
	wire w_dff_B_73vxsRqY7_2;
	wire w_dff_B_lwlF5osT4_2;
	wire w_dff_B_E2oGo5wO3_2;
	wire w_dff_B_0ECbxJA31_2;
	wire w_dff_B_X4oyjOEb6_2;
	wire w_dff_B_mhVll2lE1_2;
	wire w_dff_B_f6oVvfJU1_2;
	wire w_dff_B_kyuORWib9_2;
	wire w_dff_B_xPcuBZK88_2;
	wire w_dff_B_5PC7VOl03_2;
	wire w_dff_B_u6CBGsXu3_2;
	wire w_dff_B_Jd60A3Jd8_2;
	wire w_dff_B_4ugWdidr7_2;
	wire w_dff_B_Wv25tivg8_2;
	wire w_dff_B_Fcmq35nS5_2;
	wire w_dff_B_6bRSeZ6Y0_2;
	wire w_dff_B_k9zFCfFa8_2;
	wire w_dff_B_UIxhGLUA5_2;
	wire w_dff_B_eTtUuq7z1_2;
	wire w_dff_B_eG0Dg59U6_2;
	wire w_dff_B_QtGIqCeq3_2;
	wire w_dff_B_Vd1YzWeS3_2;
	wire w_dff_B_Eq8KXynb3_2;
	wire w_dff_B_42Kb9K9Y3_2;
	wire w_dff_B_wOQWxcFM9_2;
	wire w_dff_B_kZfnxLQn1_2;
	wire w_dff_B_XI9aL1kA6_2;
	wire w_dff_B_YZ2J9A3L8_1;
	wire w_dff_B_qmakESc91_2;
	wire w_dff_B_eu2GnKC27_2;
	wire w_dff_B_PwLcmGNU4_2;
	wire w_dff_B_WAsqVksa8_2;
	wire w_dff_B_6WIRJcBQ2_2;
	wire w_dff_B_BhEidsID0_2;
	wire w_dff_B_GbCx0CF75_2;
	wire w_dff_B_PLhHUix31_2;
	wire w_dff_B_Gu0HUX2A1_2;
	wire w_dff_B_Sn5Vhz4B5_2;
	wire w_dff_B_FuwVTXdU6_2;
	wire w_dff_B_1rVF39iu2_2;
	wire w_dff_B_KsixzHA04_2;
	wire w_dff_B_fYltOazL9_2;
	wire w_dff_B_GK1aQCcu0_2;
	wire w_dff_B_eMqGJ8F13_2;
	wire w_dff_B_3zEYds2h1_2;
	wire w_dff_B_gcFnD3vg5_2;
	wire w_dff_B_rgjRzDTl7_2;
	wire w_dff_B_FGUL7rSd9_2;
	wire w_dff_B_AE4XgTMc7_2;
	wire w_dff_B_OpgnOYYm3_2;
	wire w_dff_B_GLwLq8Om5_2;
	wire w_dff_B_8IGFw4n75_2;
	wire w_dff_B_o3nhPfho0_2;
	wire w_dff_B_aBT5OuNh7_2;
	wire w_dff_B_NS0kfxfQ2_2;
	wire w_dff_B_emF6X8te7_2;
	wire w_dff_B_s1XKdGf11_2;
	wire w_dff_B_t5twnAwt4_2;
	wire w_dff_B_RWA8z1rd4_2;
	wire w_dff_B_tGQ1HdrO5_2;
	wire w_dff_B_cnVcqDy19_2;
	wire w_dff_B_YcoEt3Rc4_2;
	wire w_dff_B_Ke7e9Ui86_2;
	wire w_dff_B_8OtDWy1P2_2;
	wire w_dff_B_sG4f9neP9_2;
	wire w_dff_B_JRXAlELz5_2;
	wire w_dff_B_XoZAkpvS4_2;
	wire w_dff_B_LWMAvW8f8_2;
	wire w_dff_B_32XNziaG7_2;
	wire w_dff_B_zULAgVPI8_2;
	wire w_dff_B_Dc2eUq571_2;
	wire w_dff_B_9yEx8lTI4_2;
	wire w_dff_B_7wcgc0jE1_2;
	wire w_dff_B_R2b2iea10_2;
	wire w_dff_B_9JNkZehn3_2;
	wire w_dff_B_qIxe3vd75_1;
	wire w_dff_B_NVfbZG8w5_2;
	wire w_dff_B_q31nTGiS3_2;
	wire w_dff_B_yj1Oysll0_2;
	wire w_dff_B_NNh7bi0w6_2;
	wire w_dff_B_OMaqo4Ru2_2;
	wire w_dff_B_XHID7XCf1_2;
	wire w_dff_B_MOkMZ7Md9_2;
	wire w_dff_B_s9qYIOlf6_2;
	wire w_dff_B_9wN18sTM0_2;
	wire w_dff_B_nAWgq8vi1_2;
	wire w_dff_B_ZGYvdwqG6_2;
	wire w_dff_B_BwM7BUln4_2;
	wire w_dff_B_3DYt0mkP2_2;
	wire w_dff_B_TjitmiLP6_2;
	wire w_dff_B_B6KatWc69_2;
	wire w_dff_B_jJyY4cTE7_2;
	wire w_dff_B_ZDJN93Bu5_2;
	wire w_dff_B_4ybuubSP4_2;
	wire w_dff_B_qYAC7WbY1_2;
	wire w_dff_B_HYOiJHHU0_2;
	wire w_dff_B_slKoBVAO3_2;
	wire w_dff_B_v73g2qe33_2;
	wire w_dff_B_RRwZcDg88_2;
	wire w_dff_B_v7PMVfU24_2;
	wire w_dff_B_Ig3GQaC66_2;
	wire w_dff_B_UH5SJ1ty1_2;
	wire w_dff_B_gbY1j1Mp7_2;
	wire w_dff_B_Nan30Hjt2_2;
	wire w_dff_B_9PByZS5W8_2;
	wire w_dff_B_qwSj470X6_2;
	wire w_dff_B_9MKSPDSP3_2;
	wire w_dff_B_u8vTxEML2_2;
	wire w_dff_B_YXpqEmOj2_2;
	wire w_dff_B_9j7eYWqM0_2;
	wire w_dff_B_I7XImHNI4_2;
	wire w_dff_B_z9Rgkd8u4_2;
	wire w_dff_B_0pDl5VBX2_2;
	wire w_dff_B_ZkHN4mcn7_2;
	wire w_dff_B_JfmcWgGP3_2;
	wire w_dff_B_R82lrEbb0_2;
	wire w_dff_B_VDz2SiDw3_2;
	wire w_dff_B_QBDy5FYn6_2;
	wire w_dff_B_uQ6Ji3YS2_2;
	wire w_dff_B_2UH6Sju27_1;
	wire w_dff_B_KPqezL1z7_2;
	wire w_dff_B_LKVCHkt39_2;
	wire w_dff_B_Kub1RPoA5_2;
	wire w_dff_B_KxCVWRow4_2;
	wire w_dff_B_CCr9oJcR6_2;
	wire w_dff_B_BgfVez5E5_2;
	wire w_dff_B_JvFE5xG48_2;
	wire w_dff_B_wAeifTfD6_2;
	wire w_dff_B_r7SEr9GN3_2;
	wire w_dff_B_iWc8oDqp6_2;
	wire w_dff_B_PjOst9vO6_2;
	wire w_dff_B_KFSz1UYg8_2;
	wire w_dff_B_stk4p4U24_2;
	wire w_dff_B_LzvV4MbZ0_2;
	wire w_dff_B_SZIE7ewA0_2;
	wire w_dff_B_PSpzbNGq7_2;
	wire w_dff_B_6wEnHQ3O8_2;
	wire w_dff_B_9rBjxFsq1_2;
	wire w_dff_B_3QJIp8YZ9_2;
	wire w_dff_B_Yjt6tcos6_2;
	wire w_dff_B_nc5pdmiF8_2;
	wire w_dff_B_QDHaZHBr1_2;
	wire w_dff_B_g9QSn8kA9_2;
	wire w_dff_B_zzJ2wYow2_2;
	wire w_dff_B_xJW8AOW98_2;
	wire w_dff_B_YLOkRTk84_2;
	wire w_dff_B_c8afeDPF4_2;
	wire w_dff_B_6qhEYN629_2;
	wire w_dff_B_8L7B1R8z3_2;
	wire w_dff_B_MvYxJbrD3_2;
	wire w_dff_B_0hN6HVNw3_2;
	wire w_dff_B_MjmfVJrZ1_2;
	wire w_dff_B_ybvTQLDj6_2;
	wire w_dff_B_NBui3msE9_2;
	wire w_dff_B_b7o55a3V5_2;
	wire w_dff_B_bYHH4Yfc8_2;
	wire w_dff_B_N9AL9DrK6_2;
	wire w_dff_B_g4sqGszj0_2;
	wire w_dff_B_YuhbQnDV1_2;
	wire w_dff_B_QaZA6LOD3_1;
	wire w_dff_B_RzWB5iSg2_2;
	wire w_dff_B_NdfeGn7z7_2;
	wire w_dff_B_I4ubmTIl0_2;
	wire w_dff_B_iWz0g9oD4_2;
	wire w_dff_B_CjGinJYp1_2;
	wire w_dff_B_BLnkTZ9F0_2;
	wire w_dff_B_V1dW6LMn0_2;
	wire w_dff_B_UlYrC57j3_2;
	wire w_dff_B_oKIsmv7I1_2;
	wire w_dff_B_s0T3wLst3_2;
	wire w_dff_B_DsevGJRv5_2;
	wire w_dff_B_3HG2h4uj7_2;
	wire w_dff_B_bl2F6YaM6_2;
	wire w_dff_B_jW8y2dBd1_2;
	wire w_dff_B_XHAP7rNe0_2;
	wire w_dff_B_j5ZlGhP52_2;
	wire w_dff_B_7Nc3XTFA8_2;
	wire w_dff_B_5TvAHopH4_2;
	wire w_dff_B_uJ0AlV0R0_2;
	wire w_dff_B_c1mHGTGw3_2;
	wire w_dff_B_P2x1g1VB8_2;
	wire w_dff_B_T6aPQNht1_2;
	wire w_dff_B_70n6rwZV7_2;
	wire w_dff_B_YNZMNGWQ8_2;
	wire w_dff_B_dDnYqVIC0_2;
	wire w_dff_B_LCP5en5G1_2;
	wire w_dff_B_UDmQUMAb0_2;
	wire w_dff_B_1Rf4n2bq3_2;
	wire w_dff_B_KQuy6tPL7_2;
	wire w_dff_B_2SX8haRQ9_2;
	wire w_dff_B_kZx66CwO6_2;
	wire w_dff_B_5ix9SUyF4_2;
	wire w_dff_B_g8O4kjua5_2;
	wire w_dff_B_8XvW1uyN8_2;
	wire w_dff_B_mKfxyogV8_2;
	wire w_dff_B_iQ0mUJQH6_1;
	wire w_dff_B_dQdqVN723_2;
	wire w_dff_B_NTPd2rSh2_2;
	wire w_dff_B_zqV67sBM5_2;
	wire w_dff_B_n099u9Pv0_2;
	wire w_dff_B_6Sab7Gvb9_2;
	wire w_dff_B_gLeGkFh78_2;
	wire w_dff_B_ddkL6cTG5_2;
	wire w_dff_B_XCUWzEbc6_2;
	wire w_dff_B_UrPrCatm2_2;
	wire w_dff_B_eu3o8Ibq0_2;
	wire w_dff_B_hzY9z3lZ4_2;
	wire w_dff_B_n2NpeEVV3_2;
	wire w_dff_B_mNy4Cxjq4_2;
	wire w_dff_B_xZQFpAmx4_2;
	wire w_dff_B_HsqbjUEV3_2;
	wire w_dff_B_wCzqPmun3_2;
	wire w_dff_B_u0zIWOXM2_2;
	wire w_dff_B_UEzWtuxx1_2;
	wire w_dff_B_O71PxFAS5_2;
	wire w_dff_B_wIaZn0DU1_2;
	wire w_dff_B_s7c5mmix7_2;
	wire w_dff_B_G4522sUc5_2;
	wire w_dff_B_9Q1p4yba0_2;
	wire w_dff_B_jhCC9DdC0_2;
	wire w_dff_B_c6yzg8PN3_2;
	wire w_dff_B_LCNauuFj0_2;
	wire w_dff_B_xLJgt0sl3_2;
	wire w_dff_B_jx55aJCp5_2;
	wire w_dff_B_84X8Q3Iq5_2;
	wire w_dff_B_qrmTfwrb9_2;
	wire w_dff_B_KkbJhSEQ3_2;
	wire w_dff_B_ho8lWHFt5_1;
	wire w_dff_B_S58oYmMa0_2;
	wire w_dff_B_IKGTS3zP1_2;
	wire w_dff_B_DUCn5t4Q7_2;
	wire w_dff_B_1MiFA5151_2;
	wire w_dff_B_C6Zyxbbl3_2;
	wire w_dff_B_ZGPI2EY02_2;
	wire w_dff_B_DkH4Sp0K4_2;
	wire w_dff_B_BciaIpX67_2;
	wire w_dff_B_hPADyZlN8_2;
	wire w_dff_B_uN7n0fjF1_2;
	wire w_dff_B_LEEUnOa70_2;
	wire w_dff_B_KhVTjsAB2_2;
	wire w_dff_B_GcII21Rg3_2;
	wire w_dff_B_U71n6pbz7_2;
	wire w_dff_B_XulHHwSR3_2;
	wire w_dff_B_KpREJOeS1_2;
	wire w_dff_B_jTA3M3jC7_2;
	wire w_dff_B_vyF548bN1_2;
	wire w_dff_B_OMv3a6iv1_2;
	wire w_dff_B_Z8u58FAa3_2;
	wire w_dff_B_5p5T4rIz2_2;
	wire w_dff_B_vtpdGxVm4_2;
	wire w_dff_B_KMI7p34y5_2;
	wire w_dff_B_QH1yS4HV2_2;
	wire w_dff_B_AHxknJIR7_2;
	wire w_dff_B_1BL8Ahqj1_2;
	wire w_dff_B_XCPKuwD08_1;
	wire w_dff_B_8fWD4FDZ5_2;
	wire w_dff_B_0bmhFsBP2_2;
	wire w_dff_B_L8tmRKeS6_2;
	wire w_dff_B_Zq0PgvtI0_2;
	wire w_dff_B_bh9e0hKE9_2;
	wire w_dff_B_gvCo8ja90_2;
	wire w_dff_B_vPabyj2N4_2;
	wire w_dff_B_C4KObj3N2_2;
	wire w_dff_B_6tM6Bikm2_2;
	wire w_dff_B_Fxh8FrRE8_2;
	wire w_dff_B_1eMWfmE62_2;
	wire w_dff_B_iLlOrbvU8_2;
	wire w_dff_B_LoGDqp0X6_2;
	wire w_dff_B_24k2RjLd8_2;
	wire w_dff_B_2fR7Wl904_2;
	wire w_dff_B_k1RGTAP00_2;
	wire w_dff_B_ccpovmWP2_2;
	wire w_dff_B_fyHA7Bdf4_2;
	wire w_dff_B_fu7MWsCY7_2;
	wire w_dff_B_i43YjZIH4_2;
	wire w_dff_B_Wv5N0oYO3_2;
	wire w_dff_B_cb5H1mkX6_2;
	wire w_dff_B_QDSLTbY30_2;
	wire w_dff_B_HCQgwVJi0_2;
	wire w_dff_B_JqAWgDf77_1;
	wire w_dff_B_cjg5O9F09_2;
	wire w_dff_B_eD6PzqY11_2;
	wire w_dff_B_0mU4iFnm1_2;
	wire w_dff_B_sXGLcywk4_2;
	wire w_dff_B_83KL4U2s0_2;
	wire w_dff_B_qnPe1rC34_2;
	wire w_dff_B_FjH128Yc7_2;
	wire w_dff_B_3MVQSV9i7_2;
	wire w_dff_B_7RFmhv6M5_2;
	wire w_dff_B_9bqj45Az9_2;
	wire w_dff_B_jcI5yAf75_2;
	wire w_dff_B_e3mmbSYq6_2;
	wire w_dff_B_jtjhHmXu3_2;
	wire w_dff_B_BQSGshNK2_2;
	wire w_dff_B_hiE1BAur6_2;
	wire w_dff_B_PBJpxvx89_2;
	wire w_dff_B_2sugV3bU7_2;
	wire w_dff_B_xIxdlzct2_2;
	wire w_dff_B_swwuuHOT8_2;
	wire w_dff_B_f1fCDRhk4_2;
	wire w_dff_B_Xe6He2ej0_2;
	wire w_dff_B_bVIrtuqp5_1;
	wire w_dff_B_6m1xM35V8_2;
	wire w_dff_B_Cg7d4s2f6_2;
	wire w_dff_B_WXTTm8Gk6_2;
	wire w_dff_B_QmjzsAcW2_2;
	wire w_dff_B_LtJR30tu6_2;
	wire w_dff_B_Nsc63dWk3_2;
	wire w_dff_B_DompU1Mn5_2;
	wire w_dff_B_qNgr9wnv7_2;
	wire w_dff_B_7qLpwFRF7_2;
	wire w_dff_B_FMwohWg13_2;
	wire w_dff_B_sm3ZAiPd7_2;
	wire w_dff_B_PGvRhzpx8_2;
	wire w_dff_B_Ff6loTOH1_2;
	wire w_dff_B_JGntCBvc0_2;
	wire w_dff_B_tgJVvPhR1_2;
	wire w_dff_B_fYzdwXKl8_2;
	wire w_dff_B_n2dKzKE83_2;
	wire w_dff_B_I90VvDvk6_2;
	wire w_dff_B_RyEVqxOx9_1;
	wire w_dff_B_5y5m7if40_2;
	wire w_dff_B_C7NOqQmo0_2;
	wire w_dff_B_nOiyILY67_2;
	wire w_dff_B_Nr3nNIHK5_2;
	wire w_dff_B_Sldwm07Z4_2;
	wire w_dff_B_696ONaBT7_2;
	wire w_dff_B_5WJOaiIf6_2;
	wire w_dff_B_owGEMTNz7_2;
	wire w_dff_B_MTvfbLHM2_2;
	wire w_dff_B_QejiHL5P1_2;
	wire w_dff_B_blyeLdE39_2;
	wire w_dff_B_ftThUZDC8_2;
	wire w_dff_B_1OYb2m226_2;
	wire w_dff_B_Ci9wtgQJ5_2;
	wire w_dff_B_smVEtmv42_2;
	wire w_dff_B_zrwX1Wfj8_1;
	wire w_dff_B_Vyrvde2k7_2;
	wire w_dff_B_7dHNVaiX3_2;
	wire w_dff_B_Z07SO9pK4_2;
	wire w_dff_B_CU3VdFFs7_2;
	wire w_dff_B_1pRFknuG1_2;
	wire w_dff_B_pDyPHFbo8_2;
	wire w_dff_B_hW581FkD7_2;
	wire w_dff_B_ax2HaJUt4_2;
	wire w_dff_B_XyB4ET0e1_2;
	wire w_dff_B_7FkRkUes7_2;
	wire w_dff_B_imKGIIwC7_2;
	wire w_dff_B_NGWTcjpH5_2;
	wire w_dff_B_4oC1homs9_1;
	wire w_dff_B_aWKR5lhH0_2;
	wire w_dff_B_AciXEQ3X1_2;
	wire w_dff_B_RC2f9G3l3_2;
	wire w_dff_B_EuFkQLMU9_2;
	wire w_dff_B_d7qrxhmy8_2;
	wire w_dff_B_lKZInh7R6_2;
	wire w_dff_B_lvn5e4YR2_2;
	wire w_dff_B_wSpih1Qt8_2;
	wire w_dff_B_9x4o2KCf7_2;
	wire w_dff_B_OzCmzcbf7_2;
	wire w_dff_B_aL4m3DRC6_2;
	wire w_dff_B_9hdXcse39_1;
	wire w_dff_B_IPyqcC861_1;
	wire w_dff_B_U4bDjFzh5_2;
	wire w_dff_B_LYiWz5wH8_2;
	wire w_dff_B_BUBibZu93_2;
	wire w_dff_B_A0THsbh72_0;
	wire w_dff_A_sRUxz9k22_0;
	wire w_dff_A_sb8ifWuf6_0;
	wire w_dff_A_v5IQem1f2_1;
	wire w_dff_A_YptSCDAG8_1;
	wire w_dff_B_3khtPMZW2_1;
	wire w_dff_B_9DLV4WV10_1;
	wire w_dff_B_faZ3ZuPl5_1;
	wire w_dff_B_MfPpxzJJ9_2;
	wire w_dff_B_wqld1sS99_2;
	wire w_dff_B_TFMUueFe3_2;
	wire w_dff_B_meT1L5XU9_2;
	wire w_dff_B_eIGPAlFf5_2;
	wire w_dff_B_GYFatfmk0_2;
	wire w_dff_B_UFZSArsj2_2;
	wire w_dff_B_brlA7cSV0_2;
	wire w_dff_B_m91rymN61_2;
	wire w_dff_B_bZPLzYsL4_2;
	wire w_dff_B_g3fF2vhK7_2;
	wire w_dff_B_NSDCk7Dd7_2;
	wire w_dff_B_GX258PLG1_2;
	wire w_dff_B_GlgEY3dY5_2;
	wire w_dff_B_w9khd0Be5_2;
	wire w_dff_B_2lfrzC9f1_2;
	wire w_dff_B_9PLjGxQl9_2;
	wire w_dff_B_LiCwUIuV8_2;
	wire w_dff_B_hYnWIWjr6_2;
	wire w_dff_B_Xmzl4cMp4_2;
	wire w_dff_B_NoZ2XuEd6_2;
	wire w_dff_B_uHW3695z4_2;
	wire w_dff_B_YYFN2Zed4_2;
	wire w_dff_B_yYEalvjV5_2;
	wire w_dff_B_NvM6fDmN8_2;
	wire w_dff_B_BuhkKyiz1_2;
	wire w_dff_B_USWE1dzW0_2;
	wire w_dff_B_HpAjlrzA1_2;
	wire w_dff_B_vYBqpBVu4_2;
	wire w_dff_B_UJbJAONb9_2;
	wire w_dff_B_PHo3CXyP2_2;
	wire w_dff_B_mcM7JGJ51_2;
	wire w_dff_B_fdrUX4wB3_2;
	wire w_dff_B_s1gwsI996_2;
	wire w_dff_B_FQBwSGez0_2;
	wire w_dff_B_sHeUz6nC6_2;
	wire w_dff_B_cOsl4YVb1_2;
	wire w_dff_B_fTwFTflT5_2;
	wire w_dff_B_H5yL1yby8_2;
	wire w_dff_B_a8SEDwBz6_2;
	wire w_dff_B_TwxTjr6m7_2;
	wire w_dff_B_Yxnipmd05_2;
	wire w_dff_B_0gvTZBI68_2;
	wire w_dff_B_PB7KWXqT8_2;
	wire w_dff_B_Lko5MVvg3_2;
	wire w_dff_B_HSCpKC7y0_2;
	wire w_dff_B_OrMGwLI38_2;
	wire w_dff_B_uTO94k8z0_2;
	wire w_dff_B_Jj1COXCJ9_2;
	wire w_dff_B_Ar2B9dB93_2;
	wire w_dff_B_fkpKJ1nu2_2;
	wire w_dff_B_77zVpOrb5_2;
	wire w_dff_B_6aixUHpW2_2;
	wire w_dff_B_IGeMV9ib9_2;
	wire w_dff_B_1hXPoMWS8_2;
	wire w_dff_B_hTm9IOLP4_2;
	wire w_dff_B_lUSdTHp65_2;
	wire w_dff_B_nkhFoypa0_2;
	wire w_dff_B_hFKUTLDw7_2;
	wire w_dff_B_OlSnPDNG8_2;
	wire w_dff_B_MJVdG18b0_2;
	wire w_dff_B_uHrKPwcu2_2;
	wire w_dff_B_ARfFCk4c8_2;
	wire w_dff_B_0uOtnRUs4_2;
	wire w_dff_B_GgziSO107_2;
	wire w_dff_B_f2H1AQPX8_2;
	wire w_dff_B_Wbda1GtI8_2;
	wire w_dff_B_YzgAQTqb6_2;
	wire w_dff_B_5a1WIX7l3_2;
	wire w_dff_B_DGGBXSaQ6_2;
	wire w_dff_B_zKSRgERY3_2;
	wire w_dff_B_ZH41LcwF6_2;
	wire w_dff_B_JxGqPK4N2_2;
	wire w_dff_B_vdOInZ5o7_2;
	wire w_dff_B_wq5U4Wf54_2;
	wire w_dff_B_8DNgGRHO6_2;
	wire w_dff_B_hBdRicXW5_2;
	wire w_dff_B_y05gS8lc0_2;
	wire w_dff_B_CKs8n0Ga0_2;
	wire w_dff_B_QSqeWaxf5_2;
	wire w_dff_B_vkXyBreC2_2;
	wire w_dff_B_RH3bIGlB7_2;
	wire w_dff_B_nkG0x9KF5_2;
	wire w_dff_B_99JDZfRv1_2;
	wire w_dff_B_gC5WPp5f2_2;
	wire w_dff_B_9gwnppzM2_2;
	wire w_dff_B_UGPfeOys5_2;
	wire w_dff_B_1p3qAfnr3_2;
	wire w_dff_B_nzqDpM5g9_2;
	wire w_dff_B_j2gRuAmv6_2;
	wire w_dff_B_qjyyVmx96_2;
	wire w_dff_B_MOd2wavx1_2;
	wire w_dff_B_edEKACBM9_2;
	wire w_dff_B_iMCb9WWC1_2;
	wire w_dff_B_2EolgRcV6_2;
	wire w_dff_B_eQikfSyF9_2;
	wire w_dff_B_zZP6iBpU1_2;
	wire w_dff_B_sxPkbQoA5_2;
	wire w_dff_B_UVizJ9OA6_2;
	wire w_dff_B_Qmo4U34Y5_2;
	wire w_dff_B_PxKGak9c1_2;
	wire w_dff_B_bZvZbHM05_2;
	wire w_dff_B_BTIdkmGU8_2;
	wire w_dff_B_LjShF65B1_2;
	wire w_dff_B_Sx5j2Lhm8_2;
	wire w_dff_B_wGYfX4iD3_2;
	wire w_dff_B_77mgntCa2_2;
	wire w_dff_B_JTBAVYp00_2;
	wire w_dff_A_kIMEJZuV4_1;
	wire w_dff_B_kLCCYxg90_1;
	wire w_dff_B_6WvChU4n7_2;
	wire w_dff_B_VeE8k1Js9_2;
	wire w_dff_B_b0ffJJZ37_2;
	wire w_dff_B_qUAGjAFZ7_2;
	wire w_dff_B_HbUZ7giP6_2;
	wire w_dff_B_225T9Tfg2_2;
	wire w_dff_B_2Ebq5G2f8_2;
	wire w_dff_B_qLonYJt09_2;
	wire w_dff_B_rW4he9le3_2;
	wire w_dff_B_WltqSuis1_2;
	wire w_dff_B_WH1ZPVG68_2;
	wire w_dff_B_JxdmMQdi8_2;
	wire w_dff_B_YtQ5t4BL2_2;
	wire w_dff_B_9cMtjPah8_2;
	wire w_dff_B_T714fXWc2_2;
	wire w_dff_B_5ehTGXKN0_2;
	wire w_dff_B_U3HENvgj9_2;
	wire w_dff_B_sale1tLe9_2;
	wire w_dff_B_uG6YmGoK2_2;
	wire w_dff_B_ucI4AD7R8_2;
	wire w_dff_B_2AtVjVru3_2;
	wire w_dff_B_wi2x7uf67_2;
	wire w_dff_B_oWb3rbPn0_2;
	wire w_dff_B_GAs5Apbm0_2;
	wire w_dff_B_89P7xuT70_2;
	wire w_dff_B_UzxMRUuo1_2;
	wire w_dff_B_UtvfWYMs8_2;
	wire w_dff_B_vTVOUeVN0_2;
	wire w_dff_B_tnw1i2EO3_2;
	wire w_dff_B_utnlB5gF5_2;
	wire w_dff_B_0jtgF9Pa2_2;
	wire w_dff_B_ToWwYuCP9_2;
	wire w_dff_B_3ElCogYp8_2;
	wire w_dff_B_da2by9p20_2;
	wire w_dff_B_XiqeBoTE8_2;
	wire w_dff_B_7PW0mHnc6_2;
	wire w_dff_B_LvrPfIdk7_2;
	wire w_dff_B_DFZ8lVSh3_2;
	wire w_dff_B_pXOmb06k6_2;
	wire w_dff_B_FrGaBkqP7_2;
	wire w_dff_B_DRKSCwm95_2;
	wire w_dff_B_CfL2HHFE9_2;
	wire w_dff_B_R1wbpUy81_2;
	wire w_dff_B_u2A0zG2l8_2;
	wire w_dff_B_bGYF4gsT3_2;
	wire w_dff_B_5DYZp9407_2;
	wire w_dff_B_n49NGnNO7_2;
	wire w_dff_B_0p1ewIGR8_2;
	wire w_dff_B_pee5vlDs6_2;
	wire w_dff_B_Nu1GZGt17_2;
	wire w_dff_B_04UzHpm74_2;
	wire w_dff_B_vc5rPiNp8_2;
	wire w_dff_B_IIrK9S8e4_1;
	wire w_dff_B_KInWw2Ze8_1;
	wire w_dff_B_NvrZTT2W4_2;
	wire w_dff_B_De0raXHb8_2;
	wire w_dff_B_8ufEoUho1_2;
	wire w_dff_B_WfiKk9ED1_2;
	wire w_dff_B_RR8CyNt29_2;
	wire w_dff_B_fwbLCIO69_2;
	wire w_dff_B_bIZv65pX6_2;
	wire w_dff_B_WlTNzLHA3_2;
	wire w_dff_B_bZc4q3YB1_2;
	wire w_dff_B_IhhxcOd89_2;
	wire w_dff_B_bvdpctnm3_2;
	wire w_dff_B_GHdlnLmj6_2;
	wire w_dff_B_mtzGz4AY3_2;
	wire w_dff_B_QGx8HGMa5_2;
	wire w_dff_B_L91D3la25_2;
	wire w_dff_B_CZ8Y5NwY2_2;
	wire w_dff_B_tpEbFM308_2;
	wire w_dff_B_9NpQc4t86_2;
	wire w_dff_B_YCFMKMzF9_2;
	wire w_dff_B_B3EHuTda0_2;
	wire w_dff_B_JhLcc2yb1_2;
	wire w_dff_B_mquBrRvZ8_2;
	wire w_dff_B_QaQo3S3Q2_2;
	wire w_dff_B_3VG0ynRn9_2;
	wire w_dff_B_t2D9BH491_2;
	wire w_dff_B_wZwMO1n63_2;
	wire w_dff_B_CSEUDD1e1_2;
	wire w_dff_B_saawBkeW2_2;
	wire w_dff_B_UemBGa1j1_2;
	wire w_dff_B_98nErRHJ8_2;
	wire w_dff_B_11LC3EgX4_2;
	wire w_dff_B_MjhrhxhZ0_2;
	wire w_dff_B_EZjFtKMT9_2;
	wire w_dff_B_jdkNWGqi4_2;
	wire w_dff_B_BQuO9eMB8_2;
	wire w_dff_B_qwHNU55a6_2;
	wire w_dff_B_iciNOIY51_2;
	wire w_dff_B_S48muyIX0_2;
	wire w_dff_B_K7cPHnl28_2;
	wire w_dff_B_f6nEfctv1_2;
	wire w_dff_B_IDk7U9bE4_2;
	wire w_dff_B_e6LfYu1o8_2;
	wire w_dff_B_NxnBI4752_2;
	wire w_dff_B_ExZacyRm6_2;
	wire w_dff_B_x5WR6gah7_2;
	wire w_dff_B_PaHaOLhD0_2;
	wire w_dff_B_0IALB7UA1_2;
	wire w_dff_B_NBVbAG3x8_2;
	wire w_dff_B_PIWEmWL32_2;
	wire w_dff_B_iImEmESC3_2;
	wire w_dff_B_ioW0lsdf2_2;
	wire w_dff_B_b8avPETQ4_2;
	wire w_dff_B_Gl93NYTU5_2;
	wire w_dff_B_Bv4Iw56G1_2;
	wire w_dff_B_NFDbYbnJ8_2;
	wire w_dff_B_ZHjLGGQq6_2;
	wire w_dff_B_vHlc8EKC4_2;
	wire w_dff_B_aN7Pusvh5_2;
	wire w_dff_B_ZJeEpx7f1_2;
	wire w_dff_B_hNeWZUh13_2;
	wire w_dff_B_Wv0oDHv37_2;
	wire w_dff_B_DY2AlFEn3_2;
	wire w_dff_B_AxjmYavE4_2;
	wire w_dff_B_OFJpi7aV4_2;
	wire w_dff_B_viHaDg3n8_2;
	wire w_dff_B_6KAxKkF52_2;
	wire w_dff_B_WvUy9Xgj7_2;
	wire w_dff_B_yjPwEgj65_2;
	wire w_dff_B_ceBBZEjj7_2;
	wire w_dff_B_xn6GsXHo8_2;
	wire w_dff_B_cGsJNLJ77_2;
	wire w_dff_B_dibxXs7f9_2;
	wire w_dff_B_BVXcjW8O3_2;
	wire w_dff_B_WHKlnkAW0_2;
	wire w_dff_B_JS1aW1tV3_2;
	wire w_dff_B_TOrT2Hal9_2;
	wire w_dff_B_edlU4s8A5_2;
	wire w_dff_B_N2b6l1Lb9_2;
	wire w_dff_B_1Q8PyZCg0_2;
	wire w_dff_B_Ryb6VMY08_2;
	wire w_dff_B_mL8KOsxt8_2;
	wire w_dff_B_Lqpb9cmN6_2;
	wire w_dff_B_we1dICRd6_2;
	wire w_dff_B_hlQ9slZK8_2;
	wire w_dff_B_OTAyjO1U2_2;
	wire w_dff_B_0t2RPjdF7_2;
	wire w_dff_B_VNckG46C8_2;
	wire w_dff_B_5AnD0mq88_2;
	wire w_dff_B_64R7jRtM0_2;
	wire w_dff_B_yZFX5zYs1_2;
	wire w_dff_B_rat0vrnm5_2;
	wire w_dff_B_cjrXDAJm2_2;
	wire w_dff_B_SX2lUEYc6_2;
	wire w_dff_B_fP9B9w7o9_2;
	wire w_dff_B_YdQuE3et0_2;
	wire w_dff_B_mDd0gWwf2_2;
	wire w_dff_B_hEINZUw46_2;
	wire w_dff_B_4S6Z5FUH4_2;
	wire w_dff_B_GAvzG52H4_2;
	wire w_dff_B_Lam9kCm25_2;
	wire w_dff_B_962kAxAN4_2;
	wire w_dff_B_w3zmnl6r0_1;
	wire w_dff_B_doL0YCC16_2;
	wire w_dff_B_PO80Hljs3_2;
	wire w_dff_B_tAoJnxxI7_2;
	wire w_dff_B_I9tNYdXt6_2;
	wire w_dff_B_xVYa1lsO8_2;
	wire w_dff_B_eGZKkaC31_2;
	wire w_dff_B_ag97yKCq3_2;
	wire w_dff_B_r5LZPEN60_2;
	wire w_dff_B_8GMA7ssn8_2;
	wire w_dff_B_HZSYmuGw2_2;
	wire w_dff_B_zpNYHYiv5_2;
	wire w_dff_B_GK7qFWiW3_2;
	wire w_dff_B_Tv4ccQm50_2;
	wire w_dff_B_lx9X790e1_2;
	wire w_dff_B_69GtdHYW0_2;
	wire w_dff_B_H8BvjoBO4_2;
	wire w_dff_B_U0rRh0O24_2;
	wire w_dff_B_Yft8nIWx2_2;
	wire w_dff_B_TULcQlcD6_2;
	wire w_dff_B_I6nnn3an5_2;
	wire w_dff_B_4UavkAXR7_2;
	wire w_dff_B_meDrfdmn5_2;
	wire w_dff_B_mZmAkMTK6_2;
	wire w_dff_B_DWy7vFSZ3_2;
	wire w_dff_B_u9cOpx384_2;
	wire w_dff_B_PrUIrbZJ0_2;
	wire w_dff_B_d0RyFGEL1_2;
	wire w_dff_B_w4FEVQiI4_2;
	wire w_dff_B_2V7g2ufw7_2;
	wire w_dff_B_qmcX0Slb6_2;
	wire w_dff_B_bi3efb5G8_2;
	wire w_dff_B_GGyeunjO4_2;
	wire w_dff_B_YYY4kqJg7_2;
	wire w_dff_B_c2rmAP3l6_2;
	wire w_dff_B_usUNnHza6_2;
	wire w_dff_B_P4zJadhL9_2;
	wire w_dff_B_cc8eC8nn5_2;
	wire w_dff_B_A6n8MjoI5_2;
	wire w_dff_B_meZHDjPW6_2;
	wire w_dff_B_hYYQqhYG9_2;
	wire w_dff_B_h5C3FUQk0_2;
	wire w_dff_B_hgpcHUij2_2;
	wire w_dff_B_waOVNIE37_2;
	wire w_dff_B_xnqK7Byh6_2;
	wire w_dff_B_p7B7sbbP7_2;
	wire w_dff_B_DcLUZTiI2_2;
	wire w_dff_B_G20dCVcg1_2;
	wire w_dff_B_Gqhqk55Q6_2;
	wire w_dff_B_KSBx9hgd8_1;
	wire w_dff_B_HuYfgTST5_1;
	wire w_dff_B_NRarIm481_2;
	wire w_dff_B_bNkLPfhj3_2;
	wire w_dff_B_HsTrgkDH7_2;
	wire w_dff_B_WJ1K3ROM2_2;
	wire w_dff_B_Sy2gkp6g9_2;
	wire w_dff_B_vQw3N8xP1_2;
	wire w_dff_B_hu3d0up95_2;
	wire w_dff_B_bwTsxGle8_2;
	wire w_dff_B_ZVHMzRyU3_2;
	wire w_dff_B_Aa3Ruav88_2;
	wire w_dff_B_1hOm2KMg3_2;
	wire w_dff_B_PstwEAOL5_2;
	wire w_dff_B_SBC3Jut87_2;
	wire w_dff_B_1x4BOWQm9_2;
	wire w_dff_B_FPk5bM1R3_2;
	wire w_dff_B_AZNJ5v4x4_2;
	wire w_dff_B_TCdxf6yk6_2;
	wire w_dff_B_13eA2AlI8_2;
	wire w_dff_B_BneWj0V76_2;
	wire w_dff_B_4GUV5hjH8_2;
	wire w_dff_B_GytnC5GA3_2;
	wire w_dff_B_vgouNKQR2_2;
	wire w_dff_B_ARMT9Ao40_2;
	wire w_dff_B_KyBIYozU9_2;
	wire w_dff_B_EnifDq9L0_2;
	wire w_dff_B_6uVhiURb5_2;
	wire w_dff_B_doFOBq3C3_2;
	wire w_dff_B_PiALsGyr0_2;
	wire w_dff_B_edLLhkFo3_2;
	wire w_dff_B_SCokj42K4_2;
	wire w_dff_B_1UDNjSQa5_2;
	wire w_dff_B_RcZVIRtI1_2;
	wire w_dff_B_l14ZrkSU1_2;
	wire w_dff_B_nsUfkMOK9_2;
	wire w_dff_B_iYkn4oJr6_2;
	wire w_dff_B_qY0Midl32_2;
	wire w_dff_B_YrCBHve83_2;
	wire w_dff_B_RzP8ufSE6_2;
	wire w_dff_B_3OaYdXdL7_2;
	wire w_dff_B_sIdjzXAe4_2;
	wire w_dff_B_iNTIn2dh8_2;
	wire w_dff_B_eJivWHm39_2;
	wire w_dff_B_OsKF9fUF4_2;
	wire w_dff_B_7atpzyXC7_2;
	wire w_dff_B_f45WlC394_2;
	wire w_dff_B_hbLmOOlo1_2;
	wire w_dff_B_YjCazqQQ3_2;
	wire w_dff_B_t1xsbvDJ0_2;
	wire w_dff_B_ZgDqR1Pc8_2;
	wire w_dff_B_jC8a5Z0i6_2;
	wire w_dff_B_CtOC030R1_2;
	wire w_dff_B_KvAkGQWQ1_2;
	wire w_dff_B_GxhBTZam8_2;
	wire w_dff_B_hmvdfGcC1_2;
	wire w_dff_B_WofEt4Ay7_2;
	wire w_dff_B_Dq5naBde3_2;
	wire w_dff_B_tM7YFD2G3_2;
	wire w_dff_B_ES7BqhXo1_2;
	wire w_dff_B_04aS6UYb8_2;
	wire w_dff_B_bdSMKOBd5_2;
	wire w_dff_B_mF38fRtk7_2;
	wire w_dff_B_CutgmOio5_2;
	wire w_dff_B_SjFGFVOn6_2;
	wire w_dff_B_L0kR6tUv3_2;
	wire w_dff_B_KI5fYqMu0_2;
	wire w_dff_B_iX5CW8J70_2;
	wire w_dff_B_YDENOHEJ1_2;
	wire w_dff_B_0aMEzOUL1_2;
	wire w_dff_B_xbVwIZ758_2;
	wire w_dff_B_uCaqHB5Y1_2;
	wire w_dff_B_lnPNylQo6_2;
	wire w_dff_B_0edCn8cW7_2;
	wire w_dff_B_tlPVmLpa7_2;
	wire w_dff_B_CrNf6jlH1_2;
	wire w_dff_B_5uTOTLMr7_2;
	wire w_dff_B_ayMTJqjq5_2;
	wire w_dff_B_ZJSE5A6u8_2;
	wire w_dff_B_JOaVQVlj1_2;
	wire w_dff_B_87GpAEat4_2;
	wire w_dff_B_R4e1XHKk7_2;
	wire w_dff_B_acDlqHo75_2;
	wire w_dff_B_tzmShRyT4_2;
	wire w_dff_B_5gTMTT226_2;
	wire w_dff_B_qf7enKqJ3_2;
	wire w_dff_B_SjS9F0V23_2;
	wire w_dff_B_81SDYdzI1_2;
	wire w_dff_B_r6NlxRvS2_2;
	wire w_dff_B_honvnWC47_2;
	wire w_dff_B_Pm4lz2TE6_2;
	wire w_dff_B_qNm5DonE1_2;
	wire w_dff_B_SV2kvBoR0_2;
	wire w_dff_B_EBIpuuQR8_2;
	wire w_dff_B_WeM40RcL6_2;
	wire w_dff_B_ntpkS7Lg8_1;
	wire w_dff_B_lG7B0dfC4_2;
	wire w_dff_B_KJecEGLT1_2;
	wire w_dff_B_5mxEd2ES5_2;
	wire w_dff_B_p5mWZGv34_2;
	wire w_dff_B_ojpNVx150_2;
	wire w_dff_B_si9fCXoa2_2;
	wire w_dff_B_OCgk9N5P9_2;
	wire w_dff_B_WnmibGQH6_2;
	wire w_dff_B_ph9dCYgJ7_2;
	wire w_dff_B_5VGsv4e43_2;
	wire w_dff_B_XZbLP5Lf1_2;
	wire w_dff_B_MNC0GTuQ2_2;
	wire w_dff_B_JbaTNY7h6_2;
	wire w_dff_B_HQyyC0Ks2_2;
	wire w_dff_B_vY6PerlF7_2;
	wire w_dff_B_1hAp9e208_2;
	wire w_dff_B_XlhxLxdf4_2;
	wire w_dff_B_ya1aadhD8_2;
	wire w_dff_B_6b2jPVpP9_2;
	wire w_dff_B_ls1Z6PYf3_2;
	wire w_dff_B_Q32PWZgJ5_2;
	wire w_dff_B_nOu8jI8L3_2;
	wire w_dff_B_ThscDitp7_2;
	wire w_dff_B_RJkYcvaE6_2;
	wire w_dff_B_XxLkv4WB8_2;
	wire w_dff_B_4a0Znj3O4_2;
	wire w_dff_B_j9tULFLz3_2;
	wire w_dff_B_n8hs05Cd5_2;
	wire w_dff_B_LPoWhfUl3_2;
	wire w_dff_B_j1zwFrvm4_2;
	wire w_dff_B_xtrKM9KJ5_2;
	wire w_dff_B_gStlqySk1_2;
	wire w_dff_B_m1XEFau04_2;
	wire w_dff_B_rgFpqpQt5_2;
	wire w_dff_B_pJTzBIea4_2;
	wire w_dff_B_VmGD0QdK1_2;
	wire w_dff_B_tL8n37lo1_2;
	wire w_dff_B_1EEhgPRe6_2;
	wire w_dff_B_W2gLu4uP4_2;
	wire w_dff_B_zrvBGAS09_2;
	wire w_dff_B_k9bITiLT4_2;
	wire w_dff_B_BamoOFI32_2;
	wire w_dff_B_kY5qNx0X4_2;
	wire w_dff_B_hc8D6Meq7_2;
	wire w_dff_B_WENRyFSp3_1;
	wire w_dff_B_dofnAvnv2_1;
	wire w_dff_B_pSBUtnzf2_2;
	wire w_dff_B_O3wxnIq12_2;
	wire w_dff_B_14OyNwMz8_2;
	wire w_dff_B_R2UkBLZN6_2;
	wire w_dff_B_Ir5t8v328_2;
	wire w_dff_B_vvhWlZZ94_2;
	wire w_dff_B_p3wJfSXo4_2;
	wire w_dff_B_FI3lRxcy8_2;
	wire w_dff_B_hUfJYE093_2;
	wire w_dff_B_GnXh7Pqn2_2;
	wire w_dff_B_98zCHcyQ2_2;
	wire w_dff_B_e1qiWSwR7_2;
	wire w_dff_B_SOnsn3GE9_2;
	wire w_dff_B_S6xX9IMr5_2;
	wire w_dff_B_U2PTNmWC1_2;
	wire w_dff_B_HhKI1uqI6_2;
	wire w_dff_B_AuJP7aRH3_2;
	wire w_dff_B_E4oFzWpb5_2;
	wire w_dff_B_hR4v2NY77_2;
	wire w_dff_B_vFwUmgL80_2;
	wire w_dff_B_CUYVvrqS3_2;
	wire w_dff_B_C5fZiopT0_2;
	wire w_dff_B_QuAmi1I34_2;
	wire w_dff_B_vr3iXH2W2_2;
	wire w_dff_B_HotQv0NS4_2;
	wire w_dff_B_HCGhOKUu4_2;
	wire w_dff_B_1MuYgIjq2_2;
	wire w_dff_B_MB9s2mwy8_2;
	wire w_dff_B_g3DZWlK20_2;
	wire w_dff_B_Q1XIJ01N1_2;
	wire w_dff_B_pl1VKKq94_2;
	wire w_dff_B_6M08i3Rs0_2;
	wire w_dff_B_ueYOJYnk6_2;
	wire w_dff_B_RMmkhvFz7_2;
	wire w_dff_B_m1BpQfr49_2;
	wire w_dff_B_ScpP36Ta3_2;
	wire w_dff_B_y7uob3vh7_2;
	wire w_dff_B_cSZHN7Iz6_2;
	wire w_dff_B_T0aF33hJ2_2;
	wire w_dff_B_8V6d5mBP2_2;
	wire w_dff_B_qvorlkVc9_2;
	wire w_dff_B_ORVskRRL0_2;
	wire w_dff_B_uFLbA16n0_2;
	wire w_dff_B_hPPU42YS7_2;
	wire w_dff_B_zSHorKoy5_2;
	wire w_dff_B_Dsq5ntar3_2;
	wire w_dff_B_hkowsfGn2_2;
	wire w_dff_B_zzUlKvej9_2;
	wire w_dff_B_nlG2aPkr8_2;
	wire w_dff_B_hpD5bY4P9_2;
	wire w_dff_B_lwvS4Zqz8_2;
	wire w_dff_B_h47sk5SR6_2;
	wire w_dff_B_z07UA75T7_2;
	wire w_dff_B_hoiRqGj51_2;
	wire w_dff_B_BU8PtD0b4_2;
	wire w_dff_B_ruquY5fG5_2;
	wire w_dff_B_ZoTcBwNy0_2;
	wire w_dff_B_zHr4kXGj1_2;
	wire w_dff_B_ACzXzg0L4_2;
	wire w_dff_B_rP9G3l960_2;
	wire w_dff_B_Rp6DzqGG0_2;
	wire w_dff_B_GBP0cfjm9_2;
	wire w_dff_B_MVtfaO6K0_2;
	wire w_dff_B_QXqo12Wh5_2;
	wire w_dff_B_X11AiJN49_2;
	wire w_dff_B_rSkWizs21_2;
	wire w_dff_B_GbEMdghI6_2;
	wire w_dff_B_CghXusbL2_2;
	wire w_dff_B_AHRYWI4h6_2;
	wire w_dff_B_b10RUB805_2;
	wire w_dff_B_E0DuHRWX5_2;
	wire w_dff_B_DQki4TfN8_2;
	wire w_dff_B_BJxRN4Rq8_2;
	wire w_dff_B_gUA60vJn9_2;
	wire w_dff_B_NKbBbhAo5_2;
	wire w_dff_B_OY1yIeMD6_2;
	wire w_dff_B_1AsiLKXu0_2;
	wire w_dff_B_YOk2K5Xj7_2;
	wire w_dff_B_5QgVmLnI6_2;
	wire w_dff_B_6Qk5svwe4_2;
	wire w_dff_B_V6ItlT3I2_2;
	wire w_dff_B_82aBdxM65_2;
	wire w_dff_B_GZT2zF813_2;
	wire w_dff_B_Iwu0JBoY1_2;
	wire w_dff_B_fSAmthdF5_2;
	wire w_dff_B_so3bvXCA9_1;
	wire w_dff_B_vtEi4Kpz3_2;
	wire w_dff_B_rMh5kDWf4_2;
	wire w_dff_B_W3huiePw8_2;
	wire w_dff_B_GmeMhhA71_2;
	wire w_dff_B_C7QERlP91_2;
	wire w_dff_B_84s5c5Nz2_2;
	wire w_dff_B_7ZW0x3g02_2;
	wire w_dff_B_aPDhGeFP9_2;
	wire w_dff_B_KaUutlwy9_2;
	wire w_dff_B_bySvzJn36_2;
	wire w_dff_B_O66wpek53_2;
	wire w_dff_B_aizqsT1X0_2;
	wire w_dff_B_aiutfzTc1_2;
	wire w_dff_B_12oASWHn1_2;
	wire w_dff_B_alXqnom34_2;
	wire w_dff_B_ONerYRmf7_2;
	wire w_dff_B_Rrpl6yNC2_2;
	wire w_dff_B_ix0Gi1mB1_2;
	wire w_dff_B_zNqUTJr67_2;
	wire w_dff_B_EmUI2uyv6_2;
	wire w_dff_B_x5jrItde3_2;
	wire w_dff_B_PvovAB4y7_2;
	wire w_dff_B_Bh9Ch4t81_2;
	wire w_dff_B_i92uPmxT6_2;
	wire w_dff_B_raTTTJJC9_2;
	wire w_dff_B_niThLe7M3_2;
	wire w_dff_B_JuaK0qrj5_2;
	wire w_dff_B_NBcwkllt8_2;
	wire w_dff_B_aYlYT9TL0_2;
	wire w_dff_B_0rHLpv2Q3_2;
	wire w_dff_B_aspizn5w9_2;
	wire w_dff_B_Lh31jnUz8_2;
	wire w_dff_B_tQKoUhBA2_2;
	wire w_dff_B_BaVR6MCD1_2;
	wire w_dff_B_Eq2yXbdA5_2;
	wire w_dff_B_EW9AYF2q3_2;
	wire w_dff_B_rjDBiP412_2;
	wire w_dff_B_VlbZDsvX9_2;
	wire w_dff_B_EZofrVWs8_2;
	wire w_dff_B_YSlYmL2F6_2;
	wire w_dff_B_Jfqm8b2C2_1;
	wire w_dff_B_XGro1DDU8_1;
	wire w_dff_B_DCt7W3KY5_2;
	wire w_dff_B_Ze1Gbbtc4_2;
	wire w_dff_B_afN3qDdr6_2;
	wire w_dff_B_zNipOtPz0_2;
	wire w_dff_B_T48beAEl9_2;
	wire w_dff_B_zanLY2pj5_2;
	wire w_dff_B_o3WkWxfY1_2;
	wire w_dff_B_4ODzqni49_2;
	wire w_dff_B_Nd0ab4CN2_2;
	wire w_dff_B_ZQLpiDU95_2;
	wire w_dff_B_mGISbn4m9_2;
	wire w_dff_B_lSaa4y9E0_2;
	wire w_dff_B_bMaQ7bwB8_2;
	wire w_dff_B_V7dQB2OC2_2;
	wire w_dff_B_cyHswZPc6_2;
	wire w_dff_B_24iqTy5j5_2;
	wire w_dff_B_8xclsG7e0_2;
	wire w_dff_B_wOx0yO1d7_2;
	wire w_dff_B_HnLvbag86_2;
	wire w_dff_B_1dpNgc582_2;
	wire w_dff_B_inlD8xDw3_2;
	wire w_dff_B_rpjd2GH41_2;
	wire w_dff_B_DjxsCOey1_2;
	wire w_dff_B_EF4Ictk27_2;
	wire w_dff_B_Mbcn8u8I1_2;
	wire w_dff_B_KZy9Wzyl2_2;
	wire w_dff_B_oTyIkkL54_2;
	wire w_dff_B_2Eqq8dfa6_2;
	wire w_dff_B_RplELcYv5_2;
	wire w_dff_B_Mpd7KjoO9_2;
	wire w_dff_B_6ZIO1vSb3_2;
	wire w_dff_B_r1Iwv30N4_2;
	wire w_dff_B_7LBpGpU68_2;
	wire w_dff_B_jrTO1hzs4_2;
	wire w_dff_B_0dPZOt1m0_2;
	wire w_dff_B_Xqy7mTJH3_2;
	wire w_dff_B_nLDF5s0E1_2;
	wire w_dff_B_Gn5z5N8B7_2;
	wire w_dff_B_oxrMN8Kh5_2;
	wire w_dff_B_4Na5e2Ve2_2;
	wire w_dff_B_mqT7sGcI9_2;
	wire w_dff_B_I0wq4VfE7_2;
	wire w_dff_B_4p7ifI9w6_2;
	wire w_dff_B_8KitNCqB3_2;
	wire w_dff_B_E8h5qvUD1_2;
	wire w_dff_B_wDljcrXF6_2;
	wire w_dff_B_FGQZMneQ8_2;
	wire w_dff_B_S4IAZWVB1_2;
	wire w_dff_B_2Kh34KYl0_2;
	wire w_dff_B_ZPGuMP478_2;
	wire w_dff_B_xxvAtJO13_2;
	wire w_dff_B_w8vxuQ7V0_2;
	wire w_dff_B_IG7nORry1_2;
	wire w_dff_B_PSJ3wbRG5_2;
	wire w_dff_B_IwR4VEJz9_2;
	wire w_dff_B_0AN5FYnj7_2;
	wire w_dff_B_rUYiWd898_2;
	wire w_dff_B_YAml3ti30_2;
	wire w_dff_B_KXMdH0Dv1_2;
	wire w_dff_B_GoOFHact8_2;
	wire w_dff_B_y1NWIWDG0_2;
	wire w_dff_B_2PNBIXAu4_2;
	wire w_dff_B_rqmfBGFq8_2;
	wire w_dff_B_LlQ4oQ0Q5_2;
	wire w_dff_B_zXddmIFX4_2;
	wire w_dff_B_VMphltbY0_2;
	wire w_dff_B_mcgQLaqK0_2;
	wire w_dff_B_islzgUuV1_2;
	wire w_dff_B_HzXEvtSl7_2;
	wire w_dff_B_90Nz1PCK0_2;
	wire w_dff_B_QcZsuWx58_2;
	wire w_dff_B_qpxyykvy9_2;
	wire w_dff_B_tjsDtm5i5_2;
	wire w_dff_B_PwJXIweD9_2;
	wire w_dff_B_f2N7aWOk5_2;
	wire w_dff_B_SKoI0v3m4_2;
	wire w_dff_B_GhTEZuUV2_2;
	wire w_dff_B_egK88UFU6_1;
	wire w_dff_B_nuPRXyN19_2;
	wire w_dff_B_OV3k2TzR9_2;
	wire w_dff_B_AkPfrcEy4_2;
	wire w_dff_B_B9JU5BK58_2;
	wire w_dff_B_95thr4gk8_2;
	wire w_dff_B_3Qn4gqZ09_2;
	wire w_dff_B_5GvkDcz38_2;
	wire w_dff_B_EPcGO0WF1_2;
	wire w_dff_B_bnL5c9sb2_2;
	wire w_dff_B_T8XW9peQ7_2;
	wire w_dff_B_9Yad3EFy0_2;
	wire w_dff_B_zn8z2mBb6_2;
	wire w_dff_B_h4DXpltR5_2;
	wire w_dff_B_lKBVVANg4_2;
	wire w_dff_B_ENot0orb1_2;
	wire w_dff_B_D09HICv27_2;
	wire w_dff_B_OAfFfalN6_2;
	wire w_dff_B_nMq9dOsC3_2;
	wire w_dff_B_K0ZaFbJq8_2;
	wire w_dff_B_uvcL2WJG4_2;
	wire w_dff_B_CZZznmh27_2;
	wire w_dff_B_OhNPlfJw6_2;
	wire w_dff_B_kW2INgSM3_2;
	wire w_dff_B_9bj1JdwC4_2;
	wire w_dff_B_KpoYko7H8_2;
	wire w_dff_B_x6RjqWcj0_2;
	wire w_dff_B_HKZYHUZX9_2;
	wire w_dff_B_nGncQTUi1_2;
	wire w_dff_B_rwrnzylx8_2;
	wire w_dff_B_5rPQpd1L3_2;
	wire w_dff_B_bExroYum5_2;
	wire w_dff_B_yxQpWcGX6_2;
	wire w_dff_B_higTDy5o0_2;
	wire w_dff_B_lL1HJHi17_2;
	wire w_dff_B_uqQT0TR96_2;
	wire w_dff_B_MoL9CwpP0_2;
	wire w_dff_B_N4JfSr7n1_1;
	wire w_dff_B_5qq234Sr4_1;
	wire w_dff_B_K68rkaQn9_2;
	wire w_dff_B_CiM7q6Xq9_2;
	wire w_dff_B_dkzLxwFq0_2;
	wire w_dff_B_uDDFTSOm6_2;
	wire w_dff_B_mgJMzQa61_2;
	wire w_dff_B_VrpVDPnN9_2;
	wire w_dff_B_G4RSUY8j0_2;
	wire w_dff_B_4cME2GAL0_2;
	wire w_dff_B_ez5PiuDK8_2;
	wire w_dff_B_LLI0imW92_2;
	wire w_dff_B_QmHDANHS5_2;
	wire w_dff_B_kI9ytiqq9_2;
	wire w_dff_B_rjTU1pez0_2;
	wire w_dff_B_lpMXW1jg1_2;
	wire w_dff_B_hoUfVHa60_2;
	wire w_dff_B_j0iP1Hub7_2;
	wire w_dff_B_aLBmGYDK6_2;
	wire w_dff_B_fzDOd8fJ1_2;
	wire w_dff_B_TpOVAHZl7_2;
	wire w_dff_B_NKzhgmlF2_2;
	wire w_dff_B_bncAS4Pf5_2;
	wire w_dff_B_LlbdaGVx6_2;
	wire w_dff_B_u1oLIKQV6_2;
	wire w_dff_B_uq7RaOV39_2;
	wire w_dff_B_auCKxZI85_2;
	wire w_dff_B_X5V6IUaz7_2;
	wire w_dff_B_eiviAIJK3_2;
	wire w_dff_B_BGC8ItBU0_2;
	wire w_dff_B_K35cnsZx0_2;
	wire w_dff_B_WaZa6cDR7_2;
	wire w_dff_B_hvBdxNAh1_2;
	wire w_dff_B_1Bs6bCOl1_2;
	wire w_dff_B_3fu1YQq02_2;
	wire w_dff_B_R9BpI6KK7_2;
	wire w_dff_B_rgqCiTNK7_2;
	wire w_dff_B_pW0QKm1x8_2;
	wire w_dff_B_xg1axJwk5_2;
	wire w_dff_B_z8qdQBbT6_2;
	wire w_dff_B_xn1SH1mG0_2;
	wire w_dff_B_0A83RMKG1_2;
	wire w_dff_B_rb4pol9V8_2;
	wire w_dff_B_Ih7bEQca3_2;
	wire w_dff_B_CXOJ9m5j8_2;
	wire w_dff_B_AKdxi1Rf0_2;
	wire w_dff_B_dHN7jQjp8_2;
	wire w_dff_B_mcPNcui82_2;
	wire w_dff_B_rzKFESw93_2;
	wire w_dff_B_UhrocrFL1_2;
	wire w_dff_B_RU89xR409_2;
	wire w_dff_B_fHbRt2Nq6_2;
	wire w_dff_B_QJgFrR4p9_2;
	wire w_dff_B_Sxvk3fOd2_2;
	wire w_dff_B_pMUf683H6_2;
	wire w_dff_B_2pLBPppL5_2;
	wire w_dff_B_jsv79wMI0_2;
	wire w_dff_B_8vTgenk18_2;
	wire w_dff_B_V1SX7UNt0_2;
	wire w_dff_B_31X9wV946_2;
	wire w_dff_B_3NQYAGCw8_2;
	wire w_dff_B_zSEpyaj96_2;
	wire w_dff_B_HKUMPwgn9_2;
	wire w_dff_B_o7bljNKx1_2;
	wire w_dff_B_vBkPOOmw4_2;
	wire w_dff_B_QtazNloG8_2;
	wire w_dff_B_rRJOtmUo5_2;
	wire w_dff_B_tid6EDcB4_2;
	wire w_dff_B_ThuaIvl45_2;
	wire w_dff_B_UxFdy8pr2_2;
	wire w_dff_B_S9b9GWiV5_2;
	wire w_dff_B_HJZteJoN3_1;
	wire w_dff_B_OmvMAqTT0_2;
	wire w_dff_B_pvsZFsx15_2;
	wire w_dff_B_AXr4O4ty0_2;
	wire w_dff_B_862N7lLh1_2;
	wire w_dff_B_P7AhAO7I5_2;
	wire w_dff_B_x1kZzuYt4_2;
	wire w_dff_B_XKApxCph2_2;
	wire w_dff_B_JaHfiVvu5_2;
	wire w_dff_B_yvXraZ4b0_2;
	wire w_dff_B_osxJEzY77_2;
	wire w_dff_B_gtYJYOf66_2;
	wire w_dff_B_XqkQqxjt0_2;
	wire w_dff_B_Oh9Z1gqE0_2;
	wire w_dff_B_sJ956VoH2_2;
	wire w_dff_B_NFSfL3w03_2;
	wire w_dff_B_bhMsQ0N37_2;
	wire w_dff_B_dWoWhe207_2;
	wire w_dff_B_7FrM7QSE4_2;
	wire w_dff_B_jp38REXl8_2;
	wire w_dff_B_JVrL0fzG6_2;
	wire w_dff_B_rgx8hFa92_2;
	wire w_dff_B_mqpK7Xad6_2;
	wire w_dff_B_zeToHgRv0_2;
	wire w_dff_B_EbJNOq1D7_2;
	wire w_dff_B_ZIMh5qSI7_2;
	wire w_dff_B_Ln9EsESf0_2;
	wire w_dff_B_trsadETY7_2;
	wire w_dff_B_xqcF2OXE4_2;
	wire w_dff_B_LCJfPLE72_2;
	wire w_dff_B_snsH9h506_2;
	wire w_dff_B_If3bHUL46_2;
	wire w_dff_B_vCWHOO814_2;
	wire w_dff_B_lyZCPGs11_1;
	wire w_dff_B_R8uxWo708_1;
	wire w_dff_B_46WPqBBn2_2;
	wire w_dff_B_1XWtqaD66_2;
	wire w_dff_B_knW16qmU7_2;
	wire w_dff_B_4GCSMxTt4_2;
	wire w_dff_B_bcXDzk9i8_2;
	wire w_dff_B_ssevscCk1_2;
	wire w_dff_B_t9CUpARs6_2;
	wire w_dff_B_PKkvjSv16_2;
	wire w_dff_B_1tQLeOoh5_2;
	wire w_dff_B_iQ0u0b7B8_2;
	wire w_dff_B_2HVBPVYn0_2;
	wire w_dff_B_Tmz9uCix5_2;
	wire w_dff_B_1a7KvG528_2;
	wire w_dff_B_Y5s6eiW44_2;
	wire w_dff_B_kqvOaVKo7_2;
	wire w_dff_B_r9B0GuIM5_2;
	wire w_dff_B_ostB113k4_2;
	wire w_dff_B_ivdue0726_2;
	wire w_dff_B_SbTmByqZ9_2;
	wire w_dff_B_UpzIo9X63_2;
	wire w_dff_B_9M1mJqd92_2;
	wire w_dff_B_1jWpo7Xj0_2;
	wire w_dff_B_AGK4g5ti1_2;
	wire w_dff_B_vcJ09U567_2;
	wire w_dff_B_uhJs6o5p9_2;
	wire w_dff_B_ZgdaOcBh9_2;
	wire w_dff_B_N5MWngKd2_2;
	wire w_dff_B_BtMKTer00_2;
	wire w_dff_B_00H811zv5_2;
	wire w_dff_B_XI8wn8Uu3_2;
	wire w_dff_B_7BwIwi7Z2_2;
	wire w_dff_B_K3tdjOh04_2;
	wire w_dff_B_nluhx48n8_2;
	wire w_dff_B_NZIDjwhe7_2;
	wire w_dff_B_Zffxkm2s6_2;
	wire w_dff_B_1phQhY8Q9_2;
	wire w_dff_B_xKjVvZqP4_2;
	wire w_dff_B_l0ZUqaLf9_2;
	wire w_dff_B_MWaep3iz6_2;
	wire w_dff_B_hU9AkzUJ6_2;
	wire w_dff_B_AjQpZnQL2_2;
	wire w_dff_B_JC37OW3r9_2;
	wire w_dff_B_hXM82lQv5_2;
	wire w_dff_B_TVfRBuFz0_2;
	wire w_dff_B_4bp5GJi99_2;
	wire w_dff_B_a1Q1jioX6_2;
	wire w_dff_B_lUUGNdUr8_2;
	wire w_dff_B_fLdWDGxq5_2;
	wire w_dff_B_2m5bpYii5_2;
	wire w_dff_B_NTT9AYFE1_2;
	wire w_dff_B_g3vSHVBW2_2;
	wire w_dff_B_f1BJmZyr2_2;
	wire w_dff_B_ZJaPvM3o5_2;
	wire w_dff_B_KDPqWNWF0_2;
	wire w_dff_B_kTuf7nG95_2;
	wire w_dff_B_lCJyOdvc2_2;
	wire w_dff_B_IH3DPNQ59_2;
	wire w_dff_B_dymqQGsn2_2;
	wire w_dff_B_6ELLYYeu3_2;
	wire w_dff_B_VtqpH4MQ5_2;
	wire w_dff_B_ipKRWSpy6_2;
	wire w_dff_B_plcpmFsX2_1;
	wire w_dff_B_Av03ybjv7_2;
	wire w_dff_B_TOXOZ8v72_2;
	wire w_dff_B_8NNliQ6X1_2;
	wire w_dff_B_zKqFceEj0_2;
	wire w_dff_B_u8HlRG636_2;
	wire w_dff_B_1CTfZ9rO2_2;
	wire w_dff_B_NFOgvyNk0_2;
	wire w_dff_B_l4BH1Z9j0_2;
	wire w_dff_B_ps38PL8f9_2;
	wire w_dff_B_3yStKIJO4_2;
	wire w_dff_B_vekcYn1c4_2;
	wire w_dff_B_rUxGzJKf2_2;
	wire w_dff_B_0GKuh1zB5_2;
	wire w_dff_B_8JPsKB0k2_2;
	wire w_dff_B_dx6bcf6z5_2;
	wire w_dff_B_O1DiOXmJ6_2;
	wire w_dff_B_vkte66X21_2;
	wire w_dff_B_aDINbv7V1_2;
	wire w_dff_B_WzghUl385_2;
	wire w_dff_B_z03Ap8BX4_2;
	wire w_dff_B_WwKReFR89_2;
	wire w_dff_B_0huAPqU41_2;
	wire w_dff_B_ucANHPEB7_2;
	wire w_dff_B_ULZfgP8H2_2;
	wire w_dff_B_hsgHv1xE6_2;
	wire w_dff_B_aIIDjXAm4_2;
	wire w_dff_B_9CVhahh19_2;
	wire w_dff_B_B2JJaT8Y1_2;
	wire w_dff_B_YFMKMXf99_1;
	wire w_dff_B_zBIB7LIv3_1;
	wire w_dff_B_2lupi1eT7_2;
	wire w_dff_B_lDeJkaEL8_2;
	wire w_dff_B_m2ps2aC25_2;
	wire w_dff_B_QmTK3o6b0_2;
	wire w_dff_B_Z0VOmMi61_2;
	wire w_dff_B_XLWiyqa95_2;
	wire w_dff_B_EA0yKMqT5_2;
	wire w_dff_B_uYntsCLe6_2;
	wire w_dff_B_W7xGSPqc6_2;
	wire w_dff_B_8BqnZydY8_2;
	wire w_dff_B_KTe0YBW91_2;
	wire w_dff_B_TDNCuHUh6_2;
	wire w_dff_B_F7zplMgm0_2;
	wire w_dff_B_7ziRD5KS4_2;
	wire w_dff_B_Zhr77VUE0_2;
	wire w_dff_B_HvIRCMU08_2;
	wire w_dff_B_Pak5dTBC9_2;
	wire w_dff_B_s7w1pX6x4_2;
	wire w_dff_B_rlNnwseh7_2;
	wire w_dff_B_0GkVLFEq5_2;
	wire w_dff_B_I4XY41NH0_2;
	wire w_dff_B_8NyDsdmn2_2;
	wire w_dff_B_8Ql4FxcU6_2;
	wire w_dff_B_l6HYqmoc5_2;
	wire w_dff_B_7pxHhch97_2;
	wire w_dff_B_A2NDWBwO0_2;
	wire w_dff_B_YNYkrfAJ7_2;
	wire w_dff_B_bN5RRWSv1_2;
	wire w_dff_B_QlHe1He51_2;
	wire w_dff_B_g9NgCkTW4_2;
	wire w_dff_B_A4GuylTi0_2;
	wire w_dff_B_U0GPJpZ77_2;
	wire w_dff_B_fZoFfEII8_2;
	wire w_dff_B_HUKTMELg4_2;
	wire w_dff_B_jqEcdhi14_2;
	wire w_dff_B_z3aWz5gU4_2;
	wire w_dff_B_GoEvd0vC6_2;
	wire w_dff_B_AYPZjyLs3_2;
	wire w_dff_B_YE4EL8mj1_2;
	wire w_dff_B_WzOT6QaG6_2;
	wire w_dff_B_efoCT5ku6_2;
	wire w_dff_B_jD55L0qG7_2;
	wire w_dff_B_QFmHvdPf5_2;
	wire w_dff_B_VOFMawPP0_2;
	wire w_dff_B_iiUpzoe22_2;
	wire w_dff_B_Y30VZ7cH5_2;
	wire w_dff_B_wgDX7S5p8_2;
	wire w_dff_B_uOzOINEo1_2;
	wire w_dff_B_pmP1MQka3_2;
	wire w_dff_B_lCFVNw2c2_2;
	wire w_dff_B_Jm9w6RiA2_2;
	wire w_dff_B_2BeACS201_2;
	wire w_dff_B_8HqNMCiP7_2;
	wire w_dff_B_S026EZg56_1;
	wire w_dff_B_II4gFpzY7_2;
	wire w_dff_B_p6KibwD58_2;
	wire w_dff_B_0NSAln6R0_2;
	wire w_dff_B_6GJH66ZJ3_2;
	wire w_dff_B_arL3XSj35_2;
	wire w_dff_B_uXKY5agJ5_2;
	wire w_dff_B_C1ODHJfy8_2;
	wire w_dff_B_YPbSpx0w3_2;
	wire w_dff_B_GS2BtMHa6_2;
	wire w_dff_B_3S7Xee543_2;
	wire w_dff_B_YIlu3IVC2_2;
	wire w_dff_B_mJEY2d3L8_2;
	wire w_dff_B_BBMuspAo1_2;
	wire w_dff_B_FUoJSM8P2_2;
	wire w_dff_B_FarZG3x59_2;
	wire w_dff_B_D1blQciI4_2;
	wire w_dff_B_PSLsGNfR4_2;
	wire w_dff_B_GkV0GfZV3_2;
	wire w_dff_B_e2573Xix1_2;
	wire w_dff_B_S29BS6Mz3_2;
	wire w_dff_B_SLJeWLzc9_2;
	wire w_dff_B_6IidSZij5_2;
	wire w_dff_B_Yun8i6zT6_2;
	wire w_dff_B_uNJ5Rqbx3_2;
	wire w_dff_B_dfts3IKL9_1;
	wire w_dff_B_L7a03A1l4_1;
	wire w_dff_B_t5tatHDx5_2;
	wire w_dff_B_R4NCvGAC8_2;
	wire w_dff_B_iXGGVD222_2;
	wire w_dff_B_VcZm2RMr9_2;
	wire w_dff_B_7DCWxgRP0_2;
	wire w_dff_B_FfpEEnUS0_2;
	wire w_dff_B_bFwnEhbF0_2;
	wire w_dff_B_xAT24ykD2_2;
	wire w_dff_B_l9Ht3rWf6_2;
	wire w_dff_B_OhHNcRaJ6_2;
	wire w_dff_B_w8ltom5m9_2;
	wire w_dff_B_KRVmArpG9_2;
	wire w_dff_B_icWNlMFz9_2;
	wire w_dff_B_y7zRgHsx7_2;
	wire w_dff_B_292f23vW9_2;
	wire w_dff_B_lMtldrk21_2;
	wire w_dff_B_V0PjiF4E6_2;
	wire w_dff_B_JCtWA6Zp9_2;
	wire w_dff_B_6Kx7oBwQ2_2;
	wire w_dff_B_AjSzTbXd6_2;
	wire w_dff_B_KO8C55j57_2;
	wire w_dff_B_iHBpOj256_2;
	wire w_dff_B_aHWJISxO2_2;
	wire w_dff_B_figRRYyU9_2;
	wire w_dff_B_3ALz3QFj1_2;
	wire w_dff_B_ylZUh7nx1_2;
	wire w_dff_B_uJHYtz8k2_2;
	wire w_dff_B_RA6k6S0C9_2;
	wire w_dff_B_lllBzQUj4_2;
	wire w_dff_B_o1bQoWKX9_2;
	wire w_dff_B_qxNWYZJC9_2;
	wire w_dff_B_R9FC6olV1_2;
	wire w_dff_B_NUWo2WtU2_2;
	wire w_dff_B_IXZKlPZk1_2;
	wire w_dff_B_28AxlOWV2_2;
	wire w_dff_B_gvtEs4qI3_2;
	wire w_dff_B_n0tCGg293_2;
	wire w_dff_B_dfRpefxj8_2;
	wire w_dff_B_HKAXMSIQ3_2;
	wire w_dff_B_4lF1Wtn35_2;
	wire w_dff_B_Ywg0Cgk01_2;
	wire w_dff_B_qDAYAYTz6_2;
	wire w_dff_B_V6JVcxgo2_2;
	wire w_dff_B_oHPukJZ31_2;
	wire w_dff_B_q8jcn1tp2_2;
	wire w_dff_B_Ep9cpCXH0_1;
	wire w_dff_B_3ltbbv398_2;
	wire w_dff_B_bocfXfef2_2;
	wire w_dff_B_GaYdGWsG5_2;
	wire w_dff_B_q9gaTcDu3_2;
	wire w_dff_B_0QW5N3qY0_2;
	wire w_dff_B_Aowu6DMd5_2;
	wire w_dff_B_GvFDmbse0_2;
	wire w_dff_B_HdTcVjcR1_2;
	wire w_dff_B_0JOnG4MU9_2;
	wire w_dff_B_yVQYx5ct9_2;
	wire w_dff_B_pMrb1zjr9_2;
	wire w_dff_B_w9qkHa0X9_2;
	wire w_dff_B_0wIZXfFx6_2;
	wire w_dff_B_htGTtLG31_2;
	wire w_dff_B_SMleNtAW7_2;
	wire w_dff_B_E2neHheu8_2;
	wire w_dff_B_Rmk0nzYJ5_2;
	wire w_dff_B_4zsRuMEd9_2;
	wire w_dff_B_qy0GjkrA5_2;
	wire w_dff_B_9qLTKO0M8_2;
	wire w_dff_B_c8bSl9KV5_1;
	wire w_dff_B_niqKiDNW8_1;
	wire w_dff_B_p0P3BqH15_2;
	wire w_dff_B_I62c8JQI2_2;
	wire w_dff_B_28qhwm4P8_2;
	wire w_dff_B_D3dcFmjD0_2;
	wire w_dff_B_C1Fw9SYq6_2;
	wire w_dff_B_CEKibw6u6_2;
	wire w_dff_B_36SM1F5p9_2;
	wire w_dff_B_UVad4XiN1_2;
	wire w_dff_B_pX10OgSl7_2;
	wire w_dff_B_7Ffryffh8_2;
	wire w_dff_B_f6WdYUHc7_2;
	wire w_dff_B_P76XU3xn8_2;
	wire w_dff_B_WGSPOU760_2;
	wire w_dff_B_Nbcylzl11_2;
	wire w_dff_B_nI0JwNwB0_2;
	wire w_dff_B_NAIdpmZ68_2;
	wire w_dff_B_6BAj7eS14_2;
	wire w_dff_B_YNZ0gsHV9_2;
	wire w_dff_B_C5oaDWd87_2;
	wire w_dff_B_sTy8tjPG0_2;
	wire w_dff_B_oGCyOuvB8_2;
	wire w_dff_B_dWMT7Lpx4_2;
	wire w_dff_B_EfmG8clW0_2;
	wire w_dff_B_qAGUZoC20_2;
	wire w_dff_B_M8j8a8cD8_2;
	wire w_dff_B_6vxfeEe18_2;
	wire w_dff_B_HnYbGdPz3_2;
	wire w_dff_B_rMASGJuo7_2;
	wire w_dff_B_qFvWF0m06_2;
	wire w_dff_B_Y2SThVqk4_2;
	wire w_dff_B_xGwlfjck2_2;
	wire w_dff_B_QP6s4kkk8_2;
	wire w_dff_B_5g7jLAsm7_2;
	wire w_dff_B_djCIo45C6_2;
	wire w_dff_B_EiNPJyiw2_2;
	wire w_dff_B_5rhA6zGm7_2;
	wire w_dff_B_AqizxOau4_1;
	wire w_dff_B_nz9DrSU60_2;
	wire w_dff_B_ntXv2OJM3_2;
	wire w_dff_B_PG7YBjra7_2;
	wire w_dff_B_5aRFOs3S3_2;
	wire w_dff_B_VoPP6YrR0_2;
	wire w_dff_B_vEotDmyG3_2;
	wire w_dff_B_Yq6fbw8A8_2;
	wire w_dff_B_LZG5QkFe4_2;
	wire w_dff_B_YLNYEWHh0_2;
	wire w_dff_B_6ywo4OgW3_2;
	wire w_dff_B_wsuBI3Td1_2;
	wire w_dff_B_jt55LJ7J9_2;
	wire w_dff_B_1vZzD2DW9_2;
	wire w_dff_B_wxBL12NL9_2;
	wire w_dff_B_Hw4blZWM1_2;
	wire w_dff_B_dS6gl4Jj2_2;
	wire w_dff_B_YDaxvvi08_2;
	wire w_dff_B_PgfjzkDW5_2;
	wire w_dff_B_w3UW7JaH0_1;
	wire w_dff_B_DIHpMLGD7_1;
	wire w_dff_B_S7miAAlE2_2;
	wire w_dff_B_IUVelolb2_2;
	wire w_dff_B_BtC00bdT3_2;
	wire w_dff_B_EZgn3QZ04_2;
	wire w_dff_B_eLLo6tPw3_2;
	wire w_dff_B_24l28blo8_2;
	wire w_dff_B_nbQo6sYz5_2;
	wire w_dff_B_vAaQu0rq1_2;
	wire w_dff_B_ZRGZ9G752_2;
	wire w_dff_B_siqKQiPV5_2;
	wire w_dff_B_jOZ1XtX40_2;
	wire w_dff_B_kHxt7nel9_2;
	wire w_dff_B_HYsBGq0B0_2;
	wire w_dff_B_tkPmTYjn8_2;
	wire w_dff_B_BxPtfmVg5_2;
	wire w_dff_B_XquK6lfj3_2;
	wire w_dff_B_pgm5CIOg2_2;
	wire w_dff_B_q5f0g6KW4_2;
	wire w_dff_B_JlVxxxPi2_2;
	wire w_dff_B_GJtcJ5q20_2;
	wire w_dff_B_BNAFJrX09_2;
	wire w_dff_B_Zaa1qRCy2_2;
	wire w_dff_B_rpMtXSaV3_2;
	wire w_dff_B_GHJChAcJ6_2;
	wire w_dff_B_WpxNynRH4_2;
	wire w_dff_B_tYLlUs1z0_2;
	wire w_dff_B_Iu5vrsMQ1_2;
	wire w_dff_B_BP1LWsrF9_2;
	wire w_dff_B_aeNosS844_1;
	wire w_dff_B_gz4ugIcs0_2;
	wire w_dff_B_0ZlW6rUd3_2;
	wire w_dff_B_iij9tUrU4_2;
	wire w_dff_B_4vgmQj8H5_2;
	wire w_dff_B_zejx364E6_2;
	wire w_dff_B_mLmBGkIA4_2;
	wire w_dff_B_oY9Nxm7D8_2;
	wire w_dff_B_gK4EYb8k8_2;
	wire w_dff_B_vpbQY6bd2_2;
	wire w_dff_B_ruSHOu9E3_2;
	wire w_dff_B_PMHAVfwd9_2;
	wire w_dff_B_LU2xYyHE0_2;
	wire w_dff_B_u6FExlep8_2;
	wire w_dff_B_DnRcI9J06_2;
	wire w_dff_B_vLBFI7kX2_2;
	wire w_dff_B_OJa5jAA83_2;
	wire w_dff_B_OFzGlZfO7_1;
	wire w_dff_B_SD9sF0Cs1_1;
	wire w_dff_B_QaLurC0e0_2;
	wire w_dff_B_bpSmEV1q8_2;
	wire w_dff_B_J7EFGDsQ1_2;
	wire w_dff_B_OX3vOu7t7_2;
	wire w_dff_B_7bXp8v1W7_2;
	wire w_dff_B_37Ba0chz7_2;
	wire w_dff_B_2KlZSCcS2_2;
	wire w_dff_B_TbL9iLmj7_2;
	wire w_dff_B_0k8pGfeg4_2;
	wire w_dff_B_mPD3MaaR6_2;
	wire w_dff_B_HvS5g1lJ0_2;
	wire w_dff_B_7IvXLYJf4_2;
	wire w_dff_B_APs3vc0s8_2;
	wire w_dff_B_CIjp0FNg9_2;
	wire w_dff_B_yr5QtQdn2_2;
	wire w_dff_B_ucHTXldm6_2;
	wire w_dff_B_R6DVXZaE2_2;
	wire w_dff_B_qGvxvP9i8_2;
	wire w_dff_B_QVDCbL2V2_2;
	wire w_dff_B_VjTNHORE0_2;
	wire w_dff_B_5fzawKms6_1;
	wire w_dff_B_wsTcT6Du0_2;
	wire w_dff_B_7r0mPeHX4_2;
	wire w_dff_B_N2I7r5sW2_2;
	wire w_dff_B_UF2C35uT0_2;
	wire w_dff_B_aCqy50DP1_2;
	wire w_dff_B_JOJvbckc7_2;
	wire w_dff_B_pdwwQ1TC8_2;
	wire w_dff_B_gN1PgTyV2_2;
	wire w_dff_B_LoTTiBbr1_2;
	wire w_dff_B_lBt4bscN8_2;
	wire w_dff_B_dsSb6e5W5_2;
	wire w_dff_B_1KLaqIJr5_2;
	wire w_dff_B_RbHQ6WDG5_2;
	wire w_dff_B_gbsWdu792_2;
	wire w_dff_B_xBcfH5Hk6_2;
	wire w_dff_B_SmC5t9hb1_2;
	wire w_dff_B_VHvBBpfl8_2;
	wire w_dff_B_k7SHEqls8_2;
	wire w_dff_B_PJgaHfRU1_2;
	wire w_dff_B_NO34ytKQ1_2;
	wire w_dff_B_UIoTEzfY3_2;
	wire w_dff_B_Hs3Qj9xI6_2;
	wire w_dff_B_dj0bbnkz3_2;
	wire w_dff_B_w1LqP5Ba0_2;
	wire w_dff_B_9AOZzDh31_2;
	wire w_dff_B_nWASdzTi0_2;
	wire w_dff_B_Kvu2NZ8E1_1;
	wire w_dff_B_b7VkWaVq0_2;
	wire w_dff_B_mkivJK7r1_2;
	wire w_dff_B_VUMyWcSP6_2;
	wire w_dff_B_5JAcsR253_2;
	wire w_dff_B_jomUdwLt9_2;
	wire w_dff_B_XFWsS37N1_2;
	wire w_dff_B_WfJUC5Th7_2;
	wire w_dff_B_rHluWfOf0_2;
	wire w_dff_B_PuzwdCvi4_2;
	wire w_dff_B_pUoWxrfk5_2;
	wire w_dff_B_P1VSDqeu3_2;
	wire w_dff_B_uSkMMjTT2_2;
	wire w_dff_B_zSwb67hh5_2;
	wire w_dff_B_4QMQO2HH8_2;
	wire w_dff_B_lQTeKuBM6_2;
	wire w_dff_A_FudOx7h20_0;
	wire w_dff_A_4HSIEWTC5_0;
	wire w_dff_A_CQ0L2kB03_0;
	wire w_dff_B_pWjCZ7xu6_2;
	wire w_dff_A_UzGkmPuH7_0;
	wire w_dff_A_MSQpi08P7_0;
	wire w_dff_A_kM3WLGk62_0;
	wire w_dff_B_4DEEQ4gN5_2;
	wire w_dff_A_cIGZ47B76_0;
	wire w_dff_A_ZGZ8rWrU5_0;
	wire w_dff_B_rJjPETkF3_2;
	wire w_dff_B_iwILiT0Z8_2;
	wire w_dff_B_6xdhJ48v5_2;
	wire w_dff_A_SBHDbXIx1_1;
	wire w_dff_A_4gQ9ZUKu3_0;
	wire w_dff_A_pPQigq9M5_0;
	wire w_dff_A_eI17mUKL4_0;
	wire w_dff_A_PdpyK4ry0_0;
	wire w_dff_A_LljHSyni0_0;
	wire w_dff_A_YeHL9aIy8_0;
	wire w_dff_A_7Y8JO7ZJ2_0;
	wire w_dff_A_iPlPA2Ip5_0;
	wire w_dff_A_zo0549vH2_0;
	wire w_dff_A_QYQci1fk0_0;
	wire w_dff_A_OiAZEN2v0_0;
	wire w_dff_A_vDxG6o7n8_0;
	wire w_dff_A_kBEVpuim4_0;
	wire w_dff_A_nhrO4Cok2_0;
	wire w_dff_A_IcvCZ8672_0;
	wire w_dff_A_tltlAlJX5_0;
	wire w_dff_A_8G0ZVXKd4_0;
	wire w_dff_A_vb3okClZ5_0;
	wire w_dff_A_vQku3r5r0_0;
	wire w_dff_A_8rg70ohz8_0;
	wire w_dff_A_3n7Q4p9d4_0;
	wire w_dff_A_y7Vu8jfj0_0;
	wire w_dff_A_9Eor3Hjo5_0;
	wire w_dff_A_1otuXqZt4_0;
	wire w_dff_A_6VIoMdNo0_0;
	wire w_dff_A_xhkOA6d50_0;
	wire w_dff_A_OlotAoqD8_0;
	wire w_dff_A_Fj4mPkYJ5_0;
	wire w_dff_A_dd4IHaLo4_0;
	wire w_dff_A_vttlEuDG3_0;
	wire w_dff_A_XFPGfoyo9_0;
	wire w_dff_A_0GuCBN7h6_0;
	wire w_dff_A_fzMSTGnW4_0;
	wire w_dff_A_Lq5pI89p4_0;
	wire w_dff_A_3aywD2BY3_0;
	wire w_dff_A_BvpnkpUv4_0;
	wire w_dff_A_p8qqB4hC7_0;
	wire w_dff_A_MWZThVTg6_0;
	wire w_dff_A_OW6khchs0_0;
	wire w_dff_A_LD4LPZq52_0;
	wire w_dff_A_u9QVAb9v2_0;
	wire w_dff_A_JoN3L7Ym8_0;
	wire w_dff_A_wn67Koel0_0;
	wire w_dff_A_80IDQ1SK6_0;
	wire w_dff_A_lJavKu555_0;
	wire w_dff_A_IhD23cpZ7_0;
	wire w_dff_A_GkZLiVdJ6_0;
	wire w_dff_A_PJj3rKIH7_0;
	wire w_dff_A_0vxVuywM2_0;
	wire w_dff_A_IsojOi9V4_0;
	wire w_dff_A_RBtRBIYw7_0;
	wire w_dff_A_DxGRfkrQ7_0;
	wire w_dff_A_er8aXkTg5_0;
	wire w_dff_A_6ntCjEA50_0;
	wire w_dff_A_WxxUDhz89_0;
	wire w_dff_A_AsbJXWKL8_0;
	wire w_dff_A_xIqktCFN7_0;
	wire w_dff_A_MKLHHGtO8_0;
	wire w_dff_A_15MuG5kP2_0;
	wire w_dff_A_oOvTVNbi6_0;
	wire w_dff_A_y0Lfbng75_0;
	wire w_dff_A_pw8NBRHb1_0;
	wire w_dff_A_h5p1L6Im0_0;
	wire w_dff_A_SXdZkzCK8_0;
	wire w_dff_A_WHkIXC9S7_0;
	wire w_dff_A_PRlghX754_0;
	wire w_dff_A_890P4iKA2_0;
	wire w_dff_A_rDYz4CU07_0;
	wire w_dff_A_5GQGx5pO5_0;
	wire w_dff_A_ooBTxhM42_0;
	wire w_dff_A_ohbgeCYa9_0;
	wire w_dff_A_JVsAVccg2_0;
	wire w_dff_A_tJS67BLc6_0;
	wire w_dff_A_TXpAQk9U3_2;
	wire w_dff_A_vRJlwoKH4_0;
	wire w_dff_A_C73LlL5J4_0;
	wire w_dff_A_yFw1wAaJ8_0;
	wire w_dff_A_rw9zDxdR1_0;
	wire w_dff_A_6hyZpext7_0;
	wire w_dff_A_Sbe3YF118_0;
	wire w_dff_A_KQCOlCla5_0;
	wire w_dff_A_2TrdDXiy6_0;
	wire w_dff_A_NWvETIUF0_0;
	wire w_dff_A_T1wKX3wU2_0;
	wire w_dff_A_NAQK3TVa0_0;
	wire w_dff_A_cszTkADn4_0;
	wire w_dff_A_unkegTzu8_0;
	wire w_dff_A_jSaQJkPg7_0;
	wire w_dff_A_tew7kQNq2_0;
	wire w_dff_A_7HqJiyOl4_0;
	wire w_dff_A_ZwjQEB1m5_0;
	wire w_dff_A_ke1r9i094_0;
	wire w_dff_A_csbgERdT2_0;
	wire w_dff_A_Evb8SzQx3_0;
	wire w_dff_A_F6cmjWKV8_0;
	wire w_dff_A_AiXJQjp85_0;
	wire w_dff_A_tuzudz8Y8_0;
	wire w_dff_A_0ExLSiUF7_0;
	wire w_dff_A_P4W3ewrv5_0;
	wire w_dff_A_HJyifzUq5_0;
	wire w_dff_A_GtoYfMj76_0;
	wire w_dff_A_V3EB6ZcX4_0;
	wire w_dff_A_W1dEsIh73_0;
	wire w_dff_A_CkV3fprj9_0;
	wire w_dff_A_20HUvyKL2_0;
	wire w_dff_A_htP9gWyX3_0;
	wire w_dff_A_PhEvehmV8_0;
	wire w_dff_A_sMZeNh7a9_0;
	wire w_dff_A_Fv68ae0f3_0;
	wire w_dff_A_D6UvXoZM2_0;
	wire w_dff_A_1EVHpBAP4_0;
	wire w_dff_A_mniHZ3B98_0;
	wire w_dff_A_Eb114fix2_0;
	wire w_dff_A_K5RERxYj4_0;
	wire w_dff_A_KUtIuPcF4_0;
	wire w_dff_A_RS0rcUYA9_0;
	wire w_dff_A_lAIycoQE7_0;
	wire w_dff_A_7gBGe5ps6_0;
	wire w_dff_A_BdaQd5Rb9_0;
	wire w_dff_A_dbATNVWm6_0;
	wire w_dff_A_tBVi5mJQ8_0;
	wire w_dff_A_INDGoFkg3_0;
	wire w_dff_A_2tnSaPAX0_0;
	wire w_dff_A_epFCYmGl7_0;
	wire w_dff_A_EsqYMR8O7_0;
	wire w_dff_A_zs9xhk1c1_0;
	wire w_dff_A_SShDmPL80_0;
	wire w_dff_A_UXcMNORi3_0;
	wire w_dff_A_T0mmnZeG6_0;
	wire w_dff_A_EEkZZj2h4_0;
	wire w_dff_A_rOD5n1Y23_0;
	wire w_dff_A_VBddhrBH2_0;
	wire w_dff_A_rOO9VspZ6_0;
	wire w_dff_A_CPjkiGVQ2_0;
	wire w_dff_A_AL20DwRz2_0;
	wire w_dff_A_vwszhUu81_0;
	wire w_dff_A_81v8lyms0_0;
	wire w_dff_A_WLCOgiXJ7_0;
	wire w_dff_A_0Lq0JNAS8_0;
	wire w_dff_A_vRK7OhD86_0;
	wire w_dff_A_q6O0bSP29_0;
	wire w_dff_A_lamaJPT51_0;
	wire w_dff_A_blGfFtq53_0;
	wire w_dff_A_buo4FdL10_2;
	wire w_dff_A_TXQDmXQu9_0;
	wire w_dff_A_poLHy51T9_0;
	wire w_dff_A_G7Yi1Tj75_0;
	wire w_dff_A_JBM5vqQf6_0;
	wire w_dff_A_WaoXTjPl0_0;
	wire w_dff_A_WOiBWxin6_0;
	wire w_dff_A_X7s0jOUv1_0;
	wire w_dff_A_NBJwJOM78_0;
	wire w_dff_A_7Q7l75KR3_0;
	wire w_dff_A_95RTOtd64_0;
	wire w_dff_A_smRvgRlM3_0;
	wire w_dff_A_IScTT8RI7_0;
	wire w_dff_A_kwZ2gT2t5_0;
	wire w_dff_A_zbTTgX4P1_0;
	wire w_dff_A_WijUF9467_0;
	wire w_dff_A_g0eAg3Co1_0;
	wire w_dff_A_57ZLz1p54_0;
	wire w_dff_A_Ie2YxNOe9_0;
	wire w_dff_A_rmuaJVc84_0;
	wire w_dff_A_kW8m9Uc21_0;
	wire w_dff_A_7hQEarXC6_0;
	wire w_dff_A_NsfJuRvx0_0;
	wire w_dff_A_lySbVBV65_0;
	wire w_dff_A_AhkEpVkb3_0;
	wire w_dff_A_AARyv2OZ4_0;
	wire w_dff_A_nv6ZFavq7_0;
	wire w_dff_A_fIYMeOPI7_0;
	wire w_dff_A_FMlrkncn3_0;
	wire w_dff_A_seEZ09Bf8_0;
	wire w_dff_A_XvhIP3zA9_0;
	wire w_dff_A_CqixKKVX0_0;
	wire w_dff_A_gz1GsxHp5_0;
	wire w_dff_A_Tyj5oO2W9_0;
	wire w_dff_A_R7C45UMu6_0;
	wire w_dff_A_kyvCI4jS6_0;
	wire w_dff_A_hdGFVPii0_0;
	wire w_dff_A_mAfEbpZI0_0;
	wire w_dff_A_CoeC1kwg1_0;
	wire w_dff_A_IGxYFOR93_0;
	wire w_dff_A_Vw5fECnz2_0;
	wire w_dff_A_WpnxNDUE8_0;
	wire w_dff_A_1YDCgfkD9_0;
	wire w_dff_A_OLAfH0io7_0;
	wire w_dff_A_jBE172ew3_0;
	wire w_dff_A_LmlYMnMJ8_0;
	wire w_dff_A_Gr02eWPc5_0;
	wire w_dff_A_l8jeQ4254_0;
	wire w_dff_A_JBUAY8Fw0_0;
	wire w_dff_A_6zutFgaU6_0;
	wire w_dff_A_rp2XgVWh3_0;
	wire w_dff_A_6wZbilJl2_0;
	wire w_dff_A_GnMpStnz1_0;
	wire w_dff_A_cMcUBohz8_0;
	wire w_dff_A_UI1R9Le08_0;
	wire w_dff_A_w8sKohNk5_0;
	wire w_dff_A_zlcWMyib6_0;
	wire w_dff_A_O0SO8ROF3_0;
	wire w_dff_A_MdHWVO2B3_0;
	wire w_dff_A_paKgfGkd1_0;
	wire w_dff_A_c4TVz89o2_0;
	wire w_dff_A_wGpiu0r74_0;
	wire w_dff_A_U6lDBDTs0_0;
	wire w_dff_A_ZI9Vowwm3_0;
	wire w_dff_A_DHpCUB6Q1_0;
	wire w_dff_A_yKS96IHA5_0;
	wire w_dff_A_yyGiPMnY0_0;
	wire w_dff_A_vUbw6a1X3_0;
	wire w_dff_A_5QNzbAT64_0;
	wire w_dff_A_dMBLpPmk9_2;
	wire w_dff_A_w7Qg4Ogm6_0;
	wire w_dff_A_aAxv4qMc1_0;
	wire w_dff_A_ItSyCivU4_0;
	wire w_dff_A_KceAzcYC0_0;
	wire w_dff_A_DJaz2nfu9_0;
	wire w_dff_A_DL4jujl76_0;
	wire w_dff_A_M7REda1w2_0;
	wire w_dff_A_T7K3CaY87_0;
	wire w_dff_A_hmRtgyuR3_0;
	wire w_dff_A_0sdC5CQt8_0;
	wire w_dff_A_3ho92WB04_0;
	wire w_dff_A_Ytp4l8vM7_0;
	wire w_dff_A_mEgezkWX4_0;
	wire w_dff_A_n0dU0Hwf3_0;
	wire w_dff_A_sANRdrOi4_0;
	wire w_dff_A_VoeJeHDR0_0;
	wire w_dff_A_R5d8JNCG8_0;
	wire w_dff_A_LkTXmiTN2_0;
	wire w_dff_A_44b5Za3q0_0;
	wire w_dff_A_65S7st0f9_0;
	wire w_dff_A_qez06FdT3_0;
	wire w_dff_A_jIfjbs3p4_0;
	wire w_dff_A_Lp23YidW0_0;
	wire w_dff_A_liEFXoqg6_0;
	wire w_dff_A_iSUWP2vl4_0;
	wire w_dff_A_0VBGkh5x9_0;
	wire w_dff_A_shQg4kMP0_0;
	wire w_dff_A_i74p85CP1_0;
	wire w_dff_A_htM5lZks8_0;
	wire w_dff_A_6VIPgpEI3_0;
	wire w_dff_A_mpJjQPkg4_0;
	wire w_dff_A_OO8pCVS49_0;
	wire w_dff_A_mSmIWK7j9_0;
	wire w_dff_A_u0gJUiq52_0;
	wire w_dff_A_y9xN8TYu4_0;
	wire w_dff_A_Sr626VtM9_0;
	wire w_dff_A_adCT9SwV1_0;
	wire w_dff_A_79qyOkIc4_0;
	wire w_dff_A_yWsc2FG58_0;
	wire w_dff_A_XvVgFn9P0_0;
	wire w_dff_A_pBRyccUm1_0;
	wire w_dff_A_urcuM0of9_0;
	wire w_dff_A_YsSHIPp28_0;
	wire w_dff_A_vL4YCkmB6_0;
	wire w_dff_A_7ao35V7m9_0;
	wire w_dff_A_KPVd0E3G7_0;
	wire w_dff_A_C84v9WI28_0;
	wire w_dff_A_merpgjMT5_0;
	wire w_dff_A_i29UEyo96_0;
	wire w_dff_A_6Ljx9aGY4_0;
	wire w_dff_A_8WYA2Jd19_0;
	wire w_dff_A_waG2YfAb8_0;
	wire w_dff_A_MZG1aCZA7_0;
	wire w_dff_A_sqbHbFPC4_0;
	wire w_dff_A_LS7bFTju7_0;
	wire w_dff_A_RZtG7oBe2_0;
	wire w_dff_A_Lo4r26GP1_0;
	wire w_dff_A_XNimF5mI3_0;
	wire w_dff_A_48zxiKJh3_0;
	wire w_dff_A_HXAkp2Hr2_0;
	wire w_dff_A_D98vrOpP9_0;
	wire w_dff_A_SbpdLbA98_0;
	wire w_dff_A_vjiFzC1H3_0;
	wire w_dff_A_O6hg4Dry9_0;
	wire w_dff_A_7yE0NEGK3_0;
	wire w_dff_A_gefk1wav5_2;
	wire w_dff_A_DWMixp4U9_0;
	wire w_dff_A_yy540UXo8_0;
	wire w_dff_A_qRfJJhsW8_0;
	wire w_dff_A_oTtkERGX3_0;
	wire w_dff_A_5waJCCo93_0;
	wire w_dff_A_9QY3BGhr5_0;
	wire w_dff_A_U5OLYsr97_0;
	wire w_dff_A_pRcNIFEJ4_0;
	wire w_dff_A_ABzoDVs39_0;
	wire w_dff_A_pFZUHEKQ7_0;
	wire w_dff_A_w4Aj6XlB2_0;
	wire w_dff_A_yIzZqKfb5_0;
	wire w_dff_A_kTaoyh0S4_0;
	wire w_dff_A_BHdxHAt01_0;
	wire w_dff_A_EErckhbs1_0;
	wire w_dff_A_5n9ZpK7C5_0;
	wire w_dff_A_vDpKBRS55_0;
	wire w_dff_A_xY2YEdT17_0;
	wire w_dff_A_O1FQhSMu2_0;
	wire w_dff_A_KwVgtCfR3_0;
	wire w_dff_A_X8hL8fkt7_0;
	wire w_dff_A_UJpwuqi06_0;
	wire w_dff_A_KPqNtckk9_0;
	wire w_dff_A_Zuq8soWV9_0;
	wire w_dff_A_aVzL60u73_0;
	wire w_dff_A_2XcVAt7h1_0;
	wire w_dff_A_vi7yjqHw6_0;
	wire w_dff_A_IOKbtvmm5_0;
	wire w_dff_A_nValV1yi1_0;
	wire w_dff_A_cYohB2Ig3_0;
	wire w_dff_A_fcy7mX9L5_0;
	wire w_dff_A_rV90dYuF4_0;
	wire w_dff_A_IS1vNVL88_0;
	wire w_dff_A_8ObDaeqV8_0;
	wire w_dff_A_NJuuxCSy0_0;
	wire w_dff_A_tExBP91x7_0;
	wire w_dff_A_fK22dD7y6_0;
	wire w_dff_A_kQuEI4zD7_0;
	wire w_dff_A_WdTMREwU5_0;
	wire w_dff_A_fbPW6fY64_0;
	wire w_dff_A_I40QanF71_0;
	wire w_dff_A_KHz6G9TZ1_0;
	wire w_dff_A_EDJQ5LCw3_0;
	wire w_dff_A_UaAQEaEB1_0;
	wire w_dff_A_cKcQoA330_0;
	wire w_dff_A_xLl8ZBKx4_0;
	wire w_dff_A_Hy0Ia5YF8_0;
	wire w_dff_A_MiTYFQNb2_0;
	wire w_dff_A_ej3NMY796_0;
	wire w_dff_A_zQLlC5Jg5_0;
	wire w_dff_A_vGJVRWXF6_0;
	wire w_dff_A_dbq52p2K5_0;
	wire w_dff_A_wtIb7jUO1_0;
	wire w_dff_A_aODrlKhT3_0;
	wire w_dff_A_v01lq88z1_0;
	wire w_dff_A_iVSpAhTK7_0;
	wire w_dff_A_7WfemrKq0_0;
	wire w_dff_A_IgrKJTUo6_0;
	wire w_dff_A_8ZFaHYJb2_0;
	wire w_dff_A_Z8lnYFP37_0;
	wire w_dff_A_x5RKSedm6_0;
	wire w_dff_A_YIn3qLDg7_0;
	wire w_dff_A_4JhpDJQk1_2;
	wire w_dff_A_nscWjhLV4_0;
	wire w_dff_A_QQtvKVR79_0;
	wire w_dff_A_zwrkMT7A1_0;
	wire w_dff_A_QwIXjRXM8_0;
	wire w_dff_A_CQnTGkZN9_0;
	wire w_dff_A_FF4UYeuX9_0;
	wire w_dff_A_bo9Idjg63_0;
	wire w_dff_A_alVAfPKn5_0;
	wire w_dff_A_0B793M7y4_0;
	wire w_dff_A_hmCun4bB8_0;
	wire w_dff_A_05M9lXxp1_0;
	wire w_dff_A_CIi0AJt59_0;
	wire w_dff_A_7tYKSSNk7_0;
	wire w_dff_A_AH7xB5E76_0;
	wire w_dff_A_K7xAnZbI1_0;
	wire w_dff_A_2MQGX1sc5_0;
	wire w_dff_A_BXAf8yXK6_0;
	wire w_dff_A_NSmRaWpA6_0;
	wire w_dff_A_6S5w8DWx4_0;
	wire w_dff_A_bLq4l5x63_0;
	wire w_dff_A_15wk6lWG7_0;
	wire w_dff_A_npCZH30I8_0;
	wire w_dff_A_lEqnh4SU5_0;
	wire w_dff_A_pqHE9Al20_0;
	wire w_dff_A_xRpkV9632_0;
	wire w_dff_A_vCbl7ueO9_0;
	wire w_dff_A_MDG60FCl4_0;
	wire w_dff_A_3ohWSRwp6_0;
	wire w_dff_A_JpKvjN0Q8_0;
	wire w_dff_A_8ctyCZPs9_0;
	wire w_dff_A_dQW0Y0CM0_0;
	wire w_dff_A_lIMMJ4mF0_0;
	wire w_dff_A_X3aSuwpr7_0;
	wire w_dff_A_So9rCyCz4_0;
	wire w_dff_A_0UJhvR7F7_0;
	wire w_dff_A_XMy9xEqY6_0;
	wire w_dff_A_mKHUZWye9_0;
	wire w_dff_A_wWWm1iD94_0;
	wire w_dff_A_lzbFtxis8_0;
	wire w_dff_A_LcacxyjB4_0;
	wire w_dff_A_pajuTJ4l9_0;
	wire w_dff_A_gajrwyFc3_0;
	wire w_dff_A_UbCLgaYO7_0;
	wire w_dff_A_XSaSblFD4_0;
	wire w_dff_A_q5LOD2tg7_0;
	wire w_dff_A_diZSij045_0;
	wire w_dff_A_Ah9bIosR8_0;
	wire w_dff_A_X2xmfMcN5_0;
	wire w_dff_A_2stJmJAI3_0;
	wire w_dff_A_C3F1ytOH2_0;
	wire w_dff_A_IRQLmgfl1_0;
	wire w_dff_A_33pAvLiG4_0;
	wire w_dff_A_VDOZAGKJ3_0;
	wire w_dff_A_D67H8ryT4_0;
	wire w_dff_A_ZcD82bRK2_0;
	wire w_dff_A_gffDqlbO2_0;
	wire w_dff_A_jMtAlfG86_0;
	wire w_dff_A_PIQxSxvV7_0;
	wire w_dff_A_V5ARinu60_0;
	wire w_dff_A_fzty24Fg7_2;
	wire w_dff_A_6iTRBODh0_0;
	wire w_dff_A_m3ufP3LF0_0;
	wire w_dff_A_22qSoX7d0_0;
	wire w_dff_A_ijIFejDa8_0;
	wire w_dff_A_RMJAOgWq7_0;
	wire w_dff_A_OOkiQ2DN0_0;
	wire w_dff_A_1nyx4VDY1_0;
	wire w_dff_A_gKZFgW2Y3_0;
	wire w_dff_A_bSzpXqiR9_0;
	wire w_dff_A_vxA7COBK1_0;
	wire w_dff_A_AGXvGq6D7_0;
	wire w_dff_A_KINI6req8_0;
	wire w_dff_A_EAgXLHIO1_0;
	wire w_dff_A_2KUCl9DI3_0;
	wire w_dff_A_8NgEBRJE8_0;
	wire w_dff_A_R16Af9wA2_0;
	wire w_dff_A_dlri9R6W5_0;
	wire w_dff_A_uXKjIZUZ8_0;
	wire w_dff_A_ocPFOu4n9_0;
	wire w_dff_A_3GNKu7tj4_0;
	wire w_dff_A_6Klz3CAM9_0;
	wire w_dff_A_d9dXtT5D1_0;
	wire w_dff_A_Y45WbqMa1_0;
	wire w_dff_A_94PULiMl6_0;
	wire w_dff_A_VnGbh9Xj3_0;
	wire w_dff_A_wRWZrKDl9_0;
	wire w_dff_A_rTm3ETE66_0;
	wire w_dff_A_cMnCFvqz6_0;
	wire w_dff_A_EqIcwaNl4_0;
	wire w_dff_A_PYTHsVSV6_0;
	wire w_dff_A_zW3StyU38_0;
	wire w_dff_A_TiiRIfM07_0;
	wire w_dff_A_Z8m1LNur4_0;
	wire w_dff_A_pDxQtBqK4_0;
	wire w_dff_A_Xxxmtu9M9_0;
	wire w_dff_A_v1i21oW54_0;
	wire w_dff_A_Q3nwZ8B10_0;
	wire w_dff_A_SxpUWssj6_0;
	wire w_dff_A_8oG1HlPz7_0;
	wire w_dff_A_XuZzfXVF6_0;
	wire w_dff_A_Pwa9WOzs5_0;
	wire w_dff_A_PfzGn3X40_0;
	wire w_dff_A_BfQIop7N9_0;
	wire w_dff_A_3Wp3jCBv0_0;
	wire w_dff_A_zOl2rtiz9_0;
	wire w_dff_A_yjXakVSd2_0;
	wire w_dff_A_uAUxLrQH5_0;
	wire w_dff_A_ySqeQT9u0_0;
	wire w_dff_A_tTPD9ViQ9_0;
	wire w_dff_A_S5aMvSkZ1_0;
	wire w_dff_A_Aj89iEXp0_0;
	wire w_dff_A_i15bLFzL8_0;
	wire w_dff_A_r47pQr0d3_0;
	wire w_dff_A_DcnzQsiz7_0;
	wire w_dff_A_9mk7is8K3_0;
	wire w_dff_A_68phYQ4d9_0;
	wire w_dff_A_1S7EK9uC0_2;
	wire w_dff_A_HPUO8x400_0;
	wire w_dff_A_WC9m3MTH6_0;
	wire w_dff_A_yV6upp311_0;
	wire w_dff_A_NkTNLiv69_0;
	wire w_dff_A_TEWSREFY8_0;
	wire w_dff_A_hahDbAXu3_0;
	wire w_dff_A_QqVaIVsn3_0;
	wire w_dff_A_kPlYeg6T3_0;
	wire w_dff_A_88CXVLny9_0;
	wire w_dff_A_pln3Ak7p8_0;
	wire w_dff_A_C6QyKAcU4_0;
	wire w_dff_A_V3wRKQ6T0_0;
	wire w_dff_A_vspatCTH4_0;
	wire w_dff_A_ONKKmu3q0_0;
	wire w_dff_A_dFA43SZV8_0;
	wire w_dff_A_zgdFauPo1_0;
	wire w_dff_A_2gmMJMzL1_0;
	wire w_dff_A_V79hsKxC5_0;
	wire w_dff_A_swYR5ZIm2_0;
	wire w_dff_A_1QJpCATX3_0;
	wire w_dff_A_RN94JaGJ7_0;
	wire w_dff_A_UAPm7bfk6_0;
	wire w_dff_A_rfc8MkMO1_0;
	wire w_dff_A_8kmJIDCC6_0;
	wire w_dff_A_vnxznyvI0_0;
	wire w_dff_A_w36IsMES2_0;
	wire w_dff_A_J0AoCJDc7_0;
	wire w_dff_A_GLZ5Xeui5_0;
	wire w_dff_A_Wc3AONrK4_0;
	wire w_dff_A_DRa0OLxR4_0;
	wire w_dff_A_btiNppzx2_0;
	wire w_dff_A_DFFZ0xWL5_0;
	wire w_dff_A_5xZ55Ezy0_0;
	wire w_dff_A_ubRN5I0d2_0;
	wire w_dff_A_48kgtEq73_0;
	wire w_dff_A_Mo7K6gIZ5_0;
	wire w_dff_A_2EloxUDu8_0;
	wire w_dff_A_7gmrsr0L6_0;
	wire w_dff_A_BTqd9MWm2_0;
	wire w_dff_A_XzN1SUH75_0;
	wire w_dff_A_CI30zncL7_0;
	wire w_dff_A_cTzWC01n7_0;
	wire w_dff_A_nCyqUpG01_0;
	wire w_dff_A_IAwfR51o0_0;
	wire w_dff_A_mhy64e4S5_0;
	wire w_dff_A_KJnPgomu6_0;
	wire w_dff_A_Xhq0SttG8_0;
	wire w_dff_A_7uhaWb3b0_0;
	wire w_dff_A_c2T70DH62_0;
	wire w_dff_A_0NeDqDHN7_0;
	wire w_dff_A_N1CbjniU6_0;
	wire w_dff_A_RaSdH8Ma7_0;
	wire w_dff_A_uZFEBlv00_0;
	wire w_dff_A_fdK3GZD42_2;
	wire w_dff_A_D1ljxla53_0;
	wire w_dff_A_tEARLD7D6_0;
	wire w_dff_A_76c5jxDK0_0;
	wire w_dff_A_zBD61QgE5_0;
	wire w_dff_A_ztwIVD195_0;
	wire w_dff_A_46XjdZOD8_0;
	wire w_dff_A_ubCCc7Ut7_0;
	wire w_dff_A_19AlYVxb6_0;
	wire w_dff_A_7nhZJRs75_0;
	wire w_dff_A_o7mc7g1c8_0;
	wire w_dff_A_PNytZXnZ6_0;
	wire w_dff_A_pYQCQtA32_0;
	wire w_dff_A_KD3YEOd65_0;
	wire w_dff_A_EGwqlcHe5_0;
	wire w_dff_A_EoZBtHPh3_0;
	wire w_dff_A_AYNaDx281_0;
	wire w_dff_A_UMl2PSNY9_0;
	wire w_dff_A_MvOEAy0u1_0;
	wire w_dff_A_5g1JbNwe1_0;
	wire w_dff_A_UvrOH25s6_0;
	wire w_dff_A_MQ0iiGvh3_0;
	wire w_dff_A_EDcfrQLi4_0;
	wire w_dff_A_pqKVAr1L2_0;
	wire w_dff_A_h48HmMfn9_0;
	wire w_dff_A_FciaFmtN9_0;
	wire w_dff_A_Q3yKlTyM2_0;
	wire w_dff_A_jyS6FEhA3_0;
	wire w_dff_A_c87I8tIR1_0;
	wire w_dff_A_HcoYOmkU1_0;
	wire w_dff_A_dbNCtryU3_0;
	wire w_dff_A_8aYcfREe7_0;
	wire w_dff_A_0W8NKevD2_0;
	wire w_dff_A_fvZktCYV2_0;
	wire w_dff_A_d4PDu5js1_0;
	wire w_dff_A_emgBjAc66_0;
	wire w_dff_A_IcrTRLzk1_0;
	wire w_dff_A_EmEDWUDA7_0;
	wire w_dff_A_ppQja7TY5_0;
	wire w_dff_A_IBxT8tdI5_0;
	wire w_dff_A_fum6iNeP8_0;
	wire w_dff_A_JaRRQPGI6_0;
	wire w_dff_A_q1dML4Pk2_0;
	wire w_dff_A_2Jk1u5j47_0;
	wire w_dff_A_PzDEvjIy5_0;
	wire w_dff_A_IBHNEwXx5_0;
	wire w_dff_A_ksiK7KtB0_0;
	wire w_dff_A_nbbZbNnd3_0;
	wire w_dff_A_cd5jhFgd7_0;
	wire w_dff_A_yKbQ2N8Z4_0;
	wire w_dff_A_pWkdBPgJ1_0;
	wire w_dff_A_rFD3ruyP8_2;
	wire w_dff_A_wCy1wkOG8_0;
	wire w_dff_A_f8dCr8qN6_0;
	wire w_dff_A_kG6bMXmL9_0;
	wire w_dff_A_nE69rSCD7_0;
	wire w_dff_A_liYaWvap4_0;
	wire w_dff_A_YZwxnTFa8_0;
	wire w_dff_A_HYrZCvr05_0;
	wire w_dff_A_H1MTa1pn2_0;
	wire w_dff_A_WJWPnB9Q8_0;
	wire w_dff_A_2eYmAzvl3_0;
	wire w_dff_A_Lerj2lpD7_0;
	wire w_dff_A_p8WJsDxe2_0;
	wire w_dff_A_BtXZHzpo6_0;
	wire w_dff_A_T2pNZOI31_0;
	wire w_dff_A_S5XawaYp1_0;
	wire w_dff_A_AdmSjIPk7_0;
	wire w_dff_A_Rz9JcqBr3_0;
	wire w_dff_A_3R3qCcjJ9_0;
	wire w_dff_A_lTAA7f5n6_0;
	wire w_dff_A_sfwro9XK1_0;
	wire w_dff_A_OWnu9flQ8_0;
	wire w_dff_A_ueVP981F2_0;
	wire w_dff_A_t339kxfb7_0;
	wire w_dff_A_ZcDslSaE2_0;
	wire w_dff_A_kIFd3SPK5_0;
	wire w_dff_A_HtpdOZjk3_0;
	wire w_dff_A_ffaHNuvX1_0;
	wire w_dff_A_el1TYYkf6_0;
	wire w_dff_A_VXlBulOn1_0;
	wire w_dff_A_ftGxvHZw6_0;
	wire w_dff_A_jVvIQzwF0_0;
	wire w_dff_A_fnJRMVzh6_0;
	wire w_dff_A_fioCgruU3_0;
	wire w_dff_A_HcBfl0mh6_0;
	wire w_dff_A_hBewRon32_0;
	wire w_dff_A_46sTgkrF7_0;
	wire w_dff_A_ahm8CCsf0_0;
	wire w_dff_A_SitAz65p3_0;
	wire w_dff_A_wuCqWLwH1_0;
	wire w_dff_A_1OeTwyEH9_0;
	wire w_dff_A_jWvUl0xN3_0;
	wire w_dff_A_v0BdXfzU6_0;
	wire w_dff_A_yFAQckSv6_0;
	wire w_dff_A_KXkzmyTm3_0;
	wire w_dff_A_LXNOeWHW9_0;
	wire w_dff_A_YFPYsXl46_0;
	wire w_dff_A_HLXQTx3j8_0;
	wire w_dff_A_xANsDdVz6_2;
	wire w_dff_A_pXTROB3q9_0;
	wire w_dff_A_jTOenI3v4_0;
	wire w_dff_A_r8okHQLl2_0;
	wire w_dff_A_fM681KaE7_0;
	wire w_dff_A_jHmMc3Ki1_0;
	wire w_dff_A_fLjFoE160_0;
	wire w_dff_A_h0g5HjaA9_0;
	wire w_dff_A_aS2bhrfJ1_0;
	wire w_dff_A_GL7PML9S7_0;
	wire w_dff_A_obzNNO2M9_0;
	wire w_dff_A_rC9QR0lC5_0;
	wire w_dff_A_G3oFA62V3_0;
	wire w_dff_A_gPMwZevJ4_0;
	wire w_dff_A_Ahq83ELf3_0;
	wire w_dff_A_3Gxy1OxP4_0;
	wire w_dff_A_tsng1w7b9_0;
	wire w_dff_A_e9OojFyN1_0;
	wire w_dff_A_lhRRBONw1_0;
	wire w_dff_A_9K9WqwCv8_0;
	wire w_dff_A_JQlLSURC0_0;
	wire w_dff_A_fQm5pxXj3_0;
	wire w_dff_A_jgkdZ4zw3_0;
	wire w_dff_A_2UBEBqK12_0;
	wire w_dff_A_TECjVfwv6_0;
	wire w_dff_A_nSqJEH3d4_0;
	wire w_dff_A_SN8bqs2Q8_0;
	wire w_dff_A_T5LinO5h6_0;
	wire w_dff_A_IM87GUaO0_0;
	wire w_dff_A_FySOt3Ij6_0;
	wire w_dff_A_Sid51fXI9_0;
	wire w_dff_A_tcKMdUFV7_0;
	wire w_dff_A_Z1MctO2O6_0;
	wire w_dff_A_RIlCVX171_0;
	wire w_dff_A_y0kfxqN95_0;
	wire w_dff_A_YZlIMUAR2_0;
	wire w_dff_A_uMQoYzc75_0;
	wire w_dff_A_ATFtiSAo6_0;
	wire w_dff_A_9vqiQXsy9_0;
	wire w_dff_A_B3kiD3K41_0;
	wire w_dff_A_J7KP6UIZ4_0;
	wire w_dff_A_KlfMuHA29_0;
	wire w_dff_A_pIiXC78S0_0;
	wire w_dff_A_uHFALARi1_0;
	wire w_dff_A_sCnUazWe3_0;
	wire w_dff_A_k3iKXLIe4_2;
	wire w_dff_A_Aglkn81E6_0;
	wire w_dff_A_XL6evCQi0_0;
	wire w_dff_A_u11dQkLr8_0;
	wire w_dff_A_XnWeIXQY3_0;
	wire w_dff_A_VZNs2JDX5_0;
	wire w_dff_A_6aVrzrep2_0;
	wire w_dff_A_ljf05tGS0_0;
	wire w_dff_A_UrPv5nGB4_0;
	wire w_dff_A_5VnNimcs2_0;
	wire w_dff_A_Hrg1rnYa5_0;
	wire w_dff_A_QcnA24mZ2_0;
	wire w_dff_A_J2rQYll28_0;
	wire w_dff_A_n7I5sYsL8_0;
	wire w_dff_A_S9hkccD34_0;
	wire w_dff_A_lpelPjES3_0;
	wire w_dff_A_YzZJmEw44_0;
	wire w_dff_A_9lcWTbCJ1_0;
	wire w_dff_A_Ov99oSIH4_0;
	wire w_dff_A_D0caj4ux5_0;
	wire w_dff_A_bsshSqi58_0;
	wire w_dff_A_Nda5H63m0_0;
	wire w_dff_A_buRSM4VA9_0;
	wire w_dff_A_HePwnezM4_0;
	wire w_dff_A_gc1VAXFE5_0;
	wire w_dff_A_fgwJtztX6_0;
	wire w_dff_A_l2OkezNQ1_0;
	wire w_dff_A_V4m9BGio9_0;
	wire w_dff_A_WoDYBINQ3_0;
	wire w_dff_A_RwfZcAnT6_0;
	wire w_dff_A_iervmNT84_0;
	wire w_dff_A_sbxqpdEo3_0;
	wire w_dff_A_Lw05cSSz2_0;
	wire w_dff_A_GmhKQyBS2_0;
	wire w_dff_A_8zV5OEf07_0;
	wire w_dff_A_77moib451_0;
	wire w_dff_A_DOBWTF6i9_0;
	wire w_dff_A_JODvmQXA8_0;
	wire w_dff_A_J58U6LNq4_0;
	wire w_dff_A_0SptStsj3_0;
	wire w_dff_A_CXuqsHmV8_0;
	wire w_dff_A_akbihhF17_0;
	wire w_dff_A_Whz6y90z4_2;
	wire w_dff_A_HZt5ri3T9_0;
	wire w_dff_A_MjSvTIG88_0;
	wire w_dff_A_JrxqGUmX7_0;
	wire w_dff_A_42z0BhHr9_0;
	wire w_dff_A_WA9QuyfT8_0;
	wire w_dff_A_hV3B999W1_0;
	wire w_dff_A_yw5RLx8R4_0;
	wire w_dff_A_GlRNSy3p5_0;
	wire w_dff_A_Ifjcdlbu3_0;
	wire w_dff_A_sSoUT4GB2_0;
	wire w_dff_A_7z4bE0cu6_0;
	wire w_dff_A_fBj8Bayd6_0;
	wire w_dff_A_ARnkUL2z7_0;
	wire w_dff_A_phchnPF09_0;
	wire w_dff_A_AbD197dt4_0;
	wire w_dff_A_qZU0jvS74_0;
	wire w_dff_A_AC60Ks0n6_0;
	wire w_dff_A_zowmw9a57_0;
	wire w_dff_A_fwwJw1VS2_0;
	wire w_dff_A_8Kb0HGMS8_0;
	wire w_dff_A_GawTFX1o1_0;
	wire w_dff_A_1QWCMiNR1_0;
	wire w_dff_A_jCTNTG1a6_0;
	wire w_dff_A_KI8nbasE7_0;
	wire w_dff_A_wRVKJ3jY9_0;
	wire w_dff_A_4k8yGm471_0;
	wire w_dff_A_dYamHiU94_0;
	wire w_dff_A_Hb5cXusa5_0;
	wire w_dff_A_EGGfkYTS7_0;
	wire w_dff_A_T5g9g3CF7_0;
	wire w_dff_A_BPTIuZLw0_0;
	wire w_dff_A_CYdXihWS8_0;
	wire w_dff_A_JfbYWNPY1_0;
	wire w_dff_A_uYc1LZQA9_0;
	wire w_dff_A_5JzA5IOY5_0;
	wire w_dff_A_zlYlzgot0_0;
	wire w_dff_A_J77gEn0R7_0;
	wire w_dff_A_IOeZXjCa0_0;
	wire w_dff_A_dSuBmHpc5_2;
	wire w_dff_A_mdoLfKW24_0;
	wire w_dff_A_fdPLxgoC7_0;
	wire w_dff_A_p0IlcEKG9_0;
	wire w_dff_A_3Pq8IOer9_0;
	wire w_dff_A_EopLJP5f8_0;
	wire w_dff_A_aZpy6ceA4_0;
	wire w_dff_A_u2yetZ701_0;
	wire w_dff_A_XRjeNN6X4_0;
	wire w_dff_A_J9I248Jp1_0;
	wire w_dff_A_htZXRUfj3_0;
	wire w_dff_A_U4JsR3Uq9_0;
	wire w_dff_A_p6E1KrtO2_0;
	wire w_dff_A_Q1tb5loz6_0;
	wire w_dff_A_h2AvVCpa7_0;
	wire w_dff_A_bzvuPIrZ7_0;
	wire w_dff_A_yy7jIqcN3_0;
	wire w_dff_A_JlQ5wT8n6_0;
	wire w_dff_A_yxNV3cxa8_0;
	wire w_dff_A_9VucbSb85_0;
	wire w_dff_A_s7UaRNx12_0;
	wire w_dff_A_9shebP5b4_0;
	wire w_dff_A_BphnsUee2_0;
	wire w_dff_A_7MN3KpQd6_0;
	wire w_dff_A_vw1RV2NV0_0;
	wire w_dff_A_SHwyh0c18_0;
	wire w_dff_A_DDAQjcyZ1_0;
	wire w_dff_A_Dg9NJat15_0;
	wire w_dff_A_2CJ6JoJ82_0;
	wire w_dff_A_cJ2U47NJ9_0;
	wire w_dff_A_w16I4wIA3_0;
	wire w_dff_A_zwpytITb0_0;
	wire w_dff_A_EgeqZIwH2_0;
	wire w_dff_A_tjFBlMny9_0;
	wire w_dff_A_iKzjfTVX4_0;
	wire w_dff_A_6VkxC2es4_0;
	wire w_dff_A_GrvPvRzD1_2;
	wire w_dff_A_pqB8Fko46_0;
	wire w_dff_A_3f80n6Gs2_0;
	wire w_dff_A_Udra6jHd0_0;
	wire w_dff_A_034Fj5gR5_0;
	wire w_dff_A_we1nG2fK9_0;
	wire w_dff_A_8uBpOEXy0_0;
	wire w_dff_A_AFM0uJ5l6_0;
	wire w_dff_A_tqQXvXDU0_0;
	wire w_dff_A_w1ApzctC7_0;
	wire w_dff_A_ztgUPg7q4_0;
	wire w_dff_A_XwcQiECs5_0;
	wire w_dff_A_vvzIJkBd2_0;
	wire w_dff_A_ujjTKTyt5_0;
	wire w_dff_A_0To7aDDQ0_0;
	wire w_dff_A_PNOJfyzw4_0;
	wire w_dff_A_fP7OT9lk4_0;
	wire w_dff_A_v2uaTy926_0;
	wire w_dff_A_wfeZErTh7_0;
	wire w_dff_A_7m7ZrYDo0_0;
	wire w_dff_A_IIEnOhAI5_0;
	wire w_dff_A_BdpJywMH1_0;
	wire w_dff_A_OeX0mVef4_0;
	wire w_dff_A_dCOIv1RO8_0;
	wire w_dff_A_gilxwOXP8_0;
	wire w_dff_A_9s0IZ3cU9_0;
	wire w_dff_A_nd2IUhhm0_0;
	wire w_dff_A_B55TaYlr1_0;
	wire w_dff_A_hwYXCZVQ2_0;
	wire w_dff_A_K83xiXkF9_0;
	wire w_dff_A_rL6AXHc15_0;
	wire w_dff_A_kD19nGPu9_0;
	wire w_dff_A_QAAJOoP98_0;
	wire w_dff_A_b9xSmEOi6_2;
	wire w_dff_A_Xgwsrhnl1_0;
	wire w_dff_A_RzkSdMIb4_0;
	wire w_dff_A_zaboybat2_0;
	wire w_dff_A_ZlJw7U003_0;
	wire w_dff_A_ieo9pNzn8_0;
	wire w_dff_A_vrhsss888_0;
	wire w_dff_A_woTG74pO7_0;
	wire w_dff_A_72D0u0by4_0;
	wire w_dff_A_PLOyHNKq5_0;
	wire w_dff_A_29S28ue60_0;
	wire w_dff_A_keZsIW5T0_0;
	wire w_dff_A_Q8l7aJsV0_0;
	wire w_dff_A_OhTY83Rd8_0;
	wire w_dff_A_kM3AliSJ6_0;
	wire w_dff_A_86whUlow5_0;
	wire w_dff_A_8UlC83LO4_0;
	wire w_dff_A_iKGDNwfx3_0;
	wire w_dff_A_hN7dwSJE8_0;
	wire w_dff_A_TnokJ5nQ7_0;
	wire w_dff_A_m86Z4tSp8_0;
	wire w_dff_A_02Bq87UL8_0;
	wire w_dff_A_WUnYuut38_0;
	wire w_dff_A_cBWohS1Z9_0;
	wire w_dff_A_5sxAXsZZ2_0;
	wire w_dff_A_NqQJ7Q9N7_0;
	wire w_dff_A_edrMVVhI0_0;
	wire w_dff_A_mc2ocRHi5_0;
	wire w_dff_A_ClIG4uEj0_0;
	wire w_dff_A_qTqooJ4g5_0;
	wire w_dff_A_okMi2w5I6_2;
	wire w_dff_A_mmqCAwQQ0_0;
	wire w_dff_A_jqnpxvNa9_0;
	wire w_dff_A_D4aIypSf1_0;
	wire w_dff_A_9F7A4NHn8_0;
	wire w_dff_A_vSOF2bZ24_0;
	wire w_dff_A_uNXe2iYU3_0;
	wire w_dff_A_lRk8e8la5_0;
	wire w_dff_A_cHwFbjZE0_0;
	wire w_dff_A_lgumkYTG3_0;
	wire w_dff_A_eb5JBGlA6_0;
	wire w_dff_A_oic7v7yG5_0;
	wire w_dff_A_FORKC9420_0;
	wire w_dff_A_gfUeqGK95_0;
	wire w_dff_A_Q7M2dmfq1_0;
	wire w_dff_A_hGO9D4ZK3_0;
	wire w_dff_A_eMN0Lyhf3_0;
	wire w_dff_A_IcRl3GVm5_0;
	wire w_dff_A_d4vweEuQ4_0;
	wire w_dff_A_fhHm3dOI4_0;
	wire w_dff_A_TjnycSFa1_0;
	wire w_dff_A_XenvYTYa7_0;
	wire w_dff_A_3hJ0cqb57_0;
	wire w_dff_A_qvypK3uu5_0;
	wire w_dff_A_TjEhGHcb0_0;
	wire w_dff_A_uQZ1sL6C8_0;
	wire w_dff_A_ShKNXAb48_0;
	wire w_dff_A_hT8zARTA3_0;
	wire w_dff_A_3iIVPtIy0_2;
	wire w_dff_A_TH0McGuv2_0;
	wire w_dff_A_1tBOBIB03_0;
	wire w_dff_A_Qeapd9vl1_0;
	wire w_dff_A_xWsUKLVc5_0;
	wire w_dff_A_EO82gKr26_0;
	wire w_dff_A_cGcdneVv0_0;
	wire w_dff_A_OXZH8Ev40_0;
	wire w_dff_A_ScY5LJbO9_0;
	wire w_dff_A_t9AJSCtL8_0;
	wire w_dff_A_8RJtbIcx6_0;
	wire w_dff_A_wkmvjhQv7_0;
	wire w_dff_A_MFUeYaer4_0;
	wire w_dff_A_2r97kzzL1_0;
	wire w_dff_A_SZPHObf33_0;
	wire w_dff_A_m7XT8p5y2_0;
	wire w_dff_A_Cqeo3oVs2_0;
	wire w_dff_A_yFybcONs6_0;
	wire w_dff_A_Cpf0AO8S8_0;
	wire w_dff_A_mIDikPEU3_0;
	wire w_dff_A_8CQWHjB58_0;
	wire w_dff_A_2kzLPTvc2_0;
	wire w_dff_A_CnQxLwoq5_0;
	wire w_dff_A_NM6yUNZu4_0;
	wire w_dff_A_QvzwaO3j7_0;
	wire w_dff_A_nESaPY9Y1_0;
	wire w_dff_A_UyaYymEo5_2;
	wire w_dff_A_CLR1cD3l5_0;
	wire w_dff_A_qbNEzUsY4_0;
	wire w_dff_A_7RC0Upu28_0;
	wire w_dff_A_LZyI69R21_0;
	wire w_dff_A_NpWq06f96_0;
	wire w_dff_A_jGs2LuPI6_0;
	wire w_dff_A_xvfqY82a2_0;
	wire w_dff_A_7wOeM5Yg7_0;
	wire w_dff_A_a4aepqnD1_0;
	wire w_dff_A_N30RBU3j1_0;
	wire w_dff_A_H0X0Wm9v6_0;
	wire w_dff_A_c5N44hHk3_0;
	wire w_dff_A_JkVAFg4G2_0;
	wire w_dff_A_T5wClN0H7_0;
	wire w_dff_A_SE7CBLWH4_0;
	wire w_dff_A_gS5j8tEI6_0;
	wire w_dff_A_oUED2Fr67_0;
	wire w_dff_A_sQEAefrg6_0;
	wire w_dff_A_j1s66bpE5_0;
	wire w_dff_A_qXI94FpI0_0;
	wire w_dff_A_K7faFUhy4_0;
	wire w_dff_A_72L7YKCR9_0;
	wire w_dff_A_3MmwWSic9_0;
	wire w_dff_A_nCWPNuLc1_0;
	wire w_dff_A_5lkC1ky40_2;
	wire w_dff_A_OISVg6qP5_0;
	wire w_dff_A_y9lT7fhQ5_0;
	wire w_dff_A_2oxaerVo3_0;
	wire w_dff_A_dk5s9Qxe5_0;
	wire w_dff_A_LEc3BTSR4_0;
	wire w_dff_A_1Jc7roqJ1_0;
	wire w_dff_A_3sKt7CUo6_0;
	wire w_dff_A_olkl87Jj3_0;
	wire w_dff_A_wsZ5ojC10_0;
	wire w_dff_A_Sb09y2jW7_0;
	wire w_dff_A_QtSPrnah2_0;
	wire w_dff_A_dV7twkBH2_0;
	wire w_dff_A_A4pMx8fq4_0;
	wire w_dff_A_hSmILgKU8_0;
	wire w_dff_A_HIv5fYST7_0;
	wire w_dff_A_zWlbSlYz7_0;
	wire w_dff_A_lInS9lwp3_0;
	wire w_dff_A_PKjcF8ZR7_0;
	wire w_dff_A_sezIkoQa5_0;
	wire w_dff_A_5hturpCd7_0;
	wire w_dff_A_HeJUNTxn5_0;
	wire w_dff_A_ZzX8KFrT7_0;
	wire w_dff_A_yzVOykgA5_2;
	wire w_dff_A_nYyHfqI36_0;
	wire w_dff_A_t3iTvneP3_0;
	wire w_dff_A_I70Es19W1_0;
	wire w_dff_A_V1TQ6Yxg8_0;
	wire w_dff_A_KJIJFdNi3_0;
	wire w_dff_A_ou10IiEt3_0;
	wire w_dff_A_EuHGMMbj1_0;
	wire w_dff_A_dv9MIYmE0_0;
	wire w_dff_A_wU7Ypb4D1_0;
	wire w_dff_A_y3QdUFRR8_0;
	wire w_dff_A_uXi4uYz30_0;
	wire w_dff_A_nmauDiGY8_0;
	wire w_dff_A_nvlstr0F3_0;
	wire w_dff_A_uK05PgXN7_0;
	wire w_dff_A_2gUMQ6Ez8_0;
	wire w_dff_A_hz74bhKB2_0;
	wire w_dff_A_Fkys4IKG2_0;
	wire w_dff_A_oVAjaGor1_0;
	wire w_dff_A_mMZtzphy0_0;
	wire w_dff_A_upFUzfVE3_0;
	wire w_dff_A_CdP4FEpr4_2;
	wire w_dff_A_YmJQOPXe6_0;
	wire w_dff_A_dZ5hM3BL9_0;
	wire w_dff_A_zMy2P6rC1_0;
	wire w_dff_A_GThilhKC2_0;
	wire w_dff_A_ZlkLXRqS6_0;
	wire w_dff_A_0gGD8cSC0_0;
	wire w_dff_A_z6O5gkmr2_0;
	wire w_dff_A_KDyyAq3I6_0;
	wire w_dff_A_ENYoDgN90_0;
	wire w_dff_A_giftbn219_0;
	wire w_dff_A_pA2bGjJH7_0;
	wire w_dff_A_hwvQOeus6_0;
	wire w_dff_A_snNeLaxx7_0;
	wire w_dff_A_XRf37nWQ7_0;
	wire w_dff_A_oOspxazI5_0;
	wire w_dff_A_105n3lWY2_0;
	wire w_dff_A_l2BaYcZ29_0;
	wire w_dff_A_euOPKNzS4_0;
	wire w_dff_A_HN7yDTv85_2;
	wire w_dff_A_RpX5OA6x2_0;
	wire w_dff_A_jmf8UfBV6_0;
	wire w_dff_A_6ivIQwPA9_0;
	wire w_dff_A_JNkMfS620_0;
	wire w_dff_A_hkNq3aHH0_0;
	wire w_dff_A_kM1wyV0K5_0;
	wire w_dff_A_RyDYXRC51_0;
	wire w_dff_A_3GSiUFl94_0;
	wire w_dff_A_Qm70PGdU8_0;
	wire w_dff_A_EAGjHtSv9_0;
	wire w_dff_A_kD5VZRvd3_0;
	wire w_dff_A_HaGpOdSV0_0;
	wire w_dff_A_MSuQjyhW9_0;
	wire w_dff_A_QYdJGrRl3_0;
	wire w_dff_A_WU8237Lx4_0;
	wire w_dff_A_uQFiSjFw0_0;
	wire w_dff_A_5arqhEZw5_2;
	wire w_dff_A_9CKZi3AS6_0;
	wire w_dff_A_8al8690v7_0;
	wire w_dff_A_CL7wU4204_0;
	wire w_dff_A_Bi1nK5XC8_0;
	wire w_dff_A_9sFUi5mS4_0;
	wire w_dff_A_cfkZlF4D1_0;
	wire w_dff_A_vM5byLDi9_0;
	wire w_dff_A_f1KZGQfn5_0;
	wire w_dff_A_MaLPbrWR8_0;
	wire w_dff_A_EbVELEbw0_0;
	wire w_dff_A_5CXZnEeV2_0;
	wire w_dff_A_ZJxOxn1Z9_0;
	wire w_dff_A_cW4hY6gH8_0;
	wire w_dff_A_VtS6o35P7_0;
	wire w_dff_A_OWGNsutV7_2;
	wire w_dff_A_H03cf2lL9_0;
	wire w_dff_A_5lHIJwDH5_0;
	wire w_dff_A_j2EuERaM6_0;
	wire w_dff_A_CG92fvNm1_0;
	wire w_dff_A_P87da74r3_0;
	wire w_dff_A_XTmRmp8A1_0;
	wire w_dff_A_GgkbaN2K3_0;
	wire w_dff_A_DKlpFjiM6_0;
	wire w_dff_A_Cv8Wk0hu7_0;
	wire w_dff_A_uD06ZPIu0_0;
	wire w_dff_A_PM8G6V623_0;
	wire w_dff_A_ldmD4Pg34_0;
	wire w_dff_A_FgSjYYdM3_2;
	wire w_dff_A_tJmfc1aX8_0;
	wire w_dff_A_esA7WomA6_0;
	wire w_dff_A_bV8WZ6pc6_0;
	wire w_dff_A_Tyex67UV2_0;
	wire w_dff_A_tBkbXq5g4_0;
	wire w_dff_A_udNx3lHZ0_0;
	wire w_dff_A_4PmcjKeH8_0;
	wire w_dff_A_b1vuRf3a4_0;
	wire w_dff_A_dua3Bi0M8_0;
	wire w_dff_A_vcl3bDJl7_0;
	wire w_dff_A_c6Fm6OCo3_2;
	wire w_dff_A_x8t5Shk49_0;
	wire w_dff_A_wDfxn7zY6_0;
	wire w_dff_A_AjLI4VpR0_0;
	wire w_dff_A_r3sMAMPb3_0;
	wire w_dff_A_WR9E9Aag2_0;
	wire w_dff_A_kuq4Pi7Z7_0;
	wire w_dff_A_ytZxEyU76_0;
	wire w_dff_A_JW9f4wSa2_0;
	wire w_dff_A_cTXjgFSt7_2;
	wire w_dff_A_zgz3aUWA5_0;
	wire w_dff_A_AvJiQkvT6_0;
	wire w_dff_A_apui6QwY8_0;
	wire w_dff_A_QWaLqLGT0_0;
	wire w_dff_A_7HV5KXse8_0;
	wire w_dff_A_OnBH3vUl3_0;
	wire w_dff_A_MtaWg8ib7_2;
	wire w_dff_A_KzyXslny6_0;
	wire w_dff_A_wSRmAakt8_0;
	wire w_dff_A_ZVdSCnXX0_0;
	wire w_dff_A_j9NUrqag8_0;
	wire w_dff_A_GvGhDXPx3_2;
	wire w_dff_A_PAyX2J2a8_0;
	wire w_dff_A_N2tTzVE14_0;
	wire w_dff_A_l6uLDiYR0_2;
	jand g0000(.dina(w_G273gat_7[1]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G290gat_7[2]),.dinb(w_G18gat_7[1]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_n65_0[1]),.dinb(w_G545gat_0),.dout(n66),.clk(gclk));
	jnot g0003(.din(w_n66_0[1]),.dout(n67),.clk(gclk));
	jnot g0004(.din(w_G18gat_7[0]),.dout(n68),.clk(gclk));
	jnot g0005(.din(w_G273gat_7[0]),.dout(n69),.clk(gclk));
	jor g0006(.dina(w_n69_0[1]),.dinb(n68),.dout(n70),.clk(gclk));
	jnot g0007(.din(w_n70_0[1]),.dout(n71),.clk(gclk));
	jand g0008(.dina(w_G290gat_7[1]),.dinb(w_G1gat_7[0]),.dout(n72),.clk(gclk));
	jor g0009(.dina(w_dff_B_lEuxbv5F0_0),.dinb(n71),.dout(n73),.clk(gclk));
	jand g0010(.dina(n73),.dinb(w_n67_0[1]),.dout(w_dff_A_TXpAQk9U3_2),.clk(gclk));
	jand g0011(.dina(w_G307gat_7[1]),.dinb(w_G1gat_6[2]),.dout(n75),.clk(gclk));
	jnot g0012(.din(w_n75_0[1]),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G290gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jor g0016(.dina(n79),.dinb(w_n70_0[0]),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G273gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jor g0018(.dina(n81),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jand g0019(.dina(w_dff_B_QKLZD07U2_0),.dinb(w_n80_0[2]),.dout(n83),.clk(gclk));
	jxor g0020(.dina(w_n83_0[1]),.dinb(w_n67_0[0]),.dout(n84),.clk(gclk));
	jxor g0021(.dina(w_n84_0[1]),.dinb(w_dff_B_5LuDeCfj3_1),.dout(w_dff_A_buo4FdL10_2),.clk(gclk));
	jand g0022(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n86),.clk(gclk));
	jnot g0023(.din(w_n86_0[1]),.dout(n87),.clk(gclk));
	jor g0024(.dina(w_n83_0[0]),.dinb(w_n66_0[0]),.dout(n88),.clk(gclk));
	jor g0025(.dina(w_n84_0[0]),.dinb(w_n75_0[0]),.dout(n89),.clk(gclk));
	jand g0026(.dina(n89),.dinb(w_dff_B_bRNIW5P95_1),.dout(n90),.clk(gclk));
	jand g0027(.dina(w_G307gat_7[0]),.dinb(w_G18gat_6[2]),.dout(n91),.clk(gclk));
	jnot g0028(.din(w_n91_0[1]),.dout(n92),.clk(gclk));
	jnot g0029(.din(w_n80_0[1]),.dout(n93),.clk(gclk));
	jor g0030(.dina(w_n69_0[0]),.dinb(w_n77_0[0]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_G52gat_7[2]),.dout(n95),.clk(gclk));
	jor g0032(.dina(w_n78_0[0]),.dinb(n95),.dout(n96),.clk(gclk));
	jor g0033(.dina(n96),.dinb(n94),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G273gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jor g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jand g0037(.dina(w_dff_B_AsRBWcbj0_0),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g0038(.dina(w_n101_0[2]),.dinb(w_n93_0[1]),.dout(n102),.clk(gclk));
	jxor g0039(.dina(n102),.dinb(w_dff_B_cXBzVoJC3_1),.dout(n103),.clk(gclk));
	jxor g0040(.dina(w_n103_0[1]),.dinb(w_n90_0[1]),.dout(n104),.clk(gclk));
	jxor g0041(.dina(w_n104_0[1]),.dinb(w_dff_B_HfeP3lcw0_1),.dout(w_dff_A_dMBLpPmk9_2),.clk(gclk));
	jand g0042(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n106),.clk(gclk));
	jnot g0043(.din(w_n106_0[1]),.dout(n107),.clk(gclk));
	jnot g0044(.din(w_n103_0[0]),.dout(n108),.clk(gclk));
	jor g0045(.dina(n108),.dinb(w_n90_0[0]),.dout(n109),.clk(gclk));
	jor g0046(.dina(w_n104_0[0]),.dinb(w_n86_0[0]),.dout(n110),.clk(gclk));
	jand g0047(.dina(n110),.dinb(w_dff_B_wzAgij7Z4_1),.dout(n111),.clk(gclk));
	jand g0048(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n112),.clk(gclk));
	jnot g0049(.din(w_n112_0[1]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n101_0[1]),.dinb(w_n93_0[0]),.dout(n114),.clk(gclk));
	jxor g0051(.dina(w_n101_0[0]),.dinb(w_n80_0[0]),.dout(n115),.clk(gclk));
	jor g0052(.dina(n115),.dinb(w_n91_0[0]),.dout(n116),.clk(gclk));
	jand g0053(.dina(n116),.dinb(w_dff_B_lka824er8_1),.dout(n117),.clk(gclk));
	jand g0054(.dina(w_G307gat_6[2]),.dinb(w_G35gat_6[2]),.dout(n118),.clk(gclk));
	jnot g0055(.din(n118),.dout(n119),.clk(gclk));
	jnot g0056(.din(w_n97_0[0]),.dout(n120),.clk(gclk));
	jand g0057(.dina(w_G290gat_6[1]),.dinb(w_G69gat_7[1]),.dout(n121),.clk(gclk));
	jand g0058(.dina(w_n121_0[1]),.dinb(w_n99_0[0]),.dout(n122),.clk(gclk));
	jnot g0059(.din(w_n122_0[1]),.dout(n123),.clk(gclk));
	jand g0060(.dina(w_G290gat_6[0]),.dinb(w_G52gat_7[0]),.dout(n124),.clk(gclk));
	jand g0061(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n125),.clk(gclk));
	jor g0062(.dina(w_n125_0[1]),.dinb(n124),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_dff_B_dzB81Hgh7_0),.dinb(w_n123_0[1]),.dout(n127),.clk(gclk));
	jxor g0064(.dina(w_n127_0[1]),.dinb(w_n120_0[1]),.dout(n128),.clk(gclk));
	jxor g0065(.dina(w_n128_0[1]),.dinb(w_n119_0[1]),.dout(n129),.clk(gclk));
	jnot g0066(.din(w_n129_0[1]),.dout(n130),.clk(gclk));
	jxor g0067(.dina(w_n130_0[1]),.dinb(w_n117_0[2]),.dout(n131),.clk(gclk));
	jxor g0068(.dina(n131),.dinb(w_dff_B_Su360Bny1_1),.dout(n132),.clk(gclk));
	jxor g0069(.dina(w_n132_0[1]),.dinb(w_n111_0[1]),.dout(n133),.clk(gclk));
	jxor g0070(.dina(w_n133_0[1]),.dinb(w_dff_B_k71p4s1n3_1),.dout(w_dff_A_gefk1wav5_2),.clk(gclk));
	jand g0071(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n135),.clk(gclk));
	jnot g0072(.din(w_n135_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(w_n132_0[0]),.dout(n137),.clk(gclk));
	jor g0074(.dina(n137),.dinb(w_n111_0[0]),.dout(n138),.clk(gclk));
	jor g0075(.dina(w_n133_0[0]),.dinb(w_n106_0[0]),.dout(n139),.clk(gclk));
	jand g0076(.dina(n139),.dinb(w_dff_B_gf04LRoR5_1),.dout(n140),.clk(gclk));
	jand g0077(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n141),.clk(gclk));
	jnot g0078(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jor g0079(.dina(w_n130_0[0]),.dinb(w_n117_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n129_0[0]),.dinb(w_n117_0[0]),.dout(n144),.clk(gclk));
	jor g0081(.dina(n144),.dinb(w_n112_0[0]),.dout(n145),.clk(gclk));
	jand g0082(.dina(n145),.dinb(w_dff_B_BZ4iv02w0_1),.dout(n146),.clk(gclk));
	jand g0083(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n147),.clk(gclk));
	jnot g0084(.din(n147),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n127_0[0]),.dinb(w_n120_0[0]),.dout(n149),.clk(gclk));
	jnot g0086(.din(n149),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_n128_0[0]),.dinb(w_n119_0[0]),.dout(n151),.clk(gclk));
	jor g0088(.dina(n151),.dinb(n150),.dout(n152),.clk(gclk));
	jand g0089(.dina(w_G307gat_6[1]),.dinb(w_G52gat_6[2]),.dout(n153),.clk(gclk));
	jnot g0090(.din(n153),.dout(n154),.clk(gclk));
	jand g0091(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n155),.clk(gclk));
	jand g0092(.dina(w_n155_0[1]),.dinb(w_n125_0[0]),.dout(n156),.clk(gclk));
	jnot g0093(.din(w_n156_0[1]),.dout(n157),.clk(gclk));
	jand g0094(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n158),.clk(gclk));
	jor g0095(.dina(w_n158_0[1]),.dinb(w_n121_0[0]),.dout(n159),.clk(gclk));
	jand g0096(.dina(w_dff_B_p96wqOZf1_0),.dinb(w_n157_0[1]),.dout(n160),.clk(gclk));
	jxor g0097(.dina(w_n160_0[1]),.dinb(w_n122_0[0]),.dout(n161),.clk(gclk));
	jxor g0098(.dina(w_n161_0[1]),.dinb(w_n154_0[1]),.dout(n162),.clk(gclk));
	jxor g0099(.dina(w_n162_0[1]),.dinb(w_n152_0[1]),.dout(n163),.clk(gclk));
	jxor g0100(.dina(w_n163_0[1]),.dinb(w_n148_0[1]),.dout(n164),.clk(gclk));
	jnot g0101(.din(w_n164_0[1]),.dout(n165),.clk(gclk));
	jxor g0102(.dina(w_n165_0[1]),.dinb(w_n146_0[2]),.dout(n166),.clk(gclk));
	jxor g0103(.dina(n166),.dinb(w_dff_B_kHBgj2ct0_1),.dout(n167),.clk(gclk));
	jxor g0104(.dina(w_n167_0[1]),.dinb(w_n140_0[1]),.dout(n168),.clk(gclk));
	jxor g0105(.dina(w_n168_0[1]),.dinb(w_dff_B_PcDM2u6M1_1),.dout(w_dff_A_4JhpDJQk1_2),.clk(gclk));
	jand g0106(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n170),.clk(gclk));
	jnot g0107(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jnot g0108(.din(w_n167_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(n172),.dinb(w_n140_0[0]),.dout(n173),.clk(gclk));
	jor g0110(.dina(w_n168_0[0]),.dinb(w_n135_0[0]),.dout(n174),.clk(gclk));
	jand g0111(.dina(n174),.dinb(w_dff_B_mivY9yYO3_1),.dout(n175),.clk(gclk));
	jand g0112(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n176),.clk(gclk));
	jnot g0113(.din(w_n176_0[1]),.dout(n177),.clk(gclk));
	jor g0114(.dina(w_n165_0[0]),.dinb(w_n146_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n164_0[0]),.dinb(w_n146_0[0]),.dout(n179),.clk(gclk));
	jor g0116(.dina(n179),.dinb(w_n141_0[0]),.dout(n180),.clk(gclk));
	jand g0117(.dina(n180),.dinb(w_dff_B_HfKmuf415_1),.dout(n181),.clk(gclk));
	jand g0118(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n182),.clk(gclk));
	jnot g0119(.din(n182),.dout(n183),.clk(gclk));
	jand g0120(.dina(w_n162_0[0]),.dinb(w_n152_0[0]),.dout(n184),.clk(gclk));
	jand g0121(.dina(w_n163_0[0]),.dinb(w_n148_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(w_dff_B_APnmgULd0_1),.dout(n186),.clk(gclk));
	jand g0123(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n187),.clk(gclk));
	jnot g0124(.din(n187),.dout(n188),.clk(gclk));
	jnot g0125(.din(w_n160_0[0]),.dout(n189),.clk(gclk));
	jand g0126(.dina(n189),.dinb(w_n123_0[0]),.dout(n190),.clk(gclk));
	jand g0127(.dina(w_n161_0[0]),.dinb(w_n154_0[0]),.dout(n191),.clk(gclk));
	jor g0128(.dina(n191),.dinb(n190),.dout(n192),.clk(gclk));
	jand g0129(.dina(w_G307gat_6[0]),.dinb(w_G69gat_6[2]),.dout(n193),.clk(gclk));
	jnot g0130(.din(n193),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n195),.clk(gclk));
	jand g0132(.dina(w_n195_0[1]),.dinb(w_n158_0[0]),.dout(n196),.clk(gclk));
	jnot g0133(.din(w_n196_0[2]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(w_n198_0[1]),.dinb(w_n155_0[0]),.dout(n199),.clk(gclk));
	jand g0136(.dina(w_dff_B_Bo96JeWH4_0),.dinb(n197),.dout(n200),.clk(gclk));
	jxor g0137(.dina(w_n200_0[1]),.dinb(w_n156_0[0]),.dout(n201),.clk(gclk));
	jxor g0138(.dina(w_n201_0[1]),.dinb(w_n194_0[1]),.dout(n202),.clk(gclk));
	jxor g0139(.dina(w_n202_0[1]),.dinb(w_n192_0[1]),.dout(n203),.clk(gclk));
	jxor g0140(.dina(w_n203_0[1]),.dinb(w_n188_0[1]),.dout(n204),.clk(gclk));
	jxor g0141(.dina(w_n204_0[1]),.dinb(w_n186_0[1]),.dout(n205),.clk(gclk));
	jxor g0142(.dina(w_n205_0[1]),.dinb(w_n183_0[1]),.dout(n206),.clk(gclk));
	jnot g0143(.din(w_n206_0[1]),.dout(n207),.clk(gclk));
	jxor g0144(.dina(w_n207_0[1]),.dinb(w_n181_0[2]),.dout(n208),.clk(gclk));
	jxor g0145(.dina(n208),.dinb(w_dff_B_223yyBnc1_1),.dout(n209),.clk(gclk));
	jxor g0146(.dina(w_n209_0[1]),.dinb(w_n175_0[1]),.dout(n210),.clk(gclk));
	jxor g0147(.dina(w_n210_0[1]),.dinb(w_dff_B_5lzuWr6g6_1),.dout(w_dff_A_fzty24Fg7_2),.clk(gclk));
	jand g0148(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n212),.clk(gclk));
	jnot g0149(.din(w_n212_0[1]),.dout(n213),.clk(gclk));
	jnot g0150(.din(w_n209_0[0]),.dout(n214),.clk(gclk));
	jor g0151(.dina(n214),.dinb(w_n175_0[0]),.dout(n215),.clk(gclk));
	jor g0152(.dina(w_n210_0[0]),.dinb(w_n170_0[0]),.dout(n216),.clk(gclk));
	jand g0153(.dina(n216),.dinb(w_dff_B_e2lxoe595_1),.dout(n217),.clk(gclk));
	jand g0154(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n218),.clk(gclk));
	jnot g0155(.din(w_n218_0[1]),.dout(n219),.clk(gclk));
	jor g0156(.dina(w_n207_0[0]),.dinb(w_n181_0[1]),.dout(n220),.clk(gclk));
	jxor g0157(.dina(w_n206_0[0]),.dinb(w_n181_0[0]),.dout(n221),.clk(gclk));
	jor g0158(.dina(n221),.dinb(w_n176_0[0]),.dout(n222),.clk(gclk));
	jand g0159(.dina(n222),.dinb(w_dff_B_3vhxBByS6_1),.dout(n223),.clk(gclk));
	jand g0160(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n224),.clk(gclk));
	jnot g0161(.din(n224),.dout(n225),.clk(gclk));
	jand g0162(.dina(w_n204_0[0]),.dinb(w_n186_0[0]),.dout(n226),.clk(gclk));
	jand g0163(.dina(w_n205_0[0]),.dinb(w_n183_0[0]),.dout(n227),.clk(gclk));
	jor g0164(.dina(n227),.dinb(w_dff_B_wrVJX94M6_1),.dout(n228),.clk(gclk));
	jand g0165(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n229),.clk(gclk));
	jnot g0166(.din(n229),.dout(n230),.clk(gclk));
	jand g0167(.dina(w_n202_0[0]),.dinb(w_n192_0[0]),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_n203_0[0]),.dinb(w_n188_0[0]),.dout(n232),.clk(gclk));
	jor g0169(.dina(n232),.dinb(w_dff_B_FHDfKqcc2_1),.dout(n233),.clk(gclk));
	jand g0170(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n234),.clk(gclk));
	jnot g0171(.din(n234),.dout(n235),.clk(gclk));
	jnot g0172(.din(w_n200_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_n157_0[0]),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_n201_0[0]),.dinb(w_n194_0[0]),.dout(n238),.clk(gclk));
	jor g0175(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_G307gat_5[2]),.dinb(w_G86gat_6[2]),.dout(n240),.clk(gclk));
	jnot g0177(.din(n240),.dout(n241),.clk(gclk));
	jand g0178(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_n242_0[1]),.dinb(w_n198_0[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(w_n243_0[2]),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n245),.clk(gclk));
	jor g0182(.dina(w_n245_0[1]),.dinb(w_n195_0[0]),.dout(n246),.clk(gclk));
	jand g0183(.dina(w_dff_B_GV8eUhdT1_0),.dinb(n244),.dout(n247),.clk(gclk));
	jxor g0184(.dina(w_n247_0[1]),.dinb(w_n196_0[1]),.dout(n248),.clk(gclk));
	jxor g0185(.dina(w_n248_0[1]),.dinb(w_n241_0[1]),.dout(n249),.clk(gclk));
	jxor g0186(.dina(w_n249_0[1]),.dinb(w_n239_0[1]),.dout(n250),.clk(gclk));
	jxor g0187(.dina(w_n250_0[1]),.dinb(w_n235_0[1]),.dout(n251),.clk(gclk));
	jxor g0188(.dina(w_n251_0[1]),.dinb(w_n233_0[1]),.dout(n252),.clk(gclk));
	jxor g0189(.dina(w_n252_0[1]),.dinb(w_n230_0[1]),.dout(n253),.clk(gclk));
	jxor g0190(.dina(w_n253_0[1]),.dinb(w_n228_0[1]),.dout(n254),.clk(gclk));
	jxor g0191(.dina(w_n254_0[1]),.dinb(w_n225_0[1]),.dout(n255),.clk(gclk));
	jnot g0192(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jxor g0193(.dina(w_n256_0[1]),.dinb(w_n223_0[2]),.dout(n257),.clk(gclk));
	jxor g0194(.dina(n257),.dinb(w_dff_B_aBcORKe87_1),.dout(n258),.clk(gclk));
	jxor g0195(.dina(w_n258_0[1]),.dinb(w_n217_0[1]),.dout(n259),.clk(gclk));
	jxor g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_so7U7eC87_1),.dout(w_dff_A_1S7EK9uC0_2),.clk(gclk));
	jand g0197(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n261),.clk(gclk));
	jnot g0198(.din(w_n261_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(w_n258_0[0]),.dout(n263),.clk(gclk));
	jor g0200(.dina(n263),.dinb(w_n217_0[0]),.dout(n264),.clk(gclk));
	jor g0201(.dina(w_n259_0[0]),.dinb(w_n212_0[0]),.dout(n265),.clk(gclk));
	jand g0202(.dina(n265),.dinb(w_dff_B_adsMT2n22_1),.dout(n266),.clk(gclk));
	jand g0203(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n267),.clk(gclk));
	jnot g0204(.din(w_n267_0[1]),.dout(n268),.clk(gclk));
	jor g0205(.dina(w_n256_0[0]),.dinb(w_n223_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n255_0[0]),.dinb(w_n223_0[0]),.dout(n270),.clk(gclk));
	jor g0207(.dina(n270),.dinb(w_n218_0[0]),.dout(n271),.clk(gclk));
	jand g0208(.dina(n271),.dinb(w_dff_B_r4hNDjzn8_1),.dout(n272),.clk(gclk));
	jand g0209(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n273),.clk(gclk));
	jnot g0210(.din(n273),.dout(n274),.clk(gclk));
	jand g0211(.dina(w_n253_0[0]),.dinb(w_n228_0[0]),.dout(n275),.clk(gclk));
	jand g0212(.dina(w_n254_0[0]),.dinb(w_n225_0[0]),.dout(n276),.clk(gclk));
	jor g0213(.dina(n276),.dinb(w_dff_B_genMed2k6_1),.dout(n277),.clk(gclk));
	jand g0214(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n278),.clk(gclk));
	jnot g0215(.din(n278),.dout(n279),.clk(gclk));
	jand g0216(.dina(w_n251_0[0]),.dinb(w_n233_0[0]),.dout(n280),.clk(gclk));
	jand g0217(.dina(w_n252_0[0]),.dinb(w_n230_0[0]),.dout(n281),.clk(gclk));
	jor g0218(.dina(n281),.dinb(w_dff_B_Y4Mwki8N8_1),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(n283),.dout(n284),.clk(gclk));
	jand g0221(.dina(w_n249_0[0]),.dinb(w_n239_0[0]),.dout(n285),.clk(gclk));
	jand g0222(.dina(w_n250_0[0]),.dinb(w_n235_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(w_dff_B_bwQLdsF85_1),.dout(n287),.clk(gclk));
	jand g0224(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n288),.clk(gclk));
	jnot g0225(.din(n288),.dout(n289),.clk(gclk));
	jor g0226(.dina(w_n247_0[0]),.dinb(w_n196_0[0]),.dout(n290),.clk(gclk));
	jnot g0227(.din(n290),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n248_0[0]),.dinb(w_n241_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(n291),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G307gat_5[1]),.dinb(w_G103gat_6[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n296_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g0234(.din(w_n297_0[2]),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n299),.clk(gclk));
	jor g0236(.dina(w_n299_0[1]),.dinb(w_n242_0[0]),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_dff_B_z4cPPlU19_0),.dinb(n298),.dout(n301),.clk(gclk));
	jxor g0238(.dina(w_n301_0[1]),.dinb(w_n243_0[1]),.dout(n302),.clk(gclk));
	jxor g0239(.dina(w_n302_0[1]),.dinb(w_n295_0[1]),.dout(n303),.clk(gclk));
	jxor g0240(.dina(w_n303_0[1]),.dinb(w_n293_0[1]),.dout(n304),.clk(gclk));
	jxor g0241(.dina(w_n304_0[1]),.dinb(w_n289_0[1]),.dout(n305),.clk(gclk));
	jxor g0242(.dina(w_n305_0[1]),.dinb(w_n287_0[1]),.dout(n306),.clk(gclk));
	jxor g0243(.dina(w_n306_0[1]),.dinb(w_n284_0[1]),.dout(n307),.clk(gclk));
	jxor g0244(.dina(w_n307_0[1]),.dinb(w_n282_0[1]),.dout(n308),.clk(gclk));
	jxor g0245(.dina(w_n308_0[1]),.dinb(w_n279_0[1]),.dout(n309),.clk(gclk));
	jxor g0246(.dina(w_n309_0[1]),.dinb(w_n277_0[1]),.dout(n310),.clk(gclk));
	jxor g0247(.dina(w_n310_0[1]),.dinb(w_n274_0[1]),.dout(n311),.clk(gclk));
	jnot g0248(.din(w_n311_0[1]),.dout(n312),.clk(gclk));
	jxor g0249(.dina(w_n312_0[1]),.dinb(w_n272_0[2]),.dout(n313),.clk(gclk));
	jxor g0250(.dina(n313),.dinb(w_dff_B_vzXoSk9X4_1),.dout(n314),.clk(gclk));
	jxor g0251(.dina(w_n314_0[1]),.dinb(w_n266_0[1]),.dout(n315),.clk(gclk));
	jxor g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_m3PEL1Gm3_1),.dout(w_dff_A_fdK3GZD42_2),.clk(gclk));
	jand g0253(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n317),.clk(gclk));
	jnot g0254(.din(w_n317_0[1]),.dout(n318),.clk(gclk));
	jnot g0255(.din(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g0256(.dina(n319),.dinb(w_n266_0[0]),.dout(n320),.clk(gclk));
	jor g0257(.dina(w_n315_0[0]),.dinb(w_n261_0[0]),.dout(n321),.clk(gclk));
	jand g0258(.dina(n321),.dinb(w_dff_B_P7NpbNA11_1),.dout(n322),.clk(gclk));
	jand g0259(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n323),.clk(gclk));
	jnot g0260(.din(w_n323_0[1]),.dout(n324),.clk(gclk));
	jor g0261(.dina(w_n312_0[0]),.dinb(w_n272_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n311_0[0]),.dinb(w_n272_0[0]),.dout(n326),.clk(gclk));
	jor g0263(.dina(n326),.dinb(w_n267_0[0]),.dout(n327),.clk(gclk));
	jand g0264(.dina(n327),.dinb(w_dff_B_qxEaHlTH9_1),.dout(n328),.clk(gclk));
	jand g0265(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n329),.clk(gclk));
	jnot g0266(.din(n329),.dout(n330),.clk(gclk));
	jand g0267(.dina(w_n309_0[0]),.dinb(w_n277_0[0]),.dout(n331),.clk(gclk));
	jand g0268(.dina(w_n310_0[0]),.dinb(w_n274_0[0]),.dout(n332),.clk(gclk));
	jor g0269(.dina(n332),.dinb(w_dff_B_TLyREf666_1),.dout(n333),.clk(gclk));
	jand g0270(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n334),.clk(gclk));
	jnot g0271(.din(n334),.dout(n335),.clk(gclk));
	jand g0272(.dina(w_n307_0[0]),.dinb(w_n282_0[0]),.dout(n336),.clk(gclk));
	jand g0273(.dina(w_n308_0[0]),.dinb(w_n279_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(w_dff_B_npBmo3FI2_1),.dout(n338),.clk(gclk));
	jand g0275(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n339),.clk(gclk));
	jnot g0276(.din(n339),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_n305_0[0]),.dinb(w_n287_0[0]),.dout(n341),.clk(gclk));
	jand g0278(.dina(w_n306_0[0]),.dinb(w_n284_0[0]),.dout(n342),.clk(gclk));
	jor g0279(.dina(n342),.dinb(w_dff_B_7jaHZNBo7_1),.dout(n343),.clk(gclk));
	jand g0280(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n344),.clk(gclk));
	jnot g0281(.din(n344),.dout(n345),.clk(gclk));
	jand g0282(.dina(w_n303_0[0]),.dinb(w_n293_0[0]),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_n304_0[0]),.dinb(w_n289_0[0]),.dout(n347),.clk(gclk));
	jor g0284(.dina(n347),.dinb(w_dff_B_vTLeOGiF5_1),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n349),.clk(gclk));
	jnot g0286(.din(n349),.dout(n350),.clk(gclk));
	jor g0287(.dina(w_n301_0[0]),.dinb(w_n243_0[0]),.dout(n351),.clk(gclk));
	jnot g0288(.din(n351),.dout(n352),.clk(gclk));
	jand g0289(.dina(w_n302_0[0]),.dinb(w_n295_0[0]),.dout(n353),.clk(gclk));
	jor g0290(.dina(n353),.dinb(n352),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_G307gat_5[0]),.dinb(w_G120gat_6[2]),.dout(n355),.clk(gclk));
	jnot g0292(.din(n355),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n357),.clk(gclk));
	jand g0294(.dina(w_n357_0[1]),.dinb(w_n299_0[0]),.dout(n358),.clk(gclk));
	jnot g0295(.din(w_n358_0[2]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(w_n360_0[1]),.dinb(w_n296_0[0]),.dout(n361),.clk(gclk));
	jand g0298(.dina(w_dff_B_wHOweIil2_0),.dinb(n359),.dout(n362),.clk(gclk));
	jxor g0299(.dina(w_n362_0[1]),.dinb(w_n297_0[1]),.dout(n363),.clk(gclk));
	jxor g0300(.dina(w_n363_0[1]),.dinb(w_n356_0[1]),.dout(n364),.clk(gclk));
	jxor g0301(.dina(w_n364_0[1]),.dinb(w_n354_0[1]),.dout(n365),.clk(gclk));
	jxor g0302(.dina(w_n365_0[1]),.dinb(w_n350_0[1]),.dout(n366),.clk(gclk));
	jxor g0303(.dina(w_n366_0[1]),.dinb(w_n348_0[1]),.dout(n367),.clk(gclk));
	jxor g0304(.dina(w_n367_0[1]),.dinb(w_n345_0[1]),.dout(n368),.clk(gclk));
	jxor g0305(.dina(w_n368_0[1]),.dinb(w_n343_0[1]),.dout(n369),.clk(gclk));
	jxor g0306(.dina(w_n369_0[1]),.dinb(w_n340_0[1]),.dout(n370),.clk(gclk));
	jxor g0307(.dina(w_n370_0[1]),.dinb(w_n338_0[1]),.dout(n371),.clk(gclk));
	jxor g0308(.dina(w_n371_0[1]),.dinb(w_n335_0[1]),.dout(n372),.clk(gclk));
	jxor g0309(.dina(w_n372_0[1]),.dinb(w_n333_0[1]),.dout(n373),.clk(gclk));
	jxor g0310(.dina(w_n373_0[1]),.dinb(w_n330_0[1]),.dout(n374),.clk(gclk));
	jnot g0311(.din(w_n374_0[1]),.dout(n375),.clk(gclk));
	jxor g0312(.dina(w_n375_0[1]),.dinb(w_n328_0[2]),.dout(n376),.clk(gclk));
	jxor g0313(.dina(n376),.dinb(w_dff_B_Y7eTPMcT7_1),.dout(n377),.clk(gclk));
	jxor g0314(.dina(w_n377_0[1]),.dinb(w_n322_0[1]),.dout(n378),.clk(gclk));
	jxor g0315(.dina(w_n378_0[1]),.dinb(w_dff_B_vGQOMZBB4_1),.dout(w_dff_A_rFD3ruyP8_2),.clk(gclk));
	jand g0316(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n380),.clk(gclk));
	jnot g0317(.din(w_n380_0[1]),.dout(n381),.clk(gclk));
	jnot g0318(.din(w_n377_0[0]),.dout(n382),.clk(gclk));
	jor g0319(.dina(n382),.dinb(w_n322_0[0]),.dout(n383),.clk(gclk));
	jor g0320(.dina(w_n378_0[0]),.dinb(w_n317_0[0]),.dout(n384),.clk(gclk));
	jand g0321(.dina(n384),.dinb(w_dff_B_qUFUEihJ6_1),.dout(n385),.clk(gclk));
	jand g0322(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n386),.clk(gclk));
	jnot g0323(.din(w_n386_0[1]),.dout(n387),.clk(gclk));
	jor g0324(.dina(w_n375_0[0]),.dinb(w_n328_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n374_0[0]),.dinb(w_n328_0[0]),.dout(n389),.clk(gclk));
	jor g0326(.dina(n389),.dinb(w_n323_0[0]),.dout(n390),.clk(gclk));
	jand g0327(.dina(n390),.dinb(w_dff_B_XzZDx8md5_1),.dout(n391),.clk(gclk));
	jand g0328(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n392),.clk(gclk));
	jnot g0329(.din(n392),.dout(n393),.clk(gclk));
	jand g0330(.dina(w_n372_0[0]),.dinb(w_n333_0[0]),.dout(n394),.clk(gclk));
	jand g0331(.dina(w_n373_0[0]),.dinb(w_n330_0[0]),.dout(n395),.clk(gclk));
	jor g0332(.dina(n395),.dinb(w_dff_B_ZPrv69rY1_1),.dout(n396),.clk(gclk));
	jand g0333(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n397),.clk(gclk));
	jnot g0334(.din(n397),.dout(n398),.clk(gclk));
	jand g0335(.dina(w_n370_0[0]),.dinb(w_n338_0[0]),.dout(n399),.clk(gclk));
	jand g0336(.dina(w_n371_0[0]),.dinb(w_n335_0[0]),.dout(n400),.clk(gclk));
	jor g0337(.dina(n400),.dinb(w_dff_B_8KXdKmmc6_1),.dout(n401),.clk(gclk));
	jand g0338(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n402),.clk(gclk));
	jnot g0339(.din(n402),.dout(n403),.clk(gclk));
	jand g0340(.dina(w_n368_0[0]),.dinb(w_n343_0[0]),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_n369_0[0]),.dinb(w_n340_0[0]),.dout(n405),.clk(gclk));
	jor g0342(.dina(n405),.dinb(w_dff_B_SU23IKnx1_1),.dout(n406),.clk(gclk));
	jand g0343(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n407),.clk(gclk));
	jnot g0344(.din(n407),.dout(n408),.clk(gclk));
	jand g0345(.dina(w_n366_0[0]),.dinb(w_n348_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(w_n367_0[0]),.dinb(w_n345_0[0]),.dout(n410),.clk(gclk));
	jor g0347(.dina(n410),.dinb(w_dff_B_NBaNDCuu2_1),.dout(n411),.clk(gclk));
	jand g0348(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n412),.clk(gclk));
	jnot g0349(.din(n412),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n364_0[0]),.dinb(w_n354_0[0]),.dout(n414),.clk(gclk));
	jand g0351(.dina(w_n365_0[0]),.dinb(w_n350_0[0]),.dout(n415),.clk(gclk));
	jor g0352(.dina(n415),.dinb(w_dff_B_thuy0MMT4_1),.dout(n416),.clk(gclk));
	jand g0353(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n417),.clk(gclk));
	jnot g0354(.din(n417),.dout(n418),.clk(gclk));
	jor g0355(.dina(w_n362_0[0]),.dinb(w_n297_0[0]),.dout(n419),.clk(gclk));
	jand g0356(.dina(w_n363_0[0]),.dinb(w_n356_0[0]),.dout(n420),.clk(gclk));
	jnot g0357(.din(n420),.dout(n421),.clk(gclk));
	jand g0358(.dina(n421),.dinb(w_dff_B_LhXZKNt04_1),.dout(n422),.clk(gclk));
	jnot g0359(.din(n422),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_G307gat_4[2]),.dinb(w_G137gat_6[2]),.dout(n424),.clk(gclk));
	jnot g0361(.din(n424),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n426),.clk(gclk));
	jand g0363(.dina(w_n426_0[1]),.dinb(w_n360_0[0]),.dout(n427),.clk(gclk));
	jnot g0364(.din(w_n427_0[2]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(w_n429_0[1]),.dinb(w_n357_0[0]),.dout(n430),.clk(gclk));
	jand g0367(.dina(w_dff_B_tFhInTpS8_0),.dinb(n428),.dout(n431),.clk(gclk));
	jxor g0368(.dina(w_n431_0[1]),.dinb(w_n358_0[1]),.dout(n432),.clk(gclk));
	jxor g0369(.dina(w_n432_0[1]),.dinb(w_n425_0[1]),.dout(n433),.clk(gclk));
	jxor g0370(.dina(w_n433_0[1]),.dinb(w_n423_0[1]),.dout(n434),.clk(gclk));
	jxor g0371(.dina(w_n434_0[1]),.dinb(w_n418_0[1]),.dout(n435),.clk(gclk));
	jxor g0372(.dina(w_n435_0[1]),.dinb(w_n416_0[1]),.dout(n436),.clk(gclk));
	jxor g0373(.dina(w_n436_0[1]),.dinb(w_n413_0[1]),.dout(n437),.clk(gclk));
	jxor g0374(.dina(w_n437_0[1]),.dinb(w_n411_0[1]),.dout(n438),.clk(gclk));
	jxor g0375(.dina(w_n438_0[1]),.dinb(w_n408_0[1]),.dout(n439),.clk(gclk));
	jxor g0376(.dina(w_n439_0[1]),.dinb(w_n406_0[1]),.dout(n440),.clk(gclk));
	jxor g0377(.dina(w_n440_0[1]),.dinb(w_n403_0[1]),.dout(n441),.clk(gclk));
	jxor g0378(.dina(w_n441_0[1]),.dinb(w_n401_0[1]),.dout(n442),.clk(gclk));
	jxor g0379(.dina(w_n442_0[1]),.dinb(w_n398_0[1]),.dout(n443),.clk(gclk));
	jxor g0380(.dina(w_n443_0[1]),.dinb(w_n396_0[1]),.dout(n444),.clk(gclk));
	jxor g0381(.dina(w_n444_0[1]),.dinb(w_n393_0[1]),.dout(n445),.clk(gclk));
	jnot g0382(.din(w_n445_0[1]),.dout(n446),.clk(gclk));
	jxor g0383(.dina(w_n446_0[1]),.dinb(w_n391_0[2]),.dout(n447),.clk(gclk));
	jxor g0384(.dina(n447),.dinb(w_dff_B_o39bPTKi1_1),.dout(n448),.clk(gclk));
	jxor g0385(.dina(w_n448_0[1]),.dinb(w_n385_0[1]),.dout(n449),.clk(gclk));
	jxor g0386(.dina(w_n449_0[1]),.dinb(w_dff_B_0X766xLg1_1),.dout(w_dff_A_xANsDdVz6_2),.clk(gclk));
	jand g0387(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n451),.clk(gclk));
	jnot g0388(.din(w_n451_0[1]),.dout(n452),.clk(gclk));
	jnot g0389(.din(w_n448_0[0]),.dout(n453),.clk(gclk));
	jor g0390(.dina(n453),.dinb(w_n385_0[0]),.dout(n454),.clk(gclk));
	jor g0391(.dina(w_n449_0[0]),.dinb(w_n380_0[0]),.dout(n455),.clk(gclk));
	jand g0392(.dina(n455),.dinb(w_dff_B_LJWEIvt20_1),.dout(n456),.clk(gclk));
	jand g0393(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n457),.clk(gclk));
	jnot g0394(.din(w_n457_0[1]),.dout(n458),.clk(gclk));
	jor g0395(.dina(w_n446_0[0]),.dinb(w_n391_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n445_0[0]),.dinb(w_n391_0[0]),.dout(n460),.clk(gclk));
	jor g0397(.dina(n460),.dinb(w_n386_0[0]),.dout(n461),.clk(gclk));
	jand g0398(.dina(n461),.dinb(w_dff_B_n8ulN2hL2_1),.dout(n462),.clk(gclk));
	jand g0399(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n463),.clk(gclk));
	jnot g0400(.din(n463),.dout(n464),.clk(gclk));
	jand g0401(.dina(w_n443_0[0]),.dinb(w_n396_0[0]),.dout(n465),.clk(gclk));
	jand g0402(.dina(w_n444_0[0]),.dinb(w_n393_0[0]),.dout(n466),.clk(gclk));
	jor g0403(.dina(n466),.dinb(w_dff_B_Jh6lq4521_1),.dout(n467),.clk(gclk));
	jand g0404(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n468),.clk(gclk));
	jnot g0405(.din(n468),.dout(n469),.clk(gclk));
	jand g0406(.dina(w_n441_0[0]),.dinb(w_n401_0[0]),.dout(n470),.clk(gclk));
	jand g0407(.dina(w_n442_0[0]),.dinb(w_n398_0[0]),.dout(n471),.clk(gclk));
	jor g0408(.dina(n471),.dinb(w_dff_B_dbiXsX4n4_1),.dout(n472),.clk(gclk));
	jand g0409(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n473),.clk(gclk));
	jnot g0410(.din(n473),.dout(n474),.clk(gclk));
	jand g0411(.dina(w_n439_0[0]),.dinb(w_n406_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(w_n440_0[0]),.dinb(w_n403_0[0]),.dout(n476),.clk(gclk));
	jor g0413(.dina(n476),.dinb(w_dff_B_OJBqW99N0_1),.dout(n477),.clk(gclk));
	jand g0414(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n478),.clk(gclk));
	jnot g0415(.din(n478),.dout(n479),.clk(gclk));
	jand g0416(.dina(w_n437_0[0]),.dinb(w_n411_0[0]),.dout(n480),.clk(gclk));
	jand g0417(.dina(w_n438_0[0]),.dinb(w_n408_0[0]),.dout(n481),.clk(gclk));
	jor g0418(.dina(n481),.dinb(w_dff_B_AwApN28D3_1),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n435_0[0]),.dinb(w_n416_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n436_0[0]),.dinb(w_n413_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(w_dff_B_w72PYw6U1_1),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n433_0[0]),.dinb(w_n423_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n434_0[0]),.dinb(w_n418_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(w_dff_B_TG7ggu479_1),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jor g0431(.dina(w_n431_0[0]),.dinb(w_n358_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n432_0[0]),.dinb(w_n425_0[0]),.dout(n496),.clk(gclk));
	jnot g0433(.din(n496),.dout(n497),.clk(gclk));
	jand g0434(.dina(n497),.dinb(w_dff_B_UTv53eIV5_1),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_G307gat_4[1]),.dinb(w_G154gat_6[2]),.dout(n500),.clk(gclk));
	jnot g0437(.din(n500),.dout(n501),.clk(gclk));
	jand g0438(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_n502_0[1]),.dinb(w_n429_0[0]),.dout(n503),.clk(gclk));
	jnot g0440(.din(w_n503_0[2]),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n505),.clk(gclk));
	jor g0442(.dina(w_n505_0[1]),.dinb(w_n426_0[0]),.dout(n506),.clk(gclk));
	jand g0443(.dina(w_dff_B_pZTOoJE89_0),.dinb(n504),.dout(n507),.clk(gclk));
	jxor g0444(.dina(w_n507_0[1]),.dinb(w_n427_0[1]),.dout(n508),.clk(gclk));
	jxor g0445(.dina(w_n508_0[1]),.dinb(w_n501_0[1]),.dout(n509),.clk(gclk));
	jxor g0446(.dina(w_n509_0[1]),.dinb(w_n499_0[1]),.dout(n510),.clk(gclk));
	jxor g0447(.dina(w_n510_0[1]),.dinb(w_n494_0[1]),.dout(n511),.clk(gclk));
	jxor g0448(.dina(w_n511_0[1]),.dinb(w_n492_0[1]),.dout(n512),.clk(gclk));
	jxor g0449(.dina(w_n512_0[1]),.dinb(w_n489_0[1]),.dout(n513),.clk(gclk));
	jxor g0450(.dina(w_n513_0[1]),.dinb(w_n487_0[1]),.dout(n514),.clk(gclk));
	jxor g0451(.dina(w_n514_0[1]),.dinb(w_n484_0[1]),.dout(n515),.clk(gclk));
	jxor g0452(.dina(w_n515_0[1]),.dinb(w_n482_0[1]),.dout(n516),.clk(gclk));
	jxor g0453(.dina(w_n516_0[1]),.dinb(w_n479_0[1]),.dout(n517),.clk(gclk));
	jxor g0454(.dina(w_n517_0[1]),.dinb(w_n477_0[1]),.dout(n518),.clk(gclk));
	jxor g0455(.dina(w_n518_0[1]),.dinb(w_n474_0[1]),.dout(n519),.clk(gclk));
	jxor g0456(.dina(w_n519_0[1]),.dinb(w_n472_0[1]),.dout(n520),.clk(gclk));
	jxor g0457(.dina(w_n520_0[1]),.dinb(w_n469_0[1]),.dout(n521),.clk(gclk));
	jxor g0458(.dina(w_n521_0[1]),.dinb(w_n467_0[1]),.dout(n522),.clk(gclk));
	jxor g0459(.dina(w_n522_0[1]),.dinb(w_n464_0[1]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[1]),.dout(n524),.clk(gclk));
	jxor g0461(.dina(w_n524_0[1]),.dinb(w_n462_0[2]),.dout(n525),.clk(gclk));
	jxor g0462(.dina(n525),.dinb(w_dff_B_YUvxqxm79_1),.dout(n526),.clk(gclk));
	jxor g0463(.dina(w_n526_0[1]),.dinb(w_n456_0[1]),.dout(n527),.clk(gclk));
	jxor g0464(.dina(w_n527_0[1]),.dinb(w_dff_B_1Aoe1Zp02_1),.dout(w_dff_A_k3iKXLIe4_2),.clk(gclk));
	jand g0465(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n529),.clk(gclk));
	jnot g0466(.din(w_n529_0[1]),.dout(n530),.clk(gclk));
	jnot g0467(.din(w_n526_0[0]),.dout(n531),.clk(gclk));
	jor g0468(.dina(n531),.dinb(w_n456_0[0]),.dout(n532),.clk(gclk));
	jor g0469(.dina(w_n527_0[0]),.dinb(w_n451_0[0]),.dout(n533),.clk(gclk));
	jand g0470(.dina(n533),.dinb(w_dff_B_VXK70yMo3_1),.dout(n534),.clk(gclk));
	jand g0471(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n535),.clk(gclk));
	jnot g0472(.din(w_n535_0[1]),.dout(n536),.clk(gclk));
	jor g0473(.dina(w_n524_0[0]),.dinb(w_n462_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n523_0[0]),.dinb(w_n462_0[0]),.dout(n538),.clk(gclk));
	jor g0475(.dina(n538),.dinb(w_n457_0[0]),.dout(n539),.clk(gclk));
	jand g0476(.dina(n539),.dinb(w_dff_B_25LyZmhv8_1),.dout(n540),.clk(gclk));
	jand g0477(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n541),.clk(gclk));
	jnot g0478(.din(n541),.dout(n542),.clk(gclk));
	jand g0479(.dina(w_n521_0[0]),.dinb(w_n467_0[0]),.dout(n543),.clk(gclk));
	jand g0480(.dina(w_n522_0[0]),.dinb(w_n464_0[0]),.dout(n544),.clk(gclk));
	jor g0481(.dina(n544),.dinb(w_dff_B_E0zn4wyP8_1),.dout(n545),.clk(gclk));
	jand g0482(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n546),.clk(gclk));
	jnot g0483(.din(n546),.dout(n547),.clk(gclk));
	jand g0484(.dina(w_n519_0[0]),.dinb(w_n472_0[0]),.dout(n548),.clk(gclk));
	jand g0485(.dina(w_n520_0[0]),.dinb(w_n469_0[0]),.dout(n549),.clk(gclk));
	jor g0486(.dina(n549),.dinb(w_dff_B_TF5vSIb98_1),.dout(n550),.clk(gclk));
	jand g0487(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n551),.clk(gclk));
	jnot g0488(.din(n551),.dout(n552),.clk(gclk));
	jand g0489(.dina(w_n517_0[0]),.dinb(w_n477_0[0]),.dout(n553),.clk(gclk));
	jand g0490(.dina(w_n518_0[0]),.dinb(w_n474_0[0]),.dout(n554),.clk(gclk));
	jor g0491(.dina(n554),.dinb(w_dff_B_5tQ7JrXv8_1),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n556),.clk(gclk));
	jnot g0493(.din(n556),.dout(n557),.clk(gclk));
	jand g0494(.dina(w_n515_0[0]),.dinb(w_n482_0[0]),.dout(n558),.clk(gclk));
	jand g0495(.dina(w_n516_0[0]),.dinb(w_n479_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(w_dff_B_yLerp6T52_1),.dout(n560),.clk(gclk));
	jand g0497(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n561),.clk(gclk));
	jnot g0498(.din(n561),.dout(n562),.clk(gclk));
	jand g0499(.dina(w_n513_0[0]),.dinb(w_n487_0[0]),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n514_0[0]),.dinb(w_n484_0[0]),.dout(n564),.clk(gclk));
	jor g0501(.dina(n564),.dinb(w_dff_B_sw5cd2Qe4_1),.dout(n565),.clk(gclk));
	jand g0502(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n566),.clk(gclk));
	jnot g0503(.din(n566),.dout(n567),.clk(gclk));
	jand g0504(.dina(w_n511_0[0]),.dinb(w_n492_0[0]),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n512_0[0]),.dinb(w_n489_0[0]),.dout(n569),.clk(gclk));
	jor g0506(.dina(n569),.dinb(w_dff_B_5W1HNHhA0_1),.dout(n570),.clk(gclk));
	jand g0507(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n571),.clk(gclk));
	jnot g0508(.din(n571),.dout(n572),.clk(gclk));
	jand g0509(.dina(w_n509_0[0]),.dinb(w_n499_0[0]),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n510_0[0]),.dinb(w_n494_0[0]),.dout(n574),.clk(gclk));
	jor g0511(.dina(n574),.dinb(w_dff_B_xDE2wZ4o5_1),.dout(n575),.clk(gclk));
	jand g0512(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n576),.clk(gclk));
	jnot g0513(.din(n576),.dout(n577),.clk(gclk));
	jor g0514(.dina(w_n507_0[0]),.dinb(w_n427_0[0]),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n508_0[0]),.dinb(w_n501_0[0]),.dout(n579),.clk(gclk));
	jnot g0516(.din(n579),.dout(n580),.clk(gclk));
	jand g0517(.dina(n580),.dinb(w_dff_B_Zdg8hQQA3_1),.dout(n581),.clk(gclk));
	jnot g0518(.din(n581),.dout(n582),.clk(gclk));
	jand g0519(.dina(w_G307gat_4[0]),.dinb(w_G171gat_6[2]),.dout(n583),.clk(gclk));
	jnot g0520(.din(n583),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n585),.clk(gclk));
	jand g0522(.dina(w_n585_0[1]),.dinb(w_n505_0[0]),.dout(n586),.clk(gclk));
	jnot g0523(.din(w_n586_0[2]),.dout(n587),.clk(gclk));
	jand g0524(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n588),.clk(gclk));
	jor g0525(.dina(w_n588_0[1]),.dinb(w_n502_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_dff_B_vPj7a03l5_0),.dinb(n587),.dout(n590),.clk(gclk));
	jxor g0527(.dina(w_n590_0[1]),.dinb(w_n503_0[1]),.dout(n591),.clk(gclk));
	jxor g0528(.dina(w_n591_0[1]),.dinb(w_n584_0[1]),.dout(n592),.clk(gclk));
	jxor g0529(.dina(w_n592_0[1]),.dinb(w_n582_0[1]),.dout(n593),.clk(gclk));
	jxor g0530(.dina(w_n593_0[1]),.dinb(w_n577_0[1]),.dout(n594),.clk(gclk));
	jxor g0531(.dina(w_n594_0[1]),.dinb(w_n575_0[1]),.dout(n595),.clk(gclk));
	jxor g0532(.dina(w_n595_0[1]),.dinb(w_n572_0[1]),.dout(n596),.clk(gclk));
	jxor g0533(.dina(w_n596_0[1]),.dinb(w_n570_0[1]),.dout(n597),.clk(gclk));
	jxor g0534(.dina(w_n597_0[1]),.dinb(w_n567_0[1]),.dout(n598),.clk(gclk));
	jxor g0535(.dina(w_n598_0[1]),.dinb(w_n565_0[1]),.dout(n599),.clk(gclk));
	jxor g0536(.dina(w_n599_0[1]),.dinb(w_n562_0[1]),.dout(n600),.clk(gclk));
	jxor g0537(.dina(w_n600_0[1]),.dinb(w_n560_0[1]),.dout(n601),.clk(gclk));
	jxor g0538(.dina(w_n601_0[1]),.dinb(w_n557_0[1]),.dout(n602),.clk(gclk));
	jxor g0539(.dina(w_n602_0[1]),.dinb(w_n555_0[1]),.dout(n603),.clk(gclk));
	jxor g0540(.dina(w_n603_0[1]),.dinb(w_n552_0[1]),.dout(n604),.clk(gclk));
	jxor g0541(.dina(w_n604_0[1]),.dinb(w_n550_0[1]),.dout(n605),.clk(gclk));
	jxor g0542(.dina(w_n605_0[1]),.dinb(w_n547_0[1]),.dout(n606),.clk(gclk));
	jxor g0543(.dina(w_n606_0[1]),.dinb(w_n545_0[1]),.dout(n607),.clk(gclk));
	jxor g0544(.dina(w_n607_0[1]),.dinb(w_n542_0[1]),.dout(n608),.clk(gclk));
	jnot g0545(.din(w_n608_0[1]),.dout(n609),.clk(gclk));
	jxor g0546(.dina(w_n609_0[1]),.dinb(w_n540_0[2]),.dout(n610),.clk(gclk));
	jxor g0547(.dina(n610),.dinb(w_dff_B_vR0plZ4L4_1),.dout(n611),.clk(gclk));
	jxor g0548(.dina(w_n611_0[1]),.dinb(w_n534_0[1]),.dout(n612),.clk(gclk));
	jxor g0549(.dina(w_n612_0[1]),.dinb(w_dff_B_EMXdE2Dp7_1),.dout(w_dff_A_Whz6y90z4_2),.clk(gclk));
	jand g0550(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n614),.clk(gclk));
	jnot g0551(.din(w_n614_0[1]),.dout(n615),.clk(gclk));
	jnot g0552(.din(w_n611_0[0]),.dout(n616),.clk(gclk));
	jor g0553(.dina(n616),.dinb(w_n534_0[0]),.dout(n617),.clk(gclk));
	jor g0554(.dina(w_n612_0[0]),.dinb(w_n529_0[0]),.dout(n618),.clk(gclk));
	jand g0555(.dina(n618),.dinb(w_dff_B_ZVITaAWb1_1),.dout(n619),.clk(gclk));
	jand g0556(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n620),.clk(gclk));
	jnot g0557(.din(w_n620_0[1]),.dout(n621),.clk(gclk));
	jor g0558(.dina(w_n609_0[0]),.dinb(w_n540_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n608_0[0]),.dinb(w_n540_0[0]),.dout(n623),.clk(gclk));
	jor g0560(.dina(n623),.dinb(w_n535_0[0]),.dout(n624),.clk(gclk));
	jand g0561(.dina(n624),.dinb(w_dff_B_L54OtKa01_1),.dout(n625),.clk(gclk));
	jand g0562(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n626),.clk(gclk));
	jnot g0563(.din(n626),.dout(n627),.clk(gclk));
	jand g0564(.dina(w_n606_0[0]),.dinb(w_n545_0[0]),.dout(n628),.clk(gclk));
	jand g0565(.dina(w_n607_0[0]),.dinb(w_n542_0[0]),.dout(n629),.clk(gclk));
	jor g0566(.dina(n629),.dinb(w_dff_B_AAk7rBFR0_1),.dout(n630),.clk(gclk));
	jand g0567(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n631),.clk(gclk));
	jnot g0568(.din(n631),.dout(n632),.clk(gclk));
	jand g0569(.dina(w_n604_0[0]),.dinb(w_n550_0[0]),.dout(n633),.clk(gclk));
	jand g0570(.dina(w_n605_0[0]),.dinb(w_n547_0[0]),.dout(n634),.clk(gclk));
	jor g0571(.dina(n634),.dinb(w_dff_B_pzUmcCNM8_1),.dout(n635),.clk(gclk));
	jand g0572(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n636),.clk(gclk));
	jnot g0573(.din(n636),.dout(n637),.clk(gclk));
	jand g0574(.dina(w_n602_0[0]),.dinb(w_n555_0[0]),.dout(n638),.clk(gclk));
	jand g0575(.dina(w_n603_0[0]),.dinb(w_n552_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(n639),.dinb(w_dff_B_zA1fVh209_1),.dout(n640),.clk(gclk));
	jand g0577(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n641),.clk(gclk));
	jnot g0578(.din(n641),.dout(n642),.clk(gclk));
	jand g0579(.dina(w_n600_0[0]),.dinb(w_n560_0[0]),.dout(n643),.clk(gclk));
	jand g0580(.dina(w_n601_0[0]),.dinb(w_n557_0[0]),.dout(n644),.clk(gclk));
	jor g0581(.dina(n644),.dinb(w_dff_B_tzp9z56e2_1),.dout(n645),.clk(gclk));
	jand g0582(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n646),.clk(gclk));
	jnot g0583(.din(n646),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_n598_0[0]),.dinb(w_n565_0[0]),.dout(n648),.clk(gclk));
	jand g0585(.dina(w_n599_0[0]),.dinb(w_n562_0[0]),.dout(n649),.clk(gclk));
	jor g0586(.dina(n649),.dinb(w_dff_B_C3gKgd3D9_1),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n651),.clk(gclk));
	jnot g0588(.din(n651),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_n596_0[0]),.dinb(w_n570_0[0]),.dout(n653),.clk(gclk));
	jand g0590(.dina(w_n597_0[0]),.dinb(w_n567_0[0]),.dout(n654),.clk(gclk));
	jor g0591(.dina(n654),.dinb(w_dff_B_3HGlLHHK0_1),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n656),.clk(gclk));
	jnot g0593(.din(n656),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_n594_0[0]),.dinb(w_n575_0[0]),.dout(n658),.clk(gclk));
	jand g0595(.dina(w_n595_0[0]),.dinb(w_n572_0[0]),.dout(n659),.clk(gclk));
	jor g0596(.dina(n659),.dinb(w_dff_B_2TtZjgDR4_1),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n661),.clk(gclk));
	jnot g0598(.din(n661),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_n592_0[0]),.dinb(w_n582_0[0]),.dout(n663),.clk(gclk));
	jand g0600(.dina(w_n593_0[0]),.dinb(w_n577_0[0]),.dout(n664),.clk(gclk));
	jor g0601(.dina(n664),.dinb(w_dff_B_fhsB5pI32_1),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n666),.clk(gclk));
	jnot g0603(.din(n666),.dout(n667),.clk(gclk));
	jor g0604(.dina(w_n590_0[0]),.dinb(w_n503_0[0]),.dout(n668),.clk(gclk));
	jand g0605(.dina(w_n591_0[0]),.dinb(w_n584_0[0]),.dout(n669),.clk(gclk));
	jnot g0606(.din(n669),.dout(n670),.clk(gclk));
	jand g0607(.dina(n670),.dinb(w_dff_B_Q8Jhx20V3_1),.dout(n671),.clk(gclk));
	jnot g0608(.din(n671),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G307gat_3[2]),.dinb(w_G188gat_6[2]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n675_0[1]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jnot g0613(.din(w_n676_0[2]),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n678),.clk(gclk));
	jor g0615(.dina(w_n678_0[1]),.dinb(w_n585_0[0]),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_dff_B_P53qelmo0_0),.dinb(n677),.dout(n680),.clk(gclk));
	jxor g0617(.dina(w_n680_0[1]),.dinb(w_n586_0[1]),.dout(n681),.clk(gclk));
	jxor g0618(.dina(w_n681_0[1]),.dinb(w_n674_0[1]),.dout(n682),.clk(gclk));
	jxor g0619(.dina(w_n682_0[1]),.dinb(w_n672_0[1]),.dout(n683),.clk(gclk));
	jxor g0620(.dina(w_n683_0[1]),.dinb(w_n667_0[1]),.dout(n684),.clk(gclk));
	jxor g0621(.dina(w_n684_0[1]),.dinb(w_n665_0[1]),.dout(n685),.clk(gclk));
	jxor g0622(.dina(w_n685_0[1]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jxor g0623(.dina(w_n686_0[1]),.dinb(w_n660_0[1]),.dout(n687),.clk(gclk));
	jxor g0624(.dina(w_n687_0[1]),.dinb(w_n657_0[1]),.dout(n688),.clk(gclk));
	jxor g0625(.dina(w_n688_0[1]),.dinb(w_n655_0[1]),.dout(n689),.clk(gclk));
	jxor g0626(.dina(w_n689_0[1]),.dinb(w_n652_0[1]),.dout(n690),.clk(gclk));
	jxor g0627(.dina(w_n690_0[1]),.dinb(w_n650_0[1]),.dout(n691),.clk(gclk));
	jxor g0628(.dina(w_n691_0[1]),.dinb(w_n647_0[1]),.dout(n692),.clk(gclk));
	jxor g0629(.dina(w_n692_0[1]),.dinb(w_n645_0[1]),.dout(n693),.clk(gclk));
	jxor g0630(.dina(w_n693_0[1]),.dinb(w_n642_0[1]),.dout(n694),.clk(gclk));
	jxor g0631(.dina(w_n694_0[1]),.dinb(w_n640_0[1]),.dout(n695),.clk(gclk));
	jxor g0632(.dina(w_n695_0[1]),.dinb(w_n637_0[1]),.dout(n696),.clk(gclk));
	jxor g0633(.dina(w_n696_0[1]),.dinb(w_n635_0[1]),.dout(n697),.clk(gclk));
	jxor g0634(.dina(w_n697_0[1]),.dinb(w_n632_0[1]),.dout(n698),.clk(gclk));
	jxor g0635(.dina(w_n698_0[1]),.dinb(w_n630_0[1]),.dout(n699),.clk(gclk));
	jxor g0636(.dina(w_n699_0[1]),.dinb(w_n627_0[1]),.dout(n700),.clk(gclk));
	jnot g0637(.din(w_n700_0[1]),.dout(n701),.clk(gclk));
	jxor g0638(.dina(w_n701_0[1]),.dinb(w_n625_0[2]),.dout(n702),.clk(gclk));
	jxor g0639(.dina(n702),.dinb(w_dff_B_0W0p7jUR3_1),.dout(n703),.clk(gclk));
	jxor g0640(.dina(w_n703_0[1]),.dinb(w_n619_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_dff_B_g0rjQRyU7_1),.dout(w_dff_A_dSuBmHpc5_2),.clk(gclk));
	jand g0642(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n706),.clk(gclk));
	jnot g0643(.din(w_n706_0[1]),.dout(n707),.clk(gclk));
	jnot g0644(.din(w_n703_0[0]),.dout(n708),.clk(gclk));
	jor g0645(.dina(n708),.dinb(w_n619_0[0]),.dout(n709),.clk(gclk));
	jor g0646(.dina(w_n704_0[0]),.dinb(w_n614_0[0]),.dout(n710),.clk(gclk));
	jand g0647(.dina(n710),.dinb(w_dff_B_fCo7Mjhw4_1),.dout(n711),.clk(gclk));
	jand g0648(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n712),.clk(gclk));
	jnot g0649(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jor g0650(.dina(w_n701_0[0]),.dinb(w_n625_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n700_0[0]),.dinb(w_n625_0[0]),.dout(n715),.clk(gclk));
	jor g0652(.dina(n715),.dinb(w_n620_0[0]),.dout(n716),.clk(gclk));
	jand g0653(.dina(n716),.dinb(w_dff_B_BOjcivN93_1),.dout(n717),.clk(gclk));
	jand g0654(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n718),.clk(gclk));
	jnot g0655(.din(n718),.dout(n719),.clk(gclk));
	jand g0656(.dina(w_n698_0[0]),.dinb(w_n630_0[0]),.dout(n720),.clk(gclk));
	jand g0657(.dina(w_n699_0[0]),.dinb(w_n627_0[0]),.dout(n721),.clk(gclk));
	jor g0658(.dina(n721),.dinb(w_dff_B_HgCApr8i9_1),.dout(n722),.clk(gclk));
	jand g0659(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n723),.clk(gclk));
	jnot g0660(.din(n723),.dout(n724),.clk(gclk));
	jand g0661(.dina(w_n696_0[0]),.dinb(w_n635_0[0]),.dout(n725),.clk(gclk));
	jand g0662(.dina(w_n697_0[0]),.dinb(w_n632_0[0]),.dout(n726),.clk(gclk));
	jor g0663(.dina(n726),.dinb(w_dff_B_72vJHDRm4_1),.dout(n727),.clk(gclk));
	jand g0664(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n728),.clk(gclk));
	jnot g0665(.din(n728),.dout(n729),.clk(gclk));
	jand g0666(.dina(w_n694_0[0]),.dinb(w_n640_0[0]),.dout(n730),.clk(gclk));
	jand g0667(.dina(w_n695_0[0]),.dinb(w_n637_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(w_dff_B_xlYWbEmV9_1),.dout(n732),.clk(gclk));
	jand g0669(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n733),.clk(gclk));
	jnot g0670(.din(n733),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_n692_0[0]),.dinb(w_n645_0[0]),.dout(n735),.clk(gclk));
	jand g0672(.dina(w_n693_0[0]),.dinb(w_n642_0[0]),.dout(n736),.clk(gclk));
	jor g0673(.dina(n736),.dinb(w_dff_B_y8GhzqHs6_1),.dout(n737),.clk(gclk));
	jand g0674(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n738),.clk(gclk));
	jnot g0675(.din(n738),.dout(n739),.clk(gclk));
	jand g0676(.dina(w_n690_0[0]),.dinb(w_n650_0[0]),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_n691_0[0]),.dinb(w_n647_0[0]),.dout(n741),.clk(gclk));
	jor g0678(.dina(n741),.dinb(w_dff_B_fmHAL9ae8_1),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n743),.clk(gclk));
	jnot g0680(.din(n743),.dout(n744),.clk(gclk));
	jand g0681(.dina(w_n688_0[0]),.dinb(w_n655_0[0]),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_n689_0[0]),.dinb(w_n652_0[0]),.dout(n746),.clk(gclk));
	jor g0683(.dina(n746),.dinb(w_dff_B_Y00TVUep1_1),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n748),.clk(gclk));
	jnot g0685(.din(n748),.dout(n749),.clk(gclk));
	jand g0686(.dina(w_n686_0[0]),.dinb(w_n660_0[0]),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_n687_0[0]),.dinb(w_n657_0[0]),.dout(n751),.clk(gclk));
	jor g0688(.dina(n751),.dinb(w_dff_B_yZ1ZLZMX3_1),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n753),.clk(gclk));
	jnot g0690(.din(n753),.dout(n754),.clk(gclk));
	jand g0691(.dina(w_n684_0[0]),.dinb(w_n665_0[0]),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_n685_0[0]),.dinb(w_n662_0[0]),.dout(n756),.clk(gclk));
	jor g0693(.dina(n756),.dinb(w_dff_B_L9dAiNeY6_1),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n758),.clk(gclk));
	jnot g0695(.din(n758),.dout(n759),.clk(gclk));
	jand g0696(.dina(w_n682_0[0]),.dinb(w_n672_0[0]),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_n683_0[0]),.dinb(w_n667_0[0]),.dout(n761),.clk(gclk));
	jor g0698(.dina(n761),.dinb(w_dff_B_MeaEWRaU7_1),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n763),.clk(gclk));
	jnot g0700(.din(n763),.dout(n764),.clk(gclk));
	jor g0701(.dina(w_n680_0[0]),.dinb(w_n586_0[0]),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_n681_0[0]),.dinb(w_n674_0[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(n767),.dinb(w_dff_B_6JvFeimc6_1),.dout(n768),.clk(gclk));
	jnot g0705(.din(n768),.dout(n769),.clk(gclk));
	jand g0706(.dina(w_G307gat_3[1]),.dinb(w_G205gat_6[2]),.dout(n770),.clk(gclk));
	jnot g0707(.din(n770),.dout(n771),.clk(gclk));
	jand g0708(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n772_0[1]),.dinb(w_n678_0[0]),.dout(n773),.clk(gclk));
	jnot g0710(.din(w_n773_0[1]),.dout(n774),.clk(gclk));
	jand g0711(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n775),.clk(gclk));
	jor g0712(.dina(w_n775_0[1]),.dinb(w_n675_0[0]),.dout(n776),.clk(gclk));
	jand g0713(.dina(w_dff_B_A0THsbh72_0),.dinb(w_n774_0[1]),.dout(n777),.clk(gclk));
	jxor g0714(.dina(w_n777_0[1]),.dinb(w_n676_0[1]),.dout(n778),.clk(gclk));
	jxor g0715(.dina(w_n778_0[1]),.dinb(w_n771_0[1]),.dout(n779),.clk(gclk));
	jxor g0716(.dina(w_n779_0[1]),.dinb(w_n769_0[1]),.dout(n780),.clk(gclk));
	jxor g0717(.dina(w_n780_0[1]),.dinb(w_n764_0[1]),.dout(n781),.clk(gclk));
	jxor g0718(.dina(w_n781_0[1]),.dinb(w_n762_0[1]),.dout(n782),.clk(gclk));
	jxor g0719(.dina(w_n782_0[1]),.dinb(w_n759_0[1]),.dout(n783),.clk(gclk));
	jxor g0720(.dina(w_n783_0[1]),.dinb(w_n757_0[1]),.dout(n784),.clk(gclk));
	jxor g0721(.dina(w_n784_0[1]),.dinb(w_n754_0[1]),.dout(n785),.clk(gclk));
	jxor g0722(.dina(w_n785_0[1]),.dinb(w_n752_0[1]),.dout(n786),.clk(gclk));
	jxor g0723(.dina(w_n786_0[1]),.dinb(w_n749_0[1]),.dout(n787),.clk(gclk));
	jxor g0724(.dina(w_n787_0[1]),.dinb(w_n747_0[1]),.dout(n788),.clk(gclk));
	jxor g0725(.dina(w_n788_0[1]),.dinb(w_n744_0[1]),.dout(n789),.clk(gclk));
	jxor g0726(.dina(w_n789_0[1]),.dinb(w_n742_0[1]),.dout(n790),.clk(gclk));
	jxor g0727(.dina(w_n790_0[1]),.dinb(w_n739_0[1]),.dout(n791),.clk(gclk));
	jxor g0728(.dina(w_n791_0[1]),.dinb(w_n737_0[1]),.dout(n792),.clk(gclk));
	jxor g0729(.dina(w_n792_0[1]),.dinb(w_n734_0[1]),.dout(n793),.clk(gclk));
	jxor g0730(.dina(w_n793_0[1]),.dinb(w_n732_0[1]),.dout(n794),.clk(gclk));
	jxor g0731(.dina(w_n794_0[1]),.dinb(w_n729_0[1]),.dout(n795),.clk(gclk));
	jxor g0732(.dina(w_n795_0[1]),.dinb(w_n727_0[1]),.dout(n796),.clk(gclk));
	jxor g0733(.dina(w_n796_0[1]),.dinb(w_n724_0[1]),.dout(n797),.clk(gclk));
	jxor g0734(.dina(w_n797_0[1]),.dinb(w_n722_0[1]),.dout(n798),.clk(gclk));
	jxor g0735(.dina(w_n798_0[1]),.dinb(w_n719_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(w_n799_0[1]),.dout(n800),.clk(gclk));
	jxor g0737(.dina(w_n800_0[1]),.dinb(w_n717_0[2]),.dout(n801),.clk(gclk));
	jxor g0738(.dina(n801),.dinb(w_dff_B_BYWga9r30_1),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n711_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_dff_B_R5ONn5iw7_1),.dout(w_dff_A_GrvPvRzD1_2),.clk(gclk));
	jand g0741(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n805),.clk(gclk));
	jnot g0742(.din(w_n805_0[1]),.dout(n806),.clk(gclk));
	jnot g0743(.din(w_n802_0[0]),.dout(n807),.clk(gclk));
	jor g0744(.dina(n807),.dinb(w_n711_0[0]),.dout(n808),.clk(gclk));
	jor g0745(.dina(w_n803_0[0]),.dinb(w_n706_0[0]),.dout(n809),.clk(gclk));
	jand g0746(.dina(n809),.dinb(w_dff_B_fUgsaO6R2_1),.dout(n810),.clk(gclk));
	jand g0747(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n811),.clk(gclk));
	jor g0748(.dina(w_n800_0[0]),.dinb(w_n717_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n799_0[0]),.dinb(w_n717_0[0]),.dout(n813),.clk(gclk));
	jor g0750(.dina(n813),.dinb(w_n712_0[0]),.dout(n814),.clk(gclk));
	jand g0751(.dina(n814),.dinb(w_dff_B_Z8LzQloI7_1),.dout(n815),.clk(gclk));
	jand g0752(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n816),.clk(gclk));
	jnot g0753(.din(w_n816_0[1]),.dout(n817),.clk(gclk));
	jand g0754(.dina(w_n797_0[0]),.dinb(w_n722_0[0]),.dout(n818),.clk(gclk));
	jand g0755(.dina(w_n798_0[0]),.dinb(w_n719_0[0]),.dout(n819),.clk(gclk));
	jor g0756(.dina(n819),.dinb(w_dff_B_S4ORdUCC3_1),.dout(n820),.clk(gclk));
	jand g0757(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n821),.clk(gclk));
	jnot g0758(.din(n821),.dout(n822),.clk(gclk));
	jand g0759(.dina(w_n795_0[0]),.dinb(w_n727_0[0]),.dout(n823),.clk(gclk));
	jand g0760(.dina(w_n796_0[0]),.dinb(w_n724_0[0]),.dout(n824),.clk(gclk));
	jor g0761(.dina(n824),.dinb(w_dff_B_ga3xMME42_1),.dout(n825),.clk(gclk));
	jand g0762(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n826),.clk(gclk));
	jnot g0763(.din(n826),.dout(n827),.clk(gclk));
	jand g0764(.dina(w_n793_0[0]),.dinb(w_n732_0[0]),.dout(n828),.clk(gclk));
	jand g0765(.dina(w_n794_0[0]),.dinb(w_n729_0[0]),.dout(n829),.clk(gclk));
	jor g0766(.dina(n829),.dinb(w_dff_B_njc17Ywt8_1),.dout(n830),.clk(gclk));
	jand g0767(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n831),.clk(gclk));
	jnot g0768(.din(n831),.dout(n832),.clk(gclk));
	jand g0769(.dina(w_n791_0[0]),.dinb(w_n737_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(w_n792_0[0]),.dinb(w_n734_0[0]),.dout(n834),.clk(gclk));
	jor g0771(.dina(n834),.dinb(w_dff_B_R0z19Jep3_1),.dout(n835),.clk(gclk));
	jand g0772(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n836),.clk(gclk));
	jnot g0773(.din(n836),.dout(n837),.clk(gclk));
	jand g0774(.dina(w_n789_0[0]),.dinb(w_n742_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(w_n790_0[0]),.dinb(w_n739_0[0]),.dout(n839),.clk(gclk));
	jor g0776(.dina(n839),.dinb(w_dff_B_AojH413d8_1),.dout(n840),.clk(gclk));
	jand g0777(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n841),.clk(gclk));
	jnot g0778(.din(n841),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n787_0[0]),.dinb(w_n747_0[0]),.dout(n843),.clk(gclk));
	jand g0780(.dina(w_n788_0[0]),.dinb(w_n744_0[0]),.dout(n844),.clk(gclk));
	jor g0781(.dina(n844),.dinb(w_dff_B_yT5jobxk4_1),.dout(n845),.clk(gclk));
	jand g0782(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n846),.clk(gclk));
	jnot g0783(.din(n846),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n785_0[0]),.dinb(w_n752_0[0]),.dout(n848),.clk(gclk));
	jand g0785(.dina(w_n786_0[0]),.dinb(w_n749_0[0]),.dout(n849),.clk(gclk));
	jor g0786(.dina(n849),.dinb(w_dff_B_ze7CwRxD5_1),.dout(n850),.clk(gclk));
	jand g0787(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n851),.clk(gclk));
	jnot g0788(.din(n851),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n783_0[0]),.dinb(w_n757_0[0]),.dout(n853),.clk(gclk));
	jand g0790(.dina(w_n784_0[0]),.dinb(w_n754_0[0]),.dout(n854),.clk(gclk));
	jor g0791(.dina(n854),.dinb(w_dff_B_0SQLVANx9_1),.dout(n855),.clk(gclk));
	jand g0792(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n856),.clk(gclk));
	jnot g0793(.din(n856),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n781_0[0]),.dinb(w_n762_0[0]),.dout(n858),.clk(gclk));
	jand g0795(.dina(w_n782_0[0]),.dinb(w_n759_0[0]),.dout(n859),.clk(gclk));
	jor g0796(.dina(n859),.dinb(w_dff_B_ls7eEVDF7_1),.dout(n860),.clk(gclk));
	jand g0797(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n861),.clk(gclk));
	jnot g0798(.din(n861),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n779_0[0]),.dinb(w_n769_0[0]),.dout(n863),.clk(gclk));
	jand g0800(.dina(w_n780_0[0]),.dinb(w_n764_0[0]),.dout(n864),.clk(gclk));
	jor g0801(.dina(n864),.dinb(w_dff_B_rX2M1cWh8_1),.dout(n865),.clk(gclk));
	jand g0802(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n866),.clk(gclk));
	jnot g0803(.din(n866),.dout(n867),.clk(gclk));
	jor g0804(.dina(w_n777_0[0]),.dinb(w_n676_0[0]),.dout(n868),.clk(gclk));
	jand g0805(.dina(w_n778_0[0]),.dinb(w_n771_0[0]),.dout(n869),.clk(gclk));
	jnot g0806(.din(n869),.dout(n870),.clk(gclk));
	jand g0807(.dina(n870),.dinb(w_dff_B_IPyqcC861_1),.dout(n871),.clk(gclk));
	jnot g0808(.din(n871),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_G307gat_3[0]),.dinb(w_G222gat_6[2]),.dout(n873),.clk(gclk));
	jnot g0810(.din(n873),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n875),.clk(gclk));
	jxor g0812(.dina(w_n875_0[1]),.dinb(w_n772_0[0]),.dout(n876),.clk(gclk));
	jor g0813(.dina(n876),.dinb(w_n773_0[0]),.dout(n877),.clk(gclk));
	jor g0814(.dina(w_n875_0[0]),.dinb(w_n774_0[0]),.dout(n878),.clk(gclk));
	jand g0815(.dina(n878),.dinb(w_n877_0[1]),.dout(n879),.clk(gclk));
	jxor g0816(.dina(w_n879_0[1]),.dinb(w_n874_0[1]),.dout(n880),.clk(gclk));
	jxor g0817(.dina(w_n880_0[1]),.dinb(w_n872_0[1]),.dout(n881),.clk(gclk));
	jxor g0818(.dina(w_n881_0[1]),.dinb(w_n867_0[1]),.dout(n882),.clk(gclk));
	jxor g0819(.dina(w_n882_0[1]),.dinb(w_n865_0[1]),.dout(n883),.clk(gclk));
	jxor g0820(.dina(w_n883_0[1]),.dinb(w_n862_0[1]),.dout(n884),.clk(gclk));
	jxor g0821(.dina(w_n884_0[1]),.dinb(w_n860_0[1]),.dout(n885),.clk(gclk));
	jxor g0822(.dina(w_n885_0[1]),.dinb(w_n857_0[1]),.dout(n886),.clk(gclk));
	jxor g0823(.dina(w_n886_0[1]),.dinb(w_n855_0[1]),.dout(n887),.clk(gclk));
	jxor g0824(.dina(w_n887_0[1]),.dinb(w_n852_0[1]),.dout(n888),.clk(gclk));
	jxor g0825(.dina(w_n888_0[1]),.dinb(w_n850_0[1]),.dout(n889),.clk(gclk));
	jxor g0826(.dina(w_n889_0[1]),.dinb(w_n847_0[1]),.dout(n890),.clk(gclk));
	jxor g0827(.dina(w_n890_0[1]),.dinb(w_n845_0[1]),.dout(n891),.clk(gclk));
	jxor g0828(.dina(w_n891_0[1]),.dinb(w_n842_0[1]),.dout(n892),.clk(gclk));
	jxor g0829(.dina(w_n892_0[1]),.dinb(w_n840_0[1]),.dout(n893),.clk(gclk));
	jxor g0830(.dina(w_n893_0[1]),.dinb(w_n837_0[1]),.dout(n894),.clk(gclk));
	jxor g0831(.dina(w_n894_0[1]),.dinb(w_n835_0[1]),.dout(n895),.clk(gclk));
	jxor g0832(.dina(w_n895_0[1]),.dinb(w_n832_0[1]),.dout(n896),.clk(gclk));
	jxor g0833(.dina(w_n896_0[1]),.dinb(w_n830_0[1]),.dout(n897),.clk(gclk));
	jxor g0834(.dina(w_n897_0[1]),.dinb(w_n827_0[1]),.dout(n898),.clk(gclk));
	jxor g0835(.dina(w_n898_0[1]),.dinb(w_n825_0[1]),.dout(n899),.clk(gclk));
	jxor g0836(.dina(w_n899_0[1]),.dinb(w_n822_0[1]),.dout(n900),.clk(gclk));
	jxor g0837(.dina(w_n900_0[2]),.dinb(w_n820_0[2]),.dout(n901),.clk(gclk));
	jxor g0838(.dina(n901),.dinb(w_dff_B_i87Plare9_1),.dout(n902),.clk(gclk));
	jxor g0839(.dina(w_n902_0[1]),.dinb(w_n815_0[1]),.dout(n903),.clk(gclk));
	jxor g0840(.dina(w_n903_0[1]),.dinb(w_n811_0[1]),.dout(n904),.clk(gclk));
	jxor g0841(.dina(w_n904_0[1]),.dinb(w_n810_0[1]),.dout(n905),.clk(gclk));
	jxor g0842(.dina(w_n905_0[1]),.dinb(w_dff_B_6y3Mt8UG5_1),.dout(w_dff_A_b9xSmEOi6_2),.clk(gclk));
	jnot g0843(.din(w_n904_0[0]),.dout(n907),.clk(gclk));
	jor g0844(.dina(n907),.dinb(w_n810_0[0]),.dout(n908),.clk(gclk));
	jor g0845(.dina(w_n905_0[0]),.dinb(w_n805_0[0]),.dout(n909),.clk(gclk));
	jand g0846(.dina(n909),.dinb(w_dff_B_4xi7J29C7_1),.dout(n910),.clk(gclk));
	jand g0847(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n911),.clk(gclk));
	jnot g0848(.din(w_n902_0[0]),.dout(n912),.clk(gclk));
	jor g0849(.dina(n912),.dinb(w_n815_0[0]),.dout(n913),.clk(gclk));
	jor g0850(.dina(w_n903_0[0]),.dinb(w_n811_0[0]),.dout(n914),.clk(gclk));
	jand g0851(.dina(n914),.dinb(w_dff_B_dHhXXkpS5_1),.dout(n915),.clk(gclk));
	jand g0852(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n916),.clk(gclk));
	jand g0853(.dina(w_n900_0[1]),.dinb(w_n820_0[1]),.dout(n917),.clk(gclk));
	jnot g0854(.din(n917),.dout(n918),.clk(gclk));
	jnot g0855(.din(w_n900_0[0]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(n919),.dinb(w_n820_0[0]),.dout(n920),.clk(gclk));
	jor g0857(.dina(n920),.dinb(w_n816_0[0]),.dout(n921),.clk(gclk));
	jand g0858(.dina(n921),.dinb(n918),.dout(n922),.clk(gclk));
	jand g0859(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n923),.clk(gclk));
	jnot g0860(.din(n923),.dout(n924),.clk(gclk));
	jand g0861(.dina(w_n898_0[0]),.dinb(w_n825_0[0]),.dout(n925),.clk(gclk));
	jand g0862(.dina(w_n899_0[0]),.dinb(w_n822_0[0]),.dout(n926),.clk(gclk));
	jor g0863(.dina(n926),.dinb(w_dff_B_kcbxlRjy9_1),.dout(n927),.clk(gclk));
	jand g0864(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n928),.clk(gclk));
	jnot g0865(.din(n928),.dout(n929),.clk(gclk));
	jand g0866(.dina(w_n896_0[0]),.dinb(w_n830_0[0]),.dout(n930),.clk(gclk));
	jand g0867(.dina(w_n897_0[0]),.dinb(w_n827_0[0]),.dout(n931),.clk(gclk));
	jor g0868(.dina(n931),.dinb(w_dff_B_btAzBAx92_1),.dout(n932),.clk(gclk));
	jand g0869(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n933),.clk(gclk));
	jnot g0870(.din(n933),.dout(n934),.clk(gclk));
	jand g0871(.dina(w_n894_0[0]),.dinb(w_n835_0[0]),.dout(n935),.clk(gclk));
	jand g0872(.dina(w_n895_0[0]),.dinb(w_n832_0[0]),.dout(n936),.clk(gclk));
	jor g0873(.dina(n936),.dinb(w_dff_B_3pE5dkfD9_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n938),.clk(gclk));
	jnot g0875(.din(n938),.dout(n939),.clk(gclk));
	jand g0876(.dina(w_n892_0[0]),.dinb(w_n840_0[0]),.dout(n940),.clk(gclk));
	jand g0877(.dina(w_n893_0[0]),.dinb(w_n837_0[0]),.dout(n941),.clk(gclk));
	jor g0878(.dina(n941),.dinb(w_dff_B_70voapNf1_1),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n943),.clk(gclk));
	jnot g0880(.din(n943),.dout(n944),.clk(gclk));
	jand g0881(.dina(w_n890_0[0]),.dinb(w_n845_0[0]),.dout(n945),.clk(gclk));
	jand g0882(.dina(w_n891_0[0]),.dinb(w_n842_0[0]),.dout(n946),.clk(gclk));
	jor g0883(.dina(n946),.dinb(w_dff_B_PDENw4BN8_1),.dout(n947),.clk(gclk));
	jand g0884(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n948),.clk(gclk));
	jnot g0885(.din(n948),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_n888_0[0]),.dinb(w_n850_0[0]),.dout(n950),.clk(gclk));
	jand g0887(.dina(w_n889_0[0]),.dinb(w_n847_0[0]),.dout(n951),.clk(gclk));
	jor g0888(.dina(n951),.dinb(w_dff_B_0oMYSq0L6_1),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n953),.clk(gclk));
	jnot g0890(.din(n953),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_n886_0[0]),.dinb(w_n855_0[0]),.dout(n955),.clk(gclk));
	jand g0892(.dina(w_n887_0[0]),.dinb(w_n852_0[0]),.dout(n956),.clk(gclk));
	jor g0893(.dina(n956),.dinb(w_dff_B_UxsF3NTc2_1),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n958),.clk(gclk));
	jnot g0895(.din(n958),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_n884_0[0]),.dinb(w_n860_0[0]),.dout(n960),.clk(gclk));
	jand g0897(.dina(w_n885_0[0]),.dinb(w_n857_0[0]),.dout(n961),.clk(gclk));
	jor g0898(.dina(n961),.dinb(w_dff_B_8eTRNjEg9_1),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n963),.clk(gclk));
	jnot g0900(.din(n963),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_n882_0[0]),.dinb(w_n865_0[0]),.dout(n965),.clk(gclk));
	jand g0902(.dina(w_n883_0[0]),.dinb(w_n862_0[0]),.dout(n966),.clk(gclk));
	jor g0903(.dina(n966),.dinb(w_dff_B_dvYDu3121_1),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n968),.clk(gclk));
	jnot g0905(.din(n968),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_n880_0[0]),.dinb(w_n872_0[0]),.dout(n970),.clk(gclk));
	jand g0907(.dina(w_n881_0[0]),.dinb(w_n867_0[0]),.dout(n971),.clk(gclk));
	jor g0908(.dina(n971),.dinb(w_dff_B_4oC1homs9_1),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n973),.clk(gclk));
	jnot g0910(.din(n973),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_n879_0[0]),.dinb(w_n874_0[0]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(n976),.dinb(w_n877_0[0]),.dout(n977),.clk(gclk));
	jnot g0914(.din(n977),.dout(n978),.clk(gclk));
	jnot g0915(.din(w_n775_0[0]),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n980),.clk(gclk));
	jand g0917(.dina(w_n980_0[1]),.dinb(n979),.dout(n981),.clk(gclk));
	jnot g0918(.din(n981),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_G307gat_2[2]),.dinb(w_G239gat_6[2]),.dout(n983),.clk(gclk));
	jxor g0920(.dina(w_n983_0[1]),.dinb(w_n982_0[1]),.dout(n984),.clk(gclk));
	jxor g0921(.dina(w_n984_0[1]),.dinb(w_n978_0[1]),.dout(n985),.clk(gclk));
	jxor g0922(.dina(w_n985_0[1]),.dinb(w_n974_0[1]),.dout(n986),.clk(gclk));
	jxor g0923(.dina(w_n986_0[1]),.dinb(w_n972_0[1]),.dout(n987),.clk(gclk));
	jxor g0924(.dina(w_n987_0[1]),.dinb(w_n969_0[1]),.dout(n988),.clk(gclk));
	jxor g0925(.dina(w_n988_0[1]),.dinb(w_n967_0[1]),.dout(n989),.clk(gclk));
	jxor g0926(.dina(w_n989_0[1]),.dinb(w_n964_0[1]),.dout(n990),.clk(gclk));
	jxor g0927(.dina(w_n990_0[1]),.dinb(w_n962_0[1]),.dout(n991),.clk(gclk));
	jxor g0928(.dina(w_n991_0[1]),.dinb(w_n959_0[1]),.dout(n992),.clk(gclk));
	jxor g0929(.dina(w_n992_0[1]),.dinb(w_n957_0[1]),.dout(n993),.clk(gclk));
	jxor g0930(.dina(w_n993_0[1]),.dinb(w_n954_0[1]),.dout(n994),.clk(gclk));
	jxor g0931(.dina(w_n994_0[1]),.dinb(w_n952_0[1]),.dout(n995),.clk(gclk));
	jxor g0932(.dina(w_n995_0[1]),.dinb(w_n949_0[1]),.dout(n996),.clk(gclk));
	jxor g0933(.dina(w_n996_0[1]),.dinb(w_n947_0[1]),.dout(n997),.clk(gclk));
	jxor g0934(.dina(w_n997_0[1]),.dinb(w_n944_0[1]),.dout(n998),.clk(gclk));
	jxor g0935(.dina(w_n998_0[1]),.dinb(w_n942_0[1]),.dout(n999),.clk(gclk));
	jxor g0936(.dina(w_n999_0[1]),.dinb(w_n939_0[1]),.dout(n1000),.clk(gclk));
	jxor g0937(.dina(w_n1000_0[1]),.dinb(w_n937_0[1]),.dout(n1001),.clk(gclk));
	jxor g0938(.dina(w_n1001_0[1]),.dinb(w_n934_0[1]),.dout(n1002),.clk(gclk));
	jxor g0939(.dina(w_n1002_0[1]),.dinb(w_n932_0[1]),.dout(n1003),.clk(gclk));
	jxor g0940(.dina(w_n1003_0[1]),.dinb(w_n929_0[1]),.dout(n1004),.clk(gclk));
	jxor g0941(.dina(w_n1004_0[1]),.dinb(w_n927_0[1]),.dout(n1005),.clk(gclk));
	jxor g0942(.dina(w_n1005_0[1]),.dinb(w_n924_0[1]),.dout(n1006),.clk(gclk));
	jxor g0943(.dina(w_n1006_0[1]),.dinb(w_n922_0[1]),.dout(n1007),.clk(gclk));
	jxor g0944(.dina(w_n1007_0[1]),.dinb(w_n916_0[1]),.dout(n1008),.clk(gclk));
	jnot g0945(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n915_0[2]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(n1010),.dinb(w_n911_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n910_0[1]),.dout(w_dff_A_okMi2w5I6_2),.clk(gclk));
	jand g0949(.dina(w_n1011_0[0]),.dinb(w_n910_0[0]),.dout(n1013),.clk(gclk));
	jor g0950(.dina(w_n1009_0[0]),.dinb(w_n915_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1008_0[0]),.dinb(w_n915_0[0]),.dout(n1015),.clk(gclk));
	jor g0952(.dina(n1015),.dinb(w_n911_0[0]),.dout(n1016),.clk(gclk));
	jand g0953(.dina(n1016),.dinb(w_dff_B_ha1f2K3W5_1),.dout(n1017),.clk(gclk));
	jand g0954(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1018),.clk(gclk));
	jnot g0955(.din(w_n1006_0[0]),.dout(n1019),.clk(gclk));
	jor g0956(.dina(n1019),.dinb(w_n922_0[0]),.dout(n1020),.clk(gclk));
	jor g0957(.dina(w_n1007_0[0]),.dinb(w_n916_0[0]),.dout(n1021),.clk(gclk));
	jand g0958(.dina(n1021),.dinb(w_dff_B_YGBk4d6B0_1),.dout(n1022),.clk(gclk));
	jand g0959(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1023),.clk(gclk));
	jand g0960(.dina(w_n1004_0[0]),.dinb(w_n927_0[0]),.dout(n1024),.clk(gclk));
	jand g0961(.dina(w_n1005_0[0]),.dinb(w_n924_0[0]),.dout(n1025),.clk(gclk));
	jor g0962(.dina(n1025),.dinb(w_dff_B_hUWPJ5Ia0_1),.dout(n1026),.clk(gclk));
	jand g0963(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1027),.clk(gclk));
	jnot g0964(.din(n1027),.dout(n1028),.clk(gclk));
	jand g0965(.dina(w_n1002_0[0]),.dinb(w_n932_0[0]),.dout(n1029),.clk(gclk));
	jand g0966(.dina(w_n1003_0[0]),.dinb(w_n929_0[0]),.dout(n1030),.clk(gclk));
	jor g0967(.dina(n1030),.dinb(w_dff_B_h5RKjoXL7_1),.dout(n1031),.clk(gclk));
	jand g0968(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1032),.clk(gclk));
	jnot g0969(.din(n1032),.dout(n1033),.clk(gclk));
	jand g0970(.dina(w_n1000_0[0]),.dinb(w_n937_0[0]),.dout(n1034),.clk(gclk));
	jand g0971(.dina(w_n1001_0[0]),.dinb(w_n934_0[0]),.dout(n1035),.clk(gclk));
	jor g0972(.dina(n1035),.dinb(w_dff_B_TOvxfCyx5_1),.dout(n1036),.clk(gclk));
	jand g0973(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1037),.clk(gclk));
	jnot g0974(.din(n1037),.dout(n1038),.clk(gclk));
	jand g0975(.dina(w_n998_0[0]),.dinb(w_n942_0[0]),.dout(n1039),.clk(gclk));
	jand g0976(.dina(w_n999_0[0]),.dinb(w_n939_0[0]),.dout(n1040),.clk(gclk));
	jor g0977(.dina(n1040),.dinb(w_dff_B_X9x5eONG1_1),.dout(n1041),.clk(gclk));
	jand g0978(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1042),.clk(gclk));
	jnot g0979(.din(n1042),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_n996_0[0]),.dinb(w_n947_0[0]),.dout(n1044),.clk(gclk));
	jand g0981(.dina(w_n997_0[0]),.dinb(w_n944_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(w_dff_B_fiFeTNe63_1),.dout(n1046),.clk(gclk));
	jand g0983(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1047),.clk(gclk));
	jnot g0984(.din(n1047),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_n994_0[0]),.dinb(w_n952_0[0]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n995_0[0]),.dinb(w_n949_0[0]),.dout(n1050),.clk(gclk));
	jor g0987(.dina(n1050),.dinb(w_dff_B_VQ99M6Cp9_1),.dout(n1051),.clk(gclk));
	jand g0988(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1052),.clk(gclk));
	jnot g0989(.din(n1052),.dout(n1053),.clk(gclk));
	jand g0990(.dina(w_n992_0[0]),.dinb(w_n957_0[0]),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n993_0[0]),.dinb(w_n954_0[0]),.dout(n1055),.clk(gclk));
	jor g0992(.dina(n1055),.dinb(w_dff_B_4uKjXcCu3_1),.dout(n1056),.clk(gclk));
	jand g0993(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1057),.clk(gclk));
	jnot g0994(.din(n1057),.dout(n1058),.clk(gclk));
	jand g0995(.dina(w_n990_0[0]),.dinb(w_n962_0[0]),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n991_0[0]),.dinb(w_n959_0[0]),.dout(n1060),.clk(gclk));
	jor g0997(.dina(n1060),.dinb(w_dff_B_Fipv8Gnp4_1),.dout(n1061),.clk(gclk));
	jand g0998(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1062),.clk(gclk));
	jnot g0999(.din(n1062),.dout(n1063),.clk(gclk));
	jand g1000(.dina(w_n988_0[0]),.dinb(w_n967_0[0]),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n989_0[0]),.dinb(w_n964_0[0]),.dout(n1065),.clk(gclk));
	jor g1002(.dina(n1065),.dinb(w_dff_B_tEIsuwSY6_1),.dout(n1066),.clk(gclk));
	jand g1003(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1067),.clk(gclk));
	jnot g1004(.din(n1067),.dout(n1068),.clk(gclk));
	jand g1005(.dina(w_n986_0[0]),.dinb(w_n972_0[0]),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n987_0[0]),.dinb(w_n969_0[0]),.dout(n1070),.clk(gclk));
	jor g1007(.dina(n1070),.dinb(w_dff_B_zrwX1Wfj8_1),.dout(n1071),.clk(gclk));
	jand g1008(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1072),.clk(gclk));
	jnot g1009(.din(n1072),.dout(n1073),.clk(gclk));
	jand g1010(.dina(w_n984_0[0]),.dinb(w_n978_0[0]),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n985_0[0]),.dinb(w_n974_0[0]),.dout(n1075),.clk(gclk));
	jor g1012(.dina(n1075),.dinb(w_dff_B_Kvu2NZ8E1_1),.dout(n1076),.clk(gclk));
	jand g1013(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G307gat_2[1]),.dinb(w_G256gat_6[2]),.dout(n1078),.clk(gclk));
	jor g1015(.dina(w_n983_0[0]),.dinb(w_n982_0[0]),.dout(n1079),.clk(gclk));
	jand g1016(.dina(n1079),.dinb(w_n980_0[0]),.dout(n1080),.clk(gclk));
	jxor g1017(.dina(w_n1080_0[1]),.dinb(w_n1078_0[1]),.dout(n1081),.clk(gclk));
	jnot g1018(.din(n1081),.dout(n1082),.clk(gclk));
	jxor g1019(.dina(w_n1082_0[1]),.dinb(w_n1077_0[1]),.dout(n1083),.clk(gclk));
	jxor g1020(.dina(w_n1083_0[1]),.dinb(w_n1076_0[1]),.dout(n1084),.clk(gclk));
	jxor g1021(.dina(w_n1084_0[1]),.dinb(w_n1073_0[1]),.dout(n1085),.clk(gclk));
	jxor g1022(.dina(w_n1085_0[1]),.dinb(w_n1071_0[1]),.dout(n1086),.clk(gclk));
	jxor g1023(.dina(w_n1086_0[1]),.dinb(w_n1068_0[1]),.dout(n1087),.clk(gclk));
	jxor g1024(.dina(w_n1087_0[1]),.dinb(w_n1066_0[1]),.dout(n1088),.clk(gclk));
	jxor g1025(.dina(w_n1088_0[1]),.dinb(w_n1063_0[1]),.dout(n1089),.clk(gclk));
	jxor g1026(.dina(w_n1089_0[1]),.dinb(w_n1061_0[1]),.dout(n1090),.clk(gclk));
	jxor g1027(.dina(w_n1090_0[1]),.dinb(w_n1058_0[1]),.dout(n1091),.clk(gclk));
	jxor g1028(.dina(w_n1091_0[1]),.dinb(w_n1056_0[1]),.dout(n1092),.clk(gclk));
	jxor g1029(.dina(w_n1092_0[1]),.dinb(w_n1053_0[1]),.dout(n1093),.clk(gclk));
	jxor g1030(.dina(w_n1093_0[1]),.dinb(w_n1051_0[1]),.dout(n1094),.clk(gclk));
	jxor g1031(.dina(w_n1094_0[1]),.dinb(w_n1048_0[1]),.dout(n1095),.clk(gclk));
	jxor g1032(.dina(w_n1095_0[1]),.dinb(w_n1046_0[1]),.dout(n1096),.clk(gclk));
	jxor g1033(.dina(w_n1096_0[1]),.dinb(w_n1043_0[1]),.dout(n1097),.clk(gclk));
	jxor g1034(.dina(w_n1097_0[1]),.dinb(w_n1041_0[1]),.dout(n1098),.clk(gclk));
	jxor g1035(.dina(w_n1098_0[1]),.dinb(w_n1038_0[1]),.dout(n1099),.clk(gclk));
	jxor g1036(.dina(w_n1099_0[1]),.dinb(w_n1036_0[1]),.dout(n1100),.clk(gclk));
	jxor g1037(.dina(w_n1100_0[1]),.dinb(w_n1033_0[1]),.dout(n1101),.clk(gclk));
	jxor g1038(.dina(w_n1101_0[1]),.dinb(w_n1031_0[1]),.dout(n1102),.clk(gclk));
	jxor g1039(.dina(w_n1102_0[1]),.dinb(w_n1028_0[1]),.dout(n1103),.clk(gclk));
	jxor g1040(.dina(w_n1103_0[1]),.dinb(w_n1026_0[1]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(n1104),.dout(n1105),.clk(gclk));
	jxor g1042(.dina(w_n1105_0[1]),.dinb(w_n1023_0[1]),.dout(n1106),.clk(gclk));
	jxor g1043(.dina(w_n1106_0[1]),.dinb(w_n1022_0[1]),.dout(n1107),.clk(gclk));
	jxor g1044(.dina(w_n1107_0[1]),.dinb(w_n1018_0[1]),.dout(n1108),.clk(gclk));
	jxor g1045(.dina(w_n1108_0[1]),.dinb(w_n1017_0[1]),.dout(n1109),.clk(gclk));
	jnot g1046(.din(w_n1109_0[1]),.dout(n1110),.clk(gclk));
	jxor g1047(.dina(n1110),.dinb(w_n1013_0[1]),.dout(w_dff_A_3iIVPtIy0_2),.clk(gclk));
	jnot g1048(.din(w_n1108_0[0]),.dout(n1112),.clk(gclk));
	jor g1049(.dina(n1112),.dinb(w_n1017_0[0]),.dout(n1113),.clk(gclk));
	jor g1050(.dina(w_n1109_0[0]),.dinb(w_n1013_0[0]),.dout(n1114),.clk(gclk));
	jand g1051(.dina(n1114),.dinb(w_dff_B_RwNnqVnb6_1),.dout(n1115),.clk(gclk));
	jnot g1052(.din(w_n1106_0[0]),.dout(n1116),.clk(gclk));
	jor g1053(.dina(n1116),.dinb(w_n1022_0[0]),.dout(n1117),.clk(gclk));
	jor g1054(.dina(w_n1107_0[0]),.dinb(w_n1018_0[0]),.dout(n1118),.clk(gclk));
	jand g1055(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jand g1056(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1120),.clk(gclk));
	jand g1057(.dina(w_n1103_0[0]),.dinb(w_n1026_0[0]),.dout(n1121),.clk(gclk));
	jnot g1058(.din(n1121),.dout(n1122),.clk(gclk));
	jor g1059(.dina(w_n1105_0[0]),.dinb(w_n1023_0[0]),.dout(n1123),.clk(gclk));
	jand g1060(.dina(n1123),.dinb(w_dff_B_DqGxwHbC1_1),.dout(n1124),.clk(gclk));
	jand g1061(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1125),.clk(gclk));
	jnot g1062(.din(n1125),.dout(n1126),.clk(gclk));
	jand g1063(.dina(w_n1101_0[0]),.dinb(w_n1031_0[0]),.dout(n1127),.clk(gclk));
	jand g1064(.dina(w_n1102_0[0]),.dinb(w_n1028_0[0]),.dout(n1128),.clk(gclk));
	jor g1065(.dina(n1128),.dinb(w_dff_B_sd11iQz02_1),.dout(n1129),.clk(gclk));
	jand g1066(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1130),.clk(gclk));
	jnot g1067(.din(n1130),.dout(n1131),.clk(gclk));
	jand g1068(.dina(w_n1099_0[0]),.dinb(w_n1036_0[0]),.dout(n1132),.clk(gclk));
	jand g1069(.dina(w_n1100_0[0]),.dinb(w_n1033_0[0]),.dout(n1133),.clk(gclk));
	jor g1070(.dina(n1133),.dinb(w_dff_B_LiVhcqFl1_1),.dout(n1134),.clk(gclk));
	jand g1071(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1135),.clk(gclk));
	jnot g1072(.din(n1135),.dout(n1136),.clk(gclk));
	jand g1073(.dina(w_n1097_0[0]),.dinb(w_n1041_0[0]),.dout(n1137),.clk(gclk));
	jand g1074(.dina(w_n1098_0[0]),.dinb(w_n1038_0[0]),.dout(n1138),.clk(gclk));
	jor g1075(.dina(n1138),.dinb(w_dff_B_FmIUrn9u6_1),.dout(n1139),.clk(gclk));
	jand g1076(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1140),.clk(gclk));
	jnot g1077(.din(n1140),.dout(n1141),.clk(gclk));
	jand g1078(.dina(w_n1095_0[0]),.dinb(w_n1046_0[0]),.dout(n1142),.clk(gclk));
	jand g1079(.dina(w_n1096_0[0]),.dinb(w_n1043_0[0]),.dout(n1143),.clk(gclk));
	jor g1080(.dina(n1143),.dinb(w_dff_B_Ks3Cgzof9_1),.dout(n1144),.clk(gclk));
	jand g1081(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1145),.clk(gclk));
	jnot g1082(.din(n1145),.dout(n1146),.clk(gclk));
	jand g1083(.dina(w_n1093_0[0]),.dinb(w_n1051_0[0]),.dout(n1147),.clk(gclk));
	jand g1084(.dina(w_n1094_0[0]),.dinb(w_n1048_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(w_dff_B_LQq7XSgV1_1),.dout(n1149),.clk(gclk));
	jand g1086(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1150),.clk(gclk));
	jnot g1087(.din(n1150),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_n1091_0[0]),.dinb(w_n1056_0[0]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1092_0[0]),.dinb(w_n1053_0[0]),.dout(n1153),.clk(gclk));
	jor g1090(.dina(n1153),.dinb(w_dff_B_OjcRlY2h2_1),.dout(n1154),.clk(gclk));
	jand g1091(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1155),.clk(gclk));
	jnot g1092(.din(n1155),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_n1089_0[0]),.dinb(w_n1061_0[0]),.dout(n1157),.clk(gclk));
	jand g1094(.dina(w_n1090_0[0]),.dinb(w_n1058_0[0]),.dout(n1158),.clk(gclk));
	jor g1095(.dina(n1158),.dinb(w_dff_B_QMF8uRl06_1),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1160),.clk(gclk));
	jnot g1097(.din(n1160),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_n1087_0[0]),.dinb(w_n1066_0[0]),.dout(n1162),.clk(gclk));
	jand g1099(.dina(w_n1088_0[0]),.dinb(w_n1063_0[0]),.dout(n1163),.clk(gclk));
	jor g1100(.dina(n1163),.dinb(w_dff_B_S4B5uJt66_1),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1165),.clk(gclk));
	jnot g1102(.din(n1165),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_n1085_0[0]),.dinb(w_n1071_0[0]),.dout(n1167),.clk(gclk));
	jand g1104(.dina(w_n1086_0[0]),.dinb(w_n1068_0[0]),.dout(n1168),.clk(gclk));
	jor g1105(.dina(n1168),.dinb(w_dff_B_RyEVqxOx9_1),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1170),.clk(gclk));
	jnot g1107(.din(n1170),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_n1083_0[0]),.dinb(w_n1076_0[0]),.dout(n1172),.clk(gclk));
	jand g1109(.dina(w_n1084_0[0]),.dinb(w_n1073_0[0]),.dout(n1173),.clk(gclk));
	jor g1110(.dina(n1173),.dinb(w_dff_B_5fzawKms6_1),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1175),.clk(gclk));
	jand g1112(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1176),.clk(gclk));
	jor g1113(.dina(w_n1080_0[0]),.dinb(w_n1078_0[0]),.dout(n1177),.clk(gclk));
	jor g1114(.dina(w_n1082_0[0]),.dinb(w_n1077_0[0]),.dout(n1178),.clk(gclk));
	jand g1115(.dina(n1178),.dinb(w_dff_B_SD9sF0Cs1_1),.dout(n1179),.clk(gclk));
	jxor g1116(.dina(w_n1179_0[1]),.dinb(w_n1176_0[1]),.dout(n1180),.clk(gclk));
	jnot g1117(.din(n1180),.dout(n1181),.clk(gclk));
	jxor g1118(.dina(w_n1181_0[1]),.dinb(w_n1175_0[1]),.dout(n1182),.clk(gclk));
	jxor g1119(.dina(w_n1182_0[1]),.dinb(w_n1174_0[1]),.dout(n1183),.clk(gclk));
	jxor g1120(.dina(w_n1183_0[1]),.dinb(w_n1171_0[1]),.dout(n1184),.clk(gclk));
	jxor g1121(.dina(w_n1184_0[1]),.dinb(w_n1169_0[1]),.dout(n1185),.clk(gclk));
	jxor g1122(.dina(w_n1185_0[1]),.dinb(w_n1166_0[1]),.dout(n1186),.clk(gclk));
	jxor g1123(.dina(w_n1186_0[1]),.dinb(w_n1164_0[1]),.dout(n1187),.clk(gclk));
	jxor g1124(.dina(w_n1187_0[1]),.dinb(w_n1161_0[1]),.dout(n1188),.clk(gclk));
	jxor g1125(.dina(w_n1188_0[1]),.dinb(w_n1159_0[1]),.dout(n1189),.clk(gclk));
	jxor g1126(.dina(w_n1189_0[1]),.dinb(w_n1156_0[1]),.dout(n1190),.clk(gclk));
	jxor g1127(.dina(w_n1190_0[1]),.dinb(w_n1154_0[1]),.dout(n1191),.clk(gclk));
	jxor g1128(.dina(w_n1191_0[1]),.dinb(w_n1151_0[1]),.dout(n1192),.clk(gclk));
	jxor g1129(.dina(w_n1192_0[1]),.dinb(w_n1149_0[1]),.dout(n1193),.clk(gclk));
	jxor g1130(.dina(w_n1193_0[1]),.dinb(w_n1146_0[1]),.dout(n1194),.clk(gclk));
	jxor g1131(.dina(w_n1194_0[1]),.dinb(w_n1144_0[1]),.dout(n1195),.clk(gclk));
	jxor g1132(.dina(w_n1195_0[1]),.dinb(w_n1141_0[1]),.dout(n1196),.clk(gclk));
	jxor g1133(.dina(w_n1196_0[1]),.dinb(w_n1139_0[1]),.dout(n1197),.clk(gclk));
	jxor g1134(.dina(w_n1197_0[1]),.dinb(w_n1136_0[1]),.dout(n1198),.clk(gclk));
	jxor g1135(.dina(w_n1198_0[1]),.dinb(w_n1134_0[1]),.dout(n1199),.clk(gclk));
	jxor g1136(.dina(w_n1199_0[1]),.dinb(w_n1131_0[1]),.dout(n1200),.clk(gclk));
	jxor g1137(.dina(w_n1200_0[1]),.dinb(w_n1129_0[1]),.dout(n1201),.clk(gclk));
	jxor g1138(.dina(w_n1201_0[1]),.dinb(w_n1126_0[1]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jxor g1140(.dina(w_n1203_0[1]),.dinb(w_n1124_0[1]),.dout(n1204),.clk(gclk));
	jnot g1141(.din(n1204),.dout(n1205),.clk(gclk));
	jxor g1142(.dina(w_n1205_0[1]),.dinb(w_n1120_0[1]),.dout(n1206),.clk(gclk));
	jxor g1143(.dina(w_n1206_0[1]),.dinb(w_n1119_0[1]),.dout(n1207),.clk(gclk));
	jnot g1144(.din(w_n1207_0[1]),.dout(n1208),.clk(gclk));
	jxor g1145(.dina(n1208),.dinb(w_n1115_0[1]),.dout(w_dff_A_UyaYymEo5_2),.clk(gclk));
	jnot g1146(.din(w_n1206_0[0]),.dout(n1210),.clk(gclk));
	jor g1147(.dina(n1210),.dinb(w_n1119_0[0]),.dout(n1211),.clk(gclk));
	jor g1148(.dina(w_n1207_0[0]),.dinb(w_n1115_0[0]),.dout(n1212),.clk(gclk));
	jand g1149(.dina(n1212),.dinb(w_dff_B_4lbaaL8i8_1),.dout(n1213),.clk(gclk));
	jor g1150(.dina(w_n1203_0[0]),.dinb(w_n1124_0[0]),.dout(n1214),.clk(gclk));
	jor g1151(.dina(w_n1205_0[0]),.dinb(w_n1120_0[0]),.dout(n1215),.clk(gclk));
	jand g1152(.dina(n1215),.dinb(w_dff_B_bDw6z2Oz2_1),.dout(n1216),.clk(gclk));
	jand g1153(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1217),.clk(gclk));
	jand g1154(.dina(w_n1200_0[0]),.dinb(w_n1129_0[0]),.dout(n1218),.clk(gclk));
	jand g1155(.dina(w_n1201_0[0]),.dinb(w_n1126_0[0]),.dout(n1219),.clk(gclk));
	jor g1156(.dina(n1219),.dinb(w_dff_B_PIGqr8be1_1),.dout(n1220),.clk(gclk));
	jand g1157(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1221),.clk(gclk));
	jnot g1158(.din(n1221),.dout(n1222),.clk(gclk));
	jand g1159(.dina(w_n1198_0[0]),.dinb(w_n1134_0[0]),.dout(n1223),.clk(gclk));
	jand g1160(.dina(w_n1199_0[0]),.dinb(w_n1131_0[0]),.dout(n1224),.clk(gclk));
	jor g1161(.dina(n1224),.dinb(w_dff_B_6d1qojQz1_1),.dout(n1225),.clk(gclk));
	jand g1162(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1226),.clk(gclk));
	jnot g1163(.din(n1226),.dout(n1227),.clk(gclk));
	jand g1164(.dina(w_n1196_0[0]),.dinb(w_n1139_0[0]),.dout(n1228),.clk(gclk));
	jand g1165(.dina(w_n1197_0[0]),.dinb(w_n1136_0[0]),.dout(n1229),.clk(gclk));
	jor g1166(.dina(n1229),.dinb(w_dff_B_eWRukfmw4_1),.dout(n1230),.clk(gclk));
	jand g1167(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1231),.clk(gclk));
	jnot g1168(.din(n1231),.dout(n1232),.clk(gclk));
	jand g1169(.dina(w_n1194_0[0]),.dinb(w_n1144_0[0]),.dout(n1233),.clk(gclk));
	jand g1170(.dina(w_n1195_0[0]),.dinb(w_n1141_0[0]),.dout(n1234),.clk(gclk));
	jor g1171(.dina(n1234),.dinb(w_dff_B_wqdKiwbS9_1),.dout(n1235),.clk(gclk));
	jand g1172(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1236),.clk(gclk));
	jnot g1173(.din(n1236),.dout(n1237),.clk(gclk));
	jand g1174(.dina(w_n1192_0[0]),.dinb(w_n1149_0[0]),.dout(n1238),.clk(gclk));
	jand g1175(.dina(w_n1193_0[0]),.dinb(w_n1146_0[0]),.dout(n1239),.clk(gclk));
	jor g1176(.dina(n1239),.dinb(w_dff_B_CsyphyLd6_1),.dout(n1240),.clk(gclk));
	jand g1177(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1241),.clk(gclk));
	jnot g1178(.din(n1241),.dout(n1242),.clk(gclk));
	jand g1179(.dina(w_n1190_0[0]),.dinb(w_n1154_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(w_n1191_0[0]),.dinb(w_n1151_0[0]),.dout(n1244),.clk(gclk));
	jor g1181(.dina(n1244),.dinb(w_dff_B_kV5BDMjF1_1),.dout(n1245),.clk(gclk));
	jand g1182(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1246),.clk(gclk));
	jnot g1183(.din(n1246),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_n1188_0[0]),.dinb(w_n1159_0[0]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1189_0[0]),.dinb(w_n1156_0[0]),.dout(n1249),.clk(gclk));
	jor g1186(.dina(n1249),.dinb(w_dff_B_D0MLO62s7_1),.dout(n1250),.clk(gclk));
	jand g1187(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1251),.clk(gclk));
	jnot g1188(.din(n1251),.dout(n1252),.clk(gclk));
	jand g1189(.dina(w_n1186_0[0]),.dinb(w_n1164_0[0]),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1187_0[0]),.dinb(w_n1161_0[0]),.dout(n1254),.clk(gclk));
	jor g1191(.dina(n1254),.dinb(w_dff_B_8eTcrcM07_1),.dout(n1255),.clk(gclk));
	jand g1192(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1256),.clk(gclk));
	jnot g1193(.din(n1256),.dout(n1257),.clk(gclk));
	jand g1194(.dina(w_n1184_0[0]),.dinb(w_n1169_0[0]),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1185_0[0]),.dinb(w_n1166_0[0]),.dout(n1259),.clk(gclk));
	jor g1196(.dina(n1259),.dinb(w_dff_B_bVIrtuqp5_1),.dout(n1260),.clk(gclk));
	jand g1197(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1261),.clk(gclk));
	jnot g1198(.din(n1261),.dout(n1262),.clk(gclk));
	jand g1199(.dina(w_n1182_0[0]),.dinb(w_n1174_0[0]),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1183_0[0]),.dinb(w_n1171_0[0]),.dout(n1264),.clk(gclk));
	jor g1201(.dina(n1264),.dinb(w_dff_B_aeNosS844_1),.dout(n1265),.clk(gclk));
	jand g1202(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1267),.clk(gclk));
	jor g1204(.dina(w_n1179_0[0]),.dinb(w_n1176_0[0]),.dout(n1268),.clk(gclk));
	jor g1205(.dina(w_n1181_0[0]),.dinb(w_n1175_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(n1269),.dinb(w_dff_B_DIHpMLGD7_1),.dout(n1270),.clk(gclk));
	jxor g1207(.dina(w_n1270_0[1]),.dinb(w_n1267_0[1]),.dout(n1271),.clk(gclk));
	jnot g1208(.din(n1271),.dout(n1272),.clk(gclk));
	jxor g1209(.dina(w_n1272_0[1]),.dinb(w_n1266_0[1]),.dout(n1273),.clk(gclk));
	jxor g1210(.dina(w_n1273_0[1]),.dinb(w_n1265_0[1]),.dout(n1274),.clk(gclk));
	jxor g1211(.dina(w_n1274_0[1]),.dinb(w_n1262_0[1]),.dout(n1275),.clk(gclk));
	jxor g1212(.dina(w_n1275_0[1]),.dinb(w_n1260_0[1]),.dout(n1276),.clk(gclk));
	jxor g1213(.dina(w_n1276_0[1]),.dinb(w_n1257_0[1]),.dout(n1277),.clk(gclk));
	jxor g1214(.dina(w_n1277_0[1]),.dinb(w_n1255_0[1]),.dout(n1278),.clk(gclk));
	jxor g1215(.dina(w_n1278_0[1]),.dinb(w_n1252_0[1]),.dout(n1279),.clk(gclk));
	jxor g1216(.dina(w_n1279_0[1]),.dinb(w_n1250_0[1]),.dout(n1280),.clk(gclk));
	jxor g1217(.dina(w_n1280_0[1]),.dinb(w_n1247_0[1]),.dout(n1281),.clk(gclk));
	jxor g1218(.dina(w_n1281_0[1]),.dinb(w_n1245_0[1]),.dout(n1282),.clk(gclk));
	jxor g1219(.dina(w_n1282_0[1]),.dinb(w_n1242_0[1]),.dout(n1283),.clk(gclk));
	jxor g1220(.dina(w_n1283_0[1]),.dinb(w_n1240_0[1]),.dout(n1284),.clk(gclk));
	jxor g1221(.dina(w_n1284_0[1]),.dinb(w_n1237_0[1]),.dout(n1285),.clk(gclk));
	jxor g1222(.dina(w_n1285_0[1]),.dinb(w_n1235_0[1]),.dout(n1286),.clk(gclk));
	jxor g1223(.dina(w_n1286_0[1]),.dinb(w_n1232_0[1]),.dout(n1287),.clk(gclk));
	jxor g1224(.dina(w_n1287_0[1]),.dinb(w_n1230_0[1]),.dout(n1288),.clk(gclk));
	jxor g1225(.dina(w_n1288_0[1]),.dinb(w_n1227_0[1]),.dout(n1289),.clk(gclk));
	jxor g1226(.dina(w_n1289_0[1]),.dinb(w_n1225_0[1]),.dout(n1290),.clk(gclk));
	jxor g1227(.dina(w_n1290_0[1]),.dinb(w_n1222_0[1]),.dout(n1291),.clk(gclk));
	jxor g1228(.dina(w_n1291_0[1]),.dinb(w_n1220_0[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jxor g1230(.dina(w_n1293_0[1]),.dinb(w_n1217_0[1]),.dout(n1294),.clk(gclk));
	jxor g1231(.dina(w_n1294_0[1]),.dinb(w_n1216_0[1]),.dout(n1295),.clk(gclk));
	jnot g1232(.din(w_n1295_0[1]),.dout(n1296),.clk(gclk));
	jxor g1233(.dina(w_dff_B_z8w0zcKB8_0),.dinb(w_n1213_0[1]),.dout(w_dff_A_5lkC1ky40_2),.clk(gclk));
	jnot g1234(.din(w_n1294_0[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(w_dff_B_LoIPBci80_0),.dinb(w_n1216_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1295_0[0]),.dinb(w_n1213_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(w_dff_B_kUkGjYFU6_1),.dout(n1301),.clk(gclk));
	jnot g1238(.din(w_n1220_0[0]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(w_n1291_0[0]),.dout(n1303),.clk(gclk));
	jor g1240(.dina(w_dff_B_qZbCVfzj9_0),.dinb(n1302),.dout(n1304),.clk(gclk));
	jor g1241(.dina(w_n1293_0[0]),.dinb(w_n1217_0[0]),.dout(n1305),.clk(gclk));
	jand g1242(.dina(n1305),.dinb(w_dff_B_QzRqY8Wk5_1),.dout(n1306),.clk(gclk));
	jand g1243(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1307),.clk(gclk));
	jand g1244(.dina(w_n1289_0[0]),.dinb(w_n1225_0[0]),.dout(n1308),.clk(gclk));
	jand g1245(.dina(w_n1290_0[0]),.dinb(w_n1222_0[0]),.dout(n1309),.clk(gclk));
	jor g1246(.dina(n1309),.dinb(w_dff_B_8gNLrgrL5_1),.dout(n1310),.clk(gclk));
	jand g1247(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1311),.clk(gclk));
	jnot g1248(.din(n1311),.dout(n1312),.clk(gclk));
	jand g1249(.dina(w_n1287_0[0]),.dinb(w_n1230_0[0]),.dout(n1313),.clk(gclk));
	jand g1250(.dina(w_n1288_0[0]),.dinb(w_n1227_0[0]),.dout(n1314),.clk(gclk));
	jor g1251(.dina(n1314),.dinb(w_dff_B_GkOsAjCA5_1),.dout(n1315),.clk(gclk));
	jand g1252(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1316),.clk(gclk));
	jnot g1253(.din(n1316),.dout(n1317),.clk(gclk));
	jand g1254(.dina(w_n1285_0[0]),.dinb(w_n1235_0[0]),.dout(n1318),.clk(gclk));
	jand g1255(.dina(w_n1286_0[0]),.dinb(w_n1232_0[0]),.dout(n1319),.clk(gclk));
	jor g1256(.dina(n1319),.dinb(w_dff_B_uDtCWuTI2_1),.dout(n1320),.clk(gclk));
	jand g1257(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1321),.clk(gclk));
	jnot g1258(.din(n1321),.dout(n1322),.clk(gclk));
	jand g1259(.dina(w_n1283_0[0]),.dinb(w_n1240_0[0]),.dout(n1323),.clk(gclk));
	jand g1260(.dina(w_n1284_0[0]),.dinb(w_n1237_0[0]),.dout(n1324),.clk(gclk));
	jor g1261(.dina(n1324),.dinb(w_dff_B_8fyuWS3C8_1),.dout(n1325),.clk(gclk));
	jand g1262(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(n1326),.dout(n1327),.clk(gclk));
	jand g1264(.dina(w_n1281_0[0]),.dinb(w_n1245_0[0]),.dout(n1328),.clk(gclk));
	jand g1265(.dina(w_n1282_0[0]),.dinb(w_n1242_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(n1329),.dinb(w_dff_B_UmQpK0rO6_1),.dout(n1330),.clk(gclk));
	jand g1267(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1331),.clk(gclk));
	jnot g1268(.din(n1331),.dout(n1332),.clk(gclk));
	jand g1269(.dina(w_n1279_0[0]),.dinb(w_n1250_0[0]),.dout(n1333),.clk(gclk));
	jand g1270(.dina(w_n1280_0[0]),.dinb(w_n1247_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(n1334),.dinb(w_dff_B_sVmjXq6O1_1),.dout(n1335),.clk(gclk));
	jand g1272(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1336),.clk(gclk));
	jnot g1273(.din(n1336),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_n1277_0[0]),.dinb(w_n1255_0[0]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1278_0[0]),.dinb(w_n1252_0[0]),.dout(n1339),.clk(gclk));
	jor g1276(.dina(n1339),.dinb(w_dff_B_fvBuavZm2_1),.dout(n1340),.clk(gclk));
	jand g1277(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1341),.clk(gclk));
	jnot g1278(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1279(.dina(w_n1275_0[0]),.dinb(w_n1260_0[0]),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1276_0[0]),.dinb(w_n1257_0[0]),.dout(n1344),.clk(gclk));
	jor g1281(.dina(n1344),.dinb(w_dff_B_JqAWgDf77_1),.dout(n1345),.clk(gclk));
	jand g1282(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1346),.clk(gclk));
	jnot g1283(.din(n1346),.dout(n1347),.clk(gclk));
	jand g1284(.dina(w_n1273_0[0]),.dinb(w_n1265_0[0]),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1274_0[0]),.dinb(w_n1262_0[0]),.dout(n1349),.clk(gclk));
	jor g1286(.dina(n1349),.dinb(w_dff_B_AqizxOau4_1),.dout(n1350),.clk(gclk));
	jand g1287(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1352),.clk(gclk));
	jor g1289(.dina(w_n1270_0[0]),.dinb(w_n1267_0[0]),.dout(n1353),.clk(gclk));
	jor g1290(.dina(w_n1272_0[0]),.dinb(w_n1266_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(n1354),.dinb(w_dff_B_niqKiDNW8_1),.dout(n1355),.clk(gclk));
	jxor g1292(.dina(w_n1355_0[1]),.dinb(w_n1352_0[1]),.dout(n1356),.clk(gclk));
	jnot g1293(.din(n1356),.dout(n1357),.clk(gclk));
	jxor g1294(.dina(w_n1357_0[1]),.dinb(w_n1351_0[1]),.dout(n1358),.clk(gclk));
	jxor g1295(.dina(w_n1358_0[1]),.dinb(w_n1350_0[1]),.dout(n1359),.clk(gclk));
	jxor g1296(.dina(w_n1359_0[1]),.dinb(w_n1347_0[1]),.dout(n1360),.clk(gclk));
	jxor g1297(.dina(w_n1360_0[1]),.dinb(w_n1345_0[1]),.dout(n1361),.clk(gclk));
	jxor g1298(.dina(w_n1361_0[1]),.dinb(w_n1342_0[1]),.dout(n1362),.clk(gclk));
	jxor g1299(.dina(w_n1362_0[1]),.dinb(w_n1340_0[1]),.dout(n1363),.clk(gclk));
	jxor g1300(.dina(w_n1363_0[1]),.dinb(w_n1337_0[1]),.dout(n1364),.clk(gclk));
	jxor g1301(.dina(w_n1364_0[1]),.dinb(w_n1335_0[1]),.dout(n1365),.clk(gclk));
	jxor g1302(.dina(w_n1365_0[1]),.dinb(w_n1332_0[1]),.dout(n1366),.clk(gclk));
	jxor g1303(.dina(w_n1366_0[1]),.dinb(w_n1330_0[1]),.dout(n1367),.clk(gclk));
	jxor g1304(.dina(w_n1367_0[1]),.dinb(w_n1327_0[1]),.dout(n1368),.clk(gclk));
	jxor g1305(.dina(w_n1368_0[1]),.dinb(w_n1325_0[1]),.dout(n1369),.clk(gclk));
	jxor g1306(.dina(w_n1369_0[1]),.dinb(w_n1322_0[1]),.dout(n1370),.clk(gclk));
	jxor g1307(.dina(w_n1370_0[1]),.dinb(w_n1320_0[1]),.dout(n1371),.clk(gclk));
	jxor g1308(.dina(w_n1371_0[1]),.dinb(w_n1317_0[1]),.dout(n1372),.clk(gclk));
	jxor g1309(.dina(w_n1372_0[1]),.dinb(w_n1315_0[1]),.dout(n1373),.clk(gclk));
	jxor g1310(.dina(w_n1373_0[1]),.dinb(w_n1312_0[1]),.dout(n1374),.clk(gclk));
	jxor g1311(.dina(w_n1374_0[1]),.dinb(w_n1310_0[1]),.dout(n1375),.clk(gclk));
	jnot g1312(.din(n1375),.dout(n1376),.clk(gclk));
	jxor g1313(.dina(w_n1376_0[1]),.dinb(w_n1307_0[1]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jxor g1315(.dina(w_n1378_0[1]),.dinb(w_n1306_0[1]),.dout(n1379),.clk(gclk));
	jxor g1316(.dina(w_n1379_0[1]),.dinb(w_n1301_0[1]),.dout(w_dff_A_yzVOykgA5_2),.clk(gclk));
	jor g1317(.dina(w_n1378_0[0]),.dinb(w_n1306_0[0]),.dout(n1381),.clk(gclk));
	jnot g1318(.din(w_n1379_0[0]),.dout(n1382),.clk(gclk));
	jor g1319(.dina(w_dff_B_ZlZ6Nbus7_0),.dinb(w_n1301_0[0]),.dout(n1383),.clk(gclk));
	jand g1320(.dina(n1383),.dinb(w_dff_B_5Qqva24S8_1),.dout(n1384),.clk(gclk));
	jnot g1321(.din(w_n1310_0[0]),.dout(n1385),.clk(gclk));
	jnot g1322(.din(w_n1374_0[0]),.dout(n1386),.clk(gclk));
	jor g1323(.dina(n1386),.dinb(n1385),.dout(n1387),.clk(gclk));
	jor g1324(.dina(w_n1376_0[0]),.dinb(w_n1307_0[0]),.dout(n1388),.clk(gclk));
	jand g1325(.dina(n1388),.dinb(w_dff_B_p8CFYD8r0_1),.dout(n1389),.clk(gclk));
	jand g1326(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1390),.clk(gclk));
	jand g1327(.dina(w_n1372_0[0]),.dinb(w_n1315_0[0]),.dout(n1391),.clk(gclk));
	jand g1328(.dina(w_n1373_0[0]),.dinb(w_n1312_0[0]),.dout(n1392),.clk(gclk));
	jor g1329(.dina(n1392),.dinb(w_dff_B_okZPYfUy4_1),.dout(n1393),.clk(gclk));
	jand g1330(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1394),.clk(gclk));
	jnot g1331(.din(n1394),.dout(n1395),.clk(gclk));
	jand g1332(.dina(w_n1370_0[0]),.dinb(w_n1320_0[0]),.dout(n1396),.clk(gclk));
	jand g1333(.dina(w_n1371_0[0]),.dinb(w_n1317_0[0]),.dout(n1397),.clk(gclk));
	jor g1334(.dina(n1397),.dinb(w_dff_B_48fLUiLC1_1),.dout(n1398),.clk(gclk));
	jand g1335(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1399),.clk(gclk));
	jnot g1336(.din(n1399),.dout(n1400),.clk(gclk));
	jand g1337(.dina(w_n1368_0[0]),.dinb(w_n1325_0[0]),.dout(n1401),.clk(gclk));
	jand g1338(.dina(w_n1369_0[0]),.dinb(w_n1322_0[0]),.dout(n1402),.clk(gclk));
	jor g1339(.dina(n1402),.dinb(w_dff_B_EEFDNy893_1),.dout(n1403),.clk(gclk));
	jand g1340(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1404),.clk(gclk));
	jnot g1341(.din(n1404),.dout(n1405),.clk(gclk));
	jand g1342(.dina(w_n1366_0[0]),.dinb(w_n1330_0[0]),.dout(n1406),.clk(gclk));
	jand g1343(.dina(w_n1367_0[0]),.dinb(w_n1327_0[0]),.dout(n1407),.clk(gclk));
	jor g1344(.dina(n1407),.dinb(w_dff_B_vokYGC0b9_1),.dout(n1408),.clk(gclk));
	jand g1345(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1409),.clk(gclk));
	jnot g1346(.din(n1409),.dout(n1410),.clk(gclk));
	jand g1347(.dina(w_n1364_0[0]),.dinb(w_n1335_0[0]),.dout(n1411),.clk(gclk));
	jand g1348(.dina(w_n1365_0[0]),.dinb(w_n1332_0[0]),.dout(n1412),.clk(gclk));
	jor g1349(.dina(n1412),.dinb(w_dff_B_Np1v8xsj0_1),.dout(n1413),.clk(gclk));
	jand g1350(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1414),.clk(gclk));
	jnot g1351(.din(n1414),.dout(n1415),.clk(gclk));
	jand g1352(.dina(w_n1362_0[0]),.dinb(w_n1340_0[0]),.dout(n1416),.clk(gclk));
	jand g1353(.dina(w_n1363_0[0]),.dinb(w_n1337_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(w_dff_B_P7pV3xtN2_1),.dout(n1418),.clk(gclk));
	jand g1355(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1419),.clk(gclk));
	jnot g1356(.din(n1419),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_n1360_0[0]),.dinb(w_n1345_0[0]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1361_0[0]),.dinb(w_n1342_0[0]),.dout(n1422),.clk(gclk));
	jor g1359(.dina(n1422),.dinb(w_dff_B_XCPKuwD08_1),.dout(n1423),.clk(gclk));
	jand g1360(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1424),.clk(gclk));
	jnot g1361(.din(n1424),.dout(n1425),.clk(gclk));
	jand g1362(.dina(w_n1358_0[0]),.dinb(w_n1350_0[0]),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1359_0[0]),.dinb(w_n1347_0[0]),.dout(n1427),.clk(gclk));
	jor g1364(.dina(n1427),.dinb(w_dff_B_Ep9cpCXH0_1),.dout(n1428),.clk(gclk));
	jand g1365(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1430),.clk(gclk));
	jor g1367(.dina(w_n1355_0[0]),.dinb(w_n1352_0[0]),.dout(n1431),.clk(gclk));
	jor g1368(.dina(w_n1357_0[0]),.dinb(w_n1351_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(n1432),.dinb(w_dff_B_L7a03A1l4_1),.dout(n1433),.clk(gclk));
	jxor g1370(.dina(w_n1433_0[1]),.dinb(w_n1430_0[1]),.dout(n1434),.clk(gclk));
	jnot g1371(.din(n1434),.dout(n1435),.clk(gclk));
	jxor g1372(.dina(w_n1435_0[1]),.dinb(w_n1429_0[1]),.dout(n1436),.clk(gclk));
	jxor g1373(.dina(w_n1436_0[1]),.dinb(w_n1428_0[1]),.dout(n1437),.clk(gclk));
	jxor g1374(.dina(w_n1437_0[1]),.dinb(w_n1425_0[1]),.dout(n1438),.clk(gclk));
	jxor g1375(.dina(w_n1438_0[1]),.dinb(w_n1423_0[1]),.dout(n1439),.clk(gclk));
	jxor g1376(.dina(w_n1439_0[1]),.dinb(w_n1420_0[1]),.dout(n1440),.clk(gclk));
	jxor g1377(.dina(w_n1440_0[1]),.dinb(w_n1418_0[1]),.dout(n1441),.clk(gclk));
	jxor g1378(.dina(w_n1441_0[1]),.dinb(w_n1415_0[1]),.dout(n1442),.clk(gclk));
	jxor g1379(.dina(w_n1442_0[1]),.dinb(w_n1413_0[1]),.dout(n1443),.clk(gclk));
	jxor g1380(.dina(w_n1443_0[1]),.dinb(w_n1410_0[1]),.dout(n1444),.clk(gclk));
	jxor g1381(.dina(w_n1444_0[1]),.dinb(w_n1408_0[1]),.dout(n1445),.clk(gclk));
	jxor g1382(.dina(w_n1445_0[1]),.dinb(w_n1405_0[1]),.dout(n1446),.clk(gclk));
	jxor g1383(.dina(w_n1446_0[1]),.dinb(w_n1403_0[1]),.dout(n1447),.clk(gclk));
	jxor g1384(.dina(w_n1447_0[1]),.dinb(w_n1400_0[1]),.dout(n1448),.clk(gclk));
	jxor g1385(.dina(w_n1448_0[1]),.dinb(w_n1398_0[1]),.dout(n1449),.clk(gclk));
	jxor g1386(.dina(w_n1449_0[1]),.dinb(w_n1395_0[1]),.dout(n1450),.clk(gclk));
	jxor g1387(.dina(w_n1450_0[1]),.dinb(w_n1393_0[1]),.dout(n1451),.clk(gclk));
	jnot g1388(.din(n1451),.dout(n1452),.clk(gclk));
	jxor g1389(.dina(w_n1452_0[1]),.dinb(w_n1390_0[1]),.dout(n1453),.clk(gclk));
	jnot g1390(.din(n1453),.dout(n1454),.clk(gclk));
	jxor g1391(.dina(w_n1454_0[1]),.dinb(w_n1389_0[1]),.dout(n1455),.clk(gclk));
	jxor g1392(.dina(w_n1455_0[1]),.dinb(w_n1384_0[1]),.dout(w_dff_A_CdP4FEpr4_2),.clk(gclk));
	jor g1393(.dina(w_n1454_0[0]),.dinb(w_n1389_0[0]),.dout(n1457),.clk(gclk));
	jnot g1394(.din(w_n1455_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(w_dff_B_HRfc0iEy8_0),.dinb(w_n1384_0[0]),.dout(n1459),.clk(gclk));
	jand g1396(.dina(n1459),.dinb(w_dff_B_6M8TUMrb7_1),.dout(n1460),.clk(gclk));
	jnot g1397(.din(w_n1393_0[0]),.dout(n1461),.clk(gclk));
	jnot g1398(.din(w_n1450_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(n1462),.dinb(n1461),.dout(n1463),.clk(gclk));
	jor g1400(.dina(w_n1452_0[0]),.dinb(w_n1390_0[0]),.dout(n1464),.clk(gclk));
	jand g1401(.dina(n1464),.dinb(w_dff_B_3QFD0j615_1),.dout(n1465),.clk(gclk));
	jand g1402(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1466),.clk(gclk));
	jand g1403(.dina(w_n1448_0[0]),.dinb(w_n1398_0[0]),.dout(n1467),.clk(gclk));
	jand g1404(.dina(w_n1449_0[0]),.dinb(w_n1395_0[0]),.dout(n1468),.clk(gclk));
	jor g1405(.dina(n1468),.dinb(w_dff_B_JumOCHSu3_1),.dout(n1469),.clk(gclk));
	jand g1406(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1470),.clk(gclk));
	jnot g1407(.din(n1470),.dout(n1471),.clk(gclk));
	jand g1408(.dina(w_n1446_0[0]),.dinb(w_n1403_0[0]),.dout(n1472),.clk(gclk));
	jand g1409(.dina(w_n1447_0[0]),.dinb(w_n1400_0[0]),.dout(n1473),.clk(gclk));
	jor g1410(.dina(n1473),.dinb(w_dff_B_0Um9Rg9s4_1),.dout(n1474),.clk(gclk));
	jand g1411(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1475),.clk(gclk));
	jnot g1412(.din(n1475),.dout(n1476),.clk(gclk));
	jand g1413(.dina(w_n1444_0[0]),.dinb(w_n1408_0[0]),.dout(n1477),.clk(gclk));
	jand g1414(.dina(w_n1445_0[0]),.dinb(w_n1405_0[0]),.dout(n1478),.clk(gclk));
	jor g1415(.dina(n1478),.dinb(w_dff_B_zf6t6t9G7_1),.dout(n1479),.clk(gclk));
	jand g1416(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1480),.clk(gclk));
	jnot g1417(.din(n1480),.dout(n1481),.clk(gclk));
	jand g1418(.dina(w_n1442_0[0]),.dinb(w_n1413_0[0]),.dout(n1482),.clk(gclk));
	jand g1419(.dina(w_n1443_0[0]),.dinb(w_n1410_0[0]),.dout(n1483),.clk(gclk));
	jor g1420(.dina(n1483),.dinb(w_dff_B_ISJUd31I5_1),.dout(n1484),.clk(gclk));
	jand g1421(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1485),.clk(gclk));
	jnot g1422(.din(n1485),.dout(n1486),.clk(gclk));
	jand g1423(.dina(w_n1440_0[0]),.dinb(w_n1418_0[0]),.dout(n1487),.clk(gclk));
	jand g1424(.dina(w_n1441_0[0]),.dinb(w_n1415_0[0]),.dout(n1488),.clk(gclk));
	jor g1425(.dina(n1488),.dinb(w_dff_B_IFTw00kJ0_1),.dout(n1489),.clk(gclk));
	jand g1426(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1490),.clk(gclk));
	jnot g1427(.din(n1490),.dout(n1491),.clk(gclk));
	jand g1428(.dina(w_n1438_0[0]),.dinb(w_n1423_0[0]),.dout(n1492),.clk(gclk));
	jand g1429(.dina(w_n1439_0[0]),.dinb(w_n1420_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(w_dff_B_ho8lWHFt5_1),.dout(n1494),.clk(gclk));
	jand g1431(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1495),.clk(gclk));
	jnot g1432(.din(n1495),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_n1436_0[0]),.dinb(w_n1428_0[0]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1437_0[0]),.dinb(w_n1425_0[0]),.dout(n1498),.clk(gclk));
	jor g1435(.dina(n1498),.dinb(w_dff_B_S026EZg56_1),.dout(n1499),.clk(gclk));
	jand g1436(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1501),.clk(gclk));
	jor g1438(.dina(w_n1433_0[0]),.dinb(w_n1430_0[0]),.dout(n1502),.clk(gclk));
	jor g1439(.dina(w_n1435_0[0]),.dinb(w_n1429_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(n1503),.dinb(w_dff_B_zBIB7LIv3_1),.dout(n1504),.clk(gclk));
	jxor g1441(.dina(w_n1504_0[1]),.dinb(w_n1501_0[1]),.dout(n1505),.clk(gclk));
	jnot g1442(.din(n1505),.dout(n1506),.clk(gclk));
	jxor g1443(.dina(w_n1506_0[1]),.dinb(w_n1500_0[1]),.dout(n1507),.clk(gclk));
	jxor g1444(.dina(w_n1507_0[1]),.dinb(w_n1499_0[1]),.dout(n1508),.clk(gclk));
	jxor g1445(.dina(w_n1508_0[1]),.dinb(w_n1496_0[1]),.dout(n1509),.clk(gclk));
	jxor g1446(.dina(w_n1509_0[1]),.dinb(w_n1494_0[1]),.dout(n1510),.clk(gclk));
	jxor g1447(.dina(w_n1510_0[1]),.dinb(w_n1491_0[1]),.dout(n1511),.clk(gclk));
	jxor g1448(.dina(w_n1511_0[1]),.dinb(w_n1489_0[1]),.dout(n1512),.clk(gclk));
	jxor g1449(.dina(w_n1512_0[1]),.dinb(w_n1486_0[1]),.dout(n1513),.clk(gclk));
	jxor g1450(.dina(w_n1513_0[1]),.dinb(w_n1484_0[1]),.dout(n1514),.clk(gclk));
	jxor g1451(.dina(w_n1514_0[1]),.dinb(w_n1481_0[1]),.dout(n1515),.clk(gclk));
	jxor g1452(.dina(w_n1515_0[1]),.dinb(w_n1479_0[1]),.dout(n1516),.clk(gclk));
	jxor g1453(.dina(w_n1516_0[1]),.dinb(w_n1476_0[1]),.dout(n1517),.clk(gclk));
	jxor g1454(.dina(w_n1517_0[1]),.dinb(w_n1474_0[1]),.dout(n1518),.clk(gclk));
	jxor g1455(.dina(w_n1518_0[1]),.dinb(w_n1471_0[1]),.dout(n1519),.clk(gclk));
	jxor g1456(.dina(w_n1519_0[1]),.dinb(w_n1469_0[1]),.dout(n1520),.clk(gclk));
	jnot g1457(.din(n1520),.dout(n1521),.clk(gclk));
	jxor g1458(.dina(w_n1521_0[1]),.dinb(w_n1466_0[1]),.dout(n1522),.clk(gclk));
	jnot g1459(.din(n1522),.dout(n1523),.clk(gclk));
	jxor g1460(.dina(w_n1523_0[1]),.dinb(w_n1465_0[1]),.dout(n1524),.clk(gclk));
	jxor g1461(.dina(w_n1524_0[1]),.dinb(w_n1460_0[1]),.dout(w_dff_A_HN7yDTv85_2),.clk(gclk));
	jor g1462(.dina(w_n1523_0[0]),.dinb(w_n1465_0[0]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(w_n1524_0[0]),.dout(n1527),.clk(gclk));
	jor g1464(.dina(w_dff_B_NW2B2g9Z9_0),.dinb(w_n1460_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(n1528),.dinb(w_dff_B_la4C7ecR3_1),.dout(n1529),.clk(gclk));
	jnot g1466(.din(w_n1469_0[0]),.dout(n1530),.clk(gclk));
	jnot g1467(.din(w_n1519_0[0]),.dout(n1531),.clk(gclk));
	jor g1468(.dina(w_dff_B_xTRmInr30_0),.dinb(n1530),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1521_0[0]),.dinb(w_n1466_0[0]),.dout(n1533),.clk(gclk));
	jand g1470(.dina(n1533),.dinb(w_dff_B_QvWK9LdJ4_1),.dout(n1534),.clk(gclk));
	jand g1471(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1535),.clk(gclk));
	jand g1472(.dina(w_n1517_0[0]),.dinb(w_n1474_0[0]),.dout(n1536),.clk(gclk));
	jand g1473(.dina(w_n1518_0[0]),.dinb(w_n1471_0[0]),.dout(n1537),.clk(gclk));
	jor g1474(.dina(n1537),.dinb(w_dff_B_mEub8Cht3_1),.dout(n1538),.clk(gclk));
	jand g1475(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1539),.clk(gclk));
	jnot g1476(.din(n1539),.dout(n1540),.clk(gclk));
	jand g1477(.dina(w_n1515_0[0]),.dinb(w_n1479_0[0]),.dout(n1541),.clk(gclk));
	jand g1478(.dina(w_n1516_0[0]),.dinb(w_n1476_0[0]),.dout(n1542),.clk(gclk));
	jor g1479(.dina(n1542),.dinb(w_dff_B_nhG2MuVO0_1),.dout(n1543),.clk(gclk));
	jand g1480(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1544),.clk(gclk));
	jnot g1481(.din(n1544),.dout(n1545),.clk(gclk));
	jand g1482(.dina(w_n1513_0[0]),.dinb(w_n1484_0[0]),.dout(n1546),.clk(gclk));
	jand g1483(.dina(w_n1514_0[0]),.dinb(w_n1481_0[0]),.dout(n1547),.clk(gclk));
	jor g1484(.dina(n1547),.dinb(w_dff_B_rtoEWXzK4_1),.dout(n1548),.clk(gclk));
	jand g1485(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1549),.clk(gclk));
	jnot g1486(.din(n1549),.dout(n1550),.clk(gclk));
	jand g1487(.dina(w_n1511_0[0]),.dinb(w_n1489_0[0]),.dout(n1551),.clk(gclk));
	jand g1488(.dina(w_n1512_0[0]),.dinb(w_n1486_0[0]),.dout(n1552),.clk(gclk));
	jor g1489(.dina(n1552),.dinb(w_dff_B_kTo0wJwr9_1),.dout(n1553),.clk(gclk));
	jand g1490(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1554),.clk(gclk));
	jnot g1491(.din(n1554),.dout(n1555),.clk(gclk));
	jand g1492(.dina(w_n1509_0[0]),.dinb(w_n1494_0[0]),.dout(n1556),.clk(gclk));
	jand g1493(.dina(w_n1510_0[0]),.dinb(w_n1491_0[0]),.dout(n1557),.clk(gclk));
	jor g1494(.dina(n1557),.dinb(w_dff_B_iQ0mUJQH6_1),.dout(n1558),.clk(gclk));
	jand g1495(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1559),.clk(gclk));
	jnot g1496(.din(n1559),.dout(n1560),.clk(gclk));
	jand g1497(.dina(w_n1507_0[0]),.dinb(w_n1499_0[0]),.dout(n1561),.clk(gclk));
	jand g1498(.dina(w_n1508_0[0]),.dinb(w_n1496_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(n1562),.dinb(w_dff_B_plcpmFsX2_1),.dout(n1563),.clk(gclk));
	jand g1500(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1565),.clk(gclk));
	jor g1502(.dina(w_n1504_0[0]),.dinb(w_n1501_0[0]),.dout(n1566),.clk(gclk));
	jor g1503(.dina(w_n1506_0[0]),.dinb(w_n1500_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(n1567),.dinb(w_dff_B_R8uxWo708_1),.dout(n1568),.clk(gclk));
	jxor g1505(.dina(w_n1568_0[1]),.dinb(w_n1565_0[1]),.dout(n1569),.clk(gclk));
	jnot g1506(.din(n1569),.dout(n1570),.clk(gclk));
	jxor g1507(.dina(w_n1570_0[1]),.dinb(w_n1564_0[1]),.dout(n1571),.clk(gclk));
	jxor g1508(.dina(w_n1571_0[1]),.dinb(w_n1563_0[1]),.dout(n1572),.clk(gclk));
	jxor g1509(.dina(w_n1572_0[1]),.dinb(w_n1560_0[1]),.dout(n1573),.clk(gclk));
	jxor g1510(.dina(w_n1573_0[1]),.dinb(w_n1558_0[1]),.dout(n1574),.clk(gclk));
	jxor g1511(.dina(w_n1574_0[1]),.dinb(w_n1555_0[1]),.dout(n1575),.clk(gclk));
	jxor g1512(.dina(w_n1575_0[1]),.dinb(w_n1553_0[1]),.dout(n1576),.clk(gclk));
	jxor g1513(.dina(w_n1576_0[1]),.dinb(w_n1550_0[1]),.dout(n1577),.clk(gclk));
	jxor g1514(.dina(w_n1577_0[1]),.dinb(w_n1548_0[1]),.dout(n1578),.clk(gclk));
	jxor g1515(.dina(w_n1578_0[1]),.dinb(w_n1545_0[1]),.dout(n1579),.clk(gclk));
	jxor g1516(.dina(w_n1579_0[1]),.dinb(w_n1543_0[1]),.dout(n1580),.clk(gclk));
	jxor g1517(.dina(w_n1580_0[1]),.dinb(w_n1540_0[1]),.dout(n1581),.clk(gclk));
	jxor g1518(.dina(w_n1581_0[1]),.dinb(w_n1538_0[1]),.dout(n1582),.clk(gclk));
	jnot g1519(.din(n1582),.dout(n1583),.clk(gclk));
	jxor g1520(.dina(w_n1583_0[1]),.dinb(w_n1535_0[1]),.dout(n1584),.clk(gclk));
	jnot g1521(.din(n1584),.dout(n1585),.clk(gclk));
	jxor g1522(.dina(w_n1585_0[1]),.dinb(w_n1534_0[1]),.dout(n1586),.clk(gclk));
	jxor g1523(.dina(w_n1586_0[1]),.dinb(w_n1529_0[1]),.dout(w_dff_A_5arqhEZw5_2),.clk(gclk));
	jor g1524(.dina(w_n1585_0[0]),.dinb(w_n1534_0[0]),.dout(n1588),.clk(gclk));
	jnot g1525(.din(w_n1586_0[0]),.dout(n1589),.clk(gclk));
	jor g1526(.dina(w_dff_B_7MkU68A62_0),.dinb(w_n1529_0[0]),.dout(n1590),.clk(gclk));
	jand g1527(.dina(n1590),.dinb(w_dff_B_fPT3ph2e2_1),.dout(n1591),.clk(gclk));
	jnot g1528(.din(w_n1538_0[0]),.dout(n1592),.clk(gclk));
	jnot g1529(.din(w_n1581_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(w_dff_B_gnw9YzMm7_0),.dinb(n1592),.dout(n1594),.clk(gclk));
	jor g1531(.dina(w_n1583_0[0]),.dinb(w_n1535_0[0]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(n1595),.dinb(w_dff_B_tH64gZ2p2_1),.dout(n1596),.clk(gclk));
	jand g1533(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1597),.clk(gclk));
	jand g1534(.dina(w_n1579_0[0]),.dinb(w_n1543_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(w_n1580_0[0]),.dinb(w_n1540_0[0]),.dout(n1599),.clk(gclk));
	jor g1536(.dina(n1599),.dinb(w_dff_B_5fqpPpqw5_1),.dout(n1600),.clk(gclk));
	jand g1537(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1601),.clk(gclk));
	jnot g1538(.din(n1601),.dout(n1602),.clk(gclk));
	jand g1539(.dina(w_n1577_0[0]),.dinb(w_n1548_0[0]),.dout(n1603),.clk(gclk));
	jand g1540(.dina(w_n1578_0[0]),.dinb(w_n1545_0[0]),.dout(n1604),.clk(gclk));
	jor g1541(.dina(n1604),.dinb(w_dff_B_72FCd2WI3_1),.dout(n1605),.clk(gclk));
	jand g1542(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1606),.clk(gclk));
	jnot g1543(.din(n1606),.dout(n1607),.clk(gclk));
	jand g1544(.dina(w_n1575_0[0]),.dinb(w_n1553_0[0]),.dout(n1608),.clk(gclk));
	jand g1545(.dina(w_n1576_0[0]),.dinb(w_n1550_0[0]),.dout(n1609),.clk(gclk));
	jor g1546(.dina(n1609),.dinb(w_dff_B_EBXg5wWk4_1),.dout(n1610),.clk(gclk));
	jand g1547(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1611),.clk(gclk));
	jnot g1548(.din(n1611),.dout(n1612),.clk(gclk));
	jand g1549(.dina(w_n1573_0[0]),.dinb(w_n1558_0[0]),.dout(n1613),.clk(gclk));
	jand g1550(.dina(w_n1574_0[0]),.dinb(w_n1555_0[0]),.dout(n1614),.clk(gclk));
	jor g1551(.dina(n1614),.dinb(w_dff_B_QaZA6LOD3_1),.dout(n1615),.clk(gclk));
	jand g1552(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1616),.clk(gclk));
	jnot g1553(.din(n1616),.dout(n1617),.clk(gclk));
	jand g1554(.dina(w_n1571_0[0]),.dinb(w_n1563_0[0]),.dout(n1618),.clk(gclk));
	jand g1555(.dina(w_n1572_0[0]),.dinb(w_n1560_0[0]),.dout(n1619),.clk(gclk));
	jor g1556(.dina(n1619),.dinb(w_dff_B_HJZteJoN3_1),.dout(n1620),.clk(gclk));
	jand g1557(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1622),.clk(gclk));
	jor g1559(.dina(w_n1568_0[0]),.dinb(w_n1565_0[0]),.dout(n1623),.clk(gclk));
	jor g1560(.dina(w_n1570_0[0]),.dinb(w_n1564_0[0]),.dout(n1624),.clk(gclk));
	jand g1561(.dina(n1624),.dinb(w_dff_B_5qq234Sr4_1),.dout(n1625),.clk(gclk));
	jxor g1562(.dina(w_n1625_0[1]),.dinb(w_n1622_0[1]),.dout(n1626),.clk(gclk));
	jnot g1563(.din(n1626),.dout(n1627),.clk(gclk));
	jxor g1564(.dina(w_n1627_0[1]),.dinb(w_n1621_0[1]),.dout(n1628),.clk(gclk));
	jxor g1565(.dina(w_n1628_0[1]),.dinb(w_n1620_0[1]),.dout(n1629),.clk(gclk));
	jxor g1566(.dina(w_n1629_0[1]),.dinb(w_n1617_0[1]),.dout(n1630),.clk(gclk));
	jxor g1567(.dina(w_n1630_0[1]),.dinb(w_n1615_0[1]),.dout(n1631),.clk(gclk));
	jxor g1568(.dina(w_n1631_0[1]),.dinb(w_n1612_0[1]),.dout(n1632),.clk(gclk));
	jxor g1569(.dina(w_n1632_0[1]),.dinb(w_n1610_0[1]),.dout(n1633),.clk(gclk));
	jxor g1570(.dina(w_n1633_0[1]),.dinb(w_n1607_0[1]),.dout(n1634),.clk(gclk));
	jxor g1571(.dina(w_n1634_0[1]),.dinb(w_n1605_0[1]),.dout(n1635),.clk(gclk));
	jxor g1572(.dina(w_n1635_0[1]),.dinb(w_n1602_0[1]),.dout(n1636),.clk(gclk));
	jxor g1573(.dina(w_n1636_0[1]),.dinb(w_n1600_0[1]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jxor g1575(.dina(w_n1638_0[1]),.dinb(w_n1597_0[1]),.dout(n1639),.clk(gclk));
	jnot g1576(.din(n1639),.dout(n1640),.clk(gclk));
	jxor g1577(.dina(w_n1640_0[1]),.dinb(w_n1596_0[1]),.dout(n1641),.clk(gclk));
	jxor g1578(.dina(w_n1641_0[1]),.dinb(w_n1591_0[1]),.dout(w_dff_A_OWGNsutV7_2),.clk(gclk));
	jor g1579(.dina(w_n1640_0[0]),.dinb(w_n1596_0[0]),.dout(n1643),.clk(gclk));
	jnot g1580(.din(w_n1641_0[0]),.dout(n1644),.clk(gclk));
	jor g1581(.dina(w_dff_B_Dmfo7PaF5_0),.dinb(w_n1591_0[0]),.dout(n1645),.clk(gclk));
	jand g1582(.dina(n1645),.dinb(w_dff_B_Dr5rfgtG5_1),.dout(n1646),.clk(gclk));
	jnot g1583(.din(w_n1600_0[0]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(w_n1636_0[0]),.dout(n1648),.clk(gclk));
	jor g1585(.dina(n1648),.dinb(n1647),.dout(n1649),.clk(gclk));
	jor g1586(.dina(w_n1638_0[0]),.dinb(w_n1597_0[0]),.dout(n1650),.clk(gclk));
	jand g1587(.dina(n1650),.dinb(w_dff_B_8u82OTEk1_1),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1652),.clk(gclk));
	jnot g1589(.din(n1652),.dout(n1653),.clk(gclk));
	jand g1590(.dina(w_n1634_0[0]),.dinb(w_n1605_0[0]),.dout(n1654),.clk(gclk));
	jand g1591(.dina(w_n1635_0[0]),.dinb(w_n1602_0[0]),.dout(n1655),.clk(gclk));
	jor g1592(.dina(n1655),.dinb(w_dff_B_fL374ioq5_1),.dout(n1656),.clk(gclk));
	jand g1593(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jand g1595(.dina(w_n1632_0[0]),.dinb(w_n1610_0[0]),.dout(n1659),.clk(gclk));
	jand g1596(.dina(w_n1633_0[0]),.dinb(w_n1607_0[0]),.dout(n1660),.clk(gclk));
	jor g1597(.dina(n1660),.dinb(w_dff_B_eWtrvpIs8_1),.dout(n1661),.clk(gclk));
	jand g1598(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1662),.clk(gclk));
	jnot g1599(.din(n1662),.dout(n1663),.clk(gclk));
	jand g1600(.dina(w_n1630_0[0]),.dinb(w_n1615_0[0]),.dout(n1664),.clk(gclk));
	jand g1601(.dina(w_n1631_0[0]),.dinb(w_n1612_0[0]),.dout(n1665),.clk(gclk));
	jor g1602(.dina(n1665),.dinb(w_dff_B_2UH6Sju27_1),.dout(n1666),.clk(gclk));
	jand g1603(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1667),.clk(gclk));
	jnot g1604(.din(n1667),.dout(n1668),.clk(gclk));
	jand g1605(.dina(w_n1628_0[0]),.dinb(w_n1620_0[0]),.dout(n1669),.clk(gclk));
	jand g1606(.dina(w_n1629_0[0]),.dinb(w_n1617_0[0]),.dout(n1670),.clk(gclk));
	jor g1607(.dina(n1670),.dinb(w_dff_B_egK88UFU6_1),.dout(n1671),.clk(gclk));
	jand g1608(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1672),.clk(gclk));
	jand g1609(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1673),.clk(gclk));
	jor g1610(.dina(w_n1625_0[0]),.dinb(w_n1622_0[0]),.dout(n1674),.clk(gclk));
	jor g1611(.dina(w_n1627_0[0]),.dinb(w_n1621_0[0]),.dout(n1675),.clk(gclk));
	jand g1612(.dina(n1675),.dinb(w_dff_B_XGro1DDU8_1),.dout(n1676),.clk(gclk));
	jxor g1613(.dina(w_n1676_0[1]),.dinb(w_n1673_0[1]),.dout(n1677),.clk(gclk));
	jnot g1614(.din(n1677),.dout(n1678),.clk(gclk));
	jxor g1615(.dina(w_n1678_0[1]),.dinb(w_n1672_0[1]),.dout(n1679),.clk(gclk));
	jxor g1616(.dina(w_n1679_0[1]),.dinb(w_n1671_0[1]),.dout(n1680),.clk(gclk));
	jxor g1617(.dina(w_n1680_0[1]),.dinb(w_n1668_0[1]),.dout(n1681),.clk(gclk));
	jxor g1618(.dina(w_n1681_0[1]),.dinb(w_n1666_0[1]),.dout(n1682),.clk(gclk));
	jxor g1619(.dina(w_n1682_0[1]),.dinb(w_n1663_0[1]),.dout(n1683),.clk(gclk));
	jxor g1620(.dina(w_n1683_0[1]),.dinb(w_n1661_0[1]),.dout(n1684),.clk(gclk));
	jxor g1621(.dina(w_n1684_0[1]),.dinb(w_n1658_0[1]),.dout(n1685),.clk(gclk));
	jxor g1622(.dina(w_n1685_0[1]),.dinb(w_n1656_0[1]),.dout(n1686),.clk(gclk));
	jxor g1623(.dina(w_n1686_0[1]),.dinb(w_n1653_0[1]),.dout(n1687),.clk(gclk));
	jnot g1624(.din(n1687),.dout(n1688),.clk(gclk));
	jxor g1625(.dina(w_n1688_0[1]),.dinb(w_n1651_0[1]),.dout(n1689),.clk(gclk));
	jxor g1626(.dina(w_n1689_0[1]),.dinb(w_n1646_0[1]),.dout(w_dff_A_FgSjYYdM3_2),.clk(gclk));
	jor g1627(.dina(w_n1688_0[0]),.dinb(w_n1651_0[0]),.dout(n1691),.clk(gclk));
	jnot g1628(.din(w_n1689_0[0]),.dout(n1692),.clk(gclk));
	jor g1629(.dina(w_dff_B_OfOjkk3r2_0),.dinb(w_n1646_0[0]),.dout(n1693),.clk(gclk));
	jand g1630(.dina(n1693),.dinb(w_dff_B_BJyvovda8_1),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1685_0[0]),.dinb(w_n1656_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1686_0[0]),.dinb(w_n1653_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(w_dff_B_2BO5H3Fh3_1),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1683_0[0]),.dinb(w_n1661_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1684_0[0]),.dinb(w_n1658_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(w_dff_B_rhnCP9QY2_1),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1703),.clk(gclk));
	jnot g1640(.din(n1703),.dout(n1704),.clk(gclk));
	jand g1641(.dina(w_n1681_0[0]),.dinb(w_n1666_0[0]),.dout(n1705),.clk(gclk));
	jand g1642(.dina(w_n1682_0[0]),.dinb(w_n1663_0[0]),.dout(n1706),.clk(gclk));
	jor g1643(.dina(n1706),.dinb(w_dff_B_qIxe3vd75_1),.dout(n1707),.clk(gclk));
	jand g1644(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jand g1646(.dina(w_n1679_0[0]),.dinb(w_n1671_0[0]),.dout(n1710),.clk(gclk));
	jand g1647(.dina(w_n1680_0[0]),.dinb(w_n1668_0[0]),.dout(n1711),.clk(gclk));
	jor g1648(.dina(n1711),.dinb(w_dff_B_so3bvXCA9_1),.dout(n1712),.clk(gclk));
	jand g1649(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1713),.clk(gclk));
	jand g1650(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1714),.clk(gclk));
	jor g1651(.dina(w_n1676_0[0]),.dinb(w_n1673_0[0]),.dout(n1715),.clk(gclk));
	jor g1652(.dina(w_n1678_0[0]),.dinb(w_n1672_0[0]),.dout(n1716),.clk(gclk));
	jand g1653(.dina(n1716),.dinb(w_dff_B_dofnAvnv2_1),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1714_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1713_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1712_0[1]),.dout(n1721),.clk(gclk));
	jxor g1658(.dina(w_n1721_0[1]),.dinb(w_n1709_0[1]),.dout(n1722),.clk(gclk));
	jxor g1659(.dina(w_n1722_0[1]),.dinb(w_n1707_0[1]),.dout(n1723),.clk(gclk));
	jxor g1660(.dina(w_n1723_0[1]),.dinb(w_n1704_0[1]),.dout(n1724),.clk(gclk));
	jxor g1661(.dina(w_n1724_0[1]),.dinb(w_n1702_0[1]),.dout(n1725),.clk(gclk));
	jxor g1662(.dina(w_n1725_0[1]),.dinb(w_n1699_0[1]),.dout(n1726),.clk(gclk));
	jxor g1663(.dina(w_n1726_0[1]),.dinb(w_n1697_0[1]),.dout(n1727),.clk(gclk));
	jxor g1664(.dina(w_n1727_0[1]),.dinb(w_n1694_0[1]),.dout(w_dff_A_c6Fm6OCo3_2),.clk(gclk));
	jnot g1665(.din(w_n1697_0[0]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(w_n1726_0[0]),.dout(n1730),.clk(gclk));
	jor g1667(.dina(n1730),.dinb(w_dff_B_GwYof2122_1),.dout(n1731),.clk(gclk));
	jnot g1668(.din(w_n1727_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(w_dff_B_CZ6KcnlD1_0),.dinb(w_n1694_0[0]),.dout(n1733),.clk(gclk));
	jand g1670(.dina(n1733),.dinb(w_dff_B_gEpp6YSE9_1),.dout(n1734),.clk(gclk));
	jand g1671(.dina(w_n1724_0[0]),.dinb(w_n1702_0[0]),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1725_0[0]),.dinb(w_n1699_0[0]),.dout(n1736),.clk(gclk));
	jor g1673(.dina(n1736),.dinb(w_dff_B_iOR8SBie2_1),.dout(n1737),.clk(gclk));
	jand g1674(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1738),.clk(gclk));
	jnot g1675(.din(n1738),.dout(n1739),.clk(gclk));
	jand g1676(.dina(w_n1722_0[0]),.dinb(w_n1707_0[0]),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1723_0[0]),.dinb(w_n1704_0[0]),.dout(n1741),.clk(gclk));
	jor g1678(.dina(n1741),.dinb(w_dff_B_YZ2J9A3L8_1),.dout(n1742),.clk(gclk));
	jand g1679(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1743),.clk(gclk));
	jnot g1680(.din(n1743),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_n1720_0[0]),.dinb(w_n1712_0[0]),.dout(n1745),.clk(gclk));
	jand g1682(.dina(w_n1721_0[0]),.dinb(w_n1709_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(n1746),.dinb(w_dff_B_ntpkS7Lg8_1),.dout(n1747),.clk(gclk));
	jand g1684(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1748),.clk(gclk));
	jand g1685(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1749),.clk(gclk));
	jor g1686(.dina(w_n1717_0[0]),.dinb(w_n1714_0[0]),.dout(n1750),.clk(gclk));
	jor g1687(.dina(w_n1719_0[0]),.dinb(w_n1713_0[0]),.dout(n1751),.clk(gclk));
	jand g1688(.dina(n1751),.dinb(w_dff_B_HuYfgTST5_1),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1749_0[1]),.dout(n1753),.clk(gclk));
	jnot g1690(.din(n1753),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1748_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1747_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1744_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1742_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1739_0[1]),.dout(n1759),.clk(gclk));
	jxor g1696(.dina(w_n1759_0[1]),.dinb(w_n1737_0[1]),.dout(n1760),.clk(gclk));
	jxor g1697(.dina(w_n1760_0[1]),.dinb(w_n1734_0[1]),.dout(w_dff_A_cTXjgFSt7_2),.clk(gclk));
	jnot g1698(.din(w_n1737_0[0]),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1759_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(n1763),.dinb(w_dff_B_s9lPq6nu2_1),.dout(n1764),.clk(gclk));
	jnot g1701(.din(w_n1760_0[0]),.dout(n1765),.clk(gclk));
	jor g1702(.dina(w_dff_B_uwUQSseo9_0),.dinb(w_n1734_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(n1766),.dinb(w_dff_B_7RvKsDtP2_1),.dout(n1767),.clk(gclk));
	jand g1704(.dina(w_n1757_0[0]),.dinb(w_n1742_0[0]),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_n1758_0[0]),.dinb(w_n1739_0[0]),.dout(n1769),.clk(gclk));
	jor g1706(.dina(n1769),.dinb(w_dff_B_cNIx8qef4_1),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1771),.clk(gclk));
	jnot g1708(.din(n1771),.dout(n1772),.clk(gclk));
	jand g1709(.dina(w_n1755_0[0]),.dinb(w_n1747_0[0]),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_n1756_0[0]),.dinb(w_n1744_0[0]),.dout(n1774),.clk(gclk));
	jor g1711(.dina(n1774),.dinb(w_dff_B_w3zmnl6r0_1),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(w_n1752_0[0]),.dinb(w_n1749_0[0]),.dout(n1778),.clk(gclk));
	jor g1715(.dina(w_n1754_0[0]),.dinb(w_n1748_0[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(n1779),.dinb(w_dff_B_KInWw2Ze8_1),.dout(n1780),.clk(gclk));
	jxor g1717(.dina(w_n1780_0[1]),.dinb(w_n1777_0[1]),.dout(n1781),.clk(gclk));
	jnot g1718(.din(n1781),.dout(n1782),.clk(gclk));
	jxor g1719(.dina(w_n1782_0[1]),.dinb(w_n1776_0[1]),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1775_0[1]),.dout(n1784),.clk(gclk));
	jxor g1721(.dina(w_n1784_0[1]),.dinb(w_n1772_0[1]),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1770_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1767_0[1]),.dout(w_dff_A_MtaWg8ib7_2),.clk(gclk));
	jnot g1724(.din(w_n1770_0[0]),.dout(n1788),.clk(gclk));
	jnot g1725(.din(w_n1785_0[0]),.dout(n1789),.clk(gclk));
	jor g1726(.dina(n1789),.dinb(w_dff_B_IuxRMeHR7_1),.dout(n1790),.clk(gclk));
	jnot g1727(.din(w_n1786_0[0]),.dout(n1791),.clk(gclk));
	jor g1728(.dina(w_dff_B_ZeYPt54T0_0),.dinb(w_n1767_0[0]),.dout(n1792),.clk(gclk));
	jand g1729(.dina(n1792),.dinb(w_dff_B_yRWuqKkw5_1),.dout(n1793),.clk(gclk));
	jand g1730(.dina(w_n1783_0[0]),.dinb(w_n1775_0[0]),.dout(n1794),.clk(gclk));
	jand g1731(.dina(w_n1784_0[0]),.dinb(w_n1772_0[0]),.dout(n1795),.clk(gclk));
	jor g1732(.dina(n1795),.dinb(w_dff_B_kLCCYxg90_1),.dout(n1796),.clk(gclk));
	jand g1733(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1798),.clk(gclk));
	jor g1735(.dina(w_n1780_0[0]),.dinb(w_n1777_0[0]),.dout(n1799),.clk(gclk));
	jor g1736(.dina(w_n1782_0[0]),.dinb(w_n1776_0[0]),.dout(n1800),.clk(gclk));
	jand g1737(.dina(n1800),.dinb(w_dff_B_faZ3ZuPl5_1),.dout(n1801),.clk(gclk));
	jxor g1738(.dina(w_n1801_0[1]),.dinb(w_n1798_0[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jxor g1740(.dina(w_n1803_0[1]),.dinb(w_n1797_0[1]),.dout(n1804),.clk(gclk));
	jxor g1741(.dina(w_n1804_0[1]),.dinb(w_n1796_0[1]),.dout(n1805),.clk(gclk));
	jxor g1742(.dina(w_n1805_0[1]),.dinb(w_n1793_0[1]),.dout(w_dff_A_GvGhDXPx3_2),.clk(gclk));
	jand g1743(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1807),.clk(gclk));
	jor g1744(.dina(w_n1801_0[0]),.dinb(w_n1798_0[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1803_0[0]),.dinb(w_n1797_0[0]),.dout(n1809),.clk(gclk));
	jand g1746(.dina(n1809),.dinb(w_dff_B_JdEVAEq01_1),.dout(n1810),.clk(gclk));
	jor g1747(.dina(w_n1810_0[1]),.dinb(w_n1807_0[1]),.dout(n1811),.clk(gclk));
	jnot g1748(.din(w_n1796_0[0]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(w_n1804_0[0]),.dout(n1813),.clk(gclk));
	jor g1750(.dina(n1813),.dinb(w_dff_B_3khtPMZW2_1),.dout(n1814),.clk(gclk));
	jnot g1751(.din(w_n1805_0[0]),.dout(n1815),.clk(gclk));
	jor g1752(.dina(w_dff_B_uG0G052K0_0),.dinb(w_n1793_0[0]),.dout(n1816),.clk(gclk));
	jand g1753(.dina(n1816),.dinb(w_dff_B_rKvz3qNj9_1),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1810_0[0]),.dinb(w_n1807_0[0]),.dout(n1818),.clk(gclk));
	jnot g1755(.din(w_n1818_0[1]),.dout(n1819),.clk(gclk));
	jor g1756(.dina(w_dff_B_sQArDvcX8_0),.dinb(w_n1817_0[1]),.dout(n1820),.clk(gclk));
	jand g1757(.dina(n1820),.dinb(w_dff_B_huyM6Sbm7_1),.dout(G6287gat),.clk(gclk));
	jxor g1758(.dina(w_n1818_0[0]),.dinb(w_n1817_0[0]),.dout(w_dff_A_l6uLDiYR0_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl jspl_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl jspl_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_G307gat_2[1]),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl jspl_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_SBHDbXIx1_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n66_0(.douta(w_dff_A_eAFIM9nI2_0),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(w_dff_B_9Vf5Icva4_2));
	jspl jspl_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n75_0(.douta(w_dff_A_eQtCUR2S4_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n80_0(.douta(w_dff_A_iGsqUyTS8_0),.doutb(w_n80_0[1]),.doutc(w_n80_0[2]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_GHg8aXye0_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_dff_A_wyHhALjm2_0),.doutb(w_n91_0[1]),.din(n91));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_GQBtAAG96_1),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_dff_A_mRes1rl40_0),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl jspl_w_n112_0(.douta(w_dff_A_yz2g5o3T1_0),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(w_dff_B_O43b9nPM6_2));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n122_0(.douta(w_dff_A_VnVkTe6E1_0),.doutb(w_n122_0[1]),.din(n122));
	jspl jspl_w_n123_0(.douta(w_dff_A_uRE18QYz7_0),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n129_0(.douta(w_dff_A_OcGInJTO8_0),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n132_0(.douta(w_n132_0[0]),.doutb(w_dff_A_WxYnSB6O0_1),.din(n132));
	jspl jspl_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.din(n133));
	jspl jspl_w_n135_0(.douta(w_dff_A_vEHJDhK88_0),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_Ub9v0iXs2_0),.doutb(w_n141_0[1]),.din(n141));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.doutc(w_n146_0[2]),.din(n146));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(w_dff_B_NaR232Rg3_2));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(w_dff_B_qFMZlzBN6_2));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_dff_A_NFpSeRGc1_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_dff_A_0Gfv49f07_0),.doutb(w_n157_0[1]),.din(n157));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(n158));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl jspl_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(w_dff_B_Z5Otzmzb1_2));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n164_0(.douta(w_dff_A_uGHgRN7S4_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_RjMD47tF9_1),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl jspl_w_n170_0(.douta(w_dff_A_O45etuQo1_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n176_0(.douta(w_dff_A_Usx6TU591_0),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.din(w_dff_B_e4Sw9TXZ8_2));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(w_dff_B_Z7m1PGz53_2));
	jspl jspl_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.din(n192));
	jspl jspl_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.din(w_dff_B_cj34X8qx6_2));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_PJAIXXDw9_0),.doutb(w_dff_A_q9M9gnBA4_1),.doutc(w_n196_0[2]),.din(n196));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(w_dff_B_9pL1rP5c5_2));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(n203));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(w_dff_B_ezZqCDx86_2));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n206_0(.douta(w_dff_A_xTHqHmzl2_0),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_w1J36y282_1),.din(n209));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_dff_A_mzsbKJ0A0_0),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_dff_A_ZGD17F2e9_0),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.doutc(w_n223_0[2]),.din(n223));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(w_dff_B_4w5HXiWm6_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(w_dff_B_NoOfWuhP6_2));
	jspl jspl_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.din(n233));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.din(w_dff_B_MLy6fGzE4_2));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(w_dff_B_lTV9VUfa5_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_dff_A_OoN2Prmy8_0),.doutb(w_dff_A_U7KNUsVf3_1),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_NTfgZDis7_2));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.din(w_dff_B_uVj7vMka2_2));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(w_dff_B_tnSzTt9L3_2));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n255_0(.douta(w_dff_A_nhN25l222_0),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.din(n256));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_dff_A_mMzflZNv3_1),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_dff_A_MScdtDYV3_0),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_dff_A_07ryFYOn6_0),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.doutc(w_n272_0[2]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_DlfQu4jH3_2));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(w_dff_B_YuxiLJVP8_2));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(w_dff_B_vjmx9RdH1_2));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(w_dff_B_uIrpoRSt3_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_rXwee7iy7_2));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl3 jspl3_w_n297_0(.douta(w_dff_A_hmDCpiYY5_0),.doutb(w_dff_A_Cqil93OE8_1),.doutc(w_n297_0[2]),.din(n297));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl jspl_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.din(n301));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_n302_0[1]),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(w_dff_B_008ENNDH2_2));
	jspl jspl_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.din(n304));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(w_dff_B_waBKwR1N6_2));
	jspl jspl_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.din(n306));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(w_dff_B_FPWiNprk3_2));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(w_dff_B_jQbxvzmW2_2));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n311_0(.douta(w_dff_A_9FZh6byn6_0),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_dff_A_z1v3IO1U1_1),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_dff_A_k1BBpuyE8_0),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_dff_A_Y1PZdxHC4_0),.doutb(w_n323_0[1]),.din(n323));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(w_dff_B_ciueZflC7_2));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.din(w_dff_B_4GGfpT8Z2_2));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(w_dff_B_aXqrKbzR6_2));
	jspl jspl_w_n343_0(.douta(w_n343_0[0]),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(w_dff_B_bhrnvtsu1_2));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(w_dff_B_sUOIGnBS8_2));
	jspl jspl_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.din(n354));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(w_dff_B_XzIhFrPZ0_2));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n358_0(.douta(w_dff_A_ld5XHP2q6_0),.doutb(w_dff_A_iGOTVGdz2_1),.doutc(w_n358_0[2]),.din(n358));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(n363));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(w_dff_B_6texNomC5_2));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(w_dff_B_AZjjbSdA3_2));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(w_dff_B_wdsUzH4j4_2));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(w_dff_B_hUuxM9Cj6_2));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(w_dff_B_sqKLcQOC4_2));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n374_0(.douta(w_dff_A_pUfXEeqD8_0),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_Bovu7nZx1_1),.din(n377));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl jspl_w_n380_0(.douta(w_dff_A_mhHgcLc15_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_dff_A_9rwQQ0ko5_0),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(w_dff_B_TLAx6knM4_2));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl jspl_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.din(w_dff_B_0vg8Nkm94_2));
	jspl jspl_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.din(n401));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(w_dff_B_BS4fxE5g2_2));
	jspl jspl_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.din(n406));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(w_dff_B_4Ews6Nh30_2));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(n411));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(w_dff_B_LCG7Dk6n8_2));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(w_dff_B_JyHIx9uu1_2));
	jspl jspl_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.din(w_dff_B_a5JaWE737_2));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(w_dff_B_qT2GWI6i5_2));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl3 jspl3_w_n427_0(.douta(w_dff_A_tI7GeNyK3_0),.doutb(w_dff_A_4MM8phz66_1),.doutc(w_n427_0[2]),.din(n427));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl jspl_w_n431_0(.douta(w_n431_0[0]),.doutb(w_n431_0[1]),.din(n431));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(n432));
	jspl jspl_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.din(w_dff_B_Baav93bQ4_2));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(w_dff_B_r0V17XPo8_2));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(w_dff_B_a3vhh17j0_2));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(w_dff_B_1M3mdTob1_2));
	jspl jspl_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.din(n444));
	jspl jspl_w_n445_0(.douta(w_dff_A_WZktrhNT6_0),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_dff_A_RSzIhc3H1_1),.din(n448));
	jspl jspl_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.din(n449));
	jspl jspl_w_n451_0(.douta(w_dff_A_ERRIE9kX2_0),.doutb(w_n451_0[1]),.din(n451));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_dff_A_ufPHR4DL3_0),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(w_dff_B_q57hWTjr9_2));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(w_dff_B_1obje77m9_2));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(w_dff_B_4CxapzYz1_2));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(w_dff_B_JfRbc5xr0_2));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_jEXVVydu5_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_YFOUAA3M5_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_enx57Ify0_2));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.din(w_dff_B_7ZZLxOsm6_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl3 jspl3_w_n503_0(.douta(w_dff_A_rWc83jMO0_0),.doutb(w_dff_A_mOLit72c0_1),.doutc(w_n503_0[2]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_HmdH1K3B2_2));
	jspl jspl_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(w_dff_B_H0YJAthz5_2));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.din(n515));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(w_dff_B_4qBsAPLP7_2));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(w_dff_B_yR9CiLXM5_2));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.din(w_dff_B_0xyfVBWM7_2));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl jspl_w_n523_0(.douta(w_dff_A_ZUZuYvs31_0),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n526_0(.douta(w_n526_0[0]),.doutb(w_dff_A_kiwmOoXQ4_1),.din(n526));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_dff_A_bu9jZuxo2_0),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_dff_A_fuaXEbQU2_0),.doutb(w_n535_0[1]),.din(n535));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_SabJs8jz7_2));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(w_dff_B_uGOp2fnT2_2));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(w_dff_B_EPOCiutL4_2));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(w_dff_B_ImxTX2uV5_2));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(w_dff_B_uF078E1D9_2));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(w_dff_B_3uAKOUMy2_2));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(w_dff_B_hpCVcopu1_2));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(w_dff_B_SF8nTlbT9_2));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(w_dff_B_ts3WuSzZ2_2));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n586_0(.douta(w_dff_A_Y85roqRL0_0),.doutb(w_dff_A_as2XVWPH6_1),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(n588));
	jspl jspl_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.din(n590));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(w_dff_B_7qNLUpmv4_2));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.din(w_dff_B_N8xVdQVc1_2));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(w_dff_B_aW03qvsr3_2));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(w_dff_B_EnMmaieR2_2));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(w_dff_B_m8OWrTci8_2));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(w_dff_B_hR5poCbV0_2));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_dff_A_tK0LOVYt9_0),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n611_0(.douta(w_n611_0[0]),.doutb(w_dff_A_tWZbizCL0_1),.din(n611));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl jspl_w_n614_0(.douta(w_dff_A_QDiMJm2D6_0),.doutb(w_n614_0[1]),.din(n614));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_dff_A_z3WtrQqV4_0),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(w_dff_B_QaEcDSuD5_2));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(w_dff_B_SVn0Kq5S2_2));
	jspl jspl_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(w_dff_B_5DMS3Dqa4_2));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(w_dff_B_N8U5UmxG3_2));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(w_dff_B_XIqTUG0R2_2));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_uqRp0sXY8_2));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(w_dff_B_ZD8FogMh6_2));
	jspl jspl_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.din(n660));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(w_dff_B_RmOrkIc96_2));
	jspl jspl_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.din(n665));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(w_dff_B_KiS2yLUk1_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_3QPnI6HQ7_2));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl3 jspl3_w_n676_0(.douta(w_dff_A_sb8ifWuf6_0),.doutb(w_dff_A_YptSCDAG8_1),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(w_dff_B_BJLQn1AZ7_2));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(w_dff_B_6vOacekQ0_2));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(w_dff_B_YZpFnkvY4_2));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n688_0(.douta(w_n688_0[0]),.doutb(w_n688_0[1]),.din(w_dff_B_dnBmfhxP0_2));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.din(w_dff_B_cHYOWHXB5_2));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(w_dff_B_QMXPycXa7_2));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(w_dff_B_TJA2DPQ43_2));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n700_0(.douta(w_dff_A_UaJP31Zr4_0),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_iUY45Q7M8_1),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n706_0(.douta(w_dff_A_Evzuf2IR8_0),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_dff_A_4Ww2YHwk1_0),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.doutc(w_n717_0[2]),.din(n717));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(w_dff_B_48MqtL2S3_2));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(w_dff_B_dn6khCWy1_2));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(w_dff_B_uISdzOLI9_2));
	jspl jspl_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.din(n732));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(w_dff_B_QgQgfMTD9_2));
	jspl jspl_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.din(n737));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(w_dff_B_IUpPIGVx7_2));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl jspl_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.din(w_dff_B_QJ1fA5oe5_2));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(w_dff_B_XlNQGqbr8_2));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(w_dff_B_VRnjLZMF3_2));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(w_dff_B_L4nzzlCr2_2));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(w_dff_B_GURg5o5w9_2));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(w_dff_B_BUBibZu93_2));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(w_dff_B_9WGQxfkY6_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(w_dff_B_t4bNrN1L3_2));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.din(w_dff_B_1GKvZS0y0_2));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(w_dff_B_5kYk2Ixa5_2));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_OBfPOlGw5_2));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl jspl_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.din(n789));
	jspl jspl_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.din(n790));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl jspl_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.din(w_dff_B_xUzkRPVC2_2));
	jspl jspl_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.din(n794));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(w_dff_B_kQ3pLChE1_2));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(w_dff_B_Ch8v8ZGe5_2));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl jspl_w_n799_0(.douta(w_dff_A_CozEEMQj4_0),.doutb(w_n799_0[1]),.din(n799));
	jspl jspl_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_dff_A_8ocpneNJ7_1),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(n803));
	jspl jspl_w_n805_0(.douta(w_dff_A_fOMSH2Sk7_0),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(w_dff_B_hfAiVJWe3_2));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_dff_A_4lszyFn33_0),.doutb(w_n816_0[1]),.din(n816));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(w_dff_B_6PAvUIMV1_2));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(w_dff_B_l0x3636S9_2));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(w_dff_B_oweQ0Jal5_2));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(w_dff_B_5ffPzOR82_2));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(w_dff_B_Jyz2QApv5_2));
	jspl jspl_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.din(n845));
	jspl jspl_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.din(w_dff_B_nKiBMnI58_2));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(w_dff_B_QFBFxzKh3_2));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(w_dff_B_y521lsx49_2));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(w_dff_B_lEt3Fjqo3_2));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(w_dff_B_wSpih1Qt8_2));
	jspl jspl_w_n872_0(.douta(w_n872_0[0]),.doutb(w_n872_0[1]),.din(n872));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(w_dff_B_6xdhJ48v5_2));
	jspl jspl_w_n875_0(.douta(w_dff_A_ZGZ8rWrU5_0),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n877_0(.douta(w_dff_A_kM3WLGk62_0),.doutb(w_n877_0[1]),.din(w_dff_B_4DEEQ4gN5_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(w_dff_B_aL4m3DRC6_2));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.din(w_dff_B_Vd6fMmaD0_2));
	jspl jspl_w_n883_0(.douta(w_n883_0[0]),.doutb(w_n883_0[1]),.din(n883));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(w_dff_B_nNHk4TPi9_2));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(w_dff_B_FYrpa1pl8_2));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl jspl_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.din(w_dff_B_OuUO3ksH5_2));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(w_dff_B_JBIaOyn81_2));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(w_dff_B_8D3wYtpI7_2));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(w_dff_B_2oTC1IeI8_2));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.din(n899));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_dff_A_PaeTrKK39_1),.doutc(w_dff_A_1ezDC40J1_2),.din(n900));
	jspl jspl_w_n902_0(.douta(w_n902_0[0]),.doutb(w_dff_A_5cOfMQR71_1),.din(n902));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_dff_A_ra8b89sL4_1),.din(n904));
	jspl jspl_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.din(n905));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(w_dff_B_5PjTactY9_2));
	jspl3 jspl3_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.doutc(w_n915_0[2]),.din(n915));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(w_dff_B_h1Ll7FdX5_2));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(w_dff_B_TERMiXSN4_2));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(w_dff_B_uKmEUj662_2));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n934_0(.douta(w_n934_0[0]),.doutb(w_n934_0[1]),.din(w_dff_B_pOWat9C22_2));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(w_dff_B_VDExURbU0_2));
	jspl jspl_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.din(n942));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(w_dff_B_lZ5Qjorr3_2));
	jspl jspl_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.din(n947));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(w_dff_B_AJ278F735_2));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(w_dff_B_f5N2DkNH4_2));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(w_dff_B_vel3G9qh4_2));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(w_dff_B_0qnDpiRu7_2));
	jspl jspl_w_n967_0(.douta(w_n967_0[0]),.doutb(w_n967_0[1]),.din(n967));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(w_dff_B_imKGIIwC7_2));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(w_dff_B_rHluWfOf0_2));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl jspl_w_n980_0(.douta(w_dff_A_CQ0L2kB03_0),.doutb(w_n980_0[1]),.din(w_dff_B_pWjCZ7xu6_2));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.din(w_dff_B_lQTeKuBM6_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(w_dff_B_uSkMMjTT2_2));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_NGWTcjpH5_2));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(w_dff_B_8aMSco662_2));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(w_dff_B_BygthE7M4_2));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(w_dff_B_D286X2Hh9_2));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(w_dff_B_6UGA7hQZ1_2));
	jspl jspl_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.din(n995));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(w_dff_B_bcP0E7Hi5_2));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(w_dff_B_ZU10pe9H4_2));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.din(w_dff_B_0s0TzxQu7_2));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_hK4FPsXJ4_1),.din(n1006));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_dff_A_2JoOJDSK2_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(w_dff_B_T4lBY7sl2_2));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_dff_A_0ILHXRq21_1),.din(n1013));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(w_dff_B_SYqhYXJy0_2));
	jspl jspl_w_n1022_0(.douta(w_dff_A_pjjutMCB9_0),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(w_dff_B_73M7BQO13_2));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(w_dff_B_yxORPfpV4_2));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(w_dff_B_bJ48C7vN1_2));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.din(w_dff_B_UImGPrEg1_2));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(w_dff_B_wqQfrI6j6_2));
	jspl jspl_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.din(n1046));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(w_dff_B_NgZUA2VO6_2));
	jspl jspl_w_n1051_0(.douta(w_n1051_0[0]),.doutb(w_n1051_0[1]),.din(n1051));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(w_dff_B_tSTxillR3_2));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1058_0(.douta(w_n1058_0[0]),.doutb(w_n1058_0[1]),.din(w_dff_B_652yf0Nx1_2));
	jspl jspl_w_n1061_0(.douta(w_n1061_0[0]),.doutb(w_n1061_0[1]),.din(n1061));
	jspl jspl_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.din(w_dff_B_7weLBBiR8_2));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(w_dff_B_Ci9wtgQJ5_2));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(w_dff_B_dsSb6e5W5_2));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(w_dff_B_nWASdzTi0_2));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(w_dff_B_PJgaHfRU1_2));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(w_dff_B_gbsWdu792_2));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(n1084));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(w_dff_B_smVEtmv42_2));
	jspl jspl_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.din(n1086));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(w_dff_B_3TVnsZem2_2));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(w_dff_B_NeEOwLOI0_2));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(w_dff_B_hTlA5sbm7_2));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(w_dff_B_a8DfgMyJ2_2));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(w_dff_B_xho3upNn0_2));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1098_0(.douta(w_n1098_0[0]),.doutb(w_n1098_0[1]),.din(n1098));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.din(n1100));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(w_dff_B_kFtO13Jo8_2));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(w_dff_B_falzzeP72_2));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_n1106_0[1]),.din(n1106));
	jspl jspl_w_n1107_0(.douta(w_n1107_0[0]),.doutb(w_n1107_0[1]),.din(n1107));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_dff_A_ezmFXke16_1),.din(n1108));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1119_0(.douta(w_dff_A_kHDRHVTJ0_0),.doutb(w_n1119_0[1]),.din(w_dff_B_cMjIhJEV7_2));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(w_dff_B_wGGF3adj5_2));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(w_dff_B_b70qJSYz4_2));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(w_dff_B_K4Sn2Y1Z6_2));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_n1136_0[1]),.din(w_dff_B_2vJ0ECc04_2));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(w_dff_B_4HCmCGDr6_2));
	jspl jspl_w_n1144_0(.douta(w_n1144_0[0]),.doutb(w_n1144_0[1]),.din(n1144));
	jspl jspl_w_n1146_0(.douta(w_n1146_0[0]),.doutb(w_n1146_0[1]),.din(w_dff_B_95Ba9HeD1_2));
	jspl jspl_w_n1149_0(.douta(w_n1149_0[0]),.doutb(w_n1149_0[1]),.din(n1149));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(w_dff_B_JryGpri68_2));
	jspl jspl_w_n1154_0(.douta(w_n1154_0[0]),.doutb(w_n1154_0[1]),.din(n1154));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(w_dff_B_mNza9tcW4_2));
	jspl jspl_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(w_dff_B_sx23HeQZ2_2));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(w_dff_B_n2dKzKE83_2));
	jspl jspl_w_n1169_0(.douta(w_n1169_0[0]),.doutb(w_n1169_0[1]),.din(n1169));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(w_dff_B_DnRcI9J06_2));
	jspl jspl_w_n1174_0(.douta(w_n1174_0[0]),.doutb(w_n1174_0[1]),.din(n1174));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(w_dff_B_VjTNHORE0_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(w_dff_B_0k8pGfeg4_2));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1182_0(.douta(w_n1182_0[0]),.doutb(w_n1182_0[1]),.din(w_dff_B_OJa5jAA83_2));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(w_dff_B_I90VvDvk6_2));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(w_dff_B_aZm2xLBW4_2));
	jspl jspl_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.din(n1187));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(w_dff_B_WUYVu1hl2_2));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(w_dff_B_Plxwei5y9_2));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1192_0(.douta(w_n1192_0[0]),.doutb(w_n1192_0[1]),.din(w_dff_B_Hv6YVCsr6_2));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl jspl_w_n1194_0(.douta(w_n1194_0[0]),.doutb(w_n1194_0[1]),.din(w_dff_B_xjUxkvVQ5_2));
	jspl jspl_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.din(n1195));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.din(n1197));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl jspl_w_n1199_0(.douta(w_n1199_0[0]),.doutb(w_n1199_0[1]),.din(n1199));
	jspl jspl_w_n1200_0(.douta(w_n1200_0[0]),.doutb(w_n1200_0[1]),.din(w_dff_B_5iKIACOp3_2));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(w_dff_B_cdwtbpXo2_2));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(n1206));
	jspl jspl_w_n1207_0(.douta(w_dff_A_PYphhLrQ4_0),.doutb(w_n1207_0[1]),.din(n1207));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(w_dff_B_lMmJApGb6_2));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(w_dff_B_kISjt9Nd0_2));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(w_dff_B_yriLKFxM6_2));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(w_dff_B_1dOlMKis6_2));
	jspl jspl_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.din(n1235));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(w_dff_B_yeqhcbgU8_2));
	jspl jspl_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.din(n1240));
	jspl jspl_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.din(w_dff_B_BJnENFj11_2));
	jspl jspl_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.din(n1245));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(w_dff_B_lI9bCXDS3_2));
	jspl jspl_w_n1250_0(.douta(w_n1250_0[0]),.doutb(w_n1250_0[1]),.din(n1250));
	jspl jspl_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.din(w_dff_B_mIQobraJ3_2));
	jspl jspl_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.din(n1255));
	jspl jspl_w_n1257_0(.douta(w_n1257_0[0]),.doutb(w_n1257_0[1]),.din(w_dff_B_f1fCDRhk4_2));
	jspl jspl_w_n1260_0(.douta(w_n1260_0[0]),.doutb(w_n1260_0[1]),.din(n1260));
	jspl jspl_w_n1262_0(.douta(w_n1262_0[0]),.doutb(w_n1262_0[1]),.din(w_dff_B_YDaxvvi08_2));
	jspl jspl_w_n1265_0(.douta(w_n1265_0[0]),.doutb(w_n1265_0[1]),.din(n1265));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(w_dff_B_BP1LWsrF9_2));
	jspl jspl_w_n1267_0(.douta(w_n1267_0[0]),.doutb(w_n1267_0[1]),.din(w_dff_B_HYsBGq0B0_2));
	jspl jspl_w_n1270_0(.douta(w_n1270_0[0]),.doutb(w_n1270_0[1]),.din(n1270));
	jspl jspl_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.din(n1272));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(w_dff_B_PgfjzkDW5_2));
	jspl jspl_w_n1274_0(.douta(w_n1274_0[0]),.doutb(w_n1274_0[1]),.din(n1274));
	jspl jspl_w_n1275_0(.douta(w_n1275_0[0]),.doutb(w_n1275_0[1]),.din(w_dff_B_Xe6He2ej0_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1277_0(.douta(w_n1277_0[0]),.doutb(w_n1277_0[1]),.din(w_dff_B_FU4KmCfZ3_2));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(n1278));
	jspl jspl_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.din(w_dff_B_vcCq38sD8_2));
	jspl jspl_w_n1280_0(.douta(w_n1280_0[0]),.doutb(w_n1280_0[1]),.din(n1280));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(w_dff_B_iPNammup2_2));
	jspl jspl_w_n1282_0(.douta(w_n1282_0[0]),.doutb(w_n1282_0[1]),.din(n1282));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(w_dff_B_rRpQxRXk6_2));
	jspl jspl_w_n1284_0(.douta(w_n1284_0[0]),.doutb(w_n1284_0[1]),.din(n1284));
	jspl jspl_w_n1285_0(.douta(w_n1285_0[0]),.doutb(w_n1285_0[1]),.din(w_dff_B_Jne99qpP9_2));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1287_0(.douta(w_n1287_0[0]),.doutb(w_n1287_0[1]),.din(n1287));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1289_0(.douta(w_n1289_0[0]),.doutb(w_n1289_0[1]),.din(n1289));
	jspl jspl_w_n1290_0(.douta(w_n1290_0[0]),.doutb(w_n1290_0[1]),.din(n1290));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_dff_A_KSJU7kjs1_1),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(n1293));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_dff_A_2JNqYLSr2_1),.din(n1294));
	jspl jspl_w_n1295_0(.douta(w_dff_A_HSElSoIF5_0),.doutb(w_n1295_0[1]),.din(n1295));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(w_dff_B_RRUhEdFG0_2));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(w_dff_B_46wlq6IK4_2));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(w_dff_B_tUH2K1Kj7_2));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(w_dff_B_sJDrkbVR3_2));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1327_0(.douta(w_n1327_0[0]),.doutb(w_n1327_0[1]),.din(w_dff_B_FQxKZDL89_2));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(w_dff_B_FIqkKil95_2));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(w_dff_B_59Rap77Z8_2));
	jspl jspl_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.din(n1340));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(w_dff_B_QDSLTbY30_2));
	jspl jspl_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.din(n1345));
	jspl jspl_w_n1347_0(.douta(w_n1347_0[0]),.doutb(w_n1347_0[1]),.din(w_dff_B_9qLTKO0M8_2));
	jspl jspl_w_n1350_0(.douta(w_n1350_0[0]),.doutb(w_n1350_0[1]),.din(n1350));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(w_dff_B_5rhA6zGm7_2));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(w_dff_B_6BAj7eS14_2));
	jspl jspl_w_n1355_0(.douta(w_n1355_0[0]),.doutb(w_n1355_0[1]),.din(n1355));
	jspl jspl_w_n1357_0(.douta(w_n1357_0[0]),.doutb(w_n1357_0[1]),.din(n1357));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.din(w_dff_B_HCQgwVJi0_2));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(w_dff_B_8SaeRHr09_2));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(w_dff_B_QCqWFUuj5_2));
	jspl jspl_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.din(n1365));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(w_dff_B_Iax4cSnN7_2));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(w_dff_B_IP2xz7gk6_2));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_n1370_0[1]),.din(w_dff_B_lcTOel7j3_2));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(n1373));
	jspl jspl_w_n1374_0(.douta(w_n1374_0[0]),.doutb(w_n1374_0[1]),.din(n1374));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(n1378));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_dff_A_eCoR4Xyq0_1),.din(n1379));
	jspl jspl_w_n1384_0(.douta(w_n1384_0[0]),.doutb(w_n1384_0[1]),.din(n1384));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(w_dff_B_82kEDmpO3_2));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(w_dff_B_Jayjf1Sp4_2));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(w_dff_B_sDfgSwXx5_2));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(w_dff_B_i3Ve0M2d3_2));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(w_dff_B_S6AkPJPj3_2));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_n1408_0[1]),.din(n1408));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(w_dff_B_b6jgOv2c9_2));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(n1413));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(w_dff_B_SaWBszGf8_2));
	jspl jspl_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.din(n1418));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_1BL8Ahqj1_2));
	jspl jspl_w_n1423_0(.douta(w_n1423_0[0]),.doutb(w_n1423_0[1]),.din(n1423));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(w_dff_B_uNJ5Rqbx3_2));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(w_dff_B_q8jcn1tp2_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(w_dff_B_oHPukJZ31_2));
	jspl jspl_w_n1430_0(.douta(w_n1430_0[0]),.doutb(w_n1430_0[1]),.din(w_dff_B_KO8C55j57_2));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl jspl_w_n1437_0(.douta(w_n1437_0[0]),.doutb(w_n1437_0[1]),.din(n1437));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_n1438_0[1]),.din(n1438));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(w_dff_B_DMjZiILv3_2));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.din(w_dff_B_OMXvXjla2_2));
	jspl jspl_w_n1443_0(.douta(w_n1443_0[0]),.doutb(w_n1443_0[1]),.din(n1443));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(w_dff_B_YJTAuJ945_2));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(w_dff_B_389B8GSI6_2));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1448_0(.douta(w_n1448_0[0]),.doutb(w_n1448_0[1]),.din(w_dff_B_OeZSAjlN6_2));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(n1449));
	jspl jspl_w_n1450_0(.douta(w_n1450_0[0]),.doutb(w_n1450_0[1]),.din(n1450));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl jspl_w_n1455_0(.douta(w_n1455_0[0]),.doutb(w_dff_A_vTJCgUqr5_1),.din(n1455));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(n1460));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(w_dff_B_w8ZEJdi97_2));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(w_dff_B_bG14cOkU1_2));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(w_dff_B_q3UgyzgI7_2));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(w_dff_B_azQbmOOL5_2));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(w_dff_B_YklFauZj3_2));
	jspl jspl_w_n1484_0(.douta(w_n1484_0[0]),.doutb(w_n1484_0[1]),.din(n1484));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(w_dff_B_6ZFVxRWY6_2));
	jspl jspl_w_n1489_0(.douta(w_n1489_0[0]),.doutb(w_n1489_0[1]),.din(n1489));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(w_dff_B_qrmTfwrb9_2));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(w_dff_B_KkbJhSEQ3_2));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_B2JJaT8Y1_2));
	jspl jspl_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.din(w_dff_B_8HqNMCiP7_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(w_dff_B_2BeACS201_2));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_n1501_0[1]),.din(w_dff_B_7pxHhch97_2));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(n1507));
	jspl jspl_w_n1508_0(.douta(w_n1508_0[0]),.doutb(w_n1508_0[1]),.din(n1508));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1511_0(.douta(w_n1511_0[0]),.doutb(w_n1511_0[1]),.din(n1511));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(n1512));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(w_dff_B_p7AWjSaB0_2));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(w_dff_B_BHERS2qa9_2));
	jspl jspl_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.din(n1516));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(w_dff_B_LidCqk3d7_2));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1519_0(.douta(w_n1519_0[0]),.doutb(w_dff_A_Z1NK3AwW0_1),.din(n1519));
	jspl jspl_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.din(n1521));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl jspl_w_n1524_0(.douta(w_n1524_0[0]),.doutb(w_dff_A_G45fXfk25_1),.din(n1524));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(w_dff_B_ERHUrecI3_2));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(w_dff_B_KK9cnNdY5_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(w_dff_B_T9xSZq4u2_2));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(w_dff_B_Qs83rpz59_2));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_g95BrBah1_2));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(w_dff_B_8XvW1uyN8_2));
	jspl jspl_w_n1558_0(.douta(w_n1558_0[0]),.doutb(w_n1558_0[1]),.din(w_dff_B_mKfxyogV8_2));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(w_dff_B_vCWHOO814_2));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(w_dff_B_ipKRWSpy6_2));
	jspl jspl_w_n1564_0(.douta(w_n1564_0[0]),.doutb(w_n1564_0[1]),.din(w_dff_B_VtqpH4MQ5_2));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(w_dff_B_00H811zv5_2));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_n1568_0[1]),.din(n1568));
	jspl jspl_w_n1570_0(.douta(w_n1570_0[0]),.doutb(w_n1570_0[1]),.din(n1570));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1572_0(.douta(w_n1572_0[0]),.doutb(w_n1572_0[1]),.din(n1572));
	jspl jspl_w_n1573_0(.douta(w_n1573_0[0]),.doutb(w_n1573_0[1]),.din(n1573));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(n1576));
	jspl jspl_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.din(n1577));
	jspl jspl_w_n1578_0(.douta(w_n1578_0[0]),.doutb(w_n1578_0[1]),.din(n1578));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(w_dff_B_qGDh7Zs29_2));
	jspl jspl_w_n1580_0(.douta(w_n1580_0[0]),.doutb(w_n1580_0[1]),.din(n1580));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_dff_A_0VYyg8st6_1),.din(n1581));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl jspl_w_n1585_0(.douta(w_n1585_0[0]),.doutb(w_n1585_0[1]),.din(n1585));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_dff_A_xuraak5w1_1),.din(n1586));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(w_dff_B_r2TRi9Mw7_2));
	jspl jspl_w_n1600_0(.douta(w_n1600_0[0]),.doutb(w_n1600_0[1]),.din(n1600));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(w_dff_B_7sCSoUGO2_2));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(w_dff_B_JeVevLGF2_2));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(w_dff_B_KFTi04Gr6_2));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(w_dff_B_lTDcgB0E7_2));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(w_dff_B_g4sqGszj0_2));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(w_dff_B_YuhbQnDV1_2));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_n1617_0[1]),.din(w_dff_B_MoL9CwpP0_2));
	jspl jspl_w_n1620_0(.douta(w_n1620_0[0]),.doutb(w_n1620_0[1]),.din(w_dff_B_S9b9GWiV5_2));
	jspl jspl_w_n1621_0(.douta(w_n1621_0[0]),.doutb(w_n1621_0[1]),.din(w_dff_B_UxFdy8pr2_2));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(w_dff_B_3fu1YQq02_2));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(n1628));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1630_0(.douta(w_n1630_0[0]),.doutb(w_n1630_0[1]),.din(n1630));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1632_0(.douta(w_n1632_0[0]),.doutb(w_n1632_0[1]),.din(n1632));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(n1634));
	jspl jspl_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.din(n1635));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(n1636));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(n1638));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_dff_A_0iecNvAh2_1),.din(n1641));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(n1646));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_H4YrT5Qg7_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_nBxfy3Zo3_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(w_dff_B_toABSUla3_2));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(w_dff_B_x0b2LiBp2_2));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(w_dff_B_oh5mULbq1_2));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(w_dff_B_QBDy5FYn6_2));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(w_dff_B_uQ6Ji3YS2_2));
	jspl jspl_w_n1668_0(.douta(w_n1668_0[0]),.doutb(w_n1668_0[1]),.din(w_dff_B_YSlYmL2F6_2));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(w_dff_B_GhTEZuUV2_2));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(w_dff_B_SKoI0v3m4_2));
	jspl jspl_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.din(w_dff_B_nLDF5s0E1_2));
	jspl jspl_w_n1676_0(.douta(w_n1676_0[0]),.doutb(w_n1676_0[1]),.din(n1676));
	jspl jspl_w_n1678_0(.douta(w_n1678_0[0]),.doutb(w_n1678_0[1]),.din(n1678));
	jspl jspl_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1681_0(.douta(w_n1681_0[0]),.doutb(w_n1681_0[1]),.din(n1681));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl jspl_w_n1683_0(.douta(w_n1683_0[0]),.doutb(w_n1683_0[1]),.din(n1683));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(n1684));
	jspl jspl_w_n1685_0(.douta(w_n1685_0[0]),.doutb(w_n1685_0[1]),.din(n1685));
	jspl jspl_w_n1686_0(.douta(w_n1686_0[0]),.doutb(w_n1686_0[1]),.din(n1686));
	jspl jspl_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.din(n1688));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_dff_A_tcFSoMZz5_1),.din(n1689));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(n1694));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_dff_A_SwQ6ri8m3_1),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_4Kjf9Xzu5_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_AUJVVuZs7_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_R2b2iea10_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(w_dff_B_9JNkZehn3_2));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(w_dff_B_hc8D6Meq7_2));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(w_dff_B_fSAmthdF5_2));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(w_dff_B_Iwu0JBoY1_2));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(w_dff_B_qvorlkVc9_2));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1721_0(.douta(w_n1721_0[0]),.doutb(w_n1721_0[1]),.din(n1721));
	jspl jspl_w_n1722_0(.douta(w_n1722_0[0]),.doutb(w_n1722_0[1]),.din(n1722));
	jspl jspl_w_n1723_0(.douta(w_n1723_0[0]),.doutb(w_n1723_0[1]),.din(n1723));
	jspl jspl_w_n1724_0(.douta(w_n1724_0[0]),.doutb(w_n1724_0[1]),.din(n1724));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1726_0(.douta(w_n1726_0[0]),.doutb(w_n1726_0[1]),.din(n1726));
	jspl jspl_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_dff_A_5HE7nm6i7_1),.din(n1727));
	jspl jspl_w_n1734_0(.douta(w_n1734_0[0]),.doutb(w_n1734_0[1]),.din(n1734));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_dff_A_xWpozIyr6_1),.din(n1737));
	jspl jspl_w_n1739_0(.douta(w_n1739_0[0]),.doutb(w_n1739_0[1]),.din(w_dff_B_kZfnxLQn1_2));
	jspl jspl_w_n1742_0(.douta(w_n1742_0[0]),.doutb(w_n1742_0[1]),.din(w_dff_B_XI9aL1kA6_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_Gqhqk55Q6_2));
	jspl jspl_w_n1747_0(.douta(w_n1747_0[0]),.doutb(w_n1747_0[1]),.din(w_dff_B_WeM40RcL6_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(w_dff_B_EBIpuuQR8_2));
	jspl jspl_w_n1749_0(.douta(w_n1749_0[0]),.doutb(w_n1749_0[1]),.din(w_dff_B_f45WlC394_2));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1759_0(.douta(w_n1759_0[0]),.doutb(w_n1759_0[1]),.din(n1759));
	jspl jspl_w_n1760_0(.douta(w_n1760_0[0]),.doutb(w_dff_A_RXQQeR0j4_1),.din(n1760));
	jspl jspl_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.din(n1767));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_dff_A_XICyd0S42_1),.din(n1770));
	jspl jspl_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.din(w_dff_B_vc5rPiNp8_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_962kAxAN4_2));
	jspl jspl_w_n1776_0(.douta(w_n1776_0[0]),.doutb(w_n1776_0[1]),.din(w_dff_B_Lam9kCm25_2));
	jspl jspl_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.din(w_dff_B_PIWEmWL32_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl jspl_w_n1782_0(.douta(w_n1782_0[0]),.doutb(w_n1782_0[1]),.din(n1782));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1784_0(.douta(w_n1784_0[0]),.doutb(w_n1784_0[1]),.din(n1784));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_dff_A_7qFQCJai5_1),.din(n1786));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1796_0(.douta(w_n1796_0[0]),.doutb(w_dff_A_kIMEJZuV4_1),.din(n1796));
	jspl jspl_w_n1797_0(.douta(w_n1797_0[0]),.doutb(w_n1797_0[1]),.din(w_dff_B_JTBAVYp00_2));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(w_dff_B_6aixUHpW2_2));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_n1801_0[1]),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.din(n1804));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_dff_A_bKLg2vTL0_1),.din(n1805));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_TnNJYkFP3_2));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.din(n1817));
	jspl jspl_w_n1818_0(.douta(w_dff_A_L8ueDPvO2_0),.doutb(w_n1818_0[1]),.din(n1818));
	jdff dff_B_CQzbtU104_0(.din(n72),.dout(w_dff_B_CQzbtU104_0),.clk(gclk));
	jdff dff_B_lEuxbv5F0_0(.din(w_dff_B_CQzbtU104_0),.dout(w_dff_B_lEuxbv5F0_0),.clk(gclk));
	jdff dff_B_m2YFsOFD9_1(.din(n76),.dout(w_dff_B_m2YFsOFD9_1),.clk(gclk));
	jdff dff_B_b2YnYtSV1_1(.din(w_dff_B_m2YFsOFD9_1),.dout(w_dff_B_b2YnYtSV1_1),.clk(gclk));
	jdff dff_B_5LuDeCfj3_1(.din(w_dff_B_b2YnYtSV1_1),.dout(w_dff_B_5LuDeCfj3_1),.clk(gclk));
	jdff dff_B_WFVxcR7l8_1(.din(n87),.dout(w_dff_B_WFVxcR7l8_1),.clk(gclk));
	jdff dff_B_A4lZUm4M2_1(.din(w_dff_B_WFVxcR7l8_1),.dout(w_dff_B_A4lZUm4M2_1),.clk(gclk));
	jdff dff_B_6FQXuesw2_1(.din(w_dff_B_A4lZUm4M2_1),.dout(w_dff_B_6FQXuesw2_1),.clk(gclk));
	jdff dff_B_0gcEPcrz3_1(.din(w_dff_B_6FQXuesw2_1),.dout(w_dff_B_0gcEPcrz3_1),.clk(gclk));
	jdff dff_B_KvMrhP0T4_1(.din(w_dff_B_0gcEPcrz3_1),.dout(w_dff_B_KvMrhP0T4_1),.clk(gclk));
	jdff dff_B_HfeP3lcw0_1(.din(w_dff_B_KvMrhP0T4_1),.dout(w_dff_B_HfeP3lcw0_1),.clk(gclk));
	jdff dff_B_i8xu0OGh6_1(.din(n107),.dout(w_dff_B_i8xu0OGh6_1),.clk(gclk));
	jdff dff_B_OQQcgr6h1_1(.din(w_dff_B_i8xu0OGh6_1),.dout(w_dff_B_OQQcgr6h1_1),.clk(gclk));
	jdff dff_B_q9eLr02q1_1(.din(w_dff_B_OQQcgr6h1_1),.dout(w_dff_B_q9eLr02q1_1),.clk(gclk));
	jdff dff_B_I3Ru0P1g5_1(.din(w_dff_B_q9eLr02q1_1),.dout(w_dff_B_I3Ru0P1g5_1),.clk(gclk));
	jdff dff_B_7YBUKEnd7_1(.din(w_dff_B_I3Ru0P1g5_1),.dout(w_dff_B_7YBUKEnd7_1),.clk(gclk));
	jdff dff_B_Zkre0t9S8_1(.din(w_dff_B_7YBUKEnd7_1),.dout(w_dff_B_Zkre0t9S8_1),.clk(gclk));
	jdff dff_B_QCM5rOcm5_1(.din(w_dff_B_Zkre0t9S8_1),.dout(w_dff_B_QCM5rOcm5_1),.clk(gclk));
	jdff dff_B_vmjV8cet6_1(.din(w_dff_B_QCM5rOcm5_1),.dout(w_dff_B_vmjV8cet6_1),.clk(gclk));
	jdff dff_B_k71p4s1n3_1(.din(w_dff_B_vmjV8cet6_1),.dout(w_dff_B_k71p4s1n3_1),.clk(gclk));
	jdff dff_B_HH8HPvVI0_1(.din(n136),.dout(w_dff_B_HH8HPvVI0_1),.clk(gclk));
	jdff dff_B_QqQK8s0U3_1(.din(w_dff_B_HH8HPvVI0_1),.dout(w_dff_B_QqQK8s0U3_1),.clk(gclk));
	jdff dff_B_kCeu8XBG1_1(.din(w_dff_B_QqQK8s0U3_1),.dout(w_dff_B_kCeu8XBG1_1),.clk(gclk));
	jdff dff_B_dxQzISG90_1(.din(w_dff_B_kCeu8XBG1_1),.dout(w_dff_B_dxQzISG90_1),.clk(gclk));
	jdff dff_B_FGCQnwCp5_1(.din(w_dff_B_dxQzISG90_1),.dout(w_dff_B_FGCQnwCp5_1),.clk(gclk));
	jdff dff_B_1CSPJc2a0_1(.din(w_dff_B_FGCQnwCp5_1),.dout(w_dff_B_1CSPJc2a0_1),.clk(gclk));
	jdff dff_B_uPvNFZ5c1_1(.din(w_dff_B_1CSPJc2a0_1),.dout(w_dff_B_uPvNFZ5c1_1),.clk(gclk));
	jdff dff_B_BNbxdmAq4_1(.din(w_dff_B_uPvNFZ5c1_1),.dout(w_dff_B_BNbxdmAq4_1),.clk(gclk));
	jdff dff_B_tBwCKQwe8_1(.din(w_dff_B_BNbxdmAq4_1),.dout(w_dff_B_tBwCKQwe8_1),.clk(gclk));
	jdff dff_B_DPQZ5tvD5_1(.din(w_dff_B_tBwCKQwe8_1),.dout(w_dff_B_DPQZ5tvD5_1),.clk(gclk));
	jdff dff_B_fqpEbCij6_1(.din(w_dff_B_DPQZ5tvD5_1),.dout(w_dff_B_fqpEbCij6_1),.clk(gclk));
	jdff dff_B_PcDM2u6M1_1(.din(w_dff_B_fqpEbCij6_1),.dout(w_dff_B_PcDM2u6M1_1),.clk(gclk));
	jdff dff_B_yAJYlebs5_1(.din(n171),.dout(w_dff_B_yAJYlebs5_1),.clk(gclk));
	jdff dff_B_L9zoaLbS3_1(.din(w_dff_B_yAJYlebs5_1),.dout(w_dff_B_L9zoaLbS3_1),.clk(gclk));
	jdff dff_B_ZF4KR1sm0_1(.din(w_dff_B_L9zoaLbS3_1),.dout(w_dff_B_ZF4KR1sm0_1),.clk(gclk));
	jdff dff_B_IUAIBhO16_1(.din(w_dff_B_ZF4KR1sm0_1),.dout(w_dff_B_IUAIBhO16_1),.clk(gclk));
	jdff dff_B_zZlEm5fz8_1(.din(w_dff_B_IUAIBhO16_1),.dout(w_dff_B_zZlEm5fz8_1),.clk(gclk));
	jdff dff_B_vjaNgyfC6_1(.din(w_dff_B_zZlEm5fz8_1),.dout(w_dff_B_vjaNgyfC6_1),.clk(gclk));
	jdff dff_B_U7jcckH96_1(.din(w_dff_B_vjaNgyfC6_1),.dout(w_dff_B_U7jcckH96_1),.clk(gclk));
	jdff dff_B_kWtxciCH1_1(.din(w_dff_B_U7jcckH96_1),.dout(w_dff_B_kWtxciCH1_1),.clk(gclk));
	jdff dff_B_cL18KVjY0_1(.din(w_dff_B_kWtxciCH1_1),.dout(w_dff_B_cL18KVjY0_1),.clk(gclk));
	jdff dff_B_5OBCqHq93_1(.din(w_dff_B_cL18KVjY0_1),.dout(w_dff_B_5OBCqHq93_1),.clk(gclk));
	jdff dff_B_SFJx1Xso7_1(.din(w_dff_B_5OBCqHq93_1),.dout(w_dff_B_SFJx1Xso7_1),.clk(gclk));
	jdff dff_B_Kja5SFmP6_1(.din(w_dff_B_SFJx1Xso7_1),.dout(w_dff_B_Kja5SFmP6_1),.clk(gclk));
	jdff dff_B_tYDsVwD79_1(.din(w_dff_B_Kja5SFmP6_1),.dout(w_dff_B_tYDsVwD79_1),.clk(gclk));
	jdff dff_B_r7koO1Cd2_1(.din(w_dff_B_tYDsVwD79_1),.dout(w_dff_B_r7koO1Cd2_1),.clk(gclk));
	jdff dff_B_5lzuWr6g6_1(.din(w_dff_B_r7koO1Cd2_1),.dout(w_dff_B_5lzuWr6g6_1),.clk(gclk));
	jdff dff_B_rvQUMrX54_1(.din(n213),.dout(w_dff_B_rvQUMrX54_1),.clk(gclk));
	jdff dff_B_lXCG7Vdi4_1(.din(w_dff_B_rvQUMrX54_1),.dout(w_dff_B_lXCG7Vdi4_1),.clk(gclk));
	jdff dff_B_QcjPscN71_1(.din(w_dff_B_lXCG7Vdi4_1),.dout(w_dff_B_QcjPscN71_1),.clk(gclk));
	jdff dff_B_8Z8mEQet0_1(.din(w_dff_B_QcjPscN71_1),.dout(w_dff_B_8Z8mEQet0_1),.clk(gclk));
	jdff dff_B_vqGt22TA8_1(.din(w_dff_B_8Z8mEQet0_1),.dout(w_dff_B_vqGt22TA8_1),.clk(gclk));
	jdff dff_B_buYVPwG02_1(.din(w_dff_B_vqGt22TA8_1),.dout(w_dff_B_buYVPwG02_1),.clk(gclk));
	jdff dff_B_axfIYrza8_1(.din(w_dff_B_buYVPwG02_1),.dout(w_dff_B_axfIYrza8_1),.clk(gclk));
	jdff dff_B_GcG9iY9w2_1(.din(w_dff_B_axfIYrza8_1),.dout(w_dff_B_GcG9iY9w2_1),.clk(gclk));
	jdff dff_B_bOkHvbh19_1(.din(w_dff_B_GcG9iY9w2_1),.dout(w_dff_B_bOkHvbh19_1),.clk(gclk));
	jdff dff_B_DVNXvqNt3_1(.din(w_dff_B_bOkHvbh19_1),.dout(w_dff_B_DVNXvqNt3_1),.clk(gclk));
	jdff dff_B_HqbXxAvh1_1(.din(w_dff_B_DVNXvqNt3_1),.dout(w_dff_B_HqbXxAvh1_1),.clk(gclk));
	jdff dff_B_OAhj6Tw48_1(.din(w_dff_B_HqbXxAvh1_1),.dout(w_dff_B_OAhj6Tw48_1),.clk(gclk));
	jdff dff_B_aRs7Cx5P3_1(.din(w_dff_B_OAhj6Tw48_1),.dout(w_dff_B_aRs7Cx5P3_1),.clk(gclk));
	jdff dff_B_wZ0tyaKd6_1(.din(w_dff_B_aRs7Cx5P3_1),.dout(w_dff_B_wZ0tyaKd6_1),.clk(gclk));
	jdff dff_B_ZY3QDktq1_1(.din(w_dff_B_wZ0tyaKd6_1),.dout(w_dff_B_ZY3QDktq1_1),.clk(gclk));
	jdff dff_B_9qnEvK782_1(.din(w_dff_B_ZY3QDktq1_1),.dout(w_dff_B_9qnEvK782_1),.clk(gclk));
	jdff dff_B_gPfvKI8H1_1(.din(w_dff_B_9qnEvK782_1),.dout(w_dff_B_gPfvKI8H1_1),.clk(gclk));
	jdff dff_B_so7U7eC87_1(.din(w_dff_B_gPfvKI8H1_1),.dout(w_dff_B_so7U7eC87_1),.clk(gclk));
	jdff dff_B_BUyvwPbb1_1(.din(n262),.dout(w_dff_B_BUyvwPbb1_1),.clk(gclk));
	jdff dff_B_elVOzZ7q4_1(.din(w_dff_B_BUyvwPbb1_1),.dout(w_dff_B_elVOzZ7q4_1),.clk(gclk));
	jdff dff_B_Vh7Y9NNi4_1(.din(w_dff_B_elVOzZ7q4_1),.dout(w_dff_B_Vh7Y9NNi4_1),.clk(gclk));
	jdff dff_B_JULEhToh9_1(.din(w_dff_B_Vh7Y9NNi4_1),.dout(w_dff_B_JULEhToh9_1),.clk(gclk));
	jdff dff_B_ZH3oGxlj7_1(.din(w_dff_B_JULEhToh9_1),.dout(w_dff_B_ZH3oGxlj7_1),.clk(gclk));
	jdff dff_B_xsy6icMC9_1(.din(w_dff_B_ZH3oGxlj7_1),.dout(w_dff_B_xsy6icMC9_1),.clk(gclk));
	jdff dff_B_WTuFu6Cv4_1(.din(w_dff_B_xsy6icMC9_1),.dout(w_dff_B_WTuFu6Cv4_1),.clk(gclk));
	jdff dff_B_cRFxGYkK1_1(.din(w_dff_B_WTuFu6Cv4_1),.dout(w_dff_B_cRFxGYkK1_1),.clk(gclk));
	jdff dff_B_AgMqf6K30_1(.din(w_dff_B_cRFxGYkK1_1),.dout(w_dff_B_AgMqf6K30_1),.clk(gclk));
	jdff dff_B_XYW3L56N0_1(.din(w_dff_B_AgMqf6K30_1),.dout(w_dff_B_XYW3L56N0_1),.clk(gclk));
	jdff dff_B_lQf1FyrY4_1(.din(w_dff_B_XYW3L56N0_1),.dout(w_dff_B_lQf1FyrY4_1),.clk(gclk));
	jdff dff_B_CLGPZbuj3_1(.din(w_dff_B_lQf1FyrY4_1),.dout(w_dff_B_CLGPZbuj3_1),.clk(gclk));
	jdff dff_B_4CV3vP6I7_1(.din(w_dff_B_CLGPZbuj3_1),.dout(w_dff_B_4CV3vP6I7_1),.clk(gclk));
	jdff dff_B_RUUqzdH85_1(.din(w_dff_B_4CV3vP6I7_1),.dout(w_dff_B_RUUqzdH85_1),.clk(gclk));
	jdff dff_B_A4zxo8ba5_1(.din(w_dff_B_RUUqzdH85_1),.dout(w_dff_B_A4zxo8ba5_1),.clk(gclk));
	jdff dff_B_PkSuJ1jH0_1(.din(w_dff_B_A4zxo8ba5_1),.dout(w_dff_B_PkSuJ1jH0_1),.clk(gclk));
	jdff dff_B_IwnpOftq1_1(.din(w_dff_B_PkSuJ1jH0_1),.dout(w_dff_B_IwnpOftq1_1),.clk(gclk));
	jdff dff_B_rgS15Ok66_1(.din(w_dff_B_IwnpOftq1_1),.dout(w_dff_B_rgS15Ok66_1),.clk(gclk));
	jdff dff_B_EpuBHSCh7_1(.din(w_dff_B_rgS15Ok66_1),.dout(w_dff_B_EpuBHSCh7_1),.clk(gclk));
	jdff dff_B_0esQzCRK8_1(.din(w_dff_B_EpuBHSCh7_1),.dout(w_dff_B_0esQzCRK8_1),.clk(gclk));
	jdff dff_B_m3PEL1Gm3_1(.din(w_dff_B_0esQzCRK8_1),.dout(w_dff_B_m3PEL1Gm3_1),.clk(gclk));
	jdff dff_B_om5yi6oo6_1(.din(n318),.dout(w_dff_B_om5yi6oo6_1),.clk(gclk));
	jdff dff_B_RNaMrRvH6_1(.din(w_dff_B_om5yi6oo6_1),.dout(w_dff_B_RNaMrRvH6_1),.clk(gclk));
	jdff dff_B_SENSpIqz4_1(.din(w_dff_B_RNaMrRvH6_1),.dout(w_dff_B_SENSpIqz4_1),.clk(gclk));
	jdff dff_B_P9Uq7ySz0_1(.din(w_dff_B_SENSpIqz4_1),.dout(w_dff_B_P9Uq7ySz0_1),.clk(gclk));
	jdff dff_B_gGLWvwHE0_1(.din(w_dff_B_P9Uq7ySz0_1),.dout(w_dff_B_gGLWvwHE0_1),.clk(gclk));
	jdff dff_B_5xawmo587_1(.din(w_dff_B_gGLWvwHE0_1),.dout(w_dff_B_5xawmo587_1),.clk(gclk));
	jdff dff_B_HF85Sorq0_1(.din(w_dff_B_5xawmo587_1),.dout(w_dff_B_HF85Sorq0_1),.clk(gclk));
	jdff dff_B_McV18ixf3_1(.din(w_dff_B_HF85Sorq0_1),.dout(w_dff_B_McV18ixf3_1),.clk(gclk));
	jdff dff_B_tspBcsNe5_1(.din(w_dff_B_McV18ixf3_1),.dout(w_dff_B_tspBcsNe5_1),.clk(gclk));
	jdff dff_B_8KvmIXAE4_1(.din(w_dff_B_tspBcsNe5_1),.dout(w_dff_B_8KvmIXAE4_1),.clk(gclk));
	jdff dff_B_1PlvDrQ21_1(.din(w_dff_B_8KvmIXAE4_1),.dout(w_dff_B_1PlvDrQ21_1),.clk(gclk));
	jdff dff_B_RRqtvSfw5_1(.din(w_dff_B_1PlvDrQ21_1),.dout(w_dff_B_RRqtvSfw5_1),.clk(gclk));
	jdff dff_B_nSHEtc8K3_1(.din(w_dff_B_RRqtvSfw5_1),.dout(w_dff_B_nSHEtc8K3_1),.clk(gclk));
	jdff dff_B_p4kuG29k6_1(.din(w_dff_B_nSHEtc8K3_1),.dout(w_dff_B_p4kuG29k6_1),.clk(gclk));
	jdff dff_B_dd5qWz7c1_1(.din(w_dff_B_p4kuG29k6_1),.dout(w_dff_B_dd5qWz7c1_1),.clk(gclk));
	jdff dff_B_G8juxv5v1_1(.din(w_dff_B_dd5qWz7c1_1),.dout(w_dff_B_G8juxv5v1_1),.clk(gclk));
	jdff dff_B_s2YN9vxX1_1(.din(w_dff_B_G8juxv5v1_1),.dout(w_dff_B_s2YN9vxX1_1),.clk(gclk));
	jdff dff_B_5YcMWnSx7_1(.din(w_dff_B_s2YN9vxX1_1),.dout(w_dff_B_5YcMWnSx7_1),.clk(gclk));
	jdff dff_B_GfcNu1Pm8_1(.din(w_dff_B_5YcMWnSx7_1),.dout(w_dff_B_GfcNu1Pm8_1),.clk(gclk));
	jdff dff_B_Q0U8vNiJ5_1(.din(w_dff_B_GfcNu1Pm8_1),.dout(w_dff_B_Q0U8vNiJ5_1),.clk(gclk));
	jdff dff_B_RTNinQqY8_1(.din(w_dff_B_Q0U8vNiJ5_1),.dout(w_dff_B_RTNinQqY8_1),.clk(gclk));
	jdff dff_B_xgb81Vz88_1(.din(w_dff_B_RTNinQqY8_1),.dout(w_dff_B_xgb81Vz88_1),.clk(gclk));
	jdff dff_B_RoA3tBvL4_1(.din(w_dff_B_xgb81Vz88_1),.dout(w_dff_B_RoA3tBvL4_1),.clk(gclk));
	jdff dff_B_vGQOMZBB4_1(.din(w_dff_B_RoA3tBvL4_1),.dout(w_dff_B_vGQOMZBB4_1),.clk(gclk));
	jdff dff_B_1thrLE4J6_1(.din(n381),.dout(w_dff_B_1thrLE4J6_1),.clk(gclk));
	jdff dff_B_d6xtxwtY7_1(.din(w_dff_B_1thrLE4J6_1),.dout(w_dff_B_d6xtxwtY7_1),.clk(gclk));
	jdff dff_B_pBJyrQGT0_1(.din(w_dff_B_d6xtxwtY7_1),.dout(w_dff_B_pBJyrQGT0_1),.clk(gclk));
	jdff dff_B_zfMrTPdX8_1(.din(w_dff_B_pBJyrQGT0_1),.dout(w_dff_B_zfMrTPdX8_1),.clk(gclk));
	jdff dff_B_rqsZCN590_1(.din(w_dff_B_zfMrTPdX8_1),.dout(w_dff_B_rqsZCN590_1),.clk(gclk));
	jdff dff_B_RgPVaUv77_1(.din(w_dff_B_rqsZCN590_1),.dout(w_dff_B_RgPVaUv77_1),.clk(gclk));
	jdff dff_B_2YqoXrLH1_1(.din(w_dff_B_RgPVaUv77_1),.dout(w_dff_B_2YqoXrLH1_1),.clk(gclk));
	jdff dff_B_oRoaPbra3_1(.din(w_dff_B_2YqoXrLH1_1),.dout(w_dff_B_oRoaPbra3_1),.clk(gclk));
	jdff dff_B_xaVLPsu49_1(.din(w_dff_B_oRoaPbra3_1),.dout(w_dff_B_xaVLPsu49_1),.clk(gclk));
	jdff dff_B_wQlgNhLa9_1(.din(w_dff_B_xaVLPsu49_1),.dout(w_dff_B_wQlgNhLa9_1),.clk(gclk));
	jdff dff_B_WrfQEx1C9_1(.din(w_dff_B_wQlgNhLa9_1),.dout(w_dff_B_WrfQEx1C9_1),.clk(gclk));
	jdff dff_B_Sd5vFueX7_1(.din(w_dff_B_WrfQEx1C9_1),.dout(w_dff_B_Sd5vFueX7_1),.clk(gclk));
	jdff dff_B_SN7GOMXW4_1(.din(w_dff_B_Sd5vFueX7_1),.dout(w_dff_B_SN7GOMXW4_1),.clk(gclk));
	jdff dff_B_fK4bgWEk7_1(.din(w_dff_B_SN7GOMXW4_1),.dout(w_dff_B_fK4bgWEk7_1),.clk(gclk));
	jdff dff_B_fW7d0Ilt6_1(.din(w_dff_B_fK4bgWEk7_1),.dout(w_dff_B_fW7d0Ilt6_1),.clk(gclk));
	jdff dff_B_Uq6KDSWv2_1(.din(w_dff_B_fW7d0Ilt6_1),.dout(w_dff_B_Uq6KDSWv2_1),.clk(gclk));
	jdff dff_B_JW9BKxOH9_1(.din(w_dff_B_Uq6KDSWv2_1),.dout(w_dff_B_JW9BKxOH9_1),.clk(gclk));
	jdff dff_B_JV781Cy01_1(.din(w_dff_B_JW9BKxOH9_1),.dout(w_dff_B_JV781Cy01_1),.clk(gclk));
	jdff dff_B_bY10uaJ73_1(.din(w_dff_B_JV781Cy01_1),.dout(w_dff_B_bY10uaJ73_1),.clk(gclk));
	jdff dff_B_sgIQiEtB3_1(.din(w_dff_B_bY10uaJ73_1),.dout(w_dff_B_sgIQiEtB3_1),.clk(gclk));
	jdff dff_B_C2SNLFqJ7_1(.din(w_dff_B_sgIQiEtB3_1),.dout(w_dff_B_C2SNLFqJ7_1),.clk(gclk));
	jdff dff_B_ahZNrPcM3_1(.din(w_dff_B_C2SNLFqJ7_1),.dout(w_dff_B_ahZNrPcM3_1),.clk(gclk));
	jdff dff_B_PRVmNAZi2_1(.din(w_dff_B_ahZNrPcM3_1),.dout(w_dff_B_PRVmNAZi2_1),.clk(gclk));
	jdff dff_B_JoZcubzt1_1(.din(w_dff_B_PRVmNAZi2_1),.dout(w_dff_B_JoZcubzt1_1),.clk(gclk));
	jdff dff_B_n3g5oXJa5_1(.din(w_dff_B_JoZcubzt1_1),.dout(w_dff_B_n3g5oXJa5_1),.clk(gclk));
	jdff dff_B_BznF3FIb6_1(.din(w_dff_B_n3g5oXJa5_1),.dout(w_dff_B_BznF3FIb6_1),.clk(gclk));
	jdff dff_B_0X766xLg1_1(.din(w_dff_B_BznF3FIb6_1),.dout(w_dff_B_0X766xLg1_1),.clk(gclk));
	jdff dff_B_Ohaxnjpv1_1(.din(n452),.dout(w_dff_B_Ohaxnjpv1_1),.clk(gclk));
	jdff dff_B_Wv2zYr603_1(.din(w_dff_B_Ohaxnjpv1_1),.dout(w_dff_B_Wv2zYr603_1),.clk(gclk));
	jdff dff_B_qCibCRSU7_1(.din(w_dff_B_Wv2zYr603_1),.dout(w_dff_B_qCibCRSU7_1),.clk(gclk));
	jdff dff_B_esUgqMcf7_1(.din(w_dff_B_qCibCRSU7_1),.dout(w_dff_B_esUgqMcf7_1),.clk(gclk));
	jdff dff_B_g5YFE9H99_1(.din(w_dff_B_esUgqMcf7_1),.dout(w_dff_B_g5YFE9H99_1),.clk(gclk));
	jdff dff_B_QQv9vc7A3_1(.din(w_dff_B_g5YFE9H99_1),.dout(w_dff_B_QQv9vc7A3_1),.clk(gclk));
	jdff dff_B_QcL6UJab8_1(.din(w_dff_B_QQv9vc7A3_1),.dout(w_dff_B_QcL6UJab8_1),.clk(gclk));
	jdff dff_B_TSTDwVwp3_1(.din(w_dff_B_QcL6UJab8_1),.dout(w_dff_B_TSTDwVwp3_1),.clk(gclk));
	jdff dff_B_Uf0UaQSc9_1(.din(w_dff_B_TSTDwVwp3_1),.dout(w_dff_B_Uf0UaQSc9_1),.clk(gclk));
	jdff dff_B_xKDbCvj80_1(.din(w_dff_B_Uf0UaQSc9_1),.dout(w_dff_B_xKDbCvj80_1),.clk(gclk));
	jdff dff_B_a9NgOcio2_1(.din(w_dff_B_xKDbCvj80_1),.dout(w_dff_B_a9NgOcio2_1),.clk(gclk));
	jdff dff_B_HcrrAszy4_1(.din(w_dff_B_a9NgOcio2_1),.dout(w_dff_B_HcrrAszy4_1),.clk(gclk));
	jdff dff_B_BX3Q1osR8_1(.din(w_dff_B_HcrrAszy4_1),.dout(w_dff_B_BX3Q1osR8_1),.clk(gclk));
	jdff dff_B_b7YPd1iR0_1(.din(w_dff_B_BX3Q1osR8_1),.dout(w_dff_B_b7YPd1iR0_1),.clk(gclk));
	jdff dff_B_mKgddXPJ7_1(.din(w_dff_B_b7YPd1iR0_1),.dout(w_dff_B_mKgddXPJ7_1),.clk(gclk));
	jdff dff_B_Ul9xBQiK3_1(.din(w_dff_B_mKgddXPJ7_1),.dout(w_dff_B_Ul9xBQiK3_1),.clk(gclk));
	jdff dff_B_TpvobFwx6_1(.din(w_dff_B_Ul9xBQiK3_1),.dout(w_dff_B_TpvobFwx6_1),.clk(gclk));
	jdff dff_B_lpnll1dX3_1(.din(w_dff_B_TpvobFwx6_1),.dout(w_dff_B_lpnll1dX3_1),.clk(gclk));
	jdff dff_B_RYRal4Ol3_1(.din(w_dff_B_lpnll1dX3_1),.dout(w_dff_B_RYRal4Ol3_1),.clk(gclk));
	jdff dff_B_hHpZTndD7_1(.din(w_dff_B_RYRal4Ol3_1),.dout(w_dff_B_hHpZTndD7_1),.clk(gclk));
	jdff dff_B_3B7n4IN74_1(.din(w_dff_B_hHpZTndD7_1),.dout(w_dff_B_3B7n4IN74_1),.clk(gclk));
	jdff dff_B_x8QwSilg4_1(.din(w_dff_B_3B7n4IN74_1),.dout(w_dff_B_x8QwSilg4_1),.clk(gclk));
	jdff dff_B_apnd5IDr9_1(.din(w_dff_B_x8QwSilg4_1),.dout(w_dff_B_apnd5IDr9_1),.clk(gclk));
	jdff dff_B_IHiiTo3O6_1(.din(w_dff_B_apnd5IDr9_1),.dout(w_dff_B_IHiiTo3O6_1),.clk(gclk));
	jdff dff_B_sIpOpXkx0_1(.din(w_dff_B_IHiiTo3O6_1),.dout(w_dff_B_sIpOpXkx0_1),.clk(gclk));
	jdff dff_B_s83mAJLg8_1(.din(w_dff_B_sIpOpXkx0_1),.dout(w_dff_B_s83mAJLg8_1),.clk(gclk));
	jdff dff_B_yeVQDdmo1_1(.din(w_dff_B_s83mAJLg8_1),.dout(w_dff_B_yeVQDdmo1_1),.clk(gclk));
	jdff dff_B_zfGdRU5l7_1(.din(w_dff_B_yeVQDdmo1_1),.dout(w_dff_B_zfGdRU5l7_1),.clk(gclk));
	jdff dff_B_67DesMrR9_1(.din(w_dff_B_zfGdRU5l7_1),.dout(w_dff_B_67DesMrR9_1),.clk(gclk));
	jdff dff_B_1Aoe1Zp02_1(.din(w_dff_B_67DesMrR9_1),.dout(w_dff_B_1Aoe1Zp02_1),.clk(gclk));
	jdff dff_B_KJ8ERTgx0_1(.din(n530),.dout(w_dff_B_KJ8ERTgx0_1),.clk(gclk));
	jdff dff_B_t6pgtpSN5_1(.din(w_dff_B_KJ8ERTgx0_1),.dout(w_dff_B_t6pgtpSN5_1),.clk(gclk));
	jdff dff_B_0wvmjINJ5_1(.din(w_dff_B_t6pgtpSN5_1),.dout(w_dff_B_0wvmjINJ5_1),.clk(gclk));
	jdff dff_B_c1bT9x5k3_1(.din(w_dff_B_0wvmjINJ5_1),.dout(w_dff_B_c1bT9x5k3_1),.clk(gclk));
	jdff dff_B_4LN2QOOh6_1(.din(w_dff_B_c1bT9x5k3_1),.dout(w_dff_B_4LN2QOOh6_1),.clk(gclk));
	jdff dff_B_OfhxVnc54_1(.din(w_dff_B_4LN2QOOh6_1),.dout(w_dff_B_OfhxVnc54_1),.clk(gclk));
	jdff dff_B_tiIEoovw4_1(.din(w_dff_B_OfhxVnc54_1),.dout(w_dff_B_tiIEoovw4_1),.clk(gclk));
	jdff dff_B_b53M9FKu8_1(.din(w_dff_B_tiIEoovw4_1),.dout(w_dff_B_b53M9FKu8_1),.clk(gclk));
	jdff dff_B_XxgO3fsy4_1(.din(w_dff_B_b53M9FKu8_1),.dout(w_dff_B_XxgO3fsy4_1),.clk(gclk));
	jdff dff_B_Xlc5vSBR1_1(.din(w_dff_B_XxgO3fsy4_1),.dout(w_dff_B_Xlc5vSBR1_1),.clk(gclk));
	jdff dff_B_aoAsfADC9_1(.din(w_dff_B_Xlc5vSBR1_1),.dout(w_dff_B_aoAsfADC9_1),.clk(gclk));
	jdff dff_B_2Mb77foR9_1(.din(w_dff_B_aoAsfADC9_1),.dout(w_dff_B_2Mb77foR9_1),.clk(gclk));
	jdff dff_B_5WwukQxC4_1(.din(w_dff_B_2Mb77foR9_1),.dout(w_dff_B_5WwukQxC4_1),.clk(gclk));
	jdff dff_B_RQ5xwhgu3_1(.din(w_dff_B_5WwukQxC4_1),.dout(w_dff_B_RQ5xwhgu3_1),.clk(gclk));
	jdff dff_B_bYMdPLlh5_1(.din(w_dff_B_RQ5xwhgu3_1),.dout(w_dff_B_bYMdPLlh5_1),.clk(gclk));
	jdff dff_B_iwxCcSjO6_1(.din(w_dff_B_bYMdPLlh5_1),.dout(w_dff_B_iwxCcSjO6_1),.clk(gclk));
	jdff dff_B_fQfxNQOK0_1(.din(w_dff_B_iwxCcSjO6_1),.dout(w_dff_B_fQfxNQOK0_1),.clk(gclk));
	jdff dff_B_s8kfIGKo6_1(.din(w_dff_B_fQfxNQOK0_1),.dout(w_dff_B_s8kfIGKo6_1),.clk(gclk));
	jdff dff_B_tyYRCZIO8_1(.din(w_dff_B_s8kfIGKo6_1),.dout(w_dff_B_tyYRCZIO8_1),.clk(gclk));
	jdff dff_B_OEb6m1KX0_1(.din(w_dff_B_tyYRCZIO8_1),.dout(w_dff_B_OEb6m1KX0_1),.clk(gclk));
	jdff dff_B_Vo9cFIp64_1(.din(w_dff_B_OEb6m1KX0_1),.dout(w_dff_B_Vo9cFIp64_1),.clk(gclk));
	jdff dff_B_8y9R6sCY2_1(.din(w_dff_B_Vo9cFIp64_1),.dout(w_dff_B_8y9R6sCY2_1),.clk(gclk));
	jdff dff_B_tmAYfzY61_1(.din(w_dff_B_8y9R6sCY2_1),.dout(w_dff_B_tmAYfzY61_1),.clk(gclk));
	jdff dff_B_LL1POgVB0_1(.din(w_dff_B_tmAYfzY61_1),.dout(w_dff_B_LL1POgVB0_1),.clk(gclk));
	jdff dff_B_1ywzHM0E6_1(.din(w_dff_B_LL1POgVB0_1),.dout(w_dff_B_1ywzHM0E6_1),.clk(gclk));
	jdff dff_B_G2YRkX784_1(.din(w_dff_B_1ywzHM0E6_1),.dout(w_dff_B_G2YRkX784_1),.clk(gclk));
	jdff dff_B_euuIZCO06_1(.din(w_dff_B_G2YRkX784_1),.dout(w_dff_B_euuIZCO06_1),.clk(gclk));
	jdff dff_B_AOLl8XXU4_1(.din(w_dff_B_euuIZCO06_1),.dout(w_dff_B_AOLl8XXU4_1),.clk(gclk));
	jdff dff_B_3tJ6Ru2z1_1(.din(w_dff_B_AOLl8XXU4_1),.dout(w_dff_B_3tJ6Ru2z1_1),.clk(gclk));
	jdff dff_B_1xWW39aW4_1(.din(w_dff_B_3tJ6Ru2z1_1),.dout(w_dff_B_1xWW39aW4_1),.clk(gclk));
	jdff dff_B_igPDpLnN4_1(.din(w_dff_B_1xWW39aW4_1),.dout(w_dff_B_igPDpLnN4_1),.clk(gclk));
	jdff dff_B_BQUck8pw6_1(.din(w_dff_B_igPDpLnN4_1),.dout(w_dff_B_BQUck8pw6_1),.clk(gclk));
	jdff dff_B_EMXdE2Dp7_1(.din(w_dff_B_BQUck8pw6_1),.dout(w_dff_B_EMXdE2Dp7_1),.clk(gclk));
	jdff dff_B_o5KyN9Av8_1(.din(n615),.dout(w_dff_B_o5KyN9Av8_1),.clk(gclk));
	jdff dff_B_iRKRjkPD3_1(.din(w_dff_B_o5KyN9Av8_1),.dout(w_dff_B_iRKRjkPD3_1),.clk(gclk));
	jdff dff_B_bNiXRNEt7_1(.din(w_dff_B_iRKRjkPD3_1),.dout(w_dff_B_bNiXRNEt7_1),.clk(gclk));
	jdff dff_B_VEZuYu6E5_1(.din(w_dff_B_bNiXRNEt7_1),.dout(w_dff_B_VEZuYu6E5_1),.clk(gclk));
	jdff dff_B_b0yhfW5y1_1(.din(w_dff_B_VEZuYu6E5_1),.dout(w_dff_B_b0yhfW5y1_1),.clk(gclk));
	jdff dff_B_XmdeWYy09_1(.din(w_dff_B_b0yhfW5y1_1),.dout(w_dff_B_XmdeWYy09_1),.clk(gclk));
	jdff dff_B_RvcMJutV0_1(.din(w_dff_B_XmdeWYy09_1),.dout(w_dff_B_RvcMJutV0_1),.clk(gclk));
	jdff dff_B_q54efvMt6_1(.din(w_dff_B_RvcMJutV0_1),.dout(w_dff_B_q54efvMt6_1),.clk(gclk));
	jdff dff_B_LZfvazFs7_1(.din(w_dff_B_q54efvMt6_1),.dout(w_dff_B_LZfvazFs7_1),.clk(gclk));
	jdff dff_B_zkdoqCH55_1(.din(w_dff_B_LZfvazFs7_1),.dout(w_dff_B_zkdoqCH55_1),.clk(gclk));
	jdff dff_B_ldcZC9kl6_1(.din(w_dff_B_zkdoqCH55_1),.dout(w_dff_B_ldcZC9kl6_1),.clk(gclk));
	jdff dff_B_zyZGnLg48_1(.din(w_dff_B_ldcZC9kl6_1),.dout(w_dff_B_zyZGnLg48_1),.clk(gclk));
	jdff dff_B_6PCwuYHb9_1(.din(w_dff_B_zyZGnLg48_1),.dout(w_dff_B_6PCwuYHb9_1),.clk(gclk));
	jdff dff_B_KO4JF4GX2_1(.din(w_dff_B_6PCwuYHb9_1),.dout(w_dff_B_KO4JF4GX2_1),.clk(gclk));
	jdff dff_B_xlK0L1Ug7_1(.din(w_dff_B_KO4JF4GX2_1),.dout(w_dff_B_xlK0L1Ug7_1),.clk(gclk));
	jdff dff_B_wJjdlrfB6_1(.din(w_dff_B_xlK0L1Ug7_1),.dout(w_dff_B_wJjdlrfB6_1),.clk(gclk));
	jdff dff_B_3Ji2gMQm7_1(.din(w_dff_B_wJjdlrfB6_1),.dout(w_dff_B_3Ji2gMQm7_1),.clk(gclk));
	jdff dff_B_PfB9bUjh7_1(.din(w_dff_B_3Ji2gMQm7_1),.dout(w_dff_B_PfB9bUjh7_1),.clk(gclk));
	jdff dff_B_dC8IHqIJ1_1(.din(w_dff_B_PfB9bUjh7_1),.dout(w_dff_B_dC8IHqIJ1_1),.clk(gclk));
	jdff dff_B_HBS5AwK51_1(.din(w_dff_B_dC8IHqIJ1_1),.dout(w_dff_B_HBS5AwK51_1),.clk(gclk));
	jdff dff_B_EouPxaki8_1(.din(w_dff_B_HBS5AwK51_1),.dout(w_dff_B_EouPxaki8_1),.clk(gclk));
	jdff dff_B_RrulAtdA1_1(.din(w_dff_B_EouPxaki8_1),.dout(w_dff_B_RrulAtdA1_1),.clk(gclk));
	jdff dff_B_pF2aKIxn5_1(.din(w_dff_B_RrulAtdA1_1),.dout(w_dff_B_pF2aKIxn5_1),.clk(gclk));
	jdff dff_B_MU30OuBi8_1(.din(w_dff_B_pF2aKIxn5_1),.dout(w_dff_B_MU30OuBi8_1),.clk(gclk));
	jdff dff_B_2OfEKHBX4_1(.din(w_dff_B_MU30OuBi8_1),.dout(w_dff_B_2OfEKHBX4_1),.clk(gclk));
	jdff dff_B_LS0Nnnbe9_1(.din(w_dff_B_2OfEKHBX4_1),.dout(w_dff_B_LS0Nnnbe9_1),.clk(gclk));
	jdff dff_B_UI1ALbJ59_1(.din(w_dff_B_LS0Nnnbe9_1),.dout(w_dff_B_UI1ALbJ59_1),.clk(gclk));
	jdff dff_B_i2YItJvF0_1(.din(w_dff_B_UI1ALbJ59_1),.dout(w_dff_B_i2YItJvF0_1),.clk(gclk));
	jdff dff_B_u8OfvAuj2_1(.din(w_dff_B_i2YItJvF0_1),.dout(w_dff_B_u8OfvAuj2_1),.clk(gclk));
	jdff dff_B_46lwCQV27_1(.din(w_dff_B_u8OfvAuj2_1),.dout(w_dff_B_46lwCQV27_1),.clk(gclk));
	jdff dff_B_ieZy9wnn7_1(.din(w_dff_B_46lwCQV27_1),.dout(w_dff_B_ieZy9wnn7_1),.clk(gclk));
	jdff dff_B_UM2IZ2TQ9_1(.din(w_dff_B_ieZy9wnn7_1),.dout(w_dff_B_UM2IZ2TQ9_1),.clk(gclk));
	jdff dff_B_G7fpRx6n5_1(.din(w_dff_B_UM2IZ2TQ9_1),.dout(w_dff_B_G7fpRx6n5_1),.clk(gclk));
	jdff dff_B_lWOX5vnu7_1(.din(w_dff_B_G7fpRx6n5_1),.dout(w_dff_B_lWOX5vnu7_1),.clk(gclk));
	jdff dff_B_w8mdgQxL8_1(.din(w_dff_B_lWOX5vnu7_1),.dout(w_dff_B_w8mdgQxL8_1),.clk(gclk));
	jdff dff_B_g0rjQRyU7_1(.din(w_dff_B_w8mdgQxL8_1),.dout(w_dff_B_g0rjQRyU7_1),.clk(gclk));
	jdff dff_B_mSkAwcO57_1(.din(n707),.dout(w_dff_B_mSkAwcO57_1),.clk(gclk));
	jdff dff_B_8aKZDA7T4_1(.din(w_dff_B_mSkAwcO57_1),.dout(w_dff_B_8aKZDA7T4_1),.clk(gclk));
	jdff dff_B_qiYe6hHG4_1(.din(w_dff_B_8aKZDA7T4_1),.dout(w_dff_B_qiYe6hHG4_1),.clk(gclk));
	jdff dff_B_p2oC7vdN4_1(.din(w_dff_B_qiYe6hHG4_1),.dout(w_dff_B_p2oC7vdN4_1),.clk(gclk));
	jdff dff_B_JbZNPpgs7_1(.din(w_dff_B_p2oC7vdN4_1),.dout(w_dff_B_JbZNPpgs7_1),.clk(gclk));
	jdff dff_B_HaaH6aMG8_1(.din(w_dff_B_JbZNPpgs7_1),.dout(w_dff_B_HaaH6aMG8_1),.clk(gclk));
	jdff dff_B_J7folQdM4_1(.din(w_dff_B_HaaH6aMG8_1),.dout(w_dff_B_J7folQdM4_1),.clk(gclk));
	jdff dff_B_yizmqqar9_1(.din(w_dff_B_J7folQdM4_1),.dout(w_dff_B_yizmqqar9_1),.clk(gclk));
	jdff dff_B_35aKkuzV0_1(.din(w_dff_B_yizmqqar9_1),.dout(w_dff_B_35aKkuzV0_1),.clk(gclk));
	jdff dff_B_EHn5wVSy5_1(.din(w_dff_B_35aKkuzV0_1),.dout(w_dff_B_EHn5wVSy5_1),.clk(gclk));
	jdff dff_B_JFgDmkrW3_1(.din(w_dff_B_EHn5wVSy5_1),.dout(w_dff_B_JFgDmkrW3_1),.clk(gclk));
	jdff dff_B_uXi9tDhs3_1(.din(w_dff_B_JFgDmkrW3_1),.dout(w_dff_B_uXi9tDhs3_1),.clk(gclk));
	jdff dff_B_vdqwhCzo3_1(.din(w_dff_B_uXi9tDhs3_1),.dout(w_dff_B_vdqwhCzo3_1),.clk(gclk));
	jdff dff_B_FqzXHXep2_1(.din(w_dff_B_vdqwhCzo3_1),.dout(w_dff_B_FqzXHXep2_1),.clk(gclk));
	jdff dff_B_5UKeuiYK9_1(.din(w_dff_B_FqzXHXep2_1),.dout(w_dff_B_5UKeuiYK9_1),.clk(gclk));
	jdff dff_B_qvxQFtuE9_1(.din(w_dff_B_5UKeuiYK9_1),.dout(w_dff_B_qvxQFtuE9_1),.clk(gclk));
	jdff dff_B_bXpVsNP53_1(.din(w_dff_B_qvxQFtuE9_1),.dout(w_dff_B_bXpVsNP53_1),.clk(gclk));
	jdff dff_B_0fmmWaq16_1(.din(w_dff_B_bXpVsNP53_1),.dout(w_dff_B_0fmmWaq16_1),.clk(gclk));
	jdff dff_B_OeStJnji3_1(.din(w_dff_B_0fmmWaq16_1),.dout(w_dff_B_OeStJnji3_1),.clk(gclk));
	jdff dff_B_LDuQEcWd1_1(.din(w_dff_B_OeStJnji3_1),.dout(w_dff_B_LDuQEcWd1_1),.clk(gclk));
	jdff dff_B_xifPqPjM2_1(.din(w_dff_B_LDuQEcWd1_1),.dout(w_dff_B_xifPqPjM2_1),.clk(gclk));
	jdff dff_B_tXSItKuV4_1(.din(w_dff_B_xifPqPjM2_1),.dout(w_dff_B_tXSItKuV4_1),.clk(gclk));
	jdff dff_B_i0Qc3n010_1(.din(w_dff_B_tXSItKuV4_1),.dout(w_dff_B_i0Qc3n010_1),.clk(gclk));
	jdff dff_B_4Qc3BT602_1(.din(w_dff_B_i0Qc3n010_1),.dout(w_dff_B_4Qc3BT602_1),.clk(gclk));
	jdff dff_B_oKhZ9Px72_1(.din(w_dff_B_4Qc3BT602_1),.dout(w_dff_B_oKhZ9Px72_1),.clk(gclk));
	jdff dff_B_r7Cgy82A9_1(.din(w_dff_B_oKhZ9Px72_1),.dout(w_dff_B_r7Cgy82A9_1),.clk(gclk));
	jdff dff_B_azoRYASO7_1(.din(w_dff_B_r7Cgy82A9_1),.dout(w_dff_B_azoRYASO7_1),.clk(gclk));
	jdff dff_B_5LPQTviR3_1(.din(w_dff_B_azoRYASO7_1),.dout(w_dff_B_5LPQTviR3_1),.clk(gclk));
	jdff dff_B_oalh4PKc8_1(.din(w_dff_B_5LPQTviR3_1),.dout(w_dff_B_oalh4PKc8_1),.clk(gclk));
	jdff dff_B_VSJ31bKI6_1(.din(w_dff_B_oalh4PKc8_1),.dout(w_dff_B_VSJ31bKI6_1),.clk(gclk));
	jdff dff_B_ERF1bee34_1(.din(w_dff_B_VSJ31bKI6_1),.dout(w_dff_B_ERF1bee34_1),.clk(gclk));
	jdff dff_B_GjShUze15_1(.din(w_dff_B_ERF1bee34_1),.dout(w_dff_B_GjShUze15_1),.clk(gclk));
	jdff dff_B_xBN9sYd73_1(.din(w_dff_B_GjShUze15_1),.dout(w_dff_B_xBN9sYd73_1),.clk(gclk));
	jdff dff_B_TrtEvN463_1(.din(w_dff_B_xBN9sYd73_1),.dout(w_dff_B_TrtEvN463_1),.clk(gclk));
	jdff dff_B_Dto28vYA0_1(.din(w_dff_B_TrtEvN463_1),.dout(w_dff_B_Dto28vYA0_1),.clk(gclk));
	jdff dff_B_Wd6tI4do1_1(.din(w_dff_B_Dto28vYA0_1),.dout(w_dff_B_Wd6tI4do1_1),.clk(gclk));
	jdff dff_B_nrI87EEZ2_1(.din(w_dff_B_Wd6tI4do1_1),.dout(w_dff_B_nrI87EEZ2_1),.clk(gclk));
	jdff dff_B_WuR5d0mp4_1(.din(w_dff_B_nrI87EEZ2_1),.dout(w_dff_B_WuR5d0mp4_1),.clk(gclk));
	jdff dff_B_R5ONn5iw7_1(.din(w_dff_B_WuR5d0mp4_1),.dout(w_dff_B_R5ONn5iw7_1),.clk(gclk));
	jdff dff_B_PP0smkJr0_1(.din(n806),.dout(w_dff_B_PP0smkJr0_1),.clk(gclk));
	jdff dff_B_Z6uSNpOy7_1(.din(w_dff_B_PP0smkJr0_1),.dout(w_dff_B_Z6uSNpOy7_1),.clk(gclk));
	jdff dff_B_FkH7Nsub6_1(.din(w_dff_B_Z6uSNpOy7_1),.dout(w_dff_B_FkH7Nsub6_1),.clk(gclk));
	jdff dff_B_bMddaBju1_1(.din(w_dff_B_FkH7Nsub6_1),.dout(w_dff_B_bMddaBju1_1),.clk(gclk));
	jdff dff_B_aNQnMqfL8_1(.din(w_dff_B_bMddaBju1_1),.dout(w_dff_B_aNQnMqfL8_1),.clk(gclk));
	jdff dff_B_cfoY5vZH4_1(.din(w_dff_B_aNQnMqfL8_1),.dout(w_dff_B_cfoY5vZH4_1),.clk(gclk));
	jdff dff_B_D1TEAkdy4_1(.din(w_dff_B_cfoY5vZH4_1),.dout(w_dff_B_D1TEAkdy4_1),.clk(gclk));
	jdff dff_B_nYixf4ck7_1(.din(w_dff_B_D1TEAkdy4_1),.dout(w_dff_B_nYixf4ck7_1),.clk(gclk));
	jdff dff_B_E7GihjsA6_1(.din(w_dff_B_nYixf4ck7_1),.dout(w_dff_B_E7GihjsA6_1),.clk(gclk));
	jdff dff_B_OsmL041d6_1(.din(w_dff_B_E7GihjsA6_1),.dout(w_dff_B_OsmL041d6_1),.clk(gclk));
	jdff dff_B_H0AYqXlV5_1(.din(w_dff_B_OsmL041d6_1),.dout(w_dff_B_H0AYqXlV5_1),.clk(gclk));
	jdff dff_B_AqCS8Wmr0_1(.din(w_dff_B_H0AYqXlV5_1),.dout(w_dff_B_AqCS8Wmr0_1),.clk(gclk));
	jdff dff_B_5E5N8fbG7_1(.din(w_dff_B_AqCS8Wmr0_1),.dout(w_dff_B_5E5N8fbG7_1),.clk(gclk));
	jdff dff_B_mbyGOUyK7_1(.din(w_dff_B_5E5N8fbG7_1),.dout(w_dff_B_mbyGOUyK7_1),.clk(gclk));
	jdff dff_B_NE2Esbso4_1(.din(w_dff_B_mbyGOUyK7_1),.dout(w_dff_B_NE2Esbso4_1),.clk(gclk));
	jdff dff_B_hKZQVC1B9_1(.din(w_dff_B_NE2Esbso4_1),.dout(w_dff_B_hKZQVC1B9_1),.clk(gclk));
	jdff dff_B_OaZI88vZ2_1(.din(w_dff_B_hKZQVC1B9_1),.dout(w_dff_B_OaZI88vZ2_1),.clk(gclk));
	jdff dff_B_QS0AaBq25_1(.din(w_dff_B_OaZI88vZ2_1),.dout(w_dff_B_QS0AaBq25_1),.clk(gclk));
	jdff dff_B_nR662HS23_1(.din(w_dff_B_QS0AaBq25_1),.dout(w_dff_B_nR662HS23_1),.clk(gclk));
	jdff dff_B_fCejSuMv7_1(.din(w_dff_B_nR662HS23_1),.dout(w_dff_B_fCejSuMv7_1),.clk(gclk));
	jdff dff_B_fAWzTRaQ1_1(.din(w_dff_B_fCejSuMv7_1),.dout(w_dff_B_fAWzTRaQ1_1),.clk(gclk));
	jdff dff_B_yOrbzuPC5_1(.din(w_dff_B_fAWzTRaQ1_1),.dout(w_dff_B_yOrbzuPC5_1),.clk(gclk));
	jdff dff_B_pzsHEBWb6_1(.din(w_dff_B_yOrbzuPC5_1),.dout(w_dff_B_pzsHEBWb6_1),.clk(gclk));
	jdff dff_B_Zn469Bwc7_1(.din(w_dff_B_pzsHEBWb6_1),.dout(w_dff_B_Zn469Bwc7_1),.clk(gclk));
	jdff dff_B_VLtRZy4v3_1(.din(w_dff_B_Zn469Bwc7_1),.dout(w_dff_B_VLtRZy4v3_1),.clk(gclk));
	jdff dff_B_ptQ25fex8_1(.din(w_dff_B_VLtRZy4v3_1),.dout(w_dff_B_ptQ25fex8_1),.clk(gclk));
	jdff dff_B_jVX8F6Xl3_1(.din(w_dff_B_ptQ25fex8_1),.dout(w_dff_B_jVX8F6Xl3_1),.clk(gclk));
	jdff dff_B_CawEFLW32_1(.din(w_dff_B_jVX8F6Xl3_1),.dout(w_dff_B_CawEFLW32_1),.clk(gclk));
	jdff dff_B_6Uk0kY1J5_1(.din(w_dff_B_CawEFLW32_1),.dout(w_dff_B_6Uk0kY1J5_1),.clk(gclk));
	jdff dff_B_bbrhRmbf2_1(.din(w_dff_B_6Uk0kY1J5_1),.dout(w_dff_B_bbrhRmbf2_1),.clk(gclk));
	jdff dff_B_Z3OEavTf6_1(.din(w_dff_B_bbrhRmbf2_1),.dout(w_dff_B_Z3OEavTf6_1),.clk(gclk));
	jdff dff_B_igpowbij3_1(.din(w_dff_B_Z3OEavTf6_1),.dout(w_dff_B_igpowbij3_1),.clk(gclk));
	jdff dff_B_olWfDcaN6_1(.din(w_dff_B_igpowbij3_1),.dout(w_dff_B_olWfDcaN6_1),.clk(gclk));
	jdff dff_B_YXhLdMks0_1(.din(w_dff_B_olWfDcaN6_1),.dout(w_dff_B_YXhLdMks0_1),.clk(gclk));
	jdff dff_B_NQAj0qbZ9_1(.din(w_dff_B_YXhLdMks0_1),.dout(w_dff_B_NQAj0qbZ9_1),.clk(gclk));
	jdff dff_B_ngqDtuqD7_1(.din(w_dff_B_NQAj0qbZ9_1),.dout(w_dff_B_ngqDtuqD7_1),.clk(gclk));
	jdff dff_B_kNPbp8J69_1(.din(w_dff_B_ngqDtuqD7_1),.dout(w_dff_B_kNPbp8J69_1),.clk(gclk));
	jdff dff_B_8VV8Qc1M7_1(.din(w_dff_B_kNPbp8J69_1),.dout(w_dff_B_8VV8Qc1M7_1),.clk(gclk));
	jdff dff_B_ttafBy0w3_1(.din(w_dff_B_8VV8Qc1M7_1),.dout(w_dff_B_ttafBy0w3_1),.clk(gclk));
	jdff dff_B_bHVB0p1Z3_1(.din(w_dff_B_ttafBy0w3_1),.dout(w_dff_B_bHVB0p1Z3_1),.clk(gclk));
	jdff dff_B_AiGyld9I4_1(.din(w_dff_B_bHVB0p1Z3_1),.dout(w_dff_B_AiGyld9I4_1),.clk(gclk));
	jdff dff_B_6y3Mt8UG5_1(.din(w_dff_B_AiGyld9I4_1),.dout(w_dff_B_6y3Mt8UG5_1),.clk(gclk));
	jdff dff_B_z8w0zcKB8_0(.din(n1296),.dout(w_dff_B_z8w0zcKB8_0),.clk(gclk));
	jdff dff_B_hV2wI3hE3_1(.din(n1811),.dout(w_dff_B_hV2wI3hE3_1),.clk(gclk));
	jdff dff_B_tPuf6rMo7_1(.din(w_dff_B_hV2wI3hE3_1),.dout(w_dff_B_tPuf6rMo7_1),.clk(gclk));
	jdff dff_B_NK12tZbp3_1(.din(w_dff_B_tPuf6rMo7_1),.dout(w_dff_B_NK12tZbp3_1),.clk(gclk));
	jdff dff_B_SKk71p9z7_1(.din(w_dff_B_NK12tZbp3_1),.dout(w_dff_B_SKk71p9z7_1),.clk(gclk));
	jdff dff_B_GiwqYT4t5_1(.din(w_dff_B_SKk71p9z7_1),.dout(w_dff_B_GiwqYT4t5_1),.clk(gclk));
	jdff dff_B_gzxu1Q299_1(.din(w_dff_B_GiwqYT4t5_1),.dout(w_dff_B_gzxu1Q299_1),.clk(gclk));
	jdff dff_B_7eVcSRTQ8_1(.din(w_dff_B_gzxu1Q299_1),.dout(w_dff_B_7eVcSRTQ8_1),.clk(gclk));
	jdff dff_B_DQvoTz455_1(.din(w_dff_B_7eVcSRTQ8_1),.dout(w_dff_B_DQvoTz455_1),.clk(gclk));
	jdff dff_B_6cc3BkZ72_1(.din(w_dff_B_DQvoTz455_1),.dout(w_dff_B_6cc3BkZ72_1),.clk(gclk));
	jdff dff_B_IkXUt7xC5_1(.din(w_dff_B_6cc3BkZ72_1),.dout(w_dff_B_IkXUt7xC5_1),.clk(gclk));
	jdff dff_B_B10s512I5_1(.din(w_dff_B_IkXUt7xC5_1),.dout(w_dff_B_B10s512I5_1),.clk(gclk));
	jdff dff_B_US89lrvl8_1(.din(w_dff_B_B10s512I5_1),.dout(w_dff_B_US89lrvl8_1),.clk(gclk));
	jdff dff_B_hSmZqu2u0_1(.din(w_dff_B_US89lrvl8_1),.dout(w_dff_B_hSmZqu2u0_1),.clk(gclk));
	jdff dff_B_bJ7asy1c2_1(.din(w_dff_B_hSmZqu2u0_1),.dout(w_dff_B_bJ7asy1c2_1),.clk(gclk));
	jdff dff_B_huyM6Sbm7_1(.din(w_dff_B_bJ7asy1c2_1),.dout(w_dff_B_huyM6Sbm7_1),.clk(gclk));
	jdff dff_B_Zzjqdy094_0(.din(n1819),.dout(w_dff_B_Zzjqdy094_0),.clk(gclk));
	jdff dff_B_Lx8y4Qgd1_0(.din(w_dff_B_Zzjqdy094_0),.dout(w_dff_B_Lx8y4Qgd1_0),.clk(gclk));
	jdff dff_B_n1DYH6Eu0_0(.din(w_dff_B_Lx8y4Qgd1_0),.dout(w_dff_B_n1DYH6Eu0_0),.clk(gclk));
	jdff dff_B_BbkwgzEX7_0(.din(w_dff_B_n1DYH6Eu0_0),.dout(w_dff_B_BbkwgzEX7_0),.clk(gclk));
	jdff dff_B_AnWxIQvn7_0(.din(w_dff_B_BbkwgzEX7_0),.dout(w_dff_B_AnWxIQvn7_0),.clk(gclk));
	jdff dff_B_Cu2zUTVv4_0(.din(w_dff_B_AnWxIQvn7_0),.dout(w_dff_B_Cu2zUTVv4_0),.clk(gclk));
	jdff dff_B_fCzsxwc23_0(.din(w_dff_B_Cu2zUTVv4_0),.dout(w_dff_B_fCzsxwc23_0),.clk(gclk));
	jdff dff_B_hC0stYPe2_0(.din(w_dff_B_fCzsxwc23_0),.dout(w_dff_B_hC0stYPe2_0),.clk(gclk));
	jdff dff_B_xDjbwjZR5_0(.din(w_dff_B_hC0stYPe2_0),.dout(w_dff_B_xDjbwjZR5_0),.clk(gclk));
	jdff dff_B_22CDTs6g3_0(.din(w_dff_B_xDjbwjZR5_0),.dout(w_dff_B_22CDTs6g3_0),.clk(gclk));
	jdff dff_B_y0h7Pa8r2_0(.din(w_dff_B_22CDTs6g3_0),.dout(w_dff_B_y0h7Pa8r2_0),.clk(gclk));
	jdff dff_B_nUH4L31U6_0(.din(w_dff_B_y0h7Pa8r2_0),.dout(w_dff_B_nUH4L31U6_0),.clk(gclk));
	jdff dff_B_sQArDvcX8_0(.din(w_dff_B_nUH4L31U6_0),.dout(w_dff_B_sQArDvcX8_0),.clk(gclk));
	jdff dff_A_zNSE46Vu5_0(.dout(w_n1818_0[0]),.din(w_dff_A_zNSE46Vu5_0),.clk(gclk));
	jdff dff_A_V2Fsx7BU9_0(.dout(w_dff_A_zNSE46Vu5_0),.din(w_dff_A_V2Fsx7BU9_0),.clk(gclk));
	jdff dff_A_bvULOijl7_0(.dout(w_dff_A_V2Fsx7BU9_0),.din(w_dff_A_bvULOijl7_0),.clk(gclk));
	jdff dff_A_YY2plMGm3_0(.dout(w_dff_A_bvULOijl7_0),.din(w_dff_A_YY2plMGm3_0),.clk(gclk));
	jdff dff_A_ccwjmVMm4_0(.dout(w_dff_A_YY2plMGm3_0),.din(w_dff_A_ccwjmVMm4_0),.clk(gclk));
	jdff dff_A_AmWwTINm2_0(.dout(w_dff_A_ccwjmVMm4_0),.din(w_dff_A_AmWwTINm2_0),.clk(gclk));
	jdff dff_A_jj2KitXd6_0(.dout(w_dff_A_AmWwTINm2_0),.din(w_dff_A_jj2KitXd6_0),.clk(gclk));
	jdff dff_A_0QE3QVJE9_0(.dout(w_dff_A_jj2KitXd6_0),.din(w_dff_A_0QE3QVJE9_0),.clk(gclk));
	jdff dff_A_rZ7ONRVB7_0(.dout(w_dff_A_0QE3QVJE9_0),.din(w_dff_A_rZ7ONRVB7_0),.clk(gclk));
	jdff dff_A_WEIV3QYS9_0(.dout(w_dff_A_rZ7ONRVB7_0),.din(w_dff_A_WEIV3QYS9_0),.clk(gclk));
	jdff dff_A_rErx2SLH9_0(.dout(w_dff_A_WEIV3QYS9_0),.din(w_dff_A_rErx2SLH9_0),.clk(gclk));
	jdff dff_A_gxGqzSXs2_0(.dout(w_dff_A_rErx2SLH9_0),.din(w_dff_A_gxGqzSXs2_0),.clk(gclk));
	jdff dff_A_pgjsqp0w8_0(.dout(w_dff_A_gxGqzSXs2_0),.din(w_dff_A_pgjsqp0w8_0),.clk(gclk));
	jdff dff_A_L8ueDPvO2_0(.dout(w_dff_A_pgjsqp0w8_0),.din(w_dff_A_L8ueDPvO2_0),.clk(gclk));
	jdff dff_B_CwRSeIak2_1(.din(n1808),.dout(w_dff_B_CwRSeIak2_1),.clk(gclk));
	jdff dff_B_JdEVAEq01_1(.din(w_dff_B_CwRSeIak2_1),.dout(w_dff_B_JdEVAEq01_1),.clk(gclk));
	jdff dff_B_9c9ST8518_2(.din(n1807),.dout(w_dff_B_9c9ST8518_2),.clk(gclk));
	jdff dff_B_MdcDDMGE5_2(.din(w_dff_B_9c9ST8518_2),.dout(w_dff_B_MdcDDMGE5_2),.clk(gclk));
	jdff dff_B_oGKanOkl0_2(.din(w_dff_B_MdcDDMGE5_2),.dout(w_dff_B_oGKanOkl0_2),.clk(gclk));
	jdff dff_B_NgeIEH9P2_2(.din(w_dff_B_oGKanOkl0_2),.dout(w_dff_B_NgeIEH9P2_2),.clk(gclk));
	jdff dff_B_DzNTginG5_2(.din(w_dff_B_NgeIEH9P2_2),.dout(w_dff_B_DzNTginG5_2),.clk(gclk));
	jdff dff_B_eKoW9Bcr7_2(.din(w_dff_B_DzNTginG5_2),.dout(w_dff_B_eKoW9Bcr7_2),.clk(gclk));
	jdff dff_B_xKfx4z0l9_2(.din(w_dff_B_eKoW9Bcr7_2),.dout(w_dff_B_xKfx4z0l9_2),.clk(gclk));
	jdff dff_B_47pJCbFJ9_2(.din(w_dff_B_xKfx4z0l9_2),.dout(w_dff_B_47pJCbFJ9_2),.clk(gclk));
	jdff dff_B_md9S7CLo4_2(.din(w_dff_B_47pJCbFJ9_2),.dout(w_dff_B_md9S7CLo4_2),.clk(gclk));
	jdff dff_B_Wug8SRLh9_2(.din(w_dff_B_md9S7CLo4_2),.dout(w_dff_B_Wug8SRLh9_2),.clk(gclk));
	jdff dff_B_c5thFNV69_2(.din(w_dff_B_Wug8SRLh9_2),.dout(w_dff_B_c5thFNV69_2),.clk(gclk));
	jdff dff_B_avL0NWVT2_2(.din(w_dff_B_c5thFNV69_2),.dout(w_dff_B_avL0NWVT2_2),.clk(gclk));
	jdff dff_B_yldM4uHr4_2(.din(w_dff_B_avL0NWVT2_2),.dout(w_dff_B_yldM4uHr4_2),.clk(gclk));
	jdff dff_B_yyCtVycQ4_2(.din(w_dff_B_yldM4uHr4_2),.dout(w_dff_B_yyCtVycQ4_2),.clk(gclk));
	jdff dff_B_Fb5PdAwy2_2(.din(w_dff_B_yyCtVycQ4_2),.dout(w_dff_B_Fb5PdAwy2_2),.clk(gclk));
	jdff dff_B_4XwPFce52_2(.din(w_dff_B_Fb5PdAwy2_2),.dout(w_dff_B_4XwPFce52_2),.clk(gclk));
	jdff dff_B_SPLC5CPS6_2(.din(w_dff_B_4XwPFce52_2),.dout(w_dff_B_SPLC5CPS6_2),.clk(gclk));
	jdff dff_B_HaKW4JTM6_2(.din(w_dff_B_SPLC5CPS6_2),.dout(w_dff_B_HaKW4JTM6_2),.clk(gclk));
	jdff dff_B_88C9hQyN6_2(.din(w_dff_B_HaKW4JTM6_2),.dout(w_dff_B_88C9hQyN6_2),.clk(gclk));
	jdff dff_B_gda2oCd96_2(.din(w_dff_B_88C9hQyN6_2),.dout(w_dff_B_gda2oCd96_2),.clk(gclk));
	jdff dff_B_QoPMMl6n7_2(.din(w_dff_B_gda2oCd96_2),.dout(w_dff_B_QoPMMl6n7_2),.clk(gclk));
	jdff dff_B_1DjAqkbo8_2(.din(w_dff_B_QoPMMl6n7_2),.dout(w_dff_B_1DjAqkbo8_2),.clk(gclk));
	jdff dff_B_EaUyJfyk4_2(.din(w_dff_B_1DjAqkbo8_2),.dout(w_dff_B_EaUyJfyk4_2),.clk(gclk));
	jdff dff_B_4p0V0LEh8_2(.din(w_dff_B_EaUyJfyk4_2),.dout(w_dff_B_4p0V0LEh8_2),.clk(gclk));
	jdff dff_B_GwtcKxKR3_2(.din(w_dff_B_4p0V0LEh8_2),.dout(w_dff_B_GwtcKxKR3_2),.clk(gclk));
	jdff dff_B_8dBBk3Rk7_2(.din(w_dff_B_GwtcKxKR3_2),.dout(w_dff_B_8dBBk3Rk7_2),.clk(gclk));
	jdff dff_B_PMIi69VZ4_2(.din(w_dff_B_8dBBk3Rk7_2),.dout(w_dff_B_PMIi69VZ4_2),.clk(gclk));
	jdff dff_B_GMkvc1yV0_2(.din(w_dff_B_PMIi69VZ4_2),.dout(w_dff_B_GMkvc1yV0_2),.clk(gclk));
	jdff dff_B_jO2yocm39_2(.din(w_dff_B_GMkvc1yV0_2),.dout(w_dff_B_jO2yocm39_2),.clk(gclk));
	jdff dff_B_Tv2aRw1p4_2(.din(w_dff_B_jO2yocm39_2),.dout(w_dff_B_Tv2aRw1p4_2),.clk(gclk));
	jdff dff_B_6g1LHoz31_2(.din(w_dff_B_Tv2aRw1p4_2),.dout(w_dff_B_6g1LHoz31_2),.clk(gclk));
	jdff dff_B_dEqZoGSd7_2(.din(w_dff_B_6g1LHoz31_2),.dout(w_dff_B_dEqZoGSd7_2),.clk(gclk));
	jdff dff_B_hQI3iIFS4_2(.din(w_dff_B_dEqZoGSd7_2),.dout(w_dff_B_hQI3iIFS4_2),.clk(gclk));
	jdff dff_B_WO3SNvig4_2(.din(w_dff_B_hQI3iIFS4_2),.dout(w_dff_B_WO3SNvig4_2),.clk(gclk));
	jdff dff_B_p620AGEX3_2(.din(w_dff_B_WO3SNvig4_2),.dout(w_dff_B_p620AGEX3_2),.clk(gclk));
	jdff dff_B_UDwP52Ud7_2(.din(w_dff_B_p620AGEX3_2),.dout(w_dff_B_UDwP52Ud7_2),.clk(gclk));
	jdff dff_B_wsO7XN0l8_2(.din(w_dff_B_UDwP52Ud7_2),.dout(w_dff_B_wsO7XN0l8_2),.clk(gclk));
	jdff dff_B_TSTtLijB6_2(.din(w_dff_B_wsO7XN0l8_2),.dout(w_dff_B_TSTtLijB6_2),.clk(gclk));
	jdff dff_B_ijDm1qaW2_2(.din(w_dff_B_TSTtLijB6_2),.dout(w_dff_B_ijDm1qaW2_2),.clk(gclk));
	jdff dff_B_0EXD4U4H2_2(.din(w_dff_B_ijDm1qaW2_2),.dout(w_dff_B_0EXD4U4H2_2),.clk(gclk));
	jdff dff_B_ia58TNRU7_2(.din(w_dff_B_0EXD4U4H2_2),.dout(w_dff_B_ia58TNRU7_2),.clk(gclk));
	jdff dff_B_xNE0itga9_2(.din(w_dff_B_ia58TNRU7_2),.dout(w_dff_B_xNE0itga9_2),.clk(gclk));
	jdff dff_B_KIGMbyhU2_2(.din(w_dff_B_xNE0itga9_2),.dout(w_dff_B_KIGMbyhU2_2),.clk(gclk));
	jdff dff_B_TrggROkz2_2(.din(w_dff_B_KIGMbyhU2_2),.dout(w_dff_B_TrggROkz2_2),.clk(gclk));
	jdff dff_B_mPZEw0Sx3_2(.din(w_dff_B_TrggROkz2_2),.dout(w_dff_B_mPZEw0Sx3_2),.clk(gclk));
	jdff dff_B_2wUTUvBm1_2(.din(w_dff_B_mPZEw0Sx3_2),.dout(w_dff_B_2wUTUvBm1_2),.clk(gclk));
	jdff dff_B_Zbsd94kw5_2(.din(w_dff_B_2wUTUvBm1_2),.dout(w_dff_B_Zbsd94kw5_2),.clk(gclk));
	jdff dff_B_qUOymOHe4_2(.din(w_dff_B_Zbsd94kw5_2),.dout(w_dff_B_qUOymOHe4_2),.clk(gclk));
	jdff dff_B_bPgX9GmS9_2(.din(w_dff_B_qUOymOHe4_2),.dout(w_dff_B_bPgX9GmS9_2),.clk(gclk));
	jdff dff_B_9eiVS16e5_2(.din(w_dff_B_bPgX9GmS9_2),.dout(w_dff_B_9eiVS16e5_2),.clk(gclk));
	jdff dff_B_gdKuuyar9_2(.din(w_dff_B_9eiVS16e5_2),.dout(w_dff_B_gdKuuyar9_2),.clk(gclk));
	jdff dff_B_iT1HOUD15_2(.din(w_dff_B_gdKuuyar9_2),.dout(w_dff_B_iT1HOUD15_2),.clk(gclk));
	jdff dff_B_pls9ok3V1_2(.din(w_dff_B_iT1HOUD15_2),.dout(w_dff_B_pls9ok3V1_2),.clk(gclk));
	jdff dff_B_Ao8U18wJ8_2(.din(w_dff_B_pls9ok3V1_2),.dout(w_dff_B_Ao8U18wJ8_2),.clk(gclk));
	jdff dff_B_vA60CrKa1_2(.din(w_dff_B_Ao8U18wJ8_2),.dout(w_dff_B_vA60CrKa1_2),.clk(gclk));
	jdff dff_B_ulT9deez7_2(.din(w_dff_B_vA60CrKa1_2),.dout(w_dff_B_ulT9deez7_2),.clk(gclk));
	jdff dff_B_TnNJYkFP3_2(.din(w_dff_B_ulT9deez7_2),.dout(w_dff_B_TnNJYkFP3_2),.clk(gclk));
	jdff dff_B_7cLve7654_1(.din(n1814),.dout(w_dff_B_7cLve7654_1),.clk(gclk));
	jdff dff_B_B7AqmFwC0_1(.din(w_dff_B_7cLve7654_1),.dout(w_dff_B_B7AqmFwC0_1),.clk(gclk));
	jdff dff_B_ZBDtyjBf7_1(.din(w_dff_B_B7AqmFwC0_1),.dout(w_dff_B_ZBDtyjBf7_1),.clk(gclk));
	jdff dff_B_nfKhVY6U7_1(.din(w_dff_B_ZBDtyjBf7_1),.dout(w_dff_B_nfKhVY6U7_1),.clk(gclk));
	jdff dff_B_s2zwTIMK9_1(.din(w_dff_B_nfKhVY6U7_1),.dout(w_dff_B_s2zwTIMK9_1),.clk(gclk));
	jdff dff_B_fH90MPwb5_1(.din(w_dff_B_s2zwTIMK9_1),.dout(w_dff_B_fH90MPwb5_1),.clk(gclk));
	jdff dff_B_yYdbQXdC5_1(.din(w_dff_B_fH90MPwb5_1),.dout(w_dff_B_yYdbQXdC5_1),.clk(gclk));
	jdff dff_B_kcXlAPcu8_1(.din(w_dff_B_yYdbQXdC5_1),.dout(w_dff_B_kcXlAPcu8_1),.clk(gclk));
	jdff dff_B_hl3AyHsE8_1(.din(w_dff_B_kcXlAPcu8_1),.dout(w_dff_B_hl3AyHsE8_1),.clk(gclk));
	jdff dff_B_lViDSS2w3_1(.din(w_dff_B_hl3AyHsE8_1),.dout(w_dff_B_lViDSS2w3_1),.clk(gclk));
	jdff dff_B_TIDP2gBH7_1(.din(w_dff_B_lViDSS2w3_1),.dout(w_dff_B_TIDP2gBH7_1),.clk(gclk));
	jdff dff_B_Jif6Ryib0_1(.din(w_dff_B_TIDP2gBH7_1),.dout(w_dff_B_Jif6Ryib0_1),.clk(gclk));
	jdff dff_B_rKvz3qNj9_1(.din(w_dff_B_Jif6Ryib0_1),.dout(w_dff_B_rKvz3qNj9_1),.clk(gclk));
	jdff dff_B_NTsVBm794_0(.din(n1815),.dout(w_dff_B_NTsVBm794_0),.clk(gclk));
	jdff dff_B_X3m0Mhqr1_0(.din(w_dff_B_NTsVBm794_0),.dout(w_dff_B_X3m0Mhqr1_0),.clk(gclk));
	jdff dff_B_JJsjNdCn2_0(.din(w_dff_B_X3m0Mhqr1_0),.dout(w_dff_B_JJsjNdCn2_0),.clk(gclk));
	jdff dff_B_xpjB9u8B6_0(.din(w_dff_B_JJsjNdCn2_0),.dout(w_dff_B_xpjB9u8B6_0),.clk(gclk));
	jdff dff_B_fMFD8vZA7_0(.din(w_dff_B_xpjB9u8B6_0),.dout(w_dff_B_fMFD8vZA7_0),.clk(gclk));
	jdff dff_B_XbszIEMB1_0(.din(w_dff_B_fMFD8vZA7_0),.dout(w_dff_B_XbszIEMB1_0),.clk(gclk));
	jdff dff_B_pdpPE8Ce2_0(.din(w_dff_B_XbszIEMB1_0),.dout(w_dff_B_pdpPE8Ce2_0),.clk(gclk));
	jdff dff_B_uFpunoN25_0(.din(w_dff_B_pdpPE8Ce2_0),.dout(w_dff_B_uFpunoN25_0),.clk(gclk));
	jdff dff_B_Bz1ltoA82_0(.din(w_dff_B_uFpunoN25_0),.dout(w_dff_B_Bz1ltoA82_0),.clk(gclk));
	jdff dff_B_1vNNiMQ23_0(.din(w_dff_B_Bz1ltoA82_0),.dout(w_dff_B_1vNNiMQ23_0),.clk(gclk));
	jdff dff_B_oT7xWidf7_0(.din(w_dff_B_1vNNiMQ23_0),.dout(w_dff_B_oT7xWidf7_0),.clk(gclk));
	jdff dff_B_uG0G052K0_0(.din(w_dff_B_oT7xWidf7_0),.dout(w_dff_B_uG0G052K0_0),.clk(gclk));
	jdff dff_A_WPGvsqm03_1(.dout(w_n1805_0[1]),.din(w_dff_A_WPGvsqm03_1),.clk(gclk));
	jdff dff_A_hETNtujh0_1(.dout(w_dff_A_WPGvsqm03_1),.din(w_dff_A_hETNtujh0_1),.clk(gclk));
	jdff dff_A_78BxAME50_1(.dout(w_dff_A_hETNtujh0_1),.din(w_dff_A_78BxAME50_1),.clk(gclk));
	jdff dff_A_KFoJGfPx5_1(.dout(w_dff_A_78BxAME50_1),.din(w_dff_A_KFoJGfPx5_1),.clk(gclk));
	jdff dff_A_TzyQriov7_1(.dout(w_dff_A_KFoJGfPx5_1),.din(w_dff_A_TzyQriov7_1),.clk(gclk));
	jdff dff_A_SczVSiE31_1(.dout(w_dff_A_TzyQriov7_1),.din(w_dff_A_SczVSiE31_1),.clk(gclk));
	jdff dff_A_DqlTu6MF6_1(.dout(w_dff_A_SczVSiE31_1),.din(w_dff_A_DqlTu6MF6_1),.clk(gclk));
	jdff dff_A_MSz7eijY0_1(.dout(w_dff_A_DqlTu6MF6_1),.din(w_dff_A_MSz7eijY0_1),.clk(gclk));
	jdff dff_A_yQFGxJ9h3_1(.dout(w_dff_A_MSz7eijY0_1),.din(w_dff_A_yQFGxJ9h3_1),.clk(gclk));
	jdff dff_A_Mgt8YJNu3_1(.dout(w_dff_A_yQFGxJ9h3_1),.din(w_dff_A_Mgt8YJNu3_1),.clk(gclk));
	jdff dff_A_hP7rHZ7F3_1(.dout(w_dff_A_Mgt8YJNu3_1),.din(w_dff_A_hP7rHZ7F3_1),.clk(gclk));
	jdff dff_A_rstKqXmV5_1(.dout(w_dff_A_hP7rHZ7F3_1),.din(w_dff_A_rstKqXmV5_1),.clk(gclk));
	jdff dff_A_bKLg2vTL0_1(.dout(w_dff_A_rstKqXmV5_1),.din(w_dff_A_bKLg2vTL0_1),.clk(gclk));
	jdff dff_B_YmazJ7807_1(.din(n1790),.dout(w_dff_B_YmazJ7807_1),.clk(gclk));
	jdff dff_B_bGUZDYX04_1(.din(w_dff_B_YmazJ7807_1),.dout(w_dff_B_bGUZDYX04_1),.clk(gclk));
	jdff dff_B_LjhZY2LC8_1(.din(w_dff_B_bGUZDYX04_1),.dout(w_dff_B_LjhZY2LC8_1),.clk(gclk));
	jdff dff_B_LrYV5Ntu7_1(.din(w_dff_B_LjhZY2LC8_1),.dout(w_dff_B_LrYV5Ntu7_1),.clk(gclk));
	jdff dff_B_oawRA7Kw5_1(.din(w_dff_B_LrYV5Ntu7_1),.dout(w_dff_B_oawRA7Kw5_1),.clk(gclk));
	jdff dff_B_8vfzK27C1_1(.din(w_dff_B_oawRA7Kw5_1),.dout(w_dff_B_8vfzK27C1_1),.clk(gclk));
	jdff dff_B_aKUpKm3y4_1(.din(w_dff_B_8vfzK27C1_1),.dout(w_dff_B_aKUpKm3y4_1),.clk(gclk));
	jdff dff_B_RFLUSRNx9_1(.din(w_dff_B_aKUpKm3y4_1),.dout(w_dff_B_RFLUSRNx9_1),.clk(gclk));
	jdff dff_B_iDbRK6Ty8_1(.din(w_dff_B_RFLUSRNx9_1),.dout(w_dff_B_iDbRK6Ty8_1),.clk(gclk));
	jdff dff_B_ix4VJOmh3_1(.din(w_dff_B_iDbRK6Ty8_1),.dout(w_dff_B_ix4VJOmh3_1),.clk(gclk));
	jdff dff_B_JpgOkr6L9_1(.din(w_dff_B_ix4VJOmh3_1),.dout(w_dff_B_JpgOkr6L9_1),.clk(gclk));
	jdff dff_B_mwwiw5lE1_1(.din(w_dff_B_JpgOkr6L9_1),.dout(w_dff_B_mwwiw5lE1_1),.clk(gclk));
	jdff dff_B_yRWuqKkw5_1(.din(w_dff_B_mwwiw5lE1_1),.dout(w_dff_B_yRWuqKkw5_1),.clk(gclk));
	jdff dff_B_GnbcdT6s3_0(.din(n1791),.dout(w_dff_B_GnbcdT6s3_0),.clk(gclk));
	jdff dff_B_PQTROi1O5_0(.din(w_dff_B_GnbcdT6s3_0),.dout(w_dff_B_PQTROi1O5_0),.clk(gclk));
	jdff dff_B_fXrwwZH15_0(.din(w_dff_B_PQTROi1O5_0),.dout(w_dff_B_fXrwwZH15_0),.clk(gclk));
	jdff dff_B_2Mux3wgO2_0(.din(w_dff_B_fXrwwZH15_0),.dout(w_dff_B_2Mux3wgO2_0),.clk(gclk));
	jdff dff_B_pwpySj0Q4_0(.din(w_dff_B_2Mux3wgO2_0),.dout(w_dff_B_pwpySj0Q4_0),.clk(gclk));
	jdff dff_B_Ys9Lr5Gk2_0(.din(w_dff_B_pwpySj0Q4_0),.dout(w_dff_B_Ys9Lr5Gk2_0),.clk(gclk));
	jdff dff_B_YKptjCab5_0(.din(w_dff_B_Ys9Lr5Gk2_0),.dout(w_dff_B_YKptjCab5_0),.clk(gclk));
	jdff dff_B_8sy3xX1L0_0(.din(w_dff_B_YKptjCab5_0),.dout(w_dff_B_8sy3xX1L0_0),.clk(gclk));
	jdff dff_B_7XPHU3ij2_0(.din(w_dff_B_8sy3xX1L0_0),.dout(w_dff_B_7XPHU3ij2_0),.clk(gclk));
	jdff dff_B_6MQAk3Jk8_0(.din(w_dff_B_7XPHU3ij2_0),.dout(w_dff_B_6MQAk3Jk8_0),.clk(gclk));
	jdff dff_B_Ue28N7Wt2_0(.din(w_dff_B_6MQAk3Jk8_0),.dout(w_dff_B_Ue28N7Wt2_0),.clk(gclk));
	jdff dff_B_ZeYPt54T0_0(.din(w_dff_B_Ue28N7Wt2_0),.dout(w_dff_B_ZeYPt54T0_0),.clk(gclk));
	jdff dff_A_DRe20etP5_1(.dout(w_n1786_0[1]),.din(w_dff_A_DRe20etP5_1),.clk(gclk));
	jdff dff_A_Payo0NRM4_1(.dout(w_dff_A_DRe20etP5_1),.din(w_dff_A_Payo0NRM4_1),.clk(gclk));
	jdff dff_A_NCnB7HKx1_1(.dout(w_dff_A_Payo0NRM4_1),.din(w_dff_A_NCnB7HKx1_1),.clk(gclk));
	jdff dff_A_xtky17vQ9_1(.dout(w_dff_A_NCnB7HKx1_1),.din(w_dff_A_xtky17vQ9_1),.clk(gclk));
	jdff dff_A_76v08Zms2_1(.dout(w_dff_A_xtky17vQ9_1),.din(w_dff_A_76v08Zms2_1),.clk(gclk));
	jdff dff_A_GHVd2Zyw9_1(.dout(w_dff_A_76v08Zms2_1),.din(w_dff_A_GHVd2Zyw9_1),.clk(gclk));
	jdff dff_A_J7RdBkdz0_1(.dout(w_dff_A_GHVd2Zyw9_1),.din(w_dff_A_J7RdBkdz0_1),.clk(gclk));
	jdff dff_A_r3anLi1b9_1(.dout(w_dff_A_J7RdBkdz0_1),.din(w_dff_A_r3anLi1b9_1),.clk(gclk));
	jdff dff_A_1l4xKHte9_1(.dout(w_dff_A_r3anLi1b9_1),.din(w_dff_A_1l4xKHte9_1),.clk(gclk));
	jdff dff_A_BzNfuLlh3_1(.dout(w_dff_A_1l4xKHte9_1),.din(w_dff_A_BzNfuLlh3_1),.clk(gclk));
	jdff dff_A_9SNYp1wM0_1(.dout(w_dff_A_BzNfuLlh3_1),.din(w_dff_A_9SNYp1wM0_1),.clk(gclk));
	jdff dff_A_Rjsuyn4I3_1(.dout(w_dff_A_9SNYp1wM0_1),.din(w_dff_A_Rjsuyn4I3_1),.clk(gclk));
	jdff dff_A_7qFQCJai5_1(.dout(w_dff_A_Rjsuyn4I3_1),.din(w_dff_A_7qFQCJai5_1),.clk(gclk));
	jdff dff_B_eNlUkgVG5_1(.din(n1764),.dout(w_dff_B_eNlUkgVG5_1),.clk(gclk));
	jdff dff_B_YWAHMO8q9_1(.din(w_dff_B_eNlUkgVG5_1),.dout(w_dff_B_YWAHMO8q9_1),.clk(gclk));
	jdff dff_B_dtiGdofG0_1(.din(w_dff_B_YWAHMO8q9_1),.dout(w_dff_B_dtiGdofG0_1),.clk(gclk));
	jdff dff_B_4duU7BmE7_1(.din(w_dff_B_dtiGdofG0_1),.dout(w_dff_B_4duU7BmE7_1),.clk(gclk));
	jdff dff_B_Z8govWyO5_1(.din(w_dff_B_4duU7BmE7_1),.dout(w_dff_B_Z8govWyO5_1),.clk(gclk));
	jdff dff_B_HzdqHQ8b1_1(.din(w_dff_B_Z8govWyO5_1),.dout(w_dff_B_HzdqHQ8b1_1),.clk(gclk));
	jdff dff_B_49hZUSiv5_1(.din(w_dff_B_HzdqHQ8b1_1),.dout(w_dff_B_49hZUSiv5_1),.clk(gclk));
	jdff dff_B_yBNeNkrt9_1(.din(w_dff_B_49hZUSiv5_1),.dout(w_dff_B_yBNeNkrt9_1),.clk(gclk));
	jdff dff_B_NV8Mmotu3_1(.din(w_dff_B_yBNeNkrt9_1),.dout(w_dff_B_NV8Mmotu3_1),.clk(gclk));
	jdff dff_B_UfNvOxqL0_1(.din(w_dff_B_NV8Mmotu3_1),.dout(w_dff_B_UfNvOxqL0_1),.clk(gclk));
	jdff dff_B_DuRBjKw84_1(.din(w_dff_B_UfNvOxqL0_1),.dout(w_dff_B_DuRBjKw84_1),.clk(gclk));
	jdff dff_B_JQXNLPIO4_1(.din(w_dff_B_DuRBjKw84_1),.dout(w_dff_B_JQXNLPIO4_1),.clk(gclk));
	jdff dff_B_7RvKsDtP2_1(.din(w_dff_B_JQXNLPIO4_1),.dout(w_dff_B_7RvKsDtP2_1),.clk(gclk));
	jdff dff_B_amPhIF7z0_0(.din(n1765),.dout(w_dff_B_amPhIF7z0_0),.clk(gclk));
	jdff dff_B_0jufnKom3_0(.din(w_dff_B_amPhIF7z0_0),.dout(w_dff_B_0jufnKom3_0),.clk(gclk));
	jdff dff_B_FhmQjCn73_0(.din(w_dff_B_0jufnKom3_0),.dout(w_dff_B_FhmQjCn73_0),.clk(gclk));
	jdff dff_B_HT2msORh7_0(.din(w_dff_B_FhmQjCn73_0),.dout(w_dff_B_HT2msORh7_0),.clk(gclk));
	jdff dff_B_RkqyehRP2_0(.din(w_dff_B_HT2msORh7_0),.dout(w_dff_B_RkqyehRP2_0),.clk(gclk));
	jdff dff_B_NSVuilWk4_0(.din(w_dff_B_RkqyehRP2_0),.dout(w_dff_B_NSVuilWk4_0),.clk(gclk));
	jdff dff_B_RNWkcmDE6_0(.din(w_dff_B_NSVuilWk4_0),.dout(w_dff_B_RNWkcmDE6_0),.clk(gclk));
	jdff dff_B_mRCXoC721_0(.din(w_dff_B_RNWkcmDE6_0),.dout(w_dff_B_mRCXoC721_0),.clk(gclk));
	jdff dff_B_P1j5d9o49_0(.din(w_dff_B_mRCXoC721_0),.dout(w_dff_B_P1j5d9o49_0),.clk(gclk));
	jdff dff_B_gmYC9GAI3_0(.din(w_dff_B_P1j5d9o49_0),.dout(w_dff_B_gmYC9GAI3_0),.clk(gclk));
	jdff dff_B_DpBUIqX74_0(.din(w_dff_B_gmYC9GAI3_0),.dout(w_dff_B_DpBUIqX74_0),.clk(gclk));
	jdff dff_B_uwUQSseo9_0(.din(w_dff_B_DpBUIqX74_0),.dout(w_dff_B_uwUQSseo9_0),.clk(gclk));
	jdff dff_A_tVT1kRa81_1(.dout(w_n1760_0[1]),.din(w_dff_A_tVT1kRa81_1),.clk(gclk));
	jdff dff_A_m27y9gzO1_1(.dout(w_dff_A_tVT1kRa81_1),.din(w_dff_A_m27y9gzO1_1),.clk(gclk));
	jdff dff_A_xd4Zz27l4_1(.dout(w_dff_A_m27y9gzO1_1),.din(w_dff_A_xd4Zz27l4_1),.clk(gclk));
	jdff dff_A_Kc73B2Dy1_1(.dout(w_dff_A_xd4Zz27l4_1),.din(w_dff_A_Kc73B2Dy1_1),.clk(gclk));
	jdff dff_A_Imk16Ha12_1(.dout(w_dff_A_Kc73B2Dy1_1),.din(w_dff_A_Imk16Ha12_1),.clk(gclk));
	jdff dff_A_rcnkaNm23_1(.dout(w_dff_A_Imk16Ha12_1),.din(w_dff_A_rcnkaNm23_1),.clk(gclk));
	jdff dff_A_iChtqyvu4_1(.dout(w_dff_A_rcnkaNm23_1),.din(w_dff_A_iChtqyvu4_1),.clk(gclk));
	jdff dff_A_ThzbdRSI1_1(.dout(w_dff_A_iChtqyvu4_1),.din(w_dff_A_ThzbdRSI1_1),.clk(gclk));
	jdff dff_A_jm8Lkqrz0_1(.dout(w_dff_A_ThzbdRSI1_1),.din(w_dff_A_jm8Lkqrz0_1),.clk(gclk));
	jdff dff_A_e6Ndbnko0_1(.dout(w_dff_A_jm8Lkqrz0_1),.din(w_dff_A_e6Ndbnko0_1),.clk(gclk));
	jdff dff_A_kMsrLRUe9_1(.dout(w_dff_A_e6Ndbnko0_1),.din(w_dff_A_kMsrLRUe9_1),.clk(gclk));
	jdff dff_A_oPgmPD5s8_1(.dout(w_dff_A_kMsrLRUe9_1),.din(w_dff_A_oPgmPD5s8_1),.clk(gclk));
	jdff dff_A_RXQQeR0j4_1(.dout(w_dff_A_oPgmPD5s8_1),.din(w_dff_A_RXQQeR0j4_1),.clk(gclk));
	jdff dff_B_Nxv2lKfY3_1(.din(n1731),.dout(w_dff_B_Nxv2lKfY3_1),.clk(gclk));
	jdff dff_B_Svgiq7dL8_1(.din(w_dff_B_Nxv2lKfY3_1),.dout(w_dff_B_Svgiq7dL8_1),.clk(gclk));
	jdff dff_B_90TNmHwt5_1(.din(w_dff_B_Svgiq7dL8_1),.dout(w_dff_B_90TNmHwt5_1),.clk(gclk));
	jdff dff_B_FrOJXGS59_1(.din(w_dff_B_90TNmHwt5_1),.dout(w_dff_B_FrOJXGS59_1),.clk(gclk));
	jdff dff_B_sxy5MF9o5_1(.din(w_dff_B_FrOJXGS59_1),.dout(w_dff_B_sxy5MF9o5_1),.clk(gclk));
	jdff dff_B_Nq6ZbYhD8_1(.din(w_dff_B_sxy5MF9o5_1),.dout(w_dff_B_Nq6ZbYhD8_1),.clk(gclk));
	jdff dff_B_hj7KsYkM8_1(.din(w_dff_B_Nq6ZbYhD8_1),.dout(w_dff_B_hj7KsYkM8_1),.clk(gclk));
	jdff dff_B_EuXoRDHk3_1(.din(w_dff_B_hj7KsYkM8_1),.dout(w_dff_B_EuXoRDHk3_1),.clk(gclk));
	jdff dff_B_SD6C0Zyb9_1(.din(w_dff_B_EuXoRDHk3_1),.dout(w_dff_B_SD6C0Zyb9_1),.clk(gclk));
	jdff dff_B_N8NeO2o61_1(.din(w_dff_B_SD6C0Zyb9_1),.dout(w_dff_B_N8NeO2o61_1),.clk(gclk));
	jdff dff_B_GRBTspeu4_1(.din(w_dff_B_N8NeO2o61_1),.dout(w_dff_B_GRBTspeu4_1),.clk(gclk));
	jdff dff_B_mLqofTnu3_1(.din(w_dff_B_GRBTspeu4_1),.dout(w_dff_B_mLqofTnu3_1),.clk(gclk));
	jdff dff_B_gEpp6YSE9_1(.din(w_dff_B_mLqofTnu3_1),.dout(w_dff_B_gEpp6YSE9_1),.clk(gclk));
	jdff dff_B_5xmx5qGV8_0(.din(n1732),.dout(w_dff_B_5xmx5qGV8_0),.clk(gclk));
	jdff dff_B_eLSVE3a04_0(.din(w_dff_B_5xmx5qGV8_0),.dout(w_dff_B_eLSVE3a04_0),.clk(gclk));
	jdff dff_B_gncrlQUf1_0(.din(w_dff_B_eLSVE3a04_0),.dout(w_dff_B_gncrlQUf1_0),.clk(gclk));
	jdff dff_B_uOqhqrZZ5_0(.din(w_dff_B_gncrlQUf1_0),.dout(w_dff_B_uOqhqrZZ5_0),.clk(gclk));
	jdff dff_B_Uh3br8OP1_0(.din(w_dff_B_uOqhqrZZ5_0),.dout(w_dff_B_Uh3br8OP1_0),.clk(gclk));
	jdff dff_B_sNHTtnzO9_0(.din(w_dff_B_Uh3br8OP1_0),.dout(w_dff_B_sNHTtnzO9_0),.clk(gclk));
	jdff dff_B_BzJNnD1D7_0(.din(w_dff_B_sNHTtnzO9_0),.dout(w_dff_B_BzJNnD1D7_0),.clk(gclk));
	jdff dff_B_BH4Of6eP9_0(.din(w_dff_B_BzJNnD1D7_0),.dout(w_dff_B_BH4Of6eP9_0),.clk(gclk));
	jdff dff_B_aVgAbiVL2_0(.din(w_dff_B_BH4Of6eP9_0),.dout(w_dff_B_aVgAbiVL2_0),.clk(gclk));
	jdff dff_B_A9IBnHUG1_0(.din(w_dff_B_aVgAbiVL2_0),.dout(w_dff_B_A9IBnHUG1_0),.clk(gclk));
	jdff dff_B_CZSJDSlp4_0(.din(w_dff_B_A9IBnHUG1_0),.dout(w_dff_B_CZSJDSlp4_0),.clk(gclk));
	jdff dff_B_CZ6KcnlD1_0(.din(w_dff_B_CZSJDSlp4_0),.dout(w_dff_B_CZ6KcnlD1_0),.clk(gclk));
	jdff dff_A_Xqu6oyos0_1(.dout(w_n1727_0[1]),.din(w_dff_A_Xqu6oyos0_1),.clk(gclk));
	jdff dff_A_FZsRS98w9_1(.dout(w_dff_A_Xqu6oyos0_1),.din(w_dff_A_FZsRS98w9_1),.clk(gclk));
	jdff dff_A_c2ocHHsM0_1(.dout(w_dff_A_FZsRS98w9_1),.din(w_dff_A_c2ocHHsM0_1),.clk(gclk));
	jdff dff_A_4hJbz2qi8_1(.dout(w_dff_A_c2ocHHsM0_1),.din(w_dff_A_4hJbz2qi8_1),.clk(gclk));
	jdff dff_A_UMsmR2nH5_1(.dout(w_dff_A_4hJbz2qi8_1),.din(w_dff_A_UMsmR2nH5_1),.clk(gclk));
	jdff dff_A_XA7goTYL7_1(.dout(w_dff_A_UMsmR2nH5_1),.din(w_dff_A_XA7goTYL7_1),.clk(gclk));
	jdff dff_A_zak9b8nx1_1(.dout(w_dff_A_XA7goTYL7_1),.din(w_dff_A_zak9b8nx1_1),.clk(gclk));
	jdff dff_A_6AwDm7zx1_1(.dout(w_dff_A_zak9b8nx1_1),.din(w_dff_A_6AwDm7zx1_1),.clk(gclk));
	jdff dff_A_ZVsb9R9N5_1(.dout(w_dff_A_6AwDm7zx1_1),.din(w_dff_A_ZVsb9R9N5_1),.clk(gclk));
	jdff dff_A_3MqrD0346_1(.dout(w_dff_A_ZVsb9R9N5_1),.din(w_dff_A_3MqrD0346_1),.clk(gclk));
	jdff dff_A_y6QKNNti8_1(.dout(w_dff_A_3MqrD0346_1),.din(w_dff_A_y6QKNNti8_1),.clk(gclk));
	jdff dff_A_9f82srkK4_1(.dout(w_dff_A_y6QKNNti8_1),.din(w_dff_A_9f82srkK4_1),.clk(gclk));
	jdff dff_A_5HE7nm6i7_1(.dout(w_dff_A_9f82srkK4_1),.din(w_dff_A_5HE7nm6i7_1),.clk(gclk));
	jdff dff_B_NiDVM0IL5_1(.din(n1691),.dout(w_dff_B_NiDVM0IL5_1),.clk(gclk));
	jdff dff_B_THVXFYeH5_1(.din(w_dff_B_NiDVM0IL5_1),.dout(w_dff_B_THVXFYeH5_1),.clk(gclk));
	jdff dff_B_7I4s2tqs1_1(.din(w_dff_B_THVXFYeH5_1),.dout(w_dff_B_7I4s2tqs1_1),.clk(gclk));
	jdff dff_B_RMbF241J6_1(.din(w_dff_B_7I4s2tqs1_1),.dout(w_dff_B_RMbF241J6_1),.clk(gclk));
	jdff dff_B_BmFgoTeU9_1(.din(w_dff_B_RMbF241J6_1),.dout(w_dff_B_BmFgoTeU9_1),.clk(gclk));
	jdff dff_B_DTPtxRqV5_1(.din(w_dff_B_BmFgoTeU9_1),.dout(w_dff_B_DTPtxRqV5_1),.clk(gclk));
	jdff dff_B_U4l6Lo1O8_1(.din(w_dff_B_DTPtxRqV5_1),.dout(w_dff_B_U4l6Lo1O8_1),.clk(gclk));
	jdff dff_B_opdsPIUC0_1(.din(w_dff_B_U4l6Lo1O8_1),.dout(w_dff_B_opdsPIUC0_1),.clk(gclk));
	jdff dff_B_R2IaWWdf9_1(.din(w_dff_B_opdsPIUC0_1),.dout(w_dff_B_R2IaWWdf9_1),.clk(gclk));
	jdff dff_B_CfiCXOBP8_1(.din(w_dff_B_R2IaWWdf9_1),.dout(w_dff_B_CfiCXOBP8_1),.clk(gclk));
	jdff dff_B_d17h1mHL1_1(.din(w_dff_B_CfiCXOBP8_1),.dout(w_dff_B_d17h1mHL1_1),.clk(gclk));
	jdff dff_B_mKcOYGMj2_1(.din(w_dff_B_d17h1mHL1_1),.dout(w_dff_B_mKcOYGMj2_1),.clk(gclk));
	jdff dff_B_BJyvovda8_1(.din(w_dff_B_mKcOYGMj2_1),.dout(w_dff_B_BJyvovda8_1),.clk(gclk));
	jdff dff_B_PHS5PLeG6_0(.din(n1692),.dout(w_dff_B_PHS5PLeG6_0),.clk(gclk));
	jdff dff_B_JIpurjGO8_0(.din(w_dff_B_PHS5PLeG6_0),.dout(w_dff_B_JIpurjGO8_0),.clk(gclk));
	jdff dff_B_sG6rwZFY1_0(.din(w_dff_B_JIpurjGO8_0),.dout(w_dff_B_sG6rwZFY1_0),.clk(gclk));
	jdff dff_B_oBhBHtF84_0(.din(w_dff_B_sG6rwZFY1_0),.dout(w_dff_B_oBhBHtF84_0),.clk(gclk));
	jdff dff_B_OdtYtcLg4_0(.din(w_dff_B_oBhBHtF84_0),.dout(w_dff_B_OdtYtcLg4_0),.clk(gclk));
	jdff dff_B_xsNTFTtr1_0(.din(w_dff_B_OdtYtcLg4_0),.dout(w_dff_B_xsNTFTtr1_0),.clk(gclk));
	jdff dff_B_WNGqTnbW3_0(.din(w_dff_B_xsNTFTtr1_0),.dout(w_dff_B_WNGqTnbW3_0),.clk(gclk));
	jdff dff_B_FKsoa0ir1_0(.din(w_dff_B_WNGqTnbW3_0),.dout(w_dff_B_FKsoa0ir1_0),.clk(gclk));
	jdff dff_B_RQHNHvPB1_0(.din(w_dff_B_FKsoa0ir1_0),.dout(w_dff_B_RQHNHvPB1_0),.clk(gclk));
	jdff dff_B_hxzfebwW3_0(.din(w_dff_B_RQHNHvPB1_0),.dout(w_dff_B_hxzfebwW3_0),.clk(gclk));
	jdff dff_B_OfOjkk3r2_0(.din(w_dff_B_hxzfebwW3_0),.dout(w_dff_B_OfOjkk3r2_0),.clk(gclk));
	jdff dff_A_vpGPPpDK3_1(.dout(w_n1689_0[1]),.din(w_dff_A_vpGPPpDK3_1),.clk(gclk));
	jdff dff_A_pSKzezHl3_1(.dout(w_dff_A_vpGPPpDK3_1),.din(w_dff_A_pSKzezHl3_1),.clk(gclk));
	jdff dff_A_Rusjejt27_1(.dout(w_dff_A_pSKzezHl3_1),.din(w_dff_A_Rusjejt27_1),.clk(gclk));
	jdff dff_A_M9euufRg3_1(.dout(w_dff_A_Rusjejt27_1),.din(w_dff_A_M9euufRg3_1),.clk(gclk));
	jdff dff_A_eRHyMjoD2_1(.dout(w_dff_A_M9euufRg3_1),.din(w_dff_A_eRHyMjoD2_1),.clk(gclk));
	jdff dff_A_PVXk5nwi7_1(.dout(w_dff_A_eRHyMjoD2_1),.din(w_dff_A_PVXk5nwi7_1),.clk(gclk));
	jdff dff_A_MfpC0Ifo4_1(.dout(w_dff_A_PVXk5nwi7_1),.din(w_dff_A_MfpC0Ifo4_1),.clk(gclk));
	jdff dff_A_hMwGH2CM1_1(.dout(w_dff_A_MfpC0Ifo4_1),.din(w_dff_A_hMwGH2CM1_1),.clk(gclk));
	jdff dff_A_Ybb0AtZm0_1(.dout(w_dff_A_hMwGH2CM1_1),.din(w_dff_A_Ybb0AtZm0_1),.clk(gclk));
	jdff dff_A_aXTdrMCm9_1(.dout(w_dff_A_Ybb0AtZm0_1),.din(w_dff_A_aXTdrMCm9_1),.clk(gclk));
	jdff dff_A_S3s5DZjn4_1(.dout(w_dff_A_aXTdrMCm9_1),.din(w_dff_A_S3s5DZjn4_1),.clk(gclk));
	jdff dff_A_tcFSoMZz5_1(.dout(w_dff_A_S3s5DZjn4_1),.din(w_dff_A_tcFSoMZz5_1),.clk(gclk));
	jdff dff_B_e3ghwwLt7_1(.din(n1643),.dout(w_dff_B_e3ghwwLt7_1),.clk(gclk));
	jdff dff_B_L9j5KGTg7_1(.din(w_dff_B_e3ghwwLt7_1),.dout(w_dff_B_L9j5KGTg7_1),.clk(gclk));
	jdff dff_B_2GY2a0XT6_1(.din(w_dff_B_L9j5KGTg7_1),.dout(w_dff_B_2GY2a0XT6_1),.clk(gclk));
	jdff dff_B_HVPxgTXN8_1(.din(w_dff_B_2GY2a0XT6_1),.dout(w_dff_B_HVPxgTXN8_1),.clk(gclk));
	jdff dff_B_mJSyy9Rn2_1(.din(w_dff_B_HVPxgTXN8_1),.dout(w_dff_B_mJSyy9Rn2_1),.clk(gclk));
	jdff dff_B_Aigm1sfF2_1(.din(w_dff_B_mJSyy9Rn2_1),.dout(w_dff_B_Aigm1sfF2_1),.clk(gclk));
	jdff dff_B_s606KOLh5_1(.din(w_dff_B_Aigm1sfF2_1),.dout(w_dff_B_s606KOLh5_1),.clk(gclk));
	jdff dff_B_OF9NdZiU4_1(.din(w_dff_B_s606KOLh5_1),.dout(w_dff_B_OF9NdZiU4_1),.clk(gclk));
	jdff dff_B_xoSSOig16_1(.din(w_dff_B_OF9NdZiU4_1),.dout(w_dff_B_xoSSOig16_1),.clk(gclk));
	jdff dff_B_m1bmlMH42_1(.din(w_dff_B_xoSSOig16_1),.dout(w_dff_B_m1bmlMH42_1),.clk(gclk));
	jdff dff_B_s8cq0cag8_1(.din(w_dff_B_m1bmlMH42_1),.dout(w_dff_B_s8cq0cag8_1),.clk(gclk));
	jdff dff_B_Dr5rfgtG5_1(.din(w_dff_B_s8cq0cag8_1),.dout(w_dff_B_Dr5rfgtG5_1),.clk(gclk));
	jdff dff_B_D1a7pTL46_0(.din(n1644),.dout(w_dff_B_D1a7pTL46_0),.clk(gclk));
	jdff dff_B_OyFgyPyf2_0(.din(w_dff_B_D1a7pTL46_0),.dout(w_dff_B_OyFgyPyf2_0),.clk(gclk));
	jdff dff_B_3Ws6aF4L7_0(.din(w_dff_B_OyFgyPyf2_0),.dout(w_dff_B_3Ws6aF4L7_0),.clk(gclk));
	jdff dff_B_ymzlpt8I1_0(.din(w_dff_B_3Ws6aF4L7_0),.dout(w_dff_B_ymzlpt8I1_0),.clk(gclk));
	jdff dff_B_OnHE1AtY9_0(.din(w_dff_B_ymzlpt8I1_0),.dout(w_dff_B_OnHE1AtY9_0),.clk(gclk));
	jdff dff_B_1oA95bXm2_0(.din(w_dff_B_OnHE1AtY9_0),.dout(w_dff_B_1oA95bXm2_0),.clk(gclk));
	jdff dff_B_dgtYZbqV3_0(.din(w_dff_B_1oA95bXm2_0),.dout(w_dff_B_dgtYZbqV3_0),.clk(gclk));
	jdff dff_B_Jo74UEam3_0(.din(w_dff_B_dgtYZbqV3_0),.dout(w_dff_B_Jo74UEam3_0),.clk(gclk));
	jdff dff_B_0nBRYLJG4_0(.din(w_dff_B_Jo74UEam3_0),.dout(w_dff_B_0nBRYLJG4_0),.clk(gclk));
	jdff dff_B_Dmfo7PaF5_0(.din(w_dff_B_0nBRYLJG4_0),.dout(w_dff_B_Dmfo7PaF5_0),.clk(gclk));
	jdff dff_A_4gYtos4m5_1(.dout(w_n1641_0[1]),.din(w_dff_A_4gYtos4m5_1),.clk(gclk));
	jdff dff_A_FV8rHZS99_1(.dout(w_dff_A_4gYtos4m5_1),.din(w_dff_A_FV8rHZS99_1),.clk(gclk));
	jdff dff_A_ydxLPViJ9_1(.dout(w_dff_A_FV8rHZS99_1),.din(w_dff_A_ydxLPViJ9_1),.clk(gclk));
	jdff dff_A_dhhiH5bd2_1(.dout(w_dff_A_ydxLPViJ9_1),.din(w_dff_A_dhhiH5bd2_1),.clk(gclk));
	jdff dff_A_Vcc0JimF0_1(.dout(w_dff_A_dhhiH5bd2_1),.din(w_dff_A_Vcc0JimF0_1),.clk(gclk));
	jdff dff_A_V8eDVjaH6_1(.dout(w_dff_A_Vcc0JimF0_1),.din(w_dff_A_V8eDVjaH6_1),.clk(gclk));
	jdff dff_A_GwGo1QBI6_1(.dout(w_dff_A_V8eDVjaH6_1),.din(w_dff_A_GwGo1QBI6_1),.clk(gclk));
	jdff dff_A_njHiTBld0_1(.dout(w_dff_A_GwGo1QBI6_1),.din(w_dff_A_njHiTBld0_1),.clk(gclk));
	jdff dff_A_S8IsL0Ib0_1(.dout(w_dff_A_njHiTBld0_1),.din(w_dff_A_S8IsL0Ib0_1),.clk(gclk));
	jdff dff_A_DhK7EMWn8_1(.dout(w_dff_A_S8IsL0Ib0_1),.din(w_dff_A_DhK7EMWn8_1),.clk(gclk));
	jdff dff_A_0iecNvAh2_1(.dout(w_dff_A_DhK7EMWn8_1),.din(w_dff_A_0iecNvAh2_1),.clk(gclk));
	jdff dff_B_LJJlWnk41_1(.din(n1588),.dout(w_dff_B_LJJlWnk41_1),.clk(gclk));
	jdff dff_B_3piuALWv7_1(.din(w_dff_B_LJJlWnk41_1),.dout(w_dff_B_3piuALWv7_1),.clk(gclk));
	jdff dff_B_oTDNCRoU0_1(.din(w_dff_B_3piuALWv7_1),.dout(w_dff_B_oTDNCRoU0_1),.clk(gclk));
	jdff dff_B_9Cz1FamL9_1(.din(w_dff_B_oTDNCRoU0_1),.dout(w_dff_B_9Cz1FamL9_1),.clk(gclk));
	jdff dff_B_Ag025cPL1_1(.din(w_dff_B_9Cz1FamL9_1),.dout(w_dff_B_Ag025cPL1_1),.clk(gclk));
	jdff dff_B_lk0hO8Yq2_1(.din(w_dff_B_Ag025cPL1_1),.dout(w_dff_B_lk0hO8Yq2_1),.clk(gclk));
	jdff dff_B_Z6oXm97H1_1(.din(w_dff_B_lk0hO8Yq2_1),.dout(w_dff_B_Z6oXm97H1_1),.clk(gclk));
	jdff dff_B_WQEF9ekj2_1(.din(w_dff_B_Z6oXm97H1_1),.dout(w_dff_B_WQEF9ekj2_1),.clk(gclk));
	jdff dff_B_hmfNt6b79_1(.din(w_dff_B_WQEF9ekj2_1),.dout(w_dff_B_hmfNt6b79_1),.clk(gclk));
	jdff dff_B_fPT3ph2e2_1(.din(w_dff_B_hmfNt6b79_1),.dout(w_dff_B_fPT3ph2e2_1),.clk(gclk));
	jdff dff_B_lxy4xvBU3_0(.din(n1589),.dout(w_dff_B_lxy4xvBU3_0),.clk(gclk));
	jdff dff_B_zpgqweIC2_0(.din(w_dff_B_lxy4xvBU3_0),.dout(w_dff_B_zpgqweIC2_0),.clk(gclk));
	jdff dff_B_PrMF6BJ27_0(.din(w_dff_B_zpgqweIC2_0),.dout(w_dff_B_PrMF6BJ27_0),.clk(gclk));
	jdff dff_B_dNHn36ia0_0(.din(w_dff_B_PrMF6BJ27_0),.dout(w_dff_B_dNHn36ia0_0),.clk(gclk));
	jdff dff_B_dMpuQB7g0_0(.din(w_dff_B_dNHn36ia0_0),.dout(w_dff_B_dMpuQB7g0_0),.clk(gclk));
	jdff dff_B_vyKnG3id5_0(.din(w_dff_B_dMpuQB7g0_0),.dout(w_dff_B_vyKnG3id5_0),.clk(gclk));
	jdff dff_B_FU2qZ6LP7_0(.din(w_dff_B_vyKnG3id5_0),.dout(w_dff_B_FU2qZ6LP7_0),.clk(gclk));
	jdff dff_B_7MkU68A62_0(.din(w_dff_B_FU2qZ6LP7_0),.dout(w_dff_B_7MkU68A62_0),.clk(gclk));
	jdff dff_A_MRcvc1uA4_1(.dout(w_n1586_0[1]),.din(w_dff_A_MRcvc1uA4_1),.clk(gclk));
	jdff dff_A_yu7UUQFT7_1(.dout(w_dff_A_MRcvc1uA4_1),.din(w_dff_A_yu7UUQFT7_1),.clk(gclk));
	jdff dff_A_OthvHi1X1_1(.dout(w_dff_A_yu7UUQFT7_1),.din(w_dff_A_OthvHi1X1_1),.clk(gclk));
	jdff dff_A_bF84zSeK2_1(.dout(w_dff_A_OthvHi1X1_1),.din(w_dff_A_bF84zSeK2_1),.clk(gclk));
	jdff dff_A_ENBa59xu0_1(.dout(w_dff_A_bF84zSeK2_1),.din(w_dff_A_ENBa59xu0_1),.clk(gclk));
	jdff dff_A_1h5GEteT0_1(.dout(w_dff_A_ENBa59xu0_1),.din(w_dff_A_1h5GEteT0_1),.clk(gclk));
	jdff dff_A_Usz5I9JG5_1(.dout(w_dff_A_1h5GEteT0_1),.din(w_dff_A_Usz5I9JG5_1),.clk(gclk));
	jdff dff_A_2sHKpfZJ6_1(.dout(w_dff_A_Usz5I9JG5_1),.din(w_dff_A_2sHKpfZJ6_1),.clk(gclk));
	jdff dff_A_xuraak5w1_1(.dout(w_dff_A_2sHKpfZJ6_1),.din(w_dff_A_xuraak5w1_1),.clk(gclk));
	jdff dff_B_ufxgNgqS8_1(.din(n1526),.dout(w_dff_B_ufxgNgqS8_1),.clk(gclk));
	jdff dff_B_ztb9utD51_1(.din(w_dff_B_ufxgNgqS8_1),.dout(w_dff_B_ztb9utD51_1),.clk(gclk));
	jdff dff_B_kKiGYkkF8_1(.din(w_dff_B_ztb9utD51_1),.dout(w_dff_B_kKiGYkkF8_1),.clk(gclk));
	jdff dff_B_FLJ4YpMp7_1(.din(w_dff_B_kKiGYkkF8_1),.dout(w_dff_B_FLJ4YpMp7_1),.clk(gclk));
	jdff dff_B_sDoBt1Vb4_1(.din(w_dff_B_FLJ4YpMp7_1),.dout(w_dff_B_sDoBt1Vb4_1),.clk(gclk));
	jdff dff_B_pgsVoisl2_1(.din(w_dff_B_sDoBt1Vb4_1),.dout(w_dff_B_pgsVoisl2_1),.clk(gclk));
	jdff dff_B_wJdjq6UD9_1(.din(w_dff_B_pgsVoisl2_1),.dout(w_dff_B_wJdjq6UD9_1),.clk(gclk));
	jdff dff_B_la4C7ecR3_1(.din(w_dff_B_wJdjq6UD9_1),.dout(w_dff_B_la4C7ecR3_1),.clk(gclk));
	jdff dff_B_dWAYz2Rc7_0(.din(n1527),.dout(w_dff_B_dWAYz2Rc7_0),.clk(gclk));
	jdff dff_B_1epMpAng0_0(.din(w_dff_B_dWAYz2Rc7_0),.dout(w_dff_B_1epMpAng0_0),.clk(gclk));
	jdff dff_B_Bz65Kcuo5_0(.din(w_dff_B_1epMpAng0_0),.dout(w_dff_B_Bz65Kcuo5_0),.clk(gclk));
	jdff dff_B_98FrXcK27_0(.din(w_dff_B_Bz65Kcuo5_0),.dout(w_dff_B_98FrXcK27_0),.clk(gclk));
	jdff dff_B_5zVSnA2z6_0(.din(w_dff_B_98FrXcK27_0),.dout(w_dff_B_5zVSnA2z6_0),.clk(gclk));
	jdff dff_B_NW2B2g9Z9_0(.din(w_dff_B_5zVSnA2z6_0),.dout(w_dff_B_NW2B2g9Z9_0),.clk(gclk));
	jdff dff_A_XFDpb1RG5_1(.dout(w_n1524_0[1]),.din(w_dff_A_XFDpb1RG5_1),.clk(gclk));
	jdff dff_A_3JmpqIru4_1(.dout(w_dff_A_XFDpb1RG5_1),.din(w_dff_A_3JmpqIru4_1),.clk(gclk));
	jdff dff_A_xbN7cE4m9_1(.dout(w_dff_A_3JmpqIru4_1),.din(w_dff_A_xbN7cE4m9_1),.clk(gclk));
	jdff dff_A_AGCUTb3e5_1(.dout(w_dff_A_xbN7cE4m9_1),.din(w_dff_A_AGCUTb3e5_1),.clk(gclk));
	jdff dff_A_o1mjaOtS0_1(.dout(w_dff_A_AGCUTb3e5_1),.din(w_dff_A_o1mjaOtS0_1),.clk(gclk));
	jdff dff_A_CzaZjN317_1(.dout(w_dff_A_o1mjaOtS0_1),.din(w_dff_A_CzaZjN317_1),.clk(gclk));
	jdff dff_A_G45fXfk25_1(.dout(w_dff_A_CzaZjN317_1),.din(w_dff_A_G45fXfk25_1),.clk(gclk));
	jdff dff_B_99jEtv879_1(.din(n1457),.dout(w_dff_B_99jEtv879_1),.clk(gclk));
	jdff dff_B_RwJTWK5E1_1(.din(w_dff_B_99jEtv879_1),.dout(w_dff_B_RwJTWK5E1_1),.clk(gclk));
	jdff dff_B_D62o8hER1_1(.din(w_dff_B_RwJTWK5E1_1),.dout(w_dff_B_D62o8hER1_1),.clk(gclk));
	jdff dff_B_JohTtuWZ5_1(.din(w_dff_B_D62o8hER1_1),.dout(w_dff_B_JohTtuWZ5_1),.clk(gclk));
	jdff dff_B_zctOC7Yx2_1(.din(w_dff_B_JohTtuWZ5_1),.dout(w_dff_B_zctOC7Yx2_1),.clk(gclk));
	jdff dff_B_u2wEuWIl8_1(.din(w_dff_B_zctOC7Yx2_1),.dout(w_dff_B_u2wEuWIl8_1),.clk(gclk));
	jdff dff_B_6M8TUMrb7_1(.din(w_dff_B_u2wEuWIl8_1),.dout(w_dff_B_6M8TUMrb7_1),.clk(gclk));
	jdff dff_B_uzcjNXjC1_0(.din(n1458),.dout(w_dff_B_uzcjNXjC1_0),.clk(gclk));
	jdff dff_B_zq4uOzPE2_0(.din(w_dff_B_uzcjNXjC1_0),.dout(w_dff_B_zq4uOzPE2_0),.clk(gclk));
	jdff dff_B_7hI0vCHj9_0(.din(w_dff_B_zq4uOzPE2_0),.dout(w_dff_B_7hI0vCHj9_0),.clk(gclk));
	jdff dff_B_HrYEjpWa5_0(.din(w_dff_B_7hI0vCHj9_0),.dout(w_dff_B_HrYEjpWa5_0),.clk(gclk));
	jdff dff_B_HRfc0iEy8_0(.din(w_dff_B_HrYEjpWa5_0),.dout(w_dff_B_HRfc0iEy8_0),.clk(gclk));
	jdff dff_A_Lrjqb8Q71_1(.dout(w_n1455_0[1]),.din(w_dff_A_Lrjqb8Q71_1),.clk(gclk));
	jdff dff_A_ggzCto9m0_1(.dout(w_dff_A_Lrjqb8Q71_1),.din(w_dff_A_ggzCto9m0_1),.clk(gclk));
	jdff dff_A_VVPVeflc3_1(.dout(w_dff_A_ggzCto9m0_1),.din(w_dff_A_VVPVeflc3_1),.clk(gclk));
	jdff dff_A_6UoLyPy62_1(.dout(w_dff_A_VVPVeflc3_1),.din(w_dff_A_6UoLyPy62_1),.clk(gclk));
	jdff dff_A_ajr6RC2b0_1(.dout(w_dff_A_6UoLyPy62_1),.din(w_dff_A_ajr6RC2b0_1),.clk(gclk));
	jdff dff_A_vTJCgUqr5_1(.dout(w_dff_A_ajr6RC2b0_1),.din(w_dff_A_vTJCgUqr5_1),.clk(gclk));
	jdff dff_B_DtWOtbt48_1(.din(n1381),.dout(w_dff_B_DtWOtbt48_1),.clk(gclk));
	jdff dff_B_x6YGrWCP2_1(.din(w_dff_B_DtWOtbt48_1),.dout(w_dff_B_x6YGrWCP2_1),.clk(gclk));
	jdff dff_B_cgKo1uKb5_1(.din(w_dff_B_x6YGrWCP2_1),.dout(w_dff_B_cgKo1uKb5_1),.clk(gclk));
	jdff dff_B_sNmOolNm6_1(.din(w_dff_B_cgKo1uKb5_1),.dout(w_dff_B_sNmOolNm6_1),.clk(gclk));
	jdff dff_B_Ly4X3evK3_1(.din(w_dff_B_sNmOolNm6_1),.dout(w_dff_B_Ly4X3evK3_1),.clk(gclk));
	jdff dff_B_5Qqva24S8_1(.din(w_dff_B_Ly4X3evK3_1),.dout(w_dff_B_5Qqva24S8_1),.clk(gclk));
	jdff dff_B_0BX5uYEF9_0(.din(n1382),.dout(w_dff_B_0BX5uYEF9_0),.clk(gclk));
	jdff dff_B_b6oP3IBR6_0(.din(w_dff_B_0BX5uYEF9_0),.dout(w_dff_B_b6oP3IBR6_0),.clk(gclk));
	jdff dff_B_2pCn1TmJ8_0(.din(w_dff_B_b6oP3IBR6_0),.dout(w_dff_B_2pCn1TmJ8_0),.clk(gclk));
	jdff dff_B_ZlZ6Nbus7_0(.din(w_dff_B_2pCn1TmJ8_0),.dout(w_dff_B_ZlZ6Nbus7_0),.clk(gclk));
	jdff dff_A_4ONEt3wy6_1(.dout(w_n1379_0[1]),.din(w_dff_A_4ONEt3wy6_1),.clk(gclk));
	jdff dff_A_2j2h0TO31_1(.dout(w_dff_A_4ONEt3wy6_1),.din(w_dff_A_2j2h0TO31_1),.clk(gclk));
	jdff dff_A_LPtiH6V44_1(.dout(w_dff_A_2j2h0TO31_1),.din(w_dff_A_LPtiH6V44_1),.clk(gclk));
	jdff dff_A_ytACUHtR0_1(.dout(w_dff_A_LPtiH6V44_1),.din(w_dff_A_ytACUHtR0_1),.clk(gclk));
	jdff dff_A_eCoR4Xyq0_1(.dout(w_dff_A_ytACUHtR0_1),.din(w_dff_A_eCoR4Xyq0_1),.clk(gclk));
	jdff dff_B_ciEhE5oa1_1(.din(n1299),.dout(w_dff_B_ciEhE5oa1_1),.clk(gclk));
	jdff dff_B_CwNbjt9l7_1(.din(w_dff_B_ciEhE5oa1_1),.dout(w_dff_B_CwNbjt9l7_1),.clk(gclk));
	jdff dff_B_kUkGjYFU6_1(.din(w_dff_B_CwNbjt9l7_1),.dout(w_dff_B_kUkGjYFU6_1),.clk(gclk));
	jdff dff_A_LFIfuljK0_0(.dout(w_n1295_0[0]),.din(w_dff_A_LFIfuljK0_0),.clk(gclk));
	jdff dff_A_HSElSoIF5_0(.dout(w_dff_A_LFIfuljK0_0),.din(w_dff_A_HSElSoIF5_0),.clk(gclk));
	jdff dff_B_4lbaaL8i8_1(.din(n1211),.dout(w_dff_B_4lbaaL8i8_1),.clk(gclk));
	jdff dff_A_PYphhLrQ4_0(.dout(w_n1207_0[0]),.din(w_dff_A_PYphhLrQ4_0),.clk(gclk));
	jdff dff_B_RwNnqVnb6_1(.din(n1113),.dout(w_dff_B_RwNnqVnb6_1),.clk(gclk));
	jdff dff_A_0ILHXRq21_1(.dout(w_n1013_0[1]),.din(w_dff_A_0ILHXRq21_1),.clk(gclk));
	jdff dff_B_T4lBY7sl2_2(.din(n1011),.dout(w_dff_B_T4lBY7sl2_2),.clk(gclk));
	jdff dff_B_4xi7J29C7_1(.din(n908),.dout(w_dff_B_4xi7J29C7_1),.clk(gclk));
	jdff dff_A_7wZHuWQL2_0(.dout(w_n805_0[0]),.din(w_dff_A_7wZHuWQL2_0),.clk(gclk));
	jdff dff_A_6cJ0fW5k2_0(.dout(w_dff_A_7wZHuWQL2_0),.din(w_dff_A_6cJ0fW5k2_0),.clk(gclk));
	jdff dff_A_uhSwwA6H0_0(.dout(w_dff_A_6cJ0fW5k2_0),.din(w_dff_A_uhSwwA6H0_0),.clk(gclk));
	jdff dff_A_f0TEMAuq8_0(.dout(w_dff_A_uhSwwA6H0_0),.din(w_dff_A_f0TEMAuq8_0),.clk(gclk));
	jdff dff_A_h7EAVs6D4_0(.dout(w_dff_A_f0TEMAuq8_0),.din(w_dff_A_h7EAVs6D4_0),.clk(gclk));
	jdff dff_A_rq093ssw9_0(.dout(w_dff_A_h7EAVs6D4_0),.din(w_dff_A_rq093ssw9_0),.clk(gclk));
	jdff dff_A_tdctkbOV7_0(.dout(w_dff_A_rq093ssw9_0),.din(w_dff_A_tdctkbOV7_0),.clk(gclk));
	jdff dff_A_IRIJoYKg8_0(.dout(w_dff_A_tdctkbOV7_0),.din(w_dff_A_IRIJoYKg8_0),.clk(gclk));
	jdff dff_A_x3REjARl0_0(.dout(w_dff_A_IRIJoYKg8_0),.din(w_dff_A_x3REjARl0_0),.clk(gclk));
	jdff dff_A_BnG97WkD2_0(.dout(w_dff_A_x3REjARl0_0),.din(w_dff_A_BnG97WkD2_0),.clk(gclk));
	jdff dff_A_519OxtWA7_0(.dout(w_dff_A_BnG97WkD2_0),.din(w_dff_A_519OxtWA7_0),.clk(gclk));
	jdff dff_A_GUR3HTEq2_0(.dout(w_dff_A_519OxtWA7_0),.din(w_dff_A_GUR3HTEq2_0),.clk(gclk));
	jdff dff_A_Ol7f7Yt26_0(.dout(w_dff_A_GUR3HTEq2_0),.din(w_dff_A_Ol7f7Yt26_0),.clk(gclk));
	jdff dff_A_qEkqeOYb4_0(.dout(w_dff_A_Ol7f7Yt26_0),.din(w_dff_A_qEkqeOYb4_0),.clk(gclk));
	jdff dff_A_p7tFtE577_0(.dout(w_dff_A_qEkqeOYb4_0),.din(w_dff_A_p7tFtE577_0),.clk(gclk));
	jdff dff_A_ZBV2MSCJ5_0(.dout(w_dff_A_p7tFtE577_0),.din(w_dff_A_ZBV2MSCJ5_0),.clk(gclk));
	jdff dff_A_Ye1uCfar5_0(.dout(w_dff_A_ZBV2MSCJ5_0),.din(w_dff_A_Ye1uCfar5_0),.clk(gclk));
	jdff dff_A_U3V8u78H4_0(.dout(w_dff_A_Ye1uCfar5_0),.din(w_dff_A_U3V8u78H4_0),.clk(gclk));
	jdff dff_A_pvdl4QGc7_0(.dout(w_dff_A_U3V8u78H4_0),.din(w_dff_A_pvdl4QGc7_0),.clk(gclk));
	jdff dff_A_hJ8zBZk38_0(.dout(w_dff_A_pvdl4QGc7_0),.din(w_dff_A_hJ8zBZk38_0),.clk(gclk));
	jdff dff_A_UAq6hRJH3_0(.dout(w_dff_A_hJ8zBZk38_0),.din(w_dff_A_UAq6hRJH3_0),.clk(gclk));
	jdff dff_A_NGo2YtPo8_0(.dout(w_dff_A_UAq6hRJH3_0),.din(w_dff_A_NGo2YtPo8_0),.clk(gclk));
	jdff dff_A_2sVv8gC40_0(.dout(w_dff_A_NGo2YtPo8_0),.din(w_dff_A_2sVv8gC40_0),.clk(gclk));
	jdff dff_A_G5Ho0abw3_0(.dout(w_dff_A_2sVv8gC40_0),.din(w_dff_A_G5Ho0abw3_0),.clk(gclk));
	jdff dff_A_zQaSjH4w4_0(.dout(w_dff_A_G5Ho0abw3_0),.din(w_dff_A_zQaSjH4w4_0),.clk(gclk));
	jdff dff_A_6vw6P3qt7_0(.dout(w_dff_A_zQaSjH4w4_0),.din(w_dff_A_6vw6P3qt7_0),.clk(gclk));
	jdff dff_A_fSUzXhIk9_0(.dout(w_dff_A_6vw6P3qt7_0),.din(w_dff_A_fSUzXhIk9_0),.clk(gclk));
	jdff dff_A_5ulZx8a16_0(.dout(w_dff_A_fSUzXhIk9_0),.din(w_dff_A_5ulZx8a16_0),.clk(gclk));
	jdff dff_A_VItp2do45_0(.dout(w_dff_A_5ulZx8a16_0),.din(w_dff_A_VItp2do45_0),.clk(gclk));
	jdff dff_A_xLxnb5Pd4_0(.dout(w_dff_A_VItp2do45_0),.din(w_dff_A_xLxnb5Pd4_0),.clk(gclk));
	jdff dff_A_mADrcsg95_0(.dout(w_dff_A_xLxnb5Pd4_0),.din(w_dff_A_mADrcsg95_0),.clk(gclk));
	jdff dff_A_gL54cPH75_0(.dout(w_dff_A_mADrcsg95_0),.din(w_dff_A_gL54cPH75_0),.clk(gclk));
	jdff dff_A_IORHVl6G9_0(.dout(w_dff_A_gL54cPH75_0),.din(w_dff_A_IORHVl6G9_0),.clk(gclk));
	jdff dff_A_TyhxclkV9_0(.dout(w_dff_A_IORHVl6G9_0),.din(w_dff_A_TyhxclkV9_0),.clk(gclk));
	jdff dff_A_3vCRfo9D2_0(.dout(w_dff_A_TyhxclkV9_0),.din(w_dff_A_3vCRfo9D2_0),.clk(gclk));
	jdff dff_A_DWvgFadZ6_0(.dout(w_dff_A_3vCRfo9D2_0),.din(w_dff_A_DWvgFadZ6_0),.clk(gclk));
	jdff dff_A_yC5md7O78_0(.dout(w_dff_A_DWvgFadZ6_0),.din(w_dff_A_yC5md7O78_0),.clk(gclk));
	jdff dff_A_Pamahlte9_0(.dout(w_dff_A_yC5md7O78_0),.din(w_dff_A_Pamahlte9_0),.clk(gclk));
	jdff dff_A_SlVhe1Ga5_0(.dout(w_dff_A_Pamahlte9_0),.din(w_dff_A_SlVhe1Ga5_0),.clk(gclk));
	jdff dff_A_ozVsdxvV6_0(.dout(w_dff_A_SlVhe1Ga5_0),.din(w_dff_A_ozVsdxvV6_0),.clk(gclk));
	jdff dff_A_2j9truBF6_0(.dout(w_dff_A_ozVsdxvV6_0),.din(w_dff_A_2j9truBF6_0),.clk(gclk));
	jdff dff_A_nCOFFhXa2_0(.dout(w_dff_A_2j9truBF6_0),.din(w_dff_A_nCOFFhXa2_0),.clk(gclk));
	jdff dff_A_fOMSH2Sk7_0(.dout(w_dff_A_nCOFFhXa2_0),.din(w_dff_A_fOMSH2Sk7_0),.clk(gclk));
	jdff dff_A_ra8b89sL4_1(.dout(w_n904_0[1]),.din(w_dff_A_ra8b89sL4_1),.clk(gclk));
	jdff dff_B_fUgsaO6R2_1(.din(n808),.dout(w_dff_B_fUgsaO6R2_1),.clk(gclk));
	jdff dff_A_9MiIiI5w5_0(.dout(w_n706_0[0]),.din(w_dff_A_9MiIiI5w5_0),.clk(gclk));
	jdff dff_A_waEKkhjf6_0(.dout(w_dff_A_9MiIiI5w5_0),.din(w_dff_A_waEKkhjf6_0),.clk(gclk));
	jdff dff_A_69ytUQ3A2_0(.dout(w_dff_A_waEKkhjf6_0),.din(w_dff_A_69ytUQ3A2_0),.clk(gclk));
	jdff dff_A_cricFCtc1_0(.dout(w_dff_A_69ytUQ3A2_0),.din(w_dff_A_cricFCtc1_0),.clk(gclk));
	jdff dff_A_FqntZ5Tl4_0(.dout(w_dff_A_cricFCtc1_0),.din(w_dff_A_FqntZ5Tl4_0),.clk(gclk));
	jdff dff_A_BDf71oEe9_0(.dout(w_dff_A_FqntZ5Tl4_0),.din(w_dff_A_BDf71oEe9_0),.clk(gclk));
	jdff dff_A_VV4S4COs5_0(.dout(w_dff_A_BDf71oEe9_0),.din(w_dff_A_VV4S4COs5_0),.clk(gclk));
	jdff dff_A_iEuW9GLf4_0(.dout(w_dff_A_VV4S4COs5_0),.din(w_dff_A_iEuW9GLf4_0),.clk(gclk));
	jdff dff_A_wGF92iH39_0(.dout(w_dff_A_iEuW9GLf4_0),.din(w_dff_A_wGF92iH39_0),.clk(gclk));
	jdff dff_A_0cM9jCbq7_0(.dout(w_dff_A_wGF92iH39_0),.din(w_dff_A_0cM9jCbq7_0),.clk(gclk));
	jdff dff_A_1RFis5Qd1_0(.dout(w_dff_A_0cM9jCbq7_0),.din(w_dff_A_1RFis5Qd1_0),.clk(gclk));
	jdff dff_A_M7FYKQnL0_0(.dout(w_dff_A_1RFis5Qd1_0),.din(w_dff_A_M7FYKQnL0_0),.clk(gclk));
	jdff dff_A_ZuQNXriM2_0(.dout(w_dff_A_M7FYKQnL0_0),.din(w_dff_A_ZuQNXriM2_0),.clk(gclk));
	jdff dff_A_A8vXEfk04_0(.dout(w_dff_A_ZuQNXriM2_0),.din(w_dff_A_A8vXEfk04_0),.clk(gclk));
	jdff dff_A_fHoQzASn9_0(.dout(w_dff_A_A8vXEfk04_0),.din(w_dff_A_fHoQzASn9_0),.clk(gclk));
	jdff dff_A_q3L2bRJV4_0(.dout(w_dff_A_fHoQzASn9_0),.din(w_dff_A_q3L2bRJV4_0),.clk(gclk));
	jdff dff_A_BHblP0pF8_0(.dout(w_dff_A_q3L2bRJV4_0),.din(w_dff_A_BHblP0pF8_0),.clk(gclk));
	jdff dff_A_80Ax4HiU1_0(.dout(w_dff_A_BHblP0pF8_0),.din(w_dff_A_80Ax4HiU1_0),.clk(gclk));
	jdff dff_A_a7bQXuza9_0(.dout(w_dff_A_80Ax4HiU1_0),.din(w_dff_A_a7bQXuza9_0),.clk(gclk));
	jdff dff_A_d3Gl7lLy4_0(.dout(w_dff_A_a7bQXuza9_0),.din(w_dff_A_d3Gl7lLy4_0),.clk(gclk));
	jdff dff_A_meFxOqsl9_0(.dout(w_dff_A_d3Gl7lLy4_0),.din(w_dff_A_meFxOqsl9_0),.clk(gclk));
	jdff dff_A_S2lwdrPZ8_0(.dout(w_dff_A_meFxOqsl9_0),.din(w_dff_A_S2lwdrPZ8_0),.clk(gclk));
	jdff dff_A_y5gs4Hco1_0(.dout(w_dff_A_S2lwdrPZ8_0),.din(w_dff_A_y5gs4Hco1_0),.clk(gclk));
	jdff dff_A_2QmPDKaM1_0(.dout(w_dff_A_y5gs4Hco1_0),.din(w_dff_A_2QmPDKaM1_0),.clk(gclk));
	jdff dff_A_82jbZI446_0(.dout(w_dff_A_2QmPDKaM1_0),.din(w_dff_A_82jbZI446_0),.clk(gclk));
	jdff dff_A_rK3tfZIg7_0(.dout(w_dff_A_82jbZI446_0),.din(w_dff_A_rK3tfZIg7_0),.clk(gclk));
	jdff dff_A_UAWSx7hy1_0(.dout(w_dff_A_rK3tfZIg7_0),.din(w_dff_A_UAWSx7hy1_0),.clk(gclk));
	jdff dff_A_Ko96IlfN0_0(.dout(w_dff_A_UAWSx7hy1_0),.din(w_dff_A_Ko96IlfN0_0),.clk(gclk));
	jdff dff_A_j9RYdZ2H2_0(.dout(w_dff_A_Ko96IlfN0_0),.din(w_dff_A_j9RYdZ2H2_0),.clk(gclk));
	jdff dff_A_Q0cTpnbQ8_0(.dout(w_dff_A_j9RYdZ2H2_0),.din(w_dff_A_Q0cTpnbQ8_0),.clk(gclk));
	jdff dff_A_wNsxdpsx3_0(.dout(w_dff_A_Q0cTpnbQ8_0),.din(w_dff_A_wNsxdpsx3_0),.clk(gclk));
	jdff dff_A_avqQY4bb2_0(.dout(w_dff_A_wNsxdpsx3_0),.din(w_dff_A_avqQY4bb2_0),.clk(gclk));
	jdff dff_A_infK8D7j8_0(.dout(w_dff_A_avqQY4bb2_0),.din(w_dff_A_infK8D7j8_0),.clk(gclk));
	jdff dff_A_pbCOyc8h0_0(.dout(w_dff_A_infK8D7j8_0),.din(w_dff_A_pbCOyc8h0_0),.clk(gclk));
	jdff dff_A_DtMsdpwU6_0(.dout(w_dff_A_pbCOyc8h0_0),.din(w_dff_A_DtMsdpwU6_0),.clk(gclk));
	jdff dff_A_A5FpTrrD7_0(.dout(w_dff_A_DtMsdpwU6_0),.din(w_dff_A_A5FpTrrD7_0),.clk(gclk));
	jdff dff_A_CVFsShbn7_0(.dout(w_dff_A_A5FpTrrD7_0),.din(w_dff_A_CVFsShbn7_0),.clk(gclk));
	jdff dff_A_75sGKR2N7_0(.dout(w_dff_A_CVFsShbn7_0),.din(w_dff_A_75sGKR2N7_0),.clk(gclk));
	jdff dff_A_juJ0YWCi8_0(.dout(w_dff_A_75sGKR2N7_0),.din(w_dff_A_juJ0YWCi8_0),.clk(gclk));
	jdff dff_A_Evzuf2IR8_0(.dout(w_dff_A_juJ0YWCi8_0),.din(w_dff_A_Evzuf2IR8_0),.clk(gclk));
	jdff dff_A_8ocpneNJ7_1(.dout(w_n802_0[1]),.din(w_dff_A_8ocpneNJ7_1),.clk(gclk));
	jdff dff_B_f2s8ll5S7_1(.din(n713),.dout(w_dff_B_f2s8ll5S7_1),.clk(gclk));
	jdff dff_B_7zUKubWB6_1(.din(w_dff_B_f2s8ll5S7_1),.dout(w_dff_B_7zUKubWB6_1),.clk(gclk));
	jdff dff_B_g3NAIaP19_1(.din(w_dff_B_7zUKubWB6_1),.dout(w_dff_B_g3NAIaP19_1),.clk(gclk));
	jdff dff_B_zKyZ22v46_1(.din(w_dff_B_g3NAIaP19_1),.dout(w_dff_B_zKyZ22v46_1),.clk(gclk));
	jdff dff_B_mpMOliPw9_1(.din(w_dff_B_zKyZ22v46_1),.dout(w_dff_B_mpMOliPw9_1),.clk(gclk));
	jdff dff_B_bcE9CSpy9_1(.din(w_dff_B_mpMOliPw9_1),.dout(w_dff_B_bcE9CSpy9_1),.clk(gclk));
	jdff dff_B_dlzDynoQ1_1(.din(w_dff_B_bcE9CSpy9_1),.dout(w_dff_B_dlzDynoQ1_1),.clk(gclk));
	jdff dff_B_j0tIeTl78_1(.din(w_dff_B_dlzDynoQ1_1),.dout(w_dff_B_j0tIeTl78_1),.clk(gclk));
	jdff dff_B_pLlDu1QI6_1(.din(w_dff_B_j0tIeTl78_1),.dout(w_dff_B_pLlDu1QI6_1),.clk(gclk));
	jdff dff_B_IPAGpyNa0_1(.din(w_dff_B_pLlDu1QI6_1),.dout(w_dff_B_IPAGpyNa0_1),.clk(gclk));
	jdff dff_B_u30lyc8x6_1(.din(w_dff_B_IPAGpyNa0_1),.dout(w_dff_B_u30lyc8x6_1),.clk(gclk));
	jdff dff_B_g9Bj4mR33_1(.din(w_dff_B_u30lyc8x6_1),.dout(w_dff_B_g9Bj4mR33_1),.clk(gclk));
	jdff dff_B_nKzF8pWz9_1(.din(w_dff_B_g9Bj4mR33_1),.dout(w_dff_B_nKzF8pWz9_1),.clk(gclk));
	jdff dff_B_TEq6th2s5_1(.din(w_dff_B_nKzF8pWz9_1),.dout(w_dff_B_TEq6th2s5_1),.clk(gclk));
	jdff dff_B_nKuV32Vx8_1(.din(w_dff_B_TEq6th2s5_1),.dout(w_dff_B_nKuV32Vx8_1),.clk(gclk));
	jdff dff_B_h6kLfVcb0_1(.din(w_dff_B_nKuV32Vx8_1),.dout(w_dff_B_h6kLfVcb0_1),.clk(gclk));
	jdff dff_B_RiyIr1VH1_1(.din(w_dff_B_h6kLfVcb0_1),.dout(w_dff_B_RiyIr1VH1_1),.clk(gclk));
	jdff dff_B_Gympt39G8_1(.din(w_dff_B_RiyIr1VH1_1),.dout(w_dff_B_Gympt39G8_1),.clk(gclk));
	jdff dff_B_auS0WcJ65_1(.din(w_dff_B_Gympt39G8_1),.dout(w_dff_B_auS0WcJ65_1),.clk(gclk));
	jdff dff_B_uHsCIQpA1_1(.din(w_dff_B_auS0WcJ65_1),.dout(w_dff_B_uHsCIQpA1_1),.clk(gclk));
	jdff dff_B_pOAFj4aZ1_1(.din(w_dff_B_uHsCIQpA1_1),.dout(w_dff_B_pOAFj4aZ1_1),.clk(gclk));
	jdff dff_B_aYxePEI51_1(.din(w_dff_B_pOAFj4aZ1_1),.dout(w_dff_B_aYxePEI51_1),.clk(gclk));
	jdff dff_B_KW18rf0u3_1(.din(w_dff_B_aYxePEI51_1),.dout(w_dff_B_KW18rf0u3_1),.clk(gclk));
	jdff dff_B_hygbpTQG2_1(.din(w_dff_B_KW18rf0u3_1),.dout(w_dff_B_hygbpTQG2_1),.clk(gclk));
	jdff dff_B_l2DXJUKw7_1(.din(w_dff_B_hygbpTQG2_1),.dout(w_dff_B_l2DXJUKw7_1),.clk(gclk));
	jdff dff_B_bpVekJAE0_1(.din(w_dff_B_l2DXJUKw7_1),.dout(w_dff_B_bpVekJAE0_1),.clk(gclk));
	jdff dff_B_P0Vt5Ayd2_1(.din(w_dff_B_bpVekJAE0_1),.dout(w_dff_B_P0Vt5Ayd2_1),.clk(gclk));
	jdff dff_B_whaAqAAA6_1(.din(w_dff_B_P0Vt5Ayd2_1),.dout(w_dff_B_whaAqAAA6_1),.clk(gclk));
	jdff dff_B_CGGRfG9D1_1(.din(w_dff_B_whaAqAAA6_1),.dout(w_dff_B_CGGRfG9D1_1),.clk(gclk));
	jdff dff_B_jqOp89Qm7_1(.din(w_dff_B_CGGRfG9D1_1),.dout(w_dff_B_jqOp89Qm7_1),.clk(gclk));
	jdff dff_B_cPDyFdle6_1(.din(w_dff_B_jqOp89Qm7_1),.dout(w_dff_B_cPDyFdle6_1),.clk(gclk));
	jdff dff_B_vWgwoJ0C9_1(.din(w_dff_B_cPDyFdle6_1),.dout(w_dff_B_vWgwoJ0C9_1),.clk(gclk));
	jdff dff_B_WcWjvEIU6_1(.din(w_dff_B_vWgwoJ0C9_1),.dout(w_dff_B_WcWjvEIU6_1),.clk(gclk));
	jdff dff_B_gumcnGAx1_1(.din(w_dff_B_WcWjvEIU6_1),.dout(w_dff_B_gumcnGAx1_1),.clk(gclk));
	jdff dff_B_nBj5gObl3_1(.din(w_dff_B_gumcnGAx1_1),.dout(w_dff_B_nBj5gObl3_1),.clk(gclk));
	jdff dff_B_BYWga9r30_1(.din(w_dff_B_nBj5gObl3_1),.dout(w_dff_B_BYWga9r30_1),.clk(gclk));
	jdff dff_B_fCo7Mjhw4_1(.din(n709),.dout(w_dff_B_fCo7Mjhw4_1),.clk(gclk));
	jdff dff_A_ZJqsWTE38_0(.dout(w_n614_0[0]),.din(w_dff_A_ZJqsWTE38_0),.clk(gclk));
	jdff dff_A_DCweRg5G9_0(.dout(w_dff_A_ZJqsWTE38_0),.din(w_dff_A_DCweRg5G9_0),.clk(gclk));
	jdff dff_A_hX73WQSW0_0(.dout(w_dff_A_DCweRg5G9_0),.din(w_dff_A_hX73WQSW0_0),.clk(gclk));
	jdff dff_A_USYjXc4M0_0(.dout(w_dff_A_hX73WQSW0_0),.din(w_dff_A_USYjXc4M0_0),.clk(gclk));
	jdff dff_A_ixLA7BGJ6_0(.dout(w_dff_A_USYjXc4M0_0),.din(w_dff_A_ixLA7BGJ6_0),.clk(gclk));
	jdff dff_A_wxoBXF8s7_0(.dout(w_dff_A_ixLA7BGJ6_0),.din(w_dff_A_wxoBXF8s7_0),.clk(gclk));
	jdff dff_A_qEHhoYL80_0(.dout(w_dff_A_wxoBXF8s7_0),.din(w_dff_A_qEHhoYL80_0),.clk(gclk));
	jdff dff_A_cX3KY70c8_0(.dout(w_dff_A_qEHhoYL80_0),.din(w_dff_A_cX3KY70c8_0),.clk(gclk));
	jdff dff_A_ijblW0et0_0(.dout(w_dff_A_cX3KY70c8_0),.din(w_dff_A_ijblW0et0_0),.clk(gclk));
	jdff dff_A_O56tFSYs1_0(.dout(w_dff_A_ijblW0et0_0),.din(w_dff_A_O56tFSYs1_0),.clk(gclk));
	jdff dff_A_0qlK8UcB2_0(.dout(w_dff_A_O56tFSYs1_0),.din(w_dff_A_0qlK8UcB2_0),.clk(gclk));
	jdff dff_A_0ai6Xu861_0(.dout(w_dff_A_0qlK8UcB2_0),.din(w_dff_A_0ai6Xu861_0),.clk(gclk));
	jdff dff_A_c7qtzy478_0(.dout(w_dff_A_0ai6Xu861_0),.din(w_dff_A_c7qtzy478_0),.clk(gclk));
	jdff dff_A_WcqWStd04_0(.dout(w_dff_A_c7qtzy478_0),.din(w_dff_A_WcqWStd04_0),.clk(gclk));
	jdff dff_A_fdY2wFf83_0(.dout(w_dff_A_WcqWStd04_0),.din(w_dff_A_fdY2wFf83_0),.clk(gclk));
	jdff dff_A_iYs6F8116_0(.dout(w_dff_A_fdY2wFf83_0),.din(w_dff_A_iYs6F8116_0),.clk(gclk));
	jdff dff_A_T5gWcaLG1_0(.dout(w_dff_A_iYs6F8116_0),.din(w_dff_A_T5gWcaLG1_0),.clk(gclk));
	jdff dff_A_JudO6DsY1_0(.dout(w_dff_A_T5gWcaLG1_0),.din(w_dff_A_JudO6DsY1_0),.clk(gclk));
	jdff dff_A_poqCqyYs2_0(.dout(w_dff_A_JudO6DsY1_0),.din(w_dff_A_poqCqyYs2_0),.clk(gclk));
	jdff dff_A_su1z9E7p4_0(.dout(w_dff_A_poqCqyYs2_0),.din(w_dff_A_su1z9E7p4_0),.clk(gclk));
	jdff dff_A_fSXXNJlq9_0(.dout(w_dff_A_su1z9E7p4_0),.din(w_dff_A_fSXXNJlq9_0),.clk(gclk));
	jdff dff_A_wEsTfLSH6_0(.dout(w_dff_A_fSXXNJlq9_0),.din(w_dff_A_wEsTfLSH6_0),.clk(gclk));
	jdff dff_A_xCLZBxnn9_0(.dout(w_dff_A_wEsTfLSH6_0),.din(w_dff_A_xCLZBxnn9_0),.clk(gclk));
	jdff dff_A_ZGgbvMH67_0(.dout(w_dff_A_xCLZBxnn9_0),.din(w_dff_A_ZGgbvMH67_0),.clk(gclk));
	jdff dff_A_Sej4oIN88_0(.dout(w_dff_A_ZGgbvMH67_0),.din(w_dff_A_Sej4oIN88_0),.clk(gclk));
	jdff dff_A_oyV8gBJ34_0(.dout(w_dff_A_Sej4oIN88_0),.din(w_dff_A_oyV8gBJ34_0),.clk(gclk));
	jdff dff_A_l7rrKOUt6_0(.dout(w_dff_A_oyV8gBJ34_0),.din(w_dff_A_l7rrKOUt6_0),.clk(gclk));
	jdff dff_A_IM9QaROx9_0(.dout(w_dff_A_l7rrKOUt6_0),.din(w_dff_A_IM9QaROx9_0),.clk(gclk));
	jdff dff_A_g2VpbbBh7_0(.dout(w_dff_A_IM9QaROx9_0),.din(w_dff_A_g2VpbbBh7_0),.clk(gclk));
	jdff dff_A_cx1u4WQ89_0(.dout(w_dff_A_g2VpbbBh7_0),.din(w_dff_A_cx1u4WQ89_0),.clk(gclk));
	jdff dff_A_e7tTKAds4_0(.dout(w_dff_A_cx1u4WQ89_0),.din(w_dff_A_e7tTKAds4_0),.clk(gclk));
	jdff dff_A_XqkBEqQ31_0(.dout(w_dff_A_e7tTKAds4_0),.din(w_dff_A_XqkBEqQ31_0),.clk(gclk));
	jdff dff_A_PWjDeHci6_0(.dout(w_dff_A_XqkBEqQ31_0),.din(w_dff_A_PWjDeHci6_0),.clk(gclk));
	jdff dff_A_dY0r4lcd6_0(.dout(w_dff_A_PWjDeHci6_0),.din(w_dff_A_dY0r4lcd6_0),.clk(gclk));
	jdff dff_A_5BRhJD7N1_0(.dout(w_dff_A_dY0r4lcd6_0),.din(w_dff_A_5BRhJD7N1_0),.clk(gclk));
	jdff dff_A_vAxDeasC0_0(.dout(w_dff_A_5BRhJD7N1_0),.din(w_dff_A_vAxDeasC0_0),.clk(gclk));
	jdff dff_A_QDiMJm2D6_0(.dout(w_dff_A_vAxDeasC0_0),.din(w_dff_A_QDiMJm2D6_0),.clk(gclk));
	jdff dff_A_iUY45Q7M8_1(.dout(w_n703_0[1]),.din(w_dff_A_iUY45Q7M8_1),.clk(gclk));
	jdff dff_B_A9VAm78q2_1(.din(n621),.dout(w_dff_B_A9VAm78q2_1),.clk(gclk));
	jdff dff_B_LzmwLakx0_1(.din(w_dff_B_A9VAm78q2_1),.dout(w_dff_B_LzmwLakx0_1),.clk(gclk));
	jdff dff_B_ZSyUTwRc7_1(.din(w_dff_B_LzmwLakx0_1),.dout(w_dff_B_ZSyUTwRc7_1),.clk(gclk));
	jdff dff_B_42Ahjxve6_1(.din(w_dff_B_ZSyUTwRc7_1),.dout(w_dff_B_42Ahjxve6_1),.clk(gclk));
	jdff dff_B_WlzyMSi54_1(.din(w_dff_B_42Ahjxve6_1),.dout(w_dff_B_WlzyMSi54_1),.clk(gclk));
	jdff dff_B_2rCRDrJq6_1(.din(w_dff_B_WlzyMSi54_1),.dout(w_dff_B_2rCRDrJq6_1),.clk(gclk));
	jdff dff_B_L977e37d9_1(.din(w_dff_B_2rCRDrJq6_1),.dout(w_dff_B_L977e37d9_1),.clk(gclk));
	jdff dff_B_6CTHGhie9_1(.din(w_dff_B_L977e37d9_1),.dout(w_dff_B_6CTHGhie9_1),.clk(gclk));
	jdff dff_B_cZeONxXS9_1(.din(w_dff_B_6CTHGhie9_1),.dout(w_dff_B_cZeONxXS9_1),.clk(gclk));
	jdff dff_B_JNLUcxS15_1(.din(w_dff_B_cZeONxXS9_1),.dout(w_dff_B_JNLUcxS15_1),.clk(gclk));
	jdff dff_B_LogmgIUp3_1(.din(w_dff_B_JNLUcxS15_1),.dout(w_dff_B_LogmgIUp3_1),.clk(gclk));
	jdff dff_B_mgBfWcrG7_1(.din(w_dff_B_LogmgIUp3_1),.dout(w_dff_B_mgBfWcrG7_1),.clk(gclk));
	jdff dff_B_EumMpXXp3_1(.din(w_dff_B_mgBfWcrG7_1),.dout(w_dff_B_EumMpXXp3_1),.clk(gclk));
	jdff dff_B_7qv4UN6Y2_1(.din(w_dff_B_EumMpXXp3_1),.dout(w_dff_B_7qv4UN6Y2_1),.clk(gclk));
	jdff dff_B_gnVaiatE6_1(.din(w_dff_B_7qv4UN6Y2_1),.dout(w_dff_B_gnVaiatE6_1),.clk(gclk));
	jdff dff_B_mECXKtel3_1(.din(w_dff_B_gnVaiatE6_1),.dout(w_dff_B_mECXKtel3_1),.clk(gclk));
	jdff dff_B_MIaqtrIC0_1(.din(w_dff_B_mECXKtel3_1),.dout(w_dff_B_MIaqtrIC0_1),.clk(gclk));
	jdff dff_B_3oUq2jOq1_1(.din(w_dff_B_MIaqtrIC0_1),.dout(w_dff_B_3oUq2jOq1_1),.clk(gclk));
	jdff dff_B_zgz4uphr2_1(.din(w_dff_B_3oUq2jOq1_1),.dout(w_dff_B_zgz4uphr2_1),.clk(gclk));
	jdff dff_B_rd9DjhPC2_1(.din(w_dff_B_zgz4uphr2_1),.dout(w_dff_B_rd9DjhPC2_1),.clk(gclk));
	jdff dff_B_7AHnIwJO3_1(.din(w_dff_B_rd9DjhPC2_1),.dout(w_dff_B_7AHnIwJO3_1),.clk(gclk));
	jdff dff_B_V2fvPVmd2_1(.din(w_dff_B_7AHnIwJO3_1),.dout(w_dff_B_V2fvPVmd2_1),.clk(gclk));
	jdff dff_B_vCZDwaJ74_1(.din(w_dff_B_V2fvPVmd2_1),.dout(w_dff_B_vCZDwaJ74_1),.clk(gclk));
	jdff dff_B_qLM4d4355_1(.din(w_dff_B_vCZDwaJ74_1),.dout(w_dff_B_qLM4d4355_1),.clk(gclk));
	jdff dff_B_DwxN9Yr58_1(.din(w_dff_B_qLM4d4355_1),.dout(w_dff_B_DwxN9Yr58_1),.clk(gclk));
	jdff dff_B_00rLh3e55_1(.din(w_dff_B_DwxN9Yr58_1),.dout(w_dff_B_00rLh3e55_1),.clk(gclk));
	jdff dff_B_fYR1K5me0_1(.din(w_dff_B_00rLh3e55_1),.dout(w_dff_B_fYR1K5me0_1),.clk(gclk));
	jdff dff_B_KKRx64nL9_1(.din(w_dff_B_fYR1K5me0_1),.dout(w_dff_B_KKRx64nL9_1),.clk(gclk));
	jdff dff_B_eEHalRt61_1(.din(w_dff_B_KKRx64nL9_1),.dout(w_dff_B_eEHalRt61_1),.clk(gclk));
	jdff dff_B_vuomH4Em3_1(.din(w_dff_B_eEHalRt61_1),.dout(w_dff_B_vuomH4Em3_1),.clk(gclk));
	jdff dff_B_m0uvBwCu9_1(.din(w_dff_B_vuomH4Em3_1),.dout(w_dff_B_m0uvBwCu9_1),.clk(gclk));
	jdff dff_B_SoQs1uK54_1(.din(w_dff_B_m0uvBwCu9_1),.dout(w_dff_B_SoQs1uK54_1),.clk(gclk));
	jdff dff_B_0W0p7jUR3_1(.din(w_dff_B_SoQs1uK54_1),.dout(w_dff_B_0W0p7jUR3_1),.clk(gclk));
	jdff dff_B_ZVITaAWb1_1(.din(n617),.dout(w_dff_B_ZVITaAWb1_1),.clk(gclk));
	jdff dff_A_nhDvlxFe4_0(.dout(w_n529_0[0]),.din(w_dff_A_nhDvlxFe4_0),.clk(gclk));
	jdff dff_A_hEzlDyid1_0(.dout(w_dff_A_nhDvlxFe4_0),.din(w_dff_A_hEzlDyid1_0),.clk(gclk));
	jdff dff_A_LMN6QWFi3_0(.dout(w_dff_A_hEzlDyid1_0),.din(w_dff_A_LMN6QWFi3_0),.clk(gclk));
	jdff dff_A_zdwR896X3_0(.dout(w_dff_A_LMN6QWFi3_0),.din(w_dff_A_zdwR896X3_0),.clk(gclk));
	jdff dff_A_Cmglstuh2_0(.dout(w_dff_A_zdwR896X3_0),.din(w_dff_A_Cmglstuh2_0),.clk(gclk));
	jdff dff_A_Nl0zI5LZ5_0(.dout(w_dff_A_Cmglstuh2_0),.din(w_dff_A_Nl0zI5LZ5_0),.clk(gclk));
	jdff dff_A_RSNCOae38_0(.dout(w_dff_A_Nl0zI5LZ5_0),.din(w_dff_A_RSNCOae38_0),.clk(gclk));
	jdff dff_A_N1FfJhoA5_0(.dout(w_dff_A_RSNCOae38_0),.din(w_dff_A_N1FfJhoA5_0),.clk(gclk));
	jdff dff_A_HYh079cz5_0(.dout(w_dff_A_N1FfJhoA5_0),.din(w_dff_A_HYh079cz5_0),.clk(gclk));
	jdff dff_A_tZljyAks7_0(.dout(w_dff_A_HYh079cz5_0),.din(w_dff_A_tZljyAks7_0),.clk(gclk));
	jdff dff_A_8X8Jhouy3_0(.dout(w_dff_A_tZljyAks7_0),.din(w_dff_A_8X8Jhouy3_0),.clk(gclk));
	jdff dff_A_Gie4ZqOK9_0(.dout(w_dff_A_8X8Jhouy3_0),.din(w_dff_A_Gie4ZqOK9_0),.clk(gclk));
	jdff dff_A_xgNC3I4N5_0(.dout(w_dff_A_Gie4ZqOK9_0),.din(w_dff_A_xgNC3I4N5_0),.clk(gclk));
	jdff dff_A_iSccoqyV6_0(.dout(w_dff_A_xgNC3I4N5_0),.din(w_dff_A_iSccoqyV6_0),.clk(gclk));
	jdff dff_A_boqlekLb4_0(.dout(w_dff_A_iSccoqyV6_0),.din(w_dff_A_boqlekLb4_0),.clk(gclk));
	jdff dff_A_nOoTvesv8_0(.dout(w_dff_A_boqlekLb4_0),.din(w_dff_A_nOoTvesv8_0),.clk(gclk));
	jdff dff_A_OuPDWl9o5_0(.dout(w_dff_A_nOoTvesv8_0),.din(w_dff_A_OuPDWl9o5_0),.clk(gclk));
	jdff dff_A_IFEyOzj68_0(.dout(w_dff_A_OuPDWl9o5_0),.din(w_dff_A_IFEyOzj68_0),.clk(gclk));
	jdff dff_A_hu77U5f90_0(.dout(w_dff_A_IFEyOzj68_0),.din(w_dff_A_hu77U5f90_0),.clk(gclk));
	jdff dff_A_lIkyySYt0_0(.dout(w_dff_A_hu77U5f90_0),.din(w_dff_A_lIkyySYt0_0),.clk(gclk));
	jdff dff_A_atsADPc67_0(.dout(w_dff_A_lIkyySYt0_0),.din(w_dff_A_atsADPc67_0),.clk(gclk));
	jdff dff_A_6ZuKJLlt6_0(.dout(w_dff_A_atsADPc67_0),.din(w_dff_A_6ZuKJLlt6_0),.clk(gclk));
	jdff dff_A_w7li6z5p6_0(.dout(w_dff_A_6ZuKJLlt6_0),.din(w_dff_A_w7li6z5p6_0),.clk(gclk));
	jdff dff_A_DmifbVad4_0(.dout(w_dff_A_w7li6z5p6_0),.din(w_dff_A_DmifbVad4_0),.clk(gclk));
	jdff dff_A_PCxv85Wy7_0(.dout(w_dff_A_DmifbVad4_0),.din(w_dff_A_PCxv85Wy7_0),.clk(gclk));
	jdff dff_A_31BEGkBD1_0(.dout(w_dff_A_PCxv85Wy7_0),.din(w_dff_A_31BEGkBD1_0),.clk(gclk));
	jdff dff_A_CFjU7RDm6_0(.dout(w_dff_A_31BEGkBD1_0),.din(w_dff_A_CFjU7RDm6_0),.clk(gclk));
	jdff dff_A_2drIfCX83_0(.dout(w_dff_A_CFjU7RDm6_0),.din(w_dff_A_2drIfCX83_0),.clk(gclk));
	jdff dff_A_ek3ulER84_0(.dout(w_dff_A_2drIfCX83_0),.din(w_dff_A_ek3ulER84_0),.clk(gclk));
	jdff dff_A_IItxrOUx2_0(.dout(w_dff_A_ek3ulER84_0),.din(w_dff_A_IItxrOUx2_0),.clk(gclk));
	jdff dff_A_AMAesH8T0_0(.dout(w_dff_A_IItxrOUx2_0),.din(w_dff_A_AMAesH8T0_0),.clk(gclk));
	jdff dff_A_vIpGoxcf1_0(.dout(w_dff_A_AMAesH8T0_0),.din(w_dff_A_vIpGoxcf1_0),.clk(gclk));
	jdff dff_A_qHCW8PGe7_0(.dout(w_dff_A_vIpGoxcf1_0),.din(w_dff_A_qHCW8PGe7_0),.clk(gclk));
	jdff dff_A_bu9jZuxo2_0(.dout(w_dff_A_qHCW8PGe7_0),.din(w_dff_A_bu9jZuxo2_0),.clk(gclk));
	jdff dff_A_tWZbizCL0_1(.dout(w_n611_0[1]),.din(w_dff_A_tWZbizCL0_1),.clk(gclk));
	jdff dff_B_kCHBFrzY0_1(.din(n536),.dout(w_dff_B_kCHBFrzY0_1),.clk(gclk));
	jdff dff_B_Rd8TzzGj5_1(.din(w_dff_B_kCHBFrzY0_1),.dout(w_dff_B_Rd8TzzGj5_1),.clk(gclk));
	jdff dff_B_tENXyBbO8_1(.din(w_dff_B_Rd8TzzGj5_1),.dout(w_dff_B_tENXyBbO8_1),.clk(gclk));
	jdff dff_B_g6xqOmz25_1(.din(w_dff_B_tENXyBbO8_1),.dout(w_dff_B_g6xqOmz25_1),.clk(gclk));
	jdff dff_B_hrUXolzj6_1(.din(w_dff_B_g6xqOmz25_1),.dout(w_dff_B_hrUXolzj6_1),.clk(gclk));
	jdff dff_B_ugocssaZ4_1(.din(w_dff_B_hrUXolzj6_1),.dout(w_dff_B_ugocssaZ4_1),.clk(gclk));
	jdff dff_B_CSr6RIpv1_1(.din(w_dff_B_ugocssaZ4_1),.dout(w_dff_B_CSr6RIpv1_1),.clk(gclk));
	jdff dff_B_iBwWptcJ3_1(.din(w_dff_B_CSr6RIpv1_1),.dout(w_dff_B_iBwWptcJ3_1),.clk(gclk));
	jdff dff_B_Fj0Pwj9V7_1(.din(w_dff_B_iBwWptcJ3_1),.dout(w_dff_B_Fj0Pwj9V7_1),.clk(gclk));
	jdff dff_B_ER53Vsgq1_1(.din(w_dff_B_Fj0Pwj9V7_1),.dout(w_dff_B_ER53Vsgq1_1),.clk(gclk));
	jdff dff_B_uXHMzpMj3_1(.din(w_dff_B_ER53Vsgq1_1),.dout(w_dff_B_uXHMzpMj3_1),.clk(gclk));
	jdff dff_B_i2aGU7eZ7_1(.din(w_dff_B_uXHMzpMj3_1),.dout(w_dff_B_i2aGU7eZ7_1),.clk(gclk));
	jdff dff_B_Ko8H580d3_1(.din(w_dff_B_i2aGU7eZ7_1),.dout(w_dff_B_Ko8H580d3_1),.clk(gclk));
	jdff dff_B_qqmrnoyj5_1(.din(w_dff_B_Ko8H580d3_1),.dout(w_dff_B_qqmrnoyj5_1),.clk(gclk));
	jdff dff_B_M5TtD4UT8_1(.din(w_dff_B_qqmrnoyj5_1),.dout(w_dff_B_M5TtD4UT8_1),.clk(gclk));
	jdff dff_B_gEHEpSTY6_1(.din(w_dff_B_M5TtD4UT8_1),.dout(w_dff_B_gEHEpSTY6_1),.clk(gclk));
	jdff dff_B_p8LGoybh8_1(.din(w_dff_B_gEHEpSTY6_1),.dout(w_dff_B_p8LGoybh8_1),.clk(gclk));
	jdff dff_B_V5hUxEtK1_1(.din(w_dff_B_p8LGoybh8_1),.dout(w_dff_B_V5hUxEtK1_1),.clk(gclk));
	jdff dff_B_25lRxmGI1_1(.din(w_dff_B_V5hUxEtK1_1),.dout(w_dff_B_25lRxmGI1_1),.clk(gclk));
	jdff dff_B_IyNrAS8v8_1(.din(w_dff_B_25lRxmGI1_1),.dout(w_dff_B_IyNrAS8v8_1),.clk(gclk));
	jdff dff_B_y8CD5oan6_1(.din(w_dff_B_IyNrAS8v8_1),.dout(w_dff_B_y8CD5oan6_1),.clk(gclk));
	jdff dff_B_748Wehi27_1(.din(w_dff_B_y8CD5oan6_1),.dout(w_dff_B_748Wehi27_1),.clk(gclk));
	jdff dff_B_kh3cpPPq2_1(.din(w_dff_B_748Wehi27_1),.dout(w_dff_B_kh3cpPPq2_1),.clk(gclk));
	jdff dff_B_yOohTYGP9_1(.din(w_dff_B_kh3cpPPq2_1),.dout(w_dff_B_yOohTYGP9_1),.clk(gclk));
	jdff dff_B_FEgnCTD95_1(.din(w_dff_B_yOohTYGP9_1),.dout(w_dff_B_FEgnCTD95_1),.clk(gclk));
	jdff dff_B_AnnayLHC9_1(.din(w_dff_B_FEgnCTD95_1),.dout(w_dff_B_AnnayLHC9_1),.clk(gclk));
	jdff dff_B_Uyh8CFlP1_1(.din(w_dff_B_AnnayLHC9_1),.dout(w_dff_B_Uyh8CFlP1_1),.clk(gclk));
	jdff dff_B_fq7cDSzQ7_1(.din(w_dff_B_Uyh8CFlP1_1),.dout(w_dff_B_fq7cDSzQ7_1),.clk(gclk));
	jdff dff_B_9mT4DgtD6_1(.din(w_dff_B_fq7cDSzQ7_1),.dout(w_dff_B_9mT4DgtD6_1),.clk(gclk));
	jdff dff_B_vR0plZ4L4_1(.din(w_dff_B_9mT4DgtD6_1),.dout(w_dff_B_vR0plZ4L4_1),.clk(gclk));
	jdff dff_B_VXK70yMo3_1(.din(n532),.dout(w_dff_B_VXK70yMo3_1),.clk(gclk));
	jdff dff_A_OTZF4ZFo9_0(.dout(w_n451_0[0]),.din(w_dff_A_OTZF4ZFo9_0),.clk(gclk));
	jdff dff_A_Cb8ck3cf5_0(.dout(w_dff_A_OTZF4ZFo9_0),.din(w_dff_A_Cb8ck3cf5_0),.clk(gclk));
	jdff dff_A_N3kcUESC7_0(.dout(w_dff_A_Cb8ck3cf5_0),.din(w_dff_A_N3kcUESC7_0),.clk(gclk));
	jdff dff_A_fBeDrGu99_0(.dout(w_dff_A_N3kcUESC7_0),.din(w_dff_A_fBeDrGu99_0),.clk(gclk));
	jdff dff_A_hHwR3u782_0(.dout(w_dff_A_fBeDrGu99_0),.din(w_dff_A_hHwR3u782_0),.clk(gclk));
	jdff dff_A_AUvVvqXm5_0(.dout(w_dff_A_hHwR3u782_0),.din(w_dff_A_AUvVvqXm5_0),.clk(gclk));
	jdff dff_A_OSAg4mRU4_0(.dout(w_dff_A_AUvVvqXm5_0),.din(w_dff_A_OSAg4mRU4_0),.clk(gclk));
	jdff dff_A_hSXfgab13_0(.dout(w_dff_A_OSAg4mRU4_0),.din(w_dff_A_hSXfgab13_0),.clk(gclk));
	jdff dff_A_aVSZUbVy0_0(.dout(w_dff_A_hSXfgab13_0),.din(w_dff_A_aVSZUbVy0_0),.clk(gclk));
	jdff dff_A_tZZZ0Cgd1_0(.dout(w_dff_A_aVSZUbVy0_0),.din(w_dff_A_tZZZ0Cgd1_0),.clk(gclk));
	jdff dff_A_a4zs17Eo1_0(.dout(w_dff_A_tZZZ0Cgd1_0),.din(w_dff_A_a4zs17Eo1_0),.clk(gclk));
	jdff dff_A_GcPPHrYn8_0(.dout(w_dff_A_a4zs17Eo1_0),.din(w_dff_A_GcPPHrYn8_0),.clk(gclk));
	jdff dff_A_vJB0qnwq9_0(.dout(w_dff_A_GcPPHrYn8_0),.din(w_dff_A_vJB0qnwq9_0),.clk(gclk));
	jdff dff_A_pfhOpkfR0_0(.dout(w_dff_A_vJB0qnwq9_0),.din(w_dff_A_pfhOpkfR0_0),.clk(gclk));
	jdff dff_A_2QKP8nLj5_0(.dout(w_dff_A_pfhOpkfR0_0),.din(w_dff_A_2QKP8nLj5_0),.clk(gclk));
	jdff dff_A_lhi8bUCk6_0(.dout(w_dff_A_2QKP8nLj5_0),.din(w_dff_A_lhi8bUCk6_0),.clk(gclk));
	jdff dff_A_n9iK2LAY2_0(.dout(w_dff_A_lhi8bUCk6_0),.din(w_dff_A_n9iK2LAY2_0),.clk(gclk));
	jdff dff_A_pCPGAd0k0_0(.dout(w_dff_A_n9iK2LAY2_0),.din(w_dff_A_pCPGAd0k0_0),.clk(gclk));
	jdff dff_A_AdIacxm98_0(.dout(w_dff_A_pCPGAd0k0_0),.din(w_dff_A_AdIacxm98_0),.clk(gclk));
	jdff dff_A_wi5K90kP1_0(.dout(w_dff_A_AdIacxm98_0),.din(w_dff_A_wi5K90kP1_0),.clk(gclk));
	jdff dff_A_OzyeiJQp1_0(.dout(w_dff_A_wi5K90kP1_0),.din(w_dff_A_OzyeiJQp1_0),.clk(gclk));
	jdff dff_A_IzGg7SBo5_0(.dout(w_dff_A_OzyeiJQp1_0),.din(w_dff_A_IzGg7SBo5_0),.clk(gclk));
	jdff dff_A_1tXWoT3N0_0(.dout(w_dff_A_IzGg7SBo5_0),.din(w_dff_A_1tXWoT3N0_0),.clk(gclk));
	jdff dff_A_Yhmi73pX0_0(.dout(w_dff_A_1tXWoT3N0_0),.din(w_dff_A_Yhmi73pX0_0),.clk(gclk));
	jdff dff_A_HW5x8sja4_0(.dout(w_dff_A_Yhmi73pX0_0),.din(w_dff_A_HW5x8sja4_0),.clk(gclk));
	jdff dff_A_JCaxpzaX2_0(.dout(w_dff_A_HW5x8sja4_0),.din(w_dff_A_JCaxpzaX2_0),.clk(gclk));
	jdff dff_A_79MTMddy7_0(.dout(w_dff_A_JCaxpzaX2_0),.din(w_dff_A_79MTMddy7_0),.clk(gclk));
	jdff dff_A_bvmvRzxa6_0(.dout(w_dff_A_79MTMddy7_0),.din(w_dff_A_bvmvRzxa6_0),.clk(gclk));
	jdff dff_A_56tZM1Q22_0(.dout(w_dff_A_bvmvRzxa6_0),.din(w_dff_A_56tZM1Q22_0),.clk(gclk));
	jdff dff_A_90ofgxfk4_0(.dout(w_dff_A_56tZM1Q22_0),.din(w_dff_A_90ofgxfk4_0),.clk(gclk));
	jdff dff_A_ERRIE9kX2_0(.dout(w_dff_A_90ofgxfk4_0),.din(w_dff_A_ERRIE9kX2_0),.clk(gclk));
	jdff dff_A_kiwmOoXQ4_1(.dout(w_n526_0[1]),.din(w_dff_A_kiwmOoXQ4_1),.clk(gclk));
	jdff dff_B_zBMuKWgD3_1(.din(n458),.dout(w_dff_B_zBMuKWgD3_1),.clk(gclk));
	jdff dff_B_DnZAdYla3_1(.din(w_dff_B_zBMuKWgD3_1),.dout(w_dff_B_DnZAdYla3_1),.clk(gclk));
	jdff dff_B_R4Ar9KN49_1(.din(w_dff_B_DnZAdYla3_1),.dout(w_dff_B_R4Ar9KN49_1),.clk(gclk));
	jdff dff_B_KcFTeE4h5_1(.din(w_dff_B_R4Ar9KN49_1),.dout(w_dff_B_KcFTeE4h5_1),.clk(gclk));
	jdff dff_B_RXR5pRJ54_1(.din(w_dff_B_KcFTeE4h5_1),.dout(w_dff_B_RXR5pRJ54_1),.clk(gclk));
	jdff dff_B_G6ai8QNX2_1(.din(w_dff_B_RXR5pRJ54_1),.dout(w_dff_B_G6ai8QNX2_1),.clk(gclk));
	jdff dff_B_LTqYmLE73_1(.din(w_dff_B_G6ai8QNX2_1),.dout(w_dff_B_LTqYmLE73_1),.clk(gclk));
	jdff dff_B_c7cHTrDQ1_1(.din(w_dff_B_LTqYmLE73_1),.dout(w_dff_B_c7cHTrDQ1_1),.clk(gclk));
	jdff dff_B_vwTbbMfu9_1(.din(w_dff_B_c7cHTrDQ1_1),.dout(w_dff_B_vwTbbMfu9_1),.clk(gclk));
	jdff dff_B_qzxyu0aN4_1(.din(w_dff_B_vwTbbMfu9_1),.dout(w_dff_B_qzxyu0aN4_1),.clk(gclk));
	jdff dff_B_HIYPKxAn3_1(.din(w_dff_B_qzxyu0aN4_1),.dout(w_dff_B_HIYPKxAn3_1),.clk(gclk));
	jdff dff_B_jU9d4w7i2_1(.din(w_dff_B_HIYPKxAn3_1),.dout(w_dff_B_jU9d4w7i2_1),.clk(gclk));
	jdff dff_B_4z6oZ8he6_1(.din(w_dff_B_jU9d4w7i2_1),.dout(w_dff_B_4z6oZ8he6_1),.clk(gclk));
	jdff dff_B_XvF1Glm41_1(.din(w_dff_B_4z6oZ8he6_1),.dout(w_dff_B_XvF1Glm41_1),.clk(gclk));
	jdff dff_B_zXNSOptH7_1(.din(w_dff_B_XvF1Glm41_1),.dout(w_dff_B_zXNSOptH7_1),.clk(gclk));
	jdff dff_B_otfm0FSw6_1(.din(w_dff_B_zXNSOptH7_1),.dout(w_dff_B_otfm0FSw6_1),.clk(gclk));
	jdff dff_B_8O76r0r17_1(.din(w_dff_B_otfm0FSw6_1),.dout(w_dff_B_8O76r0r17_1),.clk(gclk));
	jdff dff_B_UUJVWsuS2_1(.din(w_dff_B_8O76r0r17_1),.dout(w_dff_B_UUJVWsuS2_1),.clk(gclk));
	jdff dff_B_FF4VzAs23_1(.din(w_dff_B_UUJVWsuS2_1),.dout(w_dff_B_FF4VzAs23_1),.clk(gclk));
	jdff dff_B_WsWMziBW5_1(.din(w_dff_B_FF4VzAs23_1),.dout(w_dff_B_WsWMziBW5_1),.clk(gclk));
	jdff dff_B_Hwa1W5oB3_1(.din(w_dff_B_WsWMziBW5_1),.dout(w_dff_B_Hwa1W5oB3_1),.clk(gclk));
	jdff dff_B_uyrPcFlQ2_1(.din(w_dff_B_Hwa1W5oB3_1),.dout(w_dff_B_uyrPcFlQ2_1),.clk(gclk));
	jdff dff_B_ODTl2ZlX6_1(.din(w_dff_B_uyrPcFlQ2_1),.dout(w_dff_B_ODTl2ZlX6_1),.clk(gclk));
	jdff dff_B_Ak0VIRh19_1(.din(w_dff_B_ODTl2ZlX6_1),.dout(w_dff_B_Ak0VIRh19_1),.clk(gclk));
	jdff dff_B_YezfJTEd4_1(.din(w_dff_B_Ak0VIRh19_1),.dout(w_dff_B_YezfJTEd4_1),.clk(gclk));
	jdff dff_B_YrzUY8kt2_1(.din(w_dff_B_YezfJTEd4_1),.dout(w_dff_B_YrzUY8kt2_1),.clk(gclk));
	jdff dff_B_YUvxqxm79_1(.din(w_dff_B_YrzUY8kt2_1),.dout(w_dff_B_YUvxqxm79_1),.clk(gclk));
	jdff dff_B_LJWEIvt20_1(.din(n454),.dout(w_dff_B_LJWEIvt20_1),.clk(gclk));
	jdff dff_A_xFbdq81z3_0(.dout(w_n380_0[0]),.din(w_dff_A_xFbdq81z3_0),.clk(gclk));
	jdff dff_A_FCQ7mtkf0_0(.dout(w_dff_A_xFbdq81z3_0),.din(w_dff_A_FCQ7mtkf0_0),.clk(gclk));
	jdff dff_A_FEfsb2Wf5_0(.dout(w_dff_A_FCQ7mtkf0_0),.din(w_dff_A_FEfsb2Wf5_0),.clk(gclk));
	jdff dff_A_Ri2JnhyP2_0(.dout(w_dff_A_FEfsb2Wf5_0),.din(w_dff_A_Ri2JnhyP2_0),.clk(gclk));
	jdff dff_A_RVueaT9M4_0(.dout(w_dff_A_Ri2JnhyP2_0),.din(w_dff_A_RVueaT9M4_0),.clk(gclk));
	jdff dff_A_6peDFwnx9_0(.dout(w_dff_A_RVueaT9M4_0),.din(w_dff_A_6peDFwnx9_0),.clk(gclk));
	jdff dff_A_4aofisUd7_0(.dout(w_dff_A_6peDFwnx9_0),.din(w_dff_A_4aofisUd7_0),.clk(gclk));
	jdff dff_A_7GCzgXLn8_0(.dout(w_dff_A_4aofisUd7_0),.din(w_dff_A_7GCzgXLn8_0),.clk(gclk));
	jdff dff_A_SRM2ThGz5_0(.dout(w_dff_A_7GCzgXLn8_0),.din(w_dff_A_SRM2ThGz5_0),.clk(gclk));
	jdff dff_A_Gqg9NpGL7_0(.dout(w_dff_A_SRM2ThGz5_0),.din(w_dff_A_Gqg9NpGL7_0),.clk(gclk));
	jdff dff_A_TpbmBRl95_0(.dout(w_dff_A_Gqg9NpGL7_0),.din(w_dff_A_TpbmBRl95_0),.clk(gclk));
	jdff dff_A_Nmm34HsN3_0(.dout(w_dff_A_TpbmBRl95_0),.din(w_dff_A_Nmm34HsN3_0),.clk(gclk));
	jdff dff_A_qz0O7cJg1_0(.dout(w_dff_A_Nmm34HsN3_0),.din(w_dff_A_qz0O7cJg1_0),.clk(gclk));
	jdff dff_A_t4KNzypt8_0(.dout(w_dff_A_qz0O7cJg1_0),.din(w_dff_A_t4KNzypt8_0),.clk(gclk));
	jdff dff_A_HYwUUR276_0(.dout(w_dff_A_t4KNzypt8_0),.din(w_dff_A_HYwUUR276_0),.clk(gclk));
	jdff dff_A_UADPqvIj5_0(.dout(w_dff_A_HYwUUR276_0),.din(w_dff_A_UADPqvIj5_0),.clk(gclk));
	jdff dff_A_RzRk2Cvz2_0(.dout(w_dff_A_UADPqvIj5_0),.din(w_dff_A_RzRk2Cvz2_0),.clk(gclk));
	jdff dff_A_TulId1XP1_0(.dout(w_dff_A_RzRk2Cvz2_0),.din(w_dff_A_TulId1XP1_0),.clk(gclk));
	jdff dff_A_z1uLUdZy3_0(.dout(w_dff_A_TulId1XP1_0),.din(w_dff_A_z1uLUdZy3_0),.clk(gclk));
	jdff dff_A_kiJJroz33_0(.dout(w_dff_A_z1uLUdZy3_0),.din(w_dff_A_kiJJroz33_0),.clk(gclk));
	jdff dff_A_niUUt0470_0(.dout(w_dff_A_kiJJroz33_0),.din(w_dff_A_niUUt0470_0),.clk(gclk));
	jdff dff_A_G00qHLd81_0(.dout(w_dff_A_niUUt0470_0),.din(w_dff_A_G00qHLd81_0),.clk(gclk));
	jdff dff_A_X0F482pz5_0(.dout(w_dff_A_G00qHLd81_0),.din(w_dff_A_X0F482pz5_0),.clk(gclk));
	jdff dff_A_MCwLeiD24_0(.dout(w_dff_A_X0F482pz5_0),.din(w_dff_A_MCwLeiD24_0),.clk(gclk));
	jdff dff_A_7H8fdpvx4_0(.dout(w_dff_A_MCwLeiD24_0),.din(w_dff_A_7H8fdpvx4_0),.clk(gclk));
	jdff dff_A_QCgajTaP8_0(.dout(w_dff_A_7H8fdpvx4_0),.din(w_dff_A_QCgajTaP8_0),.clk(gclk));
	jdff dff_A_Cffrl4qT1_0(.dout(w_dff_A_QCgajTaP8_0),.din(w_dff_A_Cffrl4qT1_0),.clk(gclk));
	jdff dff_A_mhHgcLc15_0(.dout(w_dff_A_Cffrl4qT1_0),.din(w_dff_A_mhHgcLc15_0),.clk(gclk));
	jdff dff_A_RSzIhc3H1_1(.dout(w_n448_0[1]),.din(w_dff_A_RSzIhc3H1_1),.clk(gclk));
	jdff dff_B_8IzsM0oD3_1(.din(n387),.dout(w_dff_B_8IzsM0oD3_1),.clk(gclk));
	jdff dff_B_jL7slHTw7_1(.din(w_dff_B_8IzsM0oD3_1),.dout(w_dff_B_jL7slHTw7_1),.clk(gclk));
	jdff dff_B_MxMOhbsl4_1(.din(w_dff_B_jL7slHTw7_1),.dout(w_dff_B_MxMOhbsl4_1),.clk(gclk));
	jdff dff_B_kYRKIEJe8_1(.din(w_dff_B_MxMOhbsl4_1),.dout(w_dff_B_kYRKIEJe8_1),.clk(gclk));
	jdff dff_B_AzhsXSAm8_1(.din(w_dff_B_kYRKIEJe8_1),.dout(w_dff_B_AzhsXSAm8_1),.clk(gclk));
	jdff dff_B_l27U4c4U9_1(.din(w_dff_B_AzhsXSAm8_1),.dout(w_dff_B_l27U4c4U9_1),.clk(gclk));
	jdff dff_B_Y2BR2rwX8_1(.din(w_dff_B_l27U4c4U9_1),.dout(w_dff_B_Y2BR2rwX8_1),.clk(gclk));
	jdff dff_B_dQ7RhL0j2_1(.din(w_dff_B_Y2BR2rwX8_1),.dout(w_dff_B_dQ7RhL0j2_1),.clk(gclk));
	jdff dff_B_M3EBURiR6_1(.din(w_dff_B_dQ7RhL0j2_1),.dout(w_dff_B_M3EBURiR6_1),.clk(gclk));
	jdff dff_B_wBDy8Uej1_1(.din(w_dff_B_M3EBURiR6_1),.dout(w_dff_B_wBDy8Uej1_1),.clk(gclk));
	jdff dff_B_DVoJ7zCR3_1(.din(w_dff_B_wBDy8Uej1_1),.dout(w_dff_B_DVoJ7zCR3_1),.clk(gclk));
	jdff dff_B_S9ZaIGoN3_1(.din(w_dff_B_DVoJ7zCR3_1),.dout(w_dff_B_S9ZaIGoN3_1),.clk(gclk));
	jdff dff_B_mc7YIRdA1_1(.din(w_dff_B_S9ZaIGoN3_1),.dout(w_dff_B_mc7YIRdA1_1),.clk(gclk));
	jdff dff_B_ci266ybB5_1(.din(w_dff_B_mc7YIRdA1_1),.dout(w_dff_B_ci266ybB5_1),.clk(gclk));
	jdff dff_B_UWT8ro7g5_1(.din(w_dff_B_ci266ybB5_1),.dout(w_dff_B_UWT8ro7g5_1),.clk(gclk));
	jdff dff_B_QskdNfw20_1(.din(w_dff_B_UWT8ro7g5_1),.dout(w_dff_B_QskdNfw20_1),.clk(gclk));
	jdff dff_B_75B13Y7W2_1(.din(w_dff_B_QskdNfw20_1),.dout(w_dff_B_75B13Y7W2_1),.clk(gclk));
	jdff dff_B_Ag1D4aU29_1(.din(w_dff_B_75B13Y7W2_1),.dout(w_dff_B_Ag1D4aU29_1),.clk(gclk));
	jdff dff_B_15cdKQOx4_1(.din(w_dff_B_Ag1D4aU29_1),.dout(w_dff_B_15cdKQOx4_1),.clk(gclk));
	jdff dff_B_5Sw6A1Cq3_1(.din(w_dff_B_15cdKQOx4_1),.dout(w_dff_B_5Sw6A1Cq3_1),.clk(gclk));
	jdff dff_B_7SAOGW3R3_1(.din(w_dff_B_5Sw6A1Cq3_1),.dout(w_dff_B_7SAOGW3R3_1),.clk(gclk));
	jdff dff_B_vMg1hHGn4_1(.din(w_dff_B_7SAOGW3R3_1),.dout(w_dff_B_vMg1hHGn4_1),.clk(gclk));
	jdff dff_B_BGqwVxJj0_1(.din(w_dff_B_vMg1hHGn4_1),.dout(w_dff_B_BGqwVxJj0_1),.clk(gclk));
	jdff dff_B_o39bPTKi1_1(.din(w_dff_B_BGqwVxJj0_1),.dout(w_dff_B_o39bPTKi1_1),.clk(gclk));
	jdff dff_B_qUFUEihJ6_1(.din(n383),.dout(w_dff_B_qUFUEihJ6_1),.clk(gclk));
	jdff dff_A_6OLEzaXf3_0(.dout(w_n317_0[0]),.din(w_dff_A_6OLEzaXf3_0),.clk(gclk));
	jdff dff_A_eY119YXw3_0(.dout(w_dff_A_6OLEzaXf3_0),.din(w_dff_A_eY119YXw3_0),.clk(gclk));
	jdff dff_A_n9av7IQb4_0(.dout(w_dff_A_eY119YXw3_0),.din(w_dff_A_n9av7IQb4_0),.clk(gclk));
	jdff dff_A_auMVzTH99_0(.dout(w_dff_A_n9av7IQb4_0),.din(w_dff_A_auMVzTH99_0),.clk(gclk));
	jdff dff_A_XrQEAPYG6_0(.dout(w_dff_A_auMVzTH99_0),.din(w_dff_A_XrQEAPYG6_0),.clk(gclk));
	jdff dff_A_0nzDlDOa0_0(.dout(w_dff_A_XrQEAPYG6_0),.din(w_dff_A_0nzDlDOa0_0),.clk(gclk));
	jdff dff_A_eSBgJxCX8_0(.dout(w_dff_A_0nzDlDOa0_0),.din(w_dff_A_eSBgJxCX8_0),.clk(gclk));
	jdff dff_A_Ila1lE2m4_0(.dout(w_dff_A_eSBgJxCX8_0),.din(w_dff_A_Ila1lE2m4_0),.clk(gclk));
	jdff dff_A_WKUXKNJR6_0(.dout(w_dff_A_Ila1lE2m4_0),.din(w_dff_A_WKUXKNJR6_0),.clk(gclk));
	jdff dff_A_8xVbUGRS1_0(.dout(w_dff_A_WKUXKNJR6_0),.din(w_dff_A_8xVbUGRS1_0),.clk(gclk));
	jdff dff_A_MJZC7UVW9_0(.dout(w_dff_A_8xVbUGRS1_0),.din(w_dff_A_MJZC7UVW9_0),.clk(gclk));
	jdff dff_A_P7rHvVYo6_0(.dout(w_dff_A_MJZC7UVW9_0),.din(w_dff_A_P7rHvVYo6_0),.clk(gclk));
	jdff dff_A_c9UHDsyl7_0(.dout(w_dff_A_P7rHvVYo6_0),.din(w_dff_A_c9UHDsyl7_0),.clk(gclk));
	jdff dff_A_ERqEylzL4_0(.dout(w_dff_A_c9UHDsyl7_0),.din(w_dff_A_ERqEylzL4_0),.clk(gclk));
	jdff dff_A_MJGTWWdj1_0(.dout(w_dff_A_ERqEylzL4_0),.din(w_dff_A_MJGTWWdj1_0),.clk(gclk));
	jdff dff_A_U95dLSqh6_0(.dout(w_dff_A_MJGTWWdj1_0),.din(w_dff_A_U95dLSqh6_0),.clk(gclk));
	jdff dff_A_G2zgbwfV5_0(.dout(w_dff_A_U95dLSqh6_0),.din(w_dff_A_G2zgbwfV5_0),.clk(gclk));
	jdff dff_A_o2RSMPzA4_0(.dout(w_dff_A_G2zgbwfV5_0),.din(w_dff_A_o2RSMPzA4_0),.clk(gclk));
	jdff dff_A_RXOCSMT92_0(.dout(w_dff_A_o2RSMPzA4_0),.din(w_dff_A_RXOCSMT92_0),.clk(gclk));
	jdff dff_A_WtEesyWf0_0(.dout(w_dff_A_RXOCSMT92_0),.din(w_dff_A_WtEesyWf0_0),.clk(gclk));
	jdff dff_A_vDLIzGEw7_0(.dout(w_dff_A_WtEesyWf0_0),.din(w_dff_A_vDLIzGEw7_0),.clk(gclk));
	jdff dff_A_WCsDVMnX1_0(.dout(w_dff_A_vDLIzGEw7_0),.din(w_dff_A_WCsDVMnX1_0),.clk(gclk));
	jdff dff_A_6vSefmfV5_0(.dout(w_dff_A_WCsDVMnX1_0),.din(w_dff_A_6vSefmfV5_0),.clk(gclk));
	jdff dff_A_7HWt21FX3_0(.dout(w_dff_A_6vSefmfV5_0),.din(w_dff_A_7HWt21FX3_0),.clk(gclk));
	jdff dff_A_k1BBpuyE8_0(.dout(w_dff_A_7HWt21FX3_0),.din(w_dff_A_k1BBpuyE8_0),.clk(gclk));
	jdff dff_A_Bovu7nZx1_1(.dout(w_n377_0[1]),.din(w_dff_A_Bovu7nZx1_1),.clk(gclk));
	jdff dff_B_e8GjJcCW9_1(.din(n324),.dout(w_dff_B_e8GjJcCW9_1),.clk(gclk));
	jdff dff_B_BuGj6LmC7_1(.din(w_dff_B_e8GjJcCW9_1),.dout(w_dff_B_BuGj6LmC7_1),.clk(gclk));
	jdff dff_B_RqGqG74g8_1(.din(w_dff_B_BuGj6LmC7_1),.dout(w_dff_B_RqGqG74g8_1),.clk(gclk));
	jdff dff_B_WImsQgUi5_1(.din(w_dff_B_RqGqG74g8_1),.dout(w_dff_B_WImsQgUi5_1),.clk(gclk));
	jdff dff_B_vF7Lls0q3_1(.din(w_dff_B_WImsQgUi5_1),.dout(w_dff_B_vF7Lls0q3_1),.clk(gclk));
	jdff dff_B_Gy6lrtYG3_1(.din(w_dff_B_vF7Lls0q3_1),.dout(w_dff_B_Gy6lrtYG3_1),.clk(gclk));
	jdff dff_B_eKfU6hzp1_1(.din(w_dff_B_Gy6lrtYG3_1),.dout(w_dff_B_eKfU6hzp1_1),.clk(gclk));
	jdff dff_B_yndFDEJi3_1(.din(w_dff_B_eKfU6hzp1_1),.dout(w_dff_B_yndFDEJi3_1),.clk(gclk));
	jdff dff_B_sbJdPLQ23_1(.din(w_dff_B_yndFDEJi3_1),.dout(w_dff_B_sbJdPLQ23_1),.clk(gclk));
	jdff dff_B_ibPIAYSx6_1(.din(w_dff_B_sbJdPLQ23_1),.dout(w_dff_B_ibPIAYSx6_1),.clk(gclk));
	jdff dff_B_feS9UsVx4_1(.din(w_dff_B_ibPIAYSx6_1),.dout(w_dff_B_feS9UsVx4_1),.clk(gclk));
	jdff dff_B_FurDQtN38_1(.din(w_dff_B_feS9UsVx4_1),.dout(w_dff_B_FurDQtN38_1),.clk(gclk));
	jdff dff_B_5HMl790y2_1(.din(w_dff_B_FurDQtN38_1),.dout(w_dff_B_5HMl790y2_1),.clk(gclk));
	jdff dff_B_jyvY51ll4_1(.din(w_dff_B_5HMl790y2_1),.dout(w_dff_B_jyvY51ll4_1),.clk(gclk));
	jdff dff_B_td2FHD193_1(.din(w_dff_B_jyvY51ll4_1),.dout(w_dff_B_td2FHD193_1),.clk(gclk));
	jdff dff_B_KbefJUfY2_1(.din(w_dff_B_td2FHD193_1),.dout(w_dff_B_KbefJUfY2_1),.clk(gclk));
	jdff dff_B_eBGwZBbY3_1(.din(w_dff_B_KbefJUfY2_1),.dout(w_dff_B_eBGwZBbY3_1),.clk(gclk));
	jdff dff_B_WzNbvo4m5_1(.din(w_dff_B_eBGwZBbY3_1),.dout(w_dff_B_WzNbvo4m5_1),.clk(gclk));
	jdff dff_B_1d3JgBps1_1(.din(w_dff_B_WzNbvo4m5_1),.dout(w_dff_B_1d3JgBps1_1),.clk(gclk));
	jdff dff_B_oEH0J9py3_1(.din(w_dff_B_1d3JgBps1_1),.dout(w_dff_B_oEH0J9py3_1),.clk(gclk));
	jdff dff_B_Y7eTPMcT7_1(.din(w_dff_B_oEH0J9py3_1),.dout(w_dff_B_Y7eTPMcT7_1),.clk(gclk));
	jdff dff_B_P7NpbNA11_1(.din(n320),.dout(w_dff_B_P7NpbNA11_1),.clk(gclk));
	jdff dff_A_D0Qidzpm9_0(.dout(w_n261_0[0]),.din(w_dff_A_D0Qidzpm9_0),.clk(gclk));
	jdff dff_A_yMczb0lx9_0(.dout(w_dff_A_D0Qidzpm9_0),.din(w_dff_A_yMczb0lx9_0),.clk(gclk));
	jdff dff_A_DMy0DIpY8_0(.dout(w_dff_A_yMczb0lx9_0),.din(w_dff_A_DMy0DIpY8_0),.clk(gclk));
	jdff dff_A_oiy70Ye71_0(.dout(w_dff_A_DMy0DIpY8_0),.din(w_dff_A_oiy70Ye71_0),.clk(gclk));
	jdff dff_A_V1h4Rjwg7_0(.dout(w_dff_A_oiy70Ye71_0),.din(w_dff_A_V1h4Rjwg7_0),.clk(gclk));
	jdff dff_A_CWeX05oF3_0(.dout(w_dff_A_V1h4Rjwg7_0),.din(w_dff_A_CWeX05oF3_0),.clk(gclk));
	jdff dff_A_5qC8yfzW7_0(.dout(w_dff_A_CWeX05oF3_0),.din(w_dff_A_5qC8yfzW7_0),.clk(gclk));
	jdff dff_A_13OJlsHp3_0(.dout(w_dff_A_5qC8yfzW7_0),.din(w_dff_A_13OJlsHp3_0),.clk(gclk));
	jdff dff_A_h5S33M530_0(.dout(w_dff_A_13OJlsHp3_0),.din(w_dff_A_h5S33M530_0),.clk(gclk));
	jdff dff_A_poXiEqOV4_0(.dout(w_dff_A_h5S33M530_0),.din(w_dff_A_poXiEqOV4_0),.clk(gclk));
	jdff dff_A_5kNhbh6y7_0(.dout(w_dff_A_poXiEqOV4_0),.din(w_dff_A_5kNhbh6y7_0),.clk(gclk));
	jdff dff_A_e8JIFoMd9_0(.dout(w_dff_A_5kNhbh6y7_0),.din(w_dff_A_e8JIFoMd9_0),.clk(gclk));
	jdff dff_A_9EEJxgeo5_0(.dout(w_dff_A_e8JIFoMd9_0),.din(w_dff_A_9EEJxgeo5_0),.clk(gclk));
	jdff dff_A_ZOgyuoVn7_0(.dout(w_dff_A_9EEJxgeo5_0),.din(w_dff_A_ZOgyuoVn7_0),.clk(gclk));
	jdff dff_A_Cf2f3QFx5_0(.dout(w_dff_A_ZOgyuoVn7_0),.din(w_dff_A_Cf2f3QFx5_0),.clk(gclk));
	jdff dff_A_zvRImTZy9_0(.dout(w_dff_A_Cf2f3QFx5_0),.din(w_dff_A_zvRImTZy9_0),.clk(gclk));
	jdff dff_A_D6LMTFrW8_0(.dout(w_dff_A_zvRImTZy9_0),.din(w_dff_A_D6LMTFrW8_0),.clk(gclk));
	jdff dff_A_k7yBVQ1b5_0(.dout(w_dff_A_D6LMTFrW8_0),.din(w_dff_A_k7yBVQ1b5_0),.clk(gclk));
	jdff dff_A_r7j8Heqh9_0(.dout(w_dff_A_k7yBVQ1b5_0),.din(w_dff_A_r7j8Heqh9_0),.clk(gclk));
	jdff dff_A_Hn8yPNAj3_0(.dout(w_dff_A_r7j8Heqh9_0),.din(w_dff_A_Hn8yPNAj3_0),.clk(gclk));
	jdff dff_A_HRlk4xJI7_0(.dout(w_dff_A_Hn8yPNAj3_0),.din(w_dff_A_HRlk4xJI7_0),.clk(gclk));
	jdff dff_A_MScdtDYV3_0(.dout(w_dff_A_HRlk4xJI7_0),.din(w_dff_A_MScdtDYV3_0),.clk(gclk));
	jdff dff_A_z1v3IO1U1_1(.dout(w_n314_0[1]),.din(w_dff_A_z1v3IO1U1_1),.clk(gclk));
	jdff dff_B_OatZHRhl5_1(.din(n268),.dout(w_dff_B_OatZHRhl5_1),.clk(gclk));
	jdff dff_B_E2m2I4tc4_1(.din(w_dff_B_OatZHRhl5_1),.dout(w_dff_B_E2m2I4tc4_1),.clk(gclk));
	jdff dff_B_chenxPSq4_1(.din(w_dff_B_E2m2I4tc4_1),.dout(w_dff_B_chenxPSq4_1),.clk(gclk));
	jdff dff_B_J1Ave9H68_1(.din(w_dff_B_chenxPSq4_1),.dout(w_dff_B_J1Ave9H68_1),.clk(gclk));
	jdff dff_B_AnLyatS00_1(.din(w_dff_B_J1Ave9H68_1),.dout(w_dff_B_AnLyatS00_1),.clk(gclk));
	jdff dff_B_FhbxRMqo2_1(.din(w_dff_B_AnLyatS00_1),.dout(w_dff_B_FhbxRMqo2_1),.clk(gclk));
	jdff dff_B_Nns16vPM0_1(.din(w_dff_B_FhbxRMqo2_1),.dout(w_dff_B_Nns16vPM0_1),.clk(gclk));
	jdff dff_B_XjGdVqET9_1(.din(w_dff_B_Nns16vPM0_1),.dout(w_dff_B_XjGdVqET9_1),.clk(gclk));
	jdff dff_B_GfNLBomx2_1(.din(w_dff_B_XjGdVqET9_1),.dout(w_dff_B_GfNLBomx2_1),.clk(gclk));
	jdff dff_B_EwLD71nM2_1(.din(w_dff_B_GfNLBomx2_1),.dout(w_dff_B_EwLD71nM2_1),.clk(gclk));
	jdff dff_B_zMiVHBW53_1(.din(w_dff_B_EwLD71nM2_1),.dout(w_dff_B_zMiVHBW53_1),.clk(gclk));
	jdff dff_B_6Z095BjI0_1(.din(w_dff_B_zMiVHBW53_1),.dout(w_dff_B_6Z095BjI0_1),.clk(gclk));
	jdff dff_B_DZPrepAl3_1(.din(w_dff_B_6Z095BjI0_1),.dout(w_dff_B_DZPrepAl3_1),.clk(gclk));
	jdff dff_B_xkW8tMkH8_1(.din(w_dff_B_DZPrepAl3_1),.dout(w_dff_B_xkW8tMkH8_1),.clk(gclk));
	jdff dff_B_ZkP7TBDr9_1(.din(w_dff_B_xkW8tMkH8_1),.dout(w_dff_B_ZkP7TBDr9_1),.clk(gclk));
	jdff dff_B_LQ6f3UFc1_1(.din(w_dff_B_ZkP7TBDr9_1),.dout(w_dff_B_LQ6f3UFc1_1),.clk(gclk));
	jdff dff_B_odZ837622_1(.din(w_dff_B_LQ6f3UFc1_1),.dout(w_dff_B_odZ837622_1),.clk(gclk));
	jdff dff_B_vzXoSk9X4_1(.din(w_dff_B_odZ837622_1),.dout(w_dff_B_vzXoSk9X4_1),.clk(gclk));
	jdff dff_B_adsMT2n22_1(.din(n264),.dout(w_dff_B_adsMT2n22_1),.clk(gclk));
	jdff dff_A_k4xenT4h7_0(.dout(w_n212_0[0]),.din(w_dff_A_k4xenT4h7_0),.clk(gclk));
	jdff dff_A_a7we9Gva3_0(.dout(w_dff_A_k4xenT4h7_0),.din(w_dff_A_a7we9Gva3_0),.clk(gclk));
	jdff dff_A_I0ImGIF14_0(.dout(w_dff_A_a7we9Gva3_0),.din(w_dff_A_I0ImGIF14_0),.clk(gclk));
	jdff dff_A_13YisptX2_0(.dout(w_dff_A_I0ImGIF14_0),.din(w_dff_A_13YisptX2_0),.clk(gclk));
	jdff dff_A_I9Lt9Vzd6_0(.dout(w_dff_A_13YisptX2_0),.din(w_dff_A_I9Lt9Vzd6_0),.clk(gclk));
	jdff dff_A_BTmGs1Yk9_0(.dout(w_dff_A_I9Lt9Vzd6_0),.din(w_dff_A_BTmGs1Yk9_0),.clk(gclk));
	jdff dff_A_tPINrfYB9_0(.dout(w_dff_A_BTmGs1Yk9_0),.din(w_dff_A_tPINrfYB9_0),.clk(gclk));
	jdff dff_A_BPjLgJLX3_0(.dout(w_dff_A_tPINrfYB9_0),.din(w_dff_A_BPjLgJLX3_0),.clk(gclk));
	jdff dff_A_ucfuI76z7_0(.dout(w_dff_A_BPjLgJLX3_0),.din(w_dff_A_ucfuI76z7_0),.clk(gclk));
	jdff dff_A_dkBXmf8y8_0(.dout(w_dff_A_ucfuI76z7_0),.din(w_dff_A_dkBXmf8y8_0),.clk(gclk));
	jdff dff_A_5HtJrMS99_0(.dout(w_dff_A_dkBXmf8y8_0),.din(w_dff_A_5HtJrMS99_0),.clk(gclk));
	jdff dff_A_5zkDC9HT5_0(.dout(w_dff_A_5HtJrMS99_0),.din(w_dff_A_5zkDC9HT5_0),.clk(gclk));
	jdff dff_A_YOSbSJAe4_0(.dout(w_dff_A_5zkDC9HT5_0),.din(w_dff_A_YOSbSJAe4_0),.clk(gclk));
	jdff dff_A_Aw2O2uyB6_0(.dout(w_dff_A_YOSbSJAe4_0),.din(w_dff_A_Aw2O2uyB6_0),.clk(gclk));
	jdff dff_A_2eztFaSA8_0(.dout(w_dff_A_Aw2O2uyB6_0),.din(w_dff_A_2eztFaSA8_0),.clk(gclk));
	jdff dff_A_6D4g2EIK1_0(.dout(w_dff_A_2eztFaSA8_0),.din(w_dff_A_6D4g2EIK1_0),.clk(gclk));
	jdff dff_A_wbKw1Hd12_0(.dout(w_dff_A_6D4g2EIK1_0),.din(w_dff_A_wbKw1Hd12_0),.clk(gclk));
	jdff dff_A_Z720XUCY7_0(.dout(w_dff_A_wbKw1Hd12_0),.din(w_dff_A_Z720XUCY7_0),.clk(gclk));
	jdff dff_A_mzsbKJ0A0_0(.dout(w_dff_A_Z720XUCY7_0),.din(w_dff_A_mzsbKJ0A0_0),.clk(gclk));
	jdff dff_A_mMzflZNv3_1(.dout(w_n258_0[1]),.din(w_dff_A_mMzflZNv3_1),.clk(gclk));
	jdff dff_B_AdKknkAd7_1(.din(n219),.dout(w_dff_B_AdKknkAd7_1),.clk(gclk));
	jdff dff_B_Ym6Vbl3d6_1(.din(w_dff_B_AdKknkAd7_1),.dout(w_dff_B_Ym6Vbl3d6_1),.clk(gclk));
	jdff dff_B_ATfipyHE7_1(.din(w_dff_B_Ym6Vbl3d6_1),.dout(w_dff_B_ATfipyHE7_1),.clk(gclk));
	jdff dff_B_psPElH7X9_1(.din(w_dff_B_ATfipyHE7_1),.dout(w_dff_B_psPElH7X9_1),.clk(gclk));
	jdff dff_B_o9LOOIpQ2_1(.din(w_dff_B_psPElH7X9_1),.dout(w_dff_B_o9LOOIpQ2_1),.clk(gclk));
	jdff dff_B_57Rkjt1g2_1(.din(w_dff_B_o9LOOIpQ2_1),.dout(w_dff_B_57Rkjt1g2_1),.clk(gclk));
	jdff dff_B_oYqScWT52_1(.din(w_dff_B_57Rkjt1g2_1),.dout(w_dff_B_oYqScWT52_1),.clk(gclk));
	jdff dff_B_lV0f9tA09_1(.din(w_dff_B_oYqScWT52_1),.dout(w_dff_B_lV0f9tA09_1),.clk(gclk));
	jdff dff_B_hVxklnD74_1(.din(w_dff_B_lV0f9tA09_1),.dout(w_dff_B_hVxklnD74_1),.clk(gclk));
	jdff dff_B_5jGr5oyl7_1(.din(w_dff_B_hVxklnD74_1),.dout(w_dff_B_5jGr5oyl7_1),.clk(gclk));
	jdff dff_B_Dcg3VGSg8_1(.din(w_dff_B_5jGr5oyl7_1),.dout(w_dff_B_Dcg3VGSg8_1),.clk(gclk));
	jdff dff_B_ptQJVMAC3_1(.din(w_dff_B_Dcg3VGSg8_1),.dout(w_dff_B_ptQJVMAC3_1),.clk(gclk));
	jdff dff_B_b6MtkQpX9_1(.din(w_dff_B_ptQJVMAC3_1),.dout(w_dff_B_b6MtkQpX9_1),.clk(gclk));
	jdff dff_B_rKwLbcEY2_1(.din(w_dff_B_b6MtkQpX9_1),.dout(w_dff_B_rKwLbcEY2_1),.clk(gclk));
	jdff dff_B_aBcORKe87_1(.din(w_dff_B_rKwLbcEY2_1),.dout(w_dff_B_aBcORKe87_1),.clk(gclk));
	jdff dff_B_e2lxoe595_1(.din(n215),.dout(w_dff_B_e2lxoe595_1),.clk(gclk));
	jdff dff_A_0pDleJ5R5_0(.dout(w_n170_0[0]),.din(w_dff_A_0pDleJ5R5_0),.clk(gclk));
	jdff dff_A_mHUCRWvC3_0(.dout(w_dff_A_0pDleJ5R5_0),.din(w_dff_A_mHUCRWvC3_0),.clk(gclk));
	jdff dff_A_KvTRu6M32_0(.dout(w_dff_A_mHUCRWvC3_0),.din(w_dff_A_KvTRu6M32_0),.clk(gclk));
	jdff dff_A_NMlXlc5E6_0(.dout(w_dff_A_KvTRu6M32_0),.din(w_dff_A_NMlXlc5E6_0),.clk(gclk));
	jdff dff_A_6Vq3yUtu1_0(.dout(w_dff_A_NMlXlc5E6_0),.din(w_dff_A_6Vq3yUtu1_0),.clk(gclk));
	jdff dff_A_EnQjXoip4_0(.dout(w_dff_A_6Vq3yUtu1_0),.din(w_dff_A_EnQjXoip4_0),.clk(gclk));
	jdff dff_A_Lr4elQOt6_0(.dout(w_dff_A_EnQjXoip4_0),.din(w_dff_A_Lr4elQOt6_0),.clk(gclk));
	jdff dff_A_8UBRyQ647_0(.dout(w_dff_A_Lr4elQOt6_0),.din(w_dff_A_8UBRyQ647_0),.clk(gclk));
	jdff dff_A_JYv7GULW8_0(.dout(w_dff_A_8UBRyQ647_0),.din(w_dff_A_JYv7GULW8_0),.clk(gclk));
	jdff dff_A_GscKWzc12_0(.dout(w_dff_A_JYv7GULW8_0),.din(w_dff_A_GscKWzc12_0),.clk(gclk));
	jdff dff_A_guE4PUy30_0(.dout(w_dff_A_GscKWzc12_0),.din(w_dff_A_guE4PUy30_0),.clk(gclk));
	jdff dff_A_Ju6eZYVy8_0(.dout(w_dff_A_guE4PUy30_0),.din(w_dff_A_Ju6eZYVy8_0),.clk(gclk));
	jdff dff_A_R1jzM2gi9_0(.dout(w_dff_A_Ju6eZYVy8_0),.din(w_dff_A_R1jzM2gi9_0),.clk(gclk));
	jdff dff_A_MElvZuSi2_0(.dout(w_dff_A_R1jzM2gi9_0),.din(w_dff_A_MElvZuSi2_0),.clk(gclk));
	jdff dff_A_8MtG78A65_0(.dout(w_dff_A_MElvZuSi2_0),.din(w_dff_A_8MtG78A65_0),.clk(gclk));
	jdff dff_A_O45etuQo1_0(.dout(w_dff_A_8MtG78A65_0),.din(w_dff_A_O45etuQo1_0),.clk(gclk));
	jdff dff_A_w1J36y282_1(.dout(w_n209_0[1]),.din(w_dff_A_w1J36y282_1),.clk(gclk));
	jdff dff_B_kMJdIi8X0_1(.din(n177),.dout(w_dff_B_kMJdIi8X0_1),.clk(gclk));
	jdff dff_B_acniKS1l7_1(.din(w_dff_B_kMJdIi8X0_1),.dout(w_dff_B_acniKS1l7_1),.clk(gclk));
	jdff dff_B_sKMPpX0Y6_1(.din(w_dff_B_acniKS1l7_1),.dout(w_dff_B_sKMPpX0Y6_1),.clk(gclk));
	jdff dff_B_lkREedsx8_1(.din(w_dff_B_sKMPpX0Y6_1),.dout(w_dff_B_lkREedsx8_1),.clk(gclk));
	jdff dff_B_LuK1vCnM8_1(.din(w_dff_B_lkREedsx8_1),.dout(w_dff_B_LuK1vCnM8_1),.clk(gclk));
	jdff dff_B_7iCANmHr3_1(.din(w_dff_B_LuK1vCnM8_1),.dout(w_dff_B_7iCANmHr3_1),.clk(gclk));
	jdff dff_B_5R1v7BSg4_1(.din(w_dff_B_7iCANmHr3_1),.dout(w_dff_B_5R1v7BSg4_1),.clk(gclk));
	jdff dff_B_lIklxeFu5_1(.din(w_dff_B_5R1v7BSg4_1),.dout(w_dff_B_lIklxeFu5_1),.clk(gclk));
	jdff dff_B_EMIjIBl47_1(.din(w_dff_B_lIklxeFu5_1),.dout(w_dff_B_EMIjIBl47_1),.clk(gclk));
	jdff dff_B_pRj0KyJu7_1(.din(w_dff_B_EMIjIBl47_1),.dout(w_dff_B_pRj0KyJu7_1),.clk(gclk));
	jdff dff_B_Zyuwm4wT3_1(.din(w_dff_B_pRj0KyJu7_1),.dout(w_dff_B_Zyuwm4wT3_1),.clk(gclk));
	jdff dff_B_223yyBnc1_1(.din(w_dff_B_Zyuwm4wT3_1),.dout(w_dff_B_223yyBnc1_1),.clk(gclk));
	jdff dff_B_mivY9yYO3_1(.din(n173),.dout(w_dff_B_mivY9yYO3_1),.clk(gclk));
	jdff dff_A_YghuRqzn2_0(.dout(w_n135_0[0]),.din(w_dff_A_YghuRqzn2_0),.clk(gclk));
	jdff dff_A_mCe75unF2_0(.dout(w_dff_A_YghuRqzn2_0),.din(w_dff_A_mCe75unF2_0),.clk(gclk));
	jdff dff_A_LLBwnret3_0(.dout(w_dff_A_mCe75unF2_0),.din(w_dff_A_LLBwnret3_0),.clk(gclk));
	jdff dff_A_A2uk5kT93_0(.dout(w_dff_A_LLBwnret3_0),.din(w_dff_A_A2uk5kT93_0),.clk(gclk));
	jdff dff_A_GRq9yJjw4_0(.dout(w_dff_A_A2uk5kT93_0),.din(w_dff_A_GRq9yJjw4_0),.clk(gclk));
	jdff dff_A_IbVR6JTN4_0(.dout(w_dff_A_GRq9yJjw4_0),.din(w_dff_A_IbVR6JTN4_0),.clk(gclk));
	jdff dff_A_Kcu7LNBs7_0(.dout(w_dff_A_IbVR6JTN4_0),.din(w_dff_A_Kcu7LNBs7_0),.clk(gclk));
	jdff dff_A_rGT5YZ3j4_0(.dout(w_dff_A_Kcu7LNBs7_0),.din(w_dff_A_rGT5YZ3j4_0),.clk(gclk));
	jdff dff_A_ApxXQGR94_0(.dout(w_dff_A_rGT5YZ3j4_0),.din(w_dff_A_ApxXQGR94_0),.clk(gclk));
	jdff dff_A_V76GR7Iw8_0(.dout(w_dff_A_ApxXQGR94_0),.din(w_dff_A_V76GR7Iw8_0),.clk(gclk));
	jdff dff_A_2TC2PRkm0_0(.dout(w_dff_A_V76GR7Iw8_0),.din(w_dff_A_2TC2PRkm0_0),.clk(gclk));
	jdff dff_A_ItZ3DfJD9_0(.dout(w_dff_A_2TC2PRkm0_0),.din(w_dff_A_ItZ3DfJD9_0),.clk(gclk));
	jdff dff_A_vEHJDhK88_0(.dout(w_dff_A_ItZ3DfJD9_0),.din(w_dff_A_vEHJDhK88_0),.clk(gclk));
	jdff dff_A_RjMD47tF9_1(.dout(w_n167_0[1]),.din(w_dff_A_RjMD47tF9_1),.clk(gclk));
	jdff dff_B_uW5YyeLi5_1(.din(n142),.dout(w_dff_B_uW5YyeLi5_1),.clk(gclk));
	jdff dff_B_F8HT6iDB7_1(.din(w_dff_B_uW5YyeLi5_1),.dout(w_dff_B_F8HT6iDB7_1),.clk(gclk));
	jdff dff_B_spgkFarl1_1(.din(w_dff_B_F8HT6iDB7_1),.dout(w_dff_B_spgkFarl1_1),.clk(gclk));
	jdff dff_B_Cl3PKAn14_1(.din(w_dff_B_spgkFarl1_1),.dout(w_dff_B_Cl3PKAn14_1),.clk(gclk));
	jdff dff_B_H0hHKyTQ3_1(.din(w_dff_B_Cl3PKAn14_1),.dout(w_dff_B_H0hHKyTQ3_1),.clk(gclk));
	jdff dff_B_3NaMh7mf2_1(.din(w_dff_B_H0hHKyTQ3_1),.dout(w_dff_B_3NaMh7mf2_1),.clk(gclk));
	jdff dff_B_8u50gTNV8_1(.din(w_dff_B_3NaMh7mf2_1),.dout(w_dff_B_8u50gTNV8_1),.clk(gclk));
	jdff dff_B_U8ykEoTV5_1(.din(w_dff_B_8u50gTNV8_1),.dout(w_dff_B_U8ykEoTV5_1),.clk(gclk));
	jdff dff_B_kHBgj2ct0_1(.din(w_dff_B_U8ykEoTV5_1),.dout(w_dff_B_kHBgj2ct0_1),.clk(gclk));
	jdff dff_B_gf04LRoR5_1(.din(n138),.dout(w_dff_B_gf04LRoR5_1),.clk(gclk));
	jdff dff_A_KFtXeObF6_0(.dout(w_n106_0[0]),.din(w_dff_A_KFtXeObF6_0),.clk(gclk));
	jdff dff_A_gDAG2uvu0_0(.dout(w_dff_A_KFtXeObF6_0),.din(w_dff_A_gDAG2uvu0_0),.clk(gclk));
	jdff dff_A_l3fN9AQo9_0(.dout(w_dff_A_gDAG2uvu0_0),.din(w_dff_A_l3fN9AQo9_0),.clk(gclk));
	jdff dff_A_zmhu8g9k0_0(.dout(w_dff_A_l3fN9AQo9_0),.din(w_dff_A_zmhu8g9k0_0),.clk(gclk));
	jdff dff_A_DlyKsRMP4_0(.dout(w_dff_A_zmhu8g9k0_0),.din(w_dff_A_DlyKsRMP4_0),.clk(gclk));
	jdff dff_A_4nmWnb527_0(.dout(w_dff_A_DlyKsRMP4_0),.din(w_dff_A_4nmWnb527_0),.clk(gclk));
	jdff dff_A_valVlmqL2_0(.dout(w_dff_A_4nmWnb527_0),.din(w_dff_A_valVlmqL2_0),.clk(gclk));
	jdff dff_A_gF5BJC1H4_0(.dout(w_dff_A_valVlmqL2_0),.din(w_dff_A_gF5BJC1H4_0),.clk(gclk));
	jdff dff_A_CxuUWjyH7_0(.dout(w_dff_A_gF5BJC1H4_0),.din(w_dff_A_CxuUWjyH7_0),.clk(gclk));
	jdff dff_A_mRes1rl40_0(.dout(w_dff_A_CxuUWjyH7_0),.din(w_dff_A_mRes1rl40_0),.clk(gclk));
	jdff dff_A_WxYnSB6O0_1(.dout(w_n132_0[1]),.din(w_dff_A_WxYnSB6O0_1),.clk(gclk));
	jdff dff_B_IuinFrhh4_1(.din(n113),.dout(w_dff_B_IuinFrhh4_1),.clk(gclk));
	jdff dff_B_BQSZpY1a8_1(.din(w_dff_B_IuinFrhh4_1),.dout(w_dff_B_BQSZpY1a8_1),.clk(gclk));
	jdff dff_B_PdmuyN320_1(.din(w_dff_B_BQSZpY1a8_1),.dout(w_dff_B_PdmuyN320_1),.clk(gclk));
	jdff dff_B_W36D3cMK6_1(.din(w_dff_B_PdmuyN320_1),.dout(w_dff_B_W36D3cMK6_1),.clk(gclk));
	jdff dff_B_NGmeOSA00_1(.din(w_dff_B_W36D3cMK6_1),.dout(w_dff_B_NGmeOSA00_1),.clk(gclk));
	jdff dff_B_Su360Bny1_1(.din(w_dff_B_NGmeOSA00_1),.dout(w_dff_B_Su360Bny1_1),.clk(gclk));
	jdff dff_B_wzAgij7Z4_1(.din(n109),.dout(w_dff_B_wzAgij7Z4_1),.clk(gclk));
	jdff dff_A_9U95j5xh3_0(.dout(w_n86_0[0]),.din(w_dff_A_9U95j5xh3_0),.clk(gclk));
	jdff dff_A_ZP3HyAxE7_0(.dout(w_dff_A_9U95j5xh3_0),.din(w_dff_A_ZP3HyAxE7_0),.clk(gclk));
	jdff dff_A_uiWKBazU3_0(.dout(w_dff_A_ZP3HyAxE7_0),.din(w_dff_A_uiWKBazU3_0),.clk(gclk));
	jdff dff_A_kFeW8RfP9_0(.dout(w_dff_A_uiWKBazU3_0),.din(w_dff_A_kFeW8RfP9_0),.clk(gclk));
	jdff dff_A_KoVx2Kan5_0(.dout(w_dff_A_kFeW8RfP9_0),.din(w_dff_A_KoVx2Kan5_0),.clk(gclk));
	jdff dff_A_Ylz2tDqD9_0(.dout(w_dff_A_KoVx2Kan5_0),.din(w_dff_A_Ylz2tDqD9_0),.clk(gclk));
	jdff dff_A_GHg8aXye0_0(.dout(w_dff_A_Ylz2tDqD9_0),.din(w_dff_A_GHg8aXye0_0),.clk(gclk));
	jdff dff_A_GQBtAAG96_1(.dout(w_n103_0[1]),.din(w_dff_A_GQBtAAG96_1),.clk(gclk));
	jdff dff_B_Uv9ReWOd9_1(.din(n92),.dout(w_dff_B_Uv9ReWOd9_1),.clk(gclk));
	jdff dff_B_NMrMQwpv2_1(.din(w_dff_B_Uv9ReWOd9_1),.dout(w_dff_B_NMrMQwpv2_1),.clk(gclk));
	jdff dff_B_cXBzVoJC3_1(.din(w_dff_B_NMrMQwpv2_1),.dout(w_dff_B_cXBzVoJC3_1),.clk(gclk));
	jdff dff_B_bRNIW5P95_1(.din(n88),.dout(w_dff_B_bRNIW5P95_1),.clk(gclk));
	jdff dff_B_9Vf5Icva4_2(.din(n67),.dout(w_dff_B_9Vf5Icva4_2),.clk(gclk));
	jdff dff_A_CH6f1AEo0_0(.dout(w_n75_0[0]),.din(w_dff_A_CH6f1AEo0_0),.clk(gclk));
	jdff dff_A_BfS0jTiv1_0(.dout(w_dff_A_CH6f1AEo0_0),.din(w_dff_A_BfS0jTiv1_0),.clk(gclk));
	jdff dff_A_HwO8AQJo2_0(.dout(w_dff_A_BfS0jTiv1_0),.din(w_dff_A_HwO8AQJo2_0),.clk(gclk));
	jdff dff_A_eQtCUR2S4_0(.dout(w_dff_A_HwO8AQJo2_0),.din(w_dff_A_eQtCUR2S4_0),.clk(gclk));
	jdff dff_B_QKLZD07U2_0(.din(n82),.dout(w_dff_B_QKLZD07U2_0),.clk(gclk));
	jdff dff_A_HWHyE6Iw3_0(.dout(w_n66_0[0]),.din(w_dff_A_HWHyE6Iw3_0),.clk(gclk));
	jdff dff_A_eAFIM9nI2_0(.dout(w_dff_A_HWHyE6Iw3_0),.din(w_dff_A_eAFIM9nI2_0),.clk(gclk));
	jdff dff_A_ezmFXke16_1(.dout(w_n1108_0[1]),.din(w_dff_A_ezmFXke16_1),.clk(gclk));
	jdff dff_B_ha1f2K3W5_1(.din(n1014),.dout(w_dff_B_ha1f2K3W5_1),.clk(gclk));
	jdff dff_B_SVlH4JPV1_2(.din(n911),.dout(w_dff_B_SVlH4JPV1_2),.clk(gclk));
	jdff dff_B_1dCmcIVs7_2(.din(w_dff_B_SVlH4JPV1_2),.dout(w_dff_B_1dCmcIVs7_2),.clk(gclk));
	jdff dff_B_HXwN8Lw13_2(.din(w_dff_B_1dCmcIVs7_2),.dout(w_dff_B_HXwN8Lw13_2),.clk(gclk));
	jdff dff_B_z04SlnyX3_2(.din(w_dff_B_HXwN8Lw13_2),.dout(w_dff_B_z04SlnyX3_2),.clk(gclk));
	jdff dff_B_Yq8ukHI04_2(.din(w_dff_B_z04SlnyX3_2),.dout(w_dff_B_Yq8ukHI04_2),.clk(gclk));
	jdff dff_B_NmQc9hKf4_2(.din(w_dff_B_Yq8ukHI04_2),.dout(w_dff_B_NmQc9hKf4_2),.clk(gclk));
	jdff dff_B_XuNwJZp97_2(.din(w_dff_B_NmQc9hKf4_2),.dout(w_dff_B_XuNwJZp97_2),.clk(gclk));
	jdff dff_B_fKhPNZ3o0_2(.din(w_dff_B_XuNwJZp97_2),.dout(w_dff_B_fKhPNZ3o0_2),.clk(gclk));
	jdff dff_B_13MhYITO2_2(.din(w_dff_B_fKhPNZ3o0_2),.dout(w_dff_B_13MhYITO2_2),.clk(gclk));
	jdff dff_B_XFPRGYNU8_2(.din(w_dff_B_13MhYITO2_2),.dout(w_dff_B_XFPRGYNU8_2),.clk(gclk));
	jdff dff_B_buTV6WBg6_2(.din(w_dff_B_XFPRGYNU8_2),.dout(w_dff_B_buTV6WBg6_2),.clk(gclk));
	jdff dff_B_UjuXZ5CJ3_2(.din(w_dff_B_buTV6WBg6_2),.dout(w_dff_B_UjuXZ5CJ3_2),.clk(gclk));
	jdff dff_B_05ly3pzf6_2(.din(w_dff_B_UjuXZ5CJ3_2),.dout(w_dff_B_05ly3pzf6_2),.clk(gclk));
	jdff dff_B_1BVgJJ1u8_2(.din(w_dff_B_05ly3pzf6_2),.dout(w_dff_B_1BVgJJ1u8_2),.clk(gclk));
	jdff dff_B_XLESq5Yo7_2(.din(w_dff_B_1BVgJJ1u8_2),.dout(w_dff_B_XLESq5Yo7_2),.clk(gclk));
	jdff dff_B_bvomDQYL5_2(.din(w_dff_B_XLESq5Yo7_2),.dout(w_dff_B_bvomDQYL5_2),.clk(gclk));
	jdff dff_B_q9w15ckF9_2(.din(w_dff_B_bvomDQYL5_2),.dout(w_dff_B_q9w15ckF9_2),.clk(gclk));
	jdff dff_B_hD4v8Ou89_2(.din(w_dff_B_q9w15ckF9_2),.dout(w_dff_B_hD4v8Ou89_2),.clk(gclk));
	jdff dff_B_X7ecC6Wd5_2(.din(w_dff_B_hD4v8Ou89_2),.dout(w_dff_B_X7ecC6Wd5_2),.clk(gclk));
	jdff dff_B_QafV0eiG5_2(.din(w_dff_B_X7ecC6Wd5_2),.dout(w_dff_B_QafV0eiG5_2),.clk(gclk));
	jdff dff_B_RrjQB6hy1_2(.din(w_dff_B_QafV0eiG5_2),.dout(w_dff_B_RrjQB6hy1_2),.clk(gclk));
	jdff dff_B_NGJoTSCz3_2(.din(w_dff_B_RrjQB6hy1_2),.dout(w_dff_B_NGJoTSCz3_2),.clk(gclk));
	jdff dff_B_ayq64um91_2(.din(w_dff_B_NGJoTSCz3_2),.dout(w_dff_B_ayq64um91_2),.clk(gclk));
	jdff dff_B_19hUALFP2_2(.din(w_dff_B_ayq64um91_2),.dout(w_dff_B_19hUALFP2_2),.clk(gclk));
	jdff dff_B_MGeJWS6N6_2(.din(w_dff_B_19hUALFP2_2),.dout(w_dff_B_MGeJWS6N6_2),.clk(gclk));
	jdff dff_B_S4elgKpK0_2(.din(w_dff_B_MGeJWS6N6_2),.dout(w_dff_B_S4elgKpK0_2),.clk(gclk));
	jdff dff_B_NUkd8ZMM3_2(.din(w_dff_B_S4elgKpK0_2),.dout(w_dff_B_NUkd8ZMM3_2),.clk(gclk));
	jdff dff_B_Pdm31MgI0_2(.din(w_dff_B_NUkd8ZMM3_2),.dout(w_dff_B_Pdm31MgI0_2),.clk(gclk));
	jdff dff_B_ST9919Fo5_2(.din(w_dff_B_Pdm31MgI0_2),.dout(w_dff_B_ST9919Fo5_2),.clk(gclk));
	jdff dff_B_rykJtCo34_2(.din(w_dff_B_ST9919Fo5_2),.dout(w_dff_B_rykJtCo34_2),.clk(gclk));
	jdff dff_B_v9OHv9Jy7_2(.din(w_dff_B_rykJtCo34_2),.dout(w_dff_B_v9OHv9Jy7_2),.clk(gclk));
	jdff dff_B_9UDA5jTH7_2(.din(w_dff_B_v9OHv9Jy7_2),.dout(w_dff_B_9UDA5jTH7_2),.clk(gclk));
	jdff dff_B_o96nVqcz0_2(.din(w_dff_B_9UDA5jTH7_2),.dout(w_dff_B_o96nVqcz0_2),.clk(gclk));
	jdff dff_B_dsntBdmM9_2(.din(w_dff_B_o96nVqcz0_2),.dout(w_dff_B_dsntBdmM9_2),.clk(gclk));
	jdff dff_B_PGcsK3oM3_2(.din(w_dff_B_dsntBdmM9_2),.dout(w_dff_B_PGcsK3oM3_2),.clk(gclk));
	jdff dff_B_DW5CnjLJ6_2(.din(w_dff_B_PGcsK3oM3_2),.dout(w_dff_B_DW5CnjLJ6_2),.clk(gclk));
	jdff dff_B_kPbPoVDA1_2(.din(w_dff_B_DW5CnjLJ6_2),.dout(w_dff_B_kPbPoVDA1_2),.clk(gclk));
	jdff dff_B_U2tUafzD3_2(.din(w_dff_B_kPbPoVDA1_2),.dout(w_dff_B_U2tUafzD3_2),.clk(gclk));
	jdff dff_B_eWjOhlCz6_2(.din(w_dff_B_U2tUafzD3_2),.dout(w_dff_B_eWjOhlCz6_2),.clk(gclk));
	jdff dff_B_n3CbNZ7m1_2(.din(w_dff_B_eWjOhlCz6_2),.dout(w_dff_B_n3CbNZ7m1_2),.clk(gclk));
	jdff dff_B_h19lBGnf6_2(.din(w_dff_B_n3CbNZ7m1_2),.dout(w_dff_B_h19lBGnf6_2),.clk(gclk));
	jdff dff_B_YmRQM7ho6_2(.din(w_dff_B_h19lBGnf6_2),.dout(w_dff_B_YmRQM7ho6_2),.clk(gclk));
	jdff dff_B_5PjTactY9_2(.din(w_dff_B_YmRQM7ho6_2),.dout(w_dff_B_5PjTactY9_2),.clk(gclk));
	jdff dff_A_2JoOJDSK2_0(.dout(w_n1008_0[0]),.din(w_dff_A_2JoOJDSK2_0),.clk(gclk));
	jdff dff_B_dHhXXkpS5_1(.din(n913),.dout(w_dff_B_dHhXXkpS5_1),.clk(gclk));
	jdff dff_B_J4iVVmD45_2(.din(n811),.dout(w_dff_B_J4iVVmD45_2),.clk(gclk));
	jdff dff_B_kRUpxviw3_2(.din(w_dff_B_J4iVVmD45_2),.dout(w_dff_B_kRUpxviw3_2),.clk(gclk));
	jdff dff_B_00tmrzpk5_2(.din(w_dff_B_kRUpxviw3_2),.dout(w_dff_B_00tmrzpk5_2),.clk(gclk));
	jdff dff_B_sX4AHlqn2_2(.din(w_dff_B_00tmrzpk5_2),.dout(w_dff_B_sX4AHlqn2_2),.clk(gclk));
	jdff dff_B_XiFH1nWY4_2(.din(w_dff_B_sX4AHlqn2_2),.dout(w_dff_B_XiFH1nWY4_2),.clk(gclk));
	jdff dff_B_JjgOmFdZ7_2(.din(w_dff_B_XiFH1nWY4_2),.dout(w_dff_B_JjgOmFdZ7_2),.clk(gclk));
	jdff dff_B_xCXM2NdE3_2(.din(w_dff_B_JjgOmFdZ7_2),.dout(w_dff_B_xCXM2NdE3_2),.clk(gclk));
	jdff dff_B_tXtJZLsf3_2(.din(w_dff_B_xCXM2NdE3_2),.dout(w_dff_B_tXtJZLsf3_2),.clk(gclk));
	jdff dff_B_C68lsUKi6_2(.din(w_dff_B_tXtJZLsf3_2),.dout(w_dff_B_C68lsUKi6_2),.clk(gclk));
	jdff dff_B_o8ytgLja9_2(.din(w_dff_B_C68lsUKi6_2),.dout(w_dff_B_o8ytgLja9_2),.clk(gclk));
	jdff dff_B_5maTWP3Q7_2(.din(w_dff_B_o8ytgLja9_2),.dout(w_dff_B_5maTWP3Q7_2),.clk(gclk));
	jdff dff_B_EOLkSml62_2(.din(w_dff_B_5maTWP3Q7_2),.dout(w_dff_B_EOLkSml62_2),.clk(gclk));
	jdff dff_B_5J2p2Z6a5_2(.din(w_dff_B_EOLkSml62_2),.dout(w_dff_B_5J2p2Z6a5_2),.clk(gclk));
	jdff dff_B_wiSXpisI5_2(.din(w_dff_B_5J2p2Z6a5_2),.dout(w_dff_B_wiSXpisI5_2),.clk(gclk));
	jdff dff_B_T20hXRdQ5_2(.din(w_dff_B_wiSXpisI5_2),.dout(w_dff_B_T20hXRdQ5_2),.clk(gclk));
	jdff dff_B_hyFsdzvO5_2(.din(w_dff_B_T20hXRdQ5_2),.dout(w_dff_B_hyFsdzvO5_2),.clk(gclk));
	jdff dff_B_ZHpLUpvA3_2(.din(w_dff_B_hyFsdzvO5_2),.dout(w_dff_B_ZHpLUpvA3_2),.clk(gclk));
	jdff dff_B_C6MODavM5_2(.din(w_dff_B_ZHpLUpvA3_2),.dout(w_dff_B_C6MODavM5_2),.clk(gclk));
	jdff dff_B_Q4GKMZ6Q8_2(.din(w_dff_B_C6MODavM5_2),.dout(w_dff_B_Q4GKMZ6Q8_2),.clk(gclk));
	jdff dff_B_yBBfHVMM8_2(.din(w_dff_B_Q4GKMZ6Q8_2),.dout(w_dff_B_yBBfHVMM8_2),.clk(gclk));
	jdff dff_B_6rFDfqKX0_2(.din(w_dff_B_yBBfHVMM8_2),.dout(w_dff_B_6rFDfqKX0_2),.clk(gclk));
	jdff dff_B_rYoQMKwM4_2(.din(w_dff_B_6rFDfqKX0_2),.dout(w_dff_B_rYoQMKwM4_2),.clk(gclk));
	jdff dff_B_mC83W5Rc5_2(.din(w_dff_B_rYoQMKwM4_2),.dout(w_dff_B_mC83W5Rc5_2),.clk(gclk));
	jdff dff_B_uJtnMJem2_2(.din(w_dff_B_mC83W5Rc5_2),.dout(w_dff_B_uJtnMJem2_2),.clk(gclk));
	jdff dff_B_QKsNVTjd3_2(.din(w_dff_B_uJtnMJem2_2),.dout(w_dff_B_QKsNVTjd3_2),.clk(gclk));
	jdff dff_B_oqvn98nS2_2(.din(w_dff_B_QKsNVTjd3_2),.dout(w_dff_B_oqvn98nS2_2),.clk(gclk));
	jdff dff_B_7BcMa4337_2(.din(w_dff_B_oqvn98nS2_2),.dout(w_dff_B_7BcMa4337_2),.clk(gclk));
	jdff dff_B_8hs0nVhs3_2(.din(w_dff_B_7BcMa4337_2),.dout(w_dff_B_8hs0nVhs3_2),.clk(gclk));
	jdff dff_B_Vc8OozMm0_2(.din(w_dff_B_8hs0nVhs3_2),.dout(w_dff_B_Vc8OozMm0_2),.clk(gclk));
	jdff dff_B_PYBsMJ9P9_2(.din(w_dff_B_Vc8OozMm0_2),.dout(w_dff_B_PYBsMJ9P9_2),.clk(gclk));
	jdff dff_B_xMXPbBb82_2(.din(w_dff_B_PYBsMJ9P9_2),.dout(w_dff_B_xMXPbBb82_2),.clk(gclk));
	jdff dff_B_p2nWBI8F7_2(.din(w_dff_B_xMXPbBb82_2),.dout(w_dff_B_p2nWBI8F7_2),.clk(gclk));
	jdff dff_B_ddwJvNLP0_2(.din(w_dff_B_p2nWBI8F7_2),.dout(w_dff_B_ddwJvNLP0_2),.clk(gclk));
	jdff dff_B_KjfHu9ii9_2(.din(w_dff_B_ddwJvNLP0_2),.dout(w_dff_B_KjfHu9ii9_2),.clk(gclk));
	jdff dff_B_0AxgoCU34_2(.din(w_dff_B_KjfHu9ii9_2),.dout(w_dff_B_0AxgoCU34_2),.clk(gclk));
	jdff dff_B_FGlZw0UB6_2(.din(w_dff_B_0AxgoCU34_2),.dout(w_dff_B_FGlZw0UB6_2),.clk(gclk));
	jdff dff_B_apCgWL839_2(.din(w_dff_B_FGlZw0UB6_2),.dout(w_dff_B_apCgWL839_2),.clk(gclk));
	jdff dff_B_AgWRX1l88_2(.din(w_dff_B_apCgWL839_2),.dout(w_dff_B_AgWRX1l88_2),.clk(gclk));
	jdff dff_B_WQwPjHer9_2(.din(w_dff_B_AgWRX1l88_2),.dout(w_dff_B_WQwPjHer9_2),.clk(gclk));
	jdff dff_B_hfAiVJWe3_2(.din(w_dff_B_WQwPjHer9_2),.dout(w_dff_B_hfAiVJWe3_2),.clk(gclk));
	jdff dff_A_5cOfMQR71_1(.dout(w_n902_0[1]),.din(w_dff_A_5cOfMQR71_1),.clk(gclk));
	jdff dff_B_RNAk0Tkx4_1(.din(n817),.dout(w_dff_B_RNAk0Tkx4_1),.clk(gclk));
	jdff dff_B_PhiVPLAi5_1(.din(w_dff_B_RNAk0Tkx4_1),.dout(w_dff_B_PhiVPLAi5_1),.clk(gclk));
	jdff dff_B_InFZxYzN7_1(.din(w_dff_B_PhiVPLAi5_1),.dout(w_dff_B_InFZxYzN7_1),.clk(gclk));
	jdff dff_B_oBaMsv0G5_1(.din(w_dff_B_InFZxYzN7_1),.dout(w_dff_B_oBaMsv0G5_1),.clk(gclk));
	jdff dff_B_jMryvljm0_1(.din(w_dff_B_oBaMsv0G5_1),.dout(w_dff_B_jMryvljm0_1),.clk(gclk));
	jdff dff_B_jMceVpjg0_1(.din(w_dff_B_jMryvljm0_1),.dout(w_dff_B_jMceVpjg0_1),.clk(gclk));
	jdff dff_B_heRGCE8B9_1(.din(w_dff_B_jMceVpjg0_1),.dout(w_dff_B_heRGCE8B9_1),.clk(gclk));
	jdff dff_B_GaBfpLVx4_1(.din(w_dff_B_heRGCE8B9_1),.dout(w_dff_B_GaBfpLVx4_1),.clk(gclk));
	jdff dff_B_9uO6NMfn0_1(.din(w_dff_B_GaBfpLVx4_1),.dout(w_dff_B_9uO6NMfn0_1),.clk(gclk));
	jdff dff_B_x3ieAqcX2_1(.din(w_dff_B_9uO6NMfn0_1),.dout(w_dff_B_x3ieAqcX2_1),.clk(gclk));
	jdff dff_B_7IiFwS3P8_1(.din(w_dff_B_x3ieAqcX2_1),.dout(w_dff_B_7IiFwS3P8_1),.clk(gclk));
	jdff dff_B_MMbV8bfs2_1(.din(w_dff_B_7IiFwS3P8_1),.dout(w_dff_B_MMbV8bfs2_1),.clk(gclk));
	jdff dff_B_EwlDGIH42_1(.din(w_dff_B_MMbV8bfs2_1),.dout(w_dff_B_EwlDGIH42_1),.clk(gclk));
	jdff dff_B_cdFzpImB1_1(.din(w_dff_B_EwlDGIH42_1),.dout(w_dff_B_cdFzpImB1_1),.clk(gclk));
	jdff dff_B_dl5NeYNR9_1(.din(w_dff_B_cdFzpImB1_1),.dout(w_dff_B_dl5NeYNR9_1),.clk(gclk));
	jdff dff_B_5vqpXoGX5_1(.din(w_dff_B_dl5NeYNR9_1),.dout(w_dff_B_5vqpXoGX5_1),.clk(gclk));
	jdff dff_B_ZjGfVioi1_1(.din(w_dff_B_5vqpXoGX5_1),.dout(w_dff_B_ZjGfVioi1_1),.clk(gclk));
	jdff dff_B_0q1L5jKI0_1(.din(w_dff_B_ZjGfVioi1_1),.dout(w_dff_B_0q1L5jKI0_1),.clk(gclk));
	jdff dff_B_G80Po5kR9_1(.din(w_dff_B_0q1L5jKI0_1),.dout(w_dff_B_G80Po5kR9_1),.clk(gclk));
	jdff dff_B_huyKn8U95_1(.din(w_dff_B_G80Po5kR9_1),.dout(w_dff_B_huyKn8U95_1),.clk(gclk));
	jdff dff_B_VSsqfEtz9_1(.din(w_dff_B_huyKn8U95_1),.dout(w_dff_B_VSsqfEtz9_1),.clk(gclk));
	jdff dff_B_fHp5JBK31_1(.din(w_dff_B_VSsqfEtz9_1),.dout(w_dff_B_fHp5JBK31_1),.clk(gclk));
	jdff dff_B_Y50gPpK19_1(.din(w_dff_B_fHp5JBK31_1),.dout(w_dff_B_Y50gPpK19_1),.clk(gclk));
	jdff dff_B_3ivmdiVg8_1(.din(w_dff_B_Y50gPpK19_1),.dout(w_dff_B_3ivmdiVg8_1),.clk(gclk));
	jdff dff_B_iX1uKm0m5_1(.din(w_dff_B_3ivmdiVg8_1),.dout(w_dff_B_iX1uKm0m5_1),.clk(gclk));
	jdff dff_B_SyEwpmjE0_1(.din(w_dff_B_iX1uKm0m5_1),.dout(w_dff_B_SyEwpmjE0_1),.clk(gclk));
	jdff dff_B_lZFbIdAi7_1(.din(w_dff_B_SyEwpmjE0_1),.dout(w_dff_B_lZFbIdAi7_1),.clk(gclk));
	jdff dff_B_p6NBbtwH1_1(.din(w_dff_B_lZFbIdAi7_1),.dout(w_dff_B_p6NBbtwH1_1),.clk(gclk));
	jdff dff_B_yEzUR16l3_1(.din(w_dff_B_p6NBbtwH1_1),.dout(w_dff_B_yEzUR16l3_1),.clk(gclk));
	jdff dff_B_BVIuilGA2_1(.din(w_dff_B_yEzUR16l3_1),.dout(w_dff_B_BVIuilGA2_1),.clk(gclk));
	jdff dff_B_9Dp1CswD9_1(.din(w_dff_B_BVIuilGA2_1),.dout(w_dff_B_9Dp1CswD9_1),.clk(gclk));
	jdff dff_B_0UZTnRyO1_1(.din(w_dff_B_9Dp1CswD9_1),.dout(w_dff_B_0UZTnRyO1_1),.clk(gclk));
	jdff dff_B_mGM3q0Vz8_1(.din(w_dff_B_0UZTnRyO1_1),.dout(w_dff_B_mGM3q0Vz8_1),.clk(gclk));
	jdff dff_B_KUOq6v4B6_1(.din(w_dff_B_mGM3q0Vz8_1),.dout(w_dff_B_KUOq6v4B6_1),.clk(gclk));
	jdff dff_B_Ga6U3ZaT1_1(.din(w_dff_B_KUOq6v4B6_1),.dout(w_dff_B_Ga6U3ZaT1_1),.clk(gclk));
	jdff dff_B_i87Plare9_1(.din(w_dff_B_Ga6U3ZaT1_1),.dout(w_dff_B_i87Plare9_1),.clk(gclk));
	jdff dff_B_Z8LzQloI7_1(.din(n812),.dout(w_dff_B_Z8LzQloI7_1),.clk(gclk));
	jdff dff_A_nvzMUPSq9_0(.dout(w_n712_0[0]),.din(w_dff_A_nvzMUPSq9_0),.clk(gclk));
	jdff dff_A_mFVKxGu34_0(.dout(w_dff_A_nvzMUPSq9_0),.din(w_dff_A_mFVKxGu34_0),.clk(gclk));
	jdff dff_A_irLXAV5G9_0(.dout(w_dff_A_mFVKxGu34_0),.din(w_dff_A_irLXAV5G9_0),.clk(gclk));
	jdff dff_A_RyDPdlYE3_0(.dout(w_dff_A_irLXAV5G9_0),.din(w_dff_A_RyDPdlYE3_0),.clk(gclk));
	jdff dff_A_cE9ToscC4_0(.dout(w_dff_A_RyDPdlYE3_0),.din(w_dff_A_cE9ToscC4_0),.clk(gclk));
	jdff dff_A_E4D3sfKA6_0(.dout(w_dff_A_cE9ToscC4_0),.din(w_dff_A_E4D3sfKA6_0),.clk(gclk));
	jdff dff_A_Jk9NLDmv1_0(.dout(w_dff_A_E4D3sfKA6_0),.din(w_dff_A_Jk9NLDmv1_0),.clk(gclk));
	jdff dff_A_MX7Ewhas0_0(.dout(w_dff_A_Jk9NLDmv1_0),.din(w_dff_A_MX7Ewhas0_0),.clk(gclk));
	jdff dff_A_B8nYgEY25_0(.dout(w_dff_A_MX7Ewhas0_0),.din(w_dff_A_B8nYgEY25_0),.clk(gclk));
	jdff dff_A_eZzfNJOH7_0(.dout(w_dff_A_B8nYgEY25_0),.din(w_dff_A_eZzfNJOH7_0),.clk(gclk));
	jdff dff_A_UsNuXq1X7_0(.dout(w_dff_A_eZzfNJOH7_0),.din(w_dff_A_UsNuXq1X7_0),.clk(gclk));
	jdff dff_A_MXIAfFn31_0(.dout(w_dff_A_UsNuXq1X7_0),.din(w_dff_A_MXIAfFn31_0),.clk(gclk));
	jdff dff_A_yO15gPJr5_0(.dout(w_dff_A_MXIAfFn31_0),.din(w_dff_A_yO15gPJr5_0),.clk(gclk));
	jdff dff_A_vP0gkV1y6_0(.dout(w_dff_A_yO15gPJr5_0),.din(w_dff_A_vP0gkV1y6_0),.clk(gclk));
	jdff dff_A_kdFHnUVh3_0(.dout(w_dff_A_vP0gkV1y6_0),.din(w_dff_A_kdFHnUVh3_0),.clk(gclk));
	jdff dff_A_Lm5Gs0yh8_0(.dout(w_dff_A_kdFHnUVh3_0),.din(w_dff_A_Lm5Gs0yh8_0),.clk(gclk));
	jdff dff_A_TOM3HrQ90_0(.dout(w_dff_A_Lm5Gs0yh8_0),.din(w_dff_A_TOM3HrQ90_0),.clk(gclk));
	jdff dff_A_dViOtFSk2_0(.dout(w_dff_A_TOM3HrQ90_0),.din(w_dff_A_dViOtFSk2_0),.clk(gclk));
	jdff dff_A_AZWB3P7r5_0(.dout(w_dff_A_dViOtFSk2_0),.din(w_dff_A_AZWB3P7r5_0),.clk(gclk));
	jdff dff_A_60ukqH3e5_0(.dout(w_dff_A_AZWB3P7r5_0),.din(w_dff_A_60ukqH3e5_0),.clk(gclk));
	jdff dff_A_k9uGuW0y1_0(.dout(w_dff_A_60ukqH3e5_0),.din(w_dff_A_k9uGuW0y1_0),.clk(gclk));
	jdff dff_A_aJjaHec75_0(.dout(w_dff_A_k9uGuW0y1_0),.din(w_dff_A_aJjaHec75_0),.clk(gclk));
	jdff dff_A_DnOZtxGb6_0(.dout(w_dff_A_aJjaHec75_0),.din(w_dff_A_DnOZtxGb6_0),.clk(gclk));
	jdff dff_A_KYdOX3r87_0(.dout(w_dff_A_DnOZtxGb6_0),.din(w_dff_A_KYdOX3r87_0),.clk(gclk));
	jdff dff_A_h8Kp11Vq8_0(.dout(w_dff_A_KYdOX3r87_0),.din(w_dff_A_h8Kp11Vq8_0),.clk(gclk));
	jdff dff_A_Bt6sxac45_0(.dout(w_dff_A_h8Kp11Vq8_0),.din(w_dff_A_Bt6sxac45_0),.clk(gclk));
	jdff dff_A_BPXW0qTw3_0(.dout(w_dff_A_Bt6sxac45_0),.din(w_dff_A_BPXW0qTw3_0),.clk(gclk));
	jdff dff_A_t55fvk2X7_0(.dout(w_dff_A_BPXW0qTw3_0),.din(w_dff_A_t55fvk2X7_0),.clk(gclk));
	jdff dff_A_MaHfv1FW1_0(.dout(w_dff_A_t55fvk2X7_0),.din(w_dff_A_MaHfv1FW1_0),.clk(gclk));
	jdff dff_A_Y7GbduvZ9_0(.dout(w_dff_A_MaHfv1FW1_0),.din(w_dff_A_Y7GbduvZ9_0),.clk(gclk));
	jdff dff_A_14xhSJk46_0(.dout(w_dff_A_Y7GbduvZ9_0),.din(w_dff_A_14xhSJk46_0),.clk(gclk));
	jdff dff_A_ImEE9lU15_0(.dout(w_dff_A_14xhSJk46_0),.din(w_dff_A_ImEE9lU15_0),.clk(gclk));
	jdff dff_A_iLKi4kvh6_0(.dout(w_dff_A_ImEE9lU15_0),.din(w_dff_A_iLKi4kvh6_0),.clk(gclk));
	jdff dff_A_9KENl70F9_0(.dout(w_dff_A_iLKi4kvh6_0),.din(w_dff_A_9KENl70F9_0),.clk(gclk));
	jdff dff_A_4Rx08WPt0_0(.dout(w_dff_A_9KENl70F9_0),.din(w_dff_A_4Rx08WPt0_0),.clk(gclk));
	jdff dff_A_RF7ZFcvi5_0(.dout(w_dff_A_4Rx08WPt0_0),.din(w_dff_A_RF7ZFcvi5_0),.clk(gclk));
	jdff dff_A_4Ww2YHwk1_0(.dout(w_dff_A_RF7ZFcvi5_0),.din(w_dff_A_4Ww2YHwk1_0),.clk(gclk));
	jdff dff_A_CozEEMQj4_0(.dout(w_n799_0[0]),.din(w_dff_A_CozEEMQj4_0),.clk(gclk));
	jdff dff_B_BOjcivN93_1(.din(n714),.dout(w_dff_B_BOjcivN93_1),.clk(gclk));
	jdff dff_A_BxerMc0E2_0(.dout(w_n620_0[0]),.din(w_dff_A_BxerMc0E2_0),.clk(gclk));
	jdff dff_A_cimKIYuX4_0(.dout(w_dff_A_BxerMc0E2_0),.din(w_dff_A_cimKIYuX4_0),.clk(gclk));
	jdff dff_A_WayADUjb1_0(.dout(w_dff_A_cimKIYuX4_0),.din(w_dff_A_WayADUjb1_0),.clk(gclk));
	jdff dff_A_KuDZC9I02_0(.dout(w_dff_A_WayADUjb1_0),.din(w_dff_A_KuDZC9I02_0),.clk(gclk));
	jdff dff_A_08M9oir51_0(.dout(w_dff_A_KuDZC9I02_0),.din(w_dff_A_08M9oir51_0),.clk(gclk));
	jdff dff_A_tL04Z9ZC3_0(.dout(w_dff_A_08M9oir51_0),.din(w_dff_A_tL04Z9ZC3_0),.clk(gclk));
	jdff dff_A_lQBRQG533_0(.dout(w_dff_A_tL04Z9ZC3_0),.din(w_dff_A_lQBRQG533_0),.clk(gclk));
	jdff dff_A_yc2Ulbxy7_0(.dout(w_dff_A_lQBRQG533_0),.din(w_dff_A_yc2Ulbxy7_0),.clk(gclk));
	jdff dff_A_WALWMKSr5_0(.dout(w_dff_A_yc2Ulbxy7_0),.din(w_dff_A_WALWMKSr5_0),.clk(gclk));
	jdff dff_A_kTz6nelh8_0(.dout(w_dff_A_WALWMKSr5_0),.din(w_dff_A_kTz6nelh8_0),.clk(gclk));
	jdff dff_A_CBnURHp55_0(.dout(w_dff_A_kTz6nelh8_0),.din(w_dff_A_CBnURHp55_0),.clk(gclk));
	jdff dff_A_FbDy6Hqa8_0(.dout(w_dff_A_CBnURHp55_0),.din(w_dff_A_FbDy6Hqa8_0),.clk(gclk));
	jdff dff_A_wE4lDe5G2_0(.dout(w_dff_A_FbDy6Hqa8_0),.din(w_dff_A_wE4lDe5G2_0),.clk(gclk));
	jdff dff_A_6gPJGe730_0(.dout(w_dff_A_wE4lDe5G2_0),.din(w_dff_A_6gPJGe730_0),.clk(gclk));
	jdff dff_A_VhV8I7eJ5_0(.dout(w_dff_A_6gPJGe730_0),.din(w_dff_A_VhV8I7eJ5_0),.clk(gclk));
	jdff dff_A_gzDa1RYH1_0(.dout(w_dff_A_VhV8I7eJ5_0),.din(w_dff_A_gzDa1RYH1_0),.clk(gclk));
	jdff dff_A_nwetkaC47_0(.dout(w_dff_A_gzDa1RYH1_0),.din(w_dff_A_nwetkaC47_0),.clk(gclk));
	jdff dff_A_9EQNKs7y2_0(.dout(w_dff_A_nwetkaC47_0),.din(w_dff_A_9EQNKs7y2_0),.clk(gclk));
	jdff dff_A_0n1Cb1087_0(.dout(w_dff_A_9EQNKs7y2_0),.din(w_dff_A_0n1Cb1087_0),.clk(gclk));
	jdff dff_A_0CZJAKpG5_0(.dout(w_dff_A_0n1Cb1087_0),.din(w_dff_A_0CZJAKpG5_0),.clk(gclk));
	jdff dff_A_X2SkhwMt9_0(.dout(w_dff_A_0CZJAKpG5_0),.din(w_dff_A_X2SkhwMt9_0),.clk(gclk));
	jdff dff_A_F5OZ1ssi3_0(.dout(w_dff_A_X2SkhwMt9_0),.din(w_dff_A_F5OZ1ssi3_0),.clk(gclk));
	jdff dff_A_f3oK9d4V5_0(.dout(w_dff_A_F5OZ1ssi3_0),.din(w_dff_A_f3oK9d4V5_0),.clk(gclk));
	jdff dff_A_lOdRId168_0(.dout(w_dff_A_f3oK9d4V5_0),.din(w_dff_A_lOdRId168_0),.clk(gclk));
	jdff dff_A_SyaBC5oX3_0(.dout(w_dff_A_lOdRId168_0),.din(w_dff_A_SyaBC5oX3_0),.clk(gclk));
	jdff dff_A_PNUyjw2S6_0(.dout(w_dff_A_SyaBC5oX3_0),.din(w_dff_A_PNUyjw2S6_0),.clk(gclk));
	jdff dff_A_VHH0K7Fk1_0(.dout(w_dff_A_PNUyjw2S6_0),.din(w_dff_A_VHH0K7Fk1_0),.clk(gclk));
	jdff dff_A_I0vO1TjO2_0(.dout(w_dff_A_VHH0K7Fk1_0),.din(w_dff_A_I0vO1TjO2_0),.clk(gclk));
	jdff dff_A_QcxV2Gco2_0(.dout(w_dff_A_I0vO1TjO2_0),.din(w_dff_A_QcxV2Gco2_0),.clk(gclk));
	jdff dff_A_Uz29G7AQ7_0(.dout(w_dff_A_QcxV2Gco2_0),.din(w_dff_A_Uz29G7AQ7_0),.clk(gclk));
	jdff dff_A_AALeN3uJ1_0(.dout(w_dff_A_Uz29G7AQ7_0),.din(w_dff_A_AALeN3uJ1_0),.clk(gclk));
	jdff dff_A_VUxJTziZ8_0(.dout(w_dff_A_AALeN3uJ1_0),.din(w_dff_A_VUxJTziZ8_0),.clk(gclk));
	jdff dff_A_8AzY1BgI9_0(.dout(w_dff_A_VUxJTziZ8_0),.din(w_dff_A_8AzY1BgI9_0),.clk(gclk));
	jdff dff_A_z3WtrQqV4_0(.dout(w_dff_A_8AzY1BgI9_0),.din(w_dff_A_z3WtrQqV4_0),.clk(gclk));
	jdff dff_A_UaJP31Zr4_0(.dout(w_n700_0[0]),.din(w_dff_A_UaJP31Zr4_0),.clk(gclk));
	jdff dff_B_L54OtKa01_1(.din(n622),.dout(w_dff_B_L54OtKa01_1),.clk(gclk));
	jdff dff_A_j5LpYyAI9_0(.dout(w_n535_0[0]),.din(w_dff_A_j5LpYyAI9_0),.clk(gclk));
	jdff dff_A_4GuMcs7N8_0(.dout(w_dff_A_j5LpYyAI9_0),.din(w_dff_A_4GuMcs7N8_0),.clk(gclk));
	jdff dff_A_p0kP9c4r6_0(.dout(w_dff_A_4GuMcs7N8_0),.din(w_dff_A_p0kP9c4r6_0),.clk(gclk));
	jdff dff_A_za4cIv037_0(.dout(w_dff_A_p0kP9c4r6_0),.din(w_dff_A_za4cIv037_0),.clk(gclk));
	jdff dff_A_wAJFscVw8_0(.dout(w_dff_A_za4cIv037_0),.din(w_dff_A_wAJFscVw8_0),.clk(gclk));
	jdff dff_A_b7g7ZcYN2_0(.dout(w_dff_A_wAJFscVw8_0),.din(w_dff_A_b7g7ZcYN2_0),.clk(gclk));
	jdff dff_A_z2ZGlGEA4_0(.dout(w_dff_A_b7g7ZcYN2_0),.din(w_dff_A_z2ZGlGEA4_0),.clk(gclk));
	jdff dff_A_umsH6zCL8_0(.dout(w_dff_A_z2ZGlGEA4_0),.din(w_dff_A_umsH6zCL8_0),.clk(gclk));
	jdff dff_A_JLlDFbRd2_0(.dout(w_dff_A_umsH6zCL8_0),.din(w_dff_A_JLlDFbRd2_0),.clk(gclk));
	jdff dff_A_x5KzGJFz5_0(.dout(w_dff_A_JLlDFbRd2_0),.din(w_dff_A_x5KzGJFz5_0),.clk(gclk));
	jdff dff_A_NdGpRJNo7_0(.dout(w_dff_A_x5KzGJFz5_0),.din(w_dff_A_NdGpRJNo7_0),.clk(gclk));
	jdff dff_A_MvVhzOVP0_0(.dout(w_dff_A_NdGpRJNo7_0),.din(w_dff_A_MvVhzOVP0_0),.clk(gclk));
	jdff dff_A_mh6JhjAo7_0(.dout(w_dff_A_MvVhzOVP0_0),.din(w_dff_A_mh6JhjAo7_0),.clk(gclk));
	jdff dff_A_7hFL9iPU2_0(.dout(w_dff_A_mh6JhjAo7_0),.din(w_dff_A_7hFL9iPU2_0),.clk(gclk));
	jdff dff_A_zEVAQUr66_0(.dout(w_dff_A_7hFL9iPU2_0),.din(w_dff_A_zEVAQUr66_0),.clk(gclk));
	jdff dff_A_SnifY13u4_0(.dout(w_dff_A_zEVAQUr66_0),.din(w_dff_A_SnifY13u4_0),.clk(gclk));
	jdff dff_A_k3fn1NIj1_0(.dout(w_dff_A_SnifY13u4_0),.din(w_dff_A_k3fn1NIj1_0),.clk(gclk));
	jdff dff_A_6zqEzYZu6_0(.dout(w_dff_A_k3fn1NIj1_0),.din(w_dff_A_6zqEzYZu6_0),.clk(gclk));
	jdff dff_A_7XWCDsIC5_0(.dout(w_dff_A_6zqEzYZu6_0),.din(w_dff_A_7XWCDsIC5_0),.clk(gclk));
	jdff dff_A_fNutgw799_0(.dout(w_dff_A_7XWCDsIC5_0),.din(w_dff_A_fNutgw799_0),.clk(gclk));
	jdff dff_A_rUtuXh2z2_0(.dout(w_dff_A_fNutgw799_0),.din(w_dff_A_rUtuXh2z2_0),.clk(gclk));
	jdff dff_A_X6Mg3W7K6_0(.dout(w_dff_A_rUtuXh2z2_0),.din(w_dff_A_X6Mg3W7K6_0),.clk(gclk));
	jdff dff_A_WuETERNJ9_0(.dout(w_dff_A_X6Mg3W7K6_0),.din(w_dff_A_WuETERNJ9_0),.clk(gclk));
	jdff dff_A_m8Rt0BIM9_0(.dout(w_dff_A_WuETERNJ9_0),.din(w_dff_A_m8Rt0BIM9_0),.clk(gclk));
	jdff dff_A_ZhwonHSi7_0(.dout(w_dff_A_m8Rt0BIM9_0),.din(w_dff_A_ZhwonHSi7_0),.clk(gclk));
	jdff dff_A_CULjJBlH4_0(.dout(w_dff_A_ZhwonHSi7_0),.din(w_dff_A_CULjJBlH4_0),.clk(gclk));
	jdff dff_A_TdxwIVvD1_0(.dout(w_dff_A_CULjJBlH4_0),.din(w_dff_A_TdxwIVvD1_0),.clk(gclk));
	jdff dff_A_HfS7QI0y6_0(.dout(w_dff_A_TdxwIVvD1_0),.din(w_dff_A_HfS7QI0y6_0),.clk(gclk));
	jdff dff_A_bim36IMe0_0(.dout(w_dff_A_HfS7QI0y6_0),.din(w_dff_A_bim36IMe0_0),.clk(gclk));
	jdff dff_A_PDCWZ8WG3_0(.dout(w_dff_A_bim36IMe0_0),.din(w_dff_A_PDCWZ8WG3_0),.clk(gclk));
	jdff dff_A_fuaXEbQU2_0(.dout(w_dff_A_PDCWZ8WG3_0),.din(w_dff_A_fuaXEbQU2_0),.clk(gclk));
	jdff dff_A_tK0LOVYt9_0(.dout(w_n608_0[0]),.din(w_dff_A_tK0LOVYt9_0),.clk(gclk));
	jdff dff_B_25LyZmhv8_1(.din(n537),.dout(w_dff_B_25LyZmhv8_1),.clk(gclk));
	jdff dff_A_1DTD4n8o4_0(.dout(w_n457_0[0]),.din(w_dff_A_1DTD4n8o4_0),.clk(gclk));
	jdff dff_A_27Vjn8E55_0(.dout(w_dff_A_1DTD4n8o4_0),.din(w_dff_A_27Vjn8E55_0),.clk(gclk));
	jdff dff_A_BliCZHBw1_0(.dout(w_dff_A_27Vjn8E55_0),.din(w_dff_A_BliCZHBw1_0),.clk(gclk));
	jdff dff_A_fXjxcnL24_0(.dout(w_dff_A_BliCZHBw1_0),.din(w_dff_A_fXjxcnL24_0),.clk(gclk));
	jdff dff_A_HOjB8P6M0_0(.dout(w_dff_A_fXjxcnL24_0),.din(w_dff_A_HOjB8P6M0_0),.clk(gclk));
	jdff dff_A_1EmnySFl3_0(.dout(w_dff_A_HOjB8P6M0_0),.din(w_dff_A_1EmnySFl3_0),.clk(gclk));
	jdff dff_A_FuMXZAhx2_0(.dout(w_dff_A_1EmnySFl3_0),.din(w_dff_A_FuMXZAhx2_0),.clk(gclk));
	jdff dff_A_UxwMdAWx5_0(.dout(w_dff_A_FuMXZAhx2_0),.din(w_dff_A_UxwMdAWx5_0),.clk(gclk));
	jdff dff_A_pWCk4pl57_0(.dout(w_dff_A_UxwMdAWx5_0),.din(w_dff_A_pWCk4pl57_0),.clk(gclk));
	jdff dff_A_VAfjNRrt7_0(.dout(w_dff_A_pWCk4pl57_0),.din(w_dff_A_VAfjNRrt7_0),.clk(gclk));
	jdff dff_A_fOvk9cU14_0(.dout(w_dff_A_VAfjNRrt7_0),.din(w_dff_A_fOvk9cU14_0),.clk(gclk));
	jdff dff_A_wAk2BdGn2_0(.dout(w_dff_A_fOvk9cU14_0),.din(w_dff_A_wAk2BdGn2_0),.clk(gclk));
	jdff dff_A_Zz4QNO8u9_0(.dout(w_dff_A_wAk2BdGn2_0),.din(w_dff_A_Zz4QNO8u9_0),.clk(gclk));
	jdff dff_A_kqjg2sC43_0(.dout(w_dff_A_Zz4QNO8u9_0),.din(w_dff_A_kqjg2sC43_0),.clk(gclk));
	jdff dff_A_bHnznFdG8_0(.dout(w_dff_A_kqjg2sC43_0),.din(w_dff_A_bHnznFdG8_0),.clk(gclk));
	jdff dff_A_aVJMZtkD3_0(.dout(w_dff_A_bHnznFdG8_0),.din(w_dff_A_aVJMZtkD3_0),.clk(gclk));
	jdff dff_A_TliCd5nd7_0(.dout(w_dff_A_aVJMZtkD3_0),.din(w_dff_A_TliCd5nd7_0),.clk(gclk));
	jdff dff_A_vgzIR9E05_0(.dout(w_dff_A_TliCd5nd7_0),.din(w_dff_A_vgzIR9E05_0),.clk(gclk));
	jdff dff_A_86JmCiBZ5_0(.dout(w_dff_A_vgzIR9E05_0),.din(w_dff_A_86JmCiBZ5_0),.clk(gclk));
	jdff dff_A_z9Z0vJC13_0(.dout(w_dff_A_86JmCiBZ5_0),.din(w_dff_A_z9Z0vJC13_0),.clk(gclk));
	jdff dff_A_bVLbzTMZ9_0(.dout(w_dff_A_z9Z0vJC13_0),.din(w_dff_A_bVLbzTMZ9_0),.clk(gclk));
	jdff dff_A_OanEgcdL1_0(.dout(w_dff_A_bVLbzTMZ9_0),.din(w_dff_A_OanEgcdL1_0),.clk(gclk));
	jdff dff_A_ZQtBZvJU8_0(.dout(w_dff_A_OanEgcdL1_0),.din(w_dff_A_ZQtBZvJU8_0),.clk(gclk));
	jdff dff_A_qfSXjFBA6_0(.dout(w_dff_A_ZQtBZvJU8_0),.din(w_dff_A_qfSXjFBA6_0),.clk(gclk));
	jdff dff_A_L6IHRjm13_0(.dout(w_dff_A_qfSXjFBA6_0),.din(w_dff_A_L6IHRjm13_0),.clk(gclk));
	jdff dff_A_4Wo6oDnA2_0(.dout(w_dff_A_L6IHRjm13_0),.din(w_dff_A_4Wo6oDnA2_0),.clk(gclk));
	jdff dff_A_CqY9cvf81_0(.dout(w_dff_A_4Wo6oDnA2_0),.din(w_dff_A_CqY9cvf81_0),.clk(gclk));
	jdff dff_A_ufPHR4DL3_0(.dout(w_dff_A_CqY9cvf81_0),.din(w_dff_A_ufPHR4DL3_0),.clk(gclk));
	jdff dff_A_ZUZuYvs31_0(.dout(w_n523_0[0]),.din(w_dff_A_ZUZuYvs31_0),.clk(gclk));
	jdff dff_B_n8ulN2hL2_1(.din(n459),.dout(w_dff_B_n8ulN2hL2_1),.clk(gclk));
	jdff dff_A_xjivaEHV1_0(.dout(w_n386_0[0]),.din(w_dff_A_xjivaEHV1_0),.clk(gclk));
	jdff dff_A_ZvFdidse1_0(.dout(w_dff_A_xjivaEHV1_0),.din(w_dff_A_ZvFdidse1_0),.clk(gclk));
	jdff dff_A_xFCNRFwu0_0(.dout(w_dff_A_ZvFdidse1_0),.din(w_dff_A_xFCNRFwu0_0),.clk(gclk));
	jdff dff_A_Kua27kwP5_0(.dout(w_dff_A_xFCNRFwu0_0),.din(w_dff_A_Kua27kwP5_0),.clk(gclk));
	jdff dff_A_1FeNvmBt3_0(.dout(w_dff_A_Kua27kwP5_0),.din(w_dff_A_1FeNvmBt3_0),.clk(gclk));
	jdff dff_A_IxzFZAqA6_0(.dout(w_dff_A_1FeNvmBt3_0),.din(w_dff_A_IxzFZAqA6_0),.clk(gclk));
	jdff dff_A_2qGJEOFE4_0(.dout(w_dff_A_IxzFZAqA6_0),.din(w_dff_A_2qGJEOFE4_0),.clk(gclk));
	jdff dff_A_kaogT0kH7_0(.dout(w_dff_A_2qGJEOFE4_0),.din(w_dff_A_kaogT0kH7_0),.clk(gclk));
	jdff dff_A_bKpgsxEn1_0(.dout(w_dff_A_kaogT0kH7_0),.din(w_dff_A_bKpgsxEn1_0),.clk(gclk));
	jdff dff_A_NZwXKZmx8_0(.dout(w_dff_A_bKpgsxEn1_0),.din(w_dff_A_NZwXKZmx8_0),.clk(gclk));
	jdff dff_A_KHPVtjxh0_0(.dout(w_dff_A_NZwXKZmx8_0),.din(w_dff_A_KHPVtjxh0_0),.clk(gclk));
	jdff dff_A_xrEJUqYf1_0(.dout(w_dff_A_KHPVtjxh0_0),.din(w_dff_A_xrEJUqYf1_0),.clk(gclk));
	jdff dff_A_jY8NaeET5_0(.dout(w_dff_A_xrEJUqYf1_0),.din(w_dff_A_jY8NaeET5_0),.clk(gclk));
	jdff dff_A_POqxp1OC9_0(.dout(w_dff_A_jY8NaeET5_0),.din(w_dff_A_POqxp1OC9_0),.clk(gclk));
	jdff dff_A_cgWZzR0d5_0(.dout(w_dff_A_POqxp1OC9_0),.din(w_dff_A_cgWZzR0d5_0),.clk(gclk));
	jdff dff_A_e5NLw3368_0(.dout(w_dff_A_cgWZzR0d5_0),.din(w_dff_A_e5NLw3368_0),.clk(gclk));
	jdff dff_A_L0BiFdBL6_0(.dout(w_dff_A_e5NLw3368_0),.din(w_dff_A_L0BiFdBL6_0),.clk(gclk));
	jdff dff_A_iW3Ri9iE7_0(.dout(w_dff_A_L0BiFdBL6_0),.din(w_dff_A_iW3Ri9iE7_0),.clk(gclk));
	jdff dff_A_xoUAkCg02_0(.dout(w_dff_A_iW3Ri9iE7_0),.din(w_dff_A_xoUAkCg02_0),.clk(gclk));
	jdff dff_A_K3HezAHJ7_0(.dout(w_dff_A_xoUAkCg02_0),.din(w_dff_A_K3HezAHJ7_0),.clk(gclk));
	jdff dff_A_HGeg1hHW6_0(.dout(w_dff_A_K3HezAHJ7_0),.din(w_dff_A_HGeg1hHW6_0),.clk(gclk));
	jdff dff_A_gL9w6xVe1_0(.dout(w_dff_A_HGeg1hHW6_0),.din(w_dff_A_gL9w6xVe1_0),.clk(gclk));
	jdff dff_A_w2bfYK5X3_0(.dout(w_dff_A_gL9w6xVe1_0),.din(w_dff_A_w2bfYK5X3_0),.clk(gclk));
	jdff dff_A_rkplaC5G5_0(.dout(w_dff_A_w2bfYK5X3_0),.din(w_dff_A_rkplaC5G5_0),.clk(gclk));
	jdff dff_A_9rwQQ0ko5_0(.dout(w_dff_A_rkplaC5G5_0),.din(w_dff_A_9rwQQ0ko5_0),.clk(gclk));
	jdff dff_A_WZktrhNT6_0(.dout(w_n445_0[0]),.din(w_dff_A_WZktrhNT6_0),.clk(gclk));
	jdff dff_B_XzZDx8md5_1(.din(n388),.dout(w_dff_B_XzZDx8md5_1),.clk(gclk));
	jdff dff_A_S8SNoUsr9_0(.dout(w_n323_0[0]),.din(w_dff_A_S8SNoUsr9_0),.clk(gclk));
	jdff dff_A_wpuGUwG39_0(.dout(w_dff_A_S8SNoUsr9_0),.din(w_dff_A_wpuGUwG39_0),.clk(gclk));
	jdff dff_A_FvzflmIP5_0(.dout(w_dff_A_wpuGUwG39_0),.din(w_dff_A_FvzflmIP5_0),.clk(gclk));
	jdff dff_A_X1Fed3WN2_0(.dout(w_dff_A_FvzflmIP5_0),.din(w_dff_A_X1Fed3WN2_0),.clk(gclk));
	jdff dff_A_4EEzFBoY1_0(.dout(w_dff_A_X1Fed3WN2_0),.din(w_dff_A_4EEzFBoY1_0),.clk(gclk));
	jdff dff_A_4guQfGBD0_0(.dout(w_dff_A_4EEzFBoY1_0),.din(w_dff_A_4guQfGBD0_0),.clk(gclk));
	jdff dff_A_wS0E1z5y9_0(.dout(w_dff_A_4guQfGBD0_0),.din(w_dff_A_wS0E1z5y9_0),.clk(gclk));
	jdff dff_A_YrXEYsNd4_0(.dout(w_dff_A_wS0E1z5y9_0),.din(w_dff_A_YrXEYsNd4_0),.clk(gclk));
	jdff dff_A_OjWPk9ni2_0(.dout(w_dff_A_YrXEYsNd4_0),.din(w_dff_A_OjWPk9ni2_0),.clk(gclk));
	jdff dff_A_YignJEAz3_0(.dout(w_dff_A_OjWPk9ni2_0),.din(w_dff_A_YignJEAz3_0),.clk(gclk));
	jdff dff_A_UPRj53l43_0(.dout(w_dff_A_YignJEAz3_0),.din(w_dff_A_UPRj53l43_0),.clk(gclk));
	jdff dff_A_RHGOpSsd7_0(.dout(w_dff_A_UPRj53l43_0),.din(w_dff_A_RHGOpSsd7_0),.clk(gclk));
	jdff dff_A_4aoOijak7_0(.dout(w_dff_A_RHGOpSsd7_0),.din(w_dff_A_4aoOijak7_0),.clk(gclk));
	jdff dff_A_6Ja7ZXuS3_0(.dout(w_dff_A_4aoOijak7_0),.din(w_dff_A_6Ja7ZXuS3_0),.clk(gclk));
	jdff dff_A_pWKTwEMx6_0(.dout(w_dff_A_6Ja7ZXuS3_0),.din(w_dff_A_pWKTwEMx6_0),.clk(gclk));
	jdff dff_A_7gdt2f474_0(.dout(w_dff_A_pWKTwEMx6_0),.din(w_dff_A_7gdt2f474_0),.clk(gclk));
	jdff dff_A_4U1aKAbU6_0(.dout(w_dff_A_7gdt2f474_0),.din(w_dff_A_4U1aKAbU6_0),.clk(gclk));
	jdff dff_A_28mJBR7X3_0(.dout(w_dff_A_4U1aKAbU6_0),.din(w_dff_A_28mJBR7X3_0),.clk(gclk));
	jdff dff_A_0vlo5Euv3_0(.dout(w_dff_A_28mJBR7X3_0),.din(w_dff_A_0vlo5Euv3_0),.clk(gclk));
	jdff dff_A_b3Uh1PC65_0(.dout(w_dff_A_0vlo5Euv3_0),.din(w_dff_A_b3Uh1PC65_0),.clk(gclk));
	jdff dff_A_GzMRwxlk0_0(.dout(w_dff_A_b3Uh1PC65_0),.din(w_dff_A_GzMRwxlk0_0),.clk(gclk));
	jdff dff_A_Y1PZdxHC4_0(.dout(w_dff_A_GzMRwxlk0_0),.din(w_dff_A_Y1PZdxHC4_0),.clk(gclk));
	jdff dff_A_pUfXEeqD8_0(.dout(w_n374_0[0]),.din(w_dff_A_pUfXEeqD8_0),.clk(gclk));
	jdff dff_B_qxEaHlTH9_1(.din(n325),.dout(w_dff_B_qxEaHlTH9_1),.clk(gclk));
	jdff dff_A_TgP2QZxM9_0(.dout(w_n267_0[0]),.din(w_dff_A_TgP2QZxM9_0),.clk(gclk));
	jdff dff_A_0OEhDnkf8_0(.dout(w_dff_A_TgP2QZxM9_0),.din(w_dff_A_0OEhDnkf8_0),.clk(gclk));
	jdff dff_A_OZmavzp60_0(.dout(w_dff_A_0OEhDnkf8_0),.din(w_dff_A_OZmavzp60_0),.clk(gclk));
	jdff dff_A_dUy6AJW28_0(.dout(w_dff_A_OZmavzp60_0),.din(w_dff_A_dUy6AJW28_0),.clk(gclk));
	jdff dff_A_eGm3zfLS4_0(.dout(w_dff_A_dUy6AJW28_0),.din(w_dff_A_eGm3zfLS4_0),.clk(gclk));
	jdff dff_A_Z04TkIfy3_0(.dout(w_dff_A_eGm3zfLS4_0),.din(w_dff_A_Z04TkIfy3_0),.clk(gclk));
	jdff dff_A_we4WEDFt3_0(.dout(w_dff_A_Z04TkIfy3_0),.din(w_dff_A_we4WEDFt3_0),.clk(gclk));
	jdff dff_A_KjXsNrp10_0(.dout(w_dff_A_we4WEDFt3_0),.din(w_dff_A_KjXsNrp10_0),.clk(gclk));
	jdff dff_A_rjJE9DLc2_0(.dout(w_dff_A_KjXsNrp10_0),.din(w_dff_A_rjJE9DLc2_0),.clk(gclk));
	jdff dff_A_glNc0pJw3_0(.dout(w_dff_A_rjJE9DLc2_0),.din(w_dff_A_glNc0pJw3_0),.clk(gclk));
	jdff dff_A_BEOL1gef2_0(.dout(w_dff_A_glNc0pJw3_0),.din(w_dff_A_BEOL1gef2_0),.clk(gclk));
	jdff dff_A_617rBd9v6_0(.dout(w_dff_A_BEOL1gef2_0),.din(w_dff_A_617rBd9v6_0),.clk(gclk));
	jdff dff_A_gUGhPz4P7_0(.dout(w_dff_A_617rBd9v6_0),.din(w_dff_A_gUGhPz4P7_0),.clk(gclk));
	jdff dff_A_SIE3Puh01_0(.dout(w_dff_A_gUGhPz4P7_0),.din(w_dff_A_SIE3Puh01_0),.clk(gclk));
	jdff dff_A_DuFthvhz9_0(.dout(w_dff_A_SIE3Puh01_0),.din(w_dff_A_DuFthvhz9_0),.clk(gclk));
	jdff dff_A_byQnZsMu2_0(.dout(w_dff_A_DuFthvhz9_0),.din(w_dff_A_byQnZsMu2_0),.clk(gclk));
	jdff dff_A_ggmsijOl8_0(.dout(w_dff_A_byQnZsMu2_0),.din(w_dff_A_ggmsijOl8_0),.clk(gclk));
	jdff dff_A_HEERYzqX3_0(.dout(w_dff_A_ggmsijOl8_0),.din(w_dff_A_HEERYzqX3_0),.clk(gclk));
	jdff dff_A_07ryFYOn6_0(.dout(w_dff_A_HEERYzqX3_0),.din(w_dff_A_07ryFYOn6_0),.clk(gclk));
	jdff dff_A_9FZh6byn6_0(.dout(w_n311_0[0]),.din(w_dff_A_9FZh6byn6_0),.clk(gclk));
	jdff dff_B_r4hNDjzn8_1(.din(n269),.dout(w_dff_B_r4hNDjzn8_1),.clk(gclk));
	jdff dff_A_I8DUMGoX0_0(.dout(w_n218_0[0]),.din(w_dff_A_I8DUMGoX0_0),.clk(gclk));
	jdff dff_A_Lq53wyEv9_0(.dout(w_dff_A_I8DUMGoX0_0),.din(w_dff_A_Lq53wyEv9_0),.clk(gclk));
	jdff dff_A_ZDDJNgU28_0(.dout(w_dff_A_Lq53wyEv9_0),.din(w_dff_A_ZDDJNgU28_0),.clk(gclk));
	jdff dff_A_lIx0bLKJ0_0(.dout(w_dff_A_ZDDJNgU28_0),.din(w_dff_A_lIx0bLKJ0_0),.clk(gclk));
	jdff dff_A_MfRrB5g66_0(.dout(w_dff_A_lIx0bLKJ0_0),.din(w_dff_A_MfRrB5g66_0),.clk(gclk));
	jdff dff_A_Y63wSNTp3_0(.dout(w_dff_A_MfRrB5g66_0),.din(w_dff_A_Y63wSNTp3_0),.clk(gclk));
	jdff dff_A_iwE2BmLL0_0(.dout(w_dff_A_Y63wSNTp3_0),.din(w_dff_A_iwE2BmLL0_0),.clk(gclk));
	jdff dff_A_I1qV6Jaa1_0(.dout(w_dff_A_iwE2BmLL0_0),.din(w_dff_A_I1qV6Jaa1_0),.clk(gclk));
	jdff dff_A_yRNag3fp1_0(.dout(w_dff_A_I1qV6Jaa1_0),.din(w_dff_A_yRNag3fp1_0),.clk(gclk));
	jdff dff_A_RlUYuPSY5_0(.dout(w_dff_A_yRNag3fp1_0),.din(w_dff_A_RlUYuPSY5_0),.clk(gclk));
	jdff dff_A_rAoiwxM79_0(.dout(w_dff_A_RlUYuPSY5_0),.din(w_dff_A_rAoiwxM79_0),.clk(gclk));
	jdff dff_A_k0fiZLEa3_0(.dout(w_dff_A_rAoiwxM79_0),.din(w_dff_A_k0fiZLEa3_0),.clk(gclk));
	jdff dff_A_aFVBh2xO5_0(.dout(w_dff_A_k0fiZLEa3_0),.din(w_dff_A_aFVBh2xO5_0),.clk(gclk));
	jdff dff_A_9jfXyD3y3_0(.dout(w_dff_A_aFVBh2xO5_0),.din(w_dff_A_9jfXyD3y3_0),.clk(gclk));
	jdff dff_A_U1tuxpQ13_0(.dout(w_dff_A_9jfXyD3y3_0),.din(w_dff_A_U1tuxpQ13_0),.clk(gclk));
	jdff dff_A_ZGD17F2e9_0(.dout(w_dff_A_U1tuxpQ13_0),.din(w_dff_A_ZGD17F2e9_0),.clk(gclk));
	jdff dff_A_nhN25l222_0(.dout(w_n255_0[0]),.din(w_dff_A_nhN25l222_0),.clk(gclk));
	jdff dff_B_3vhxBByS6_1(.din(n220),.dout(w_dff_B_3vhxBByS6_1),.clk(gclk));
	jdff dff_A_Ps0Tcvho8_0(.dout(w_n176_0[0]),.din(w_dff_A_Ps0Tcvho8_0),.clk(gclk));
	jdff dff_A_25z5P6Bh1_0(.dout(w_dff_A_Ps0Tcvho8_0),.din(w_dff_A_25z5P6Bh1_0),.clk(gclk));
	jdff dff_A_WkQvTt551_0(.dout(w_dff_A_25z5P6Bh1_0),.din(w_dff_A_WkQvTt551_0),.clk(gclk));
	jdff dff_A_npWI4njK8_0(.dout(w_dff_A_WkQvTt551_0),.din(w_dff_A_npWI4njK8_0),.clk(gclk));
	jdff dff_A_YRLimjjR8_0(.dout(w_dff_A_npWI4njK8_0),.din(w_dff_A_YRLimjjR8_0),.clk(gclk));
	jdff dff_A_jBdQNVfI9_0(.dout(w_dff_A_YRLimjjR8_0),.din(w_dff_A_jBdQNVfI9_0),.clk(gclk));
	jdff dff_A_7PdzuaE90_0(.dout(w_dff_A_jBdQNVfI9_0),.din(w_dff_A_7PdzuaE90_0),.clk(gclk));
	jdff dff_A_nA7dc5BY9_0(.dout(w_dff_A_7PdzuaE90_0),.din(w_dff_A_nA7dc5BY9_0),.clk(gclk));
	jdff dff_A_jhRbLA6Q7_0(.dout(w_dff_A_nA7dc5BY9_0),.din(w_dff_A_jhRbLA6Q7_0),.clk(gclk));
	jdff dff_A_4EuBYuut9_0(.dout(w_dff_A_jhRbLA6Q7_0),.din(w_dff_A_4EuBYuut9_0),.clk(gclk));
	jdff dff_A_yhwUhhM33_0(.dout(w_dff_A_4EuBYuut9_0),.din(w_dff_A_yhwUhhM33_0),.clk(gclk));
	jdff dff_A_m062pSjM0_0(.dout(w_dff_A_yhwUhhM33_0),.din(w_dff_A_m062pSjM0_0),.clk(gclk));
	jdff dff_A_Usx6TU591_0(.dout(w_dff_A_m062pSjM0_0),.din(w_dff_A_Usx6TU591_0),.clk(gclk));
	jdff dff_A_xTHqHmzl2_0(.dout(w_n206_0[0]),.din(w_dff_A_xTHqHmzl2_0),.clk(gclk));
	jdff dff_B_HfKmuf415_1(.din(n178),.dout(w_dff_B_HfKmuf415_1),.clk(gclk));
	jdff dff_A_0qNLck1J0_0(.dout(w_n141_0[0]),.din(w_dff_A_0qNLck1J0_0),.clk(gclk));
	jdff dff_A_17ZMACWF0_0(.dout(w_dff_A_0qNLck1J0_0),.din(w_dff_A_17ZMACWF0_0),.clk(gclk));
	jdff dff_A_Gc39vKPx9_0(.dout(w_dff_A_17ZMACWF0_0),.din(w_dff_A_Gc39vKPx9_0),.clk(gclk));
	jdff dff_A_RtNC1uB15_0(.dout(w_dff_A_Gc39vKPx9_0),.din(w_dff_A_RtNC1uB15_0),.clk(gclk));
	jdff dff_A_PV9EYaJr3_0(.dout(w_dff_A_RtNC1uB15_0),.din(w_dff_A_PV9EYaJr3_0),.clk(gclk));
	jdff dff_A_OMyJ6xQq8_0(.dout(w_dff_A_PV9EYaJr3_0),.din(w_dff_A_OMyJ6xQq8_0),.clk(gclk));
	jdff dff_A_UFZvJpGt8_0(.dout(w_dff_A_OMyJ6xQq8_0),.din(w_dff_A_UFZvJpGt8_0),.clk(gclk));
	jdff dff_A_E2NoMfwW0_0(.dout(w_dff_A_UFZvJpGt8_0),.din(w_dff_A_E2NoMfwW0_0),.clk(gclk));
	jdff dff_A_jALWbNxy6_0(.dout(w_dff_A_E2NoMfwW0_0),.din(w_dff_A_jALWbNxy6_0),.clk(gclk));
	jdff dff_A_Ub9v0iXs2_0(.dout(w_dff_A_jALWbNxy6_0),.din(w_dff_A_Ub9v0iXs2_0),.clk(gclk));
	jdff dff_A_uGHgRN7S4_0(.dout(w_n164_0[0]),.din(w_dff_A_uGHgRN7S4_0),.clk(gclk));
	jdff dff_B_BZ4iv02w0_1(.din(n143),.dout(w_dff_B_BZ4iv02w0_1),.clk(gclk));
	jdff dff_A_DMVcyFUf3_0(.dout(w_n112_0[0]),.din(w_dff_A_DMVcyFUf3_0),.clk(gclk));
	jdff dff_A_mIiBCANF5_0(.dout(w_dff_A_DMVcyFUf3_0),.din(w_dff_A_mIiBCANF5_0),.clk(gclk));
	jdff dff_A_oJ5GVM8I1_0(.dout(w_dff_A_mIiBCANF5_0),.din(w_dff_A_oJ5GVM8I1_0),.clk(gclk));
	jdff dff_A_lfYOIB5d5_0(.dout(w_dff_A_oJ5GVM8I1_0),.din(w_dff_A_lfYOIB5d5_0),.clk(gclk));
	jdff dff_A_3gPfbbnv4_0(.dout(w_dff_A_lfYOIB5d5_0),.din(w_dff_A_3gPfbbnv4_0),.clk(gclk));
	jdff dff_A_kYqYKoxr2_0(.dout(w_dff_A_3gPfbbnv4_0),.din(w_dff_A_kYqYKoxr2_0),.clk(gclk));
	jdff dff_A_yz2g5o3T1_0(.dout(w_dff_A_kYqYKoxr2_0),.din(w_dff_A_yz2g5o3T1_0),.clk(gclk));
	jdff dff_A_OcGInJTO8_0(.dout(w_n129_0[0]),.din(w_dff_A_OcGInJTO8_0),.clk(gclk));
	jdff dff_B_lka824er8_1(.din(n114),.dout(w_dff_B_lka824er8_1),.clk(gclk));
	jdff dff_A_ZdyDGYRF6_0(.dout(w_n91_0[0]),.din(w_dff_A_ZdyDGYRF6_0),.clk(gclk));
	jdff dff_A_7RScKASn6_0(.dout(w_dff_A_ZdyDGYRF6_0),.din(w_dff_A_7RScKASn6_0),.clk(gclk));
	jdff dff_A_G0LNzcrn8_0(.dout(w_dff_A_7RScKASn6_0),.din(w_dff_A_G0LNzcrn8_0),.clk(gclk));
	jdff dff_A_wyHhALjm2_0(.dout(w_dff_A_G0LNzcrn8_0),.din(w_dff_A_wyHhALjm2_0),.clk(gclk));
	jdff dff_B_AsRBWcbj0_0(.din(n100),.dout(w_dff_B_AsRBWcbj0_0),.clk(gclk));
	jdff dff_A_iGsqUyTS8_0(.dout(w_n80_0[0]),.din(w_dff_A_iGsqUyTS8_0),.clk(gclk));
	jdff dff_A_kHDRHVTJ0_0(.dout(w_n1119_0[0]),.din(w_dff_A_kHDRHVTJ0_0),.clk(gclk));
	jdff dff_B_cMjIhJEV7_2(.din(n1119),.dout(w_dff_B_cMjIhJEV7_2),.clk(gclk));
	jdff dff_B_sWP56mRH1_2(.din(n1018),.dout(w_dff_B_sWP56mRH1_2),.clk(gclk));
	jdff dff_B_z2gJh9B52_2(.din(w_dff_B_sWP56mRH1_2),.dout(w_dff_B_z2gJh9B52_2),.clk(gclk));
	jdff dff_B_s9MKeXFT0_2(.din(w_dff_B_z2gJh9B52_2),.dout(w_dff_B_s9MKeXFT0_2),.clk(gclk));
	jdff dff_B_BlJtStrS9_2(.din(w_dff_B_s9MKeXFT0_2),.dout(w_dff_B_BlJtStrS9_2),.clk(gclk));
	jdff dff_B_4ZrApfOc7_2(.din(w_dff_B_BlJtStrS9_2),.dout(w_dff_B_4ZrApfOc7_2),.clk(gclk));
	jdff dff_B_8WTIScRC8_2(.din(w_dff_B_4ZrApfOc7_2),.dout(w_dff_B_8WTIScRC8_2),.clk(gclk));
	jdff dff_B_aaE8ibXH6_2(.din(w_dff_B_8WTIScRC8_2),.dout(w_dff_B_aaE8ibXH6_2),.clk(gclk));
	jdff dff_B_p8XQ9mHl2_2(.din(w_dff_B_aaE8ibXH6_2),.dout(w_dff_B_p8XQ9mHl2_2),.clk(gclk));
	jdff dff_B_rsoZITgZ2_2(.din(w_dff_B_p8XQ9mHl2_2),.dout(w_dff_B_rsoZITgZ2_2),.clk(gclk));
	jdff dff_B_jskZ009W2_2(.din(w_dff_B_rsoZITgZ2_2),.dout(w_dff_B_jskZ009W2_2),.clk(gclk));
	jdff dff_B_xaX5NC4Z6_2(.din(w_dff_B_jskZ009W2_2),.dout(w_dff_B_xaX5NC4Z6_2),.clk(gclk));
	jdff dff_B_zVOHL91y4_2(.din(w_dff_B_xaX5NC4Z6_2),.dout(w_dff_B_zVOHL91y4_2),.clk(gclk));
	jdff dff_B_AoneoiBe9_2(.din(w_dff_B_zVOHL91y4_2),.dout(w_dff_B_AoneoiBe9_2),.clk(gclk));
	jdff dff_B_oa4YAf3i9_2(.din(w_dff_B_AoneoiBe9_2),.dout(w_dff_B_oa4YAf3i9_2),.clk(gclk));
	jdff dff_B_JsRxpWHk4_2(.din(w_dff_B_oa4YAf3i9_2),.dout(w_dff_B_JsRxpWHk4_2),.clk(gclk));
	jdff dff_B_V75BtALJ3_2(.din(w_dff_B_JsRxpWHk4_2),.dout(w_dff_B_V75BtALJ3_2),.clk(gclk));
	jdff dff_B_wMJb6RMj2_2(.din(w_dff_B_V75BtALJ3_2),.dout(w_dff_B_wMJb6RMj2_2),.clk(gclk));
	jdff dff_B_C2abLtti9_2(.din(w_dff_B_wMJb6RMj2_2),.dout(w_dff_B_C2abLtti9_2),.clk(gclk));
	jdff dff_B_aiyDfmbh1_2(.din(w_dff_B_C2abLtti9_2),.dout(w_dff_B_aiyDfmbh1_2),.clk(gclk));
	jdff dff_B_kFzdtis48_2(.din(w_dff_B_aiyDfmbh1_2),.dout(w_dff_B_kFzdtis48_2),.clk(gclk));
	jdff dff_B_9puinoJx4_2(.din(w_dff_B_kFzdtis48_2),.dout(w_dff_B_9puinoJx4_2),.clk(gclk));
	jdff dff_B_PJWfu2Pf8_2(.din(w_dff_B_9puinoJx4_2),.dout(w_dff_B_PJWfu2Pf8_2),.clk(gclk));
	jdff dff_B_DYGmZ1rB0_2(.din(w_dff_B_PJWfu2Pf8_2),.dout(w_dff_B_DYGmZ1rB0_2),.clk(gclk));
	jdff dff_B_9ImUXCEc7_2(.din(w_dff_B_DYGmZ1rB0_2),.dout(w_dff_B_9ImUXCEc7_2),.clk(gclk));
	jdff dff_B_AqnN7G0m1_2(.din(w_dff_B_9ImUXCEc7_2),.dout(w_dff_B_AqnN7G0m1_2),.clk(gclk));
	jdff dff_B_AGVbdhUS4_2(.din(w_dff_B_AqnN7G0m1_2),.dout(w_dff_B_AGVbdhUS4_2),.clk(gclk));
	jdff dff_B_ItjhBvyb7_2(.din(w_dff_B_AGVbdhUS4_2),.dout(w_dff_B_ItjhBvyb7_2),.clk(gclk));
	jdff dff_B_q11eEC790_2(.din(w_dff_B_ItjhBvyb7_2),.dout(w_dff_B_q11eEC790_2),.clk(gclk));
	jdff dff_B_GlJLWQMp1_2(.din(w_dff_B_q11eEC790_2),.dout(w_dff_B_GlJLWQMp1_2),.clk(gclk));
	jdff dff_B_w76aUxrT4_2(.din(w_dff_B_GlJLWQMp1_2),.dout(w_dff_B_w76aUxrT4_2),.clk(gclk));
	jdff dff_B_0gDijboI2_2(.din(w_dff_B_w76aUxrT4_2),.dout(w_dff_B_0gDijboI2_2),.clk(gclk));
	jdff dff_B_jGYKGauk4_2(.din(w_dff_B_0gDijboI2_2),.dout(w_dff_B_jGYKGauk4_2),.clk(gclk));
	jdff dff_B_rLjNOMb91_2(.din(w_dff_B_jGYKGauk4_2),.dout(w_dff_B_rLjNOMb91_2),.clk(gclk));
	jdff dff_B_zAdSHiSq5_2(.din(w_dff_B_rLjNOMb91_2),.dout(w_dff_B_zAdSHiSq5_2),.clk(gclk));
	jdff dff_B_2emaucSo3_2(.din(w_dff_B_zAdSHiSq5_2),.dout(w_dff_B_2emaucSo3_2),.clk(gclk));
	jdff dff_B_Eevua5uk6_2(.din(w_dff_B_2emaucSo3_2),.dout(w_dff_B_Eevua5uk6_2),.clk(gclk));
	jdff dff_B_shMmYz582_2(.din(w_dff_B_Eevua5uk6_2),.dout(w_dff_B_shMmYz582_2),.clk(gclk));
	jdff dff_B_NZ4Gurnf1_2(.din(w_dff_B_shMmYz582_2),.dout(w_dff_B_NZ4Gurnf1_2),.clk(gclk));
	jdff dff_B_htANaIDt2_2(.din(w_dff_B_NZ4Gurnf1_2),.dout(w_dff_B_htANaIDt2_2),.clk(gclk));
	jdff dff_B_lJ5FMkbB7_2(.din(w_dff_B_htANaIDt2_2),.dout(w_dff_B_lJ5FMkbB7_2),.clk(gclk));
	jdff dff_B_F9pzeo6i8_2(.din(w_dff_B_lJ5FMkbB7_2),.dout(w_dff_B_F9pzeo6i8_2),.clk(gclk));
	jdff dff_B_eu71PbNQ2_2(.din(w_dff_B_F9pzeo6i8_2),.dout(w_dff_B_eu71PbNQ2_2),.clk(gclk));
	jdff dff_B_SYqhYXJy0_2(.din(w_dff_B_eu71PbNQ2_2),.dout(w_dff_B_SYqhYXJy0_2),.clk(gclk));
	jdff dff_A_pjjutMCB9_0(.dout(w_n1022_0[0]),.din(w_dff_A_pjjutMCB9_0),.clk(gclk));
	jdff dff_B_YGBk4d6B0_1(.din(n1020),.dout(w_dff_B_YGBk4d6B0_1),.clk(gclk));
	jdff dff_B_DNzvvfS67_2(.din(n916),.dout(w_dff_B_DNzvvfS67_2),.clk(gclk));
	jdff dff_B_9PEsjT5o3_2(.din(w_dff_B_DNzvvfS67_2),.dout(w_dff_B_9PEsjT5o3_2),.clk(gclk));
	jdff dff_B_F9IZMHeN6_2(.din(w_dff_B_9PEsjT5o3_2),.dout(w_dff_B_F9IZMHeN6_2),.clk(gclk));
	jdff dff_B_n4xbpcwy0_2(.din(w_dff_B_F9IZMHeN6_2),.dout(w_dff_B_n4xbpcwy0_2),.clk(gclk));
	jdff dff_B_TX0PA1M27_2(.din(w_dff_B_n4xbpcwy0_2),.dout(w_dff_B_TX0PA1M27_2),.clk(gclk));
	jdff dff_B_s0ldgvR69_2(.din(w_dff_B_TX0PA1M27_2),.dout(w_dff_B_s0ldgvR69_2),.clk(gclk));
	jdff dff_B_ufuef6bT3_2(.din(w_dff_B_s0ldgvR69_2),.dout(w_dff_B_ufuef6bT3_2),.clk(gclk));
	jdff dff_B_AWDttdoo6_2(.din(w_dff_B_ufuef6bT3_2),.dout(w_dff_B_AWDttdoo6_2),.clk(gclk));
	jdff dff_B_46xmwMo04_2(.din(w_dff_B_AWDttdoo6_2),.dout(w_dff_B_46xmwMo04_2),.clk(gclk));
	jdff dff_B_DdNHP23u2_2(.din(w_dff_B_46xmwMo04_2),.dout(w_dff_B_DdNHP23u2_2),.clk(gclk));
	jdff dff_B_3si6Bylu5_2(.din(w_dff_B_DdNHP23u2_2),.dout(w_dff_B_3si6Bylu5_2),.clk(gclk));
	jdff dff_B_6md3Pfvk6_2(.din(w_dff_B_3si6Bylu5_2),.dout(w_dff_B_6md3Pfvk6_2),.clk(gclk));
	jdff dff_B_zMoJKukp6_2(.din(w_dff_B_6md3Pfvk6_2),.dout(w_dff_B_zMoJKukp6_2),.clk(gclk));
	jdff dff_B_T7pmnkJE6_2(.din(w_dff_B_zMoJKukp6_2),.dout(w_dff_B_T7pmnkJE6_2),.clk(gclk));
	jdff dff_B_pJFDvR551_2(.din(w_dff_B_T7pmnkJE6_2),.dout(w_dff_B_pJFDvR551_2),.clk(gclk));
	jdff dff_B_XdTbbgsw2_2(.din(w_dff_B_pJFDvR551_2),.dout(w_dff_B_XdTbbgsw2_2),.clk(gclk));
	jdff dff_B_3GcBCU8N6_2(.din(w_dff_B_XdTbbgsw2_2),.dout(w_dff_B_3GcBCU8N6_2),.clk(gclk));
	jdff dff_B_ONcR3NhH2_2(.din(w_dff_B_3GcBCU8N6_2),.dout(w_dff_B_ONcR3NhH2_2),.clk(gclk));
	jdff dff_B_mKjN1i3f4_2(.din(w_dff_B_ONcR3NhH2_2),.dout(w_dff_B_mKjN1i3f4_2),.clk(gclk));
	jdff dff_B_bLNxqumJ4_2(.din(w_dff_B_mKjN1i3f4_2),.dout(w_dff_B_bLNxqumJ4_2),.clk(gclk));
	jdff dff_B_bBPrEfQk3_2(.din(w_dff_B_bLNxqumJ4_2),.dout(w_dff_B_bBPrEfQk3_2),.clk(gclk));
	jdff dff_B_dfR48Bq79_2(.din(w_dff_B_bBPrEfQk3_2),.dout(w_dff_B_dfR48Bq79_2),.clk(gclk));
	jdff dff_B_tkF1pB0Z6_2(.din(w_dff_B_dfR48Bq79_2),.dout(w_dff_B_tkF1pB0Z6_2),.clk(gclk));
	jdff dff_B_4DlmKAeM9_2(.din(w_dff_B_tkF1pB0Z6_2),.dout(w_dff_B_4DlmKAeM9_2),.clk(gclk));
	jdff dff_B_6oKVEMCU6_2(.din(w_dff_B_4DlmKAeM9_2),.dout(w_dff_B_6oKVEMCU6_2),.clk(gclk));
	jdff dff_B_EnQPCE8p7_2(.din(w_dff_B_6oKVEMCU6_2),.dout(w_dff_B_EnQPCE8p7_2),.clk(gclk));
	jdff dff_B_cHf5ylHZ9_2(.din(w_dff_B_EnQPCE8p7_2),.dout(w_dff_B_cHf5ylHZ9_2),.clk(gclk));
	jdff dff_B_BAK4Yd0c4_2(.din(w_dff_B_cHf5ylHZ9_2),.dout(w_dff_B_BAK4Yd0c4_2),.clk(gclk));
	jdff dff_B_SlQVWnTe7_2(.din(w_dff_B_BAK4Yd0c4_2),.dout(w_dff_B_SlQVWnTe7_2),.clk(gclk));
	jdff dff_B_S8kf8kxz5_2(.din(w_dff_B_SlQVWnTe7_2),.dout(w_dff_B_S8kf8kxz5_2),.clk(gclk));
	jdff dff_B_fsWyEvLm5_2(.din(w_dff_B_S8kf8kxz5_2),.dout(w_dff_B_fsWyEvLm5_2),.clk(gclk));
	jdff dff_B_kvg1jy7G3_2(.din(w_dff_B_fsWyEvLm5_2),.dout(w_dff_B_kvg1jy7G3_2),.clk(gclk));
	jdff dff_B_zxP7er6f1_2(.din(w_dff_B_kvg1jy7G3_2),.dout(w_dff_B_zxP7er6f1_2),.clk(gclk));
	jdff dff_B_lYmcxQpE6_2(.din(w_dff_B_zxP7er6f1_2),.dout(w_dff_B_lYmcxQpE6_2),.clk(gclk));
	jdff dff_B_dDExMTO48_2(.din(w_dff_B_lYmcxQpE6_2),.dout(w_dff_B_dDExMTO48_2),.clk(gclk));
	jdff dff_B_vl2mcgNi2_2(.din(w_dff_B_dDExMTO48_2),.dout(w_dff_B_vl2mcgNi2_2),.clk(gclk));
	jdff dff_B_TgsGOfhP3_2(.din(w_dff_B_vl2mcgNi2_2),.dout(w_dff_B_TgsGOfhP3_2),.clk(gclk));
	jdff dff_B_DyxWsHIf6_2(.din(w_dff_B_TgsGOfhP3_2),.dout(w_dff_B_DyxWsHIf6_2),.clk(gclk));
	jdff dff_B_aPoveLqF9_2(.din(w_dff_B_DyxWsHIf6_2),.dout(w_dff_B_aPoveLqF9_2),.clk(gclk));
	jdff dff_B_h1Ll7FdX5_2(.din(w_dff_B_aPoveLqF9_2),.dout(w_dff_B_h1Ll7FdX5_2),.clk(gclk));
	jdff dff_A_hK4FPsXJ4_1(.dout(w_n1006_0[1]),.din(w_dff_A_hK4FPsXJ4_1),.clk(gclk));
	jdff dff_A_IkfscCdt0_0(.dout(w_n816_0[0]),.din(w_dff_A_IkfscCdt0_0),.clk(gclk));
	jdff dff_A_o7mAy3Ez9_0(.dout(w_dff_A_IkfscCdt0_0),.din(w_dff_A_o7mAy3Ez9_0),.clk(gclk));
	jdff dff_A_0GxAqjJG5_0(.dout(w_dff_A_o7mAy3Ez9_0),.din(w_dff_A_0GxAqjJG5_0),.clk(gclk));
	jdff dff_A_5SACCQAh5_0(.dout(w_dff_A_0GxAqjJG5_0),.din(w_dff_A_5SACCQAh5_0),.clk(gclk));
	jdff dff_A_Ik0Oth9e5_0(.dout(w_dff_A_5SACCQAh5_0),.din(w_dff_A_Ik0Oth9e5_0),.clk(gclk));
	jdff dff_A_nsYC6Hbg7_0(.dout(w_dff_A_Ik0Oth9e5_0),.din(w_dff_A_nsYC6Hbg7_0),.clk(gclk));
	jdff dff_A_An1SyVrE2_0(.dout(w_dff_A_nsYC6Hbg7_0),.din(w_dff_A_An1SyVrE2_0),.clk(gclk));
	jdff dff_A_M7gSdpXs0_0(.dout(w_dff_A_An1SyVrE2_0),.din(w_dff_A_M7gSdpXs0_0),.clk(gclk));
	jdff dff_A_5rpS1fqF4_0(.dout(w_dff_A_M7gSdpXs0_0),.din(w_dff_A_5rpS1fqF4_0),.clk(gclk));
	jdff dff_A_pSdRuKNy8_0(.dout(w_dff_A_5rpS1fqF4_0),.din(w_dff_A_pSdRuKNy8_0),.clk(gclk));
	jdff dff_A_XKVGVf5W9_0(.dout(w_dff_A_pSdRuKNy8_0),.din(w_dff_A_XKVGVf5W9_0),.clk(gclk));
	jdff dff_A_VWHnLsL63_0(.dout(w_dff_A_XKVGVf5W9_0),.din(w_dff_A_VWHnLsL63_0),.clk(gclk));
	jdff dff_A_WEnicOu88_0(.dout(w_dff_A_VWHnLsL63_0),.din(w_dff_A_WEnicOu88_0),.clk(gclk));
	jdff dff_A_1zrSoqdJ3_0(.dout(w_dff_A_WEnicOu88_0),.din(w_dff_A_1zrSoqdJ3_0),.clk(gclk));
	jdff dff_A_yVQzp8SB4_0(.dout(w_dff_A_1zrSoqdJ3_0),.din(w_dff_A_yVQzp8SB4_0),.clk(gclk));
	jdff dff_A_xslBY8zI0_0(.dout(w_dff_A_yVQzp8SB4_0),.din(w_dff_A_xslBY8zI0_0),.clk(gclk));
	jdff dff_A_35C7cfdF6_0(.dout(w_dff_A_xslBY8zI0_0),.din(w_dff_A_35C7cfdF6_0),.clk(gclk));
	jdff dff_A_8cBoGORk7_0(.dout(w_dff_A_35C7cfdF6_0),.din(w_dff_A_8cBoGORk7_0),.clk(gclk));
	jdff dff_A_egw93r2D5_0(.dout(w_dff_A_8cBoGORk7_0),.din(w_dff_A_egw93r2D5_0),.clk(gclk));
	jdff dff_A_WZxTySWC9_0(.dout(w_dff_A_egw93r2D5_0),.din(w_dff_A_WZxTySWC9_0),.clk(gclk));
	jdff dff_A_DZBG9ZFJ8_0(.dout(w_dff_A_WZxTySWC9_0),.din(w_dff_A_DZBG9ZFJ8_0),.clk(gclk));
	jdff dff_A_R99VK25B9_0(.dout(w_dff_A_DZBG9ZFJ8_0),.din(w_dff_A_R99VK25B9_0),.clk(gclk));
	jdff dff_A_wHvWHxvY7_0(.dout(w_dff_A_R99VK25B9_0),.din(w_dff_A_wHvWHxvY7_0),.clk(gclk));
	jdff dff_A_Q1y6kjRc2_0(.dout(w_dff_A_wHvWHxvY7_0),.din(w_dff_A_Q1y6kjRc2_0),.clk(gclk));
	jdff dff_A_JRrZcsmk8_0(.dout(w_dff_A_Q1y6kjRc2_0),.din(w_dff_A_JRrZcsmk8_0),.clk(gclk));
	jdff dff_A_LYjliNrx4_0(.dout(w_dff_A_JRrZcsmk8_0),.din(w_dff_A_LYjliNrx4_0),.clk(gclk));
	jdff dff_A_vGqp6JRk5_0(.dout(w_dff_A_LYjliNrx4_0),.din(w_dff_A_vGqp6JRk5_0),.clk(gclk));
	jdff dff_A_mR8NV3dy0_0(.dout(w_dff_A_vGqp6JRk5_0),.din(w_dff_A_mR8NV3dy0_0),.clk(gclk));
	jdff dff_A_lBdYvBH87_0(.dout(w_dff_A_mR8NV3dy0_0),.din(w_dff_A_lBdYvBH87_0),.clk(gclk));
	jdff dff_A_RC3CelW55_0(.dout(w_dff_A_lBdYvBH87_0),.din(w_dff_A_RC3CelW55_0),.clk(gclk));
	jdff dff_A_YHXS3FzX4_0(.dout(w_dff_A_RC3CelW55_0),.din(w_dff_A_YHXS3FzX4_0),.clk(gclk));
	jdff dff_A_WlHj1mDf7_0(.dout(w_dff_A_YHXS3FzX4_0),.din(w_dff_A_WlHj1mDf7_0),.clk(gclk));
	jdff dff_A_eaK2RJ0m7_0(.dout(w_dff_A_WlHj1mDf7_0),.din(w_dff_A_eaK2RJ0m7_0),.clk(gclk));
	jdff dff_A_uca9syKp0_0(.dout(w_dff_A_eaK2RJ0m7_0),.din(w_dff_A_uca9syKp0_0),.clk(gclk));
	jdff dff_A_lio901276_0(.dout(w_dff_A_uca9syKp0_0),.din(w_dff_A_lio901276_0),.clk(gclk));
	jdff dff_A_1EnTW8GZ1_0(.dout(w_dff_A_lio901276_0),.din(w_dff_A_1EnTW8GZ1_0),.clk(gclk));
	jdff dff_A_4lszyFn33_0(.dout(w_dff_A_1EnTW8GZ1_0),.din(w_dff_A_4lszyFn33_0),.clk(gclk));
	jdff dff_A_PaeTrKK39_1(.dout(w_n900_0[1]),.din(w_dff_A_PaeTrKK39_1),.clk(gclk));
	jdff dff_A_1ezDC40J1_2(.dout(w_n900_0[2]),.din(w_dff_A_1ezDC40J1_2),.clk(gclk));
	jdff dff_B_S4ORdUCC3_1(.din(n818),.dout(w_dff_B_S4ORdUCC3_1),.clk(gclk));
	jdff dff_B_OKyzk8Am3_2(.din(n719),.dout(w_dff_B_OKyzk8Am3_2),.clk(gclk));
	jdff dff_B_QrOMOxpq3_2(.din(w_dff_B_OKyzk8Am3_2),.dout(w_dff_B_QrOMOxpq3_2),.clk(gclk));
	jdff dff_B_HQ5mZaLc5_2(.din(w_dff_B_QrOMOxpq3_2),.dout(w_dff_B_HQ5mZaLc5_2),.clk(gclk));
	jdff dff_B_mWzklsGZ8_2(.din(w_dff_B_HQ5mZaLc5_2),.dout(w_dff_B_mWzklsGZ8_2),.clk(gclk));
	jdff dff_B_sPbXZwBI1_2(.din(w_dff_B_mWzklsGZ8_2),.dout(w_dff_B_sPbXZwBI1_2),.clk(gclk));
	jdff dff_B_Hy6mtHDx0_2(.din(w_dff_B_sPbXZwBI1_2),.dout(w_dff_B_Hy6mtHDx0_2),.clk(gclk));
	jdff dff_B_x3l5EV4w5_2(.din(w_dff_B_Hy6mtHDx0_2),.dout(w_dff_B_x3l5EV4w5_2),.clk(gclk));
	jdff dff_B_4cEYmsvB1_2(.din(w_dff_B_x3l5EV4w5_2),.dout(w_dff_B_4cEYmsvB1_2),.clk(gclk));
	jdff dff_B_8MIdHzbJ5_2(.din(w_dff_B_4cEYmsvB1_2),.dout(w_dff_B_8MIdHzbJ5_2),.clk(gclk));
	jdff dff_B_kdifOqQd7_2(.din(w_dff_B_8MIdHzbJ5_2),.dout(w_dff_B_kdifOqQd7_2),.clk(gclk));
	jdff dff_B_vrR4YgeA2_2(.din(w_dff_B_kdifOqQd7_2),.dout(w_dff_B_vrR4YgeA2_2),.clk(gclk));
	jdff dff_B_lJIkTdyN4_2(.din(w_dff_B_vrR4YgeA2_2),.dout(w_dff_B_lJIkTdyN4_2),.clk(gclk));
	jdff dff_B_jDm2Xwa08_2(.din(w_dff_B_lJIkTdyN4_2),.dout(w_dff_B_jDm2Xwa08_2),.clk(gclk));
	jdff dff_B_RYTP8VTC3_2(.din(w_dff_B_jDm2Xwa08_2),.dout(w_dff_B_RYTP8VTC3_2),.clk(gclk));
	jdff dff_B_HFKsYVuF3_2(.din(w_dff_B_RYTP8VTC3_2),.dout(w_dff_B_HFKsYVuF3_2),.clk(gclk));
	jdff dff_B_I4ktasz51_2(.din(w_dff_B_HFKsYVuF3_2),.dout(w_dff_B_I4ktasz51_2),.clk(gclk));
	jdff dff_B_nw3p254o3_2(.din(w_dff_B_I4ktasz51_2),.dout(w_dff_B_nw3p254o3_2),.clk(gclk));
	jdff dff_B_QimNdpqH1_2(.din(w_dff_B_nw3p254o3_2),.dout(w_dff_B_QimNdpqH1_2),.clk(gclk));
	jdff dff_B_mbMrcQet5_2(.din(w_dff_B_QimNdpqH1_2),.dout(w_dff_B_mbMrcQet5_2),.clk(gclk));
	jdff dff_B_dy8Lzjex8_2(.din(w_dff_B_mbMrcQet5_2),.dout(w_dff_B_dy8Lzjex8_2),.clk(gclk));
	jdff dff_B_30BLDKRy9_2(.din(w_dff_B_dy8Lzjex8_2),.dout(w_dff_B_30BLDKRy9_2),.clk(gclk));
	jdff dff_B_1NGgOigZ9_2(.din(w_dff_B_30BLDKRy9_2),.dout(w_dff_B_1NGgOigZ9_2),.clk(gclk));
	jdff dff_B_FN4SjH7s3_2(.din(w_dff_B_1NGgOigZ9_2),.dout(w_dff_B_FN4SjH7s3_2),.clk(gclk));
	jdff dff_B_Ppqrb9gF4_2(.din(w_dff_B_FN4SjH7s3_2),.dout(w_dff_B_Ppqrb9gF4_2),.clk(gclk));
	jdff dff_B_ikvOKAlh6_2(.din(w_dff_B_Ppqrb9gF4_2),.dout(w_dff_B_ikvOKAlh6_2),.clk(gclk));
	jdff dff_B_3TVZMWGu1_2(.din(w_dff_B_ikvOKAlh6_2),.dout(w_dff_B_3TVZMWGu1_2),.clk(gclk));
	jdff dff_B_KW8k5q2W6_2(.din(w_dff_B_3TVZMWGu1_2),.dout(w_dff_B_KW8k5q2W6_2),.clk(gclk));
	jdff dff_B_JAMLgE5S9_2(.din(w_dff_B_KW8k5q2W6_2),.dout(w_dff_B_JAMLgE5S9_2),.clk(gclk));
	jdff dff_B_xLQ3FboZ2_2(.din(w_dff_B_JAMLgE5S9_2),.dout(w_dff_B_xLQ3FboZ2_2),.clk(gclk));
	jdff dff_B_SuUU2NdK7_2(.din(w_dff_B_xLQ3FboZ2_2),.dout(w_dff_B_SuUU2NdK7_2),.clk(gclk));
	jdff dff_B_6GiWr4pP6_2(.din(w_dff_B_SuUU2NdK7_2),.dout(w_dff_B_6GiWr4pP6_2),.clk(gclk));
	jdff dff_B_iI2UZcQj6_2(.din(w_dff_B_6GiWr4pP6_2),.dout(w_dff_B_iI2UZcQj6_2),.clk(gclk));
	jdff dff_B_48MqtL2S3_2(.din(w_dff_B_iI2UZcQj6_2),.dout(w_dff_B_48MqtL2S3_2),.clk(gclk));
	jdff dff_B_Ch8v8ZGe5_2(.din(n797),.dout(w_dff_B_Ch8v8ZGe5_2),.clk(gclk));
	jdff dff_B_HgCApr8i9_1(.din(n720),.dout(w_dff_B_HgCApr8i9_1),.clk(gclk));
	jdff dff_B_7rpKxDZC5_2(.din(n627),.dout(w_dff_B_7rpKxDZC5_2),.clk(gclk));
	jdff dff_B_PA0FYVIU6_2(.din(w_dff_B_7rpKxDZC5_2),.dout(w_dff_B_PA0FYVIU6_2),.clk(gclk));
	jdff dff_B_udIlobvs4_2(.din(w_dff_B_PA0FYVIU6_2),.dout(w_dff_B_udIlobvs4_2),.clk(gclk));
	jdff dff_B_4RYQuMem5_2(.din(w_dff_B_udIlobvs4_2),.dout(w_dff_B_4RYQuMem5_2),.clk(gclk));
	jdff dff_B_CrwMvU7m9_2(.din(w_dff_B_4RYQuMem5_2),.dout(w_dff_B_CrwMvU7m9_2),.clk(gclk));
	jdff dff_B_tNMH12mS0_2(.din(w_dff_B_CrwMvU7m9_2),.dout(w_dff_B_tNMH12mS0_2),.clk(gclk));
	jdff dff_B_l5jHD8MR4_2(.din(w_dff_B_tNMH12mS0_2),.dout(w_dff_B_l5jHD8MR4_2),.clk(gclk));
	jdff dff_B_qePmiZwV4_2(.din(w_dff_B_l5jHD8MR4_2),.dout(w_dff_B_qePmiZwV4_2),.clk(gclk));
	jdff dff_B_OLuMQmi39_2(.din(w_dff_B_qePmiZwV4_2),.dout(w_dff_B_OLuMQmi39_2),.clk(gclk));
	jdff dff_B_8KIr8lb44_2(.din(w_dff_B_OLuMQmi39_2),.dout(w_dff_B_8KIr8lb44_2),.clk(gclk));
	jdff dff_B_czveACIn4_2(.din(w_dff_B_8KIr8lb44_2),.dout(w_dff_B_czveACIn4_2),.clk(gclk));
	jdff dff_B_hAZy3l651_2(.din(w_dff_B_czveACIn4_2),.dout(w_dff_B_hAZy3l651_2),.clk(gclk));
	jdff dff_B_NQ8nkmsP1_2(.din(w_dff_B_hAZy3l651_2),.dout(w_dff_B_NQ8nkmsP1_2),.clk(gclk));
	jdff dff_B_fk6Cz92y8_2(.din(w_dff_B_NQ8nkmsP1_2),.dout(w_dff_B_fk6Cz92y8_2),.clk(gclk));
	jdff dff_B_ZqHVFzJZ2_2(.din(w_dff_B_fk6Cz92y8_2),.dout(w_dff_B_ZqHVFzJZ2_2),.clk(gclk));
	jdff dff_B_mTFfpFVL5_2(.din(w_dff_B_ZqHVFzJZ2_2),.dout(w_dff_B_mTFfpFVL5_2),.clk(gclk));
	jdff dff_B_GDRo23Pv9_2(.din(w_dff_B_mTFfpFVL5_2),.dout(w_dff_B_GDRo23Pv9_2),.clk(gclk));
	jdff dff_B_QiA1G6pS1_2(.din(w_dff_B_GDRo23Pv9_2),.dout(w_dff_B_QiA1G6pS1_2),.clk(gclk));
	jdff dff_B_niBFkt3b7_2(.din(w_dff_B_QiA1G6pS1_2),.dout(w_dff_B_niBFkt3b7_2),.clk(gclk));
	jdff dff_B_QKoQBLWg2_2(.din(w_dff_B_niBFkt3b7_2),.dout(w_dff_B_QKoQBLWg2_2),.clk(gclk));
	jdff dff_B_HEmFGvd54_2(.din(w_dff_B_QKoQBLWg2_2),.dout(w_dff_B_HEmFGvd54_2),.clk(gclk));
	jdff dff_B_mKI4ZSl27_2(.din(w_dff_B_HEmFGvd54_2),.dout(w_dff_B_mKI4ZSl27_2),.clk(gclk));
	jdff dff_B_jULFZCLS9_2(.din(w_dff_B_mKI4ZSl27_2),.dout(w_dff_B_jULFZCLS9_2),.clk(gclk));
	jdff dff_B_KtQEJS3O6_2(.din(w_dff_B_jULFZCLS9_2),.dout(w_dff_B_KtQEJS3O6_2),.clk(gclk));
	jdff dff_B_IYezIVQ78_2(.din(w_dff_B_KtQEJS3O6_2),.dout(w_dff_B_IYezIVQ78_2),.clk(gclk));
	jdff dff_B_foWNZZ9p7_2(.din(w_dff_B_IYezIVQ78_2),.dout(w_dff_B_foWNZZ9p7_2),.clk(gclk));
	jdff dff_B_UZL6lfpx4_2(.din(w_dff_B_foWNZZ9p7_2),.dout(w_dff_B_UZL6lfpx4_2),.clk(gclk));
	jdff dff_B_ZPYN26713_2(.din(w_dff_B_UZL6lfpx4_2),.dout(w_dff_B_ZPYN26713_2),.clk(gclk));
	jdff dff_B_ellVHP0T5_2(.din(w_dff_B_ZPYN26713_2),.dout(w_dff_B_ellVHP0T5_2),.clk(gclk));
	jdff dff_B_QaEcDSuD5_2(.din(w_dff_B_ellVHP0T5_2),.dout(w_dff_B_QaEcDSuD5_2),.clk(gclk));
	jdff dff_B_TJA2DPQ43_2(.din(n698),.dout(w_dff_B_TJA2DPQ43_2),.clk(gclk));
	jdff dff_B_AAk7rBFR0_1(.din(n628),.dout(w_dff_B_AAk7rBFR0_1),.clk(gclk));
	jdff dff_B_ZWLLn9iO4_2(.din(n542),.dout(w_dff_B_ZWLLn9iO4_2),.clk(gclk));
	jdff dff_B_B5DJdmPx2_2(.din(w_dff_B_ZWLLn9iO4_2),.dout(w_dff_B_B5DJdmPx2_2),.clk(gclk));
	jdff dff_B_B0ltlHbD7_2(.din(w_dff_B_B5DJdmPx2_2),.dout(w_dff_B_B0ltlHbD7_2),.clk(gclk));
	jdff dff_B_rtksfZyz1_2(.din(w_dff_B_B0ltlHbD7_2),.dout(w_dff_B_rtksfZyz1_2),.clk(gclk));
	jdff dff_B_IZqBLimd3_2(.din(w_dff_B_rtksfZyz1_2),.dout(w_dff_B_IZqBLimd3_2),.clk(gclk));
	jdff dff_B_L5uThb3m5_2(.din(w_dff_B_IZqBLimd3_2),.dout(w_dff_B_L5uThb3m5_2),.clk(gclk));
	jdff dff_B_edTWyWv18_2(.din(w_dff_B_L5uThb3m5_2),.dout(w_dff_B_edTWyWv18_2),.clk(gclk));
	jdff dff_B_oXxetAOU7_2(.din(w_dff_B_edTWyWv18_2),.dout(w_dff_B_oXxetAOU7_2),.clk(gclk));
	jdff dff_B_buIo5cxD3_2(.din(w_dff_B_oXxetAOU7_2),.dout(w_dff_B_buIo5cxD3_2),.clk(gclk));
	jdff dff_B_OzSw6qXi9_2(.din(w_dff_B_buIo5cxD3_2),.dout(w_dff_B_OzSw6qXi9_2),.clk(gclk));
	jdff dff_B_TiI6N7T87_2(.din(w_dff_B_OzSw6qXi9_2),.dout(w_dff_B_TiI6N7T87_2),.clk(gclk));
	jdff dff_B_RCrHm3Xz7_2(.din(w_dff_B_TiI6N7T87_2),.dout(w_dff_B_RCrHm3Xz7_2),.clk(gclk));
	jdff dff_B_it2SQyoQ9_2(.din(w_dff_B_RCrHm3Xz7_2),.dout(w_dff_B_it2SQyoQ9_2),.clk(gclk));
	jdff dff_B_QMs1OM2m9_2(.din(w_dff_B_it2SQyoQ9_2),.dout(w_dff_B_QMs1OM2m9_2),.clk(gclk));
	jdff dff_B_ybz9E4168_2(.din(w_dff_B_QMs1OM2m9_2),.dout(w_dff_B_ybz9E4168_2),.clk(gclk));
	jdff dff_B_zgUtsPIU0_2(.din(w_dff_B_ybz9E4168_2),.dout(w_dff_B_zgUtsPIU0_2),.clk(gclk));
	jdff dff_B_95oHT9fe1_2(.din(w_dff_B_zgUtsPIU0_2),.dout(w_dff_B_95oHT9fe1_2),.clk(gclk));
	jdff dff_B_eRILAvIh6_2(.din(w_dff_B_95oHT9fe1_2),.dout(w_dff_B_eRILAvIh6_2),.clk(gclk));
	jdff dff_B_Md6ppQSk7_2(.din(w_dff_B_eRILAvIh6_2),.dout(w_dff_B_Md6ppQSk7_2),.clk(gclk));
	jdff dff_B_etzLcrmj9_2(.din(w_dff_B_Md6ppQSk7_2),.dout(w_dff_B_etzLcrmj9_2),.clk(gclk));
	jdff dff_B_SinFgzVt4_2(.din(w_dff_B_etzLcrmj9_2),.dout(w_dff_B_SinFgzVt4_2),.clk(gclk));
	jdff dff_B_SvLkIe8e0_2(.din(w_dff_B_SinFgzVt4_2),.dout(w_dff_B_SvLkIe8e0_2),.clk(gclk));
	jdff dff_B_1q12hnRw7_2(.din(w_dff_B_SvLkIe8e0_2),.dout(w_dff_B_1q12hnRw7_2),.clk(gclk));
	jdff dff_B_xBntAbYr8_2(.din(w_dff_B_1q12hnRw7_2),.dout(w_dff_B_xBntAbYr8_2),.clk(gclk));
	jdff dff_B_An2QI8fG8_2(.din(w_dff_B_xBntAbYr8_2),.dout(w_dff_B_An2QI8fG8_2),.clk(gclk));
	jdff dff_B_ehX91O2y4_2(.din(w_dff_B_An2QI8fG8_2),.dout(w_dff_B_ehX91O2y4_2),.clk(gclk));
	jdff dff_B_SabJs8jz7_2(.din(w_dff_B_ehX91O2y4_2),.dout(w_dff_B_SabJs8jz7_2),.clk(gclk));
	jdff dff_B_hR5poCbV0_2(.din(n606),.dout(w_dff_B_hR5poCbV0_2),.clk(gclk));
	jdff dff_B_E0zn4wyP8_1(.din(n543),.dout(w_dff_B_E0zn4wyP8_1),.clk(gclk));
	jdff dff_B_ZZyPhveW8_2(.din(n464),.dout(w_dff_B_ZZyPhveW8_2),.clk(gclk));
	jdff dff_B_MIqa1AyF2_2(.din(w_dff_B_ZZyPhveW8_2),.dout(w_dff_B_MIqa1AyF2_2),.clk(gclk));
	jdff dff_B_qBmtmQtj2_2(.din(w_dff_B_MIqa1AyF2_2),.dout(w_dff_B_qBmtmQtj2_2),.clk(gclk));
	jdff dff_B_rd3rvPc38_2(.din(w_dff_B_qBmtmQtj2_2),.dout(w_dff_B_rd3rvPc38_2),.clk(gclk));
	jdff dff_B_usGTkVpu1_2(.din(w_dff_B_rd3rvPc38_2),.dout(w_dff_B_usGTkVpu1_2),.clk(gclk));
	jdff dff_B_825KKHae9_2(.din(w_dff_B_usGTkVpu1_2),.dout(w_dff_B_825KKHae9_2),.clk(gclk));
	jdff dff_B_N8ROcOzd9_2(.din(w_dff_B_825KKHae9_2),.dout(w_dff_B_N8ROcOzd9_2),.clk(gclk));
	jdff dff_B_xYtmxULo3_2(.din(w_dff_B_N8ROcOzd9_2),.dout(w_dff_B_xYtmxULo3_2),.clk(gclk));
	jdff dff_B_nrQD752S8_2(.din(w_dff_B_xYtmxULo3_2),.dout(w_dff_B_nrQD752S8_2),.clk(gclk));
	jdff dff_B_EMqMMHyE5_2(.din(w_dff_B_nrQD752S8_2),.dout(w_dff_B_EMqMMHyE5_2),.clk(gclk));
	jdff dff_B_Q106ELUE1_2(.din(w_dff_B_EMqMMHyE5_2),.dout(w_dff_B_Q106ELUE1_2),.clk(gclk));
	jdff dff_B_uaLusQio5_2(.din(w_dff_B_Q106ELUE1_2),.dout(w_dff_B_uaLusQio5_2),.clk(gclk));
	jdff dff_B_q8welTEc0_2(.din(w_dff_B_uaLusQio5_2),.dout(w_dff_B_q8welTEc0_2),.clk(gclk));
	jdff dff_B_oDDvjCoj2_2(.din(w_dff_B_q8welTEc0_2),.dout(w_dff_B_oDDvjCoj2_2),.clk(gclk));
	jdff dff_B_8HwWkaG32_2(.din(w_dff_B_oDDvjCoj2_2),.dout(w_dff_B_8HwWkaG32_2),.clk(gclk));
	jdff dff_B_MIVvcWb63_2(.din(w_dff_B_8HwWkaG32_2),.dout(w_dff_B_MIVvcWb63_2),.clk(gclk));
	jdff dff_B_B0z1MmyT0_2(.din(w_dff_B_MIVvcWb63_2),.dout(w_dff_B_B0z1MmyT0_2),.clk(gclk));
	jdff dff_B_9EBzyWvx7_2(.din(w_dff_B_B0z1MmyT0_2),.dout(w_dff_B_9EBzyWvx7_2),.clk(gclk));
	jdff dff_B_5monQgmX4_2(.din(w_dff_B_9EBzyWvx7_2),.dout(w_dff_B_5monQgmX4_2),.clk(gclk));
	jdff dff_B_rmr0cjqc3_2(.din(w_dff_B_5monQgmX4_2),.dout(w_dff_B_rmr0cjqc3_2),.clk(gclk));
	jdff dff_B_ULDb7L4G2_2(.din(w_dff_B_rmr0cjqc3_2),.dout(w_dff_B_ULDb7L4G2_2),.clk(gclk));
	jdff dff_B_TtEmYi327_2(.din(w_dff_B_ULDb7L4G2_2),.dout(w_dff_B_TtEmYi327_2),.clk(gclk));
	jdff dff_B_w0Tkh8XO5_2(.din(w_dff_B_TtEmYi327_2),.dout(w_dff_B_w0Tkh8XO5_2),.clk(gclk));
	jdff dff_B_q57hWTjr9_2(.din(w_dff_B_w0Tkh8XO5_2),.dout(w_dff_B_q57hWTjr9_2),.clk(gclk));
	jdff dff_B_0xyfVBWM7_2(.din(n521),.dout(w_dff_B_0xyfVBWM7_2),.clk(gclk));
	jdff dff_B_Jh6lq4521_1(.din(n465),.dout(w_dff_B_Jh6lq4521_1),.clk(gclk));
	jdff dff_B_lANTmmel5_2(.din(n393),.dout(w_dff_B_lANTmmel5_2),.clk(gclk));
	jdff dff_B_0ZG2LOSb2_2(.din(w_dff_B_lANTmmel5_2),.dout(w_dff_B_0ZG2LOSb2_2),.clk(gclk));
	jdff dff_B_c7ztxUz32_2(.din(w_dff_B_0ZG2LOSb2_2),.dout(w_dff_B_c7ztxUz32_2),.clk(gclk));
	jdff dff_B_sXmtubWl5_2(.din(w_dff_B_c7ztxUz32_2),.dout(w_dff_B_sXmtubWl5_2),.clk(gclk));
	jdff dff_B_yb5GS2Gt2_2(.din(w_dff_B_sXmtubWl5_2),.dout(w_dff_B_yb5GS2Gt2_2),.clk(gclk));
	jdff dff_B_mtJ3BfXa4_2(.din(w_dff_B_yb5GS2Gt2_2),.dout(w_dff_B_mtJ3BfXa4_2),.clk(gclk));
	jdff dff_B_KDc0nzDV6_2(.din(w_dff_B_mtJ3BfXa4_2),.dout(w_dff_B_KDc0nzDV6_2),.clk(gclk));
	jdff dff_B_k8XBaHQ05_2(.din(w_dff_B_KDc0nzDV6_2),.dout(w_dff_B_k8XBaHQ05_2),.clk(gclk));
	jdff dff_B_lJSoHneo5_2(.din(w_dff_B_k8XBaHQ05_2),.dout(w_dff_B_lJSoHneo5_2),.clk(gclk));
	jdff dff_B_NSEFXBjI0_2(.din(w_dff_B_lJSoHneo5_2),.dout(w_dff_B_NSEFXBjI0_2),.clk(gclk));
	jdff dff_B_rMwsg27l6_2(.din(w_dff_B_NSEFXBjI0_2),.dout(w_dff_B_rMwsg27l6_2),.clk(gclk));
	jdff dff_B_BgW5oD0n5_2(.din(w_dff_B_rMwsg27l6_2),.dout(w_dff_B_BgW5oD0n5_2),.clk(gclk));
	jdff dff_B_KZPQY57t3_2(.din(w_dff_B_BgW5oD0n5_2),.dout(w_dff_B_KZPQY57t3_2),.clk(gclk));
	jdff dff_B_B70Eamoi1_2(.din(w_dff_B_KZPQY57t3_2),.dout(w_dff_B_B70Eamoi1_2),.clk(gclk));
	jdff dff_B_Jl3RscIH9_2(.din(w_dff_B_B70Eamoi1_2),.dout(w_dff_B_Jl3RscIH9_2),.clk(gclk));
	jdff dff_B_LcQSTCgc3_2(.din(w_dff_B_Jl3RscIH9_2),.dout(w_dff_B_LcQSTCgc3_2),.clk(gclk));
	jdff dff_B_UduQqCAt0_2(.din(w_dff_B_LcQSTCgc3_2),.dout(w_dff_B_UduQqCAt0_2),.clk(gclk));
	jdff dff_B_mzj2trgd0_2(.din(w_dff_B_UduQqCAt0_2),.dout(w_dff_B_mzj2trgd0_2),.clk(gclk));
	jdff dff_B_uUV632eO3_2(.din(w_dff_B_mzj2trgd0_2),.dout(w_dff_B_uUV632eO3_2),.clk(gclk));
	jdff dff_B_KPaKpPg85_2(.din(w_dff_B_uUV632eO3_2),.dout(w_dff_B_KPaKpPg85_2),.clk(gclk));
	jdff dff_B_TLAx6knM4_2(.din(w_dff_B_KPaKpPg85_2),.dout(w_dff_B_TLAx6knM4_2),.clk(gclk));
	jdff dff_B_1M3mdTob1_2(.din(n443),.dout(w_dff_B_1M3mdTob1_2),.clk(gclk));
	jdff dff_B_ZPrv69rY1_1(.din(n394),.dout(w_dff_B_ZPrv69rY1_1),.clk(gclk));
	jdff dff_B_lLyytNMO4_2(.din(n330),.dout(w_dff_B_lLyytNMO4_2),.clk(gclk));
	jdff dff_B_q9Gu2eiS7_2(.din(w_dff_B_lLyytNMO4_2),.dout(w_dff_B_q9Gu2eiS7_2),.clk(gclk));
	jdff dff_B_Qnk4Z3XI8_2(.din(w_dff_B_q9Gu2eiS7_2),.dout(w_dff_B_Qnk4Z3XI8_2),.clk(gclk));
	jdff dff_B_JDG4hyvH6_2(.din(w_dff_B_Qnk4Z3XI8_2),.dout(w_dff_B_JDG4hyvH6_2),.clk(gclk));
	jdff dff_B_YibEVKDh6_2(.din(w_dff_B_JDG4hyvH6_2),.dout(w_dff_B_YibEVKDh6_2),.clk(gclk));
	jdff dff_B_mbI4Fcqw5_2(.din(w_dff_B_YibEVKDh6_2),.dout(w_dff_B_mbI4Fcqw5_2),.clk(gclk));
	jdff dff_B_TYspeDOi8_2(.din(w_dff_B_mbI4Fcqw5_2),.dout(w_dff_B_TYspeDOi8_2),.clk(gclk));
	jdff dff_B_I7HuwlUW0_2(.din(w_dff_B_TYspeDOi8_2),.dout(w_dff_B_I7HuwlUW0_2),.clk(gclk));
	jdff dff_B_ZJeV8KQq0_2(.din(w_dff_B_I7HuwlUW0_2),.dout(w_dff_B_ZJeV8KQq0_2),.clk(gclk));
	jdff dff_B_UyzBVT2o6_2(.din(w_dff_B_ZJeV8KQq0_2),.dout(w_dff_B_UyzBVT2o6_2),.clk(gclk));
	jdff dff_B_D39Jdf8i9_2(.din(w_dff_B_UyzBVT2o6_2),.dout(w_dff_B_D39Jdf8i9_2),.clk(gclk));
	jdff dff_B_0ErRhg7G6_2(.din(w_dff_B_D39Jdf8i9_2),.dout(w_dff_B_0ErRhg7G6_2),.clk(gclk));
	jdff dff_B_V8zmzqOd3_2(.din(w_dff_B_0ErRhg7G6_2),.dout(w_dff_B_V8zmzqOd3_2),.clk(gclk));
	jdff dff_B_vlvm1FA74_2(.din(w_dff_B_V8zmzqOd3_2),.dout(w_dff_B_vlvm1FA74_2),.clk(gclk));
	jdff dff_B_Odve1Lhe6_2(.din(w_dff_B_vlvm1FA74_2),.dout(w_dff_B_Odve1Lhe6_2),.clk(gclk));
	jdff dff_B_delXOXpE8_2(.din(w_dff_B_Odve1Lhe6_2),.dout(w_dff_B_delXOXpE8_2),.clk(gclk));
	jdff dff_B_bvDYa1ZN5_2(.din(w_dff_B_delXOXpE8_2),.dout(w_dff_B_bvDYa1ZN5_2),.clk(gclk));
	jdff dff_B_ciueZflC7_2(.din(w_dff_B_bvDYa1ZN5_2),.dout(w_dff_B_ciueZflC7_2),.clk(gclk));
	jdff dff_B_sqKLcQOC4_2(.din(n372),.dout(w_dff_B_sqKLcQOC4_2),.clk(gclk));
	jdff dff_B_TLyREf666_1(.din(n331),.dout(w_dff_B_TLyREf666_1),.clk(gclk));
	jdff dff_B_IrrZjGgS5_2(.din(n274),.dout(w_dff_B_IrrZjGgS5_2),.clk(gclk));
	jdff dff_B_cGe2yHM70_2(.din(w_dff_B_IrrZjGgS5_2),.dout(w_dff_B_cGe2yHM70_2),.clk(gclk));
	jdff dff_B_1wgzXjHn1_2(.din(w_dff_B_cGe2yHM70_2),.dout(w_dff_B_1wgzXjHn1_2),.clk(gclk));
	jdff dff_B_1jjrzbDi0_2(.din(w_dff_B_1wgzXjHn1_2),.dout(w_dff_B_1jjrzbDi0_2),.clk(gclk));
	jdff dff_B_heFUKkxg4_2(.din(w_dff_B_1jjrzbDi0_2),.dout(w_dff_B_heFUKkxg4_2),.clk(gclk));
	jdff dff_B_1VszxwXr2_2(.din(w_dff_B_heFUKkxg4_2),.dout(w_dff_B_1VszxwXr2_2),.clk(gclk));
	jdff dff_B_csLb90T36_2(.din(w_dff_B_1VszxwXr2_2),.dout(w_dff_B_csLb90T36_2),.clk(gclk));
	jdff dff_B_R6PbYK4y9_2(.din(w_dff_B_csLb90T36_2),.dout(w_dff_B_R6PbYK4y9_2),.clk(gclk));
	jdff dff_B_T7akaYFz9_2(.din(w_dff_B_R6PbYK4y9_2),.dout(w_dff_B_T7akaYFz9_2),.clk(gclk));
	jdff dff_B_4HVlGHnt6_2(.din(w_dff_B_T7akaYFz9_2),.dout(w_dff_B_4HVlGHnt6_2),.clk(gclk));
	jdff dff_B_IfJ7XFg28_2(.din(w_dff_B_4HVlGHnt6_2),.dout(w_dff_B_IfJ7XFg28_2),.clk(gclk));
	jdff dff_B_YFvkUf2B4_2(.din(w_dff_B_IfJ7XFg28_2),.dout(w_dff_B_YFvkUf2B4_2),.clk(gclk));
	jdff dff_B_vQSkTbsO0_2(.din(w_dff_B_YFvkUf2B4_2),.dout(w_dff_B_vQSkTbsO0_2),.clk(gclk));
	jdff dff_B_gOonVgmw2_2(.din(w_dff_B_vQSkTbsO0_2),.dout(w_dff_B_gOonVgmw2_2),.clk(gclk));
	jdff dff_B_DlfQu4jH3_2(.din(w_dff_B_gOonVgmw2_2),.dout(w_dff_B_DlfQu4jH3_2),.clk(gclk));
	jdff dff_B_jQbxvzmW2_2(.din(n309),.dout(w_dff_B_jQbxvzmW2_2),.clk(gclk));
	jdff dff_B_genMed2k6_1(.din(n275),.dout(w_dff_B_genMed2k6_1),.clk(gclk));
	jdff dff_B_euvDCGwU1_2(.din(n225),.dout(w_dff_B_euvDCGwU1_2),.clk(gclk));
	jdff dff_B_jm1HdqEf7_2(.din(w_dff_B_euvDCGwU1_2),.dout(w_dff_B_jm1HdqEf7_2),.clk(gclk));
	jdff dff_B_PvityzRU3_2(.din(w_dff_B_jm1HdqEf7_2),.dout(w_dff_B_PvityzRU3_2),.clk(gclk));
	jdff dff_B_fbqMY5Fy7_2(.din(w_dff_B_PvityzRU3_2),.dout(w_dff_B_fbqMY5Fy7_2),.clk(gclk));
	jdff dff_B_XlrAH4nN9_2(.din(w_dff_B_fbqMY5Fy7_2),.dout(w_dff_B_XlrAH4nN9_2),.clk(gclk));
	jdff dff_B_VDOgafZk5_2(.din(w_dff_B_XlrAH4nN9_2),.dout(w_dff_B_VDOgafZk5_2),.clk(gclk));
	jdff dff_B_yIxQC1JB1_2(.din(w_dff_B_VDOgafZk5_2),.dout(w_dff_B_yIxQC1JB1_2),.clk(gclk));
	jdff dff_B_R9KdxMF81_2(.din(w_dff_B_yIxQC1JB1_2),.dout(w_dff_B_R9KdxMF81_2),.clk(gclk));
	jdff dff_B_PFtbiEVC2_2(.din(w_dff_B_R9KdxMF81_2),.dout(w_dff_B_PFtbiEVC2_2),.clk(gclk));
	jdff dff_B_qmSAHCoo1_2(.din(w_dff_B_PFtbiEVC2_2),.dout(w_dff_B_qmSAHCoo1_2),.clk(gclk));
	jdff dff_B_YeWPrfTF1_2(.din(w_dff_B_qmSAHCoo1_2),.dout(w_dff_B_YeWPrfTF1_2),.clk(gclk));
	jdff dff_B_4w5HXiWm6_2(.din(w_dff_B_YeWPrfTF1_2),.dout(w_dff_B_4w5HXiWm6_2),.clk(gclk));
	jdff dff_B_tnSzTt9L3_2(.din(n253),.dout(w_dff_B_tnSzTt9L3_2),.clk(gclk));
	jdff dff_B_wrVJX94M6_1(.din(n226),.dout(w_dff_B_wrVJX94M6_1),.clk(gclk));
	jdff dff_B_895YVFTo0_2(.din(n183),.dout(w_dff_B_895YVFTo0_2),.clk(gclk));
	jdff dff_B_4s2w8K9Y7_2(.din(w_dff_B_895YVFTo0_2),.dout(w_dff_B_4s2w8K9Y7_2),.clk(gclk));
	jdff dff_B_ZI8ipCT06_2(.din(w_dff_B_4s2w8K9Y7_2),.dout(w_dff_B_ZI8ipCT06_2),.clk(gclk));
	jdff dff_B_bX9VQi0l8_2(.din(w_dff_B_ZI8ipCT06_2),.dout(w_dff_B_bX9VQi0l8_2),.clk(gclk));
	jdff dff_B_3eTLC9ts9_2(.din(w_dff_B_bX9VQi0l8_2),.dout(w_dff_B_3eTLC9ts9_2),.clk(gclk));
	jdff dff_B_042cQft63_2(.din(w_dff_B_3eTLC9ts9_2),.dout(w_dff_B_042cQft63_2),.clk(gclk));
	jdff dff_B_Acj0Q3uf9_2(.din(w_dff_B_042cQft63_2),.dout(w_dff_B_Acj0Q3uf9_2),.clk(gclk));
	jdff dff_B_Hotdf22T6_2(.din(w_dff_B_Acj0Q3uf9_2),.dout(w_dff_B_Hotdf22T6_2),.clk(gclk));
	jdff dff_B_e4Sw9TXZ8_2(.din(w_dff_B_Hotdf22T6_2),.dout(w_dff_B_e4Sw9TXZ8_2),.clk(gclk));
	jdff dff_B_ezZqCDx86_2(.din(n204),.dout(w_dff_B_ezZqCDx86_2),.clk(gclk));
	jdff dff_B_APnmgULd0_1(.din(n184),.dout(w_dff_B_APnmgULd0_1),.clk(gclk));
	jdff dff_B_4chyMujv4_2(.din(n148),.dout(w_dff_B_4chyMujv4_2),.clk(gclk));
	jdff dff_B_OyqFo2pv3_2(.din(w_dff_B_4chyMujv4_2),.dout(w_dff_B_OyqFo2pv3_2),.clk(gclk));
	jdff dff_B_YlC1PFSL0_2(.din(w_dff_B_OyqFo2pv3_2),.dout(w_dff_B_YlC1PFSL0_2),.clk(gclk));
	jdff dff_B_hgHBTYbN4_2(.din(w_dff_B_YlC1PFSL0_2),.dout(w_dff_B_hgHBTYbN4_2),.clk(gclk));
	jdff dff_B_RwhEWNGK6_2(.din(w_dff_B_hgHBTYbN4_2),.dout(w_dff_B_RwhEWNGK6_2),.clk(gclk));
	jdff dff_B_NaR232Rg3_2(.din(w_dff_B_RwhEWNGK6_2),.dout(w_dff_B_NaR232Rg3_2),.clk(gclk));
	jdff dff_B_Z5Otzmzb1_2(.din(n162),.dout(w_dff_B_Z5Otzmzb1_2),.clk(gclk));
	jdff dff_B_577uiCVg7_2(.din(n119),.dout(w_dff_B_577uiCVg7_2),.clk(gclk));
	jdff dff_B_sx2C9rLO4_2(.din(w_dff_B_577uiCVg7_2),.dout(w_dff_B_sx2C9rLO4_2),.clk(gclk));
	jdff dff_B_O43b9nPM6_2(.din(w_dff_B_sx2C9rLO4_2),.dout(w_dff_B_O43b9nPM6_2),.clk(gclk));
	jdff dff_B_dzB81Hgh7_0(.din(n126),.dout(w_dff_B_dzB81Hgh7_0),.clk(gclk));
	jdff dff_B_LoIPBci80_0(.din(n1298),.dout(w_dff_B_LoIPBci80_0),.clk(gclk));
	jdff dff_A_qpxHJBxk7_1(.dout(w_n1294_0[1]),.din(w_dff_A_qpxHJBxk7_1),.clk(gclk));
	jdff dff_A_2JNqYLSr2_1(.dout(w_dff_A_qpxHJBxk7_1),.din(w_dff_A_2JNqYLSr2_1),.clk(gclk));
	jdff dff_B_1fupoCDN4_1(.din(n1214),.dout(w_dff_B_1fupoCDN4_1),.clk(gclk));
	jdff dff_B_bDw6z2Oz2_1(.din(w_dff_B_1fupoCDN4_1),.dout(w_dff_B_bDw6z2Oz2_1),.clk(gclk));
	jdff dff_B_agULwE7d2_2(.din(n1120),.dout(w_dff_B_agULwE7d2_2),.clk(gclk));
	jdff dff_B_9G69aGdd5_2(.din(w_dff_B_agULwE7d2_2),.dout(w_dff_B_9G69aGdd5_2),.clk(gclk));
	jdff dff_B_tKOA0cNV7_2(.din(w_dff_B_9G69aGdd5_2),.dout(w_dff_B_tKOA0cNV7_2),.clk(gclk));
	jdff dff_B_I8NQoZMb0_2(.din(w_dff_B_tKOA0cNV7_2),.dout(w_dff_B_I8NQoZMb0_2),.clk(gclk));
	jdff dff_B_3d7BK34F9_2(.din(w_dff_B_I8NQoZMb0_2),.dout(w_dff_B_3d7BK34F9_2),.clk(gclk));
	jdff dff_B_Z7r1eV5q3_2(.din(w_dff_B_3d7BK34F9_2),.dout(w_dff_B_Z7r1eV5q3_2),.clk(gclk));
	jdff dff_B_0Lb0Z4XO1_2(.din(w_dff_B_Z7r1eV5q3_2),.dout(w_dff_B_0Lb0Z4XO1_2),.clk(gclk));
	jdff dff_B_nQFnVsln3_2(.din(w_dff_B_0Lb0Z4XO1_2),.dout(w_dff_B_nQFnVsln3_2),.clk(gclk));
	jdff dff_B_Kb7Zeb3Y6_2(.din(w_dff_B_nQFnVsln3_2),.dout(w_dff_B_Kb7Zeb3Y6_2),.clk(gclk));
	jdff dff_B_2X3IdqpE8_2(.din(w_dff_B_Kb7Zeb3Y6_2),.dout(w_dff_B_2X3IdqpE8_2),.clk(gclk));
	jdff dff_B_AM3Gsmgg2_2(.din(w_dff_B_2X3IdqpE8_2),.dout(w_dff_B_AM3Gsmgg2_2),.clk(gclk));
	jdff dff_B_js2o9Z0f2_2(.din(w_dff_B_AM3Gsmgg2_2),.dout(w_dff_B_js2o9Z0f2_2),.clk(gclk));
	jdff dff_B_jABkcMLU9_2(.din(w_dff_B_js2o9Z0f2_2),.dout(w_dff_B_jABkcMLU9_2),.clk(gclk));
	jdff dff_B_GEq0rs3t1_2(.din(w_dff_B_jABkcMLU9_2),.dout(w_dff_B_GEq0rs3t1_2),.clk(gclk));
	jdff dff_B_z3jHJwCv0_2(.din(w_dff_B_GEq0rs3t1_2),.dout(w_dff_B_z3jHJwCv0_2),.clk(gclk));
	jdff dff_B_OsDbvXug6_2(.din(w_dff_B_z3jHJwCv0_2),.dout(w_dff_B_OsDbvXug6_2),.clk(gclk));
	jdff dff_B_yCyNaL3H4_2(.din(w_dff_B_OsDbvXug6_2),.dout(w_dff_B_yCyNaL3H4_2),.clk(gclk));
	jdff dff_B_qc7t4wag4_2(.din(w_dff_B_yCyNaL3H4_2),.dout(w_dff_B_qc7t4wag4_2),.clk(gclk));
	jdff dff_B_zNShhUgA5_2(.din(w_dff_B_qc7t4wag4_2),.dout(w_dff_B_zNShhUgA5_2),.clk(gclk));
	jdff dff_B_ZfHSKcpl7_2(.din(w_dff_B_zNShhUgA5_2),.dout(w_dff_B_ZfHSKcpl7_2),.clk(gclk));
	jdff dff_B_4nWPXNbs0_2(.din(w_dff_B_ZfHSKcpl7_2),.dout(w_dff_B_4nWPXNbs0_2),.clk(gclk));
	jdff dff_B_p2gXxWfN5_2(.din(w_dff_B_4nWPXNbs0_2),.dout(w_dff_B_p2gXxWfN5_2),.clk(gclk));
	jdff dff_B_zJyTFgA67_2(.din(w_dff_B_p2gXxWfN5_2),.dout(w_dff_B_zJyTFgA67_2),.clk(gclk));
	jdff dff_B_rz3cbqO80_2(.din(w_dff_B_zJyTFgA67_2),.dout(w_dff_B_rz3cbqO80_2),.clk(gclk));
	jdff dff_B_6zMnba1y1_2(.din(w_dff_B_rz3cbqO80_2),.dout(w_dff_B_6zMnba1y1_2),.clk(gclk));
	jdff dff_B_79eag0Im4_2(.din(w_dff_B_6zMnba1y1_2),.dout(w_dff_B_79eag0Im4_2),.clk(gclk));
	jdff dff_B_s7YJnI191_2(.din(w_dff_B_79eag0Im4_2),.dout(w_dff_B_s7YJnI191_2),.clk(gclk));
	jdff dff_B_QQAIagTG4_2(.din(w_dff_B_s7YJnI191_2),.dout(w_dff_B_QQAIagTG4_2),.clk(gclk));
	jdff dff_B_1lIRuHz28_2(.din(w_dff_B_QQAIagTG4_2),.dout(w_dff_B_1lIRuHz28_2),.clk(gclk));
	jdff dff_B_IidVnOHl6_2(.din(w_dff_B_1lIRuHz28_2),.dout(w_dff_B_IidVnOHl6_2),.clk(gclk));
	jdff dff_B_Tp1iF3st0_2(.din(w_dff_B_IidVnOHl6_2),.dout(w_dff_B_Tp1iF3st0_2),.clk(gclk));
	jdff dff_B_WkK6Jg3g3_2(.din(w_dff_B_Tp1iF3st0_2),.dout(w_dff_B_WkK6Jg3g3_2),.clk(gclk));
	jdff dff_B_lH4z1VnS0_2(.din(w_dff_B_WkK6Jg3g3_2),.dout(w_dff_B_lH4z1VnS0_2),.clk(gclk));
	jdff dff_B_rEbARcMs4_2(.din(w_dff_B_lH4z1VnS0_2),.dout(w_dff_B_rEbARcMs4_2),.clk(gclk));
	jdff dff_B_g7WqY3Vk1_2(.din(w_dff_B_rEbARcMs4_2),.dout(w_dff_B_g7WqY3Vk1_2),.clk(gclk));
	jdff dff_B_NUMWLlKW5_2(.din(w_dff_B_g7WqY3Vk1_2),.dout(w_dff_B_NUMWLlKW5_2),.clk(gclk));
	jdff dff_B_JrUy5QGY1_2(.din(w_dff_B_NUMWLlKW5_2),.dout(w_dff_B_JrUy5QGY1_2),.clk(gclk));
	jdff dff_B_aPPa0fvm0_2(.din(w_dff_B_JrUy5QGY1_2),.dout(w_dff_B_aPPa0fvm0_2),.clk(gclk));
	jdff dff_B_7H0YXTN93_2(.din(w_dff_B_aPPa0fvm0_2),.dout(w_dff_B_7H0YXTN93_2),.clk(gclk));
	jdff dff_B_1nH08Sja8_2(.din(w_dff_B_7H0YXTN93_2),.dout(w_dff_B_1nH08Sja8_2),.clk(gclk));
	jdff dff_B_XG3sNIfl3_2(.din(w_dff_B_1nH08Sja8_2),.dout(w_dff_B_XG3sNIfl3_2),.clk(gclk));
	jdff dff_B_yXpJVcTT4_2(.din(w_dff_B_XG3sNIfl3_2),.dout(w_dff_B_yXpJVcTT4_2),.clk(gclk));
	jdff dff_B_R2JGXC7W8_2(.din(w_dff_B_yXpJVcTT4_2),.dout(w_dff_B_R2JGXC7W8_2),.clk(gclk));
	jdff dff_B_Yl0vInWa3_2(.din(w_dff_B_R2JGXC7W8_2),.dout(w_dff_B_Yl0vInWa3_2),.clk(gclk));
	jdff dff_B_wGGF3adj5_2(.din(w_dff_B_Yl0vInWa3_2),.dout(w_dff_B_wGGF3adj5_2),.clk(gclk));
	jdff dff_B_cdwtbpXo2_2(.din(n1203),.dout(w_dff_B_cdwtbpXo2_2),.clk(gclk));
	jdff dff_B_DqGxwHbC1_1(.din(n1122),.dout(w_dff_B_DqGxwHbC1_1),.clk(gclk));
	jdff dff_B_VV78izEa9_2(.din(n1023),.dout(w_dff_B_VV78izEa9_2),.clk(gclk));
	jdff dff_B_JMfHh7yQ0_2(.din(w_dff_B_VV78izEa9_2),.dout(w_dff_B_JMfHh7yQ0_2),.clk(gclk));
	jdff dff_B_ZYCJzGjH1_2(.din(w_dff_B_JMfHh7yQ0_2),.dout(w_dff_B_ZYCJzGjH1_2),.clk(gclk));
	jdff dff_B_wf8qKgqo5_2(.din(w_dff_B_ZYCJzGjH1_2),.dout(w_dff_B_wf8qKgqo5_2),.clk(gclk));
	jdff dff_B_Ob14SXDA6_2(.din(w_dff_B_wf8qKgqo5_2),.dout(w_dff_B_Ob14SXDA6_2),.clk(gclk));
	jdff dff_B_H8wrZPF16_2(.din(w_dff_B_Ob14SXDA6_2),.dout(w_dff_B_H8wrZPF16_2),.clk(gclk));
	jdff dff_B_t6MrAjES9_2(.din(w_dff_B_H8wrZPF16_2),.dout(w_dff_B_t6MrAjES9_2),.clk(gclk));
	jdff dff_B_XnWuqa858_2(.din(w_dff_B_t6MrAjES9_2),.dout(w_dff_B_XnWuqa858_2),.clk(gclk));
	jdff dff_B_kZDBTZal0_2(.din(w_dff_B_XnWuqa858_2),.dout(w_dff_B_kZDBTZal0_2),.clk(gclk));
	jdff dff_B_6yvoHXFB8_2(.din(w_dff_B_kZDBTZal0_2),.dout(w_dff_B_6yvoHXFB8_2),.clk(gclk));
	jdff dff_B_kmO6vQG50_2(.din(w_dff_B_6yvoHXFB8_2),.dout(w_dff_B_kmO6vQG50_2),.clk(gclk));
	jdff dff_B_4k5jc4My3_2(.din(w_dff_B_kmO6vQG50_2),.dout(w_dff_B_4k5jc4My3_2),.clk(gclk));
	jdff dff_B_vr977IGf2_2(.din(w_dff_B_4k5jc4My3_2),.dout(w_dff_B_vr977IGf2_2),.clk(gclk));
	jdff dff_B_nSYaRnhO1_2(.din(w_dff_B_vr977IGf2_2),.dout(w_dff_B_nSYaRnhO1_2),.clk(gclk));
	jdff dff_B_vJ78mm8x6_2(.din(w_dff_B_nSYaRnhO1_2),.dout(w_dff_B_vJ78mm8x6_2),.clk(gclk));
	jdff dff_B_RyP6E7gn7_2(.din(w_dff_B_vJ78mm8x6_2),.dout(w_dff_B_RyP6E7gn7_2),.clk(gclk));
	jdff dff_B_Myshnbe47_2(.din(w_dff_B_RyP6E7gn7_2),.dout(w_dff_B_Myshnbe47_2),.clk(gclk));
	jdff dff_B_qKkLw8Kc0_2(.din(w_dff_B_Myshnbe47_2),.dout(w_dff_B_qKkLw8Kc0_2),.clk(gclk));
	jdff dff_B_IisZFHk28_2(.din(w_dff_B_qKkLw8Kc0_2),.dout(w_dff_B_IisZFHk28_2),.clk(gclk));
	jdff dff_B_173zE3wI9_2(.din(w_dff_B_IisZFHk28_2),.dout(w_dff_B_173zE3wI9_2),.clk(gclk));
	jdff dff_B_iRmfp9v25_2(.din(w_dff_B_173zE3wI9_2),.dout(w_dff_B_iRmfp9v25_2),.clk(gclk));
	jdff dff_B_Q9WrxAtQ0_2(.din(w_dff_B_iRmfp9v25_2),.dout(w_dff_B_Q9WrxAtQ0_2),.clk(gclk));
	jdff dff_B_IneNu71y8_2(.din(w_dff_B_Q9WrxAtQ0_2),.dout(w_dff_B_IneNu71y8_2),.clk(gclk));
	jdff dff_B_u2K4lrpV7_2(.din(w_dff_B_IneNu71y8_2),.dout(w_dff_B_u2K4lrpV7_2),.clk(gclk));
	jdff dff_B_gfMryNpa4_2(.din(w_dff_B_u2K4lrpV7_2),.dout(w_dff_B_gfMryNpa4_2),.clk(gclk));
	jdff dff_B_fRjP8YWz6_2(.din(w_dff_B_gfMryNpa4_2),.dout(w_dff_B_fRjP8YWz6_2),.clk(gclk));
	jdff dff_B_D5pOJyV48_2(.din(w_dff_B_fRjP8YWz6_2),.dout(w_dff_B_D5pOJyV48_2),.clk(gclk));
	jdff dff_B_lrRpCMSJ2_2(.din(w_dff_B_D5pOJyV48_2),.dout(w_dff_B_lrRpCMSJ2_2),.clk(gclk));
	jdff dff_B_Xvy2Y6VW9_2(.din(w_dff_B_lrRpCMSJ2_2),.dout(w_dff_B_Xvy2Y6VW9_2),.clk(gclk));
	jdff dff_B_kapuTbQO3_2(.din(w_dff_B_Xvy2Y6VW9_2),.dout(w_dff_B_kapuTbQO3_2),.clk(gclk));
	jdff dff_B_XGW6OSEY6_2(.din(w_dff_B_kapuTbQO3_2),.dout(w_dff_B_XGW6OSEY6_2),.clk(gclk));
	jdff dff_B_vCc9X8W45_2(.din(w_dff_B_XGW6OSEY6_2),.dout(w_dff_B_vCc9X8W45_2),.clk(gclk));
	jdff dff_B_it0Mh74z4_2(.din(w_dff_B_vCc9X8W45_2),.dout(w_dff_B_it0Mh74z4_2),.clk(gclk));
	jdff dff_B_hFTNOiXp8_2(.din(w_dff_B_it0Mh74z4_2),.dout(w_dff_B_hFTNOiXp8_2),.clk(gclk));
	jdff dff_B_r37wjaCq0_2(.din(w_dff_B_hFTNOiXp8_2),.dout(w_dff_B_r37wjaCq0_2),.clk(gclk));
	jdff dff_B_xdNBrZCi3_2(.din(w_dff_B_r37wjaCq0_2),.dout(w_dff_B_xdNBrZCi3_2),.clk(gclk));
	jdff dff_B_hbOlwcAs2_2(.din(w_dff_B_xdNBrZCi3_2),.dout(w_dff_B_hbOlwcAs2_2),.clk(gclk));
	jdff dff_B_czKOHofc8_2(.din(w_dff_B_hbOlwcAs2_2),.dout(w_dff_B_czKOHofc8_2),.clk(gclk));
	jdff dff_B_ygtjzrFC1_2(.din(w_dff_B_czKOHofc8_2),.dout(w_dff_B_ygtjzrFC1_2),.clk(gclk));
	jdff dff_B_QYiA9Km83_2(.din(w_dff_B_ygtjzrFC1_2),.dout(w_dff_B_QYiA9Km83_2),.clk(gclk));
	jdff dff_B_73M7BQO13_2(.din(w_dff_B_QYiA9Km83_2),.dout(w_dff_B_73M7BQO13_2),.clk(gclk));
	jdff dff_B_falzzeP72_2(.din(n1103),.dout(w_dff_B_falzzeP72_2),.clk(gclk));
	jdff dff_B_hUWPJ5Ia0_1(.din(n1024),.dout(w_dff_B_hUWPJ5Ia0_1),.clk(gclk));
	jdff dff_B_38pXlEXW0_2(.din(n924),.dout(w_dff_B_38pXlEXW0_2),.clk(gclk));
	jdff dff_B_Crpe4JDv4_2(.din(w_dff_B_38pXlEXW0_2),.dout(w_dff_B_Crpe4JDv4_2),.clk(gclk));
	jdff dff_B_97xQvbry6_2(.din(w_dff_B_Crpe4JDv4_2),.dout(w_dff_B_97xQvbry6_2),.clk(gclk));
	jdff dff_B_mrqPKc1Z9_2(.din(w_dff_B_97xQvbry6_2),.dout(w_dff_B_mrqPKc1Z9_2),.clk(gclk));
	jdff dff_B_jt0FEUrP4_2(.din(w_dff_B_mrqPKc1Z9_2),.dout(w_dff_B_jt0FEUrP4_2),.clk(gclk));
	jdff dff_B_mGJMO9eB6_2(.din(w_dff_B_jt0FEUrP4_2),.dout(w_dff_B_mGJMO9eB6_2),.clk(gclk));
	jdff dff_B_RT6MvAg04_2(.din(w_dff_B_mGJMO9eB6_2),.dout(w_dff_B_RT6MvAg04_2),.clk(gclk));
	jdff dff_B_1LtO1l2e5_2(.din(w_dff_B_RT6MvAg04_2),.dout(w_dff_B_1LtO1l2e5_2),.clk(gclk));
	jdff dff_B_Q2eDYiTU0_2(.din(w_dff_B_1LtO1l2e5_2),.dout(w_dff_B_Q2eDYiTU0_2),.clk(gclk));
	jdff dff_B_ezHkWKvm5_2(.din(w_dff_B_Q2eDYiTU0_2),.dout(w_dff_B_ezHkWKvm5_2),.clk(gclk));
	jdff dff_B_M6PcMdri6_2(.din(w_dff_B_ezHkWKvm5_2),.dout(w_dff_B_M6PcMdri6_2),.clk(gclk));
	jdff dff_B_P3VgKcs09_2(.din(w_dff_B_M6PcMdri6_2),.dout(w_dff_B_P3VgKcs09_2),.clk(gclk));
	jdff dff_B_yBk1mHDO0_2(.din(w_dff_B_P3VgKcs09_2),.dout(w_dff_B_yBk1mHDO0_2),.clk(gclk));
	jdff dff_B_BlxQOUZS7_2(.din(w_dff_B_yBk1mHDO0_2),.dout(w_dff_B_BlxQOUZS7_2),.clk(gclk));
	jdff dff_B_ltFOv6Vo1_2(.din(w_dff_B_BlxQOUZS7_2),.dout(w_dff_B_ltFOv6Vo1_2),.clk(gclk));
	jdff dff_B_4J8Yf2W26_2(.din(w_dff_B_ltFOv6Vo1_2),.dout(w_dff_B_4J8Yf2W26_2),.clk(gclk));
	jdff dff_B_BYr64GK65_2(.din(w_dff_B_4J8Yf2W26_2),.dout(w_dff_B_BYr64GK65_2),.clk(gclk));
	jdff dff_B_8rB9nKcx1_2(.din(w_dff_B_BYr64GK65_2),.dout(w_dff_B_8rB9nKcx1_2),.clk(gclk));
	jdff dff_B_wqUHvkBj8_2(.din(w_dff_B_8rB9nKcx1_2),.dout(w_dff_B_wqUHvkBj8_2),.clk(gclk));
	jdff dff_B_ywuXpUg47_2(.din(w_dff_B_wqUHvkBj8_2),.dout(w_dff_B_ywuXpUg47_2),.clk(gclk));
	jdff dff_B_8gURS7ci2_2(.din(w_dff_B_ywuXpUg47_2),.dout(w_dff_B_8gURS7ci2_2),.clk(gclk));
	jdff dff_B_7jpLkQnA1_2(.din(w_dff_B_8gURS7ci2_2),.dout(w_dff_B_7jpLkQnA1_2),.clk(gclk));
	jdff dff_B_ZxD3NAAN4_2(.din(w_dff_B_7jpLkQnA1_2),.dout(w_dff_B_ZxD3NAAN4_2),.clk(gclk));
	jdff dff_B_V06AWYwM1_2(.din(w_dff_B_ZxD3NAAN4_2),.dout(w_dff_B_V06AWYwM1_2),.clk(gclk));
	jdff dff_B_9SUaudRb2_2(.din(w_dff_B_V06AWYwM1_2),.dout(w_dff_B_9SUaudRb2_2),.clk(gclk));
	jdff dff_B_VrWv7SJo9_2(.din(w_dff_B_9SUaudRb2_2),.dout(w_dff_B_VrWv7SJo9_2),.clk(gclk));
	jdff dff_B_Apnxg2Su3_2(.din(w_dff_B_VrWv7SJo9_2),.dout(w_dff_B_Apnxg2Su3_2),.clk(gclk));
	jdff dff_B_a4hT12As6_2(.din(w_dff_B_Apnxg2Su3_2),.dout(w_dff_B_a4hT12As6_2),.clk(gclk));
	jdff dff_B_iJMMg6Ci0_2(.din(w_dff_B_a4hT12As6_2),.dout(w_dff_B_iJMMg6Ci0_2),.clk(gclk));
	jdff dff_B_udsFMJq63_2(.din(w_dff_B_iJMMg6Ci0_2),.dout(w_dff_B_udsFMJq63_2),.clk(gclk));
	jdff dff_B_nh31iq2e9_2(.din(w_dff_B_udsFMJq63_2),.dout(w_dff_B_nh31iq2e9_2),.clk(gclk));
	jdff dff_B_3OVzZOA39_2(.din(w_dff_B_nh31iq2e9_2),.dout(w_dff_B_3OVzZOA39_2),.clk(gclk));
	jdff dff_B_HTKKiomk7_2(.din(w_dff_B_3OVzZOA39_2),.dout(w_dff_B_HTKKiomk7_2),.clk(gclk));
	jdff dff_B_35qTgeS53_2(.din(w_dff_B_HTKKiomk7_2),.dout(w_dff_B_35qTgeS53_2),.clk(gclk));
	jdff dff_B_Zn1pUUIV4_2(.din(w_dff_B_35qTgeS53_2),.dout(w_dff_B_Zn1pUUIV4_2),.clk(gclk));
	jdff dff_B_TERMiXSN4_2(.din(w_dff_B_Zn1pUUIV4_2),.dout(w_dff_B_TERMiXSN4_2),.clk(gclk));
	jdff dff_B_0s0TzxQu7_2(.din(n1004),.dout(w_dff_B_0s0TzxQu7_2),.clk(gclk));
	jdff dff_B_kcbxlRjy9_1(.din(n925),.dout(w_dff_B_kcbxlRjy9_1),.clk(gclk));
	jdff dff_B_sXUB0K114_2(.din(n822),.dout(w_dff_B_sXUB0K114_2),.clk(gclk));
	jdff dff_B_YYgudbEX2_2(.din(w_dff_B_sXUB0K114_2),.dout(w_dff_B_YYgudbEX2_2),.clk(gclk));
	jdff dff_B_vJXMOotG0_2(.din(w_dff_B_YYgudbEX2_2),.dout(w_dff_B_vJXMOotG0_2),.clk(gclk));
	jdff dff_B_NTZ2dVIL2_2(.din(w_dff_B_vJXMOotG0_2),.dout(w_dff_B_NTZ2dVIL2_2),.clk(gclk));
	jdff dff_B_X4nHCl4w9_2(.din(w_dff_B_NTZ2dVIL2_2),.dout(w_dff_B_X4nHCl4w9_2),.clk(gclk));
	jdff dff_B_gAE62IgG1_2(.din(w_dff_B_X4nHCl4w9_2),.dout(w_dff_B_gAE62IgG1_2),.clk(gclk));
	jdff dff_B_aQZGDkUz8_2(.din(w_dff_B_gAE62IgG1_2),.dout(w_dff_B_aQZGDkUz8_2),.clk(gclk));
	jdff dff_B_onVMGKRj3_2(.din(w_dff_B_aQZGDkUz8_2),.dout(w_dff_B_onVMGKRj3_2),.clk(gclk));
	jdff dff_B_FgjOxEOF1_2(.din(w_dff_B_onVMGKRj3_2),.dout(w_dff_B_FgjOxEOF1_2),.clk(gclk));
	jdff dff_B_bfyIWMSJ1_2(.din(w_dff_B_FgjOxEOF1_2),.dout(w_dff_B_bfyIWMSJ1_2),.clk(gclk));
	jdff dff_B_xDZnBuEW5_2(.din(w_dff_B_bfyIWMSJ1_2),.dout(w_dff_B_xDZnBuEW5_2),.clk(gclk));
	jdff dff_B_GErPVUKH1_2(.din(w_dff_B_xDZnBuEW5_2),.dout(w_dff_B_GErPVUKH1_2),.clk(gclk));
	jdff dff_B_Gd7Hg6vj8_2(.din(w_dff_B_GErPVUKH1_2),.dout(w_dff_B_Gd7Hg6vj8_2),.clk(gclk));
	jdff dff_B_pMVFnvOx5_2(.din(w_dff_B_Gd7Hg6vj8_2),.dout(w_dff_B_pMVFnvOx5_2),.clk(gclk));
	jdff dff_B_AehMOhl39_2(.din(w_dff_B_pMVFnvOx5_2),.dout(w_dff_B_AehMOhl39_2),.clk(gclk));
	jdff dff_B_TpH9i84D8_2(.din(w_dff_B_AehMOhl39_2),.dout(w_dff_B_TpH9i84D8_2),.clk(gclk));
	jdff dff_B_AQPdMPZB4_2(.din(w_dff_B_TpH9i84D8_2),.dout(w_dff_B_AQPdMPZB4_2),.clk(gclk));
	jdff dff_B_GU4ROdY50_2(.din(w_dff_B_AQPdMPZB4_2),.dout(w_dff_B_GU4ROdY50_2),.clk(gclk));
	jdff dff_B_hoyULrMt1_2(.din(w_dff_B_GU4ROdY50_2),.dout(w_dff_B_hoyULrMt1_2),.clk(gclk));
	jdff dff_B_REC2RIuZ3_2(.din(w_dff_B_hoyULrMt1_2),.dout(w_dff_B_REC2RIuZ3_2),.clk(gclk));
	jdff dff_B_3WRI4TEW0_2(.din(w_dff_B_REC2RIuZ3_2),.dout(w_dff_B_3WRI4TEW0_2),.clk(gclk));
	jdff dff_B_AOovrG2I8_2(.din(w_dff_B_3WRI4TEW0_2),.dout(w_dff_B_AOovrG2I8_2),.clk(gclk));
	jdff dff_B_iVdF1zSj9_2(.din(w_dff_B_AOovrG2I8_2),.dout(w_dff_B_iVdF1zSj9_2),.clk(gclk));
	jdff dff_B_CSJejrr00_2(.din(w_dff_B_iVdF1zSj9_2),.dout(w_dff_B_CSJejrr00_2),.clk(gclk));
	jdff dff_B_TmgQY7aq7_2(.din(w_dff_B_CSJejrr00_2),.dout(w_dff_B_TmgQY7aq7_2),.clk(gclk));
	jdff dff_B_h0FRUO3j1_2(.din(w_dff_B_TmgQY7aq7_2),.dout(w_dff_B_h0FRUO3j1_2),.clk(gclk));
	jdff dff_B_cxljlFJk5_2(.din(w_dff_B_h0FRUO3j1_2),.dout(w_dff_B_cxljlFJk5_2),.clk(gclk));
	jdff dff_B_YT0MdckA4_2(.din(w_dff_B_cxljlFJk5_2),.dout(w_dff_B_YT0MdckA4_2),.clk(gclk));
	jdff dff_B_G4X87IfJ0_2(.din(w_dff_B_YT0MdckA4_2),.dout(w_dff_B_G4X87IfJ0_2),.clk(gclk));
	jdff dff_B_CXA7bD8E7_2(.din(w_dff_B_G4X87IfJ0_2),.dout(w_dff_B_CXA7bD8E7_2),.clk(gclk));
	jdff dff_B_Kr04a6zH7_2(.din(w_dff_B_CXA7bD8E7_2),.dout(w_dff_B_Kr04a6zH7_2),.clk(gclk));
	jdff dff_B_wiemeGC85_2(.din(w_dff_B_Kr04a6zH7_2),.dout(w_dff_B_wiemeGC85_2),.clk(gclk));
	jdff dff_B_6PAvUIMV1_2(.din(w_dff_B_wiemeGC85_2),.dout(w_dff_B_6PAvUIMV1_2),.clk(gclk));
	jdff dff_B_2oTC1IeI8_2(.din(n898),.dout(w_dff_B_2oTC1IeI8_2),.clk(gclk));
	jdff dff_B_ga3xMME42_1(.din(n823),.dout(w_dff_B_ga3xMME42_1),.clk(gclk));
	jdff dff_B_vTMbvAtu7_2(.din(n724),.dout(w_dff_B_vTMbvAtu7_2),.clk(gclk));
	jdff dff_B_G4nAPH1o3_2(.din(w_dff_B_vTMbvAtu7_2),.dout(w_dff_B_G4nAPH1o3_2),.clk(gclk));
	jdff dff_B_NnmeNfwY3_2(.din(w_dff_B_G4nAPH1o3_2),.dout(w_dff_B_NnmeNfwY3_2),.clk(gclk));
	jdff dff_B_rfwclIUl9_2(.din(w_dff_B_NnmeNfwY3_2),.dout(w_dff_B_rfwclIUl9_2),.clk(gclk));
	jdff dff_B_2qcbZqSG7_2(.din(w_dff_B_rfwclIUl9_2),.dout(w_dff_B_2qcbZqSG7_2),.clk(gclk));
	jdff dff_B_Jv9X6WHL8_2(.din(w_dff_B_2qcbZqSG7_2),.dout(w_dff_B_Jv9X6WHL8_2),.clk(gclk));
	jdff dff_B_7tMLKjnG5_2(.din(w_dff_B_Jv9X6WHL8_2),.dout(w_dff_B_7tMLKjnG5_2),.clk(gclk));
	jdff dff_B_7001iSvU5_2(.din(w_dff_B_7tMLKjnG5_2),.dout(w_dff_B_7001iSvU5_2),.clk(gclk));
	jdff dff_B_i7ycTdzN4_2(.din(w_dff_B_7001iSvU5_2),.dout(w_dff_B_i7ycTdzN4_2),.clk(gclk));
	jdff dff_B_IIDlM1ND3_2(.din(w_dff_B_i7ycTdzN4_2),.dout(w_dff_B_IIDlM1ND3_2),.clk(gclk));
	jdff dff_B_9dRHixW77_2(.din(w_dff_B_IIDlM1ND3_2),.dout(w_dff_B_9dRHixW77_2),.clk(gclk));
	jdff dff_B_PYVcYUhh0_2(.din(w_dff_B_9dRHixW77_2),.dout(w_dff_B_PYVcYUhh0_2),.clk(gclk));
	jdff dff_B_6uRsDfVo0_2(.din(w_dff_B_PYVcYUhh0_2),.dout(w_dff_B_6uRsDfVo0_2),.clk(gclk));
	jdff dff_B_bIISXcli7_2(.din(w_dff_B_6uRsDfVo0_2),.dout(w_dff_B_bIISXcli7_2),.clk(gclk));
	jdff dff_B_Et2FDZtn3_2(.din(w_dff_B_bIISXcli7_2),.dout(w_dff_B_Et2FDZtn3_2),.clk(gclk));
	jdff dff_B_8qZZ8Nt57_2(.din(w_dff_B_Et2FDZtn3_2),.dout(w_dff_B_8qZZ8Nt57_2),.clk(gclk));
	jdff dff_B_AERnxkmb3_2(.din(w_dff_B_8qZZ8Nt57_2),.dout(w_dff_B_AERnxkmb3_2),.clk(gclk));
	jdff dff_B_dpix5o353_2(.din(w_dff_B_AERnxkmb3_2),.dout(w_dff_B_dpix5o353_2),.clk(gclk));
	jdff dff_B_XSC01LDr4_2(.din(w_dff_B_dpix5o353_2),.dout(w_dff_B_XSC01LDr4_2),.clk(gclk));
	jdff dff_B_VzC8j6nj0_2(.din(w_dff_B_XSC01LDr4_2),.dout(w_dff_B_VzC8j6nj0_2),.clk(gclk));
	jdff dff_B_rXnnaJ8p2_2(.din(w_dff_B_VzC8j6nj0_2),.dout(w_dff_B_rXnnaJ8p2_2),.clk(gclk));
	jdff dff_B_99nxWuam3_2(.din(w_dff_B_rXnnaJ8p2_2),.dout(w_dff_B_99nxWuam3_2),.clk(gclk));
	jdff dff_B_7xjFRmPL5_2(.din(w_dff_B_99nxWuam3_2),.dout(w_dff_B_7xjFRmPL5_2),.clk(gclk));
	jdff dff_B_mRuCOBGJ1_2(.din(w_dff_B_7xjFRmPL5_2),.dout(w_dff_B_mRuCOBGJ1_2),.clk(gclk));
	jdff dff_B_oXeNmgWz7_2(.din(w_dff_B_mRuCOBGJ1_2),.dout(w_dff_B_oXeNmgWz7_2),.clk(gclk));
	jdff dff_B_ycWV6Zts4_2(.din(w_dff_B_oXeNmgWz7_2),.dout(w_dff_B_ycWV6Zts4_2),.clk(gclk));
	jdff dff_B_fZhepIFF1_2(.din(w_dff_B_ycWV6Zts4_2),.dout(w_dff_B_fZhepIFF1_2),.clk(gclk));
	jdff dff_B_5V2BFPIT7_2(.din(w_dff_B_fZhepIFF1_2),.dout(w_dff_B_5V2BFPIT7_2),.clk(gclk));
	jdff dff_B_MY9aCvZg6_2(.din(w_dff_B_5V2BFPIT7_2),.dout(w_dff_B_MY9aCvZg6_2),.clk(gclk));
	jdff dff_B_dn6khCWy1_2(.din(w_dff_B_MY9aCvZg6_2),.dout(w_dff_B_dn6khCWy1_2),.clk(gclk));
	jdff dff_B_kQ3pLChE1_2(.din(n795),.dout(w_dff_B_kQ3pLChE1_2),.clk(gclk));
	jdff dff_B_72vJHDRm4_1(.din(n725),.dout(w_dff_B_72vJHDRm4_1),.clk(gclk));
	jdff dff_B_WNXECbNp2_2(.din(n632),.dout(w_dff_B_WNXECbNp2_2),.clk(gclk));
	jdff dff_B_6yy8D0MW7_2(.din(w_dff_B_WNXECbNp2_2),.dout(w_dff_B_6yy8D0MW7_2),.clk(gclk));
	jdff dff_B_095mUswf9_2(.din(w_dff_B_6yy8D0MW7_2),.dout(w_dff_B_095mUswf9_2),.clk(gclk));
	jdff dff_B_ra6e7fzJ3_2(.din(w_dff_B_095mUswf9_2),.dout(w_dff_B_ra6e7fzJ3_2),.clk(gclk));
	jdff dff_B_bnGmFO3i5_2(.din(w_dff_B_ra6e7fzJ3_2),.dout(w_dff_B_bnGmFO3i5_2),.clk(gclk));
	jdff dff_B_dIlXzTbE6_2(.din(w_dff_B_bnGmFO3i5_2),.dout(w_dff_B_dIlXzTbE6_2),.clk(gclk));
	jdff dff_B_ke0Ex4BD3_2(.din(w_dff_B_dIlXzTbE6_2),.dout(w_dff_B_ke0Ex4BD3_2),.clk(gclk));
	jdff dff_B_KAHiQ5MD5_2(.din(w_dff_B_ke0Ex4BD3_2),.dout(w_dff_B_KAHiQ5MD5_2),.clk(gclk));
	jdff dff_B_bQJjeAAb6_2(.din(w_dff_B_KAHiQ5MD5_2),.dout(w_dff_B_bQJjeAAb6_2),.clk(gclk));
	jdff dff_B_S8pShqH10_2(.din(w_dff_B_bQJjeAAb6_2),.dout(w_dff_B_S8pShqH10_2),.clk(gclk));
	jdff dff_B_MxzhyBte1_2(.din(w_dff_B_S8pShqH10_2),.dout(w_dff_B_MxzhyBte1_2),.clk(gclk));
	jdff dff_B_jbY18xuA5_2(.din(w_dff_B_MxzhyBte1_2),.dout(w_dff_B_jbY18xuA5_2),.clk(gclk));
	jdff dff_B_GjZpbovM5_2(.din(w_dff_B_jbY18xuA5_2),.dout(w_dff_B_GjZpbovM5_2),.clk(gclk));
	jdff dff_B_NsfHKnrZ2_2(.din(w_dff_B_GjZpbovM5_2),.dout(w_dff_B_NsfHKnrZ2_2),.clk(gclk));
	jdff dff_B_WaTfX6FN6_2(.din(w_dff_B_NsfHKnrZ2_2),.dout(w_dff_B_WaTfX6FN6_2),.clk(gclk));
	jdff dff_B_arKz1MVK2_2(.din(w_dff_B_WaTfX6FN6_2),.dout(w_dff_B_arKz1MVK2_2),.clk(gclk));
	jdff dff_B_Ud9JqVjp2_2(.din(w_dff_B_arKz1MVK2_2),.dout(w_dff_B_Ud9JqVjp2_2),.clk(gclk));
	jdff dff_B_wf0MDSsA7_2(.din(w_dff_B_Ud9JqVjp2_2),.dout(w_dff_B_wf0MDSsA7_2),.clk(gclk));
	jdff dff_B_GvL24ZfN1_2(.din(w_dff_B_wf0MDSsA7_2),.dout(w_dff_B_GvL24ZfN1_2),.clk(gclk));
	jdff dff_B_M83a0Eab1_2(.din(w_dff_B_GvL24ZfN1_2),.dout(w_dff_B_M83a0Eab1_2),.clk(gclk));
	jdff dff_B_ME0FJdGH6_2(.din(w_dff_B_M83a0Eab1_2),.dout(w_dff_B_ME0FJdGH6_2),.clk(gclk));
	jdff dff_B_mQ5KoUqM3_2(.din(w_dff_B_ME0FJdGH6_2),.dout(w_dff_B_mQ5KoUqM3_2),.clk(gclk));
	jdff dff_B_87p6jvvS3_2(.din(w_dff_B_mQ5KoUqM3_2),.dout(w_dff_B_87p6jvvS3_2),.clk(gclk));
	jdff dff_B_0HG02Vwh6_2(.din(w_dff_B_87p6jvvS3_2),.dout(w_dff_B_0HG02Vwh6_2),.clk(gclk));
	jdff dff_B_UfNS9ONN4_2(.din(w_dff_B_0HG02Vwh6_2),.dout(w_dff_B_UfNS9ONN4_2),.clk(gclk));
	jdff dff_B_Toz374d67_2(.din(w_dff_B_UfNS9ONN4_2),.dout(w_dff_B_Toz374d67_2),.clk(gclk));
	jdff dff_B_SVn0Kq5S2_2(.din(w_dff_B_Toz374d67_2),.dout(w_dff_B_SVn0Kq5S2_2),.clk(gclk));
	jdff dff_B_QMXPycXa7_2(.din(n696),.dout(w_dff_B_QMXPycXa7_2),.clk(gclk));
	jdff dff_B_pzUmcCNM8_1(.din(n633),.dout(w_dff_B_pzUmcCNM8_1),.clk(gclk));
	jdff dff_B_C42Mg9dF7_2(.din(n547),.dout(w_dff_B_C42Mg9dF7_2),.clk(gclk));
	jdff dff_B_pVjvpTb82_2(.din(w_dff_B_C42Mg9dF7_2),.dout(w_dff_B_pVjvpTb82_2),.clk(gclk));
	jdff dff_B_QZ5Ergr54_2(.din(w_dff_B_pVjvpTb82_2),.dout(w_dff_B_QZ5Ergr54_2),.clk(gclk));
	jdff dff_B_0F1z5oQc6_2(.din(w_dff_B_QZ5Ergr54_2),.dout(w_dff_B_0F1z5oQc6_2),.clk(gclk));
	jdff dff_B_UeUDiyVH4_2(.din(w_dff_B_0F1z5oQc6_2),.dout(w_dff_B_UeUDiyVH4_2),.clk(gclk));
	jdff dff_B_LanzuH9v9_2(.din(w_dff_B_UeUDiyVH4_2),.dout(w_dff_B_LanzuH9v9_2),.clk(gclk));
	jdff dff_B_z233RMrP0_2(.din(w_dff_B_LanzuH9v9_2),.dout(w_dff_B_z233RMrP0_2),.clk(gclk));
	jdff dff_B_NqmiiqCc0_2(.din(w_dff_B_z233RMrP0_2),.dout(w_dff_B_NqmiiqCc0_2),.clk(gclk));
	jdff dff_B_FkWLYgRS5_2(.din(w_dff_B_NqmiiqCc0_2),.dout(w_dff_B_FkWLYgRS5_2),.clk(gclk));
	jdff dff_B_cGomwskl3_2(.din(w_dff_B_FkWLYgRS5_2),.dout(w_dff_B_cGomwskl3_2),.clk(gclk));
	jdff dff_B_hqs1QI3m7_2(.din(w_dff_B_cGomwskl3_2),.dout(w_dff_B_hqs1QI3m7_2),.clk(gclk));
	jdff dff_B_SMA1iwBW7_2(.din(w_dff_B_hqs1QI3m7_2),.dout(w_dff_B_SMA1iwBW7_2),.clk(gclk));
	jdff dff_B_8CGju51P5_2(.din(w_dff_B_SMA1iwBW7_2),.dout(w_dff_B_8CGju51P5_2),.clk(gclk));
	jdff dff_B_4P63Sk099_2(.din(w_dff_B_8CGju51P5_2),.dout(w_dff_B_4P63Sk099_2),.clk(gclk));
	jdff dff_B_8RovYKMb4_2(.din(w_dff_B_4P63Sk099_2),.dout(w_dff_B_8RovYKMb4_2),.clk(gclk));
	jdff dff_B_fmaC9uC59_2(.din(w_dff_B_8RovYKMb4_2),.dout(w_dff_B_fmaC9uC59_2),.clk(gclk));
	jdff dff_B_lF1rxL5v7_2(.din(w_dff_B_fmaC9uC59_2),.dout(w_dff_B_lF1rxL5v7_2),.clk(gclk));
	jdff dff_B_Cwkc5HQG3_2(.din(w_dff_B_lF1rxL5v7_2),.dout(w_dff_B_Cwkc5HQG3_2),.clk(gclk));
	jdff dff_B_aKonAQ029_2(.din(w_dff_B_Cwkc5HQG3_2),.dout(w_dff_B_aKonAQ029_2),.clk(gclk));
	jdff dff_B_qCDbyKzR8_2(.din(w_dff_B_aKonAQ029_2),.dout(w_dff_B_qCDbyKzR8_2),.clk(gclk));
	jdff dff_B_tmX8AwQQ1_2(.din(w_dff_B_qCDbyKzR8_2),.dout(w_dff_B_tmX8AwQQ1_2),.clk(gclk));
	jdff dff_B_0YCRTGia0_2(.din(w_dff_B_tmX8AwQQ1_2),.dout(w_dff_B_0YCRTGia0_2),.clk(gclk));
	jdff dff_B_dLSiwg0c4_2(.din(w_dff_B_0YCRTGia0_2),.dout(w_dff_B_dLSiwg0c4_2),.clk(gclk));
	jdff dff_B_uGOp2fnT2_2(.din(w_dff_B_dLSiwg0c4_2),.dout(w_dff_B_uGOp2fnT2_2),.clk(gclk));
	jdff dff_B_m8OWrTci8_2(.din(n604),.dout(w_dff_B_m8OWrTci8_2),.clk(gclk));
	jdff dff_B_TF5vSIb98_1(.din(n548),.dout(w_dff_B_TF5vSIb98_1),.clk(gclk));
	jdff dff_B_tQ4qXZ1x6_2(.din(n469),.dout(w_dff_B_tQ4qXZ1x6_2),.clk(gclk));
	jdff dff_B_mClwyOzS8_2(.din(w_dff_B_tQ4qXZ1x6_2),.dout(w_dff_B_mClwyOzS8_2),.clk(gclk));
	jdff dff_B_Kxlplazs1_2(.din(w_dff_B_mClwyOzS8_2),.dout(w_dff_B_Kxlplazs1_2),.clk(gclk));
	jdff dff_B_N5a60De67_2(.din(w_dff_B_Kxlplazs1_2),.dout(w_dff_B_N5a60De67_2),.clk(gclk));
	jdff dff_B_ektGJC4b7_2(.din(w_dff_B_N5a60De67_2),.dout(w_dff_B_ektGJC4b7_2),.clk(gclk));
	jdff dff_B_kUC2MXDG0_2(.din(w_dff_B_ektGJC4b7_2),.dout(w_dff_B_kUC2MXDG0_2),.clk(gclk));
	jdff dff_B_BWCi4y7u3_2(.din(w_dff_B_kUC2MXDG0_2),.dout(w_dff_B_BWCi4y7u3_2),.clk(gclk));
	jdff dff_B_yKfef8Pu0_2(.din(w_dff_B_BWCi4y7u3_2),.dout(w_dff_B_yKfef8Pu0_2),.clk(gclk));
	jdff dff_B_Fp8V6JlI0_2(.din(w_dff_B_yKfef8Pu0_2),.dout(w_dff_B_Fp8V6JlI0_2),.clk(gclk));
	jdff dff_B_DnZORb424_2(.din(w_dff_B_Fp8V6JlI0_2),.dout(w_dff_B_DnZORb424_2),.clk(gclk));
	jdff dff_B_7p2Mnrod6_2(.din(w_dff_B_DnZORb424_2),.dout(w_dff_B_7p2Mnrod6_2),.clk(gclk));
	jdff dff_B_NzmfXrmJ6_2(.din(w_dff_B_7p2Mnrod6_2),.dout(w_dff_B_NzmfXrmJ6_2),.clk(gclk));
	jdff dff_B_CkSWZqT83_2(.din(w_dff_B_NzmfXrmJ6_2),.dout(w_dff_B_CkSWZqT83_2),.clk(gclk));
	jdff dff_B_Gb3iBuFG9_2(.din(w_dff_B_CkSWZqT83_2),.dout(w_dff_B_Gb3iBuFG9_2),.clk(gclk));
	jdff dff_B_mOkqK3Gg9_2(.din(w_dff_B_Gb3iBuFG9_2),.dout(w_dff_B_mOkqK3Gg9_2),.clk(gclk));
	jdff dff_B_JWUZTMPr4_2(.din(w_dff_B_mOkqK3Gg9_2),.dout(w_dff_B_JWUZTMPr4_2),.clk(gclk));
	jdff dff_B_AyP0BeJS5_2(.din(w_dff_B_JWUZTMPr4_2),.dout(w_dff_B_AyP0BeJS5_2),.clk(gclk));
	jdff dff_B_2AWjIdOv7_2(.din(w_dff_B_AyP0BeJS5_2),.dout(w_dff_B_2AWjIdOv7_2),.clk(gclk));
	jdff dff_B_oh0qzwZ21_2(.din(w_dff_B_2AWjIdOv7_2),.dout(w_dff_B_oh0qzwZ21_2),.clk(gclk));
	jdff dff_B_2gms4NKT4_2(.din(w_dff_B_oh0qzwZ21_2),.dout(w_dff_B_2gms4NKT4_2),.clk(gclk));
	jdff dff_B_1obje77m9_2(.din(w_dff_B_2gms4NKT4_2),.dout(w_dff_B_1obje77m9_2),.clk(gclk));
	jdff dff_B_yR9CiLXM5_2(.din(n519),.dout(w_dff_B_yR9CiLXM5_2),.clk(gclk));
	jdff dff_B_dbiXsX4n4_1(.din(n470),.dout(w_dff_B_dbiXsX4n4_1),.clk(gclk));
	jdff dff_B_S6ClhJNw1_2(.din(n398),.dout(w_dff_B_S6ClhJNw1_2),.clk(gclk));
	jdff dff_B_WSKv8KBR4_2(.din(w_dff_B_S6ClhJNw1_2),.dout(w_dff_B_WSKv8KBR4_2),.clk(gclk));
	jdff dff_B_xbLX4O0F3_2(.din(w_dff_B_WSKv8KBR4_2),.dout(w_dff_B_xbLX4O0F3_2),.clk(gclk));
	jdff dff_B_S23IViRA3_2(.din(w_dff_B_xbLX4O0F3_2),.dout(w_dff_B_S23IViRA3_2),.clk(gclk));
	jdff dff_B_W2KmOD0e8_2(.din(w_dff_B_S23IViRA3_2),.dout(w_dff_B_W2KmOD0e8_2),.clk(gclk));
	jdff dff_B_8F2KyJNg0_2(.din(w_dff_B_W2KmOD0e8_2),.dout(w_dff_B_8F2KyJNg0_2),.clk(gclk));
	jdff dff_B_cCmCpYAe2_2(.din(w_dff_B_8F2KyJNg0_2),.dout(w_dff_B_cCmCpYAe2_2),.clk(gclk));
	jdff dff_B_4ViM8jpT8_2(.din(w_dff_B_cCmCpYAe2_2),.dout(w_dff_B_4ViM8jpT8_2),.clk(gclk));
	jdff dff_B_iqCsRr4K0_2(.din(w_dff_B_4ViM8jpT8_2),.dout(w_dff_B_iqCsRr4K0_2),.clk(gclk));
	jdff dff_B_b3U0LBdv4_2(.din(w_dff_B_iqCsRr4K0_2),.dout(w_dff_B_b3U0LBdv4_2),.clk(gclk));
	jdff dff_B_GxMsT4im8_2(.din(w_dff_B_b3U0LBdv4_2),.dout(w_dff_B_GxMsT4im8_2),.clk(gclk));
	jdff dff_B_esmiuX8b5_2(.din(w_dff_B_GxMsT4im8_2),.dout(w_dff_B_esmiuX8b5_2),.clk(gclk));
	jdff dff_B_3HHKbp6f0_2(.din(w_dff_B_esmiuX8b5_2),.dout(w_dff_B_3HHKbp6f0_2),.clk(gclk));
	jdff dff_B_PLmQuOCZ8_2(.din(w_dff_B_3HHKbp6f0_2),.dout(w_dff_B_PLmQuOCZ8_2),.clk(gclk));
	jdff dff_B_mkCIRXr34_2(.din(w_dff_B_PLmQuOCZ8_2),.dout(w_dff_B_mkCIRXr34_2),.clk(gclk));
	jdff dff_B_iOstxyim7_2(.din(w_dff_B_mkCIRXr34_2),.dout(w_dff_B_iOstxyim7_2),.clk(gclk));
	jdff dff_B_IV2nnOEA5_2(.din(w_dff_B_iOstxyim7_2),.dout(w_dff_B_IV2nnOEA5_2),.clk(gclk));
	jdff dff_B_0vg8Nkm94_2(.din(w_dff_B_IV2nnOEA5_2),.dout(w_dff_B_0vg8Nkm94_2),.clk(gclk));
	jdff dff_B_a3vhh17j0_2(.din(n441),.dout(w_dff_B_a3vhh17j0_2),.clk(gclk));
	jdff dff_B_8KXdKmmc6_1(.din(n399),.dout(w_dff_B_8KXdKmmc6_1),.clk(gclk));
	jdff dff_B_81DpVl7v2_2(.din(n335),.dout(w_dff_B_81DpVl7v2_2),.clk(gclk));
	jdff dff_B_kAjE0D7I4_2(.din(w_dff_B_81DpVl7v2_2),.dout(w_dff_B_kAjE0D7I4_2),.clk(gclk));
	jdff dff_B_RAeSevz53_2(.din(w_dff_B_kAjE0D7I4_2),.dout(w_dff_B_RAeSevz53_2),.clk(gclk));
	jdff dff_B_IuAArMSN9_2(.din(w_dff_B_RAeSevz53_2),.dout(w_dff_B_IuAArMSN9_2),.clk(gclk));
	jdff dff_B_DgacSUbd6_2(.din(w_dff_B_IuAArMSN9_2),.dout(w_dff_B_DgacSUbd6_2),.clk(gclk));
	jdff dff_B_N6zbtjUG2_2(.din(w_dff_B_DgacSUbd6_2),.dout(w_dff_B_N6zbtjUG2_2),.clk(gclk));
	jdff dff_B_87EYA9Y24_2(.din(w_dff_B_N6zbtjUG2_2),.dout(w_dff_B_87EYA9Y24_2),.clk(gclk));
	jdff dff_B_j7nDCuoL8_2(.din(w_dff_B_87EYA9Y24_2),.dout(w_dff_B_j7nDCuoL8_2),.clk(gclk));
	jdff dff_B_7EixtPTM1_2(.din(w_dff_B_j7nDCuoL8_2),.dout(w_dff_B_7EixtPTM1_2),.clk(gclk));
	jdff dff_B_eJVg4sHJ5_2(.din(w_dff_B_7EixtPTM1_2),.dout(w_dff_B_eJVg4sHJ5_2),.clk(gclk));
	jdff dff_B_VMoPedRs6_2(.din(w_dff_B_eJVg4sHJ5_2),.dout(w_dff_B_VMoPedRs6_2),.clk(gclk));
	jdff dff_B_01JQ4hfl9_2(.din(w_dff_B_VMoPedRs6_2),.dout(w_dff_B_01JQ4hfl9_2),.clk(gclk));
	jdff dff_B_DjleBzKY8_2(.din(w_dff_B_01JQ4hfl9_2),.dout(w_dff_B_DjleBzKY8_2),.clk(gclk));
	jdff dff_B_c9L2D4CH9_2(.din(w_dff_B_DjleBzKY8_2),.dout(w_dff_B_c9L2D4CH9_2),.clk(gclk));
	jdff dff_B_4GGfpT8Z2_2(.din(w_dff_B_c9L2D4CH9_2),.dout(w_dff_B_4GGfpT8Z2_2),.clk(gclk));
	jdff dff_B_hUuxM9Cj6_2(.din(n370),.dout(w_dff_B_hUuxM9Cj6_2),.clk(gclk));
	jdff dff_B_npBmo3FI2_1(.din(n336),.dout(w_dff_B_npBmo3FI2_1),.clk(gclk));
	jdff dff_B_RhK0niGN5_2(.din(n279),.dout(w_dff_B_RhK0niGN5_2),.clk(gclk));
	jdff dff_B_OEwf7hP66_2(.din(w_dff_B_RhK0niGN5_2),.dout(w_dff_B_OEwf7hP66_2),.clk(gclk));
	jdff dff_B_MtaKCeQ73_2(.din(w_dff_B_OEwf7hP66_2),.dout(w_dff_B_MtaKCeQ73_2),.clk(gclk));
	jdff dff_B_cqrkvAVp5_2(.din(w_dff_B_MtaKCeQ73_2),.dout(w_dff_B_cqrkvAVp5_2),.clk(gclk));
	jdff dff_B_NgYT9d8Q1_2(.din(w_dff_B_cqrkvAVp5_2),.dout(w_dff_B_NgYT9d8Q1_2),.clk(gclk));
	jdff dff_B_K1oAFODJ0_2(.din(w_dff_B_NgYT9d8Q1_2),.dout(w_dff_B_K1oAFODJ0_2),.clk(gclk));
	jdff dff_B_7lGNjVI75_2(.din(w_dff_B_K1oAFODJ0_2),.dout(w_dff_B_7lGNjVI75_2),.clk(gclk));
	jdff dff_B_kWvFYJsq6_2(.din(w_dff_B_7lGNjVI75_2),.dout(w_dff_B_kWvFYJsq6_2),.clk(gclk));
	jdff dff_B_1vqvDT3b4_2(.din(w_dff_B_kWvFYJsq6_2),.dout(w_dff_B_1vqvDT3b4_2),.clk(gclk));
	jdff dff_B_4jZlZdKo0_2(.din(w_dff_B_1vqvDT3b4_2),.dout(w_dff_B_4jZlZdKo0_2),.clk(gclk));
	jdff dff_B_eHDaJjSf8_2(.din(w_dff_B_4jZlZdKo0_2),.dout(w_dff_B_eHDaJjSf8_2),.clk(gclk));
	jdff dff_B_YuxiLJVP8_2(.din(w_dff_B_eHDaJjSf8_2),.dout(w_dff_B_YuxiLJVP8_2),.clk(gclk));
	jdff dff_B_FPWiNprk3_2(.din(n307),.dout(w_dff_B_FPWiNprk3_2),.clk(gclk));
	jdff dff_B_Y4Mwki8N8_1(.din(n280),.dout(w_dff_B_Y4Mwki8N8_1),.clk(gclk));
	jdff dff_B_buPbW46o2_2(.din(n230),.dout(w_dff_B_buPbW46o2_2),.clk(gclk));
	jdff dff_B_SDqNf5448_2(.din(w_dff_B_buPbW46o2_2),.dout(w_dff_B_SDqNf5448_2),.clk(gclk));
	jdff dff_B_jdejU4C27_2(.din(w_dff_B_SDqNf5448_2),.dout(w_dff_B_jdejU4C27_2),.clk(gclk));
	jdff dff_B_0AFkGHTD9_2(.din(w_dff_B_jdejU4C27_2),.dout(w_dff_B_0AFkGHTD9_2),.clk(gclk));
	jdff dff_B_NAGmiFYT7_2(.din(w_dff_B_0AFkGHTD9_2),.dout(w_dff_B_NAGmiFYT7_2),.clk(gclk));
	jdff dff_B_taqlKBRo7_2(.din(w_dff_B_NAGmiFYT7_2),.dout(w_dff_B_taqlKBRo7_2),.clk(gclk));
	jdff dff_B_brYJ81LH6_2(.din(w_dff_B_taqlKBRo7_2),.dout(w_dff_B_brYJ81LH6_2),.clk(gclk));
	jdff dff_B_lNswk0dg6_2(.din(w_dff_B_brYJ81LH6_2),.dout(w_dff_B_lNswk0dg6_2),.clk(gclk));
	jdff dff_B_NoOfWuhP6_2(.din(w_dff_B_lNswk0dg6_2),.dout(w_dff_B_NoOfWuhP6_2),.clk(gclk));
	jdff dff_B_uVj7vMka2_2(.din(n251),.dout(w_dff_B_uVj7vMka2_2),.clk(gclk));
	jdff dff_B_FHDfKqcc2_1(.din(n231),.dout(w_dff_B_FHDfKqcc2_1),.clk(gclk));
	jdff dff_B_fUk4hqjq2_2(.din(n188),.dout(w_dff_B_fUk4hqjq2_2),.clk(gclk));
	jdff dff_B_NMJW5qQQ6_2(.din(w_dff_B_fUk4hqjq2_2),.dout(w_dff_B_NMJW5qQQ6_2),.clk(gclk));
	jdff dff_B_p0VVpxOD7_2(.din(w_dff_B_NMJW5qQQ6_2),.dout(w_dff_B_p0VVpxOD7_2),.clk(gclk));
	jdff dff_B_fcmW6xwU6_2(.din(w_dff_B_p0VVpxOD7_2),.dout(w_dff_B_fcmW6xwU6_2),.clk(gclk));
	jdff dff_B_guLnpw2S4_2(.din(w_dff_B_fcmW6xwU6_2),.dout(w_dff_B_guLnpw2S4_2),.clk(gclk));
	jdff dff_B_Z7m1PGz53_2(.din(w_dff_B_guLnpw2S4_2),.dout(w_dff_B_Z7m1PGz53_2),.clk(gclk));
	jdff dff_B_9pL1rP5c5_2(.din(n202),.dout(w_dff_B_9pL1rP5c5_2),.clk(gclk));
	jdff dff_B_2iH3l9Ps9_2(.din(n154),.dout(w_dff_B_2iH3l9Ps9_2),.clk(gclk));
	jdff dff_B_rcPjiLWS1_2(.din(w_dff_B_2iH3l9Ps9_2),.dout(w_dff_B_rcPjiLWS1_2),.clk(gclk));
	jdff dff_B_qFMZlzBN6_2(.din(w_dff_B_rcPjiLWS1_2),.dout(w_dff_B_qFMZlzBN6_2),.clk(gclk));
	jdff dff_B_p96wqOZf1_0(.din(n159),.dout(w_dff_B_p96wqOZf1_0),.clk(gclk));
	jdff dff_A_hn2ihA4X7_0(.dout(w_n123_0[0]),.din(w_dff_A_hn2ihA4X7_0),.clk(gclk));
	jdff dff_A_uRE18QYz7_0(.dout(w_dff_A_hn2ihA4X7_0),.din(w_dff_A_uRE18QYz7_0),.clk(gclk));
	jdff dff_A_9DHjInrX5_0(.dout(w_n122_0[0]),.din(w_dff_A_9DHjInrX5_0),.clk(gclk));
	jdff dff_A_VnVkTe6E1_0(.dout(w_dff_A_9DHjInrX5_0),.din(w_dff_A_VnVkTe6E1_0),.clk(gclk));
	jdff dff_B_QzRqY8Wk5_1(.din(n1304),.dout(w_dff_B_QzRqY8Wk5_1),.clk(gclk));
	jdff dff_B_EkBsbp5C6_2(.din(n1217),.dout(w_dff_B_EkBsbp5C6_2),.clk(gclk));
	jdff dff_B_V9gy66MR8_2(.din(w_dff_B_EkBsbp5C6_2),.dout(w_dff_B_V9gy66MR8_2),.clk(gclk));
	jdff dff_B_yvxOb0tX3_2(.din(w_dff_B_V9gy66MR8_2),.dout(w_dff_B_yvxOb0tX3_2),.clk(gclk));
	jdff dff_B_0htVR8JQ3_2(.din(w_dff_B_yvxOb0tX3_2),.dout(w_dff_B_0htVR8JQ3_2),.clk(gclk));
	jdff dff_B_kgx9rspv3_2(.din(w_dff_B_0htVR8JQ3_2),.dout(w_dff_B_kgx9rspv3_2),.clk(gclk));
	jdff dff_B_wW5J3Qoh9_2(.din(w_dff_B_kgx9rspv3_2),.dout(w_dff_B_wW5J3Qoh9_2),.clk(gclk));
	jdff dff_B_soxLtRFc3_2(.din(w_dff_B_wW5J3Qoh9_2),.dout(w_dff_B_soxLtRFc3_2),.clk(gclk));
	jdff dff_B_FWVnXE4p0_2(.din(w_dff_B_soxLtRFc3_2),.dout(w_dff_B_FWVnXE4p0_2),.clk(gclk));
	jdff dff_B_WzvgQYNR4_2(.din(w_dff_B_FWVnXE4p0_2),.dout(w_dff_B_WzvgQYNR4_2),.clk(gclk));
	jdff dff_B_mAyzAEGv6_2(.din(w_dff_B_WzvgQYNR4_2),.dout(w_dff_B_mAyzAEGv6_2),.clk(gclk));
	jdff dff_B_5kND4eji3_2(.din(w_dff_B_mAyzAEGv6_2),.dout(w_dff_B_5kND4eji3_2),.clk(gclk));
	jdff dff_B_DbAaB1HS5_2(.din(w_dff_B_5kND4eji3_2),.dout(w_dff_B_DbAaB1HS5_2),.clk(gclk));
	jdff dff_B_e4KXCDof2_2(.din(w_dff_B_DbAaB1HS5_2),.dout(w_dff_B_e4KXCDof2_2),.clk(gclk));
	jdff dff_B_49mKgtxF0_2(.din(w_dff_B_e4KXCDof2_2),.dout(w_dff_B_49mKgtxF0_2),.clk(gclk));
	jdff dff_B_9CdU1SOe2_2(.din(w_dff_B_49mKgtxF0_2),.dout(w_dff_B_9CdU1SOe2_2),.clk(gclk));
	jdff dff_B_5hYqEvx10_2(.din(w_dff_B_9CdU1SOe2_2),.dout(w_dff_B_5hYqEvx10_2),.clk(gclk));
	jdff dff_B_pvutrAiR3_2(.din(w_dff_B_5hYqEvx10_2),.dout(w_dff_B_pvutrAiR3_2),.clk(gclk));
	jdff dff_B_AqLBlfe52_2(.din(w_dff_B_pvutrAiR3_2),.dout(w_dff_B_AqLBlfe52_2),.clk(gclk));
	jdff dff_B_2GA041mq3_2(.din(w_dff_B_AqLBlfe52_2),.dout(w_dff_B_2GA041mq3_2),.clk(gclk));
	jdff dff_B_C2zU20Io9_2(.din(w_dff_B_2GA041mq3_2),.dout(w_dff_B_C2zU20Io9_2),.clk(gclk));
	jdff dff_B_rU33edgr0_2(.din(w_dff_B_C2zU20Io9_2),.dout(w_dff_B_rU33edgr0_2),.clk(gclk));
	jdff dff_B_OjLXyaVm5_2(.din(w_dff_B_rU33edgr0_2),.dout(w_dff_B_OjLXyaVm5_2),.clk(gclk));
	jdff dff_B_81I1jSqI7_2(.din(w_dff_B_OjLXyaVm5_2),.dout(w_dff_B_81I1jSqI7_2),.clk(gclk));
	jdff dff_B_U93Whbfi2_2(.din(w_dff_B_81I1jSqI7_2),.dout(w_dff_B_U93Whbfi2_2),.clk(gclk));
	jdff dff_B_OyWiSILw4_2(.din(w_dff_B_U93Whbfi2_2),.dout(w_dff_B_OyWiSILw4_2),.clk(gclk));
	jdff dff_B_4PLsqf2P9_2(.din(w_dff_B_OyWiSILw4_2),.dout(w_dff_B_4PLsqf2P9_2),.clk(gclk));
	jdff dff_B_YFt1gIIa4_2(.din(w_dff_B_4PLsqf2P9_2),.dout(w_dff_B_YFt1gIIa4_2),.clk(gclk));
	jdff dff_B_v7PNWjxa0_2(.din(w_dff_B_YFt1gIIa4_2),.dout(w_dff_B_v7PNWjxa0_2),.clk(gclk));
	jdff dff_B_z7Ry1QkT6_2(.din(w_dff_B_v7PNWjxa0_2),.dout(w_dff_B_z7Ry1QkT6_2),.clk(gclk));
	jdff dff_B_cDt5Zpe71_2(.din(w_dff_B_z7Ry1QkT6_2),.dout(w_dff_B_cDt5Zpe71_2),.clk(gclk));
	jdff dff_B_OoEpJWQ75_2(.din(w_dff_B_cDt5Zpe71_2),.dout(w_dff_B_OoEpJWQ75_2),.clk(gclk));
	jdff dff_B_qZ5tv5vY1_2(.din(w_dff_B_OoEpJWQ75_2),.dout(w_dff_B_qZ5tv5vY1_2),.clk(gclk));
	jdff dff_B_kwTMnRty0_2(.din(w_dff_B_qZ5tv5vY1_2),.dout(w_dff_B_kwTMnRty0_2),.clk(gclk));
	jdff dff_B_1Xdjdf6N3_2(.din(w_dff_B_kwTMnRty0_2),.dout(w_dff_B_1Xdjdf6N3_2),.clk(gclk));
	jdff dff_B_Pmgh6Obo0_2(.din(w_dff_B_1Xdjdf6N3_2),.dout(w_dff_B_Pmgh6Obo0_2),.clk(gclk));
	jdff dff_B_AnrDfWcl1_2(.din(w_dff_B_Pmgh6Obo0_2),.dout(w_dff_B_AnrDfWcl1_2),.clk(gclk));
	jdff dff_B_cROquOB40_2(.din(w_dff_B_AnrDfWcl1_2),.dout(w_dff_B_cROquOB40_2),.clk(gclk));
	jdff dff_B_8iPXoG4N2_2(.din(w_dff_B_cROquOB40_2),.dout(w_dff_B_8iPXoG4N2_2),.clk(gclk));
	jdff dff_B_dFmAg3GA4_2(.din(w_dff_B_8iPXoG4N2_2),.dout(w_dff_B_dFmAg3GA4_2),.clk(gclk));
	jdff dff_B_MBQbCFaM1_2(.din(w_dff_B_dFmAg3GA4_2),.dout(w_dff_B_MBQbCFaM1_2),.clk(gclk));
	jdff dff_B_r03NUlUN3_2(.din(w_dff_B_MBQbCFaM1_2),.dout(w_dff_B_r03NUlUN3_2),.clk(gclk));
	jdff dff_B_XQyldepu8_2(.din(w_dff_B_r03NUlUN3_2),.dout(w_dff_B_XQyldepu8_2),.clk(gclk));
	jdff dff_B_ihKtn3974_2(.din(w_dff_B_XQyldepu8_2),.dout(w_dff_B_ihKtn3974_2),.clk(gclk));
	jdff dff_B_lMmJApGb6_2(.din(w_dff_B_ihKtn3974_2),.dout(w_dff_B_lMmJApGb6_2),.clk(gclk));
	jdff dff_B_qZbCVfzj9_0(.din(n1303),.dout(w_dff_B_qZbCVfzj9_0),.clk(gclk));
	jdff dff_A_KSJU7kjs1_1(.dout(w_n1291_0[1]),.din(w_dff_A_KSJU7kjs1_1),.clk(gclk));
	jdff dff_B_PIGqr8be1_1(.din(n1218),.dout(w_dff_B_PIGqr8be1_1),.clk(gclk));
	jdff dff_B_Ty8a6ple1_2(.din(n1126),.dout(w_dff_B_Ty8a6ple1_2),.clk(gclk));
	jdff dff_B_TgjVLXRI8_2(.din(w_dff_B_Ty8a6ple1_2),.dout(w_dff_B_TgjVLXRI8_2),.clk(gclk));
	jdff dff_B_iX1SIyCK9_2(.din(w_dff_B_TgjVLXRI8_2),.dout(w_dff_B_iX1SIyCK9_2),.clk(gclk));
	jdff dff_B_Bpbbljzn2_2(.din(w_dff_B_iX1SIyCK9_2),.dout(w_dff_B_Bpbbljzn2_2),.clk(gclk));
	jdff dff_B_BWbAjSqr9_2(.din(w_dff_B_Bpbbljzn2_2),.dout(w_dff_B_BWbAjSqr9_2),.clk(gclk));
	jdff dff_B_QiCnsXfR8_2(.din(w_dff_B_BWbAjSqr9_2),.dout(w_dff_B_QiCnsXfR8_2),.clk(gclk));
	jdff dff_B_ndOyVV2j6_2(.din(w_dff_B_QiCnsXfR8_2),.dout(w_dff_B_ndOyVV2j6_2),.clk(gclk));
	jdff dff_B_61lASTgb5_2(.din(w_dff_B_ndOyVV2j6_2),.dout(w_dff_B_61lASTgb5_2),.clk(gclk));
	jdff dff_B_5DdOldDp4_2(.din(w_dff_B_61lASTgb5_2),.dout(w_dff_B_5DdOldDp4_2),.clk(gclk));
	jdff dff_B_MW2rohRv5_2(.din(w_dff_B_5DdOldDp4_2),.dout(w_dff_B_MW2rohRv5_2),.clk(gclk));
	jdff dff_B_vw7WS6Vh2_2(.din(w_dff_B_MW2rohRv5_2),.dout(w_dff_B_vw7WS6Vh2_2),.clk(gclk));
	jdff dff_B_O72Qgpf74_2(.din(w_dff_B_vw7WS6Vh2_2),.dout(w_dff_B_O72Qgpf74_2),.clk(gclk));
	jdff dff_B_y1TaDchZ3_2(.din(w_dff_B_O72Qgpf74_2),.dout(w_dff_B_y1TaDchZ3_2),.clk(gclk));
	jdff dff_B_tUTWzf819_2(.din(w_dff_B_y1TaDchZ3_2),.dout(w_dff_B_tUTWzf819_2),.clk(gclk));
	jdff dff_B_YFiYT1dE0_2(.din(w_dff_B_tUTWzf819_2),.dout(w_dff_B_YFiYT1dE0_2),.clk(gclk));
	jdff dff_B_zvHLBJFV5_2(.din(w_dff_B_YFiYT1dE0_2),.dout(w_dff_B_zvHLBJFV5_2),.clk(gclk));
	jdff dff_B_2Mx7iK5f4_2(.din(w_dff_B_zvHLBJFV5_2),.dout(w_dff_B_2Mx7iK5f4_2),.clk(gclk));
	jdff dff_B_bRBWLhek8_2(.din(w_dff_B_2Mx7iK5f4_2),.dout(w_dff_B_bRBWLhek8_2),.clk(gclk));
	jdff dff_B_otkSlVI13_2(.din(w_dff_B_bRBWLhek8_2),.dout(w_dff_B_otkSlVI13_2),.clk(gclk));
	jdff dff_B_ENapcN2Q7_2(.din(w_dff_B_otkSlVI13_2),.dout(w_dff_B_ENapcN2Q7_2),.clk(gclk));
	jdff dff_B_wznB5eDK4_2(.din(w_dff_B_ENapcN2Q7_2),.dout(w_dff_B_wznB5eDK4_2),.clk(gclk));
	jdff dff_B_3GKlaIZe6_2(.din(w_dff_B_wznB5eDK4_2),.dout(w_dff_B_3GKlaIZe6_2),.clk(gclk));
	jdff dff_B_uoHfKMwe3_2(.din(w_dff_B_3GKlaIZe6_2),.dout(w_dff_B_uoHfKMwe3_2),.clk(gclk));
	jdff dff_B_QUFRqTmT9_2(.din(w_dff_B_uoHfKMwe3_2),.dout(w_dff_B_QUFRqTmT9_2),.clk(gclk));
	jdff dff_B_DtG11sPz5_2(.din(w_dff_B_QUFRqTmT9_2),.dout(w_dff_B_DtG11sPz5_2),.clk(gclk));
	jdff dff_B_XgtGxpl03_2(.din(w_dff_B_DtG11sPz5_2),.dout(w_dff_B_XgtGxpl03_2),.clk(gclk));
	jdff dff_B_1vmPD2DE7_2(.din(w_dff_B_XgtGxpl03_2),.dout(w_dff_B_1vmPD2DE7_2),.clk(gclk));
	jdff dff_B_YZQ42WSY0_2(.din(w_dff_B_1vmPD2DE7_2),.dout(w_dff_B_YZQ42WSY0_2),.clk(gclk));
	jdff dff_B_KYsVBEqh2_2(.din(w_dff_B_YZQ42WSY0_2),.dout(w_dff_B_KYsVBEqh2_2),.clk(gclk));
	jdff dff_B_sQAQDt9x0_2(.din(w_dff_B_KYsVBEqh2_2),.dout(w_dff_B_sQAQDt9x0_2),.clk(gclk));
	jdff dff_B_oyWSxQ8s7_2(.din(w_dff_B_sQAQDt9x0_2),.dout(w_dff_B_oyWSxQ8s7_2),.clk(gclk));
	jdff dff_B_VVkazXL08_2(.din(w_dff_B_oyWSxQ8s7_2),.dout(w_dff_B_VVkazXL08_2),.clk(gclk));
	jdff dff_B_p14iwy2s5_2(.din(w_dff_B_VVkazXL08_2),.dout(w_dff_B_p14iwy2s5_2),.clk(gclk));
	jdff dff_B_nWvH51cH1_2(.din(w_dff_B_p14iwy2s5_2),.dout(w_dff_B_nWvH51cH1_2),.clk(gclk));
	jdff dff_B_mXrTqje64_2(.din(w_dff_B_nWvH51cH1_2),.dout(w_dff_B_mXrTqje64_2),.clk(gclk));
	jdff dff_B_mMzPzBnB3_2(.din(w_dff_B_mXrTqje64_2),.dout(w_dff_B_mMzPzBnB3_2),.clk(gclk));
	jdff dff_B_pDd7DsGf2_2(.din(w_dff_B_mMzPzBnB3_2),.dout(w_dff_B_pDd7DsGf2_2),.clk(gclk));
	jdff dff_B_7UA23h9k2_2(.din(w_dff_B_pDd7DsGf2_2),.dout(w_dff_B_7UA23h9k2_2),.clk(gclk));
	jdff dff_B_b70qJSYz4_2(.din(w_dff_B_7UA23h9k2_2),.dout(w_dff_B_b70qJSYz4_2),.clk(gclk));
	jdff dff_B_5iKIACOp3_2(.din(n1200),.dout(w_dff_B_5iKIACOp3_2),.clk(gclk));
	jdff dff_B_sd11iQz02_1(.din(n1127),.dout(w_dff_B_sd11iQz02_1),.clk(gclk));
	jdff dff_B_hEbWQPmX7_2(.din(n1028),.dout(w_dff_B_hEbWQPmX7_2),.clk(gclk));
	jdff dff_B_iSAHyJDU1_2(.din(w_dff_B_hEbWQPmX7_2),.dout(w_dff_B_iSAHyJDU1_2),.clk(gclk));
	jdff dff_B_fWquE1lm3_2(.din(w_dff_B_iSAHyJDU1_2),.dout(w_dff_B_fWquE1lm3_2),.clk(gclk));
	jdff dff_B_IXoj6phy2_2(.din(w_dff_B_fWquE1lm3_2),.dout(w_dff_B_IXoj6phy2_2),.clk(gclk));
	jdff dff_B_F6nurJeV8_2(.din(w_dff_B_IXoj6phy2_2),.dout(w_dff_B_F6nurJeV8_2),.clk(gclk));
	jdff dff_B_6BhQ51V03_2(.din(w_dff_B_F6nurJeV8_2),.dout(w_dff_B_6BhQ51V03_2),.clk(gclk));
	jdff dff_B_bCwoT1087_2(.din(w_dff_B_6BhQ51V03_2),.dout(w_dff_B_bCwoT1087_2),.clk(gclk));
	jdff dff_B_63redlre2_2(.din(w_dff_B_bCwoT1087_2),.dout(w_dff_B_63redlre2_2),.clk(gclk));
	jdff dff_B_KhVip9yp2_2(.din(w_dff_B_63redlre2_2),.dout(w_dff_B_KhVip9yp2_2),.clk(gclk));
	jdff dff_B_9eFEpYFy0_2(.din(w_dff_B_KhVip9yp2_2),.dout(w_dff_B_9eFEpYFy0_2),.clk(gclk));
	jdff dff_B_IiLtqin01_2(.din(w_dff_B_9eFEpYFy0_2),.dout(w_dff_B_IiLtqin01_2),.clk(gclk));
	jdff dff_B_p2cgsK5s6_2(.din(w_dff_B_IiLtqin01_2),.dout(w_dff_B_p2cgsK5s6_2),.clk(gclk));
	jdff dff_B_of7gZplG1_2(.din(w_dff_B_p2cgsK5s6_2),.dout(w_dff_B_of7gZplG1_2),.clk(gclk));
	jdff dff_B_bs3hwhOS7_2(.din(w_dff_B_of7gZplG1_2),.dout(w_dff_B_bs3hwhOS7_2),.clk(gclk));
	jdff dff_B_eduZAaEZ4_2(.din(w_dff_B_bs3hwhOS7_2),.dout(w_dff_B_eduZAaEZ4_2),.clk(gclk));
	jdff dff_B_S0g0nGY06_2(.din(w_dff_B_eduZAaEZ4_2),.dout(w_dff_B_S0g0nGY06_2),.clk(gclk));
	jdff dff_B_3MpBENIv7_2(.din(w_dff_B_S0g0nGY06_2),.dout(w_dff_B_3MpBENIv7_2),.clk(gclk));
	jdff dff_B_wtFYxcyM4_2(.din(w_dff_B_3MpBENIv7_2),.dout(w_dff_B_wtFYxcyM4_2),.clk(gclk));
	jdff dff_B_AV4j1lCr9_2(.din(w_dff_B_wtFYxcyM4_2),.dout(w_dff_B_AV4j1lCr9_2),.clk(gclk));
	jdff dff_B_ppbbj4CA7_2(.din(w_dff_B_AV4j1lCr9_2),.dout(w_dff_B_ppbbj4CA7_2),.clk(gclk));
	jdff dff_B_CgPF2nQd7_2(.din(w_dff_B_ppbbj4CA7_2),.dout(w_dff_B_CgPF2nQd7_2),.clk(gclk));
	jdff dff_B_zHiCCIu05_2(.din(w_dff_B_CgPF2nQd7_2),.dout(w_dff_B_zHiCCIu05_2),.clk(gclk));
	jdff dff_B_LfNVZFHD4_2(.din(w_dff_B_zHiCCIu05_2),.dout(w_dff_B_LfNVZFHD4_2),.clk(gclk));
	jdff dff_B_3PL62WaT2_2(.din(w_dff_B_LfNVZFHD4_2),.dout(w_dff_B_3PL62WaT2_2),.clk(gclk));
	jdff dff_B_ZSbUGnJW2_2(.din(w_dff_B_3PL62WaT2_2),.dout(w_dff_B_ZSbUGnJW2_2),.clk(gclk));
	jdff dff_B_pWWTM2Y27_2(.din(w_dff_B_ZSbUGnJW2_2),.dout(w_dff_B_pWWTM2Y27_2),.clk(gclk));
	jdff dff_B_Al4mrGMr3_2(.din(w_dff_B_pWWTM2Y27_2),.dout(w_dff_B_Al4mrGMr3_2),.clk(gclk));
	jdff dff_B_6nyFcD707_2(.din(w_dff_B_Al4mrGMr3_2),.dout(w_dff_B_6nyFcD707_2),.clk(gclk));
	jdff dff_B_hcK1CvGR3_2(.din(w_dff_B_6nyFcD707_2),.dout(w_dff_B_hcK1CvGR3_2),.clk(gclk));
	jdff dff_B_EzUzla1W5_2(.din(w_dff_B_hcK1CvGR3_2),.dout(w_dff_B_EzUzla1W5_2),.clk(gclk));
	jdff dff_B_FmlE7YQ12_2(.din(w_dff_B_EzUzla1W5_2),.dout(w_dff_B_FmlE7YQ12_2),.clk(gclk));
	jdff dff_B_zAg5CuoL4_2(.din(w_dff_B_FmlE7YQ12_2),.dout(w_dff_B_zAg5CuoL4_2),.clk(gclk));
	jdff dff_B_cHCEvE6K0_2(.din(w_dff_B_zAg5CuoL4_2),.dout(w_dff_B_cHCEvE6K0_2),.clk(gclk));
	jdff dff_B_hiXhoUJe8_2(.din(w_dff_B_cHCEvE6K0_2),.dout(w_dff_B_hiXhoUJe8_2),.clk(gclk));
	jdff dff_B_GAIlJRWL5_2(.din(w_dff_B_hiXhoUJe8_2),.dout(w_dff_B_GAIlJRWL5_2),.clk(gclk));
	jdff dff_B_yxORPfpV4_2(.din(w_dff_B_GAIlJRWL5_2),.dout(w_dff_B_yxORPfpV4_2),.clk(gclk));
	jdff dff_B_kFtO13Jo8_2(.din(n1101),.dout(w_dff_B_kFtO13Jo8_2),.clk(gclk));
	jdff dff_B_h5RKjoXL7_1(.din(n1029),.dout(w_dff_B_h5RKjoXL7_1),.clk(gclk));
	jdff dff_B_NnjAGsoU7_2(.din(n929),.dout(w_dff_B_NnjAGsoU7_2),.clk(gclk));
	jdff dff_B_LYVkxd7D5_2(.din(w_dff_B_NnjAGsoU7_2),.dout(w_dff_B_LYVkxd7D5_2),.clk(gclk));
	jdff dff_B_VmWTAZtv4_2(.din(w_dff_B_LYVkxd7D5_2),.dout(w_dff_B_VmWTAZtv4_2),.clk(gclk));
	jdff dff_B_tnMALOZq3_2(.din(w_dff_B_VmWTAZtv4_2),.dout(w_dff_B_tnMALOZq3_2),.clk(gclk));
	jdff dff_B_d7bR3JMp8_2(.din(w_dff_B_tnMALOZq3_2),.dout(w_dff_B_d7bR3JMp8_2),.clk(gclk));
	jdff dff_B_ruUHm3AQ6_2(.din(w_dff_B_d7bR3JMp8_2),.dout(w_dff_B_ruUHm3AQ6_2),.clk(gclk));
	jdff dff_B_TC4EuuNo9_2(.din(w_dff_B_ruUHm3AQ6_2),.dout(w_dff_B_TC4EuuNo9_2),.clk(gclk));
	jdff dff_B_yM2L6Mdt9_2(.din(w_dff_B_TC4EuuNo9_2),.dout(w_dff_B_yM2L6Mdt9_2),.clk(gclk));
	jdff dff_B_0IPI0RnW8_2(.din(w_dff_B_yM2L6Mdt9_2),.dout(w_dff_B_0IPI0RnW8_2),.clk(gclk));
	jdff dff_B_Q3q1zVDc1_2(.din(w_dff_B_0IPI0RnW8_2),.dout(w_dff_B_Q3q1zVDc1_2),.clk(gclk));
	jdff dff_B_bI9xB2bZ9_2(.din(w_dff_B_Q3q1zVDc1_2),.dout(w_dff_B_bI9xB2bZ9_2),.clk(gclk));
	jdff dff_B_TjPZ7ovH1_2(.din(w_dff_B_bI9xB2bZ9_2),.dout(w_dff_B_TjPZ7ovH1_2),.clk(gclk));
	jdff dff_B_Lm9FGTjR5_2(.din(w_dff_B_TjPZ7ovH1_2),.dout(w_dff_B_Lm9FGTjR5_2),.clk(gclk));
	jdff dff_B_tZNQvoH75_2(.din(w_dff_B_Lm9FGTjR5_2),.dout(w_dff_B_tZNQvoH75_2),.clk(gclk));
	jdff dff_B_4pJm1sHH8_2(.din(w_dff_B_tZNQvoH75_2),.dout(w_dff_B_4pJm1sHH8_2),.clk(gclk));
	jdff dff_B_H4pbYAZF2_2(.din(w_dff_B_4pJm1sHH8_2),.dout(w_dff_B_H4pbYAZF2_2),.clk(gclk));
	jdff dff_B_sVdGHBeJ4_2(.din(w_dff_B_H4pbYAZF2_2),.dout(w_dff_B_sVdGHBeJ4_2),.clk(gclk));
	jdff dff_B_so5KxBVc1_2(.din(w_dff_B_sVdGHBeJ4_2),.dout(w_dff_B_so5KxBVc1_2),.clk(gclk));
	jdff dff_B_OLx5nN6y6_2(.din(w_dff_B_so5KxBVc1_2),.dout(w_dff_B_OLx5nN6y6_2),.clk(gclk));
	jdff dff_B_A6cRI4CC0_2(.din(w_dff_B_OLx5nN6y6_2),.dout(w_dff_B_A6cRI4CC0_2),.clk(gclk));
	jdff dff_B_H5aKrbt48_2(.din(w_dff_B_A6cRI4CC0_2),.dout(w_dff_B_H5aKrbt48_2),.clk(gclk));
	jdff dff_B_tQKB44Qv3_2(.din(w_dff_B_H5aKrbt48_2),.dout(w_dff_B_tQKB44Qv3_2),.clk(gclk));
	jdff dff_B_cFMP2liM2_2(.din(w_dff_B_tQKB44Qv3_2),.dout(w_dff_B_cFMP2liM2_2),.clk(gclk));
	jdff dff_B_mAIyepEz8_2(.din(w_dff_B_cFMP2liM2_2),.dout(w_dff_B_mAIyepEz8_2),.clk(gclk));
	jdff dff_B_kTr9xOqP9_2(.din(w_dff_B_mAIyepEz8_2),.dout(w_dff_B_kTr9xOqP9_2),.clk(gclk));
	jdff dff_B_vCH8Yl6s0_2(.din(w_dff_B_kTr9xOqP9_2),.dout(w_dff_B_vCH8Yl6s0_2),.clk(gclk));
	jdff dff_B_zXluw1Pn2_2(.din(w_dff_B_vCH8Yl6s0_2),.dout(w_dff_B_zXluw1Pn2_2),.clk(gclk));
	jdff dff_B_9colIbKg8_2(.din(w_dff_B_zXluw1Pn2_2),.dout(w_dff_B_9colIbKg8_2),.clk(gclk));
	jdff dff_B_ZAZGKhV92_2(.din(w_dff_B_9colIbKg8_2),.dout(w_dff_B_ZAZGKhV92_2),.clk(gclk));
	jdff dff_B_cPn2rPyx0_2(.din(w_dff_B_ZAZGKhV92_2),.dout(w_dff_B_cPn2rPyx0_2),.clk(gclk));
	jdff dff_B_cn1O666u4_2(.din(w_dff_B_cPn2rPyx0_2),.dout(w_dff_B_cn1O666u4_2),.clk(gclk));
	jdff dff_B_41p4QyuJ8_2(.din(w_dff_B_cn1O666u4_2),.dout(w_dff_B_41p4QyuJ8_2),.clk(gclk));
	jdff dff_B_uKmEUj662_2(.din(w_dff_B_41p4QyuJ8_2),.dout(w_dff_B_uKmEUj662_2),.clk(gclk));
	jdff dff_B_ZU10pe9H4_2(.din(n1002),.dout(w_dff_B_ZU10pe9H4_2),.clk(gclk));
	jdff dff_B_btAzBAx92_1(.din(n930),.dout(w_dff_B_btAzBAx92_1),.clk(gclk));
	jdff dff_B_VfH5eDLA1_2(.din(n827),.dout(w_dff_B_VfH5eDLA1_2),.clk(gclk));
	jdff dff_B_oaqYiaht3_2(.din(w_dff_B_VfH5eDLA1_2),.dout(w_dff_B_oaqYiaht3_2),.clk(gclk));
	jdff dff_B_0yXjSoOC4_2(.din(w_dff_B_oaqYiaht3_2),.dout(w_dff_B_0yXjSoOC4_2),.clk(gclk));
	jdff dff_B_0M9xiurG3_2(.din(w_dff_B_0yXjSoOC4_2),.dout(w_dff_B_0M9xiurG3_2),.clk(gclk));
	jdff dff_B_NHpPM4v32_2(.din(w_dff_B_0M9xiurG3_2),.dout(w_dff_B_NHpPM4v32_2),.clk(gclk));
	jdff dff_B_tOnSlKTU0_2(.din(w_dff_B_NHpPM4v32_2),.dout(w_dff_B_tOnSlKTU0_2),.clk(gclk));
	jdff dff_B_2ODDkCKI1_2(.din(w_dff_B_tOnSlKTU0_2),.dout(w_dff_B_2ODDkCKI1_2),.clk(gclk));
	jdff dff_B_joaL3qXE0_2(.din(w_dff_B_2ODDkCKI1_2),.dout(w_dff_B_joaL3qXE0_2),.clk(gclk));
	jdff dff_B_CLQvEiQE2_2(.din(w_dff_B_joaL3qXE0_2),.dout(w_dff_B_CLQvEiQE2_2),.clk(gclk));
	jdff dff_B_jDHRomNs2_2(.din(w_dff_B_CLQvEiQE2_2),.dout(w_dff_B_jDHRomNs2_2),.clk(gclk));
	jdff dff_B_gUogtGF26_2(.din(w_dff_B_jDHRomNs2_2),.dout(w_dff_B_gUogtGF26_2),.clk(gclk));
	jdff dff_B_OQVanudn7_2(.din(w_dff_B_gUogtGF26_2),.dout(w_dff_B_OQVanudn7_2),.clk(gclk));
	jdff dff_B_6SX5KmRQ8_2(.din(w_dff_B_OQVanudn7_2),.dout(w_dff_B_6SX5KmRQ8_2),.clk(gclk));
	jdff dff_B_yzV2Or5e4_2(.din(w_dff_B_6SX5KmRQ8_2),.dout(w_dff_B_yzV2Or5e4_2),.clk(gclk));
	jdff dff_B_tvV6kvBu0_2(.din(w_dff_B_yzV2Or5e4_2),.dout(w_dff_B_tvV6kvBu0_2),.clk(gclk));
	jdff dff_B_5K8zSqgW8_2(.din(w_dff_B_tvV6kvBu0_2),.dout(w_dff_B_5K8zSqgW8_2),.clk(gclk));
	jdff dff_B_kxCncmAs0_2(.din(w_dff_B_5K8zSqgW8_2),.dout(w_dff_B_kxCncmAs0_2),.clk(gclk));
	jdff dff_B_Ag3YV6zH0_2(.din(w_dff_B_kxCncmAs0_2),.dout(w_dff_B_Ag3YV6zH0_2),.clk(gclk));
	jdff dff_B_PlsJUzfM3_2(.din(w_dff_B_Ag3YV6zH0_2),.dout(w_dff_B_PlsJUzfM3_2),.clk(gclk));
	jdff dff_B_l2dIo4kx2_2(.din(w_dff_B_PlsJUzfM3_2),.dout(w_dff_B_l2dIo4kx2_2),.clk(gclk));
	jdff dff_B_U0akR9E61_2(.din(w_dff_B_l2dIo4kx2_2),.dout(w_dff_B_U0akR9E61_2),.clk(gclk));
	jdff dff_B_NNCM58xX8_2(.din(w_dff_B_U0akR9E61_2),.dout(w_dff_B_NNCM58xX8_2),.clk(gclk));
	jdff dff_B_oixyRztc2_2(.din(w_dff_B_NNCM58xX8_2),.dout(w_dff_B_oixyRztc2_2),.clk(gclk));
	jdff dff_B_OXM9SkIO4_2(.din(w_dff_B_oixyRztc2_2),.dout(w_dff_B_OXM9SkIO4_2),.clk(gclk));
	jdff dff_B_oC5ZLoHu2_2(.din(w_dff_B_OXM9SkIO4_2),.dout(w_dff_B_oC5ZLoHu2_2),.clk(gclk));
	jdff dff_B_mOPvEqd12_2(.din(w_dff_B_oC5ZLoHu2_2),.dout(w_dff_B_mOPvEqd12_2),.clk(gclk));
	jdff dff_B_zUZlpJFU2_2(.din(w_dff_B_mOPvEqd12_2),.dout(w_dff_B_zUZlpJFU2_2),.clk(gclk));
	jdff dff_B_5ICvawnu0_2(.din(w_dff_B_zUZlpJFU2_2),.dout(w_dff_B_5ICvawnu0_2),.clk(gclk));
	jdff dff_B_aBYRBPMW7_2(.din(w_dff_B_5ICvawnu0_2),.dout(w_dff_B_aBYRBPMW7_2),.clk(gclk));
	jdff dff_B_l0x3636S9_2(.din(w_dff_B_aBYRBPMW7_2),.dout(w_dff_B_l0x3636S9_2),.clk(gclk));
	jdff dff_B_8D3wYtpI7_2(.din(n896),.dout(w_dff_B_8D3wYtpI7_2),.clk(gclk));
	jdff dff_B_njc17Ywt8_1(.din(n828),.dout(w_dff_B_njc17Ywt8_1),.clk(gclk));
	jdff dff_B_6cC8yWm12_2(.din(n729),.dout(w_dff_B_6cC8yWm12_2),.clk(gclk));
	jdff dff_B_plZlpx0s6_2(.din(w_dff_B_6cC8yWm12_2),.dout(w_dff_B_plZlpx0s6_2),.clk(gclk));
	jdff dff_B_xb8gVmEt6_2(.din(w_dff_B_plZlpx0s6_2),.dout(w_dff_B_xb8gVmEt6_2),.clk(gclk));
	jdff dff_B_w5Xido9G2_2(.din(w_dff_B_xb8gVmEt6_2),.dout(w_dff_B_w5Xido9G2_2),.clk(gclk));
	jdff dff_B_HOPuzNZf5_2(.din(w_dff_B_w5Xido9G2_2),.dout(w_dff_B_HOPuzNZf5_2),.clk(gclk));
	jdff dff_B_Qvz7TyA18_2(.din(w_dff_B_HOPuzNZf5_2),.dout(w_dff_B_Qvz7TyA18_2),.clk(gclk));
	jdff dff_B_wuIZJW1W9_2(.din(w_dff_B_Qvz7TyA18_2),.dout(w_dff_B_wuIZJW1W9_2),.clk(gclk));
	jdff dff_B_bvELdRvx3_2(.din(w_dff_B_wuIZJW1W9_2),.dout(w_dff_B_bvELdRvx3_2),.clk(gclk));
	jdff dff_B_ceOTJzh47_2(.din(w_dff_B_bvELdRvx3_2),.dout(w_dff_B_ceOTJzh47_2),.clk(gclk));
	jdff dff_B_TKpfZjDq6_2(.din(w_dff_B_ceOTJzh47_2),.dout(w_dff_B_TKpfZjDq6_2),.clk(gclk));
	jdff dff_B_WuACwFQS9_2(.din(w_dff_B_TKpfZjDq6_2),.dout(w_dff_B_WuACwFQS9_2),.clk(gclk));
	jdff dff_B_tx0XA0783_2(.din(w_dff_B_WuACwFQS9_2),.dout(w_dff_B_tx0XA0783_2),.clk(gclk));
	jdff dff_B_NWz40CIk0_2(.din(w_dff_B_tx0XA0783_2),.dout(w_dff_B_NWz40CIk0_2),.clk(gclk));
	jdff dff_B_vIFXtAW55_2(.din(w_dff_B_NWz40CIk0_2),.dout(w_dff_B_vIFXtAW55_2),.clk(gclk));
	jdff dff_B_bzFWu4ny1_2(.din(w_dff_B_vIFXtAW55_2),.dout(w_dff_B_bzFWu4ny1_2),.clk(gclk));
	jdff dff_B_75wCUuzk0_2(.din(w_dff_B_bzFWu4ny1_2),.dout(w_dff_B_75wCUuzk0_2),.clk(gclk));
	jdff dff_B_tfdl6AfL5_2(.din(w_dff_B_75wCUuzk0_2),.dout(w_dff_B_tfdl6AfL5_2),.clk(gclk));
	jdff dff_B_YZpG7Fea5_2(.din(w_dff_B_tfdl6AfL5_2),.dout(w_dff_B_YZpG7Fea5_2),.clk(gclk));
	jdff dff_B_LaH0a9xn0_2(.din(w_dff_B_YZpG7Fea5_2),.dout(w_dff_B_LaH0a9xn0_2),.clk(gclk));
	jdff dff_B_UJ4MCAKo1_2(.din(w_dff_B_LaH0a9xn0_2),.dout(w_dff_B_UJ4MCAKo1_2),.clk(gclk));
	jdff dff_B_fOYjXp3i4_2(.din(w_dff_B_UJ4MCAKo1_2),.dout(w_dff_B_fOYjXp3i4_2),.clk(gclk));
	jdff dff_B_vJoXqYFp8_2(.din(w_dff_B_fOYjXp3i4_2),.dout(w_dff_B_vJoXqYFp8_2),.clk(gclk));
	jdff dff_B_g2y8LwN22_2(.din(w_dff_B_vJoXqYFp8_2),.dout(w_dff_B_g2y8LwN22_2),.clk(gclk));
	jdff dff_B_i2MIQDRW4_2(.din(w_dff_B_g2y8LwN22_2),.dout(w_dff_B_i2MIQDRW4_2),.clk(gclk));
	jdff dff_B_NIJGMWC59_2(.din(w_dff_B_i2MIQDRW4_2),.dout(w_dff_B_NIJGMWC59_2),.clk(gclk));
	jdff dff_B_51UgwMD87_2(.din(w_dff_B_NIJGMWC59_2),.dout(w_dff_B_51UgwMD87_2),.clk(gclk));
	jdff dff_B_uISdzOLI9_2(.din(w_dff_B_51UgwMD87_2),.dout(w_dff_B_uISdzOLI9_2),.clk(gclk));
	jdff dff_B_xUzkRPVC2_2(.din(n793),.dout(w_dff_B_xUzkRPVC2_2),.clk(gclk));
	jdff dff_B_xlYWbEmV9_1(.din(n730),.dout(w_dff_B_xlYWbEmV9_1),.clk(gclk));
	jdff dff_B_pt8vCAy86_2(.din(n637),.dout(w_dff_B_pt8vCAy86_2),.clk(gclk));
	jdff dff_B_s5txgLny6_2(.din(w_dff_B_pt8vCAy86_2),.dout(w_dff_B_s5txgLny6_2),.clk(gclk));
	jdff dff_B_t4oyNgGK6_2(.din(w_dff_B_s5txgLny6_2),.dout(w_dff_B_t4oyNgGK6_2),.clk(gclk));
	jdff dff_B_yTAOYG8R6_2(.din(w_dff_B_t4oyNgGK6_2),.dout(w_dff_B_yTAOYG8R6_2),.clk(gclk));
	jdff dff_B_qt64Ig8W3_2(.din(w_dff_B_yTAOYG8R6_2),.dout(w_dff_B_qt64Ig8W3_2),.clk(gclk));
	jdff dff_B_2Eme1FDV3_2(.din(w_dff_B_qt64Ig8W3_2),.dout(w_dff_B_2Eme1FDV3_2),.clk(gclk));
	jdff dff_B_6tjTP7AH4_2(.din(w_dff_B_2Eme1FDV3_2),.dout(w_dff_B_6tjTP7AH4_2),.clk(gclk));
	jdff dff_B_9RCxY58A2_2(.din(w_dff_B_6tjTP7AH4_2),.dout(w_dff_B_9RCxY58A2_2),.clk(gclk));
	jdff dff_B_aTQZ94k94_2(.din(w_dff_B_9RCxY58A2_2),.dout(w_dff_B_aTQZ94k94_2),.clk(gclk));
	jdff dff_B_sJyoePeo2_2(.din(w_dff_B_aTQZ94k94_2),.dout(w_dff_B_sJyoePeo2_2),.clk(gclk));
	jdff dff_B_ImeqOoTv9_2(.din(w_dff_B_sJyoePeo2_2),.dout(w_dff_B_ImeqOoTv9_2),.clk(gclk));
	jdff dff_B_1Itl3AOh3_2(.din(w_dff_B_ImeqOoTv9_2),.dout(w_dff_B_1Itl3AOh3_2),.clk(gclk));
	jdff dff_B_mZbG4vqC8_2(.din(w_dff_B_1Itl3AOh3_2),.dout(w_dff_B_mZbG4vqC8_2),.clk(gclk));
	jdff dff_B_rSfylnvx7_2(.din(w_dff_B_mZbG4vqC8_2),.dout(w_dff_B_rSfylnvx7_2),.clk(gclk));
	jdff dff_B_m61EIGg49_2(.din(w_dff_B_rSfylnvx7_2),.dout(w_dff_B_m61EIGg49_2),.clk(gclk));
	jdff dff_B_MqoDtEPs3_2(.din(w_dff_B_m61EIGg49_2),.dout(w_dff_B_MqoDtEPs3_2),.clk(gclk));
	jdff dff_B_2MiqQLhx2_2(.din(w_dff_B_MqoDtEPs3_2),.dout(w_dff_B_2MiqQLhx2_2),.clk(gclk));
	jdff dff_B_1Gyz0rPC4_2(.din(w_dff_B_2MiqQLhx2_2),.dout(w_dff_B_1Gyz0rPC4_2),.clk(gclk));
	jdff dff_B_FiWusDru0_2(.din(w_dff_B_1Gyz0rPC4_2),.dout(w_dff_B_FiWusDru0_2),.clk(gclk));
	jdff dff_B_slO8bQ4h7_2(.din(w_dff_B_FiWusDru0_2),.dout(w_dff_B_slO8bQ4h7_2),.clk(gclk));
	jdff dff_B_7A5LtFVb7_2(.din(w_dff_B_slO8bQ4h7_2),.dout(w_dff_B_7A5LtFVb7_2),.clk(gclk));
	jdff dff_B_rKjJMvQ06_2(.din(w_dff_B_7A5LtFVb7_2),.dout(w_dff_B_rKjJMvQ06_2),.clk(gclk));
	jdff dff_B_hZEEUm4Y3_2(.din(w_dff_B_rKjJMvQ06_2),.dout(w_dff_B_hZEEUm4Y3_2),.clk(gclk));
	jdff dff_B_5DMS3Dqa4_2(.din(w_dff_B_hZEEUm4Y3_2),.dout(w_dff_B_5DMS3Dqa4_2),.clk(gclk));
	jdff dff_B_cHYOWHXB5_2(.din(n694),.dout(w_dff_B_cHYOWHXB5_2),.clk(gclk));
	jdff dff_B_zA1fVh209_1(.din(n638),.dout(w_dff_B_zA1fVh209_1),.clk(gclk));
	jdff dff_B_1TX4ygRy1_2(.din(n552),.dout(w_dff_B_1TX4ygRy1_2),.clk(gclk));
	jdff dff_B_2Ap0Oqjh9_2(.din(w_dff_B_1TX4ygRy1_2),.dout(w_dff_B_2Ap0Oqjh9_2),.clk(gclk));
	jdff dff_B_fy72smUI6_2(.din(w_dff_B_2Ap0Oqjh9_2),.dout(w_dff_B_fy72smUI6_2),.clk(gclk));
	jdff dff_B_v6yxoG7W3_2(.din(w_dff_B_fy72smUI6_2),.dout(w_dff_B_v6yxoG7W3_2),.clk(gclk));
	jdff dff_B_9xjHvdEt9_2(.din(w_dff_B_v6yxoG7W3_2),.dout(w_dff_B_9xjHvdEt9_2),.clk(gclk));
	jdff dff_B_Pcfv2wn50_2(.din(w_dff_B_9xjHvdEt9_2),.dout(w_dff_B_Pcfv2wn50_2),.clk(gclk));
	jdff dff_B_XPrzWFuJ1_2(.din(w_dff_B_Pcfv2wn50_2),.dout(w_dff_B_XPrzWFuJ1_2),.clk(gclk));
	jdff dff_B_jWl5kXsp0_2(.din(w_dff_B_XPrzWFuJ1_2),.dout(w_dff_B_jWl5kXsp0_2),.clk(gclk));
	jdff dff_B_dgaqfbzw1_2(.din(w_dff_B_jWl5kXsp0_2),.dout(w_dff_B_dgaqfbzw1_2),.clk(gclk));
	jdff dff_B_moLpdjUd3_2(.din(w_dff_B_dgaqfbzw1_2),.dout(w_dff_B_moLpdjUd3_2),.clk(gclk));
	jdff dff_B_yKpLB11R7_2(.din(w_dff_B_moLpdjUd3_2),.dout(w_dff_B_yKpLB11R7_2),.clk(gclk));
	jdff dff_B_Lcg9y8Rs8_2(.din(w_dff_B_yKpLB11R7_2),.dout(w_dff_B_Lcg9y8Rs8_2),.clk(gclk));
	jdff dff_B_dYU88pkw3_2(.din(w_dff_B_Lcg9y8Rs8_2),.dout(w_dff_B_dYU88pkw3_2),.clk(gclk));
	jdff dff_B_jAOlGQVv3_2(.din(w_dff_B_dYU88pkw3_2),.dout(w_dff_B_jAOlGQVv3_2),.clk(gclk));
	jdff dff_B_anPlZ8127_2(.din(w_dff_B_jAOlGQVv3_2),.dout(w_dff_B_anPlZ8127_2),.clk(gclk));
	jdff dff_B_GHpfCaqR4_2(.din(w_dff_B_anPlZ8127_2),.dout(w_dff_B_GHpfCaqR4_2),.clk(gclk));
	jdff dff_B_RLwUrAon2_2(.din(w_dff_B_GHpfCaqR4_2),.dout(w_dff_B_RLwUrAon2_2),.clk(gclk));
	jdff dff_B_stLmgViI4_2(.din(w_dff_B_RLwUrAon2_2),.dout(w_dff_B_stLmgViI4_2),.clk(gclk));
	jdff dff_B_N3kdYXo48_2(.din(w_dff_B_stLmgViI4_2),.dout(w_dff_B_N3kdYXo48_2),.clk(gclk));
	jdff dff_B_MgyIN9sG8_2(.din(w_dff_B_N3kdYXo48_2),.dout(w_dff_B_MgyIN9sG8_2),.clk(gclk));
	jdff dff_B_EPOCiutL4_2(.din(w_dff_B_MgyIN9sG8_2),.dout(w_dff_B_EPOCiutL4_2),.clk(gclk));
	jdff dff_B_EnMmaieR2_2(.din(n602),.dout(w_dff_B_EnMmaieR2_2),.clk(gclk));
	jdff dff_B_5tQ7JrXv8_1(.din(n553),.dout(w_dff_B_5tQ7JrXv8_1),.clk(gclk));
	jdff dff_B_unxCXfma1_2(.din(n474),.dout(w_dff_B_unxCXfma1_2),.clk(gclk));
	jdff dff_B_DP6qr3E65_2(.din(w_dff_B_unxCXfma1_2),.dout(w_dff_B_DP6qr3E65_2),.clk(gclk));
	jdff dff_B_8WCx9P2a0_2(.din(w_dff_B_DP6qr3E65_2),.dout(w_dff_B_8WCx9P2a0_2),.clk(gclk));
	jdff dff_B_s9KaS7nA7_2(.din(w_dff_B_8WCx9P2a0_2),.dout(w_dff_B_s9KaS7nA7_2),.clk(gclk));
	jdff dff_B_Qk2RJZfU0_2(.din(w_dff_B_s9KaS7nA7_2),.dout(w_dff_B_Qk2RJZfU0_2),.clk(gclk));
	jdff dff_B_HucCc95M5_2(.din(w_dff_B_Qk2RJZfU0_2),.dout(w_dff_B_HucCc95M5_2),.clk(gclk));
	jdff dff_B_aEXFm0rz2_2(.din(w_dff_B_HucCc95M5_2),.dout(w_dff_B_aEXFm0rz2_2),.clk(gclk));
	jdff dff_B_8bl8lquq5_2(.din(w_dff_B_aEXFm0rz2_2),.dout(w_dff_B_8bl8lquq5_2),.clk(gclk));
	jdff dff_B_Yhzy4Ndu3_2(.din(w_dff_B_8bl8lquq5_2),.dout(w_dff_B_Yhzy4Ndu3_2),.clk(gclk));
	jdff dff_B_njnJNp6A2_2(.din(w_dff_B_Yhzy4Ndu3_2),.dout(w_dff_B_njnJNp6A2_2),.clk(gclk));
	jdff dff_B_cS8zJBEm8_2(.din(w_dff_B_njnJNp6A2_2),.dout(w_dff_B_cS8zJBEm8_2),.clk(gclk));
	jdff dff_B_5CUOBbrJ7_2(.din(w_dff_B_cS8zJBEm8_2),.dout(w_dff_B_5CUOBbrJ7_2),.clk(gclk));
	jdff dff_B_HqXxARjb4_2(.din(w_dff_B_5CUOBbrJ7_2),.dout(w_dff_B_HqXxARjb4_2),.clk(gclk));
	jdff dff_B_xOSps5fC8_2(.din(w_dff_B_HqXxARjb4_2),.dout(w_dff_B_xOSps5fC8_2),.clk(gclk));
	jdff dff_B_iZ8ykPvT0_2(.din(w_dff_B_xOSps5fC8_2),.dout(w_dff_B_iZ8ykPvT0_2),.clk(gclk));
	jdff dff_B_2ZKYKSsb9_2(.din(w_dff_B_iZ8ykPvT0_2),.dout(w_dff_B_2ZKYKSsb9_2),.clk(gclk));
	jdff dff_B_tsuREzKB2_2(.din(w_dff_B_2ZKYKSsb9_2),.dout(w_dff_B_tsuREzKB2_2),.clk(gclk));
	jdff dff_B_4CxapzYz1_2(.din(w_dff_B_tsuREzKB2_2),.dout(w_dff_B_4CxapzYz1_2),.clk(gclk));
	jdff dff_B_4qBsAPLP7_2(.din(n517),.dout(w_dff_B_4qBsAPLP7_2),.clk(gclk));
	jdff dff_B_OJBqW99N0_1(.din(n475),.dout(w_dff_B_OJBqW99N0_1),.clk(gclk));
	jdff dff_B_8TiqfJm83_2(.din(n403),.dout(w_dff_B_8TiqfJm83_2),.clk(gclk));
	jdff dff_B_spq7FsAY6_2(.din(w_dff_B_8TiqfJm83_2),.dout(w_dff_B_spq7FsAY6_2),.clk(gclk));
	jdff dff_B_iU8hxj5e1_2(.din(w_dff_B_spq7FsAY6_2),.dout(w_dff_B_iU8hxj5e1_2),.clk(gclk));
	jdff dff_B_PoU6hK8L2_2(.din(w_dff_B_iU8hxj5e1_2),.dout(w_dff_B_PoU6hK8L2_2),.clk(gclk));
	jdff dff_B_YEs4TTuI8_2(.din(w_dff_B_PoU6hK8L2_2),.dout(w_dff_B_YEs4TTuI8_2),.clk(gclk));
	jdff dff_B_aKduiEst8_2(.din(w_dff_B_YEs4TTuI8_2),.dout(w_dff_B_aKduiEst8_2),.clk(gclk));
	jdff dff_B_4qvfDN7q2_2(.din(w_dff_B_aKduiEst8_2),.dout(w_dff_B_4qvfDN7q2_2),.clk(gclk));
	jdff dff_B_8hgihRAU9_2(.din(w_dff_B_4qvfDN7q2_2),.dout(w_dff_B_8hgihRAU9_2),.clk(gclk));
	jdff dff_B_1GD3gS9O6_2(.din(w_dff_B_8hgihRAU9_2),.dout(w_dff_B_1GD3gS9O6_2),.clk(gclk));
	jdff dff_B_EOP7VZoZ8_2(.din(w_dff_B_1GD3gS9O6_2),.dout(w_dff_B_EOP7VZoZ8_2),.clk(gclk));
	jdff dff_B_lovxccja4_2(.din(w_dff_B_EOP7VZoZ8_2),.dout(w_dff_B_lovxccja4_2),.clk(gclk));
	jdff dff_B_itFyY2Vu1_2(.din(w_dff_B_lovxccja4_2),.dout(w_dff_B_itFyY2Vu1_2),.clk(gclk));
	jdff dff_B_gQntoKex1_2(.din(w_dff_B_itFyY2Vu1_2),.dout(w_dff_B_gQntoKex1_2),.clk(gclk));
	jdff dff_B_9hBpI5fz1_2(.din(w_dff_B_gQntoKex1_2),.dout(w_dff_B_9hBpI5fz1_2),.clk(gclk));
	jdff dff_B_BS4fxE5g2_2(.din(w_dff_B_9hBpI5fz1_2),.dout(w_dff_B_BS4fxE5g2_2),.clk(gclk));
	jdff dff_B_r0V17XPo8_2(.din(n439),.dout(w_dff_B_r0V17XPo8_2),.clk(gclk));
	jdff dff_B_SU23IKnx1_1(.din(n404),.dout(w_dff_B_SU23IKnx1_1),.clk(gclk));
	jdff dff_B_Qg4SlNPd6_2(.din(n340),.dout(w_dff_B_Qg4SlNPd6_2),.clk(gclk));
	jdff dff_B_mZfea7FP3_2(.din(w_dff_B_Qg4SlNPd6_2),.dout(w_dff_B_mZfea7FP3_2),.clk(gclk));
	jdff dff_B_Cq93G2qv7_2(.din(w_dff_B_mZfea7FP3_2),.dout(w_dff_B_Cq93G2qv7_2),.clk(gclk));
	jdff dff_B_kpgUEfDk0_2(.din(w_dff_B_Cq93G2qv7_2),.dout(w_dff_B_kpgUEfDk0_2),.clk(gclk));
	jdff dff_B_Kfx9Yzom1_2(.din(w_dff_B_kpgUEfDk0_2),.dout(w_dff_B_Kfx9Yzom1_2),.clk(gclk));
	jdff dff_B_FE3Gv6zn0_2(.din(w_dff_B_Kfx9Yzom1_2),.dout(w_dff_B_FE3Gv6zn0_2),.clk(gclk));
	jdff dff_B_zx2YoD5R1_2(.din(w_dff_B_FE3Gv6zn0_2),.dout(w_dff_B_zx2YoD5R1_2),.clk(gclk));
	jdff dff_B_DxyAWonr9_2(.din(w_dff_B_zx2YoD5R1_2),.dout(w_dff_B_DxyAWonr9_2),.clk(gclk));
	jdff dff_B_elgOHi1A7_2(.din(w_dff_B_DxyAWonr9_2),.dout(w_dff_B_elgOHi1A7_2),.clk(gclk));
	jdff dff_B_Hm7V5PC60_2(.din(w_dff_B_elgOHi1A7_2),.dout(w_dff_B_Hm7V5PC60_2),.clk(gclk));
	jdff dff_B_cbYwfaWm6_2(.din(w_dff_B_Hm7V5PC60_2),.dout(w_dff_B_cbYwfaWm6_2),.clk(gclk));
	jdff dff_B_aXqrKbzR6_2(.din(w_dff_B_cbYwfaWm6_2),.dout(w_dff_B_aXqrKbzR6_2),.clk(gclk));
	jdff dff_B_wdsUzH4j4_2(.din(n368),.dout(w_dff_B_wdsUzH4j4_2),.clk(gclk));
	jdff dff_B_7jaHZNBo7_1(.din(n341),.dout(w_dff_B_7jaHZNBo7_1),.clk(gclk));
	jdff dff_B_7DToSdmf9_2(.din(n284),.dout(w_dff_B_7DToSdmf9_2),.clk(gclk));
	jdff dff_B_M4yhwTvW1_2(.din(w_dff_B_7DToSdmf9_2),.dout(w_dff_B_M4yhwTvW1_2),.clk(gclk));
	jdff dff_B_lcqc8b7C2_2(.din(w_dff_B_M4yhwTvW1_2),.dout(w_dff_B_lcqc8b7C2_2),.clk(gclk));
	jdff dff_B_epfj3P5X7_2(.din(w_dff_B_lcqc8b7C2_2),.dout(w_dff_B_epfj3P5X7_2),.clk(gclk));
	jdff dff_B_MansYrIu4_2(.din(w_dff_B_epfj3P5X7_2),.dout(w_dff_B_MansYrIu4_2),.clk(gclk));
	jdff dff_B_EQiZtGhV6_2(.din(w_dff_B_MansYrIu4_2),.dout(w_dff_B_EQiZtGhV6_2),.clk(gclk));
	jdff dff_B_AdXqyWo67_2(.din(w_dff_B_EQiZtGhV6_2),.dout(w_dff_B_AdXqyWo67_2),.clk(gclk));
	jdff dff_B_JKAZmDuY8_2(.din(w_dff_B_AdXqyWo67_2),.dout(w_dff_B_JKAZmDuY8_2),.clk(gclk));
	jdff dff_B_vjmx9RdH1_2(.din(w_dff_B_JKAZmDuY8_2),.dout(w_dff_B_vjmx9RdH1_2),.clk(gclk));
	jdff dff_B_waBKwR1N6_2(.din(n305),.dout(w_dff_B_waBKwR1N6_2),.clk(gclk));
	jdff dff_B_bwQLdsF85_1(.din(n285),.dout(w_dff_B_bwQLdsF85_1),.clk(gclk));
	jdff dff_B_rWS67cWL3_2(.din(n235),.dout(w_dff_B_rWS67cWL3_2),.clk(gclk));
	jdff dff_B_eJtv3WUt9_2(.din(w_dff_B_rWS67cWL3_2),.dout(w_dff_B_eJtv3WUt9_2),.clk(gclk));
	jdff dff_B_cYqClYIx4_2(.din(w_dff_B_eJtv3WUt9_2),.dout(w_dff_B_cYqClYIx4_2),.clk(gclk));
	jdff dff_B_CV3Uu8y61_2(.din(w_dff_B_cYqClYIx4_2),.dout(w_dff_B_CV3Uu8y61_2),.clk(gclk));
	jdff dff_B_atcqW1Xi4_2(.din(w_dff_B_CV3Uu8y61_2),.dout(w_dff_B_atcqW1Xi4_2),.clk(gclk));
	jdff dff_B_MLy6fGzE4_2(.din(w_dff_B_atcqW1Xi4_2),.dout(w_dff_B_MLy6fGzE4_2),.clk(gclk));
	jdff dff_B_NTfgZDis7_2(.din(n249),.dout(w_dff_B_NTfgZDis7_2),.clk(gclk));
	jdff dff_B_pD4IhY2h2_2(.din(n194),.dout(w_dff_B_pD4IhY2h2_2),.clk(gclk));
	jdff dff_B_vgbS1Rp80_2(.din(w_dff_B_pD4IhY2h2_2),.dout(w_dff_B_vgbS1Rp80_2),.clk(gclk));
	jdff dff_B_cj34X8qx6_2(.din(w_dff_B_vgbS1Rp80_2),.dout(w_dff_B_cj34X8qx6_2),.clk(gclk));
	jdff dff_B_Bo96JeWH4_0(.din(n199),.dout(w_dff_B_Bo96JeWH4_0),.clk(gclk));
	jdff dff_A_9FnJfSj86_0(.dout(w_n157_0[0]),.din(w_dff_A_9FnJfSj86_0),.clk(gclk));
	jdff dff_A_0Gfv49f07_0(.dout(w_dff_A_9FnJfSj86_0),.din(w_dff_A_0Gfv49f07_0),.clk(gclk));
	jdff dff_A_bfPU2Rw02_0(.dout(w_n156_0[0]),.din(w_dff_A_bfPU2Rw02_0),.clk(gclk));
	jdff dff_A_NFpSeRGc1_0(.dout(w_dff_A_bfPU2Rw02_0),.din(w_dff_A_NFpSeRGc1_0),.clk(gclk));
	jdff dff_B_82kEDmpO3_2(.din(n1389),.dout(w_dff_B_82kEDmpO3_2),.clk(gclk));
	jdff dff_B_p8CFYD8r0_1(.din(n1387),.dout(w_dff_B_p8CFYD8r0_1),.clk(gclk));
	jdff dff_B_HI0qfoCK6_2(.din(n1307),.dout(w_dff_B_HI0qfoCK6_2),.clk(gclk));
	jdff dff_B_w73QtY3Q9_2(.din(w_dff_B_HI0qfoCK6_2),.dout(w_dff_B_w73QtY3Q9_2),.clk(gclk));
	jdff dff_B_LNYBxVAH7_2(.din(w_dff_B_w73QtY3Q9_2),.dout(w_dff_B_LNYBxVAH7_2),.clk(gclk));
	jdff dff_B_lPzsAtnl1_2(.din(w_dff_B_LNYBxVAH7_2),.dout(w_dff_B_lPzsAtnl1_2),.clk(gclk));
	jdff dff_B_i6rbg7Gh2_2(.din(w_dff_B_lPzsAtnl1_2),.dout(w_dff_B_i6rbg7Gh2_2),.clk(gclk));
	jdff dff_B_H2vf3QHQ9_2(.din(w_dff_B_i6rbg7Gh2_2),.dout(w_dff_B_H2vf3QHQ9_2),.clk(gclk));
	jdff dff_B_644zwNW39_2(.din(w_dff_B_H2vf3QHQ9_2),.dout(w_dff_B_644zwNW39_2),.clk(gclk));
	jdff dff_B_AUHmEi0s6_2(.din(w_dff_B_644zwNW39_2),.dout(w_dff_B_AUHmEi0s6_2),.clk(gclk));
	jdff dff_B_0XDnDoZu7_2(.din(w_dff_B_AUHmEi0s6_2),.dout(w_dff_B_0XDnDoZu7_2),.clk(gclk));
	jdff dff_B_GWh1cxgr8_2(.din(w_dff_B_0XDnDoZu7_2),.dout(w_dff_B_GWh1cxgr8_2),.clk(gclk));
	jdff dff_B_Mc1DBr5L5_2(.din(w_dff_B_GWh1cxgr8_2),.dout(w_dff_B_Mc1DBr5L5_2),.clk(gclk));
	jdff dff_B_OaBZf7ZE6_2(.din(w_dff_B_Mc1DBr5L5_2),.dout(w_dff_B_OaBZf7ZE6_2),.clk(gclk));
	jdff dff_B_58AJcBXl5_2(.din(w_dff_B_OaBZf7ZE6_2),.dout(w_dff_B_58AJcBXl5_2),.clk(gclk));
	jdff dff_B_5tmlsUO70_2(.din(w_dff_B_58AJcBXl5_2),.dout(w_dff_B_5tmlsUO70_2),.clk(gclk));
	jdff dff_B_Tmk9yV9w1_2(.din(w_dff_B_5tmlsUO70_2),.dout(w_dff_B_Tmk9yV9w1_2),.clk(gclk));
	jdff dff_B_WdOXA5mO3_2(.din(w_dff_B_Tmk9yV9w1_2),.dout(w_dff_B_WdOXA5mO3_2),.clk(gclk));
	jdff dff_B_Zs0lAgYe5_2(.din(w_dff_B_WdOXA5mO3_2),.dout(w_dff_B_Zs0lAgYe5_2),.clk(gclk));
	jdff dff_B_ZBSGuona0_2(.din(w_dff_B_Zs0lAgYe5_2),.dout(w_dff_B_ZBSGuona0_2),.clk(gclk));
	jdff dff_B_DSnE9pEi0_2(.din(w_dff_B_ZBSGuona0_2),.dout(w_dff_B_DSnE9pEi0_2),.clk(gclk));
	jdff dff_B_N3MGM5NK5_2(.din(w_dff_B_DSnE9pEi0_2),.dout(w_dff_B_N3MGM5NK5_2),.clk(gclk));
	jdff dff_B_0QJHOML52_2(.din(w_dff_B_N3MGM5NK5_2),.dout(w_dff_B_0QJHOML52_2),.clk(gclk));
	jdff dff_B_DAQtcvhJ1_2(.din(w_dff_B_0QJHOML52_2),.dout(w_dff_B_DAQtcvhJ1_2),.clk(gclk));
	jdff dff_B_JhCNHU203_2(.din(w_dff_B_DAQtcvhJ1_2),.dout(w_dff_B_JhCNHU203_2),.clk(gclk));
	jdff dff_B_iPkvAayr1_2(.din(w_dff_B_JhCNHU203_2),.dout(w_dff_B_iPkvAayr1_2),.clk(gclk));
	jdff dff_B_yIxlhDMw1_2(.din(w_dff_B_iPkvAayr1_2),.dout(w_dff_B_yIxlhDMw1_2),.clk(gclk));
	jdff dff_B_ANWPsLnT1_2(.din(w_dff_B_yIxlhDMw1_2),.dout(w_dff_B_ANWPsLnT1_2),.clk(gclk));
	jdff dff_B_8OEexEgb5_2(.din(w_dff_B_ANWPsLnT1_2),.dout(w_dff_B_8OEexEgb5_2),.clk(gclk));
	jdff dff_B_PX4UNlqr5_2(.din(w_dff_B_8OEexEgb5_2),.dout(w_dff_B_PX4UNlqr5_2),.clk(gclk));
	jdff dff_B_oa0pRPl03_2(.din(w_dff_B_PX4UNlqr5_2),.dout(w_dff_B_oa0pRPl03_2),.clk(gclk));
	jdff dff_B_FibqFtvc0_2(.din(w_dff_B_oa0pRPl03_2),.dout(w_dff_B_FibqFtvc0_2),.clk(gclk));
	jdff dff_B_zzVScD3D7_2(.din(w_dff_B_FibqFtvc0_2),.dout(w_dff_B_zzVScD3D7_2),.clk(gclk));
	jdff dff_B_luxOHkko4_2(.din(w_dff_B_zzVScD3D7_2),.dout(w_dff_B_luxOHkko4_2),.clk(gclk));
	jdff dff_B_yfR7hewW4_2(.din(w_dff_B_luxOHkko4_2),.dout(w_dff_B_yfR7hewW4_2),.clk(gclk));
	jdff dff_B_jRtBBDC25_2(.din(w_dff_B_yfR7hewW4_2),.dout(w_dff_B_jRtBBDC25_2),.clk(gclk));
	jdff dff_B_WxJYm7pB9_2(.din(w_dff_B_jRtBBDC25_2),.dout(w_dff_B_WxJYm7pB9_2),.clk(gclk));
	jdff dff_B_uMKWbvTc7_2(.din(w_dff_B_WxJYm7pB9_2),.dout(w_dff_B_uMKWbvTc7_2),.clk(gclk));
	jdff dff_B_CvaJ2SY51_2(.din(w_dff_B_uMKWbvTc7_2),.dout(w_dff_B_CvaJ2SY51_2),.clk(gclk));
	jdff dff_B_FmLZ3YRa6_2(.din(w_dff_B_CvaJ2SY51_2),.dout(w_dff_B_FmLZ3YRa6_2),.clk(gclk));
	jdff dff_B_obwItojH0_2(.din(w_dff_B_FmLZ3YRa6_2),.dout(w_dff_B_obwItojH0_2),.clk(gclk));
	jdff dff_B_bC6drbKZ5_2(.din(w_dff_B_obwItojH0_2),.dout(w_dff_B_bC6drbKZ5_2),.clk(gclk));
	jdff dff_B_2xx4hGKK8_2(.din(w_dff_B_bC6drbKZ5_2),.dout(w_dff_B_2xx4hGKK8_2),.clk(gclk));
	jdff dff_B_78y7PVT11_2(.din(w_dff_B_2xx4hGKK8_2),.dout(w_dff_B_78y7PVT11_2),.clk(gclk));
	jdff dff_B_SmH6ODnO9_2(.din(w_dff_B_78y7PVT11_2),.dout(w_dff_B_SmH6ODnO9_2),.clk(gclk));
	jdff dff_B_RRUhEdFG0_2(.din(w_dff_B_SmH6ODnO9_2),.dout(w_dff_B_RRUhEdFG0_2),.clk(gclk));
	jdff dff_B_8gNLrgrL5_1(.din(n1308),.dout(w_dff_B_8gNLrgrL5_1),.clk(gclk));
	jdff dff_B_EGvTs1xQ9_2(.din(n1222),.dout(w_dff_B_EGvTs1xQ9_2),.clk(gclk));
	jdff dff_B_vmsMTtn00_2(.din(w_dff_B_EGvTs1xQ9_2),.dout(w_dff_B_vmsMTtn00_2),.clk(gclk));
	jdff dff_B_Zzdhxzqe1_2(.din(w_dff_B_vmsMTtn00_2),.dout(w_dff_B_Zzdhxzqe1_2),.clk(gclk));
	jdff dff_B_r0mzhX8g9_2(.din(w_dff_B_Zzdhxzqe1_2),.dout(w_dff_B_r0mzhX8g9_2),.clk(gclk));
	jdff dff_B_ABwxiugB5_2(.din(w_dff_B_r0mzhX8g9_2),.dout(w_dff_B_ABwxiugB5_2),.clk(gclk));
	jdff dff_B_QmTSpFZp3_2(.din(w_dff_B_ABwxiugB5_2),.dout(w_dff_B_QmTSpFZp3_2),.clk(gclk));
	jdff dff_B_FWRpa9tG3_2(.din(w_dff_B_QmTSpFZp3_2),.dout(w_dff_B_FWRpa9tG3_2),.clk(gclk));
	jdff dff_B_CuoKJ7Sx5_2(.din(w_dff_B_FWRpa9tG3_2),.dout(w_dff_B_CuoKJ7Sx5_2),.clk(gclk));
	jdff dff_B_WowdH8jj9_2(.din(w_dff_B_CuoKJ7Sx5_2),.dout(w_dff_B_WowdH8jj9_2),.clk(gclk));
	jdff dff_B_fSLnroM98_2(.din(w_dff_B_WowdH8jj9_2),.dout(w_dff_B_fSLnroM98_2),.clk(gclk));
	jdff dff_B_SDYmAZBe9_2(.din(w_dff_B_fSLnroM98_2),.dout(w_dff_B_SDYmAZBe9_2),.clk(gclk));
	jdff dff_B_CnjXIl4S1_2(.din(w_dff_B_SDYmAZBe9_2),.dout(w_dff_B_CnjXIl4S1_2),.clk(gclk));
	jdff dff_B_RTL4yCjC8_2(.din(w_dff_B_CnjXIl4S1_2),.dout(w_dff_B_RTL4yCjC8_2),.clk(gclk));
	jdff dff_B_YEiyUClY1_2(.din(w_dff_B_RTL4yCjC8_2),.dout(w_dff_B_YEiyUClY1_2),.clk(gclk));
	jdff dff_B_M6m0kAGz4_2(.din(w_dff_B_YEiyUClY1_2),.dout(w_dff_B_M6m0kAGz4_2),.clk(gclk));
	jdff dff_B_RNWrOxw22_2(.din(w_dff_B_M6m0kAGz4_2),.dout(w_dff_B_RNWrOxw22_2),.clk(gclk));
	jdff dff_B_VZj7Jbbp9_2(.din(w_dff_B_RNWrOxw22_2),.dout(w_dff_B_VZj7Jbbp9_2),.clk(gclk));
	jdff dff_B_gL287Ds75_2(.din(w_dff_B_VZj7Jbbp9_2),.dout(w_dff_B_gL287Ds75_2),.clk(gclk));
	jdff dff_B_noyylPMX4_2(.din(w_dff_B_gL287Ds75_2),.dout(w_dff_B_noyylPMX4_2),.clk(gclk));
	jdff dff_B_GUT3ncYz4_2(.din(w_dff_B_noyylPMX4_2),.dout(w_dff_B_GUT3ncYz4_2),.clk(gclk));
	jdff dff_B_Qye8awiK7_2(.din(w_dff_B_GUT3ncYz4_2),.dout(w_dff_B_Qye8awiK7_2),.clk(gclk));
	jdff dff_B_O7kn2KFC2_2(.din(w_dff_B_Qye8awiK7_2),.dout(w_dff_B_O7kn2KFC2_2),.clk(gclk));
	jdff dff_B_xaYz8JMU4_2(.din(w_dff_B_O7kn2KFC2_2),.dout(w_dff_B_xaYz8JMU4_2),.clk(gclk));
	jdff dff_B_QzuES2Gt2_2(.din(w_dff_B_xaYz8JMU4_2),.dout(w_dff_B_QzuES2Gt2_2),.clk(gclk));
	jdff dff_B_frUWt0if3_2(.din(w_dff_B_QzuES2Gt2_2),.dout(w_dff_B_frUWt0if3_2),.clk(gclk));
	jdff dff_B_gPjMMraJ6_2(.din(w_dff_B_frUWt0if3_2),.dout(w_dff_B_gPjMMraJ6_2),.clk(gclk));
	jdff dff_B_rQAbOnRM8_2(.din(w_dff_B_gPjMMraJ6_2),.dout(w_dff_B_rQAbOnRM8_2),.clk(gclk));
	jdff dff_B_iTUhyJ955_2(.din(w_dff_B_rQAbOnRM8_2),.dout(w_dff_B_iTUhyJ955_2),.clk(gclk));
	jdff dff_B_gO1OiREC7_2(.din(w_dff_B_iTUhyJ955_2),.dout(w_dff_B_gO1OiREC7_2),.clk(gclk));
	jdff dff_B_GI2S4c4N1_2(.din(w_dff_B_gO1OiREC7_2),.dout(w_dff_B_GI2S4c4N1_2),.clk(gclk));
	jdff dff_B_PbHefd6e7_2(.din(w_dff_B_GI2S4c4N1_2),.dout(w_dff_B_PbHefd6e7_2),.clk(gclk));
	jdff dff_B_20oLcZmG6_2(.din(w_dff_B_PbHefd6e7_2),.dout(w_dff_B_20oLcZmG6_2),.clk(gclk));
	jdff dff_B_xMYI3rRT2_2(.din(w_dff_B_20oLcZmG6_2),.dout(w_dff_B_xMYI3rRT2_2),.clk(gclk));
	jdff dff_B_CSBp4CcL0_2(.din(w_dff_B_xMYI3rRT2_2),.dout(w_dff_B_CSBp4CcL0_2),.clk(gclk));
	jdff dff_B_k0b7nD5x0_2(.din(w_dff_B_CSBp4CcL0_2),.dout(w_dff_B_k0b7nD5x0_2),.clk(gclk));
	jdff dff_B_odrsetPv7_2(.din(w_dff_B_k0b7nD5x0_2),.dout(w_dff_B_odrsetPv7_2),.clk(gclk));
	jdff dff_B_CWleIVRD5_2(.din(w_dff_B_odrsetPv7_2),.dout(w_dff_B_CWleIVRD5_2),.clk(gclk));
	jdff dff_B_ZrBCp82e3_2(.din(w_dff_B_CWleIVRD5_2),.dout(w_dff_B_ZrBCp82e3_2),.clk(gclk));
	jdff dff_B_kISjt9Nd0_2(.din(w_dff_B_ZrBCp82e3_2),.dout(w_dff_B_kISjt9Nd0_2),.clk(gclk));
	jdff dff_B_6d1qojQz1_1(.din(n1223),.dout(w_dff_B_6d1qojQz1_1),.clk(gclk));
	jdff dff_B_arPmkPW94_2(.din(n1131),.dout(w_dff_B_arPmkPW94_2),.clk(gclk));
	jdff dff_B_eYb4nYSB6_2(.din(w_dff_B_arPmkPW94_2),.dout(w_dff_B_eYb4nYSB6_2),.clk(gclk));
	jdff dff_B_UA0qZu8p6_2(.din(w_dff_B_eYb4nYSB6_2),.dout(w_dff_B_UA0qZu8p6_2),.clk(gclk));
	jdff dff_B_ycShQNNf1_2(.din(w_dff_B_UA0qZu8p6_2),.dout(w_dff_B_ycShQNNf1_2),.clk(gclk));
	jdff dff_B_vwywIjc38_2(.din(w_dff_B_ycShQNNf1_2),.dout(w_dff_B_vwywIjc38_2),.clk(gclk));
	jdff dff_B_at1gFTkX8_2(.din(w_dff_B_vwywIjc38_2),.dout(w_dff_B_at1gFTkX8_2),.clk(gclk));
	jdff dff_B_cmhlqIXG9_2(.din(w_dff_B_at1gFTkX8_2),.dout(w_dff_B_cmhlqIXG9_2),.clk(gclk));
	jdff dff_B_pISZsA3N8_2(.din(w_dff_B_cmhlqIXG9_2),.dout(w_dff_B_pISZsA3N8_2),.clk(gclk));
	jdff dff_B_mMikUdx37_2(.din(w_dff_B_pISZsA3N8_2),.dout(w_dff_B_mMikUdx37_2),.clk(gclk));
	jdff dff_B_QLYrlFXX6_2(.din(w_dff_B_mMikUdx37_2),.dout(w_dff_B_QLYrlFXX6_2),.clk(gclk));
	jdff dff_B_jHcBvwUM4_2(.din(w_dff_B_QLYrlFXX6_2),.dout(w_dff_B_jHcBvwUM4_2),.clk(gclk));
	jdff dff_B_1QeLrvrj9_2(.din(w_dff_B_jHcBvwUM4_2),.dout(w_dff_B_1QeLrvrj9_2),.clk(gclk));
	jdff dff_B_y537y5px3_2(.din(w_dff_B_1QeLrvrj9_2),.dout(w_dff_B_y537y5px3_2),.clk(gclk));
	jdff dff_B_7EOGJAyi0_2(.din(w_dff_B_y537y5px3_2),.dout(w_dff_B_7EOGJAyi0_2),.clk(gclk));
	jdff dff_B_SRZiTzNW4_2(.din(w_dff_B_7EOGJAyi0_2),.dout(w_dff_B_SRZiTzNW4_2),.clk(gclk));
	jdff dff_B_BBsEUafp8_2(.din(w_dff_B_SRZiTzNW4_2),.dout(w_dff_B_BBsEUafp8_2),.clk(gclk));
	jdff dff_B_SuLWa2X11_2(.din(w_dff_B_BBsEUafp8_2),.dout(w_dff_B_SuLWa2X11_2),.clk(gclk));
	jdff dff_B_N1fq99Ep3_2(.din(w_dff_B_SuLWa2X11_2),.dout(w_dff_B_N1fq99Ep3_2),.clk(gclk));
	jdff dff_B_LbBO6qaN2_2(.din(w_dff_B_N1fq99Ep3_2),.dout(w_dff_B_LbBO6qaN2_2),.clk(gclk));
	jdff dff_B_TyOotS5b3_2(.din(w_dff_B_LbBO6qaN2_2),.dout(w_dff_B_TyOotS5b3_2),.clk(gclk));
	jdff dff_B_sG5fA6rP3_2(.din(w_dff_B_TyOotS5b3_2),.dout(w_dff_B_sG5fA6rP3_2),.clk(gclk));
	jdff dff_B_9Mr5x8V88_2(.din(w_dff_B_sG5fA6rP3_2),.dout(w_dff_B_9Mr5x8V88_2),.clk(gclk));
	jdff dff_B_5rC9Sz629_2(.din(w_dff_B_9Mr5x8V88_2),.dout(w_dff_B_5rC9Sz629_2),.clk(gclk));
	jdff dff_B_2XOD3RCs5_2(.din(w_dff_B_5rC9Sz629_2),.dout(w_dff_B_2XOD3RCs5_2),.clk(gclk));
	jdff dff_B_iUV9ddRP3_2(.din(w_dff_B_2XOD3RCs5_2),.dout(w_dff_B_iUV9ddRP3_2),.clk(gclk));
	jdff dff_B_lmhbLABn6_2(.din(w_dff_B_iUV9ddRP3_2),.dout(w_dff_B_lmhbLABn6_2),.clk(gclk));
	jdff dff_B_gd9OMT3T3_2(.din(w_dff_B_lmhbLABn6_2),.dout(w_dff_B_gd9OMT3T3_2),.clk(gclk));
	jdff dff_B_LDYzMncT7_2(.din(w_dff_B_gd9OMT3T3_2),.dout(w_dff_B_LDYzMncT7_2),.clk(gclk));
	jdff dff_B_kP9rWVYB7_2(.din(w_dff_B_LDYzMncT7_2),.dout(w_dff_B_kP9rWVYB7_2),.clk(gclk));
	jdff dff_B_0lC176QA7_2(.din(w_dff_B_kP9rWVYB7_2),.dout(w_dff_B_0lC176QA7_2),.clk(gclk));
	jdff dff_B_hQAH83qA2_2(.din(w_dff_B_0lC176QA7_2),.dout(w_dff_B_hQAH83qA2_2),.clk(gclk));
	jdff dff_B_kq3TksPn3_2(.din(w_dff_B_hQAH83qA2_2),.dout(w_dff_B_kq3TksPn3_2),.clk(gclk));
	jdff dff_B_9RGTEren2_2(.din(w_dff_B_kq3TksPn3_2),.dout(w_dff_B_9RGTEren2_2),.clk(gclk));
	jdff dff_B_eo8HzTsY9_2(.din(w_dff_B_9RGTEren2_2),.dout(w_dff_B_eo8HzTsY9_2),.clk(gclk));
	jdff dff_B_vCCULbSY1_2(.din(w_dff_B_eo8HzTsY9_2),.dout(w_dff_B_vCCULbSY1_2),.clk(gclk));
	jdff dff_B_K4Sn2Y1Z6_2(.din(w_dff_B_vCCULbSY1_2),.dout(w_dff_B_K4Sn2Y1Z6_2),.clk(gclk));
	jdff dff_B_LiVhcqFl1_1(.din(n1132),.dout(w_dff_B_LiVhcqFl1_1),.clk(gclk));
	jdff dff_B_5T1BUQmj0_2(.din(n1033),.dout(w_dff_B_5T1BUQmj0_2),.clk(gclk));
	jdff dff_B_6hDLsMDT8_2(.din(w_dff_B_5T1BUQmj0_2),.dout(w_dff_B_6hDLsMDT8_2),.clk(gclk));
	jdff dff_B_sA8hbA520_2(.din(w_dff_B_6hDLsMDT8_2),.dout(w_dff_B_sA8hbA520_2),.clk(gclk));
	jdff dff_B_THETvd4u5_2(.din(w_dff_B_sA8hbA520_2),.dout(w_dff_B_THETvd4u5_2),.clk(gclk));
	jdff dff_B_VxDt8xz84_2(.din(w_dff_B_THETvd4u5_2),.dout(w_dff_B_VxDt8xz84_2),.clk(gclk));
	jdff dff_B_xFbP1kHF3_2(.din(w_dff_B_VxDt8xz84_2),.dout(w_dff_B_xFbP1kHF3_2),.clk(gclk));
	jdff dff_B_silobUlP7_2(.din(w_dff_B_xFbP1kHF3_2),.dout(w_dff_B_silobUlP7_2),.clk(gclk));
	jdff dff_B_0jBhBDnc6_2(.din(w_dff_B_silobUlP7_2),.dout(w_dff_B_0jBhBDnc6_2),.clk(gclk));
	jdff dff_B_04O1bZi03_2(.din(w_dff_B_0jBhBDnc6_2),.dout(w_dff_B_04O1bZi03_2),.clk(gclk));
	jdff dff_B_t02yxgQk1_2(.din(w_dff_B_04O1bZi03_2),.dout(w_dff_B_t02yxgQk1_2),.clk(gclk));
	jdff dff_B_MewjG7D89_2(.din(w_dff_B_t02yxgQk1_2),.dout(w_dff_B_MewjG7D89_2),.clk(gclk));
	jdff dff_B_dFCn7i5V6_2(.din(w_dff_B_MewjG7D89_2),.dout(w_dff_B_dFCn7i5V6_2),.clk(gclk));
	jdff dff_B_aVcUdzfJ1_2(.din(w_dff_B_dFCn7i5V6_2),.dout(w_dff_B_aVcUdzfJ1_2),.clk(gclk));
	jdff dff_B_5CNxMRfU1_2(.din(w_dff_B_aVcUdzfJ1_2),.dout(w_dff_B_5CNxMRfU1_2),.clk(gclk));
	jdff dff_B_cFdAtfq98_2(.din(w_dff_B_5CNxMRfU1_2),.dout(w_dff_B_cFdAtfq98_2),.clk(gclk));
	jdff dff_B_CqDelUtY8_2(.din(w_dff_B_cFdAtfq98_2),.dout(w_dff_B_CqDelUtY8_2),.clk(gclk));
	jdff dff_B_HN26A4Ni0_2(.din(w_dff_B_CqDelUtY8_2),.dout(w_dff_B_HN26A4Ni0_2),.clk(gclk));
	jdff dff_B_ESmp7wAC2_2(.din(w_dff_B_HN26A4Ni0_2),.dout(w_dff_B_ESmp7wAC2_2),.clk(gclk));
	jdff dff_B_6SQQFuWk0_2(.din(w_dff_B_ESmp7wAC2_2),.dout(w_dff_B_6SQQFuWk0_2),.clk(gclk));
	jdff dff_B_ZdHZhSpi1_2(.din(w_dff_B_6SQQFuWk0_2),.dout(w_dff_B_ZdHZhSpi1_2),.clk(gclk));
	jdff dff_B_ydtLEszk5_2(.din(w_dff_B_ZdHZhSpi1_2),.dout(w_dff_B_ydtLEszk5_2),.clk(gclk));
	jdff dff_B_yJlNFCTq1_2(.din(w_dff_B_ydtLEszk5_2),.dout(w_dff_B_yJlNFCTq1_2),.clk(gclk));
	jdff dff_B_T9STk5IL3_2(.din(w_dff_B_yJlNFCTq1_2),.dout(w_dff_B_T9STk5IL3_2),.clk(gclk));
	jdff dff_B_jr5fRvJ45_2(.din(w_dff_B_T9STk5IL3_2),.dout(w_dff_B_jr5fRvJ45_2),.clk(gclk));
	jdff dff_B_EdQo7zSe0_2(.din(w_dff_B_jr5fRvJ45_2),.dout(w_dff_B_EdQo7zSe0_2),.clk(gclk));
	jdff dff_B_GCfu9r2u5_2(.din(w_dff_B_EdQo7zSe0_2),.dout(w_dff_B_GCfu9r2u5_2),.clk(gclk));
	jdff dff_B_GbPeGblU3_2(.din(w_dff_B_GCfu9r2u5_2),.dout(w_dff_B_GbPeGblU3_2),.clk(gclk));
	jdff dff_B_ETSuWgpd3_2(.din(w_dff_B_GbPeGblU3_2),.dout(w_dff_B_ETSuWgpd3_2),.clk(gclk));
	jdff dff_B_BBvFPJw66_2(.din(w_dff_B_ETSuWgpd3_2),.dout(w_dff_B_BBvFPJw66_2),.clk(gclk));
	jdff dff_B_ZkoKZYV51_2(.din(w_dff_B_BBvFPJw66_2),.dout(w_dff_B_ZkoKZYV51_2),.clk(gclk));
	jdff dff_B_Tv3gA1nG5_2(.din(w_dff_B_ZkoKZYV51_2),.dout(w_dff_B_Tv3gA1nG5_2),.clk(gclk));
	jdff dff_B_ExnYwyxT1_2(.din(w_dff_B_Tv3gA1nG5_2),.dout(w_dff_B_ExnYwyxT1_2),.clk(gclk));
	jdff dff_B_bJ48C7vN1_2(.din(w_dff_B_ExnYwyxT1_2),.dout(w_dff_B_bJ48C7vN1_2),.clk(gclk));
	jdff dff_B_TOvxfCyx5_1(.din(n1034),.dout(w_dff_B_TOvxfCyx5_1),.clk(gclk));
	jdff dff_B_OOBUTOR80_2(.din(n934),.dout(w_dff_B_OOBUTOR80_2),.clk(gclk));
	jdff dff_B_D8hCKFkA6_2(.din(w_dff_B_OOBUTOR80_2),.dout(w_dff_B_D8hCKFkA6_2),.clk(gclk));
	jdff dff_B_b1EnRnaB3_2(.din(w_dff_B_D8hCKFkA6_2),.dout(w_dff_B_b1EnRnaB3_2),.clk(gclk));
	jdff dff_B_BXIPDdgF9_2(.din(w_dff_B_b1EnRnaB3_2),.dout(w_dff_B_BXIPDdgF9_2),.clk(gclk));
	jdff dff_B_v2VkihFM1_2(.din(w_dff_B_BXIPDdgF9_2),.dout(w_dff_B_v2VkihFM1_2),.clk(gclk));
	jdff dff_B_AVv2Zxrm7_2(.din(w_dff_B_v2VkihFM1_2),.dout(w_dff_B_AVv2Zxrm7_2),.clk(gclk));
	jdff dff_B_MH4fLmfQ2_2(.din(w_dff_B_AVv2Zxrm7_2),.dout(w_dff_B_MH4fLmfQ2_2),.clk(gclk));
	jdff dff_B_fPbrqTmk8_2(.din(w_dff_B_MH4fLmfQ2_2),.dout(w_dff_B_fPbrqTmk8_2),.clk(gclk));
	jdff dff_B_jT1SUDCg2_2(.din(w_dff_B_fPbrqTmk8_2),.dout(w_dff_B_jT1SUDCg2_2),.clk(gclk));
	jdff dff_B_WKMyKDQw5_2(.din(w_dff_B_jT1SUDCg2_2),.dout(w_dff_B_WKMyKDQw5_2),.clk(gclk));
	jdff dff_B_mJQtkapL5_2(.din(w_dff_B_WKMyKDQw5_2),.dout(w_dff_B_mJQtkapL5_2),.clk(gclk));
	jdff dff_B_1MfXvMZP2_2(.din(w_dff_B_mJQtkapL5_2),.dout(w_dff_B_1MfXvMZP2_2),.clk(gclk));
	jdff dff_B_9DHT5X8f3_2(.din(w_dff_B_1MfXvMZP2_2),.dout(w_dff_B_9DHT5X8f3_2),.clk(gclk));
	jdff dff_B_351IfMQB1_2(.din(w_dff_B_9DHT5X8f3_2),.dout(w_dff_B_351IfMQB1_2),.clk(gclk));
	jdff dff_B_y4NHOxFn7_2(.din(w_dff_B_351IfMQB1_2),.dout(w_dff_B_y4NHOxFn7_2),.clk(gclk));
	jdff dff_B_YPCthopJ1_2(.din(w_dff_B_y4NHOxFn7_2),.dout(w_dff_B_YPCthopJ1_2),.clk(gclk));
	jdff dff_B_4awknyCS9_2(.din(w_dff_B_YPCthopJ1_2),.dout(w_dff_B_4awknyCS9_2),.clk(gclk));
	jdff dff_B_DWLC9RBZ3_2(.din(w_dff_B_4awknyCS9_2),.dout(w_dff_B_DWLC9RBZ3_2),.clk(gclk));
	jdff dff_B_OqWSA1Nw7_2(.din(w_dff_B_DWLC9RBZ3_2),.dout(w_dff_B_OqWSA1Nw7_2),.clk(gclk));
	jdff dff_B_gCtn49xw4_2(.din(w_dff_B_OqWSA1Nw7_2),.dout(w_dff_B_gCtn49xw4_2),.clk(gclk));
	jdff dff_B_Pi0nXxgR0_2(.din(w_dff_B_gCtn49xw4_2),.dout(w_dff_B_Pi0nXxgR0_2),.clk(gclk));
	jdff dff_B_8AZnS9pP3_2(.din(w_dff_B_Pi0nXxgR0_2),.dout(w_dff_B_8AZnS9pP3_2),.clk(gclk));
	jdff dff_B_Xxba8x8E1_2(.din(w_dff_B_8AZnS9pP3_2),.dout(w_dff_B_Xxba8x8E1_2),.clk(gclk));
	jdff dff_B_Ehs56RKh6_2(.din(w_dff_B_Xxba8x8E1_2),.dout(w_dff_B_Ehs56RKh6_2),.clk(gclk));
	jdff dff_B_HD4A2ZOK1_2(.din(w_dff_B_Ehs56RKh6_2),.dout(w_dff_B_HD4A2ZOK1_2),.clk(gclk));
	jdff dff_B_tGNUhpZH2_2(.din(w_dff_B_HD4A2ZOK1_2),.dout(w_dff_B_tGNUhpZH2_2),.clk(gclk));
	jdff dff_B_pfjyruZ24_2(.din(w_dff_B_tGNUhpZH2_2),.dout(w_dff_B_pfjyruZ24_2),.clk(gclk));
	jdff dff_B_JbvP0yVV6_2(.din(w_dff_B_pfjyruZ24_2),.dout(w_dff_B_JbvP0yVV6_2),.clk(gclk));
	jdff dff_B_Ob6Fd71d9_2(.din(w_dff_B_JbvP0yVV6_2),.dout(w_dff_B_Ob6Fd71d9_2),.clk(gclk));
	jdff dff_B_pOWat9C22_2(.din(w_dff_B_Ob6Fd71d9_2),.dout(w_dff_B_pOWat9C22_2),.clk(gclk));
	jdff dff_B_3pE5dkfD9_1(.din(n935),.dout(w_dff_B_3pE5dkfD9_1),.clk(gclk));
	jdff dff_B_Sdv33Ges1_2(.din(n832),.dout(w_dff_B_Sdv33Ges1_2),.clk(gclk));
	jdff dff_B_aGtrsy8H2_2(.din(w_dff_B_Sdv33Ges1_2),.dout(w_dff_B_aGtrsy8H2_2),.clk(gclk));
	jdff dff_B_gwpL6CsZ7_2(.din(w_dff_B_aGtrsy8H2_2),.dout(w_dff_B_gwpL6CsZ7_2),.clk(gclk));
	jdff dff_B_JJvg7gsc7_2(.din(w_dff_B_gwpL6CsZ7_2),.dout(w_dff_B_JJvg7gsc7_2),.clk(gclk));
	jdff dff_B_gFquDKE14_2(.din(w_dff_B_JJvg7gsc7_2),.dout(w_dff_B_gFquDKE14_2),.clk(gclk));
	jdff dff_B_IHxtHSjZ1_2(.din(w_dff_B_gFquDKE14_2),.dout(w_dff_B_IHxtHSjZ1_2),.clk(gclk));
	jdff dff_B_SP6uV0Fr4_2(.din(w_dff_B_IHxtHSjZ1_2),.dout(w_dff_B_SP6uV0Fr4_2),.clk(gclk));
	jdff dff_B_EUc7JVss8_2(.din(w_dff_B_SP6uV0Fr4_2),.dout(w_dff_B_EUc7JVss8_2),.clk(gclk));
	jdff dff_B_Gq3OZvl68_2(.din(w_dff_B_EUc7JVss8_2),.dout(w_dff_B_Gq3OZvl68_2),.clk(gclk));
	jdff dff_B_OlSijAxY2_2(.din(w_dff_B_Gq3OZvl68_2),.dout(w_dff_B_OlSijAxY2_2),.clk(gclk));
	jdff dff_B_mvxnN1Jh5_2(.din(w_dff_B_OlSijAxY2_2),.dout(w_dff_B_mvxnN1Jh5_2),.clk(gclk));
	jdff dff_B_7WigKAb76_2(.din(w_dff_B_mvxnN1Jh5_2),.dout(w_dff_B_7WigKAb76_2),.clk(gclk));
	jdff dff_B_mOah6vMx6_2(.din(w_dff_B_7WigKAb76_2),.dout(w_dff_B_mOah6vMx6_2),.clk(gclk));
	jdff dff_B_bv47knXu4_2(.din(w_dff_B_mOah6vMx6_2),.dout(w_dff_B_bv47knXu4_2),.clk(gclk));
	jdff dff_B_tujRlVA13_2(.din(w_dff_B_bv47knXu4_2),.dout(w_dff_B_tujRlVA13_2),.clk(gclk));
	jdff dff_B_ZTTkuLQJ6_2(.din(w_dff_B_tujRlVA13_2),.dout(w_dff_B_ZTTkuLQJ6_2),.clk(gclk));
	jdff dff_B_EJc5b1yF0_2(.din(w_dff_B_ZTTkuLQJ6_2),.dout(w_dff_B_EJc5b1yF0_2),.clk(gclk));
	jdff dff_B_ksKWp9c14_2(.din(w_dff_B_EJc5b1yF0_2),.dout(w_dff_B_ksKWp9c14_2),.clk(gclk));
	jdff dff_B_SERcjpHn4_2(.din(w_dff_B_ksKWp9c14_2),.dout(w_dff_B_SERcjpHn4_2),.clk(gclk));
	jdff dff_B_tvqRN6p74_2(.din(w_dff_B_SERcjpHn4_2),.dout(w_dff_B_tvqRN6p74_2),.clk(gclk));
	jdff dff_B_QfL4rNG06_2(.din(w_dff_B_tvqRN6p74_2),.dout(w_dff_B_QfL4rNG06_2),.clk(gclk));
	jdff dff_B_CZvNo3Yr6_2(.din(w_dff_B_QfL4rNG06_2),.dout(w_dff_B_CZvNo3Yr6_2),.clk(gclk));
	jdff dff_B_ucpVJGBH3_2(.din(w_dff_B_CZvNo3Yr6_2),.dout(w_dff_B_ucpVJGBH3_2),.clk(gclk));
	jdff dff_B_toF0Zfpz7_2(.din(w_dff_B_ucpVJGBH3_2),.dout(w_dff_B_toF0Zfpz7_2),.clk(gclk));
	jdff dff_B_28ZkR1Dl2_2(.din(w_dff_B_toF0Zfpz7_2),.dout(w_dff_B_28ZkR1Dl2_2),.clk(gclk));
	jdff dff_B_nS4ZgaTO2_2(.din(w_dff_B_28ZkR1Dl2_2),.dout(w_dff_B_nS4ZgaTO2_2),.clk(gclk));
	jdff dff_B_oweQ0Jal5_2(.din(w_dff_B_nS4ZgaTO2_2),.dout(w_dff_B_oweQ0Jal5_2),.clk(gclk));
	jdff dff_B_R0z19Jep3_1(.din(n833),.dout(w_dff_B_R0z19Jep3_1),.clk(gclk));
	jdff dff_B_QXRnl56v5_2(.din(n734),.dout(w_dff_B_QXRnl56v5_2),.clk(gclk));
	jdff dff_B_v8ZdHMr87_2(.din(w_dff_B_QXRnl56v5_2),.dout(w_dff_B_v8ZdHMr87_2),.clk(gclk));
	jdff dff_B_V1zqU0I55_2(.din(w_dff_B_v8ZdHMr87_2),.dout(w_dff_B_V1zqU0I55_2),.clk(gclk));
	jdff dff_B_CisTQMR80_2(.din(w_dff_B_V1zqU0I55_2),.dout(w_dff_B_CisTQMR80_2),.clk(gclk));
	jdff dff_B_fe4cb1eZ6_2(.din(w_dff_B_CisTQMR80_2),.dout(w_dff_B_fe4cb1eZ6_2),.clk(gclk));
	jdff dff_B_ijIuYNse6_2(.din(w_dff_B_fe4cb1eZ6_2),.dout(w_dff_B_ijIuYNse6_2),.clk(gclk));
	jdff dff_B_566cVKcr4_2(.din(w_dff_B_ijIuYNse6_2),.dout(w_dff_B_566cVKcr4_2),.clk(gclk));
	jdff dff_B_WqcfleWR4_2(.din(w_dff_B_566cVKcr4_2),.dout(w_dff_B_WqcfleWR4_2),.clk(gclk));
	jdff dff_B_S3eKu4XR9_2(.din(w_dff_B_WqcfleWR4_2),.dout(w_dff_B_S3eKu4XR9_2),.clk(gclk));
	jdff dff_B_pQ4tXXlM0_2(.din(w_dff_B_S3eKu4XR9_2),.dout(w_dff_B_pQ4tXXlM0_2),.clk(gclk));
	jdff dff_B_VWJBY6Ak9_2(.din(w_dff_B_pQ4tXXlM0_2),.dout(w_dff_B_VWJBY6Ak9_2),.clk(gclk));
	jdff dff_B_144ktcIl9_2(.din(w_dff_B_VWJBY6Ak9_2),.dout(w_dff_B_144ktcIl9_2),.clk(gclk));
	jdff dff_B_rTcU2Qbc6_2(.din(w_dff_B_144ktcIl9_2),.dout(w_dff_B_rTcU2Qbc6_2),.clk(gclk));
	jdff dff_B_5txrRGBZ7_2(.din(w_dff_B_rTcU2Qbc6_2),.dout(w_dff_B_5txrRGBZ7_2),.clk(gclk));
	jdff dff_B_ceTNVhgU7_2(.din(w_dff_B_5txrRGBZ7_2),.dout(w_dff_B_ceTNVhgU7_2),.clk(gclk));
	jdff dff_B_oM1CwD9C8_2(.din(w_dff_B_ceTNVhgU7_2),.dout(w_dff_B_oM1CwD9C8_2),.clk(gclk));
	jdff dff_B_FCiStozC3_2(.din(w_dff_B_oM1CwD9C8_2),.dout(w_dff_B_FCiStozC3_2),.clk(gclk));
	jdff dff_B_uCabLax15_2(.din(w_dff_B_FCiStozC3_2),.dout(w_dff_B_uCabLax15_2),.clk(gclk));
	jdff dff_B_MMFxZGqu2_2(.din(w_dff_B_uCabLax15_2),.dout(w_dff_B_MMFxZGqu2_2),.clk(gclk));
	jdff dff_B_ptfX8f457_2(.din(w_dff_B_MMFxZGqu2_2),.dout(w_dff_B_ptfX8f457_2),.clk(gclk));
	jdff dff_B_Cnn5jTTL5_2(.din(w_dff_B_ptfX8f457_2),.dout(w_dff_B_Cnn5jTTL5_2),.clk(gclk));
	jdff dff_B_2ydK2cuO5_2(.din(w_dff_B_Cnn5jTTL5_2),.dout(w_dff_B_2ydK2cuO5_2),.clk(gclk));
	jdff dff_B_ZUEycug21_2(.din(w_dff_B_2ydK2cuO5_2),.dout(w_dff_B_ZUEycug21_2),.clk(gclk));
	jdff dff_B_QgQgfMTD9_2(.din(w_dff_B_ZUEycug21_2),.dout(w_dff_B_QgQgfMTD9_2),.clk(gclk));
	jdff dff_B_y8GhzqHs6_1(.din(n735),.dout(w_dff_B_y8GhzqHs6_1),.clk(gclk));
	jdff dff_B_wKUwr2961_2(.din(n642),.dout(w_dff_B_wKUwr2961_2),.clk(gclk));
	jdff dff_B_cAHx3hjm3_2(.din(w_dff_B_wKUwr2961_2),.dout(w_dff_B_cAHx3hjm3_2),.clk(gclk));
	jdff dff_B_hZNCI5Hf4_2(.din(w_dff_B_cAHx3hjm3_2),.dout(w_dff_B_hZNCI5Hf4_2),.clk(gclk));
	jdff dff_B_sP1w03i44_2(.din(w_dff_B_hZNCI5Hf4_2),.dout(w_dff_B_sP1w03i44_2),.clk(gclk));
	jdff dff_B_9iWZnr7B6_2(.din(w_dff_B_sP1w03i44_2),.dout(w_dff_B_9iWZnr7B6_2),.clk(gclk));
	jdff dff_B_knllvzOm7_2(.din(w_dff_B_9iWZnr7B6_2),.dout(w_dff_B_knllvzOm7_2),.clk(gclk));
	jdff dff_B_8Ck0rVff5_2(.din(w_dff_B_knllvzOm7_2),.dout(w_dff_B_8Ck0rVff5_2),.clk(gclk));
	jdff dff_B_9gBWMI4B5_2(.din(w_dff_B_8Ck0rVff5_2),.dout(w_dff_B_9gBWMI4B5_2),.clk(gclk));
	jdff dff_B_rgx9td3J4_2(.din(w_dff_B_9gBWMI4B5_2),.dout(w_dff_B_rgx9td3J4_2),.clk(gclk));
	jdff dff_B_WQ171XwV0_2(.din(w_dff_B_rgx9td3J4_2),.dout(w_dff_B_WQ171XwV0_2),.clk(gclk));
	jdff dff_B_dwY2m9UF3_2(.din(w_dff_B_WQ171XwV0_2),.dout(w_dff_B_dwY2m9UF3_2),.clk(gclk));
	jdff dff_B_JUxIufPX6_2(.din(w_dff_B_dwY2m9UF3_2),.dout(w_dff_B_JUxIufPX6_2),.clk(gclk));
	jdff dff_B_PV8T9nrb8_2(.din(w_dff_B_JUxIufPX6_2),.dout(w_dff_B_PV8T9nrb8_2),.clk(gclk));
	jdff dff_B_5h6mvSNl8_2(.din(w_dff_B_PV8T9nrb8_2),.dout(w_dff_B_5h6mvSNl8_2),.clk(gclk));
	jdff dff_B_Ojy9qFaM2_2(.din(w_dff_B_5h6mvSNl8_2),.dout(w_dff_B_Ojy9qFaM2_2),.clk(gclk));
	jdff dff_B_dol2pIu93_2(.din(w_dff_B_Ojy9qFaM2_2),.dout(w_dff_B_dol2pIu93_2),.clk(gclk));
	jdff dff_B_FRJtNm0V9_2(.din(w_dff_B_dol2pIu93_2),.dout(w_dff_B_FRJtNm0V9_2),.clk(gclk));
	jdff dff_B_YOq2of3r1_2(.din(w_dff_B_FRJtNm0V9_2),.dout(w_dff_B_YOq2of3r1_2),.clk(gclk));
	jdff dff_B_IyBLy1eD9_2(.din(w_dff_B_YOq2of3r1_2),.dout(w_dff_B_IyBLy1eD9_2),.clk(gclk));
	jdff dff_B_jQaiMMzj2_2(.din(w_dff_B_IyBLy1eD9_2),.dout(w_dff_B_jQaiMMzj2_2),.clk(gclk));
	jdff dff_B_N8U5UmxG3_2(.din(w_dff_B_jQaiMMzj2_2),.dout(w_dff_B_N8U5UmxG3_2),.clk(gclk));
	jdff dff_B_tzp9z56e2_1(.din(n643),.dout(w_dff_B_tzp9z56e2_1),.clk(gclk));
	jdff dff_B_jPNCXNaj2_2(.din(n557),.dout(w_dff_B_jPNCXNaj2_2),.clk(gclk));
	jdff dff_B_Cpi0dReh1_2(.din(w_dff_B_jPNCXNaj2_2),.dout(w_dff_B_Cpi0dReh1_2),.clk(gclk));
	jdff dff_B_OWU55v149_2(.din(w_dff_B_Cpi0dReh1_2),.dout(w_dff_B_OWU55v149_2),.clk(gclk));
	jdff dff_B_wvPkt51q9_2(.din(w_dff_B_OWU55v149_2),.dout(w_dff_B_wvPkt51q9_2),.clk(gclk));
	jdff dff_B_3juSFDU49_2(.din(w_dff_B_wvPkt51q9_2),.dout(w_dff_B_3juSFDU49_2),.clk(gclk));
	jdff dff_B_Lrkf98dy0_2(.din(w_dff_B_3juSFDU49_2),.dout(w_dff_B_Lrkf98dy0_2),.clk(gclk));
	jdff dff_B_yl3iKIQG4_2(.din(w_dff_B_Lrkf98dy0_2),.dout(w_dff_B_yl3iKIQG4_2),.clk(gclk));
	jdff dff_B_yZdKaMai2_2(.din(w_dff_B_yl3iKIQG4_2),.dout(w_dff_B_yZdKaMai2_2),.clk(gclk));
	jdff dff_B_DLeQDyfQ9_2(.din(w_dff_B_yZdKaMai2_2),.dout(w_dff_B_DLeQDyfQ9_2),.clk(gclk));
	jdff dff_B_2bPKmKWU6_2(.din(w_dff_B_DLeQDyfQ9_2),.dout(w_dff_B_2bPKmKWU6_2),.clk(gclk));
	jdff dff_B_GcPNPhsu4_2(.din(w_dff_B_2bPKmKWU6_2),.dout(w_dff_B_GcPNPhsu4_2),.clk(gclk));
	jdff dff_B_rndqwl6u4_2(.din(w_dff_B_GcPNPhsu4_2),.dout(w_dff_B_rndqwl6u4_2),.clk(gclk));
	jdff dff_B_DknIx0LD7_2(.din(w_dff_B_rndqwl6u4_2),.dout(w_dff_B_DknIx0LD7_2),.clk(gclk));
	jdff dff_B_t4DhqEG94_2(.din(w_dff_B_DknIx0LD7_2),.dout(w_dff_B_t4DhqEG94_2),.clk(gclk));
	jdff dff_B_Td7YVL914_2(.din(w_dff_B_t4DhqEG94_2),.dout(w_dff_B_Td7YVL914_2),.clk(gclk));
	jdff dff_B_mlVKHcth2_2(.din(w_dff_B_Td7YVL914_2),.dout(w_dff_B_mlVKHcth2_2),.clk(gclk));
	jdff dff_B_GZaXYlnM9_2(.din(w_dff_B_mlVKHcth2_2),.dout(w_dff_B_GZaXYlnM9_2),.clk(gclk));
	jdff dff_B_ImxTX2uV5_2(.din(w_dff_B_GZaXYlnM9_2),.dout(w_dff_B_ImxTX2uV5_2),.clk(gclk));
	jdff dff_B_yLerp6T52_1(.din(n558),.dout(w_dff_B_yLerp6T52_1),.clk(gclk));
	jdff dff_B_xh23TJQr8_2(.din(n479),.dout(w_dff_B_xh23TJQr8_2),.clk(gclk));
	jdff dff_B_09jGHuYQ8_2(.din(w_dff_B_xh23TJQr8_2),.dout(w_dff_B_09jGHuYQ8_2),.clk(gclk));
	jdff dff_B_6ejMo3wB8_2(.din(w_dff_B_09jGHuYQ8_2),.dout(w_dff_B_6ejMo3wB8_2),.clk(gclk));
	jdff dff_B_c5X5DqdK8_2(.din(w_dff_B_6ejMo3wB8_2),.dout(w_dff_B_c5X5DqdK8_2),.clk(gclk));
	jdff dff_B_HGtgy4R34_2(.din(w_dff_B_c5X5DqdK8_2),.dout(w_dff_B_HGtgy4R34_2),.clk(gclk));
	jdff dff_B_yCSnzhs16_2(.din(w_dff_B_HGtgy4R34_2),.dout(w_dff_B_yCSnzhs16_2),.clk(gclk));
	jdff dff_B_SFvSsLEM0_2(.din(w_dff_B_yCSnzhs16_2),.dout(w_dff_B_SFvSsLEM0_2),.clk(gclk));
	jdff dff_B_1jqv8wRl7_2(.din(w_dff_B_SFvSsLEM0_2),.dout(w_dff_B_1jqv8wRl7_2),.clk(gclk));
	jdff dff_B_dBRo2nOc2_2(.din(w_dff_B_1jqv8wRl7_2),.dout(w_dff_B_dBRo2nOc2_2),.clk(gclk));
	jdff dff_B_ZzuDrKUA1_2(.din(w_dff_B_dBRo2nOc2_2),.dout(w_dff_B_ZzuDrKUA1_2),.clk(gclk));
	jdff dff_B_fd8RLpn81_2(.din(w_dff_B_ZzuDrKUA1_2),.dout(w_dff_B_fd8RLpn81_2),.clk(gclk));
	jdff dff_B_HZl9l0B42_2(.din(w_dff_B_fd8RLpn81_2),.dout(w_dff_B_HZl9l0B42_2),.clk(gclk));
	jdff dff_B_TcTb2V1f6_2(.din(w_dff_B_HZl9l0B42_2),.dout(w_dff_B_TcTb2V1f6_2),.clk(gclk));
	jdff dff_B_8kyQZQZ51_2(.din(w_dff_B_TcTb2V1f6_2),.dout(w_dff_B_8kyQZQZ51_2),.clk(gclk));
	jdff dff_B_JfRbc5xr0_2(.din(w_dff_B_8kyQZQZ51_2),.dout(w_dff_B_JfRbc5xr0_2),.clk(gclk));
	jdff dff_B_AwApN28D3_1(.din(n480),.dout(w_dff_B_AwApN28D3_1),.clk(gclk));
	jdff dff_B_ui3Vok8d8_2(.din(n408),.dout(w_dff_B_ui3Vok8d8_2),.clk(gclk));
	jdff dff_B_rycLXFoe9_2(.din(w_dff_B_ui3Vok8d8_2),.dout(w_dff_B_rycLXFoe9_2),.clk(gclk));
	jdff dff_B_BAIFFObf8_2(.din(w_dff_B_rycLXFoe9_2),.dout(w_dff_B_BAIFFObf8_2),.clk(gclk));
	jdff dff_B_i6dKyt5G1_2(.din(w_dff_B_BAIFFObf8_2),.dout(w_dff_B_i6dKyt5G1_2),.clk(gclk));
	jdff dff_B_zAncI7QG6_2(.din(w_dff_B_i6dKyt5G1_2),.dout(w_dff_B_zAncI7QG6_2),.clk(gclk));
	jdff dff_B_duj50ZVH5_2(.din(w_dff_B_zAncI7QG6_2),.dout(w_dff_B_duj50ZVH5_2),.clk(gclk));
	jdff dff_B_5QHiVTBT2_2(.din(w_dff_B_duj50ZVH5_2),.dout(w_dff_B_5QHiVTBT2_2),.clk(gclk));
	jdff dff_B_Eli7zVJp5_2(.din(w_dff_B_5QHiVTBT2_2),.dout(w_dff_B_Eli7zVJp5_2),.clk(gclk));
	jdff dff_B_HuYzGv3G8_2(.din(w_dff_B_Eli7zVJp5_2),.dout(w_dff_B_HuYzGv3G8_2),.clk(gclk));
	jdff dff_B_vM8hH5fA0_2(.din(w_dff_B_HuYzGv3G8_2),.dout(w_dff_B_vM8hH5fA0_2),.clk(gclk));
	jdff dff_B_2wEY9y9G1_2(.din(w_dff_B_vM8hH5fA0_2),.dout(w_dff_B_2wEY9y9G1_2),.clk(gclk));
	jdff dff_B_4Ews6Nh30_2(.din(w_dff_B_2wEY9y9G1_2),.dout(w_dff_B_4Ews6Nh30_2),.clk(gclk));
	jdff dff_B_NBaNDCuu2_1(.din(n409),.dout(w_dff_B_NBaNDCuu2_1),.clk(gclk));
	jdff dff_B_em16gT3f0_2(.din(n345),.dout(w_dff_B_em16gT3f0_2),.clk(gclk));
	jdff dff_B_UhREfVy77_2(.din(w_dff_B_em16gT3f0_2),.dout(w_dff_B_UhREfVy77_2),.clk(gclk));
	jdff dff_B_ZGV8XdVu4_2(.din(w_dff_B_UhREfVy77_2),.dout(w_dff_B_ZGV8XdVu4_2),.clk(gclk));
	jdff dff_B_FiMxoM3v3_2(.din(w_dff_B_ZGV8XdVu4_2),.dout(w_dff_B_FiMxoM3v3_2),.clk(gclk));
	jdff dff_B_NhkCPPxv1_2(.din(w_dff_B_FiMxoM3v3_2),.dout(w_dff_B_NhkCPPxv1_2),.clk(gclk));
	jdff dff_B_oWJ8I7fA0_2(.din(w_dff_B_NhkCPPxv1_2),.dout(w_dff_B_oWJ8I7fA0_2),.clk(gclk));
	jdff dff_B_U5HSUCU58_2(.din(w_dff_B_oWJ8I7fA0_2),.dout(w_dff_B_U5HSUCU58_2),.clk(gclk));
	jdff dff_B_RIt4nk6Q7_2(.din(w_dff_B_U5HSUCU58_2),.dout(w_dff_B_RIt4nk6Q7_2),.clk(gclk));
	jdff dff_B_bhrnvtsu1_2(.din(w_dff_B_RIt4nk6Q7_2),.dout(w_dff_B_bhrnvtsu1_2),.clk(gclk));
	jdff dff_B_AZjjbSdA3_2(.din(n366),.dout(w_dff_B_AZjjbSdA3_2),.clk(gclk));
	jdff dff_B_vTLeOGiF5_1(.din(n346),.dout(w_dff_B_vTLeOGiF5_1),.clk(gclk));
	jdff dff_B_96ZCAOpF3_2(.din(n289),.dout(w_dff_B_96ZCAOpF3_2),.clk(gclk));
	jdff dff_B_yrshsnC17_2(.din(w_dff_B_96ZCAOpF3_2),.dout(w_dff_B_yrshsnC17_2),.clk(gclk));
	jdff dff_B_9AaqN74H3_2(.din(w_dff_B_yrshsnC17_2),.dout(w_dff_B_9AaqN74H3_2),.clk(gclk));
	jdff dff_B_Tn8aBqFA4_2(.din(w_dff_B_9AaqN74H3_2),.dout(w_dff_B_Tn8aBqFA4_2),.clk(gclk));
	jdff dff_B_w4EXgv7l6_2(.din(w_dff_B_Tn8aBqFA4_2),.dout(w_dff_B_w4EXgv7l6_2),.clk(gclk));
	jdff dff_B_uIrpoRSt3_2(.din(w_dff_B_w4EXgv7l6_2),.dout(w_dff_B_uIrpoRSt3_2),.clk(gclk));
	jdff dff_B_008ENNDH2_2(.din(n303),.dout(w_dff_B_008ENNDH2_2),.clk(gclk));
	jdff dff_B_9mLinlEm2_2(.din(n241),.dout(w_dff_B_9mLinlEm2_2),.clk(gclk));
	jdff dff_B_lGbCP0C67_2(.din(w_dff_B_9mLinlEm2_2),.dout(w_dff_B_lGbCP0C67_2),.clk(gclk));
	jdff dff_B_lTV9VUfa5_2(.din(w_dff_B_lGbCP0C67_2),.dout(w_dff_B_lTV9VUfa5_2),.clk(gclk));
	jdff dff_B_GV8eUhdT1_0(.din(n246),.dout(w_dff_B_GV8eUhdT1_0),.clk(gclk));
	jdff dff_A_GLXUj7kV6_0(.dout(w_n196_0[0]),.din(w_dff_A_GLXUj7kV6_0),.clk(gclk));
	jdff dff_A_PJAIXXDw9_0(.dout(w_dff_A_GLXUj7kV6_0),.din(w_dff_A_PJAIXXDw9_0),.clk(gclk));
	jdff dff_A_yrorCRtU1_1(.dout(w_n196_0[1]),.din(w_dff_A_yrorCRtU1_1),.clk(gclk));
	jdff dff_A_q9M9gnBA4_1(.dout(w_dff_A_yrorCRtU1_1),.din(w_dff_A_q9M9gnBA4_1),.clk(gclk));
	jdff dff_B_w8ZEJdi97_2(.din(n1465),.dout(w_dff_B_w8ZEJdi97_2),.clk(gclk));
	jdff dff_B_3QFD0j615_1(.din(n1463),.dout(w_dff_B_3QFD0j615_1),.clk(gclk));
	jdff dff_B_k2wqKZQZ9_2(.din(n1390),.dout(w_dff_B_k2wqKZQZ9_2),.clk(gclk));
	jdff dff_B_SQ3Agozi2_2(.din(w_dff_B_k2wqKZQZ9_2),.dout(w_dff_B_SQ3Agozi2_2),.clk(gclk));
	jdff dff_B_Ub5cjh3i8_2(.din(w_dff_B_SQ3Agozi2_2),.dout(w_dff_B_Ub5cjh3i8_2),.clk(gclk));
	jdff dff_B_5c4vqkeX8_2(.din(w_dff_B_Ub5cjh3i8_2),.dout(w_dff_B_5c4vqkeX8_2),.clk(gclk));
	jdff dff_B_3Nuek61q6_2(.din(w_dff_B_5c4vqkeX8_2),.dout(w_dff_B_3Nuek61q6_2),.clk(gclk));
	jdff dff_B_sfNeiznr8_2(.din(w_dff_B_3Nuek61q6_2),.dout(w_dff_B_sfNeiznr8_2),.clk(gclk));
	jdff dff_B_Mp7ndH4q8_2(.din(w_dff_B_sfNeiznr8_2),.dout(w_dff_B_Mp7ndH4q8_2),.clk(gclk));
	jdff dff_B_ArSjtfMa1_2(.din(w_dff_B_Mp7ndH4q8_2),.dout(w_dff_B_ArSjtfMa1_2),.clk(gclk));
	jdff dff_B_wnb6lGO95_2(.din(w_dff_B_ArSjtfMa1_2),.dout(w_dff_B_wnb6lGO95_2),.clk(gclk));
	jdff dff_B_x3L7vdKr0_2(.din(w_dff_B_wnb6lGO95_2),.dout(w_dff_B_x3L7vdKr0_2),.clk(gclk));
	jdff dff_B_3pbMwHA09_2(.din(w_dff_B_x3L7vdKr0_2),.dout(w_dff_B_3pbMwHA09_2),.clk(gclk));
	jdff dff_B_CnP5aY734_2(.din(w_dff_B_3pbMwHA09_2),.dout(w_dff_B_CnP5aY734_2),.clk(gclk));
	jdff dff_B_StkDG3hZ3_2(.din(w_dff_B_CnP5aY734_2),.dout(w_dff_B_StkDG3hZ3_2),.clk(gclk));
	jdff dff_B_eybkSGqS9_2(.din(w_dff_B_StkDG3hZ3_2),.dout(w_dff_B_eybkSGqS9_2),.clk(gclk));
	jdff dff_B_AqZy4FWR8_2(.din(w_dff_B_eybkSGqS9_2),.dout(w_dff_B_AqZy4FWR8_2),.clk(gclk));
	jdff dff_B_3fuGERfV3_2(.din(w_dff_B_AqZy4FWR8_2),.dout(w_dff_B_3fuGERfV3_2),.clk(gclk));
	jdff dff_B_xO7fNMXW9_2(.din(w_dff_B_3fuGERfV3_2),.dout(w_dff_B_xO7fNMXW9_2),.clk(gclk));
	jdff dff_B_MPmlsFHX5_2(.din(w_dff_B_xO7fNMXW9_2),.dout(w_dff_B_MPmlsFHX5_2),.clk(gclk));
	jdff dff_B_QflfAzRo9_2(.din(w_dff_B_MPmlsFHX5_2),.dout(w_dff_B_QflfAzRo9_2),.clk(gclk));
	jdff dff_B_IPHjuRXg6_2(.din(w_dff_B_QflfAzRo9_2),.dout(w_dff_B_IPHjuRXg6_2),.clk(gclk));
	jdff dff_B_iNBJO3Iw4_2(.din(w_dff_B_IPHjuRXg6_2),.dout(w_dff_B_iNBJO3Iw4_2),.clk(gclk));
	jdff dff_B_p1UJ8gvY2_2(.din(w_dff_B_iNBJO3Iw4_2),.dout(w_dff_B_p1UJ8gvY2_2),.clk(gclk));
	jdff dff_B_A70XKMX65_2(.din(w_dff_B_p1UJ8gvY2_2),.dout(w_dff_B_A70XKMX65_2),.clk(gclk));
	jdff dff_B_xVATjQpv2_2(.din(w_dff_B_A70XKMX65_2),.dout(w_dff_B_xVATjQpv2_2),.clk(gclk));
	jdff dff_B_FfQGHvcz9_2(.din(w_dff_B_xVATjQpv2_2),.dout(w_dff_B_FfQGHvcz9_2),.clk(gclk));
	jdff dff_B_tpDpCILF9_2(.din(w_dff_B_FfQGHvcz9_2),.dout(w_dff_B_tpDpCILF9_2),.clk(gclk));
	jdff dff_B_y7UBxaVe9_2(.din(w_dff_B_tpDpCILF9_2),.dout(w_dff_B_y7UBxaVe9_2),.clk(gclk));
	jdff dff_B_t3zvDPvW5_2(.din(w_dff_B_y7UBxaVe9_2),.dout(w_dff_B_t3zvDPvW5_2),.clk(gclk));
	jdff dff_B_sdIisz9O7_2(.din(w_dff_B_t3zvDPvW5_2),.dout(w_dff_B_sdIisz9O7_2),.clk(gclk));
	jdff dff_B_j20DL4N69_2(.din(w_dff_B_sdIisz9O7_2),.dout(w_dff_B_j20DL4N69_2),.clk(gclk));
	jdff dff_B_8ay992s14_2(.din(w_dff_B_j20DL4N69_2),.dout(w_dff_B_8ay992s14_2),.clk(gclk));
	jdff dff_B_0a14F5911_2(.din(w_dff_B_8ay992s14_2),.dout(w_dff_B_0a14F5911_2),.clk(gclk));
	jdff dff_B_ljbBY7Lj5_2(.din(w_dff_B_0a14F5911_2),.dout(w_dff_B_ljbBY7Lj5_2),.clk(gclk));
	jdff dff_B_vAfuBllz1_2(.din(w_dff_B_ljbBY7Lj5_2),.dout(w_dff_B_vAfuBllz1_2),.clk(gclk));
	jdff dff_B_9R6hN7230_2(.din(w_dff_B_vAfuBllz1_2),.dout(w_dff_B_9R6hN7230_2),.clk(gclk));
	jdff dff_B_6eoxZfhQ4_2(.din(w_dff_B_9R6hN7230_2),.dout(w_dff_B_6eoxZfhQ4_2),.clk(gclk));
	jdff dff_B_6LRWDamo4_2(.din(w_dff_B_6eoxZfhQ4_2),.dout(w_dff_B_6LRWDamo4_2),.clk(gclk));
	jdff dff_B_8fNPFrdf1_2(.din(w_dff_B_6LRWDamo4_2),.dout(w_dff_B_8fNPFrdf1_2),.clk(gclk));
	jdff dff_B_aapST4Cv0_2(.din(w_dff_B_8fNPFrdf1_2),.dout(w_dff_B_aapST4Cv0_2),.clk(gclk));
	jdff dff_B_UJh4Cvpm5_2(.din(w_dff_B_aapST4Cv0_2),.dout(w_dff_B_UJh4Cvpm5_2),.clk(gclk));
	jdff dff_B_3Rj94cVZ0_2(.din(w_dff_B_UJh4Cvpm5_2),.dout(w_dff_B_3Rj94cVZ0_2),.clk(gclk));
	jdff dff_B_xrHz6jpY7_2(.din(w_dff_B_3Rj94cVZ0_2),.dout(w_dff_B_xrHz6jpY7_2),.clk(gclk));
	jdff dff_B_UUKJBab72_2(.din(w_dff_B_xrHz6jpY7_2),.dout(w_dff_B_UUKJBab72_2),.clk(gclk));
	jdff dff_B_bWkcc7Z69_2(.din(w_dff_B_UUKJBab72_2),.dout(w_dff_B_bWkcc7Z69_2),.clk(gclk));
	jdff dff_B_Jayjf1Sp4_2(.din(w_dff_B_bWkcc7Z69_2),.dout(w_dff_B_Jayjf1Sp4_2),.clk(gclk));
	jdff dff_B_okZPYfUy4_1(.din(n1391),.dout(w_dff_B_okZPYfUy4_1),.clk(gclk));
	jdff dff_B_2FHgVOBY5_2(.din(n1312),.dout(w_dff_B_2FHgVOBY5_2),.clk(gclk));
	jdff dff_B_AiUKz9DE9_2(.din(w_dff_B_2FHgVOBY5_2),.dout(w_dff_B_AiUKz9DE9_2),.clk(gclk));
	jdff dff_B_GxH1MmvG7_2(.din(w_dff_B_AiUKz9DE9_2),.dout(w_dff_B_GxH1MmvG7_2),.clk(gclk));
	jdff dff_B_m4tnjpuY3_2(.din(w_dff_B_GxH1MmvG7_2),.dout(w_dff_B_m4tnjpuY3_2),.clk(gclk));
	jdff dff_B_cfai8G0e3_2(.din(w_dff_B_m4tnjpuY3_2),.dout(w_dff_B_cfai8G0e3_2),.clk(gclk));
	jdff dff_B_KKUPwmjX8_2(.din(w_dff_B_cfai8G0e3_2),.dout(w_dff_B_KKUPwmjX8_2),.clk(gclk));
	jdff dff_B_aDOm0Xx91_2(.din(w_dff_B_KKUPwmjX8_2),.dout(w_dff_B_aDOm0Xx91_2),.clk(gclk));
	jdff dff_B_Rj9sCT1D3_2(.din(w_dff_B_aDOm0Xx91_2),.dout(w_dff_B_Rj9sCT1D3_2),.clk(gclk));
	jdff dff_B_CPqFrG2y8_2(.din(w_dff_B_Rj9sCT1D3_2),.dout(w_dff_B_CPqFrG2y8_2),.clk(gclk));
	jdff dff_B_3tQuH77c7_2(.din(w_dff_B_CPqFrG2y8_2),.dout(w_dff_B_3tQuH77c7_2),.clk(gclk));
	jdff dff_B_0e7vG31u5_2(.din(w_dff_B_3tQuH77c7_2),.dout(w_dff_B_0e7vG31u5_2),.clk(gclk));
	jdff dff_B_TdBal9S57_2(.din(w_dff_B_0e7vG31u5_2),.dout(w_dff_B_TdBal9S57_2),.clk(gclk));
	jdff dff_B_ft8Dn88k7_2(.din(w_dff_B_TdBal9S57_2),.dout(w_dff_B_ft8Dn88k7_2),.clk(gclk));
	jdff dff_B_e01OjxXX3_2(.din(w_dff_B_ft8Dn88k7_2),.dout(w_dff_B_e01OjxXX3_2),.clk(gclk));
	jdff dff_B_AW0MOot52_2(.din(w_dff_B_e01OjxXX3_2),.dout(w_dff_B_AW0MOot52_2),.clk(gclk));
	jdff dff_B_jl81WEhp0_2(.din(w_dff_B_AW0MOot52_2),.dout(w_dff_B_jl81WEhp0_2),.clk(gclk));
	jdff dff_B_rBITXdHJ1_2(.din(w_dff_B_jl81WEhp0_2),.dout(w_dff_B_rBITXdHJ1_2),.clk(gclk));
	jdff dff_B_RMp93ep76_2(.din(w_dff_B_rBITXdHJ1_2),.dout(w_dff_B_RMp93ep76_2),.clk(gclk));
	jdff dff_B_Pq315Gmc5_2(.din(w_dff_B_RMp93ep76_2),.dout(w_dff_B_Pq315Gmc5_2),.clk(gclk));
	jdff dff_B_GjW8idSO6_2(.din(w_dff_B_Pq315Gmc5_2),.dout(w_dff_B_GjW8idSO6_2),.clk(gclk));
	jdff dff_B_PcNx6c0N0_2(.din(w_dff_B_GjW8idSO6_2),.dout(w_dff_B_PcNx6c0N0_2),.clk(gclk));
	jdff dff_B_7AyP6H7O7_2(.din(w_dff_B_PcNx6c0N0_2),.dout(w_dff_B_7AyP6H7O7_2),.clk(gclk));
	jdff dff_B_rY2At0qi5_2(.din(w_dff_B_7AyP6H7O7_2),.dout(w_dff_B_rY2At0qi5_2),.clk(gclk));
	jdff dff_B_uQXcYRnD8_2(.din(w_dff_B_rY2At0qi5_2),.dout(w_dff_B_uQXcYRnD8_2),.clk(gclk));
	jdff dff_B_3HOUjZ767_2(.din(w_dff_B_uQXcYRnD8_2),.dout(w_dff_B_3HOUjZ767_2),.clk(gclk));
	jdff dff_B_Q8KQnlZG4_2(.din(w_dff_B_3HOUjZ767_2),.dout(w_dff_B_Q8KQnlZG4_2),.clk(gclk));
	jdff dff_B_BfZmWP7T6_2(.din(w_dff_B_Q8KQnlZG4_2),.dout(w_dff_B_BfZmWP7T6_2),.clk(gclk));
	jdff dff_B_TsQO7Wvf1_2(.din(w_dff_B_BfZmWP7T6_2),.dout(w_dff_B_TsQO7Wvf1_2),.clk(gclk));
	jdff dff_B_zzPrbLCm3_2(.din(w_dff_B_TsQO7Wvf1_2),.dout(w_dff_B_zzPrbLCm3_2),.clk(gclk));
	jdff dff_B_Te1i66hV5_2(.din(w_dff_B_zzPrbLCm3_2),.dout(w_dff_B_Te1i66hV5_2),.clk(gclk));
	jdff dff_B_htUOUhmr2_2(.din(w_dff_B_Te1i66hV5_2),.dout(w_dff_B_htUOUhmr2_2),.clk(gclk));
	jdff dff_B_SvxBL2CX5_2(.din(w_dff_B_htUOUhmr2_2),.dout(w_dff_B_SvxBL2CX5_2),.clk(gclk));
	jdff dff_B_XFH8kGgb9_2(.din(w_dff_B_SvxBL2CX5_2),.dout(w_dff_B_XFH8kGgb9_2),.clk(gclk));
	jdff dff_B_Eat20wwF4_2(.din(w_dff_B_XFH8kGgb9_2),.dout(w_dff_B_Eat20wwF4_2),.clk(gclk));
	jdff dff_B_p53BAToJ1_2(.din(w_dff_B_Eat20wwF4_2),.dout(w_dff_B_p53BAToJ1_2),.clk(gclk));
	jdff dff_B_1If2QCPg3_2(.din(w_dff_B_p53BAToJ1_2),.dout(w_dff_B_1If2QCPg3_2),.clk(gclk));
	jdff dff_B_QzXJUNAG0_2(.din(w_dff_B_1If2QCPg3_2),.dout(w_dff_B_QzXJUNAG0_2),.clk(gclk));
	jdff dff_B_Yt2BTntV6_2(.din(w_dff_B_QzXJUNAG0_2),.dout(w_dff_B_Yt2BTntV6_2),.clk(gclk));
	jdff dff_B_5Tscc3mU5_2(.din(w_dff_B_Yt2BTntV6_2),.dout(w_dff_B_5Tscc3mU5_2),.clk(gclk));
	jdff dff_B_46wlq6IK4_2(.din(w_dff_B_5Tscc3mU5_2),.dout(w_dff_B_46wlq6IK4_2),.clk(gclk));
	jdff dff_B_GkOsAjCA5_1(.din(n1313),.dout(w_dff_B_GkOsAjCA5_1),.clk(gclk));
	jdff dff_B_qCfy96cX7_2(.din(n1227),.dout(w_dff_B_qCfy96cX7_2),.clk(gclk));
	jdff dff_B_qWFkwedW8_2(.din(w_dff_B_qCfy96cX7_2),.dout(w_dff_B_qWFkwedW8_2),.clk(gclk));
	jdff dff_B_ETqTeCqg5_2(.din(w_dff_B_qWFkwedW8_2),.dout(w_dff_B_ETqTeCqg5_2),.clk(gclk));
	jdff dff_B_mrs8oaK01_2(.din(w_dff_B_ETqTeCqg5_2),.dout(w_dff_B_mrs8oaK01_2),.clk(gclk));
	jdff dff_B_Ym8bGeRl2_2(.din(w_dff_B_mrs8oaK01_2),.dout(w_dff_B_Ym8bGeRl2_2),.clk(gclk));
	jdff dff_B_DsylCa3W7_2(.din(w_dff_B_Ym8bGeRl2_2),.dout(w_dff_B_DsylCa3W7_2),.clk(gclk));
	jdff dff_B_ij8RsBNT2_2(.din(w_dff_B_DsylCa3W7_2),.dout(w_dff_B_ij8RsBNT2_2),.clk(gclk));
	jdff dff_B_s822BQXD2_2(.din(w_dff_B_ij8RsBNT2_2),.dout(w_dff_B_s822BQXD2_2),.clk(gclk));
	jdff dff_B_4LJR26Zz4_2(.din(w_dff_B_s822BQXD2_2),.dout(w_dff_B_4LJR26Zz4_2),.clk(gclk));
	jdff dff_B_I8FsOP383_2(.din(w_dff_B_4LJR26Zz4_2),.dout(w_dff_B_I8FsOP383_2),.clk(gclk));
	jdff dff_B_4TyCm9ea4_2(.din(w_dff_B_I8FsOP383_2),.dout(w_dff_B_4TyCm9ea4_2),.clk(gclk));
	jdff dff_B_jNm1oBz20_2(.din(w_dff_B_4TyCm9ea4_2),.dout(w_dff_B_jNm1oBz20_2),.clk(gclk));
	jdff dff_B_yDvWNEvw1_2(.din(w_dff_B_jNm1oBz20_2),.dout(w_dff_B_yDvWNEvw1_2),.clk(gclk));
	jdff dff_B_jQSi0nhl7_2(.din(w_dff_B_yDvWNEvw1_2),.dout(w_dff_B_jQSi0nhl7_2),.clk(gclk));
	jdff dff_B_zYfO4QD10_2(.din(w_dff_B_jQSi0nhl7_2),.dout(w_dff_B_zYfO4QD10_2),.clk(gclk));
	jdff dff_B_npo0KMU07_2(.din(w_dff_B_zYfO4QD10_2),.dout(w_dff_B_npo0KMU07_2),.clk(gclk));
	jdff dff_B_zNGsRY8g2_2(.din(w_dff_B_npo0KMU07_2),.dout(w_dff_B_zNGsRY8g2_2),.clk(gclk));
	jdff dff_B_rm5N9AZt7_2(.din(w_dff_B_zNGsRY8g2_2),.dout(w_dff_B_rm5N9AZt7_2),.clk(gclk));
	jdff dff_B_wgWjRY6A8_2(.din(w_dff_B_rm5N9AZt7_2),.dout(w_dff_B_wgWjRY6A8_2),.clk(gclk));
	jdff dff_B_BOFFIOU05_2(.din(w_dff_B_wgWjRY6A8_2),.dout(w_dff_B_BOFFIOU05_2),.clk(gclk));
	jdff dff_B_Gxmvnb5R5_2(.din(w_dff_B_BOFFIOU05_2),.dout(w_dff_B_Gxmvnb5R5_2),.clk(gclk));
	jdff dff_B_XvF3he9e9_2(.din(w_dff_B_Gxmvnb5R5_2),.dout(w_dff_B_XvF3he9e9_2),.clk(gclk));
	jdff dff_B_3LlcdKAo3_2(.din(w_dff_B_XvF3he9e9_2),.dout(w_dff_B_3LlcdKAo3_2),.clk(gclk));
	jdff dff_B_a6VJsaRx5_2(.din(w_dff_B_3LlcdKAo3_2),.dout(w_dff_B_a6VJsaRx5_2),.clk(gclk));
	jdff dff_B_fj0iVqtX8_2(.din(w_dff_B_a6VJsaRx5_2),.dout(w_dff_B_fj0iVqtX8_2),.clk(gclk));
	jdff dff_B_fhlgibW17_2(.din(w_dff_B_fj0iVqtX8_2),.dout(w_dff_B_fhlgibW17_2),.clk(gclk));
	jdff dff_B_Cp7XneBh6_2(.din(w_dff_B_fhlgibW17_2),.dout(w_dff_B_Cp7XneBh6_2),.clk(gclk));
	jdff dff_B_5IhKFno72_2(.din(w_dff_B_Cp7XneBh6_2),.dout(w_dff_B_5IhKFno72_2),.clk(gclk));
	jdff dff_B_SDTPaPew4_2(.din(w_dff_B_5IhKFno72_2),.dout(w_dff_B_SDTPaPew4_2),.clk(gclk));
	jdff dff_B_LosGJHyD2_2(.din(w_dff_B_SDTPaPew4_2),.dout(w_dff_B_LosGJHyD2_2),.clk(gclk));
	jdff dff_B_olGrOOJb1_2(.din(w_dff_B_LosGJHyD2_2),.dout(w_dff_B_olGrOOJb1_2),.clk(gclk));
	jdff dff_B_2MIsppXc9_2(.din(w_dff_B_olGrOOJb1_2),.dout(w_dff_B_2MIsppXc9_2),.clk(gclk));
	jdff dff_B_t4jWqFVG6_2(.din(w_dff_B_2MIsppXc9_2),.dout(w_dff_B_t4jWqFVG6_2),.clk(gclk));
	jdff dff_B_OZ6qpPTy4_2(.din(w_dff_B_t4jWqFVG6_2),.dout(w_dff_B_OZ6qpPTy4_2),.clk(gclk));
	jdff dff_B_wnkFhy2N6_2(.din(w_dff_B_OZ6qpPTy4_2),.dout(w_dff_B_wnkFhy2N6_2),.clk(gclk));
	jdff dff_B_XlSilwFu7_2(.din(w_dff_B_wnkFhy2N6_2),.dout(w_dff_B_XlSilwFu7_2),.clk(gclk));
	jdff dff_B_yriLKFxM6_2(.din(w_dff_B_XlSilwFu7_2),.dout(w_dff_B_yriLKFxM6_2),.clk(gclk));
	jdff dff_B_eWRukfmw4_1(.din(n1228),.dout(w_dff_B_eWRukfmw4_1),.clk(gclk));
	jdff dff_B_ydnRlVpB3_2(.din(n1136),.dout(w_dff_B_ydnRlVpB3_2),.clk(gclk));
	jdff dff_B_w7fsqj4P0_2(.din(w_dff_B_ydnRlVpB3_2),.dout(w_dff_B_w7fsqj4P0_2),.clk(gclk));
	jdff dff_B_ObquUWuS3_2(.din(w_dff_B_w7fsqj4P0_2),.dout(w_dff_B_ObquUWuS3_2),.clk(gclk));
	jdff dff_B_HB8JQfSM1_2(.din(w_dff_B_ObquUWuS3_2),.dout(w_dff_B_HB8JQfSM1_2),.clk(gclk));
	jdff dff_B_F02MSOvL3_2(.din(w_dff_B_HB8JQfSM1_2),.dout(w_dff_B_F02MSOvL3_2),.clk(gclk));
	jdff dff_B_FGbvqy2Q7_2(.din(w_dff_B_F02MSOvL3_2),.dout(w_dff_B_FGbvqy2Q7_2),.clk(gclk));
	jdff dff_B_QQupTRmD1_2(.din(w_dff_B_FGbvqy2Q7_2),.dout(w_dff_B_QQupTRmD1_2),.clk(gclk));
	jdff dff_B_71fpE7MR4_2(.din(w_dff_B_QQupTRmD1_2),.dout(w_dff_B_71fpE7MR4_2),.clk(gclk));
	jdff dff_B_NauiZ4Fy0_2(.din(w_dff_B_71fpE7MR4_2),.dout(w_dff_B_NauiZ4Fy0_2),.clk(gclk));
	jdff dff_B_RX9WqM9h0_2(.din(w_dff_B_NauiZ4Fy0_2),.dout(w_dff_B_RX9WqM9h0_2),.clk(gclk));
	jdff dff_B_XI0Fftw28_2(.din(w_dff_B_RX9WqM9h0_2),.dout(w_dff_B_XI0Fftw28_2),.clk(gclk));
	jdff dff_B_JPYRxwGb9_2(.din(w_dff_B_XI0Fftw28_2),.dout(w_dff_B_JPYRxwGb9_2),.clk(gclk));
	jdff dff_B_5PY4syl25_2(.din(w_dff_B_JPYRxwGb9_2),.dout(w_dff_B_5PY4syl25_2),.clk(gclk));
	jdff dff_B_rM1B12IR7_2(.din(w_dff_B_5PY4syl25_2),.dout(w_dff_B_rM1B12IR7_2),.clk(gclk));
	jdff dff_B_kzbweZEn4_2(.din(w_dff_B_rM1B12IR7_2),.dout(w_dff_B_kzbweZEn4_2),.clk(gclk));
	jdff dff_B_hPe3EIBr9_2(.din(w_dff_B_kzbweZEn4_2),.dout(w_dff_B_hPe3EIBr9_2),.clk(gclk));
	jdff dff_B_jlKiSpEy3_2(.din(w_dff_B_hPe3EIBr9_2),.dout(w_dff_B_jlKiSpEy3_2),.clk(gclk));
	jdff dff_B_SvRxmqY43_2(.din(w_dff_B_jlKiSpEy3_2),.dout(w_dff_B_SvRxmqY43_2),.clk(gclk));
	jdff dff_B_sVpnHyj48_2(.din(w_dff_B_SvRxmqY43_2),.dout(w_dff_B_sVpnHyj48_2),.clk(gclk));
	jdff dff_B_ZtETKS3z6_2(.din(w_dff_B_sVpnHyj48_2),.dout(w_dff_B_ZtETKS3z6_2),.clk(gclk));
	jdff dff_B_moEckjPF2_2(.din(w_dff_B_ZtETKS3z6_2),.dout(w_dff_B_moEckjPF2_2),.clk(gclk));
	jdff dff_B_go3ZHA9c7_2(.din(w_dff_B_moEckjPF2_2),.dout(w_dff_B_go3ZHA9c7_2),.clk(gclk));
	jdff dff_B_nbiclrTt7_2(.din(w_dff_B_go3ZHA9c7_2),.dout(w_dff_B_nbiclrTt7_2),.clk(gclk));
	jdff dff_B_ZGsriYPt7_2(.din(w_dff_B_nbiclrTt7_2),.dout(w_dff_B_ZGsriYPt7_2),.clk(gclk));
	jdff dff_B_H2jBMIvq9_2(.din(w_dff_B_ZGsriYPt7_2),.dout(w_dff_B_H2jBMIvq9_2),.clk(gclk));
	jdff dff_B_RGsD2Ahi9_2(.din(w_dff_B_H2jBMIvq9_2),.dout(w_dff_B_RGsD2Ahi9_2),.clk(gclk));
	jdff dff_B_3h3hCPL00_2(.din(w_dff_B_RGsD2Ahi9_2),.dout(w_dff_B_3h3hCPL00_2),.clk(gclk));
	jdff dff_B_MAN844QY8_2(.din(w_dff_B_3h3hCPL00_2),.dout(w_dff_B_MAN844QY8_2),.clk(gclk));
	jdff dff_B_iHtcMqOh4_2(.din(w_dff_B_MAN844QY8_2),.dout(w_dff_B_iHtcMqOh4_2),.clk(gclk));
	jdff dff_B_KCXcFZxf4_2(.din(w_dff_B_iHtcMqOh4_2),.dout(w_dff_B_KCXcFZxf4_2),.clk(gclk));
	jdff dff_B_Ba1c2bqR6_2(.din(w_dff_B_KCXcFZxf4_2),.dout(w_dff_B_Ba1c2bqR6_2),.clk(gclk));
	jdff dff_B_nAh4pjQW7_2(.din(w_dff_B_Ba1c2bqR6_2),.dout(w_dff_B_nAh4pjQW7_2),.clk(gclk));
	jdff dff_B_L0ho2uIT0_2(.din(w_dff_B_nAh4pjQW7_2),.dout(w_dff_B_L0ho2uIT0_2),.clk(gclk));
	jdff dff_B_2vJ0ECc04_2(.din(w_dff_B_L0ho2uIT0_2),.dout(w_dff_B_2vJ0ECc04_2),.clk(gclk));
	jdff dff_B_FmIUrn9u6_1(.din(n1137),.dout(w_dff_B_FmIUrn9u6_1),.clk(gclk));
	jdff dff_B_YhOheFMg0_2(.din(n1038),.dout(w_dff_B_YhOheFMg0_2),.clk(gclk));
	jdff dff_B_5cIrRVT33_2(.din(w_dff_B_YhOheFMg0_2),.dout(w_dff_B_5cIrRVT33_2),.clk(gclk));
	jdff dff_B_kOYBXiHE9_2(.din(w_dff_B_5cIrRVT33_2),.dout(w_dff_B_kOYBXiHE9_2),.clk(gclk));
	jdff dff_B_M6Wwa9E80_2(.din(w_dff_B_kOYBXiHE9_2),.dout(w_dff_B_M6Wwa9E80_2),.clk(gclk));
	jdff dff_B_IbJm1Q2G1_2(.din(w_dff_B_M6Wwa9E80_2),.dout(w_dff_B_IbJm1Q2G1_2),.clk(gclk));
	jdff dff_B_o65yV4W44_2(.din(w_dff_B_IbJm1Q2G1_2),.dout(w_dff_B_o65yV4W44_2),.clk(gclk));
	jdff dff_B_oq3h95fv5_2(.din(w_dff_B_o65yV4W44_2),.dout(w_dff_B_oq3h95fv5_2),.clk(gclk));
	jdff dff_B_YPRjFFTg2_2(.din(w_dff_B_oq3h95fv5_2),.dout(w_dff_B_YPRjFFTg2_2),.clk(gclk));
	jdff dff_B_9jWxiIwf0_2(.din(w_dff_B_YPRjFFTg2_2),.dout(w_dff_B_9jWxiIwf0_2),.clk(gclk));
	jdff dff_B_9oihohtO2_2(.din(w_dff_B_9jWxiIwf0_2),.dout(w_dff_B_9oihohtO2_2),.clk(gclk));
	jdff dff_B_3L40jCqf7_2(.din(w_dff_B_9oihohtO2_2),.dout(w_dff_B_3L40jCqf7_2),.clk(gclk));
	jdff dff_B_zL8YWxPk1_2(.din(w_dff_B_3L40jCqf7_2),.dout(w_dff_B_zL8YWxPk1_2),.clk(gclk));
	jdff dff_B_5xWILhr79_2(.din(w_dff_B_zL8YWxPk1_2),.dout(w_dff_B_5xWILhr79_2),.clk(gclk));
	jdff dff_B_gRWqRPTD8_2(.din(w_dff_B_5xWILhr79_2),.dout(w_dff_B_gRWqRPTD8_2),.clk(gclk));
	jdff dff_B_Xvrm9jtV6_2(.din(w_dff_B_gRWqRPTD8_2),.dout(w_dff_B_Xvrm9jtV6_2),.clk(gclk));
	jdff dff_B_M2GUvrHP8_2(.din(w_dff_B_Xvrm9jtV6_2),.dout(w_dff_B_M2GUvrHP8_2),.clk(gclk));
	jdff dff_B_ezwzdqy06_2(.din(w_dff_B_M2GUvrHP8_2),.dout(w_dff_B_ezwzdqy06_2),.clk(gclk));
	jdff dff_B_UTwgntyC9_2(.din(w_dff_B_ezwzdqy06_2),.dout(w_dff_B_UTwgntyC9_2),.clk(gclk));
	jdff dff_B_SyqnNlG53_2(.din(w_dff_B_UTwgntyC9_2),.dout(w_dff_B_SyqnNlG53_2),.clk(gclk));
	jdff dff_B_dXG8MYI47_2(.din(w_dff_B_SyqnNlG53_2),.dout(w_dff_B_dXG8MYI47_2),.clk(gclk));
	jdff dff_B_bivUJdQg9_2(.din(w_dff_B_dXG8MYI47_2),.dout(w_dff_B_bivUJdQg9_2),.clk(gclk));
	jdff dff_B_0hyWc2yJ5_2(.din(w_dff_B_bivUJdQg9_2),.dout(w_dff_B_0hyWc2yJ5_2),.clk(gclk));
	jdff dff_B_YkUMhdsQ6_2(.din(w_dff_B_0hyWc2yJ5_2),.dout(w_dff_B_YkUMhdsQ6_2),.clk(gclk));
	jdff dff_B_ALrXiQfO9_2(.din(w_dff_B_YkUMhdsQ6_2),.dout(w_dff_B_ALrXiQfO9_2),.clk(gclk));
	jdff dff_B_3o62TwvU7_2(.din(w_dff_B_ALrXiQfO9_2),.dout(w_dff_B_3o62TwvU7_2),.clk(gclk));
	jdff dff_B_hv9kSpGt7_2(.din(w_dff_B_3o62TwvU7_2),.dout(w_dff_B_hv9kSpGt7_2),.clk(gclk));
	jdff dff_B_Cl89ITno8_2(.din(w_dff_B_hv9kSpGt7_2),.dout(w_dff_B_Cl89ITno8_2),.clk(gclk));
	jdff dff_B_bvYFSfcm1_2(.din(w_dff_B_Cl89ITno8_2),.dout(w_dff_B_bvYFSfcm1_2),.clk(gclk));
	jdff dff_B_4xLBcRnD9_2(.din(w_dff_B_bvYFSfcm1_2),.dout(w_dff_B_4xLBcRnD9_2),.clk(gclk));
	jdff dff_B_pMWVECVB6_2(.din(w_dff_B_4xLBcRnD9_2),.dout(w_dff_B_pMWVECVB6_2),.clk(gclk));
	jdff dff_B_UImGPrEg1_2(.din(w_dff_B_pMWVECVB6_2),.dout(w_dff_B_UImGPrEg1_2),.clk(gclk));
	jdff dff_B_X9x5eONG1_1(.din(n1039),.dout(w_dff_B_X9x5eONG1_1),.clk(gclk));
	jdff dff_B_lfBrzUrz6_2(.din(n939),.dout(w_dff_B_lfBrzUrz6_2),.clk(gclk));
	jdff dff_B_I4gDPI392_2(.din(w_dff_B_lfBrzUrz6_2),.dout(w_dff_B_I4gDPI392_2),.clk(gclk));
	jdff dff_B_BYaGUQBu7_2(.din(w_dff_B_I4gDPI392_2),.dout(w_dff_B_BYaGUQBu7_2),.clk(gclk));
	jdff dff_B_4SEIkHOT4_2(.din(w_dff_B_BYaGUQBu7_2),.dout(w_dff_B_4SEIkHOT4_2),.clk(gclk));
	jdff dff_B_FoWaM2DB1_2(.din(w_dff_B_4SEIkHOT4_2),.dout(w_dff_B_FoWaM2DB1_2),.clk(gclk));
	jdff dff_B_vtqDLHrl3_2(.din(w_dff_B_FoWaM2DB1_2),.dout(w_dff_B_vtqDLHrl3_2),.clk(gclk));
	jdff dff_B_qlO9WPcz7_2(.din(w_dff_B_vtqDLHrl3_2),.dout(w_dff_B_qlO9WPcz7_2),.clk(gclk));
	jdff dff_B_Gv3WRA0O5_2(.din(w_dff_B_qlO9WPcz7_2),.dout(w_dff_B_Gv3WRA0O5_2),.clk(gclk));
	jdff dff_B_Hym1lT2v2_2(.din(w_dff_B_Gv3WRA0O5_2),.dout(w_dff_B_Hym1lT2v2_2),.clk(gclk));
	jdff dff_B_QnELvtVC3_2(.din(w_dff_B_Hym1lT2v2_2),.dout(w_dff_B_QnELvtVC3_2),.clk(gclk));
	jdff dff_B_z5fmOBeh4_2(.din(w_dff_B_QnELvtVC3_2),.dout(w_dff_B_z5fmOBeh4_2),.clk(gclk));
	jdff dff_B_xfTH8nsm5_2(.din(w_dff_B_z5fmOBeh4_2),.dout(w_dff_B_xfTH8nsm5_2),.clk(gclk));
	jdff dff_B_PwRJ4YaM8_2(.din(w_dff_B_xfTH8nsm5_2),.dout(w_dff_B_PwRJ4YaM8_2),.clk(gclk));
	jdff dff_B_VIYUXkdD6_2(.din(w_dff_B_PwRJ4YaM8_2),.dout(w_dff_B_VIYUXkdD6_2),.clk(gclk));
	jdff dff_B_c2ygEIGp6_2(.din(w_dff_B_VIYUXkdD6_2),.dout(w_dff_B_c2ygEIGp6_2),.clk(gclk));
	jdff dff_B_8K4SJKp38_2(.din(w_dff_B_c2ygEIGp6_2),.dout(w_dff_B_8K4SJKp38_2),.clk(gclk));
	jdff dff_B_8WTgtnfC7_2(.din(w_dff_B_8K4SJKp38_2),.dout(w_dff_B_8WTgtnfC7_2),.clk(gclk));
	jdff dff_B_URCHDs8v9_2(.din(w_dff_B_8WTgtnfC7_2),.dout(w_dff_B_URCHDs8v9_2),.clk(gclk));
	jdff dff_B_y35Sv2AP7_2(.din(w_dff_B_URCHDs8v9_2),.dout(w_dff_B_y35Sv2AP7_2),.clk(gclk));
	jdff dff_B_Oyr3oh2T5_2(.din(w_dff_B_y35Sv2AP7_2),.dout(w_dff_B_Oyr3oh2T5_2),.clk(gclk));
	jdff dff_B_kj4TQQJI6_2(.din(w_dff_B_Oyr3oh2T5_2),.dout(w_dff_B_kj4TQQJI6_2),.clk(gclk));
	jdff dff_B_U5nNO81N0_2(.din(w_dff_B_kj4TQQJI6_2),.dout(w_dff_B_U5nNO81N0_2),.clk(gclk));
	jdff dff_B_W06xmaZP0_2(.din(w_dff_B_U5nNO81N0_2),.dout(w_dff_B_W06xmaZP0_2),.clk(gclk));
	jdff dff_B_gq6YKjlZ3_2(.din(w_dff_B_W06xmaZP0_2),.dout(w_dff_B_gq6YKjlZ3_2),.clk(gclk));
	jdff dff_B_bm1ZlNgl4_2(.din(w_dff_B_gq6YKjlZ3_2),.dout(w_dff_B_bm1ZlNgl4_2),.clk(gclk));
	jdff dff_B_HD6R4fCa1_2(.din(w_dff_B_bm1ZlNgl4_2),.dout(w_dff_B_HD6R4fCa1_2),.clk(gclk));
	jdff dff_B_GZNE8dma7_2(.din(w_dff_B_HD6R4fCa1_2),.dout(w_dff_B_GZNE8dma7_2),.clk(gclk));
	jdff dff_B_VDExURbU0_2(.din(w_dff_B_GZNE8dma7_2),.dout(w_dff_B_VDExURbU0_2),.clk(gclk));
	jdff dff_B_70voapNf1_1(.din(n940),.dout(w_dff_B_70voapNf1_1),.clk(gclk));
	jdff dff_B_TnajQOjF5_2(.din(n837),.dout(w_dff_B_TnajQOjF5_2),.clk(gclk));
	jdff dff_B_nX7Vn4xJ0_2(.din(w_dff_B_TnajQOjF5_2),.dout(w_dff_B_nX7Vn4xJ0_2),.clk(gclk));
	jdff dff_B_T0Uzh5Y36_2(.din(w_dff_B_nX7Vn4xJ0_2),.dout(w_dff_B_T0Uzh5Y36_2),.clk(gclk));
	jdff dff_B_x0u8nhnw7_2(.din(w_dff_B_T0Uzh5Y36_2),.dout(w_dff_B_x0u8nhnw7_2),.clk(gclk));
	jdff dff_B_jaIlhc4N4_2(.din(w_dff_B_x0u8nhnw7_2),.dout(w_dff_B_jaIlhc4N4_2),.clk(gclk));
	jdff dff_B_e4TP2vWq7_2(.din(w_dff_B_jaIlhc4N4_2),.dout(w_dff_B_e4TP2vWq7_2),.clk(gclk));
	jdff dff_B_nxV8kibe6_2(.din(w_dff_B_e4TP2vWq7_2),.dout(w_dff_B_nxV8kibe6_2),.clk(gclk));
	jdff dff_B_c0u3t53e8_2(.din(w_dff_B_nxV8kibe6_2),.dout(w_dff_B_c0u3t53e8_2),.clk(gclk));
	jdff dff_B_PIbZcqUT2_2(.din(w_dff_B_c0u3t53e8_2),.dout(w_dff_B_PIbZcqUT2_2),.clk(gclk));
	jdff dff_B_91UUNVtU3_2(.din(w_dff_B_PIbZcqUT2_2),.dout(w_dff_B_91UUNVtU3_2),.clk(gclk));
	jdff dff_B_wFMIMidM1_2(.din(w_dff_B_91UUNVtU3_2),.dout(w_dff_B_wFMIMidM1_2),.clk(gclk));
	jdff dff_B_8t7O4wBV8_2(.din(w_dff_B_wFMIMidM1_2),.dout(w_dff_B_8t7O4wBV8_2),.clk(gclk));
	jdff dff_B_tRlUm20j6_2(.din(w_dff_B_8t7O4wBV8_2),.dout(w_dff_B_tRlUm20j6_2),.clk(gclk));
	jdff dff_B_QyVkVUSp4_2(.din(w_dff_B_tRlUm20j6_2),.dout(w_dff_B_QyVkVUSp4_2),.clk(gclk));
	jdff dff_B_YymKICMc9_2(.din(w_dff_B_QyVkVUSp4_2),.dout(w_dff_B_YymKICMc9_2),.clk(gclk));
	jdff dff_B_aCMHH9qC4_2(.din(w_dff_B_YymKICMc9_2),.dout(w_dff_B_aCMHH9qC4_2),.clk(gclk));
	jdff dff_B_hwY2v7cA7_2(.din(w_dff_B_aCMHH9qC4_2),.dout(w_dff_B_hwY2v7cA7_2),.clk(gclk));
	jdff dff_B_vVhDKRVx4_2(.din(w_dff_B_hwY2v7cA7_2),.dout(w_dff_B_vVhDKRVx4_2),.clk(gclk));
	jdff dff_B_6WwIKGxL4_2(.din(w_dff_B_vVhDKRVx4_2),.dout(w_dff_B_6WwIKGxL4_2),.clk(gclk));
	jdff dff_B_TRxvA4oM1_2(.din(w_dff_B_6WwIKGxL4_2),.dout(w_dff_B_TRxvA4oM1_2),.clk(gclk));
	jdff dff_B_QFo2R29W7_2(.din(w_dff_B_TRxvA4oM1_2),.dout(w_dff_B_QFo2R29W7_2),.clk(gclk));
	jdff dff_B_lWDsRKFF7_2(.din(w_dff_B_QFo2R29W7_2),.dout(w_dff_B_lWDsRKFF7_2),.clk(gclk));
	jdff dff_B_Wa67a40Z2_2(.din(w_dff_B_lWDsRKFF7_2),.dout(w_dff_B_Wa67a40Z2_2),.clk(gclk));
	jdff dff_B_2mA5JmjA2_2(.din(w_dff_B_Wa67a40Z2_2),.dout(w_dff_B_2mA5JmjA2_2),.clk(gclk));
	jdff dff_B_5ffPzOR82_2(.din(w_dff_B_2mA5JmjA2_2),.dout(w_dff_B_5ffPzOR82_2),.clk(gclk));
	jdff dff_B_AojH413d8_1(.din(n838),.dout(w_dff_B_AojH413d8_1),.clk(gclk));
	jdff dff_B_bojL8AXu1_2(.din(n739),.dout(w_dff_B_bojL8AXu1_2),.clk(gclk));
	jdff dff_B_SFc7Rnd68_2(.din(w_dff_B_bojL8AXu1_2),.dout(w_dff_B_SFc7Rnd68_2),.clk(gclk));
	jdff dff_B_UEQUFxnz8_2(.din(w_dff_B_SFc7Rnd68_2),.dout(w_dff_B_UEQUFxnz8_2),.clk(gclk));
	jdff dff_B_5pgdEYHc1_2(.din(w_dff_B_UEQUFxnz8_2),.dout(w_dff_B_5pgdEYHc1_2),.clk(gclk));
	jdff dff_B_Ek4SrkcL4_2(.din(w_dff_B_5pgdEYHc1_2),.dout(w_dff_B_Ek4SrkcL4_2),.clk(gclk));
	jdff dff_B_Ykuj1MrY5_2(.din(w_dff_B_Ek4SrkcL4_2),.dout(w_dff_B_Ykuj1MrY5_2),.clk(gclk));
	jdff dff_B_Z8op9tpd0_2(.din(w_dff_B_Ykuj1MrY5_2),.dout(w_dff_B_Z8op9tpd0_2),.clk(gclk));
	jdff dff_B_5E3MbnFt2_2(.din(w_dff_B_Z8op9tpd0_2),.dout(w_dff_B_5E3MbnFt2_2),.clk(gclk));
	jdff dff_B_WVyxDF8I4_2(.din(w_dff_B_5E3MbnFt2_2),.dout(w_dff_B_WVyxDF8I4_2),.clk(gclk));
	jdff dff_B_b1NwTAOJ4_2(.din(w_dff_B_WVyxDF8I4_2),.dout(w_dff_B_b1NwTAOJ4_2),.clk(gclk));
	jdff dff_B_lNHeQRKb6_2(.din(w_dff_B_b1NwTAOJ4_2),.dout(w_dff_B_lNHeQRKb6_2),.clk(gclk));
	jdff dff_B_VAyTxHL41_2(.din(w_dff_B_lNHeQRKb6_2),.dout(w_dff_B_VAyTxHL41_2),.clk(gclk));
	jdff dff_B_fTBCHUgh1_2(.din(w_dff_B_VAyTxHL41_2),.dout(w_dff_B_fTBCHUgh1_2),.clk(gclk));
	jdff dff_B_DQMvKJ7t2_2(.din(w_dff_B_fTBCHUgh1_2),.dout(w_dff_B_DQMvKJ7t2_2),.clk(gclk));
	jdff dff_B_g8yulbvU8_2(.din(w_dff_B_DQMvKJ7t2_2),.dout(w_dff_B_g8yulbvU8_2),.clk(gclk));
	jdff dff_B_H6I1go5J2_2(.din(w_dff_B_g8yulbvU8_2),.dout(w_dff_B_H6I1go5J2_2),.clk(gclk));
	jdff dff_B_DWQ0Z7NF1_2(.din(w_dff_B_H6I1go5J2_2),.dout(w_dff_B_DWQ0Z7NF1_2),.clk(gclk));
	jdff dff_B_3naLMSS43_2(.din(w_dff_B_DWQ0Z7NF1_2),.dout(w_dff_B_3naLMSS43_2),.clk(gclk));
	jdff dff_B_LKYOLMbw2_2(.din(w_dff_B_3naLMSS43_2),.dout(w_dff_B_LKYOLMbw2_2),.clk(gclk));
	jdff dff_B_Xe8hfpQ35_2(.din(w_dff_B_LKYOLMbw2_2),.dout(w_dff_B_Xe8hfpQ35_2),.clk(gclk));
	jdff dff_B_djo0VUY31_2(.din(w_dff_B_Xe8hfpQ35_2),.dout(w_dff_B_djo0VUY31_2),.clk(gclk));
	jdff dff_B_IUpPIGVx7_2(.din(w_dff_B_djo0VUY31_2),.dout(w_dff_B_IUpPIGVx7_2),.clk(gclk));
	jdff dff_B_fmHAL9ae8_1(.din(n740),.dout(w_dff_B_fmHAL9ae8_1),.clk(gclk));
	jdff dff_B_p0tE444d6_2(.din(n647),.dout(w_dff_B_p0tE444d6_2),.clk(gclk));
	jdff dff_B_K7UTe42L6_2(.din(w_dff_B_p0tE444d6_2),.dout(w_dff_B_K7UTe42L6_2),.clk(gclk));
	jdff dff_B_usZ9fHwx7_2(.din(w_dff_B_K7UTe42L6_2),.dout(w_dff_B_usZ9fHwx7_2),.clk(gclk));
	jdff dff_B_CbklaxfM4_2(.din(w_dff_B_usZ9fHwx7_2),.dout(w_dff_B_CbklaxfM4_2),.clk(gclk));
	jdff dff_B_nYoSMv0S4_2(.din(w_dff_B_CbklaxfM4_2),.dout(w_dff_B_nYoSMv0S4_2),.clk(gclk));
	jdff dff_B_Y01bI1t40_2(.din(w_dff_B_nYoSMv0S4_2),.dout(w_dff_B_Y01bI1t40_2),.clk(gclk));
	jdff dff_B_lyYWGvSQ6_2(.din(w_dff_B_Y01bI1t40_2),.dout(w_dff_B_lyYWGvSQ6_2),.clk(gclk));
	jdff dff_B_SpMFarON3_2(.din(w_dff_B_lyYWGvSQ6_2),.dout(w_dff_B_SpMFarON3_2),.clk(gclk));
	jdff dff_B_wHlfpW2R6_2(.din(w_dff_B_SpMFarON3_2),.dout(w_dff_B_wHlfpW2R6_2),.clk(gclk));
	jdff dff_B_2SCrIjwV1_2(.din(w_dff_B_wHlfpW2R6_2),.dout(w_dff_B_2SCrIjwV1_2),.clk(gclk));
	jdff dff_B_DAxOj5kw2_2(.din(w_dff_B_2SCrIjwV1_2),.dout(w_dff_B_DAxOj5kw2_2),.clk(gclk));
	jdff dff_B_F5LGktB03_2(.din(w_dff_B_DAxOj5kw2_2),.dout(w_dff_B_F5LGktB03_2),.clk(gclk));
	jdff dff_B_dL8pwDjZ5_2(.din(w_dff_B_F5LGktB03_2),.dout(w_dff_B_dL8pwDjZ5_2),.clk(gclk));
	jdff dff_B_4125E9pF6_2(.din(w_dff_B_dL8pwDjZ5_2),.dout(w_dff_B_4125E9pF6_2),.clk(gclk));
	jdff dff_B_ouX0EVPl2_2(.din(w_dff_B_4125E9pF6_2),.dout(w_dff_B_ouX0EVPl2_2),.clk(gclk));
	jdff dff_B_cMnm8UwX8_2(.din(w_dff_B_ouX0EVPl2_2),.dout(w_dff_B_cMnm8UwX8_2),.clk(gclk));
	jdff dff_B_YZicZTeH6_2(.din(w_dff_B_cMnm8UwX8_2),.dout(w_dff_B_YZicZTeH6_2),.clk(gclk));
	jdff dff_B_JOVUyAjR9_2(.din(w_dff_B_YZicZTeH6_2),.dout(w_dff_B_JOVUyAjR9_2),.clk(gclk));
	jdff dff_B_XIqTUG0R2_2(.din(w_dff_B_JOVUyAjR9_2),.dout(w_dff_B_XIqTUG0R2_2),.clk(gclk));
	jdff dff_B_C3gKgd3D9_1(.din(n648),.dout(w_dff_B_C3gKgd3D9_1),.clk(gclk));
	jdff dff_B_UIQ4Tq8K0_2(.din(n562),.dout(w_dff_B_UIQ4Tq8K0_2),.clk(gclk));
	jdff dff_B_xZKQC6Z66_2(.din(w_dff_B_UIQ4Tq8K0_2),.dout(w_dff_B_xZKQC6Z66_2),.clk(gclk));
	jdff dff_B_lNb5zbNw0_2(.din(w_dff_B_xZKQC6Z66_2),.dout(w_dff_B_lNb5zbNw0_2),.clk(gclk));
	jdff dff_B_ga64F56D5_2(.din(w_dff_B_lNb5zbNw0_2),.dout(w_dff_B_ga64F56D5_2),.clk(gclk));
	jdff dff_B_d7xdTB787_2(.din(w_dff_B_ga64F56D5_2),.dout(w_dff_B_d7xdTB787_2),.clk(gclk));
	jdff dff_B_2feWtac50_2(.din(w_dff_B_d7xdTB787_2),.dout(w_dff_B_2feWtac50_2),.clk(gclk));
	jdff dff_B_WQK4Y9oX0_2(.din(w_dff_B_2feWtac50_2),.dout(w_dff_B_WQK4Y9oX0_2),.clk(gclk));
	jdff dff_B_Yk8M5kI21_2(.din(w_dff_B_WQK4Y9oX0_2),.dout(w_dff_B_Yk8M5kI21_2),.clk(gclk));
	jdff dff_B_f4xQt3x57_2(.din(w_dff_B_Yk8M5kI21_2),.dout(w_dff_B_f4xQt3x57_2),.clk(gclk));
	jdff dff_B_eYPa24kv9_2(.din(w_dff_B_f4xQt3x57_2),.dout(w_dff_B_eYPa24kv9_2),.clk(gclk));
	jdff dff_B_5xrQ4LJY0_2(.din(w_dff_B_eYPa24kv9_2),.dout(w_dff_B_5xrQ4LJY0_2),.clk(gclk));
	jdff dff_B_fErRU8Wa4_2(.din(w_dff_B_5xrQ4LJY0_2),.dout(w_dff_B_fErRU8Wa4_2),.clk(gclk));
	jdff dff_B_Bd6Lq7wK7_2(.din(w_dff_B_fErRU8Wa4_2),.dout(w_dff_B_Bd6Lq7wK7_2),.clk(gclk));
	jdff dff_B_x36fGRs87_2(.din(w_dff_B_Bd6Lq7wK7_2),.dout(w_dff_B_x36fGRs87_2),.clk(gclk));
	jdff dff_B_D8eIa9Ef0_2(.din(w_dff_B_x36fGRs87_2),.dout(w_dff_B_D8eIa9Ef0_2),.clk(gclk));
	jdff dff_B_uF078E1D9_2(.din(w_dff_B_D8eIa9Ef0_2),.dout(w_dff_B_uF078E1D9_2),.clk(gclk));
	jdff dff_B_sw5cd2Qe4_1(.din(n563),.dout(w_dff_B_sw5cd2Qe4_1),.clk(gclk));
	jdff dff_B_FGIlsyaX8_2(.din(n484),.dout(w_dff_B_FGIlsyaX8_2),.clk(gclk));
	jdff dff_B_n0mfdLxC7_2(.din(w_dff_B_FGIlsyaX8_2),.dout(w_dff_B_n0mfdLxC7_2),.clk(gclk));
	jdff dff_B_62jIwzj55_2(.din(w_dff_B_n0mfdLxC7_2),.dout(w_dff_B_62jIwzj55_2),.clk(gclk));
	jdff dff_B_XhVzmfEv7_2(.din(w_dff_B_62jIwzj55_2),.dout(w_dff_B_XhVzmfEv7_2),.clk(gclk));
	jdff dff_B_5eJCXF1s5_2(.din(w_dff_B_XhVzmfEv7_2),.dout(w_dff_B_5eJCXF1s5_2),.clk(gclk));
	jdff dff_B_NOQRRBaB4_2(.din(w_dff_B_5eJCXF1s5_2),.dout(w_dff_B_NOQRRBaB4_2),.clk(gclk));
	jdff dff_B_kHeG3J936_2(.din(w_dff_B_NOQRRBaB4_2),.dout(w_dff_B_kHeG3J936_2),.clk(gclk));
	jdff dff_B_YZ9xqlzj5_2(.din(w_dff_B_kHeG3J936_2),.dout(w_dff_B_YZ9xqlzj5_2),.clk(gclk));
	jdff dff_B_iHiiKhso8_2(.din(w_dff_B_YZ9xqlzj5_2),.dout(w_dff_B_iHiiKhso8_2),.clk(gclk));
	jdff dff_B_1lthIbJN1_2(.din(w_dff_B_iHiiKhso8_2),.dout(w_dff_B_1lthIbJN1_2),.clk(gclk));
	jdff dff_B_ZEY1crJr7_2(.din(w_dff_B_1lthIbJN1_2),.dout(w_dff_B_ZEY1crJr7_2),.clk(gclk));
	jdff dff_B_54IVPH8S9_2(.din(w_dff_B_ZEY1crJr7_2),.dout(w_dff_B_54IVPH8S9_2),.clk(gclk));
	jdff dff_B_jEXVVydu5_2(.din(w_dff_B_54IVPH8S9_2),.dout(w_dff_B_jEXVVydu5_2),.clk(gclk));
	jdff dff_B_w72PYw6U1_1(.din(n485),.dout(w_dff_B_w72PYw6U1_1),.clk(gclk));
	jdff dff_B_GVirOKkz8_2(.din(n413),.dout(w_dff_B_GVirOKkz8_2),.clk(gclk));
	jdff dff_B_8VwgNTfV6_2(.din(w_dff_B_GVirOKkz8_2),.dout(w_dff_B_8VwgNTfV6_2),.clk(gclk));
	jdff dff_B_LGWtgeBN4_2(.din(w_dff_B_8VwgNTfV6_2),.dout(w_dff_B_LGWtgeBN4_2),.clk(gclk));
	jdff dff_B_p1Qsan2p5_2(.din(w_dff_B_LGWtgeBN4_2),.dout(w_dff_B_p1Qsan2p5_2),.clk(gclk));
	jdff dff_B_KAxhzIm75_2(.din(w_dff_B_p1Qsan2p5_2),.dout(w_dff_B_KAxhzIm75_2),.clk(gclk));
	jdff dff_B_FNNwejJq3_2(.din(w_dff_B_KAxhzIm75_2),.dout(w_dff_B_FNNwejJq3_2),.clk(gclk));
	jdff dff_B_BMlDPU3H2_2(.din(w_dff_B_FNNwejJq3_2),.dout(w_dff_B_BMlDPU3H2_2),.clk(gclk));
	jdff dff_B_j38HnXvi8_2(.din(w_dff_B_BMlDPU3H2_2),.dout(w_dff_B_j38HnXvi8_2),.clk(gclk));
	jdff dff_B_LmNVtie13_2(.din(w_dff_B_j38HnXvi8_2),.dout(w_dff_B_LmNVtie13_2),.clk(gclk));
	jdff dff_B_LCG7Dk6n8_2(.din(w_dff_B_LmNVtie13_2),.dout(w_dff_B_LCG7Dk6n8_2),.clk(gclk));
	jdff dff_B_JyHIx9uu1_2(.din(n416),.dout(w_dff_B_JyHIx9uu1_2),.clk(gclk));
	jdff dff_B_thuy0MMT4_1(.din(n414),.dout(w_dff_B_thuy0MMT4_1),.clk(gclk));
	jdff dff_B_ljJHdLN36_2(.din(n350),.dout(w_dff_B_ljJHdLN36_2),.clk(gclk));
	jdff dff_B_h6o6Ds5F7_2(.din(w_dff_B_ljJHdLN36_2),.dout(w_dff_B_h6o6Ds5F7_2),.clk(gclk));
	jdff dff_B_YtVsayaB5_2(.din(w_dff_B_h6o6Ds5F7_2),.dout(w_dff_B_YtVsayaB5_2),.clk(gclk));
	jdff dff_B_cjpEUtrF4_2(.din(w_dff_B_YtVsayaB5_2),.dout(w_dff_B_cjpEUtrF4_2),.clk(gclk));
	jdff dff_B_5WzQe57n6_2(.din(w_dff_B_cjpEUtrF4_2),.dout(w_dff_B_5WzQe57n6_2),.clk(gclk));
	jdff dff_B_sUOIGnBS8_2(.din(w_dff_B_5WzQe57n6_2),.dout(w_dff_B_sUOIGnBS8_2),.clk(gclk));
	jdff dff_B_6texNomC5_2(.din(n364),.dout(w_dff_B_6texNomC5_2),.clk(gclk));
	jdff dff_B_q5ZAGjY43_2(.din(n295),.dout(w_dff_B_q5ZAGjY43_2),.clk(gclk));
	jdff dff_B_ZYfDr3Pu6_2(.din(w_dff_B_q5ZAGjY43_2),.dout(w_dff_B_ZYfDr3Pu6_2),.clk(gclk));
	jdff dff_B_rXwee7iy7_2(.din(w_dff_B_ZYfDr3Pu6_2),.dout(w_dff_B_rXwee7iy7_2),.clk(gclk));
	jdff dff_B_z4cPPlU19_0(.din(n300),.dout(w_dff_B_z4cPPlU19_0),.clk(gclk));
	jdff dff_A_UHb6hdmf2_0(.dout(w_n243_0[0]),.din(w_dff_A_UHb6hdmf2_0),.clk(gclk));
	jdff dff_A_OoN2Prmy8_0(.dout(w_dff_A_UHb6hdmf2_0),.din(w_dff_A_OoN2Prmy8_0),.clk(gclk));
	jdff dff_A_xqfz72US4_1(.dout(w_n243_0[1]),.din(w_dff_A_xqfz72US4_1),.clk(gclk));
	jdff dff_A_U7KNUsVf3_1(.dout(w_dff_A_xqfz72US4_1),.din(w_dff_A_U7KNUsVf3_1),.clk(gclk));
	jdff dff_B_QvWK9LdJ4_1(.din(n1532),.dout(w_dff_B_QvWK9LdJ4_1),.clk(gclk));
	jdff dff_B_ppWMHWH82_2(.din(n1466),.dout(w_dff_B_ppWMHWH82_2),.clk(gclk));
	jdff dff_B_Du9yRvuv4_2(.din(w_dff_B_ppWMHWH82_2),.dout(w_dff_B_Du9yRvuv4_2),.clk(gclk));
	jdff dff_B_rfOzPZWh0_2(.din(w_dff_B_Du9yRvuv4_2),.dout(w_dff_B_rfOzPZWh0_2),.clk(gclk));
	jdff dff_B_YRD4GLRA9_2(.din(w_dff_B_rfOzPZWh0_2),.dout(w_dff_B_YRD4GLRA9_2),.clk(gclk));
	jdff dff_B_qtVBLd7Y9_2(.din(w_dff_B_YRD4GLRA9_2),.dout(w_dff_B_qtVBLd7Y9_2),.clk(gclk));
	jdff dff_B_xXxxeo2k8_2(.din(w_dff_B_qtVBLd7Y9_2),.dout(w_dff_B_xXxxeo2k8_2),.clk(gclk));
	jdff dff_B_d8ZyoDXL4_2(.din(w_dff_B_xXxxeo2k8_2),.dout(w_dff_B_d8ZyoDXL4_2),.clk(gclk));
	jdff dff_B_ZSyl96Lv8_2(.din(w_dff_B_d8ZyoDXL4_2),.dout(w_dff_B_ZSyl96Lv8_2),.clk(gclk));
	jdff dff_B_ty4Ue4Zf2_2(.din(w_dff_B_ZSyl96Lv8_2),.dout(w_dff_B_ty4Ue4Zf2_2),.clk(gclk));
	jdff dff_B_QUKVixNC3_2(.din(w_dff_B_ty4Ue4Zf2_2),.dout(w_dff_B_QUKVixNC3_2),.clk(gclk));
	jdff dff_B_EAF4somy5_2(.din(w_dff_B_QUKVixNC3_2),.dout(w_dff_B_EAF4somy5_2),.clk(gclk));
	jdff dff_B_C9a3ZSxp0_2(.din(w_dff_B_EAF4somy5_2),.dout(w_dff_B_C9a3ZSxp0_2),.clk(gclk));
	jdff dff_B_tNmU4ROw3_2(.din(w_dff_B_C9a3ZSxp0_2),.dout(w_dff_B_tNmU4ROw3_2),.clk(gclk));
	jdff dff_B_8gGogAKO4_2(.din(w_dff_B_tNmU4ROw3_2),.dout(w_dff_B_8gGogAKO4_2),.clk(gclk));
	jdff dff_B_iHw0yWVS2_2(.din(w_dff_B_8gGogAKO4_2),.dout(w_dff_B_iHw0yWVS2_2),.clk(gclk));
	jdff dff_B_BfLDeT4F0_2(.din(w_dff_B_iHw0yWVS2_2),.dout(w_dff_B_BfLDeT4F0_2),.clk(gclk));
	jdff dff_B_HHnTZyAA9_2(.din(w_dff_B_BfLDeT4F0_2),.dout(w_dff_B_HHnTZyAA9_2),.clk(gclk));
	jdff dff_B_6myBpVsI6_2(.din(w_dff_B_HHnTZyAA9_2),.dout(w_dff_B_6myBpVsI6_2),.clk(gclk));
	jdff dff_B_RKm6MBC72_2(.din(w_dff_B_6myBpVsI6_2),.dout(w_dff_B_RKm6MBC72_2),.clk(gclk));
	jdff dff_B_CYVv1W5i4_2(.din(w_dff_B_RKm6MBC72_2),.dout(w_dff_B_CYVv1W5i4_2),.clk(gclk));
	jdff dff_B_l3al1kNK2_2(.din(w_dff_B_CYVv1W5i4_2),.dout(w_dff_B_l3al1kNK2_2),.clk(gclk));
	jdff dff_B_6DiyvSLa4_2(.din(w_dff_B_l3al1kNK2_2),.dout(w_dff_B_6DiyvSLa4_2),.clk(gclk));
	jdff dff_B_coAxeVZi2_2(.din(w_dff_B_6DiyvSLa4_2),.dout(w_dff_B_coAxeVZi2_2),.clk(gclk));
	jdff dff_B_Bm9ZbwX94_2(.din(w_dff_B_coAxeVZi2_2),.dout(w_dff_B_Bm9ZbwX94_2),.clk(gclk));
	jdff dff_B_DSTJ5NN37_2(.din(w_dff_B_Bm9ZbwX94_2),.dout(w_dff_B_DSTJ5NN37_2),.clk(gclk));
	jdff dff_B_bvZFtliG9_2(.din(w_dff_B_DSTJ5NN37_2),.dout(w_dff_B_bvZFtliG9_2),.clk(gclk));
	jdff dff_B_U2I4LaUO3_2(.din(w_dff_B_bvZFtliG9_2),.dout(w_dff_B_U2I4LaUO3_2),.clk(gclk));
	jdff dff_B_3EmoHhCN9_2(.din(w_dff_B_U2I4LaUO3_2),.dout(w_dff_B_3EmoHhCN9_2),.clk(gclk));
	jdff dff_B_vpWzQMEl9_2(.din(w_dff_B_3EmoHhCN9_2),.dout(w_dff_B_vpWzQMEl9_2),.clk(gclk));
	jdff dff_B_RaFgWQMW8_2(.din(w_dff_B_vpWzQMEl9_2),.dout(w_dff_B_RaFgWQMW8_2),.clk(gclk));
	jdff dff_B_85e4b9YS0_2(.din(w_dff_B_RaFgWQMW8_2),.dout(w_dff_B_85e4b9YS0_2),.clk(gclk));
	jdff dff_B_TwqKLTjI6_2(.din(w_dff_B_85e4b9YS0_2),.dout(w_dff_B_TwqKLTjI6_2),.clk(gclk));
	jdff dff_B_IJpz2FlE4_2(.din(w_dff_B_TwqKLTjI6_2),.dout(w_dff_B_IJpz2FlE4_2),.clk(gclk));
	jdff dff_B_RXGS2Cq57_2(.din(w_dff_B_IJpz2FlE4_2),.dout(w_dff_B_RXGS2Cq57_2),.clk(gclk));
	jdff dff_B_NqeVhiCF4_2(.din(w_dff_B_RXGS2Cq57_2),.dout(w_dff_B_NqeVhiCF4_2),.clk(gclk));
	jdff dff_B_KE23DJSF1_2(.din(w_dff_B_NqeVhiCF4_2),.dout(w_dff_B_KE23DJSF1_2),.clk(gclk));
	jdff dff_B_27oEDSQy4_2(.din(w_dff_B_KE23DJSF1_2),.dout(w_dff_B_27oEDSQy4_2),.clk(gclk));
	jdff dff_B_WcwpsT4j7_2(.din(w_dff_B_27oEDSQy4_2),.dout(w_dff_B_WcwpsT4j7_2),.clk(gclk));
	jdff dff_B_OhiqQqoW1_2(.din(w_dff_B_WcwpsT4j7_2),.dout(w_dff_B_OhiqQqoW1_2),.clk(gclk));
	jdff dff_B_e4TzaCi25_2(.din(w_dff_B_OhiqQqoW1_2),.dout(w_dff_B_e4TzaCi25_2),.clk(gclk));
	jdff dff_B_zgaLzjm17_2(.din(w_dff_B_e4TzaCi25_2),.dout(w_dff_B_zgaLzjm17_2),.clk(gclk));
	jdff dff_B_ufmkUT7W0_2(.din(w_dff_B_zgaLzjm17_2),.dout(w_dff_B_ufmkUT7W0_2),.clk(gclk));
	jdff dff_B_OfDykzgp6_2(.din(w_dff_B_ufmkUT7W0_2),.dout(w_dff_B_OfDykzgp6_2),.clk(gclk));
	jdff dff_B_769FflUu8_2(.din(w_dff_B_OfDykzgp6_2),.dout(w_dff_B_769FflUu8_2),.clk(gclk));
	jdff dff_B_cWIKRbme5_2(.din(w_dff_B_769FflUu8_2),.dout(w_dff_B_cWIKRbme5_2),.clk(gclk));
	jdff dff_B_bG14cOkU1_2(.din(w_dff_B_cWIKRbme5_2),.dout(w_dff_B_bG14cOkU1_2),.clk(gclk));
	jdff dff_B_xTRmInr30_0(.din(n1531),.dout(w_dff_B_xTRmInr30_0),.clk(gclk));
	jdff dff_A_Z1NK3AwW0_1(.dout(w_n1519_0[1]),.din(w_dff_A_Z1NK3AwW0_1),.clk(gclk));
	jdff dff_B_JumOCHSu3_1(.din(n1467),.dout(w_dff_B_JumOCHSu3_1),.clk(gclk));
	jdff dff_B_djXDBNZ67_2(.din(n1395),.dout(w_dff_B_djXDBNZ67_2),.clk(gclk));
	jdff dff_B_rgShl3M96_2(.din(w_dff_B_djXDBNZ67_2),.dout(w_dff_B_rgShl3M96_2),.clk(gclk));
	jdff dff_B_MbQSwguy8_2(.din(w_dff_B_rgShl3M96_2),.dout(w_dff_B_MbQSwguy8_2),.clk(gclk));
	jdff dff_B_rTXAzY9u6_2(.din(w_dff_B_MbQSwguy8_2),.dout(w_dff_B_rTXAzY9u6_2),.clk(gclk));
	jdff dff_B_TAxIsREk8_2(.din(w_dff_B_rTXAzY9u6_2),.dout(w_dff_B_TAxIsREk8_2),.clk(gclk));
	jdff dff_B_SWI5FPZO2_2(.din(w_dff_B_TAxIsREk8_2),.dout(w_dff_B_SWI5FPZO2_2),.clk(gclk));
	jdff dff_B_nES1lzeJ1_2(.din(w_dff_B_SWI5FPZO2_2),.dout(w_dff_B_nES1lzeJ1_2),.clk(gclk));
	jdff dff_B_6yVykT7u9_2(.din(w_dff_B_nES1lzeJ1_2),.dout(w_dff_B_6yVykT7u9_2),.clk(gclk));
	jdff dff_B_X9DvH45u2_2(.din(w_dff_B_6yVykT7u9_2),.dout(w_dff_B_X9DvH45u2_2),.clk(gclk));
	jdff dff_B_TOFT54Yp0_2(.din(w_dff_B_X9DvH45u2_2),.dout(w_dff_B_TOFT54Yp0_2),.clk(gclk));
	jdff dff_B_OdCsBtY38_2(.din(w_dff_B_TOFT54Yp0_2),.dout(w_dff_B_OdCsBtY38_2),.clk(gclk));
	jdff dff_B_g10y2h3c7_2(.din(w_dff_B_OdCsBtY38_2),.dout(w_dff_B_g10y2h3c7_2),.clk(gclk));
	jdff dff_B_f3DeNnlr7_2(.din(w_dff_B_g10y2h3c7_2),.dout(w_dff_B_f3DeNnlr7_2),.clk(gclk));
	jdff dff_B_SxCiQWFo4_2(.din(w_dff_B_f3DeNnlr7_2),.dout(w_dff_B_SxCiQWFo4_2),.clk(gclk));
	jdff dff_B_v9SIsnLb9_2(.din(w_dff_B_SxCiQWFo4_2),.dout(w_dff_B_v9SIsnLb9_2),.clk(gclk));
	jdff dff_B_ZNzTCBjo3_2(.din(w_dff_B_v9SIsnLb9_2),.dout(w_dff_B_ZNzTCBjo3_2),.clk(gclk));
	jdff dff_B_egjYoBMq4_2(.din(w_dff_B_ZNzTCBjo3_2),.dout(w_dff_B_egjYoBMq4_2),.clk(gclk));
	jdff dff_B_k4CU2HWw1_2(.din(w_dff_B_egjYoBMq4_2),.dout(w_dff_B_k4CU2HWw1_2),.clk(gclk));
	jdff dff_B_faOXZq9f7_2(.din(w_dff_B_k4CU2HWw1_2),.dout(w_dff_B_faOXZq9f7_2),.clk(gclk));
	jdff dff_B_Ztrfcz5F5_2(.din(w_dff_B_faOXZq9f7_2),.dout(w_dff_B_Ztrfcz5F5_2),.clk(gclk));
	jdff dff_B_an9KytBv9_2(.din(w_dff_B_Ztrfcz5F5_2),.dout(w_dff_B_an9KytBv9_2),.clk(gclk));
	jdff dff_B_LTd2AH0n9_2(.din(w_dff_B_an9KytBv9_2),.dout(w_dff_B_LTd2AH0n9_2),.clk(gclk));
	jdff dff_B_vd0NwYDS0_2(.din(w_dff_B_LTd2AH0n9_2),.dout(w_dff_B_vd0NwYDS0_2),.clk(gclk));
	jdff dff_B_jpAy5BiJ6_2(.din(w_dff_B_vd0NwYDS0_2),.dout(w_dff_B_jpAy5BiJ6_2),.clk(gclk));
	jdff dff_B_Jx3w7Wv96_2(.din(w_dff_B_jpAy5BiJ6_2),.dout(w_dff_B_Jx3w7Wv96_2),.clk(gclk));
	jdff dff_B_mx0KoNRe1_2(.din(w_dff_B_Jx3w7Wv96_2),.dout(w_dff_B_mx0KoNRe1_2),.clk(gclk));
	jdff dff_B_Lrim48jw3_2(.din(w_dff_B_mx0KoNRe1_2),.dout(w_dff_B_Lrim48jw3_2),.clk(gclk));
	jdff dff_B_Gywrwyt91_2(.din(w_dff_B_Lrim48jw3_2),.dout(w_dff_B_Gywrwyt91_2),.clk(gclk));
	jdff dff_B_4stycAfw9_2(.din(w_dff_B_Gywrwyt91_2),.dout(w_dff_B_4stycAfw9_2),.clk(gclk));
	jdff dff_B_5v1tJlmS4_2(.din(w_dff_B_4stycAfw9_2),.dout(w_dff_B_5v1tJlmS4_2),.clk(gclk));
	jdff dff_B_o9DQ50o20_2(.din(w_dff_B_5v1tJlmS4_2),.dout(w_dff_B_o9DQ50o20_2),.clk(gclk));
	jdff dff_B_EMoVDda25_2(.din(w_dff_B_o9DQ50o20_2),.dout(w_dff_B_EMoVDda25_2),.clk(gclk));
	jdff dff_B_480Yo4J14_2(.din(w_dff_B_EMoVDda25_2),.dout(w_dff_B_480Yo4J14_2),.clk(gclk));
	jdff dff_B_KftfVnJe9_2(.din(w_dff_B_480Yo4J14_2),.dout(w_dff_B_KftfVnJe9_2),.clk(gclk));
	jdff dff_B_6Q6U5BxS6_2(.din(w_dff_B_KftfVnJe9_2),.dout(w_dff_B_6Q6U5BxS6_2),.clk(gclk));
	jdff dff_B_lgHEpE4d0_2(.din(w_dff_B_6Q6U5BxS6_2),.dout(w_dff_B_lgHEpE4d0_2),.clk(gclk));
	jdff dff_B_KgXNBHXA8_2(.din(w_dff_B_lgHEpE4d0_2),.dout(w_dff_B_KgXNBHXA8_2),.clk(gclk));
	jdff dff_B_0qqmCVOu2_2(.din(w_dff_B_KgXNBHXA8_2),.dout(w_dff_B_0qqmCVOu2_2),.clk(gclk));
	jdff dff_B_cyDokG0S9_2(.din(w_dff_B_0qqmCVOu2_2),.dout(w_dff_B_cyDokG0S9_2),.clk(gclk));
	jdff dff_B_GRujP2cX2_2(.din(w_dff_B_cyDokG0S9_2),.dout(w_dff_B_GRujP2cX2_2),.clk(gclk));
	jdff dff_B_sDfgSwXx5_2(.din(w_dff_B_GRujP2cX2_2),.dout(w_dff_B_sDfgSwXx5_2),.clk(gclk));
	jdff dff_B_OeZSAjlN6_2(.din(n1448),.dout(w_dff_B_OeZSAjlN6_2),.clk(gclk));
	jdff dff_B_48fLUiLC1_1(.din(n1396),.dout(w_dff_B_48fLUiLC1_1),.clk(gclk));
	jdff dff_B_Ze3kLx3K1_2(.din(n1317),.dout(w_dff_B_Ze3kLx3K1_2),.clk(gclk));
	jdff dff_B_D0RzeeaR9_2(.din(w_dff_B_Ze3kLx3K1_2),.dout(w_dff_B_D0RzeeaR9_2),.clk(gclk));
	jdff dff_B_uvEPI7238_2(.din(w_dff_B_D0RzeeaR9_2),.dout(w_dff_B_uvEPI7238_2),.clk(gclk));
	jdff dff_B_1GtuQFdD7_2(.din(w_dff_B_uvEPI7238_2),.dout(w_dff_B_1GtuQFdD7_2),.clk(gclk));
	jdff dff_B_6I9bN3aj2_2(.din(w_dff_B_1GtuQFdD7_2),.dout(w_dff_B_6I9bN3aj2_2),.clk(gclk));
	jdff dff_B_pDkBuq3W4_2(.din(w_dff_B_6I9bN3aj2_2),.dout(w_dff_B_pDkBuq3W4_2),.clk(gclk));
	jdff dff_B_l6egQqTq1_2(.din(w_dff_B_pDkBuq3W4_2),.dout(w_dff_B_l6egQqTq1_2),.clk(gclk));
	jdff dff_B_EeIx6lWu5_2(.din(w_dff_B_l6egQqTq1_2),.dout(w_dff_B_EeIx6lWu5_2),.clk(gclk));
	jdff dff_B_ZKzze1G45_2(.din(w_dff_B_EeIx6lWu5_2),.dout(w_dff_B_ZKzze1G45_2),.clk(gclk));
	jdff dff_B_5EIQBByw2_2(.din(w_dff_B_ZKzze1G45_2),.dout(w_dff_B_5EIQBByw2_2),.clk(gclk));
	jdff dff_B_WnUd9fAB9_2(.din(w_dff_B_5EIQBByw2_2),.dout(w_dff_B_WnUd9fAB9_2),.clk(gclk));
	jdff dff_B_XJ7ye8VP4_2(.din(w_dff_B_WnUd9fAB9_2),.dout(w_dff_B_XJ7ye8VP4_2),.clk(gclk));
	jdff dff_B_iATijlvg3_2(.din(w_dff_B_XJ7ye8VP4_2),.dout(w_dff_B_iATijlvg3_2),.clk(gclk));
	jdff dff_B_WJsVMLVr2_2(.din(w_dff_B_iATijlvg3_2),.dout(w_dff_B_WJsVMLVr2_2),.clk(gclk));
	jdff dff_B_SoQN8u6O6_2(.din(w_dff_B_WJsVMLVr2_2),.dout(w_dff_B_SoQN8u6O6_2),.clk(gclk));
	jdff dff_B_WMpKEzfw9_2(.din(w_dff_B_SoQN8u6O6_2),.dout(w_dff_B_WMpKEzfw9_2),.clk(gclk));
	jdff dff_B_VyaUp4V64_2(.din(w_dff_B_WMpKEzfw9_2),.dout(w_dff_B_VyaUp4V64_2),.clk(gclk));
	jdff dff_B_eOWDQZM86_2(.din(w_dff_B_VyaUp4V64_2),.dout(w_dff_B_eOWDQZM86_2),.clk(gclk));
	jdff dff_B_9fiXV1DK3_2(.din(w_dff_B_eOWDQZM86_2),.dout(w_dff_B_9fiXV1DK3_2),.clk(gclk));
	jdff dff_B_cVKcOvl73_2(.din(w_dff_B_9fiXV1DK3_2),.dout(w_dff_B_cVKcOvl73_2),.clk(gclk));
	jdff dff_B_2cCtsE6g0_2(.din(w_dff_B_cVKcOvl73_2),.dout(w_dff_B_2cCtsE6g0_2),.clk(gclk));
	jdff dff_B_QFeoGzuf5_2(.din(w_dff_B_2cCtsE6g0_2),.dout(w_dff_B_QFeoGzuf5_2),.clk(gclk));
	jdff dff_B_MpVpW8QW2_2(.din(w_dff_B_QFeoGzuf5_2),.dout(w_dff_B_MpVpW8QW2_2),.clk(gclk));
	jdff dff_B_9I3MpTzM1_2(.din(w_dff_B_MpVpW8QW2_2),.dout(w_dff_B_9I3MpTzM1_2),.clk(gclk));
	jdff dff_B_FsC1pxoD0_2(.din(w_dff_B_9I3MpTzM1_2),.dout(w_dff_B_FsC1pxoD0_2),.clk(gclk));
	jdff dff_B_npHzAUx52_2(.din(w_dff_B_FsC1pxoD0_2),.dout(w_dff_B_npHzAUx52_2),.clk(gclk));
	jdff dff_B_lmkokJKy3_2(.din(w_dff_B_npHzAUx52_2),.dout(w_dff_B_lmkokJKy3_2),.clk(gclk));
	jdff dff_B_Nla71nIv1_2(.din(w_dff_B_lmkokJKy3_2),.dout(w_dff_B_Nla71nIv1_2),.clk(gclk));
	jdff dff_B_rBTTfBLi3_2(.din(w_dff_B_Nla71nIv1_2),.dout(w_dff_B_rBTTfBLi3_2),.clk(gclk));
	jdff dff_B_OsS6zM8y5_2(.din(w_dff_B_rBTTfBLi3_2),.dout(w_dff_B_OsS6zM8y5_2),.clk(gclk));
	jdff dff_B_j7TGoQOg7_2(.din(w_dff_B_OsS6zM8y5_2),.dout(w_dff_B_j7TGoQOg7_2),.clk(gclk));
	jdff dff_B_1xncBhks8_2(.din(w_dff_B_j7TGoQOg7_2),.dout(w_dff_B_1xncBhks8_2),.clk(gclk));
	jdff dff_B_aauT4CO23_2(.din(w_dff_B_1xncBhks8_2),.dout(w_dff_B_aauT4CO23_2),.clk(gclk));
	jdff dff_B_hK8ZzDrd1_2(.din(w_dff_B_aauT4CO23_2),.dout(w_dff_B_hK8ZzDrd1_2),.clk(gclk));
	jdff dff_B_OzuIHOuw2_2(.din(w_dff_B_hK8ZzDrd1_2),.dout(w_dff_B_OzuIHOuw2_2),.clk(gclk));
	jdff dff_B_SyOUUt9X8_2(.din(w_dff_B_OzuIHOuw2_2),.dout(w_dff_B_SyOUUt9X8_2),.clk(gclk));
	jdff dff_B_yX9rmHxl6_2(.din(w_dff_B_SyOUUt9X8_2),.dout(w_dff_B_yX9rmHxl6_2),.clk(gclk));
	jdff dff_B_tUH2K1Kj7_2(.din(w_dff_B_yX9rmHxl6_2),.dout(w_dff_B_tUH2K1Kj7_2),.clk(gclk));
	jdff dff_B_lcTOel7j3_2(.din(n1370),.dout(w_dff_B_lcTOel7j3_2),.clk(gclk));
	jdff dff_B_uDtCWuTI2_1(.din(n1318),.dout(w_dff_B_uDtCWuTI2_1),.clk(gclk));
	jdff dff_B_6Yaw6uqx5_2(.din(n1232),.dout(w_dff_B_6Yaw6uqx5_2),.clk(gclk));
	jdff dff_B_LKpBOd4S8_2(.din(w_dff_B_6Yaw6uqx5_2),.dout(w_dff_B_LKpBOd4S8_2),.clk(gclk));
	jdff dff_B_yJLB6yw02_2(.din(w_dff_B_LKpBOd4S8_2),.dout(w_dff_B_yJLB6yw02_2),.clk(gclk));
	jdff dff_B_GsbWfNwj8_2(.din(w_dff_B_yJLB6yw02_2),.dout(w_dff_B_GsbWfNwj8_2),.clk(gclk));
	jdff dff_B_z9ITqEVW7_2(.din(w_dff_B_GsbWfNwj8_2),.dout(w_dff_B_z9ITqEVW7_2),.clk(gclk));
	jdff dff_B_p9IB5jVJ4_2(.din(w_dff_B_z9ITqEVW7_2),.dout(w_dff_B_p9IB5jVJ4_2),.clk(gclk));
	jdff dff_B_EDkMg6i13_2(.din(w_dff_B_p9IB5jVJ4_2),.dout(w_dff_B_EDkMg6i13_2),.clk(gclk));
	jdff dff_B_lP6sjAII6_2(.din(w_dff_B_EDkMg6i13_2),.dout(w_dff_B_lP6sjAII6_2),.clk(gclk));
	jdff dff_B_8h7NaPld4_2(.din(w_dff_B_lP6sjAII6_2),.dout(w_dff_B_8h7NaPld4_2),.clk(gclk));
	jdff dff_B_J6f9wVXD2_2(.din(w_dff_B_8h7NaPld4_2),.dout(w_dff_B_J6f9wVXD2_2),.clk(gclk));
	jdff dff_B_KD3qxIVs4_2(.din(w_dff_B_J6f9wVXD2_2),.dout(w_dff_B_KD3qxIVs4_2),.clk(gclk));
	jdff dff_B_txNDtw8o4_2(.din(w_dff_B_KD3qxIVs4_2),.dout(w_dff_B_txNDtw8o4_2),.clk(gclk));
	jdff dff_B_GpM0pypo0_2(.din(w_dff_B_txNDtw8o4_2),.dout(w_dff_B_GpM0pypo0_2),.clk(gclk));
	jdff dff_B_iCeFsNNo9_2(.din(w_dff_B_GpM0pypo0_2),.dout(w_dff_B_iCeFsNNo9_2),.clk(gclk));
	jdff dff_B_CUFHkhrZ5_2(.din(w_dff_B_iCeFsNNo9_2),.dout(w_dff_B_CUFHkhrZ5_2),.clk(gclk));
	jdff dff_B_GIlZr1Dv9_2(.din(w_dff_B_CUFHkhrZ5_2),.dout(w_dff_B_GIlZr1Dv9_2),.clk(gclk));
	jdff dff_B_DEd7KeBy8_2(.din(w_dff_B_GIlZr1Dv9_2),.dout(w_dff_B_DEd7KeBy8_2),.clk(gclk));
	jdff dff_B_NrOlrH518_2(.din(w_dff_B_DEd7KeBy8_2),.dout(w_dff_B_NrOlrH518_2),.clk(gclk));
	jdff dff_B_Lth8MXWF7_2(.din(w_dff_B_NrOlrH518_2),.dout(w_dff_B_Lth8MXWF7_2),.clk(gclk));
	jdff dff_B_GH5mXvln3_2(.din(w_dff_B_Lth8MXWF7_2),.dout(w_dff_B_GH5mXvln3_2),.clk(gclk));
	jdff dff_B_nWFoS2jl6_2(.din(w_dff_B_GH5mXvln3_2),.dout(w_dff_B_nWFoS2jl6_2),.clk(gclk));
	jdff dff_B_xiXCikwH9_2(.din(w_dff_B_nWFoS2jl6_2),.dout(w_dff_B_xiXCikwH9_2),.clk(gclk));
	jdff dff_B_jQFxVyoR7_2(.din(w_dff_B_xiXCikwH9_2),.dout(w_dff_B_jQFxVyoR7_2),.clk(gclk));
	jdff dff_B_i0DgvZ6z9_2(.din(w_dff_B_jQFxVyoR7_2),.dout(w_dff_B_i0DgvZ6z9_2),.clk(gclk));
	jdff dff_B_psaKYNCg1_2(.din(w_dff_B_i0DgvZ6z9_2),.dout(w_dff_B_psaKYNCg1_2),.clk(gclk));
	jdff dff_B_zO67d4XR7_2(.din(w_dff_B_psaKYNCg1_2),.dout(w_dff_B_zO67d4XR7_2),.clk(gclk));
	jdff dff_B_PchzTo831_2(.din(w_dff_B_zO67d4XR7_2),.dout(w_dff_B_PchzTo831_2),.clk(gclk));
	jdff dff_B_FhYYglJE0_2(.din(w_dff_B_PchzTo831_2),.dout(w_dff_B_FhYYglJE0_2),.clk(gclk));
	jdff dff_B_0Z8dxuCq2_2(.din(w_dff_B_FhYYglJE0_2),.dout(w_dff_B_0Z8dxuCq2_2),.clk(gclk));
	jdff dff_B_raInsWt43_2(.din(w_dff_B_0Z8dxuCq2_2),.dout(w_dff_B_raInsWt43_2),.clk(gclk));
	jdff dff_B_xjhE7TFx1_2(.din(w_dff_B_raInsWt43_2),.dout(w_dff_B_xjhE7TFx1_2),.clk(gclk));
	jdff dff_B_wtkhyI6N7_2(.din(w_dff_B_xjhE7TFx1_2),.dout(w_dff_B_wtkhyI6N7_2),.clk(gclk));
	jdff dff_B_MB2L94Ng8_2(.din(w_dff_B_wtkhyI6N7_2),.dout(w_dff_B_MB2L94Ng8_2),.clk(gclk));
	jdff dff_B_Jhi8veVz7_2(.din(w_dff_B_MB2L94Ng8_2),.dout(w_dff_B_Jhi8veVz7_2),.clk(gclk));
	jdff dff_B_1dOlMKis6_2(.din(w_dff_B_Jhi8veVz7_2),.dout(w_dff_B_1dOlMKis6_2),.clk(gclk));
	jdff dff_B_Jne99qpP9_2(.din(n1285),.dout(w_dff_B_Jne99qpP9_2),.clk(gclk));
	jdff dff_B_wqdKiwbS9_1(.din(n1233),.dout(w_dff_B_wqdKiwbS9_1),.clk(gclk));
	jdff dff_B_CHpjLhuk3_2(.din(n1141),.dout(w_dff_B_CHpjLhuk3_2),.clk(gclk));
	jdff dff_B_LpyoHiG38_2(.din(w_dff_B_CHpjLhuk3_2),.dout(w_dff_B_LpyoHiG38_2),.clk(gclk));
	jdff dff_B_oT9evhYB1_2(.din(w_dff_B_LpyoHiG38_2),.dout(w_dff_B_oT9evhYB1_2),.clk(gclk));
	jdff dff_B_YfPu9CoH1_2(.din(w_dff_B_oT9evhYB1_2),.dout(w_dff_B_YfPu9CoH1_2),.clk(gclk));
	jdff dff_B_58QxJlSM5_2(.din(w_dff_B_YfPu9CoH1_2),.dout(w_dff_B_58QxJlSM5_2),.clk(gclk));
	jdff dff_B_zteXz2tj4_2(.din(w_dff_B_58QxJlSM5_2),.dout(w_dff_B_zteXz2tj4_2),.clk(gclk));
	jdff dff_B_tzSbd6xs9_2(.din(w_dff_B_zteXz2tj4_2),.dout(w_dff_B_tzSbd6xs9_2),.clk(gclk));
	jdff dff_B_QoKpxNwm7_2(.din(w_dff_B_tzSbd6xs9_2),.dout(w_dff_B_QoKpxNwm7_2),.clk(gclk));
	jdff dff_B_1HGe7cXS1_2(.din(w_dff_B_QoKpxNwm7_2),.dout(w_dff_B_1HGe7cXS1_2),.clk(gclk));
	jdff dff_B_btzooBeW8_2(.din(w_dff_B_1HGe7cXS1_2),.dout(w_dff_B_btzooBeW8_2),.clk(gclk));
	jdff dff_B_pWBrxOSL1_2(.din(w_dff_B_btzooBeW8_2),.dout(w_dff_B_pWBrxOSL1_2),.clk(gclk));
	jdff dff_B_DPu6pGJB2_2(.din(w_dff_B_pWBrxOSL1_2),.dout(w_dff_B_DPu6pGJB2_2),.clk(gclk));
	jdff dff_B_AzLLaukc4_2(.din(w_dff_B_DPu6pGJB2_2),.dout(w_dff_B_AzLLaukc4_2),.clk(gclk));
	jdff dff_B_9VsHYNVU5_2(.din(w_dff_B_AzLLaukc4_2),.dout(w_dff_B_9VsHYNVU5_2),.clk(gclk));
	jdff dff_B_R2wqIfy29_2(.din(w_dff_B_9VsHYNVU5_2),.dout(w_dff_B_R2wqIfy29_2),.clk(gclk));
	jdff dff_B_61Mi9vDS6_2(.din(w_dff_B_R2wqIfy29_2),.dout(w_dff_B_61Mi9vDS6_2),.clk(gclk));
	jdff dff_B_m9xDWTid6_2(.din(w_dff_B_61Mi9vDS6_2),.dout(w_dff_B_m9xDWTid6_2),.clk(gclk));
	jdff dff_B_CcgNIaTM2_2(.din(w_dff_B_m9xDWTid6_2),.dout(w_dff_B_CcgNIaTM2_2),.clk(gclk));
	jdff dff_B_h5OAkxsp3_2(.din(w_dff_B_CcgNIaTM2_2),.dout(w_dff_B_h5OAkxsp3_2),.clk(gclk));
	jdff dff_B_HEGYzhwY5_2(.din(w_dff_B_h5OAkxsp3_2),.dout(w_dff_B_HEGYzhwY5_2),.clk(gclk));
	jdff dff_B_kfbk9PY04_2(.din(w_dff_B_HEGYzhwY5_2),.dout(w_dff_B_kfbk9PY04_2),.clk(gclk));
	jdff dff_B_jmaO7NWx0_2(.din(w_dff_B_kfbk9PY04_2),.dout(w_dff_B_jmaO7NWx0_2),.clk(gclk));
	jdff dff_B_TShXzsna3_2(.din(w_dff_B_jmaO7NWx0_2),.dout(w_dff_B_TShXzsna3_2),.clk(gclk));
	jdff dff_B_pNS8rVN69_2(.din(w_dff_B_TShXzsna3_2),.dout(w_dff_B_pNS8rVN69_2),.clk(gclk));
	jdff dff_B_hFPCJFyh2_2(.din(w_dff_B_pNS8rVN69_2),.dout(w_dff_B_hFPCJFyh2_2),.clk(gclk));
	jdff dff_B_A0tafV0w9_2(.din(w_dff_B_hFPCJFyh2_2),.dout(w_dff_B_A0tafV0w9_2),.clk(gclk));
	jdff dff_B_AEbfou5c6_2(.din(w_dff_B_A0tafV0w9_2),.dout(w_dff_B_AEbfou5c6_2),.clk(gclk));
	jdff dff_B_K75tx89b6_2(.din(w_dff_B_AEbfou5c6_2),.dout(w_dff_B_K75tx89b6_2),.clk(gclk));
	jdff dff_B_wzPUwsfF3_2(.din(w_dff_B_K75tx89b6_2),.dout(w_dff_B_wzPUwsfF3_2),.clk(gclk));
	jdff dff_B_ZZcJZLBn4_2(.din(w_dff_B_wzPUwsfF3_2),.dout(w_dff_B_ZZcJZLBn4_2),.clk(gclk));
	jdff dff_B_4VF6pijT7_2(.din(w_dff_B_ZZcJZLBn4_2),.dout(w_dff_B_4VF6pijT7_2),.clk(gclk));
	jdff dff_B_4HCmCGDr6_2(.din(w_dff_B_4VF6pijT7_2),.dout(w_dff_B_4HCmCGDr6_2),.clk(gclk));
	jdff dff_B_xjUxkvVQ5_2(.din(n1194),.dout(w_dff_B_xjUxkvVQ5_2),.clk(gclk));
	jdff dff_B_Ks3Cgzof9_1(.din(n1142),.dout(w_dff_B_Ks3Cgzof9_1),.clk(gclk));
	jdff dff_B_LotTPgHT2_2(.din(n1043),.dout(w_dff_B_LotTPgHT2_2),.clk(gclk));
	jdff dff_B_eiVwXRlF0_2(.din(w_dff_B_LotTPgHT2_2),.dout(w_dff_B_eiVwXRlF0_2),.clk(gclk));
	jdff dff_B_GApNkSkT3_2(.din(w_dff_B_eiVwXRlF0_2),.dout(w_dff_B_GApNkSkT3_2),.clk(gclk));
	jdff dff_B_0UPiT9ic9_2(.din(w_dff_B_GApNkSkT3_2),.dout(w_dff_B_0UPiT9ic9_2),.clk(gclk));
	jdff dff_B_Il2GKSpk7_2(.din(w_dff_B_0UPiT9ic9_2),.dout(w_dff_B_Il2GKSpk7_2),.clk(gclk));
	jdff dff_B_lUTGmdDb2_2(.din(w_dff_B_Il2GKSpk7_2),.dout(w_dff_B_lUTGmdDb2_2),.clk(gclk));
	jdff dff_B_xuW5NKz55_2(.din(w_dff_B_lUTGmdDb2_2),.dout(w_dff_B_xuW5NKz55_2),.clk(gclk));
	jdff dff_B_w1R3Xp8i3_2(.din(w_dff_B_xuW5NKz55_2),.dout(w_dff_B_w1R3Xp8i3_2),.clk(gclk));
	jdff dff_B_DQw6JW6I5_2(.din(w_dff_B_w1R3Xp8i3_2),.dout(w_dff_B_DQw6JW6I5_2),.clk(gclk));
	jdff dff_B_ThdgcyjF7_2(.din(w_dff_B_DQw6JW6I5_2),.dout(w_dff_B_ThdgcyjF7_2),.clk(gclk));
	jdff dff_B_Fm0jZ2AS0_2(.din(w_dff_B_ThdgcyjF7_2),.dout(w_dff_B_Fm0jZ2AS0_2),.clk(gclk));
	jdff dff_B_9hfurshI2_2(.din(w_dff_B_Fm0jZ2AS0_2),.dout(w_dff_B_9hfurshI2_2),.clk(gclk));
	jdff dff_B_fFRCeOFU6_2(.din(w_dff_B_9hfurshI2_2),.dout(w_dff_B_fFRCeOFU6_2),.clk(gclk));
	jdff dff_B_sL9yCUtx2_2(.din(w_dff_B_fFRCeOFU6_2),.dout(w_dff_B_sL9yCUtx2_2),.clk(gclk));
	jdff dff_B_zBNIm5ku7_2(.din(w_dff_B_sL9yCUtx2_2),.dout(w_dff_B_zBNIm5ku7_2),.clk(gclk));
	jdff dff_B_35zlfNO25_2(.din(w_dff_B_zBNIm5ku7_2),.dout(w_dff_B_35zlfNO25_2),.clk(gclk));
	jdff dff_B_ozIz7hsk9_2(.din(w_dff_B_35zlfNO25_2),.dout(w_dff_B_ozIz7hsk9_2),.clk(gclk));
	jdff dff_B_iBDx4kTa8_2(.din(w_dff_B_ozIz7hsk9_2),.dout(w_dff_B_iBDx4kTa8_2),.clk(gclk));
	jdff dff_B_FRqwOUtL0_2(.din(w_dff_B_iBDx4kTa8_2),.dout(w_dff_B_FRqwOUtL0_2),.clk(gclk));
	jdff dff_B_5SioB8bi0_2(.din(w_dff_B_FRqwOUtL0_2),.dout(w_dff_B_5SioB8bi0_2),.clk(gclk));
	jdff dff_B_dRfhkIXO6_2(.din(w_dff_B_5SioB8bi0_2),.dout(w_dff_B_dRfhkIXO6_2),.clk(gclk));
	jdff dff_B_meGfJ4Ml7_2(.din(w_dff_B_dRfhkIXO6_2),.dout(w_dff_B_meGfJ4Ml7_2),.clk(gclk));
	jdff dff_B_THRXSfUE3_2(.din(w_dff_B_meGfJ4Ml7_2),.dout(w_dff_B_THRXSfUE3_2),.clk(gclk));
	jdff dff_B_djv53PIm9_2(.din(w_dff_B_THRXSfUE3_2),.dout(w_dff_B_djv53PIm9_2),.clk(gclk));
	jdff dff_B_EQBEhJzu3_2(.din(w_dff_B_djv53PIm9_2),.dout(w_dff_B_EQBEhJzu3_2),.clk(gclk));
	jdff dff_B_SbD6dXDL5_2(.din(w_dff_B_EQBEhJzu3_2),.dout(w_dff_B_SbD6dXDL5_2),.clk(gclk));
	jdff dff_B_PZcz0VKj4_2(.din(w_dff_B_SbD6dXDL5_2),.dout(w_dff_B_PZcz0VKj4_2),.clk(gclk));
	jdff dff_B_Vv5vw15y6_2(.din(w_dff_B_PZcz0VKj4_2),.dout(w_dff_B_Vv5vw15y6_2),.clk(gclk));
	jdff dff_B_wqQfrI6j6_2(.din(w_dff_B_Vv5vw15y6_2),.dout(w_dff_B_wqQfrI6j6_2),.clk(gclk));
	jdff dff_B_xho3upNn0_2(.din(n1095),.dout(w_dff_B_xho3upNn0_2),.clk(gclk));
	jdff dff_B_fiFeTNe63_1(.din(n1044),.dout(w_dff_B_fiFeTNe63_1),.clk(gclk));
	jdff dff_B_9HwILk8E8_2(.din(n944),.dout(w_dff_B_9HwILk8E8_2),.clk(gclk));
	jdff dff_B_BmLP96EL6_2(.din(w_dff_B_9HwILk8E8_2),.dout(w_dff_B_BmLP96EL6_2),.clk(gclk));
	jdff dff_B_95OsEaqm3_2(.din(w_dff_B_BmLP96EL6_2),.dout(w_dff_B_95OsEaqm3_2),.clk(gclk));
	jdff dff_B_u1vD9SdR2_2(.din(w_dff_B_95OsEaqm3_2),.dout(w_dff_B_u1vD9SdR2_2),.clk(gclk));
	jdff dff_B_iyhTj8nm2_2(.din(w_dff_B_u1vD9SdR2_2),.dout(w_dff_B_iyhTj8nm2_2),.clk(gclk));
	jdff dff_B_M4IeJZNd0_2(.din(w_dff_B_iyhTj8nm2_2),.dout(w_dff_B_M4IeJZNd0_2),.clk(gclk));
	jdff dff_B_ZEyAsnHN7_2(.din(w_dff_B_M4IeJZNd0_2),.dout(w_dff_B_ZEyAsnHN7_2),.clk(gclk));
	jdff dff_B_4WlfT4Mr9_2(.din(w_dff_B_ZEyAsnHN7_2),.dout(w_dff_B_4WlfT4Mr9_2),.clk(gclk));
	jdff dff_B_tbs6DpMD0_2(.din(w_dff_B_4WlfT4Mr9_2),.dout(w_dff_B_tbs6DpMD0_2),.clk(gclk));
	jdff dff_B_L8MrorfR3_2(.din(w_dff_B_tbs6DpMD0_2),.dout(w_dff_B_L8MrorfR3_2),.clk(gclk));
	jdff dff_B_u8g5p00Q1_2(.din(w_dff_B_L8MrorfR3_2),.dout(w_dff_B_u8g5p00Q1_2),.clk(gclk));
	jdff dff_B_5dMGJnKw8_2(.din(w_dff_B_u8g5p00Q1_2),.dout(w_dff_B_5dMGJnKw8_2),.clk(gclk));
	jdff dff_B_auTy16xV2_2(.din(w_dff_B_5dMGJnKw8_2),.dout(w_dff_B_auTy16xV2_2),.clk(gclk));
	jdff dff_B_jzl2WbeF3_2(.din(w_dff_B_auTy16xV2_2),.dout(w_dff_B_jzl2WbeF3_2),.clk(gclk));
	jdff dff_B_VAok8B1c7_2(.din(w_dff_B_jzl2WbeF3_2),.dout(w_dff_B_VAok8B1c7_2),.clk(gclk));
	jdff dff_B_UYzEA5X27_2(.din(w_dff_B_VAok8B1c7_2),.dout(w_dff_B_UYzEA5X27_2),.clk(gclk));
	jdff dff_B_d2Gkv2e39_2(.din(w_dff_B_UYzEA5X27_2),.dout(w_dff_B_d2Gkv2e39_2),.clk(gclk));
	jdff dff_B_0eXg0p0U9_2(.din(w_dff_B_d2Gkv2e39_2),.dout(w_dff_B_0eXg0p0U9_2),.clk(gclk));
	jdff dff_B_xiRj92M16_2(.din(w_dff_B_0eXg0p0U9_2),.dout(w_dff_B_xiRj92M16_2),.clk(gclk));
	jdff dff_B_u6oZYj6j5_2(.din(w_dff_B_xiRj92M16_2),.dout(w_dff_B_u6oZYj6j5_2),.clk(gclk));
	jdff dff_B_TnozkIyp2_2(.din(w_dff_B_u6oZYj6j5_2),.dout(w_dff_B_TnozkIyp2_2),.clk(gclk));
	jdff dff_B_qnhEsylH2_2(.din(w_dff_B_TnozkIyp2_2),.dout(w_dff_B_qnhEsylH2_2),.clk(gclk));
	jdff dff_B_qkhO7al72_2(.din(w_dff_B_qnhEsylH2_2),.dout(w_dff_B_qkhO7al72_2),.clk(gclk));
	jdff dff_B_y6kwC2sf6_2(.din(w_dff_B_qkhO7al72_2),.dout(w_dff_B_y6kwC2sf6_2),.clk(gclk));
	jdff dff_B_vV0bDt1L1_2(.din(w_dff_B_y6kwC2sf6_2),.dout(w_dff_B_vV0bDt1L1_2),.clk(gclk));
	jdff dff_B_lZ5Qjorr3_2(.din(w_dff_B_vV0bDt1L1_2),.dout(w_dff_B_lZ5Qjorr3_2),.clk(gclk));
	jdff dff_B_bcP0E7Hi5_2(.din(n996),.dout(w_dff_B_bcP0E7Hi5_2),.clk(gclk));
	jdff dff_B_PDENw4BN8_1(.din(n945),.dout(w_dff_B_PDENw4BN8_1),.clk(gclk));
	jdff dff_B_hNgHePwe0_2(.din(n842),.dout(w_dff_B_hNgHePwe0_2),.clk(gclk));
	jdff dff_B_LygJ5N0O7_2(.din(w_dff_B_hNgHePwe0_2),.dout(w_dff_B_LygJ5N0O7_2),.clk(gclk));
	jdff dff_B_vLA6d5pQ6_2(.din(w_dff_B_LygJ5N0O7_2),.dout(w_dff_B_vLA6d5pQ6_2),.clk(gclk));
	jdff dff_B_Cgfh33L38_2(.din(w_dff_B_vLA6d5pQ6_2),.dout(w_dff_B_Cgfh33L38_2),.clk(gclk));
	jdff dff_B_SlTnutle6_2(.din(w_dff_B_Cgfh33L38_2),.dout(w_dff_B_SlTnutle6_2),.clk(gclk));
	jdff dff_B_piViiJcf3_2(.din(w_dff_B_SlTnutle6_2),.dout(w_dff_B_piViiJcf3_2),.clk(gclk));
	jdff dff_B_o90DMMD02_2(.din(w_dff_B_piViiJcf3_2),.dout(w_dff_B_o90DMMD02_2),.clk(gclk));
	jdff dff_B_4XRK2MfO1_2(.din(w_dff_B_o90DMMD02_2),.dout(w_dff_B_4XRK2MfO1_2),.clk(gclk));
	jdff dff_B_Umx2e0Ti1_2(.din(w_dff_B_4XRK2MfO1_2),.dout(w_dff_B_Umx2e0Ti1_2),.clk(gclk));
	jdff dff_B_V9ZXbxxY2_2(.din(w_dff_B_Umx2e0Ti1_2),.dout(w_dff_B_V9ZXbxxY2_2),.clk(gclk));
	jdff dff_B_ptmoT6kf6_2(.din(w_dff_B_V9ZXbxxY2_2),.dout(w_dff_B_ptmoT6kf6_2),.clk(gclk));
	jdff dff_B_uyGMp8xf6_2(.din(w_dff_B_ptmoT6kf6_2),.dout(w_dff_B_uyGMp8xf6_2),.clk(gclk));
	jdff dff_B_0aqzSceQ4_2(.din(w_dff_B_uyGMp8xf6_2),.dout(w_dff_B_0aqzSceQ4_2),.clk(gclk));
	jdff dff_B_WfaHkpyi8_2(.din(w_dff_B_0aqzSceQ4_2),.dout(w_dff_B_WfaHkpyi8_2),.clk(gclk));
	jdff dff_B_FQgo4IeQ5_2(.din(w_dff_B_WfaHkpyi8_2),.dout(w_dff_B_FQgo4IeQ5_2),.clk(gclk));
	jdff dff_B_aHhwdnR76_2(.din(w_dff_B_FQgo4IeQ5_2),.dout(w_dff_B_aHhwdnR76_2),.clk(gclk));
	jdff dff_B_EZTUX7EG6_2(.din(w_dff_B_aHhwdnR76_2),.dout(w_dff_B_EZTUX7EG6_2),.clk(gclk));
	jdff dff_B_11je3hXV5_2(.din(w_dff_B_EZTUX7EG6_2),.dout(w_dff_B_11je3hXV5_2),.clk(gclk));
	jdff dff_B_dNzfvh2j6_2(.din(w_dff_B_11je3hXV5_2),.dout(w_dff_B_dNzfvh2j6_2),.clk(gclk));
	jdff dff_B_ii4FWdKs3_2(.din(w_dff_B_dNzfvh2j6_2),.dout(w_dff_B_ii4FWdKs3_2),.clk(gclk));
	jdff dff_B_PMTWwnZD2_2(.din(w_dff_B_ii4FWdKs3_2),.dout(w_dff_B_PMTWwnZD2_2),.clk(gclk));
	jdff dff_B_2R7uQTqB7_2(.din(w_dff_B_PMTWwnZD2_2),.dout(w_dff_B_2R7uQTqB7_2),.clk(gclk));
	jdff dff_B_Jyz2QApv5_2(.din(w_dff_B_2R7uQTqB7_2),.dout(w_dff_B_Jyz2QApv5_2),.clk(gclk));
	jdff dff_B_JBIaOyn81_2(.din(n890),.dout(w_dff_B_JBIaOyn81_2),.clk(gclk));
	jdff dff_B_yT5jobxk4_1(.din(n843),.dout(w_dff_B_yT5jobxk4_1),.clk(gclk));
	jdff dff_B_7JAqNfso5_2(.din(n744),.dout(w_dff_B_7JAqNfso5_2),.clk(gclk));
	jdff dff_B_retg5sal1_2(.din(w_dff_B_7JAqNfso5_2),.dout(w_dff_B_retg5sal1_2),.clk(gclk));
	jdff dff_B_A4vrtnSH3_2(.din(w_dff_B_retg5sal1_2),.dout(w_dff_B_A4vrtnSH3_2),.clk(gclk));
	jdff dff_B_qlYry9lt8_2(.din(w_dff_B_A4vrtnSH3_2),.dout(w_dff_B_qlYry9lt8_2),.clk(gclk));
	jdff dff_B_r1y2DTad6_2(.din(w_dff_B_qlYry9lt8_2),.dout(w_dff_B_r1y2DTad6_2),.clk(gclk));
	jdff dff_B_IpJS6Yjr3_2(.din(w_dff_B_r1y2DTad6_2),.dout(w_dff_B_IpJS6Yjr3_2),.clk(gclk));
	jdff dff_B_aSytTE3v5_2(.din(w_dff_B_IpJS6Yjr3_2),.dout(w_dff_B_aSytTE3v5_2),.clk(gclk));
	jdff dff_B_eA3eVsOS5_2(.din(w_dff_B_aSytTE3v5_2),.dout(w_dff_B_eA3eVsOS5_2),.clk(gclk));
	jdff dff_B_NmyyoUbH7_2(.din(w_dff_B_eA3eVsOS5_2),.dout(w_dff_B_NmyyoUbH7_2),.clk(gclk));
	jdff dff_B_N30qgxtY5_2(.din(w_dff_B_NmyyoUbH7_2),.dout(w_dff_B_N30qgxtY5_2),.clk(gclk));
	jdff dff_B_sBD5fOAS7_2(.din(w_dff_B_N30qgxtY5_2),.dout(w_dff_B_sBD5fOAS7_2),.clk(gclk));
	jdff dff_B_ROiWYELl3_2(.din(w_dff_B_sBD5fOAS7_2),.dout(w_dff_B_ROiWYELl3_2),.clk(gclk));
	jdff dff_B_JwGCPUiN1_2(.din(w_dff_B_ROiWYELl3_2),.dout(w_dff_B_JwGCPUiN1_2),.clk(gclk));
	jdff dff_B_QP6oDmvm3_2(.din(w_dff_B_JwGCPUiN1_2),.dout(w_dff_B_QP6oDmvm3_2),.clk(gclk));
	jdff dff_B_IrJyoUG20_2(.din(w_dff_B_QP6oDmvm3_2),.dout(w_dff_B_IrJyoUG20_2),.clk(gclk));
	jdff dff_B_Vh5xl8JH8_2(.din(w_dff_B_IrJyoUG20_2),.dout(w_dff_B_Vh5xl8JH8_2),.clk(gclk));
	jdff dff_B_uhyn0yt57_2(.din(w_dff_B_Vh5xl8JH8_2),.dout(w_dff_B_uhyn0yt57_2),.clk(gclk));
	jdff dff_B_8vJAl03n1_2(.din(w_dff_B_uhyn0yt57_2),.dout(w_dff_B_8vJAl03n1_2),.clk(gclk));
	jdff dff_B_3r6Rjrm44_2(.din(w_dff_B_8vJAl03n1_2),.dout(w_dff_B_3r6Rjrm44_2),.clk(gclk));
	jdff dff_B_QJ1fA5oe5_2(.din(w_dff_B_3r6Rjrm44_2),.dout(w_dff_B_QJ1fA5oe5_2),.clk(gclk));
	jdff dff_B_OBfPOlGw5_2(.din(n787),.dout(w_dff_B_OBfPOlGw5_2),.clk(gclk));
	jdff dff_B_Y00TVUep1_1(.din(n745),.dout(w_dff_B_Y00TVUep1_1),.clk(gclk));
	jdff dff_B_GBVQ5kQi4_2(.din(n652),.dout(w_dff_B_GBVQ5kQi4_2),.clk(gclk));
	jdff dff_B_emarn5hR8_2(.din(w_dff_B_GBVQ5kQi4_2),.dout(w_dff_B_emarn5hR8_2),.clk(gclk));
	jdff dff_B_xo7lOydL0_2(.din(w_dff_B_emarn5hR8_2),.dout(w_dff_B_xo7lOydL0_2),.clk(gclk));
	jdff dff_B_1y3bl1DT5_2(.din(w_dff_B_xo7lOydL0_2),.dout(w_dff_B_1y3bl1DT5_2),.clk(gclk));
	jdff dff_B_S8pJRnZ08_2(.din(w_dff_B_1y3bl1DT5_2),.dout(w_dff_B_S8pJRnZ08_2),.clk(gclk));
	jdff dff_B_zyBgXcK69_2(.din(w_dff_B_S8pJRnZ08_2),.dout(w_dff_B_zyBgXcK69_2),.clk(gclk));
	jdff dff_B_2l6JgLO20_2(.din(w_dff_B_zyBgXcK69_2),.dout(w_dff_B_2l6JgLO20_2),.clk(gclk));
	jdff dff_B_vvGstb3u6_2(.din(w_dff_B_2l6JgLO20_2),.dout(w_dff_B_vvGstb3u6_2),.clk(gclk));
	jdff dff_B_Ojxe2w5V1_2(.din(w_dff_B_vvGstb3u6_2),.dout(w_dff_B_Ojxe2w5V1_2),.clk(gclk));
	jdff dff_B_NJQC5RLN1_2(.din(w_dff_B_Ojxe2w5V1_2),.dout(w_dff_B_NJQC5RLN1_2),.clk(gclk));
	jdff dff_B_xkyLc5QC5_2(.din(w_dff_B_NJQC5RLN1_2),.dout(w_dff_B_xkyLc5QC5_2),.clk(gclk));
	jdff dff_B_g4Xk05fy1_2(.din(w_dff_B_xkyLc5QC5_2),.dout(w_dff_B_g4Xk05fy1_2),.clk(gclk));
	jdff dff_B_LojWqOlZ3_2(.din(w_dff_B_g4Xk05fy1_2),.dout(w_dff_B_LojWqOlZ3_2),.clk(gclk));
	jdff dff_B_B9DS5n4x2_2(.din(w_dff_B_LojWqOlZ3_2),.dout(w_dff_B_B9DS5n4x2_2),.clk(gclk));
	jdff dff_B_UzAZefYP7_2(.din(w_dff_B_B9DS5n4x2_2),.dout(w_dff_B_UzAZefYP7_2),.clk(gclk));
	jdff dff_B_zRtuluKM3_2(.din(w_dff_B_UzAZefYP7_2),.dout(w_dff_B_zRtuluKM3_2),.clk(gclk));
	jdff dff_B_uqRp0sXY8_2(.din(w_dff_B_zRtuluKM3_2),.dout(w_dff_B_uqRp0sXY8_2),.clk(gclk));
	jdff dff_B_dnBmfhxP0_2(.din(n688),.dout(w_dff_B_dnBmfhxP0_2),.clk(gclk));
	jdff dff_B_3HGlLHHK0_1(.din(n653),.dout(w_dff_B_3HGlLHHK0_1),.clk(gclk));
	jdff dff_B_YfSYz0J25_2(.din(n567),.dout(w_dff_B_YfSYz0J25_2),.clk(gclk));
	jdff dff_B_zRZmOvmZ9_2(.din(w_dff_B_YfSYz0J25_2),.dout(w_dff_B_zRZmOvmZ9_2),.clk(gclk));
	jdff dff_B_vHLmVdCp7_2(.din(w_dff_B_zRZmOvmZ9_2),.dout(w_dff_B_vHLmVdCp7_2),.clk(gclk));
	jdff dff_B_WeDC8Aqf4_2(.din(w_dff_B_vHLmVdCp7_2),.dout(w_dff_B_WeDC8Aqf4_2),.clk(gclk));
	jdff dff_B_pCDmsHui1_2(.din(w_dff_B_WeDC8Aqf4_2),.dout(w_dff_B_pCDmsHui1_2),.clk(gclk));
	jdff dff_B_A5EVWbOE0_2(.din(w_dff_B_pCDmsHui1_2),.dout(w_dff_B_A5EVWbOE0_2),.clk(gclk));
	jdff dff_B_ygM08s7E1_2(.din(w_dff_B_A5EVWbOE0_2),.dout(w_dff_B_ygM08s7E1_2),.clk(gclk));
	jdff dff_B_IIZZ6ubz3_2(.din(w_dff_B_ygM08s7E1_2),.dout(w_dff_B_IIZZ6ubz3_2),.clk(gclk));
	jdff dff_B_rCEn5z0B8_2(.din(w_dff_B_IIZZ6ubz3_2),.dout(w_dff_B_rCEn5z0B8_2),.clk(gclk));
	jdff dff_B_Xo7uSpIc3_2(.din(w_dff_B_rCEn5z0B8_2),.dout(w_dff_B_Xo7uSpIc3_2),.clk(gclk));
	jdff dff_B_AUIvz5kU7_2(.din(w_dff_B_Xo7uSpIc3_2),.dout(w_dff_B_AUIvz5kU7_2),.clk(gclk));
	jdff dff_B_6J6Zapwv8_2(.din(w_dff_B_AUIvz5kU7_2),.dout(w_dff_B_6J6Zapwv8_2),.clk(gclk));
	jdff dff_B_Qds8q9tS3_2(.din(w_dff_B_6J6Zapwv8_2),.dout(w_dff_B_Qds8q9tS3_2),.clk(gclk));
	jdff dff_B_3uAKOUMy2_2(.din(w_dff_B_Qds8q9tS3_2),.dout(w_dff_B_3uAKOUMy2_2),.clk(gclk));
	jdff dff_B_aW03qvsr3_2(.din(n596),.dout(w_dff_B_aW03qvsr3_2),.clk(gclk));
	jdff dff_B_5W1HNHhA0_1(.din(n568),.dout(w_dff_B_5W1HNHhA0_1),.clk(gclk));
	jdff dff_B_zeqJF3l42_2(.din(n489),.dout(w_dff_B_zeqJF3l42_2),.clk(gclk));
	jdff dff_B_EX0KBTux0_2(.din(w_dff_B_zeqJF3l42_2),.dout(w_dff_B_EX0KBTux0_2),.clk(gclk));
	jdff dff_B_40DQ05gC1_2(.din(w_dff_B_EX0KBTux0_2),.dout(w_dff_B_40DQ05gC1_2),.clk(gclk));
	jdff dff_B_ispNmflQ4_2(.din(w_dff_B_40DQ05gC1_2),.dout(w_dff_B_ispNmflQ4_2),.clk(gclk));
	jdff dff_B_SUYk7Gpm9_2(.din(w_dff_B_ispNmflQ4_2),.dout(w_dff_B_SUYk7Gpm9_2),.clk(gclk));
	jdff dff_B_0wiadfvI9_2(.din(w_dff_B_SUYk7Gpm9_2),.dout(w_dff_B_0wiadfvI9_2),.clk(gclk));
	jdff dff_B_wCwrZ7sT0_2(.din(w_dff_B_0wiadfvI9_2),.dout(w_dff_B_wCwrZ7sT0_2),.clk(gclk));
	jdff dff_B_Ez6ZSNkI5_2(.din(w_dff_B_wCwrZ7sT0_2),.dout(w_dff_B_Ez6ZSNkI5_2),.clk(gclk));
	jdff dff_B_9qG03qPU5_2(.din(w_dff_B_Ez6ZSNkI5_2),.dout(w_dff_B_9qG03qPU5_2),.clk(gclk));
	jdff dff_B_lFuhzVqH5_2(.din(w_dff_B_9qG03qPU5_2),.dout(w_dff_B_lFuhzVqH5_2),.clk(gclk));
	jdff dff_B_YFOUAA3M5_2(.din(w_dff_B_lFuhzVqH5_2),.dout(w_dff_B_YFOUAA3M5_2),.clk(gclk));
	jdff dff_B_H0YJAthz5_2(.din(n511),.dout(w_dff_B_H0YJAthz5_2),.clk(gclk));
	jdff dff_B_TG7ggu479_1(.din(n490),.dout(w_dff_B_TG7ggu479_1),.clk(gclk));
	jdff dff_B_gICaoszp8_2(.din(n418),.dout(w_dff_B_gICaoszp8_2),.clk(gclk));
	jdff dff_B_AQ3BNbBd1_2(.din(w_dff_B_gICaoszp8_2),.dout(w_dff_B_AQ3BNbBd1_2),.clk(gclk));
	jdff dff_B_LpODIpdX2_2(.din(w_dff_B_AQ3BNbBd1_2),.dout(w_dff_B_LpODIpdX2_2),.clk(gclk));
	jdff dff_B_qCK0mbns7_2(.din(w_dff_B_LpODIpdX2_2),.dout(w_dff_B_qCK0mbns7_2),.clk(gclk));
	jdff dff_B_yM5iZlxK9_2(.din(w_dff_B_qCK0mbns7_2),.dout(w_dff_B_yM5iZlxK9_2),.clk(gclk));
	jdff dff_B_dE0RJCMY2_2(.din(w_dff_B_yM5iZlxK9_2),.dout(w_dff_B_dE0RJCMY2_2),.clk(gclk));
	jdff dff_B_BnSvBPJn0_2(.din(w_dff_B_dE0RJCMY2_2),.dout(w_dff_B_BnSvBPJn0_2),.clk(gclk));
	jdff dff_B_a5JaWE737_2(.din(w_dff_B_BnSvBPJn0_2),.dout(w_dff_B_a5JaWE737_2),.clk(gclk));
	jdff dff_B_StYRvpWz0_2(.din(n433),.dout(w_dff_B_StYRvpWz0_2),.clk(gclk));
	jdff dff_B_xBcKVmxU9_2(.din(w_dff_B_StYRvpWz0_2),.dout(w_dff_B_xBcKVmxU9_2),.clk(gclk));
	jdff dff_B_Baav93bQ4_2(.din(w_dff_B_xBcKVmxU9_2),.dout(w_dff_B_Baav93bQ4_2),.clk(gclk));
	jdff dff_B_Cecb2C139_1(.din(n419),.dout(w_dff_B_Cecb2C139_1),.clk(gclk));
	jdff dff_B_LhXZKNt04_1(.din(w_dff_B_Cecb2C139_1),.dout(w_dff_B_LhXZKNt04_1),.clk(gclk));
	jdff dff_B_GQQ7GrVa6_2(.din(n356),.dout(w_dff_B_GQQ7GrVa6_2),.clk(gclk));
	jdff dff_B_tssskMr49_2(.din(w_dff_B_GQQ7GrVa6_2),.dout(w_dff_B_tssskMr49_2),.clk(gclk));
	jdff dff_B_XzIhFrPZ0_2(.din(w_dff_B_tssskMr49_2),.dout(w_dff_B_XzIhFrPZ0_2),.clk(gclk));
	jdff dff_B_wHOweIil2_0(.din(n361),.dout(w_dff_B_wHOweIil2_0),.clk(gclk));
	jdff dff_A_kPRBdduK3_0(.dout(w_n297_0[0]),.din(w_dff_A_kPRBdduK3_0),.clk(gclk));
	jdff dff_A_hmDCpiYY5_0(.dout(w_dff_A_kPRBdduK3_0),.din(w_dff_A_hmDCpiYY5_0),.clk(gclk));
	jdff dff_A_ONStMVIT2_1(.dout(w_n297_0[1]),.din(w_dff_A_ONStMVIT2_1),.clk(gclk));
	jdff dff_A_Cqil93OE8_1(.dout(w_dff_A_ONStMVIT2_1),.din(w_dff_A_Cqil93OE8_1),.clk(gclk));
	jdff dff_B_tH64gZ2p2_1(.din(n1594),.dout(w_dff_B_tH64gZ2p2_1),.clk(gclk));
	jdff dff_B_vsBkSVvQ9_2(.din(n1535),.dout(w_dff_B_vsBkSVvQ9_2),.clk(gclk));
	jdff dff_B_YDKIcx736_2(.din(w_dff_B_vsBkSVvQ9_2),.dout(w_dff_B_YDKIcx736_2),.clk(gclk));
	jdff dff_B_wiQ12gCq0_2(.din(w_dff_B_YDKIcx736_2),.dout(w_dff_B_wiQ12gCq0_2),.clk(gclk));
	jdff dff_B_bc7mP5u12_2(.din(w_dff_B_wiQ12gCq0_2),.dout(w_dff_B_bc7mP5u12_2),.clk(gclk));
	jdff dff_B_pJwiY3L16_2(.din(w_dff_B_bc7mP5u12_2),.dout(w_dff_B_pJwiY3L16_2),.clk(gclk));
	jdff dff_B_CfVTyzbr7_2(.din(w_dff_B_pJwiY3L16_2),.dout(w_dff_B_CfVTyzbr7_2),.clk(gclk));
	jdff dff_B_3nC7AJco0_2(.din(w_dff_B_CfVTyzbr7_2),.dout(w_dff_B_3nC7AJco0_2),.clk(gclk));
	jdff dff_B_z5Zy6f9Q3_2(.din(w_dff_B_3nC7AJco0_2),.dout(w_dff_B_z5Zy6f9Q3_2),.clk(gclk));
	jdff dff_B_JiiRaLyT6_2(.din(w_dff_B_z5Zy6f9Q3_2),.dout(w_dff_B_JiiRaLyT6_2),.clk(gclk));
	jdff dff_B_dWWWBkCr0_2(.din(w_dff_B_JiiRaLyT6_2),.dout(w_dff_B_dWWWBkCr0_2),.clk(gclk));
	jdff dff_B_hVJNX2qw9_2(.din(w_dff_B_dWWWBkCr0_2),.dout(w_dff_B_hVJNX2qw9_2),.clk(gclk));
	jdff dff_B_8JGAj5iT2_2(.din(w_dff_B_hVJNX2qw9_2),.dout(w_dff_B_8JGAj5iT2_2),.clk(gclk));
	jdff dff_B_b6KKmoqP2_2(.din(w_dff_B_8JGAj5iT2_2),.dout(w_dff_B_b6KKmoqP2_2),.clk(gclk));
	jdff dff_B_p2xCU6m46_2(.din(w_dff_B_b6KKmoqP2_2),.dout(w_dff_B_p2xCU6m46_2),.clk(gclk));
	jdff dff_B_uJrcZC8F0_2(.din(w_dff_B_p2xCU6m46_2),.dout(w_dff_B_uJrcZC8F0_2),.clk(gclk));
	jdff dff_B_g1fcwlwt0_2(.din(w_dff_B_uJrcZC8F0_2),.dout(w_dff_B_g1fcwlwt0_2),.clk(gclk));
	jdff dff_B_gBggXZDR0_2(.din(w_dff_B_g1fcwlwt0_2),.dout(w_dff_B_gBggXZDR0_2),.clk(gclk));
	jdff dff_B_qYAFNbPN4_2(.din(w_dff_B_gBggXZDR0_2),.dout(w_dff_B_qYAFNbPN4_2),.clk(gclk));
	jdff dff_B_LXBC5JLy0_2(.din(w_dff_B_qYAFNbPN4_2),.dout(w_dff_B_LXBC5JLy0_2),.clk(gclk));
	jdff dff_B_BEpY2dra0_2(.din(w_dff_B_LXBC5JLy0_2),.dout(w_dff_B_BEpY2dra0_2),.clk(gclk));
	jdff dff_B_oNRq0rgT5_2(.din(w_dff_B_BEpY2dra0_2),.dout(w_dff_B_oNRq0rgT5_2),.clk(gclk));
	jdff dff_B_FUrM4H2e0_2(.din(w_dff_B_oNRq0rgT5_2),.dout(w_dff_B_FUrM4H2e0_2),.clk(gclk));
	jdff dff_B_hE4UHJNO5_2(.din(w_dff_B_FUrM4H2e0_2),.dout(w_dff_B_hE4UHJNO5_2),.clk(gclk));
	jdff dff_B_XpKPpW862_2(.din(w_dff_B_hE4UHJNO5_2),.dout(w_dff_B_XpKPpW862_2),.clk(gclk));
	jdff dff_B_Pukwssw95_2(.din(w_dff_B_XpKPpW862_2),.dout(w_dff_B_Pukwssw95_2),.clk(gclk));
	jdff dff_B_iDh9LQAv8_2(.din(w_dff_B_Pukwssw95_2),.dout(w_dff_B_iDh9LQAv8_2),.clk(gclk));
	jdff dff_B_zZ0kqyn91_2(.din(w_dff_B_iDh9LQAv8_2),.dout(w_dff_B_zZ0kqyn91_2),.clk(gclk));
	jdff dff_B_91ISSEBv4_2(.din(w_dff_B_zZ0kqyn91_2),.dout(w_dff_B_91ISSEBv4_2),.clk(gclk));
	jdff dff_B_qPa29pS04_2(.din(w_dff_B_91ISSEBv4_2),.dout(w_dff_B_qPa29pS04_2),.clk(gclk));
	jdff dff_B_kfwyd9nP9_2(.din(w_dff_B_qPa29pS04_2),.dout(w_dff_B_kfwyd9nP9_2),.clk(gclk));
	jdff dff_B_yrxVOoOE8_2(.din(w_dff_B_kfwyd9nP9_2),.dout(w_dff_B_yrxVOoOE8_2),.clk(gclk));
	jdff dff_B_AY7lYIUV9_2(.din(w_dff_B_yrxVOoOE8_2),.dout(w_dff_B_AY7lYIUV9_2),.clk(gclk));
	jdff dff_B_mrrtY6pt7_2(.din(w_dff_B_AY7lYIUV9_2),.dout(w_dff_B_mrrtY6pt7_2),.clk(gclk));
	jdff dff_B_LKQUuxjj8_2(.din(w_dff_B_mrrtY6pt7_2),.dout(w_dff_B_LKQUuxjj8_2),.clk(gclk));
	jdff dff_B_1kTDukAs5_2(.din(w_dff_B_LKQUuxjj8_2),.dout(w_dff_B_1kTDukAs5_2),.clk(gclk));
	jdff dff_B_hUXzn7KH6_2(.din(w_dff_B_1kTDukAs5_2),.dout(w_dff_B_hUXzn7KH6_2),.clk(gclk));
	jdff dff_B_njlmG7O59_2(.din(w_dff_B_hUXzn7KH6_2),.dout(w_dff_B_njlmG7O59_2),.clk(gclk));
	jdff dff_B_POyDQKv68_2(.din(w_dff_B_njlmG7O59_2),.dout(w_dff_B_POyDQKv68_2),.clk(gclk));
	jdff dff_B_4EvScwfw9_2(.din(w_dff_B_POyDQKv68_2),.dout(w_dff_B_4EvScwfw9_2),.clk(gclk));
	jdff dff_B_Th3njhLC2_2(.din(w_dff_B_4EvScwfw9_2),.dout(w_dff_B_Th3njhLC2_2),.clk(gclk));
	jdff dff_B_w1gSjeAf4_2(.din(w_dff_B_Th3njhLC2_2),.dout(w_dff_B_w1gSjeAf4_2),.clk(gclk));
	jdff dff_B_OsKlf9aE8_2(.din(w_dff_B_w1gSjeAf4_2),.dout(w_dff_B_OsKlf9aE8_2),.clk(gclk));
	jdff dff_B_2lysxwuL8_2(.din(w_dff_B_OsKlf9aE8_2),.dout(w_dff_B_2lysxwuL8_2),.clk(gclk));
	jdff dff_B_NUZsT6f97_2(.din(w_dff_B_2lysxwuL8_2),.dout(w_dff_B_NUZsT6f97_2),.clk(gclk));
	jdff dff_B_ulbJp4165_2(.din(w_dff_B_NUZsT6f97_2),.dout(w_dff_B_ulbJp4165_2),.clk(gclk));
	jdff dff_B_ERHUrecI3_2(.din(w_dff_B_ulbJp4165_2),.dout(w_dff_B_ERHUrecI3_2),.clk(gclk));
	jdff dff_B_gnw9YzMm7_0(.din(n1593),.dout(w_dff_B_gnw9YzMm7_0),.clk(gclk));
	jdff dff_A_0VYyg8st6_1(.dout(w_n1581_0[1]),.din(w_dff_A_0VYyg8st6_1),.clk(gclk));
	jdff dff_B_mEub8Cht3_1(.din(n1536),.dout(w_dff_B_mEub8Cht3_1),.clk(gclk));
	jdff dff_B_04aaA9Pj2_2(.din(n1471),.dout(w_dff_B_04aaA9Pj2_2),.clk(gclk));
	jdff dff_B_uGPEyDWy3_2(.din(w_dff_B_04aaA9Pj2_2),.dout(w_dff_B_uGPEyDWy3_2),.clk(gclk));
	jdff dff_B_Jw4gCK698_2(.din(w_dff_B_uGPEyDWy3_2),.dout(w_dff_B_Jw4gCK698_2),.clk(gclk));
	jdff dff_B_4MHLehCB7_2(.din(w_dff_B_Jw4gCK698_2),.dout(w_dff_B_4MHLehCB7_2),.clk(gclk));
	jdff dff_B_mho9pv3N5_2(.din(w_dff_B_4MHLehCB7_2),.dout(w_dff_B_mho9pv3N5_2),.clk(gclk));
	jdff dff_B_9cKZPClz3_2(.din(w_dff_B_mho9pv3N5_2),.dout(w_dff_B_9cKZPClz3_2),.clk(gclk));
	jdff dff_B_aL7DujUi5_2(.din(w_dff_B_9cKZPClz3_2),.dout(w_dff_B_aL7DujUi5_2),.clk(gclk));
	jdff dff_B_WNed0ixx4_2(.din(w_dff_B_aL7DujUi5_2),.dout(w_dff_B_WNed0ixx4_2),.clk(gclk));
	jdff dff_B_RlHJfAZj3_2(.din(w_dff_B_WNed0ixx4_2),.dout(w_dff_B_RlHJfAZj3_2),.clk(gclk));
	jdff dff_B_OXey3Q4g5_2(.din(w_dff_B_RlHJfAZj3_2),.dout(w_dff_B_OXey3Q4g5_2),.clk(gclk));
	jdff dff_B_Fb4TIpvM9_2(.din(w_dff_B_OXey3Q4g5_2),.dout(w_dff_B_Fb4TIpvM9_2),.clk(gclk));
	jdff dff_B_hvDhxpSV8_2(.din(w_dff_B_Fb4TIpvM9_2),.dout(w_dff_B_hvDhxpSV8_2),.clk(gclk));
	jdff dff_B_IlmlciXJ9_2(.din(w_dff_B_hvDhxpSV8_2),.dout(w_dff_B_IlmlciXJ9_2),.clk(gclk));
	jdff dff_B_NU3PDFub9_2(.din(w_dff_B_IlmlciXJ9_2),.dout(w_dff_B_NU3PDFub9_2),.clk(gclk));
	jdff dff_B_kjDWGwKC5_2(.din(w_dff_B_NU3PDFub9_2),.dout(w_dff_B_kjDWGwKC5_2),.clk(gclk));
	jdff dff_B_5EXv2p1d4_2(.din(w_dff_B_kjDWGwKC5_2),.dout(w_dff_B_5EXv2p1d4_2),.clk(gclk));
	jdff dff_B_f1JfoURg7_2(.din(w_dff_B_5EXv2p1d4_2),.dout(w_dff_B_f1JfoURg7_2),.clk(gclk));
	jdff dff_B_VRDgX8f18_2(.din(w_dff_B_f1JfoURg7_2),.dout(w_dff_B_VRDgX8f18_2),.clk(gclk));
	jdff dff_B_GZkdl9En5_2(.din(w_dff_B_VRDgX8f18_2),.dout(w_dff_B_GZkdl9En5_2),.clk(gclk));
	jdff dff_B_I8KzF8wc2_2(.din(w_dff_B_GZkdl9En5_2),.dout(w_dff_B_I8KzF8wc2_2),.clk(gclk));
	jdff dff_B_gaRqe6bL1_2(.din(w_dff_B_I8KzF8wc2_2),.dout(w_dff_B_gaRqe6bL1_2),.clk(gclk));
	jdff dff_B_kkHFDaT97_2(.din(w_dff_B_gaRqe6bL1_2),.dout(w_dff_B_kkHFDaT97_2),.clk(gclk));
	jdff dff_B_SLCXx6yq3_2(.din(w_dff_B_kkHFDaT97_2),.dout(w_dff_B_SLCXx6yq3_2),.clk(gclk));
	jdff dff_B_CIHttLD85_2(.din(w_dff_B_SLCXx6yq3_2),.dout(w_dff_B_CIHttLD85_2),.clk(gclk));
	jdff dff_B_LAMs7jrJ3_2(.din(w_dff_B_CIHttLD85_2),.dout(w_dff_B_LAMs7jrJ3_2),.clk(gclk));
	jdff dff_B_Qp8Tv7Y91_2(.din(w_dff_B_LAMs7jrJ3_2),.dout(w_dff_B_Qp8Tv7Y91_2),.clk(gclk));
	jdff dff_B_oeu70c2d3_2(.din(w_dff_B_Qp8Tv7Y91_2),.dout(w_dff_B_oeu70c2d3_2),.clk(gclk));
	jdff dff_B_QyTblDHL5_2(.din(w_dff_B_oeu70c2d3_2),.dout(w_dff_B_QyTblDHL5_2),.clk(gclk));
	jdff dff_B_YqwMphmv2_2(.din(w_dff_B_QyTblDHL5_2),.dout(w_dff_B_YqwMphmv2_2),.clk(gclk));
	jdff dff_B_pC1cg0cG3_2(.din(w_dff_B_YqwMphmv2_2),.dout(w_dff_B_pC1cg0cG3_2),.clk(gclk));
	jdff dff_B_D3KQpFdg0_2(.din(w_dff_B_pC1cg0cG3_2),.dout(w_dff_B_D3KQpFdg0_2),.clk(gclk));
	jdff dff_B_gDvfvCPO2_2(.din(w_dff_B_D3KQpFdg0_2),.dout(w_dff_B_gDvfvCPO2_2),.clk(gclk));
	jdff dff_B_zJAf4Cmw7_2(.din(w_dff_B_gDvfvCPO2_2),.dout(w_dff_B_zJAf4Cmw7_2),.clk(gclk));
	jdff dff_B_IpZCzPRt6_2(.din(w_dff_B_zJAf4Cmw7_2),.dout(w_dff_B_IpZCzPRt6_2),.clk(gclk));
	jdff dff_B_en0pEEKL1_2(.din(w_dff_B_IpZCzPRt6_2),.dout(w_dff_B_en0pEEKL1_2),.clk(gclk));
	jdff dff_B_wsaxXHHs7_2(.din(w_dff_B_en0pEEKL1_2),.dout(w_dff_B_wsaxXHHs7_2),.clk(gclk));
	jdff dff_B_IUhOhLE62_2(.din(w_dff_B_wsaxXHHs7_2),.dout(w_dff_B_IUhOhLE62_2),.clk(gclk));
	jdff dff_B_jTOsY1Br4_2(.din(w_dff_B_IUhOhLE62_2),.dout(w_dff_B_jTOsY1Br4_2),.clk(gclk));
	jdff dff_B_t6m14mr58_2(.din(w_dff_B_jTOsY1Br4_2),.dout(w_dff_B_t6m14mr58_2),.clk(gclk));
	jdff dff_B_7I4L68L81_2(.din(w_dff_B_t6m14mr58_2),.dout(w_dff_B_7I4L68L81_2),.clk(gclk));
	jdff dff_B_q3UgyzgI7_2(.din(w_dff_B_7I4L68L81_2),.dout(w_dff_B_q3UgyzgI7_2),.clk(gclk));
	jdff dff_B_LidCqk3d7_2(.din(n1517),.dout(w_dff_B_LidCqk3d7_2),.clk(gclk));
	jdff dff_B_0Um9Rg9s4_1(.din(n1472),.dout(w_dff_B_0Um9Rg9s4_1),.clk(gclk));
	jdff dff_B_FYeqss1r8_2(.din(n1400),.dout(w_dff_B_FYeqss1r8_2),.clk(gclk));
	jdff dff_B_0W5GxR8j8_2(.din(w_dff_B_FYeqss1r8_2),.dout(w_dff_B_0W5GxR8j8_2),.clk(gclk));
	jdff dff_B_NEVodtvL7_2(.din(w_dff_B_0W5GxR8j8_2),.dout(w_dff_B_NEVodtvL7_2),.clk(gclk));
	jdff dff_B_dS7nhfoN4_2(.din(w_dff_B_NEVodtvL7_2),.dout(w_dff_B_dS7nhfoN4_2),.clk(gclk));
	jdff dff_B_DxMaCaeA6_2(.din(w_dff_B_dS7nhfoN4_2),.dout(w_dff_B_DxMaCaeA6_2),.clk(gclk));
	jdff dff_B_4DuoXHBK1_2(.din(w_dff_B_DxMaCaeA6_2),.dout(w_dff_B_4DuoXHBK1_2),.clk(gclk));
	jdff dff_B_xnHIWkkX9_2(.din(w_dff_B_4DuoXHBK1_2),.dout(w_dff_B_xnHIWkkX9_2),.clk(gclk));
	jdff dff_B_OguhmY5w5_2(.din(w_dff_B_xnHIWkkX9_2),.dout(w_dff_B_OguhmY5w5_2),.clk(gclk));
	jdff dff_B_lrRq2WNd1_2(.din(w_dff_B_OguhmY5w5_2),.dout(w_dff_B_lrRq2WNd1_2),.clk(gclk));
	jdff dff_B_LUS16xPf8_2(.din(w_dff_B_lrRq2WNd1_2),.dout(w_dff_B_LUS16xPf8_2),.clk(gclk));
	jdff dff_B_0c9zDrv27_2(.din(w_dff_B_LUS16xPf8_2),.dout(w_dff_B_0c9zDrv27_2),.clk(gclk));
	jdff dff_B_2lR4bZBX6_2(.din(w_dff_B_0c9zDrv27_2),.dout(w_dff_B_2lR4bZBX6_2),.clk(gclk));
	jdff dff_B_KgCCofJ52_2(.din(w_dff_B_2lR4bZBX6_2),.dout(w_dff_B_KgCCofJ52_2),.clk(gclk));
	jdff dff_B_VJZliVqm8_2(.din(w_dff_B_KgCCofJ52_2),.dout(w_dff_B_VJZliVqm8_2),.clk(gclk));
	jdff dff_B_pbKSCjGs5_2(.din(w_dff_B_VJZliVqm8_2),.dout(w_dff_B_pbKSCjGs5_2),.clk(gclk));
	jdff dff_B_XnRPovyT7_2(.din(w_dff_B_pbKSCjGs5_2),.dout(w_dff_B_XnRPovyT7_2),.clk(gclk));
	jdff dff_B_u0kxdFDU7_2(.din(w_dff_B_XnRPovyT7_2),.dout(w_dff_B_u0kxdFDU7_2),.clk(gclk));
	jdff dff_B_MNcbHyEE3_2(.din(w_dff_B_u0kxdFDU7_2),.dout(w_dff_B_MNcbHyEE3_2),.clk(gclk));
	jdff dff_B_Q4OwdjlL3_2(.din(w_dff_B_MNcbHyEE3_2),.dout(w_dff_B_Q4OwdjlL3_2),.clk(gclk));
	jdff dff_B_o4bAO1UA8_2(.din(w_dff_B_Q4OwdjlL3_2),.dout(w_dff_B_o4bAO1UA8_2),.clk(gclk));
	jdff dff_B_bBxnxwqF7_2(.din(w_dff_B_o4bAO1UA8_2),.dout(w_dff_B_bBxnxwqF7_2),.clk(gclk));
	jdff dff_B_nCngdcef7_2(.din(w_dff_B_bBxnxwqF7_2),.dout(w_dff_B_nCngdcef7_2),.clk(gclk));
	jdff dff_B_b1sbFnIp3_2(.din(w_dff_B_nCngdcef7_2),.dout(w_dff_B_b1sbFnIp3_2),.clk(gclk));
	jdff dff_B_Z51BpY3j1_2(.din(w_dff_B_b1sbFnIp3_2),.dout(w_dff_B_Z51BpY3j1_2),.clk(gclk));
	jdff dff_B_g0EJDHDJ5_2(.din(w_dff_B_Z51BpY3j1_2),.dout(w_dff_B_g0EJDHDJ5_2),.clk(gclk));
	jdff dff_B_4gtwUJOe7_2(.din(w_dff_B_g0EJDHDJ5_2),.dout(w_dff_B_4gtwUJOe7_2),.clk(gclk));
	jdff dff_B_XGXJ9S162_2(.din(w_dff_B_4gtwUJOe7_2),.dout(w_dff_B_XGXJ9S162_2),.clk(gclk));
	jdff dff_B_lqSVTLqO9_2(.din(w_dff_B_XGXJ9S162_2),.dout(w_dff_B_lqSVTLqO9_2),.clk(gclk));
	jdff dff_B_1ccNLfBt2_2(.din(w_dff_B_lqSVTLqO9_2),.dout(w_dff_B_1ccNLfBt2_2),.clk(gclk));
	jdff dff_B_ySeAm6lW3_2(.din(w_dff_B_1ccNLfBt2_2),.dout(w_dff_B_ySeAm6lW3_2),.clk(gclk));
	jdff dff_B_Tma7Mkyr4_2(.din(w_dff_B_ySeAm6lW3_2),.dout(w_dff_B_Tma7Mkyr4_2),.clk(gclk));
	jdff dff_B_ry4mptlp7_2(.din(w_dff_B_Tma7Mkyr4_2),.dout(w_dff_B_ry4mptlp7_2),.clk(gclk));
	jdff dff_B_Y7zLzYTy3_2(.din(w_dff_B_ry4mptlp7_2),.dout(w_dff_B_Y7zLzYTy3_2),.clk(gclk));
	jdff dff_B_20eYAsih1_2(.din(w_dff_B_Y7zLzYTy3_2),.dout(w_dff_B_20eYAsih1_2),.clk(gclk));
	jdff dff_B_WyUNR5Ew3_2(.din(w_dff_B_20eYAsih1_2),.dout(w_dff_B_WyUNR5Ew3_2),.clk(gclk));
	jdff dff_B_P6uXQ72v4_2(.din(w_dff_B_WyUNR5Ew3_2),.dout(w_dff_B_P6uXQ72v4_2),.clk(gclk));
	jdff dff_B_oSg6BDzv9_2(.din(w_dff_B_P6uXQ72v4_2),.dout(w_dff_B_oSg6BDzv9_2),.clk(gclk));
	jdff dff_B_i3Ve0M2d3_2(.din(w_dff_B_oSg6BDzv9_2),.dout(w_dff_B_i3Ve0M2d3_2),.clk(gclk));
	jdff dff_B_389B8GSI6_2(.din(n1446),.dout(w_dff_B_389B8GSI6_2),.clk(gclk));
	jdff dff_B_EEFDNy893_1(.din(n1401),.dout(w_dff_B_EEFDNy893_1),.clk(gclk));
	jdff dff_B_9McnlYsm1_2(.din(n1322),.dout(w_dff_B_9McnlYsm1_2),.clk(gclk));
	jdff dff_B_pKf1HR1x4_2(.din(w_dff_B_9McnlYsm1_2),.dout(w_dff_B_pKf1HR1x4_2),.clk(gclk));
	jdff dff_B_ZzQzMXrZ2_2(.din(w_dff_B_pKf1HR1x4_2),.dout(w_dff_B_ZzQzMXrZ2_2),.clk(gclk));
	jdff dff_B_rFb84YWB2_2(.din(w_dff_B_ZzQzMXrZ2_2),.dout(w_dff_B_rFb84YWB2_2),.clk(gclk));
	jdff dff_B_7nHviEfH9_2(.din(w_dff_B_rFb84YWB2_2),.dout(w_dff_B_7nHviEfH9_2),.clk(gclk));
	jdff dff_B_81ooFWeb5_2(.din(w_dff_B_7nHviEfH9_2),.dout(w_dff_B_81ooFWeb5_2),.clk(gclk));
	jdff dff_B_YoHzIqbB8_2(.din(w_dff_B_81ooFWeb5_2),.dout(w_dff_B_YoHzIqbB8_2),.clk(gclk));
	jdff dff_B_1ydIIUHn3_2(.din(w_dff_B_YoHzIqbB8_2),.dout(w_dff_B_1ydIIUHn3_2),.clk(gclk));
	jdff dff_B_s5ig4Y2j8_2(.din(w_dff_B_1ydIIUHn3_2),.dout(w_dff_B_s5ig4Y2j8_2),.clk(gclk));
	jdff dff_B_rNt2kuqR7_2(.din(w_dff_B_s5ig4Y2j8_2),.dout(w_dff_B_rNt2kuqR7_2),.clk(gclk));
	jdff dff_B_CgeR1ohU2_2(.din(w_dff_B_rNt2kuqR7_2),.dout(w_dff_B_CgeR1ohU2_2),.clk(gclk));
	jdff dff_B_0kXB4qhL2_2(.din(w_dff_B_CgeR1ohU2_2),.dout(w_dff_B_0kXB4qhL2_2),.clk(gclk));
	jdff dff_B_KB8LWmM05_2(.din(w_dff_B_0kXB4qhL2_2),.dout(w_dff_B_KB8LWmM05_2),.clk(gclk));
	jdff dff_B_WiRQ99eB1_2(.din(w_dff_B_KB8LWmM05_2),.dout(w_dff_B_WiRQ99eB1_2),.clk(gclk));
	jdff dff_B_suPLVpzt2_2(.din(w_dff_B_WiRQ99eB1_2),.dout(w_dff_B_suPLVpzt2_2),.clk(gclk));
	jdff dff_B_XNBJe3SD3_2(.din(w_dff_B_suPLVpzt2_2),.dout(w_dff_B_XNBJe3SD3_2),.clk(gclk));
	jdff dff_B_2Jcdb9cm1_2(.din(w_dff_B_XNBJe3SD3_2),.dout(w_dff_B_2Jcdb9cm1_2),.clk(gclk));
	jdff dff_B_SxIBpEx52_2(.din(w_dff_B_2Jcdb9cm1_2),.dout(w_dff_B_SxIBpEx52_2),.clk(gclk));
	jdff dff_B_xp7BD0NP4_2(.din(w_dff_B_SxIBpEx52_2),.dout(w_dff_B_xp7BD0NP4_2),.clk(gclk));
	jdff dff_B_fKc2By9A8_2(.din(w_dff_B_xp7BD0NP4_2),.dout(w_dff_B_fKc2By9A8_2),.clk(gclk));
	jdff dff_B_x1gpd9tU7_2(.din(w_dff_B_fKc2By9A8_2),.dout(w_dff_B_x1gpd9tU7_2),.clk(gclk));
	jdff dff_B_KWAnneZX5_2(.din(w_dff_B_x1gpd9tU7_2),.dout(w_dff_B_KWAnneZX5_2),.clk(gclk));
	jdff dff_B_pK1bjzOe0_2(.din(w_dff_B_KWAnneZX5_2),.dout(w_dff_B_pK1bjzOe0_2),.clk(gclk));
	jdff dff_B_qKvLM4Iq3_2(.din(w_dff_B_pK1bjzOe0_2),.dout(w_dff_B_qKvLM4Iq3_2),.clk(gclk));
	jdff dff_B_nhlIYQLz9_2(.din(w_dff_B_qKvLM4Iq3_2),.dout(w_dff_B_nhlIYQLz9_2),.clk(gclk));
	jdff dff_B_JB3bG6Ez7_2(.din(w_dff_B_nhlIYQLz9_2),.dout(w_dff_B_JB3bG6Ez7_2),.clk(gclk));
	jdff dff_B_rE2btYBL6_2(.din(w_dff_B_JB3bG6Ez7_2),.dout(w_dff_B_rE2btYBL6_2),.clk(gclk));
	jdff dff_B_jamFC7LZ3_2(.din(w_dff_B_rE2btYBL6_2),.dout(w_dff_B_jamFC7LZ3_2),.clk(gclk));
	jdff dff_B_4FG32wZ97_2(.din(w_dff_B_jamFC7LZ3_2),.dout(w_dff_B_4FG32wZ97_2),.clk(gclk));
	jdff dff_B_sh2kcuiY3_2(.din(w_dff_B_4FG32wZ97_2),.dout(w_dff_B_sh2kcuiY3_2),.clk(gclk));
	jdff dff_B_Cwv5OEyC3_2(.din(w_dff_B_sh2kcuiY3_2),.dout(w_dff_B_Cwv5OEyC3_2),.clk(gclk));
	jdff dff_B_E6RTjQmc2_2(.din(w_dff_B_Cwv5OEyC3_2),.dout(w_dff_B_E6RTjQmc2_2),.clk(gclk));
	jdff dff_B_b5uOftRa7_2(.din(w_dff_B_E6RTjQmc2_2),.dout(w_dff_B_b5uOftRa7_2),.clk(gclk));
	jdff dff_B_m4B0bsaM0_2(.din(w_dff_B_b5uOftRa7_2),.dout(w_dff_B_m4B0bsaM0_2),.clk(gclk));
	jdff dff_B_sJDrkbVR3_2(.din(w_dff_B_m4B0bsaM0_2),.dout(w_dff_B_sJDrkbVR3_2),.clk(gclk));
	jdff dff_B_IP2xz7gk6_2(.din(n1368),.dout(w_dff_B_IP2xz7gk6_2),.clk(gclk));
	jdff dff_B_8fyuWS3C8_1(.din(n1323),.dout(w_dff_B_8fyuWS3C8_1),.clk(gclk));
	jdff dff_B_CZ4lnBnU4_2(.din(n1237),.dout(w_dff_B_CZ4lnBnU4_2),.clk(gclk));
	jdff dff_B_uJTWmKKg9_2(.din(w_dff_B_CZ4lnBnU4_2),.dout(w_dff_B_uJTWmKKg9_2),.clk(gclk));
	jdff dff_B_W8kdiqNn7_2(.din(w_dff_B_uJTWmKKg9_2),.dout(w_dff_B_W8kdiqNn7_2),.clk(gclk));
	jdff dff_B_DMpF30di2_2(.din(w_dff_B_W8kdiqNn7_2),.dout(w_dff_B_DMpF30di2_2),.clk(gclk));
	jdff dff_B_jObhIa4m8_2(.din(w_dff_B_DMpF30di2_2),.dout(w_dff_B_jObhIa4m8_2),.clk(gclk));
	jdff dff_B_DkXtiUhh5_2(.din(w_dff_B_jObhIa4m8_2),.dout(w_dff_B_DkXtiUhh5_2),.clk(gclk));
	jdff dff_B_3AZzWK5K9_2(.din(w_dff_B_DkXtiUhh5_2),.dout(w_dff_B_3AZzWK5K9_2),.clk(gclk));
	jdff dff_B_RB8EGyzc3_2(.din(w_dff_B_3AZzWK5K9_2),.dout(w_dff_B_RB8EGyzc3_2),.clk(gclk));
	jdff dff_B_2Rkc27738_2(.din(w_dff_B_RB8EGyzc3_2),.dout(w_dff_B_2Rkc27738_2),.clk(gclk));
	jdff dff_B_8bct5HR39_2(.din(w_dff_B_2Rkc27738_2),.dout(w_dff_B_8bct5HR39_2),.clk(gclk));
	jdff dff_B_TTeqG0FQ9_2(.din(w_dff_B_8bct5HR39_2),.dout(w_dff_B_TTeqG0FQ9_2),.clk(gclk));
	jdff dff_B_blGsaODc0_2(.din(w_dff_B_TTeqG0FQ9_2),.dout(w_dff_B_blGsaODc0_2),.clk(gclk));
	jdff dff_B_dC8F7YR52_2(.din(w_dff_B_blGsaODc0_2),.dout(w_dff_B_dC8F7YR52_2),.clk(gclk));
	jdff dff_B_0CWn7SjJ2_2(.din(w_dff_B_dC8F7YR52_2),.dout(w_dff_B_0CWn7SjJ2_2),.clk(gclk));
	jdff dff_B_nwh0I2Wz3_2(.din(w_dff_B_0CWn7SjJ2_2),.dout(w_dff_B_nwh0I2Wz3_2),.clk(gclk));
	jdff dff_B_RUdayj0h1_2(.din(w_dff_B_nwh0I2Wz3_2),.dout(w_dff_B_RUdayj0h1_2),.clk(gclk));
	jdff dff_B_0taMoH0W1_2(.din(w_dff_B_RUdayj0h1_2),.dout(w_dff_B_0taMoH0W1_2),.clk(gclk));
	jdff dff_B_N06HOcfl0_2(.din(w_dff_B_0taMoH0W1_2),.dout(w_dff_B_N06HOcfl0_2),.clk(gclk));
	jdff dff_B_S6kSeQDQ7_2(.din(w_dff_B_N06HOcfl0_2),.dout(w_dff_B_S6kSeQDQ7_2),.clk(gclk));
	jdff dff_B_TnDkHids0_2(.din(w_dff_B_S6kSeQDQ7_2),.dout(w_dff_B_TnDkHids0_2),.clk(gclk));
	jdff dff_B_QcMnnVQb5_2(.din(w_dff_B_TnDkHids0_2),.dout(w_dff_B_QcMnnVQb5_2),.clk(gclk));
	jdff dff_B_LZyd5xTg3_2(.din(w_dff_B_QcMnnVQb5_2),.dout(w_dff_B_LZyd5xTg3_2),.clk(gclk));
	jdff dff_B_jpyCYVHf7_2(.din(w_dff_B_LZyd5xTg3_2),.dout(w_dff_B_jpyCYVHf7_2),.clk(gclk));
	jdff dff_B_clxmQnR12_2(.din(w_dff_B_jpyCYVHf7_2),.dout(w_dff_B_clxmQnR12_2),.clk(gclk));
	jdff dff_B_tSSBfNa53_2(.din(w_dff_B_clxmQnR12_2),.dout(w_dff_B_tSSBfNa53_2),.clk(gclk));
	jdff dff_B_EMA8cHjx2_2(.din(w_dff_B_tSSBfNa53_2),.dout(w_dff_B_EMA8cHjx2_2),.clk(gclk));
	jdff dff_B_vPuxReyu7_2(.din(w_dff_B_EMA8cHjx2_2),.dout(w_dff_B_vPuxReyu7_2),.clk(gclk));
	jdff dff_B_WpTXQUJm7_2(.din(w_dff_B_vPuxReyu7_2),.dout(w_dff_B_WpTXQUJm7_2),.clk(gclk));
	jdff dff_B_ZwD6HCR57_2(.din(w_dff_B_WpTXQUJm7_2),.dout(w_dff_B_ZwD6HCR57_2),.clk(gclk));
	jdff dff_B_ywKQgdwa4_2(.din(w_dff_B_ZwD6HCR57_2),.dout(w_dff_B_ywKQgdwa4_2),.clk(gclk));
	jdff dff_B_j0Buq58s5_2(.din(w_dff_B_ywKQgdwa4_2),.dout(w_dff_B_j0Buq58s5_2),.clk(gclk));
	jdff dff_B_yeqhcbgU8_2(.din(w_dff_B_j0Buq58s5_2),.dout(w_dff_B_yeqhcbgU8_2),.clk(gclk));
	jdff dff_B_rRpQxRXk6_2(.din(n1283),.dout(w_dff_B_rRpQxRXk6_2),.clk(gclk));
	jdff dff_B_CsyphyLd6_1(.din(n1238),.dout(w_dff_B_CsyphyLd6_1),.clk(gclk));
	jdff dff_B_hwIpHyGz5_2(.din(n1146),.dout(w_dff_B_hwIpHyGz5_2),.clk(gclk));
	jdff dff_B_JaLNPF1R5_2(.din(w_dff_B_hwIpHyGz5_2),.dout(w_dff_B_JaLNPF1R5_2),.clk(gclk));
	jdff dff_B_Zoz5qMIX0_2(.din(w_dff_B_JaLNPF1R5_2),.dout(w_dff_B_Zoz5qMIX0_2),.clk(gclk));
	jdff dff_B_3WYuB6Xe5_2(.din(w_dff_B_Zoz5qMIX0_2),.dout(w_dff_B_3WYuB6Xe5_2),.clk(gclk));
	jdff dff_B_O26byoBL3_2(.din(w_dff_B_3WYuB6Xe5_2),.dout(w_dff_B_O26byoBL3_2),.clk(gclk));
	jdff dff_B_Wq22OHV66_2(.din(w_dff_B_O26byoBL3_2),.dout(w_dff_B_Wq22OHV66_2),.clk(gclk));
	jdff dff_B_OMek1LYa7_2(.din(w_dff_B_Wq22OHV66_2),.dout(w_dff_B_OMek1LYa7_2),.clk(gclk));
	jdff dff_B_umbRiCSr6_2(.din(w_dff_B_OMek1LYa7_2),.dout(w_dff_B_umbRiCSr6_2),.clk(gclk));
	jdff dff_B_rLrmj8R86_2(.din(w_dff_B_umbRiCSr6_2),.dout(w_dff_B_rLrmj8R86_2),.clk(gclk));
	jdff dff_B_TGZvNaf38_2(.din(w_dff_B_rLrmj8R86_2),.dout(w_dff_B_TGZvNaf38_2),.clk(gclk));
	jdff dff_B_L6VddQaT1_2(.din(w_dff_B_TGZvNaf38_2),.dout(w_dff_B_L6VddQaT1_2),.clk(gclk));
	jdff dff_B_IeuTQqpa0_2(.din(w_dff_B_L6VddQaT1_2),.dout(w_dff_B_IeuTQqpa0_2),.clk(gclk));
	jdff dff_B_bMmCb6Ng6_2(.din(w_dff_B_IeuTQqpa0_2),.dout(w_dff_B_bMmCb6Ng6_2),.clk(gclk));
	jdff dff_B_3ObcaEG11_2(.din(w_dff_B_bMmCb6Ng6_2),.dout(w_dff_B_3ObcaEG11_2),.clk(gclk));
	jdff dff_B_1Nz5Iy0p0_2(.din(w_dff_B_3ObcaEG11_2),.dout(w_dff_B_1Nz5Iy0p0_2),.clk(gclk));
	jdff dff_B_I8eRL6Ot3_2(.din(w_dff_B_1Nz5Iy0p0_2),.dout(w_dff_B_I8eRL6Ot3_2),.clk(gclk));
	jdff dff_B_tlWbOF6S3_2(.din(w_dff_B_I8eRL6Ot3_2),.dout(w_dff_B_tlWbOF6S3_2),.clk(gclk));
	jdff dff_B_JkJ5zbY76_2(.din(w_dff_B_tlWbOF6S3_2),.dout(w_dff_B_JkJ5zbY76_2),.clk(gclk));
	jdff dff_B_vJoA67bg3_2(.din(w_dff_B_JkJ5zbY76_2),.dout(w_dff_B_vJoA67bg3_2),.clk(gclk));
	jdff dff_B_8zk7mE1u7_2(.din(w_dff_B_vJoA67bg3_2),.dout(w_dff_B_8zk7mE1u7_2),.clk(gclk));
	jdff dff_B_4XKKqanO3_2(.din(w_dff_B_8zk7mE1u7_2),.dout(w_dff_B_4XKKqanO3_2),.clk(gclk));
	jdff dff_B_4rGBuJul6_2(.din(w_dff_B_4XKKqanO3_2),.dout(w_dff_B_4rGBuJul6_2),.clk(gclk));
	jdff dff_B_bEemoxrx1_2(.din(w_dff_B_4rGBuJul6_2),.dout(w_dff_B_bEemoxrx1_2),.clk(gclk));
	jdff dff_B_xrQzQvAZ3_2(.din(w_dff_B_bEemoxrx1_2),.dout(w_dff_B_xrQzQvAZ3_2),.clk(gclk));
	jdff dff_B_gtHlNTOL7_2(.din(w_dff_B_xrQzQvAZ3_2),.dout(w_dff_B_gtHlNTOL7_2),.clk(gclk));
	jdff dff_B_mwnWALYY4_2(.din(w_dff_B_gtHlNTOL7_2),.dout(w_dff_B_mwnWALYY4_2),.clk(gclk));
	jdff dff_B_6rzBcZzE7_2(.din(w_dff_B_mwnWALYY4_2),.dout(w_dff_B_6rzBcZzE7_2),.clk(gclk));
	jdff dff_B_eGjzVzzH4_2(.din(w_dff_B_6rzBcZzE7_2),.dout(w_dff_B_eGjzVzzH4_2),.clk(gclk));
	jdff dff_B_95Ba9HeD1_2(.din(w_dff_B_eGjzVzzH4_2),.dout(w_dff_B_95Ba9HeD1_2),.clk(gclk));
	jdff dff_B_Hv6YVCsr6_2(.din(n1192),.dout(w_dff_B_Hv6YVCsr6_2),.clk(gclk));
	jdff dff_B_LQq7XSgV1_1(.din(n1147),.dout(w_dff_B_LQq7XSgV1_1),.clk(gclk));
	jdff dff_B_vcJIzG6e5_2(.din(n1048),.dout(w_dff_B_vcJIzG6e5_2),.clk(gclk));
	jdff dff_B_KyAy0u7z2_2(.din(w_dff_B_vcJIzG6e5_2),.dout(w_dff_B_KyAy0u7z2_2),.clk(gclk));
	jdff dff_B_bwFVgsCd8_2(.din(w_dff_B_KyAy0u7z2_2),.dout(w_dff_B_bwFVgsCd8_2),.clk(gclk));
	jdff dff_B_ryv10emY7_2(.din(w_dff_B_bwFVgsCd8_2),.dout(w_dff_B_ryv10emY7_2),.clk(gclk));
	jdff dff_B_QLutS9cy4_2(.din(w_dff_B_ryv10emY7_2),.dout(w_dff_B_QLutS9cy4_2),.clk(gclk));
	jdff dff_B_v9840jYK1_2(.din(w_dff_B_QLutS9cy4_2),.dout(w_dff_B_v9840jYK1_2),.clk(gclk));
	jdff dff_B_BrCgUxQT1_2(.din(w_dff_B_v9840jYK1_2),.dout(w_dff_B_BrCgUxQT1_2),.clk(gclk));
	jdff dff_B_93aRqduI4_2(.din(w_dff_B_BrCgUxQT1_2),.dout(w_dff_B_93aRqduI4_2),.clk(gclk));
	jdff dff_B_PNnW47wB3_2(.din(w_dff_B_93aRqduI4_2),.dout(w_dff_B_PNnW47wB3_2),.clk(gclk));
	jdff dff_B_rbEFlcNa3_2(.din(w_dff_B_PNnW47wB3_2),.dout(w_dff_B_rbEFlcNa3_2),.clk(gclk));
	jdff dff_B_wvnIlnOQ6_2(.din(w_dff_B_rbEFlcNa3_2),.dout(w_dff_B_wvnIlnOQ6_2),.clk(gclk));
	jdff dff_B_Dr87KwPU9_2(.din(w_dff_B_wvnIlnOQ6_2),.dout(w_dff_B_Dr87KwPU9_2),.clk(gclk));
	jdff dff_B_iVVXmieo7_2(.din(w_dff_B_Dr87KwPU9_2),.dout(w_dff_B_iVVXmieo7_2),.clk(gclk));
	jdff dff_B_XlvhNH716_2(.din(w_dff_B_iVVXmieo7_2),.dout(w_dff_B_XlvhNH716_2),.clk(gclk));
	jdff dff_B_AgCiMPqe9_2(.din(w_dff_B_XlvhNH716_2),.dout(w_dff_B_AgCiMPqe9_2),.clk(gclk));
	jdff dff_B_7texvTvg8_2(.din(w_dff_B_AgCiMPqe9_2),.dout(w_dff_B_7texvTvg8_2),.clk(gclk));
	jdff dff_B_hYW46rO79_2(.din(w_dff_B_7texvTvg8_2),.dout(w_dff_B_hYW46rO79_2),.clk(gclk));
	jdff dff_B_tfZRLX5F1_2(.din(w_dff_B_hYW46rO79_2),.dout(w_dff_B_tfZRLX5F1_2),.clk(gclk));
	jdff dff_B_fdfRDlZi0_2(.din(w_dff_B_tfZRLX5F1_2),.dout(w_dff_B_fdfRDlZi0_2),.clk(gclk));
	jdff dff_B_KkekWbYD4_2(.din(w_dff_B_fdfRDlZi0_2),.dout(w_dff_B_KkekWbYD4_2),.clk(gclk));
	jdff dff_B_DA453B0D7_2(.din(w_dff_B_KkekWbYD4_2),.dout(w_dff_B_DA453B0D7_2),.clk(gclk));
	jdff dff_B_Tsr0aNow7_2(.din(w_dff_B_DA453B0D7_2),.dout(w_dff_B_Tsr0aNow7_2),.clk(gclk));
	jdff dff_B_bbOFfDPy5_2(.din(w_dff_B_Tsr0aNow7_2),.dout(w_dff_B_bbOFfDPy5_2),.clk(gclk));
	jdff dff_B_XGlQejHS2_2(.din(w_dff_B_bbOFfDPy5_2),.dout(w_dff_B_XGlQejHS2_2),.clk(gclk));
	jdff dff_B_tpqpxOud6_2(.din(w_dff_B_XGlQejHS2_2),.dout(w_dff_B_tpqpxOud6_2),.clk(gclk));
	jdff dff_B_NgZUA2VO6_2(.din(w_dff_B_tpqpxOud6_2),.dout(w_dff_B_NgZUA2VO6_2),.clk(gclk));
	jdff dff_B_a8DfgMyJ2_2(.din(n1093),.dout(w_dff_B_a8DfgMyJ2_2),.clk(gclk));
	jdff dff_B_VQ99M6Cp9_1(.din(n1049),.dout(w_dff_B_VQ99M6Cp9_1),.clk(gclk));
	jdff dff_B_fLOEm6OU5_2(.din(n949),.dout(w_dff_B_fLOEm6OU5_2),.clk(gclk));
	jdff dff_B_b7EgqpGf5_2(.din(w_dff_B_fLOEm6OU5_2),.dout(w_dff_B_b7EgqpGf5_2),.clk(gclk));
	jdff dff_B_IsKYsYA35_2(.din(w_dff_B_b7EgqpGf5_2),.dout(w_dff_B_IsKYsYA35_2),.clk(gclk));
	jdff dff_B_mmaiWdOm9_2(.din(w_dff_B_IsKYsYA35_2),.dout(w_dff_B_mmaiWdOm9_2),.clk(gclk));
	jdff dff_B_uifbmBo90_2(.din(w_dff_B_mmaiWdOm9_2),.dout(w_dff_B_uifbmBo90_2),.clk(gclk));
	jdff dff_B_VPp2sZDf3_2(.din(w_dff_B_uifbmBo90_2),.dout(w_dff_B_VPp2sZDf3_2),.clk(gclk));
	jdff dff_B_qSggmim50_2(.din(w_dff_B_VPp2sZDf3_2),.dout(w_dff_B_qSggmim50_2),.clk(gclk));
	jdff dff_B_mvAoWqJI4_2(.din(w_dff_B_qSggmim50_2),.dout(w_dff_B_mvAoWqJI4_2),.clk(gclk));
	jdff dff_B_QYgGxJNT9_2(.din(w_dff_B_mvAoWqJI4_2),.dout(w_dff_B_QYgGxJNT9_2),.clk(gclk));
	jdff dff_B_OjC2kcUA2_2(.din(w_dff_B_QYgGxJNT9_2),.dout(w_dff_B_OjC2kcUA2_2),.clk(gclk));
	jdff dff_B_ihnlVSrx3_2(.din(w_dff_B_OjC2kcUA2_2),.dout(w_dff_B_ihnlVSrx3_2),.clk(gclk));
	jdff dff_B_MMmXR79t3_2(.din(w_dff_B_ihnlVSrx3_2),.dout(w_dff_B_MMmXR79t3_2),.clk(gclk));
	jdff dff_B_YZu4mbko4_2(.din(w_dff_B_MMmXR79t3_2),.dout(w_dff_B_YZu4mbko4_2),.clk(gclk));
	jdff dff_B_R2YHob0V1_2(.din(w_dff_B_YZu4mbko4_2),.dout(w_dff_B_R2YHob0V1_2),.clk(gclk));
	jdff dff_B_HGKn9FQW3_2(.din(w_dff_B_R2YHob0V1_2),.dout(w_dff_B_HGKn9FQW3_2),.clk(gclk));
	jdff dff_B_KHbhU1An3_2(.din(w_dff_B_HGKn9FQW3_2),.dout(w_dff_B_KHbhU1An3_2),.clk(gclk));
	jdff dff_B_dfrDS8QZ4_2(.din(w_dff_B_KHbhU1An3_2),.dout(w_dff_B_dfrDS8QZ4_2),.clk(gclk));
	jdff dff_B_VpsGrLNj7_2(.din(w_dff_B_dfrDS8QZ4_2),.dout(w_dff_B_VpsGrLNj7_2),.clk(gclk));
	jdff dff_B_1iysCM1M1_2(.din(w_dff_B_VpsGrLNj7_2),.dout(w_dff_B_1iysCM1M1_2),.clk(gclk));
	jdff dff_B_dbbJhbRE7_2(.din(w_dff_B_1iysCM1M1_2),.dout(w_dff_B_dbbJhbRE7_2),.clk(gclk));
	jdff dff_B_m9jNYSza4_2(.din(w_dff_B_dbbJhbRE7_2),.dout(w_dff_B_m9jNYSza4_2),.clk(gclk));
	jdff dff_B_fYo9iQxr0_2(.din(w_dff_B_m9jNYSza4_2),.dout(w_dff_B_fYo9iQxr0_2),.clk(gclk));
	jdff dff_B_AJ278F735_2(.din(w_dff_B_fYo9iQxr0_2),.dout(w_dff_B_AJ278F735_2),.clk(gclk));
	jdff dff_B_6UGA7hQZ1_2(.din(n994),.dout(w_dff_B_6UGA7hQZ1_2),.clk(gclk));
	jdff dff_B_0oMYSq0L6_1(.din(n950),.dout(w_dff_B_0oMYSq0L6_1),.clk(gclk));
	jdff dff_B_loGNozgi9_2(.din(n847),.dout(w_dff_B_loGNozgi9_2),.clk(gclk));
	jdff dff_B_WwYCtl412_2(.din(w_dff_B_loGNozgi9_2),.dout(w_dff_B_WwYCtl412_2),.clk(gclk));
	jdff dff_B_0n1Jadz66_2(.din(w_dff_B_WwYCtl412_2),.dout(w_dff_B_0n1Jadz66_2),.clk(gclk));
	jdff dff_B_PVehoIcG1_2(.din(w_dff_B_0n1Jadz66_2),.dout(w_dff_B_PVehoIcG1_2),.clk(gclk));
	jdff dff_B_vgegI7jV3_2(.din(w_dff_B_PVehoIcG1_2),.dout(w_dff_B_vgegI7jV3_2),.clk(gclk));
	jdff dff_B_1Pkxkatc6_2(.din(w_dff_B_vgegI7jV3_2),.dout(w_dff_B_1Pkxkatc6_2),.clk(gclk));
	jdff dff_B_8YPRvzTG9_2(.din(w_dff_B_1Pkxkatc6_2),.dout(w_dff_B_8YPRvzTG9_2),.clk(gclk));
	jdff dff_B_5BL8usaY8_2(.din(w_dff_B_8YPRvzTG9_2),.dout(w_dff_B_5BL8usaY8_2),.clk(gclk));
	jdff dff_B_5Wt5ibDr7_2(.din(w_dff_B_5BL8usaY8_2),.dout(w_dff_B_5Wt5ibDr7_2),.clk(gclk));
	jdff dff_B_HGp057y16_2(.din(w_dff_B_5Wt5ibDr7_2),.dout(w_dff_B_HGp057y16_2),.clk(gclk));
	jdff dff_B_N3HA4PbK2_2(.din(w_dff_B_HGp057y16_2),.dout(w_dff_B_N3HA4PbK2_2),.clk(gclk));
	jdff dff_B_YP7WalGR7_2(.din(w_dff_B_N3HA4PbK2_2),.dout(w_dff_B_YP7WalGR7_2),.clk(gclk));
	jdff dff_B_xXCczbKI4_2(.din(w_dff_B_YP7WalGR7_2),.dout(w_dff_B_xXCczbKI4_2),.clk(gclk));
	jdff dff_B_GG2LoV179_2(.din(w_dff_B_xXCczbKI4_2),.dout(w_dff_B_GG2LoV179_2),.clk(gclk));
	jdff dff_B_7rTj1hxk0_2(.din(w_dff_B_GG2LoV179_2),.dout(w_dff_B_7rTj1hxk0_2),.clk(gclk));
	jdff dff_B_CU0GAnsS0_2(.din(w_dff_B_7rTj1hxk0_2),.dout(w_dff_B_CU0GAnsS0_2),.clk(gclk));
	jdff dff_B_lOPgQupd8_2(.din(w_dff_B_CU0GAnsS0_2),.dout(w_dff_B_lOPgQupd8_2),.clk(gclk));
	jdff dff_B_r7yNn4561_2(.din(w_dff_B_lOPgQupd8_2),.dout(w_dff_B_r7yNn4561_2),.clk(gclk));
	jdff dff_B_U5REUEV02_2(.din(w_dff_B_r7yNn4561_2),.dout(w_dff_B_U5REUEV02_2),.clk(gclk));
	jdff dff_B_nKiBMnI58_2(.din(w_dff_B_U5REUEV02_2),.dout(w_dff_B_nKiBMnI58_2),.clk(gclk));
	jdff dff_B_OuUO3ksH5_2(.din(n888),.dout(w_dff_B_OuUO3ksH5_2),.clk(gclk));
	jdff dff_B_ze7CwRxD5_1(.din(n848),.dout(w_dff_B_ze7CwRxD5_1),.clk(gclk));
	jdff dff_B_t2qiqlq82_2(.din(n749),.dout(w_dff_B_t2qiqlq82_2),.clk(gclk));
	jdff dff_B_hO8a1Kat6_2(.din(w_dff_B_t2qiqlq82_2),.dout(w_dff_B_hO8a1Kat6_2),.clk(gclk));
	jdff dff_B_vIvEHoZA5_2(.din(w_dff_B_hO8a1Kat6_2),.dout(w_dff_B_vIvEHoZA5_2),.clk(gclk));
	jdff dff_B_M4VIBpVI8_2(.din(w_dff_B_vIvEHoZA5_2),.dout(w_dff_B_M4VIBpVI8_2),.clk(gclk));
	jdff dff_B_rie1OaCW6_2(.din(w_dff_B_M4VIBpVI8_2),.dout(w_dff_B_rie1OaCW6_2),.clk(gclk));
	jdff dff_B_Q64ShAcO6_2(.din(w_dff_B_rie1OaCW6_2),.dout(w_dff_B_Q64ShAcO6_2),.clk(gclk));
	jdff dff_B_0aDQFoDM4_2(.din(w_dff_B_Q64ShAcO6_2),.dout(w_dff_B_0aDQFoDM4_2),.clk(gclk));
	jdff dff_B_LU8Dum5u8_2(.din(w_dff_B_0aDQFoDM4_2),.dout(w_dff_B_LU8Dum5u8_2),.clk(gclk));
	jdff dff_B_cM3drlQI4_2(.din(w_dff_B_LU8Dum5u8_2),.dout(w_dff_B_cM3drlQI4_2),.clk(gclk));
	jdff dff_B_Vl92Qsgo9_2(.din(w_dff_B_cM3drlQI4_2),.dout(w_dff_B_Vl92Qsgo9_2),.clk(gclk));
	jdff dff_B_uEBfFmQA5_2(.din(w_dff_B_Vl92Qsgo9_2),.dout(w_dff_B_uEBfFmQA5_2),.clk(gclk));
	jdff dff_B_1JArMmMc1_2(.din(w_dff_B_uEBfFmQA5_2),.dout(w_dff_B_1JArMmMc1_2),.clk(gclk));
	jdff dff_B_i5U1hvRO7_2(.din(w_dff_B_1JArMmMc1_2),.dout(w_dff_B_i5U1hvRO7_2),.clk(gclk));
	jdff dff_B_SGnsI4oE7_2(.din(w_dff_B_i5U1hvRO7_2),.dout(w_dff_B_SGnsI4oE7_2),.clk(gclk));
	jdff dff_B_zEE62LWO5_2(.din(w_dff_B_SGnsI4oE7_2),.dout(w_dff_B_zEE62LWO5_2),.clk(gclk));
	jdff dff_B_Y9rOaHPJ9_2(.din(w_dff_B_zEE62LWO5_2),.dout(w_dff_B_Y9rOaHPJ9_2),.clk(gclk));
	jdff dff_B_XlNQGqbr8_2(.din(w_dff_B_Y9rOaHPJ9_2),.dout(w_dff_B_XlNQGqbr8_2),.clk(gclk));
	jdff dff_B_5kYk2Ixa5_2(.din(n785),.dout(w_dff_B_5kYk2Ixa5_2),.clk(gclk));
	jdff dff_B_yZ1ZLZMX3_1(.din(n750),.dout(w_dff_B_yZ1ZLZMX3_1),.clk(gclk));
	jdff dff_B_9aoLueLy1_2(.din(n657),.dout(w_dff_B_9aoLueLy1_2),.clk(gclk));
	jdff dff_B_NKCKydGn2_2(.din(w_dff_B_9aoLueLy1_2),.dout(w_dff_B_NKCKydGn2_2),.clk(gclk));
	jdff dff_B_EnS2MZHq4_2(.din(w_dff_B_NKCKydGn2_2),.dout(w_dff_B_EnS2MZHq4_2),.clk(gclk));
	jdff dff_B_H4nkGOZq9_2(.din(w_dff_B_EnS2MZHq4_2),.dout(w_dff_B_H4nkGOZq9_2),.clk(gclk));
	jdff dff_B_I65d36uz4_2(.din(w_dff_B_H4nkGOZq9_2),.dout(w_dff_B_I65d36uz4_2),.clk(gclk));
	jdff dff_B_ODDEud1P6_2(.din(w_dff_B_I65d36uz4_2),.dout(w_dff_B_ODDEud1P6_2),.clk(gclk));
	jdff dff_B_YOraFkZV4_2(.din(w_dff_B_ODDEud1P6_2),.dout(w_dff_B_YOraFkZV4_2),.clk(gclk));
	jdff dff_B_Do3QMKhj3_2(.din(w_dff_B_YOraFkZV4_2),.dout(w_dff_B_Do3QMKhj3_2),.clk(gclk));
	jdff dff_B_5ngNZ9rE4_2(.din(w_dff_B_Do3QMKhj3_2),.dout(w_dff_B_5ngNZ9rE4_2),.clk(gclk));
	jdff dff_B_MMv7rcA25_2(.din(w_dff_B_5ngNZ9rE4_2),.dout(w_dff_B_MMv7rcA25_2),.clk(gclk));
	jdff dff_B_PfO4DHBQ4_2(.din(w_dff_B_MMv7rcA25_2),.dout(w_dff_B_PfO4DHBQ4_2),.clk(gclk));
	jdff dff_B_LksThUh49_2(.din(w_dff_B_PfO4DHBQ4_2),.dout(w_dff_B_LksThUh49_2),.clk(gclk));
	jdff dff_B_o4GO084i3_2(.din(w_dff_B_LksThUh49_2),.dout(w_dff_B_o4GO084i3_2),.clk(gclk));
	jdff dff_B_ZD8FogMh6_2(.din(w_dff_B_o4GO084i3_2),.dout(w_dff_B_ZD8FogMh6_2),.clk(gclk));
	jdff dff_B_YZpFnkvY4_2(.din(n686),.dout(w_dff_B_YZpFnkvY4_2),.clk(gclk));
	jdff dff_B_2TtZjgDR4_1(.din(n658),.dout(w_dff_B_2TtZjgDR4_1),.clk(gclk));
	jdff dff_B_Fjt8NB8M0_2(.din(n572),.dout(w_dff_B_Fjt8NB8M0_2),.clk(gclk));
	jdff dff_B_u3Ye1c305_2(.din(w_dff_B_Fjt8NB8M0_2),.dout(w_dff_B_u3Ye1c305_2),.clk(gclk));
	jdff dff_B_gUTxaUXY9_2(.din(w_dff_B_u3Ye1c305_2),.dout(w_dff_B_gUTxaUXY9_2),.clk(gclk));
	jdff dff_B_oevza0wB1_2(.din(w_dff_B_gUTxaUXY9_2),.dout(w_dff_B_oevza0wB1_2),.clk(gclk));
	jdff dff_B_a5k7dsn76_2(.din(w_dff_B_oevza0wB1_2),.dout(w_dff_B_a5k7dsn76_2),.clk(gclk));
	jdff dff_B_jd9iXizh0_2(.din(w_dff_B_a5k7dsn76_2),.dout(w_dff_B_jd9iXizh0_2),.clk(gclk));
	jdff dff_B_Gg90a2hp3_2(.din(w_dff_B_jd9iXizh0_2),.dout(w_dff_B_Gg90a2hp3_2),.clk(gclk));
	jdff dff_B_3CvsAI2d8_2(.din(w_dff_B_Gg90a2hp3_2),.dout(w_dff_B_3CvsAI2d8_2),.clk(gclk));
	jdff dff_B_yuFhykAK8_2(.din(w_dff_B_3CvsAI2d8_2),.dout(w_dff_B_yuFhykAK8_2),.clk(gclk));
	jdff dff_B_7cHnDViy2_2(.din(w_dff_B_yuFhykAK8_2),.dout(w_dff_B_7cHnDViy2_2),.clk(gclk));
	jdff dff_B_hpCVcopu1_2(.din(w_dff_B_7cHnDViy2_2),.dout(w_dff_B_hpCVcopu1_2),.clk(gclk));
	jdff dff_B_N8xVdQVc1_2(.din(n594),.dout(w_dff_B_N8xVdQVc1_2),.clk(gclk));
	jdff dff_B_xDE2wZ4o5_1(.din(n573),.dout(w_dff_B_xDE2wZ4o5_1),.clk(gclk));
	jdff dff_B_RVTKO89N5_2(.din(n494),.dout(w_dff_B_RVTKO89N5_2),.clk(gclk));
	jdff dff_B_A9ghjFdp7_2(.din(w_dff_B_RVTKO89N5_2),.dout(w_dff_B_A9ghjFdp7_2),.clk(gclk));
	jdff dff_B_WMQLPQZL3_2(.din(w_dff_B_A9ghjFdp7_2),.dout(w_dff_B_WMQLPQZL3_2),.clk(gclk));
	jdff dff_B_aFF7X2kQ6_2(.din(w_dff_B_WMQLPQZL3_2),.dout(w_dff_B_aFF7X2kQ6_2),.clk(gclk));
	jdff dff_B_XU1FHgmb0_2(.din(w_dff_B_aFF7X2kQ6_2),.dout(w_dff_B_XU1FHgmb0_2),.clk(gclk));
	jdff dff_B_DxLwwvlN7_2(.din(w_dff_B_XU1FHgmb0_2),.dout(w_dff_B_DxLwwvlN7_2),.clk(gclk));
	jdff dff_B_T9Gfyxhh1_2(.din(w_dff_B_DxLwwvlN7_2),.dout(w_dff_B_T9Gfyxhh1_2),.clk(gclk));
	jdff dff_B_enx57Ify0_2(.din(w_dff_B_T9Gfyxhh1_2),.dout(w_dff_B_enx57Ify0_2),.clk(gclk));
	jdff dff_B_NtmhkJ5H6_2(.din(n509),.dout(w_dff_B_NtmhkJ5H6_2),.clk(gclk));
	jdff dff_B_s5WQ3C6t1_2(.din(w_dff_B_NtmhkJ5H6_2),.dout(w_dff_B_s5WQ3C6t1_2),.clk(gclk));
	jdff dff_B_HmdH1K3B2_2(.din(w_dff_B_s5WQ3C6t1_2),.dout(w_dff_B_HmdH1K3B2_2),.clk(gclk));
	jdff dff_B_9yuZU2o59_1(.din(n495),.dout(w_dff_B_9yuZU2o59_1),.clk(gclk));
	jdff dff_B_UTv53eIV5_1(.din(w_dff_B_9yuZU2o59_1),.dout(w_dff_B_UTv53eIV5_1),.clk(gclk));
	jdff dff_B_tWtgbXPF4_2(.din(n425),.dout(w_dff_B_tWtgbXPF4_2),.clk(gclk));
	jdff dff_B_ac57eWrJ6_2(.din(w_dff_B_tWtgbXPF4_2),.dout(w_dff_B_ac57eWrJ6_2),.clk(gclk));
	jdff dff_B_qT2GWI6i5_2(.din(w_dff_B_ac57eWrJ6_2),.dout(w_dff_B_qT2GWI6i5_2),.clk(gclk));
	jdff dff_B_tFhInTpS8_0(.din(n430),.dout(w_dff_B_tFhInTpS8_0),.clk(gclk));
	jdff dff_A_Nr7FDlQy8_0(.dout(w_n358_0[0]),.din(w_dff_A_Nr7FDlQy8_0),.clk(gclk));
	jdff dff_A_ld5XHP2q6_0(.dout(w_dff_A_Nr7FDlQy8_0),.din(w_dff_A_ld5XHP2q6_0),.clk(gclk));
	jdff dff_A_eYh6xHTD4_1(.dout(w_n358_0[1]),.din(w_dff_A_eYh6xHTD4_1),.clk(gclk));
	jdff dff_A_iGOTVGdz2_1(.dout(w_dff_A_eYh6xHTD4_1),.din(w_dff_A_iGOTVGdz2_1),.clk(gclk));
	jdff dff_B_H4YrT5Qg7_2(.din(n1651),.dout(w_dff_B_H4YrT5Qg7_2),.clk(gclk));
	jdff dff_B_8u82OTEk1_1(.din(n1649),.dout(w_dff_B_8u82OTEk1_1),.clk(gclk));
	jdff dff_B_FGBf8jTf5_2(.din(n1597),.dout(w_dff_B_FGBf8jTf5_2),.clk(gclk));
	jdff dff_B_U6B4oF6j0_2(.din(w_dff_B_FGBf8jTf5_2),.dout(w_dff_B_U6B4oF6j0_2),.clk(gclk));
	jdff dff_B_3fEIf1bE7_2(.din(w_dff_B_U6B4oF6j0_2),.dout(w_dff_B_3fEIf1bE7_2),.clk(gclk));
	jdff dff_B_yMlOjoPT8_2(.din(w_dff_B_3fEIf1bE7_2),.dout(w_dff_B_yMlOjoPT8_2),.clk(gclk));
	jdff dff_B_kCyg5rZc0_2(.din(w_dff_B_yMlOjoPT8_2),.dout(w_dff_B_kCyg5rZc0_2),.clk(gclk));
	jdff dff_B_ss9DrP9Y1_2(.din(w_dff_B_kCyg5rZc0_2),.dout(w_dff_B_ss9DrP9Y1_2),.clk(gclk));
	jdff dff_B_dvk5yyze7_2(.din(w_dff_B_ss9DrP9Y1_2),.dout(w_dff_B_dvk5yyze7_2),.clk(gclk));
	jdff dff_B_4ywqs0yT2_2(.din(w_dff_B_dvk5yyze7_2),.dout(w_dff_B_4ywqs0yT2_2),.clk(gclk));
	jdff dff_B_Gh7a08yD4_2(.din(w_dff_B_4ywqs0yT2_2),.dout(w_dff_B_Gh7a08yD4_2),.clk(gclk));
	jdff dff_B_JdaNaoCJ2_2(.din(w_dff_B_Gh7a08yD4_2),.dout(w_dff_B_JdaNaoCJ2_2),.clk(gclk));
	jdff dff_B_pectrKqf5_2(.din(w_dff_B_JdaNaoCJ2_2),.dout(w_dff_B_pectrKqf5_2),.clk(gclk));
	jdff dff_B_3R9HEZGO0_2(.din(w_dff_B_pectrKqf5_2),.dout(w_dff_B_3R9HEZGO0_2),.clk(gclk));
	jdff dff_B_9ygUsPbc1_2(.din(w_dff_B_3R9HEZGO0_2),.dout(w_dff_B_9ygUsPbc1_2),.clk(gclk));
	jdff dff_B_bOpPDq8M7_2(.din(w_dff_B_9ygUsPbc1_2),.dout(w_dff_B_bOpPDq8M7_2),.clk(gclk));
	jdff dff_B_Yj0muCWl6_2(.din(w_dff_B_bOpPDq8M7_2),.dout(w_dff_B_Yj0muCWl6_2),.clk(gclk));
	jdff dff_B_se3wxhWY6_2(.din(w_dff_B_Yj0muCWl6_2),.dout(w_dff_B_se3wxhWY6_2),.clk(gclk));
	jdff dff_B_F3XBj8p07_2(.din(w_dff_B_se3wxhWY6_2),.dout(w_dff_B_F3XBj8p07_2),.clk(gclk));
	jdff dff_B_VVdkneR19_2(.din(w_dff_B_F3XBj8p07_2),.dout(w_dff_B_VVdkneR19_2),.clk(gclk));
	jdff dff_B_LpBLNGRS6_2(.din(w_dff_B_VVdkneR19_2),.dout(w_dff_B_LpBLNGRS6_2),.clk(gclk));
	jdff dff_B_2VuZlde11_2(.din(w_dff_B_LpBLNGRS6_2),.dout(w_dff_B_2VuZlde11_2),.clk(gclk));
	jdff dff_B_nFCJ8jKP4_2(.din(w_dff_B_2VuZlde11_2),.dout(w_dff_B_nFCJ8jKP4_2),.clk(gclk));
	jdff dff_B_KJT6IcWt6_2(.din(w_dff_B_nFCJ8jKP4_2),.dout(w_dff_B_KJT6IcWt6_2),.clk(gclk));
	jdff dff_B_yRnuStW29_2(.din(w_dff_B_KJT6IcWt6_2),.dout(w_dff_B_yRnuStW29_2),.clk(gclk));
	jdff dff_B_f7ZKQCdD4_2(.din(w_dff_B_yRnuStW29_2),.dout(w_dff_B_f7ZKQCdD4_2),.clk(gclk));
	jdff dff_B_cXNZhmIG1_2(.din(w_dff_B_f7ZKQCdD4_2),.dout(w_dff_B_cXNZhmIG1_2),.clk(gclk));
	jdff dff_B_crvvGL4B9_2(.din(w_dff_B_cXNZhmIG1_2),.dout(w_dff_B_crvvGL4B9_2),.clk(gclk));
	jdff dff_B_UhOpIEwD0_2(.din(w_dff_B_crvvGL4B9_2),.dout(w_dff_B_UhOpIEwD0_2),.clk(gclk));
	jdff dff_B_ORNnKSAZ3_2(.din(w_dff_B_UhOpIEwD0_2),.dout(w_dff_B_ORNnKSAZ3_2),.clk(gclk));
	jdff dff_B_O8kLOrDs2_2(.din(w_dff_B_ORNnKSAZ3_2),.dout(w_dff_B_O8kLOrDs2_2),.clk(gclk));
	jdff dff_B_uDZeASMP8_2(.din(w_dff_B_O8kLOrDs2_2),.dout(w_dff_B_uDZeASMP8_2),.clk(gclk));
	jdff dff_B_7PCcJPzQ8_2(.din(w_dff_B_uDZeASMP8_2),.dout(w_dff_B_7PCcJPzQ8_2),.clk(gclk));
	jdff dff_B_Wr61stAb9_2(.din(w_dff_B_7PCcJPzQ8_2),.dout(w_dff_B_Wr61stAb9_2),.clk(gclk));
	jdff dff_B_QiQR7aMu3_2(.din(w_dff_B_Wr61stAb9_2),.dout(w_dff_B_QiQR7aMu3_2),.clk(gclk));
	jdff dff_B_i18PVtYj0_2(.din(w_dff_B_QiQR7aMu3_2),.dout(w_dff_B_i18PVtYj0_2),.clk(gclk));
	jdff dff_B_CaZbuqti0_2(.din(w_dff_B_i18PVtYj0_2),.dout(w_dff_B_CaZbuqti0_2),.clk(gclk));
	jdff dff_B_KjIXxOAI4_2(.din(w_dff_B_CaZbuqti0_2),.dout(w_dff_B_KjIXxOAI4_2),.clk(gclk));
	jdff dff_B_yNlJaCvY2_2(.din(w_dff_B_KjIXxOAI4_2),.dout(w_dff_B_yNlJaCvY2_2),.clk(gclk));
	jdff dff_B_0vT1vTWF3_2(.din(w_dff_B_yNlJaCvY2_2),.dout(w_dff_B_0vT1vTWF3_2),.clk(gclk));
	jdff dff_B_txootfBz2_2(.din(w_dff_B_0vT1vTWF3_2),.dout(w_dff_B_txootfBz2_2),.clk(gclk));
	jdff dff_B_kNuXWdfu9_2(.din(w_dff_B_txootfBz2_2),.dout(w_dff_B_kNuXWdfu9_2),.clk(gclk));
	jdff dff_B_detvEDeQ7_2(.din(w_dff_B_kNuXWdfu9_2),.dout(w_dff_B_detvEDeQ7_2),.clk(gclk));
	jdff dff_B_sWByKdUo7_2(.din(w_dff_B_detvEDeQ7_2),.dout(w_dff_B_sWByKdUo7_2),.clk(gclk));
	jdff dff_B_2AclVfkZ8_2(.din(w_dff_B_sWByKdUo7_2),.dout(w_dff_B_2AclVfkZ8_2),.clk(gclk));
	jdff dff_B_q3Jkis7o0_2(.din(w_dff_B_2AclVfkZ8_2),.dout(w_dff_B_q3Jkis7o0_2),.clk(gclk));
	jdff dff_B_Atz20Po82_2(.din(w_dff_B_q3Jkis7o0_2),.dout(w_dff_B_Atz20Po82_2),.clk(gclk));
	jdff dff_B_r2TRi9Mw7_2(.din(w_dff_B_Atz20Po82_2),.dout(w_dff_B_r2TRi9Mw7_2),.clk(gclk));
	jdff dff_B_5fqpPpqw5_1(.din(n1598),.dout(w_dff_B_5fqpPpqw5_1),.clk(gclk));
	jdff dff_B_QrfLMSFN7_2(.din(n1540),.dout(w_dff_B_QrfLMSFN7_2),.clk(gclk));
	jdff dff_B_SwO2J2EG7_2(.din(w_dff_B_QrfLMSFN7_2),.dout(w_dff_B_SwO2J2EG7_2),.clk(gclk));
	jdff dff_B_Dhp19eWZ8_2(.din(w_dff_B_SwO2J2EG7_2),.dout(w_dff_B_Dhp19eWZ8_2),.clk(gclk));
	jdff dff_B_oEFFDRTh8_2(.din(w_dff_B_Dhp19eWZ8_2),.dout(w_dff_B_oEFFDRTh8_2),.clk(gclk));
	jdff dff_B_n4yAV2wC8_2(.din(w_dff_B_oEFFDRTh8_2),.dout(w_dff_B_n4yAV2wC8_2),.clk(gclk));
	jdff dff_B_3SGtO3pG8_2(.din(w_dff_B_n4yAV2wC8_2),.dout(w_dff_B_3SGtO3pG8_2),.clk(gclk));
	jdff dff_B_WPmYJb8g0_2(.din(w_dff_B_3SGtO3pG8_2),.dout(w_dff_B_WPmYJb8g0_2),.clk(gclk));
	jdff dff_B_vamdq46V0_2(.din(w_dff_B_WPmYJb8g0_2),.dout(w_dff_B_vamdq46V0_2),.clk(gclk));
	jdff dff_B_2c0lb1Bf7_2(.din(w_dff_B_vamdq46V0_2),.dout(w_dff_B_2c0lb1Bf7_2),.clk(gclk));
	jdff dff_B_Sm94U7RC0_2(.din(w_dff_B_2c0lb1Bf7_2),.dout(w_dff_B_Sm94U7RC0_2),.clk(gclk));
	jdff dff_B_tovPr3Gj6_2(.din(w_dff_B_Sm94U7RC0_2),.dout(w_dff_B_tovPr3Gj6_2),.clk(gclk));
	jdff dff_B_zPC9L6st9_2(.din(w_dff_B_tovPr3Gj6_2),.dout(w_dff_B_zPC9L6st9_2),.clk(gclk));
	jdff dff_B_sTXdIzQA2_2(.din(w_dff_B_zPC9L6st9_2),.dout(w_dff_B_sTXdIzQA2_2),.clk(gclk));
	jdff dff_B_x1NngZmO0_2(.din(w_dff_B_sTXdIzQA2_2),.dout(w_dff_B_x1NngZmO0_2),.clk(gclk));
	jdff dff_B_azJUgKoO7_2(.din(w_dff_B_x1NngZmO0_2),.dout(w_dff_B_azJUgKoO7_2),.clk(gclk));
	jdff dff_B_u3P2LWv37_2(.din(w_dff_B_azJUgKoO7_2),.dout(w_dff_B_u3P2LWv37_2),.clk(gclk));
	jdff dff_B_cdPaMq575_2(.din(w_dff_B_u3P2LWv37_2),.dout(w_dff_B_cdPaMq575_2),.clk(gclk));
	jdff dff_B_Zq5If9UR2_2(.din(w_dff_B_cdPaMq575_2),.dout(w_dff_B_Zq5If9UR2_2),.clk(gclk));
	jdff dff_B_w6kQEEtk9_2(.din(w_dff_B_Zq5If9UR2_2),.dout(w_dff_B_w6kQEEtk9_2),.clk(gclk));
	jdff dff_B_fbeGPNnm0_2(.din(w_dff_B_w6kQEEtk9_2),.dout(w_dff_B_fbeGPNnm0_2),.clk(gclk));
	jdff dff_B_BkEWtN9y7_2(.din(w_dff_B_fbeGPNnm0_2),.dout(w_dff_B_BkEWtN9y7_2),.clk(gclk));
	jdff dff_B_lvhUxNJ98_2(.din(w_dff_B_BkEWtN9y7_2),.dout(w_dff_B_lvhUxNJ98_2),.clk(gclk));
	jdff dff_B_ecqrKTUu2_2(.din(w_dff_B_lvhUxNJ98_2),.dout(w_dff_B_ecqrKTUu2_2),.clk(gclk));
	jdff dff_B_Y5dEumy19_2(.din(w_dff_B_ecqrKTUu2_2),.dout(w_dff_B_Y5dEumy19_2),.clk(gclk));
	jdff dff_B_s2o6rmh26_2(.din(w_dff_B_Y5dEumy19_2),.dout(w_dff_B_s2o6rmh26_2),.clk(gclk));
	jdff dff_B_NMEG0RSD1_2(.din(w_dff_B_s2o6rmh26_2),.dout(w_dff_B_NMEG0RSD1_2),.clk(gclk));
	jdff dff_B_JC3shGiu0_2(.din(w_dff_B_NMEG0RSD1_2),.dout(w_dff_B_JC3shGiu0_2),.clk(gclk));
	jdff dff_B_pXr7CSBT4_2(.din(w_dff_B_JC3shGiu0_2),.dout(w_dff_B_pXr7CSBT4_2),.clk(gclk));
	jdff dff_B_8w5qjcmb8_2(.din(w_dff_B_pXr7CSBT4_2),.dout(w_dff_B_8w5qjcmb8_2),.clk(gclk));
	jdff dff_B_z0CxYak16_2(.din(w_dff_B_8w5qjcmb8_2),.dout(w_dff_B_z0CxYak16_2),.clk(gclk));
	jdff dff_B_n8slCP0C6_2(.din(w_dff_B_z0CxYak16_2),.dout(w_dff_B_n8slCP0C6_2),.clk(gclk));
	jdff dff_B_VT0uZWCC8_2(.din(w_dff_B_n8slCP0C6_2),.dout(w_dff_B_VT0uZWCC8_2),.clk(gclk));
	jdff dff_B_bADfbBni1_2(.din(w_dff_B_VT0uZWCC8_2),.dout(w_dff_B_bADfbBni1_2),.clk(gclk));
	jdff dff_B_4BIGkTLY9_2(.din(w_dff_B_bADfbBni1_2),.dout(w_dff_B_4BIGkTLY9_2),.clk(gclk));
	jdff dff_B_4emyKrqa6_2(.din(w_dff_B_4BIGkTLY9_2),.dout(w_dff_B_4emyKrqa6_2),.clk(gclk));
	jdff dff_B_m5RFnYi50_2(.din(w_dff_B_4emyKrqa6_2),.dout(w_dff_B_m5RFnYi50_2),.clk(gclk));
	jdff dff_B_HUgFLPur3_2(.din(w_dff_B_m5RFnYi50_2),.dout(w_dff_B_HUgFLPur3_2),.clk(gclk));
	jdff dff_B_a4usGJD99_2(.din(w_dff_B_HUgFLPur3_2),.dout(w_dff_B_a4usGJD99_2),.clk(gclk));
	jdff dff_B_74qhYA3S4_2(.din(w_dff_B_a4usGJD99_2),.dout(w_dff_B_74qhYA3S4_2),.clk(gclk));
	jdff dff_B_K35Yb9Sz9_2(.din(w_dff_B_74qhYA3S4_2),.dout(w_dff_B_K35Yb9Sz9_2),.clk(gclk));
	jdff dff_B_KK9cnNdY5_2(.din(w_dff_B_K35Yb9Sz9_2),.dout(w_dff_B_KK9cnNdY5_2),.clk(gclk));
	jdff dff_B_qGDh7Zs29_2(.din(n1579),.dout(w_dff_B_qGDh7Zs29_2),.clk(gclk));
	jdff dff_B_nhG2MuVO0_1(.din(n1541),.dout(w_dff_B_nhG2MuVO0_1),.clk(gclk));
	jdff dff_B_a1J0J8zG7_2(.din(n1476),.dout(w_dff_B_a1J0J8zG7_2),.clk(gclk));
	jdff dff_B_sLsiD19P3_2(.din(w_dff_B_a1J0J8zG7_2),.dout(w_dff_B_sLsiD19P3_2),.clk(gclk));
	jdff dff_B_kZurIMWo1_2(.din(w_dff_B_sLsiD19P3_2),.dout(w_dff_B_kZurIMWo1_2),.clk(gclk));
	jdff dff_B_v1clK4ii3_2(.din(w_dff_B_kZurIMWo1_2),.dout(w_dff_B_v1clK4ii3_2),.clk(gclk));
	jdff dff_B_kbrYLWt37_2(.din(w_dff_B_v1clK4ii3_2),.dout(w_dff_B_kbrYLWt37_2),.clk(gclk));
	jdff dff_B_C1Pb4Yuh2_2(.din(w_dff_B_kbrYLWt37_2),.dout(w_dff_B_C1Pb4Yuh2_2),.clk(gclk));
	jdff dff_B_Dut4g0gZ1_2(.din(w_dff_B_C1Pb4Yuh2_2),.dout(w_dff_B_Dut4g0gZ1_2),.clk(gclk));
	jdff dff_B_MpKWRWAR2_2(.din(w_dff_B_Dut4g0gZ1_2),.dout(w_dff_B_MpKWRWAR2_2),.clk(gclk));
	jdff dff_B_Fql4Qd7Y3_2(.din(w_dff_B_MpKWRWAR2_2),.dout(w_dff_B_Fql4Qd7Y3_2),.clk(gclk));
	jdff dff_B_HHxpagHl6_2(.din(w_dff_B_Fql4Qd7Y3_2),.dout(w_dff_B_HHxpagHl6_2),.clk(gclk));
	jdff dff_B_PZ1KQNwm2_2(.din(w_dff_B_HHxpagHl6_2),.dout(w_dff_B_PZ1KQNwm2_2),.clk(gclk));
	jdff dff_B_nKl0y47p4_2(.din(w_dff_B_PZ1KQNwm2_2),.dout(w_dff_B_nKl0y47p4_2),.clk(gclk));
	jdff dff_B_OYBpVMMG4_2(.din(w_dff_B_nKl0y47p4_2),.dout(w_dff_B_OYBpVMMG4_2),.clk(gclk));
	jdff dff_B_DhW66jAU8_2(.din(w_dff_B_OYBpVMMG4_2),.dout(w_dff_B_DhW66jAU8_2),.clk(gclk));
	jdff dff_B_PKuxjvw20_2(.din(w_dff_B_DhW66jAU8_2),.dout(w_dff_B_PKuxjvw20_2),.clk(gclk));
	jdff dff_B_XO8h7PGg5_2(.din(w_dff_B_PKuxjvw20_2),.dout(w_dff_B_XO8h7PGg5_2),.clk(gclk));
	jdff dff_B_6upL2GWj7_2(.din(w_dff_B_XO8h7PGg5_2),.dout(w_dff_B_6upL2GWj7_2),.clk(gclk));
	jdff dff_B_GFhoQmhn0_2(.din(w_dff_B_6upL2GWj7_2),.dout(w_dff_B_GFhoQmhn0_2),.clk(gclk));
	jdff dff_B_SY94yo6c3_2(.din(w_dff_B_GFhoQmhn0_2),.dout(w_dff_B_SY94yo6c3_2),.clk(gclk));
	jdff dff_B_usDLdEv52_2(.din(w_dff_B_SY94yo6c3_2),.dout(w_dff_B_usDLdEv52_2),.clk(gclk));
	jdff dff_B_sQZJRW9M8_2(.din(w_dff_B_usDLdEv52_2),.dout(w_dff_B_sQZJRW9M8_2),.clk(gclk));
	jdff dff_B_RS1zbws18_2(.din(w_dff_B_sQZJRW9M8_2),.dout(w_dff_B_RS1zbws18_2),.clk(gclk));
	jdff dff_B_oizmTqgH0_2(.din(w_dff_B_RS1zbws18_2),.dout(w_dff_B_oizmTqgH0_2),.clk(gclk));
	jdff dff_B_7PiZW7l29_2(.din(w_dff_B_oizmTqgH0_2),.dout(w_dff_B_7PiZW7l29_2),.clk(gclk));
	jdff dff_B_A6TJtnUN1_2(.din(w_dff_B_7PiZW7l29_2),.dout(w_dff_B_A6TJtnUN1_2),.clk(gclk));
	jdff dff_B_ohZEdczW6_2(.din(w_dff_B_A6TJtnUN1_2),.dout(w_dff_B_ohZEdczW6_2),.clk(gclk));
	jdff dff_B_qy9MKSzC9_2(.din(w_dff_B_ohZEdczW6_2),.dout(w_dff_B_qy9MKSzC9_2),.clk(gclk));
	jdff dff_B_iIQ3jMah6_2(.din(w_dff_B_qy9MKSzC9_2),.dout(w_dff_B_iIQ3jMah6_2),.clk(gclk));
	jdff dff_B_R38DuS625_2(.din(w_dff_B_iIQ3jMah6_2),.dout(w_dff_B_R38DuS625_2),.clk(gclk));
	jdff dff_B_vIsaCBPL2_2(.din(w_dff_B_R38DuS625_2),.dout(w_dff_B_vIsaCBPL2_2),.clk(gclk));
	jdff dff_B_cUbWS54X7_2(.din(w_dff_B_vIsaCBPL2_2),.dout(w_dff_B_cUbWS54X7_2),.clk(gclk));
	jdff dff_B_eOyqHQmx1_2(.din(w_dff_B_cUbWS54X7_2),.dout(w_dff_B_eOyqHQmx1_2),.clk(gclk));
	jdff dff_B_i0NGRoIy4_2(.din(w_dff_B_eOyqHQmx1_2),.dout(w_dff_B_i0NGRoIy4_2),.clk(gclk));
	jdff dff_B_QUAW3t0y8_2(.din(w_dff_B_i0NGRoIy4_2),.dout(w_dff_B_QUAW3t0y8_2),.clk(gclk));
	jdff dff_B_fLeIxoKr1_2(.din(w_dff_B_QUAW3t0y8_2),.dout(w_dff_B_fLeIxoKr1_2),.clk(gclk));
	jdff dff_B_hKsMYOUV6_2(.din(w_dff_B_fLeIxoKr1_2),.dout(w_dff_B_hKsMYOUV6_2),.clk(gclk));
	jdff dff_B_9uGbm21M2_2(.din(w_dff_B_hKsMYOUV6_2),.dout(w_dff_B_9uGbm21M2_2),.clk(gclk));
	jdff dff_B_azQbmOOL5_2(.din(w_dff_B_9uGbm21M2_2),.dout(w_dff_B_azQbmOOL5_2),.clk(gclk));
	jdff dff_B_BHERS2qa9_2(.din(n1515),.dout(w_dff_B_BHERS2qa9_2),.clk(gclk));
	jdff dff_B_zf6t6t9G7_1(.din(n1477),.dout(w_dff_B_zf6t6t9G7_1),.clk(gclk));
	jdff dff_B_dHAvEPUM8_2(.din(n1405),.dout(w_dff_B_dHAvEPUM8_2),.clk(gclk));
	jdff dff_B_9vA585IV4_2(.din(w_dff_B_dHAvEPUM8_2),.dout(w_dff_B_9vA585IV4_2),.clk(gclk));
	jdff dff_B_5Ot79jrZ1_2(.din(w_dff_B_9vA585IV4_2),.dout(w_dff_B_5Ot79jrZ1_2),.clk(gclk));
	jdff dff_B_bQt6pq1O5_2(.din(w_dff_B_5Ot79jrZ1_2),.dout(w_dff_B_bQt6pq1O5_2),.clk(gclk));
	jdff dff_B_aCRvs3vO8_2(.din(w_dff_B_bQt6pq1O5_2),.dout(w_dff_B_aCRvs3vO8_2),.clk(gclk));
	jdff dff_B_OuMRJDx00_2(.din(w_dff_B_aCRvs3vO8_2),.dout(w_dff_B_OuMRJDx00_2),.clk(gclk));
	jdff dff_B_7rnNunb37_2(.din(w_dff_B_OuMRJDx00_2),.dout(w_dff_B_7rnNunb37_2),.clk(gclk));
	jdff dff_B_UNyA0LNQ6_2(.din(w_dff_B_7rnNunb37_2),.dout(w_dff_B_UNyA0LNQ6_2),.clk(gclk));
	jdff dff_B_NkuPCib06_2(.din(w_dff_B_UNyA0LNQ6_2),.dout(w_dff_B_NkuPCib06_2),.clk(gclk));
	jdff dff_B_HrWAqTVg2_2(.din(w_dff_B_NkuPCib06_2),.dout(w_dff_B_HrWAqTVg2_2),.clk(gclk));
	jdff dff_B_jr0H6M1h2_2(.din(w_dff_B_HrWAqTVg2_2),.dout(w_dff_B_jr0H6M1h2_2),.clk(gclk));
	jdff dff_B_SWrWulLa4_2(.din(w_dff_B_jr0H6M1h2_2),.dout(w_dff_B_SWrWulLa4_2),.clk(gclk));
	jdff dff_B_Jct4dJkK5_2(.din(w_dff_B_SWrWulLa4_2),.dout(w_dff_B_Jct4dJkK5_2),.clk(gclk));
	jdff dff_B_gvxPh2zu3_2(.din(w_dff_B_Jct4dJkK5_2),.dout(w_dff_B_gvxPh2zu3_2),.clk(gclk));
	jdff dff_B_irv6qS638_2(.din(w_dff_B_gvxPh2zu3_2),.dout(w_dff_B_irv6qS638_2),.clk(gclk));
	jdff dff_B_77RqiY8q1_2(.din(w_dff_B_irv6qS638_2),.dout(w_dff_B_77RqiY8q1_2),.clk(gclk));
	jdff dff_B_4vLrbhgG4_2(.din(w_dff_B_77RqiY8q1_2),.dout(w_dff_B_4vLrbhgG4_2),.clk(gclk));
	jdff dff_B_oshIgT4C9_2(.din(w_dff_B_4vLrbhgG4_2),.dout(w_dff_B_oshIgT4C9_2),.clk(gclk));
	jdff dff_B_m3SBlrPt7_2(.din(w_dff_B_oshIgT4C9_2),.dout(w_dff_B_m3SBlrPt7_2),.clk(gclk));
	jdff dff_B_tfumFg1C3_2(.din(w_dff_B_m3SBlrPt7_2),.dout(w_dff_B_tfumFg1C3_2),.clk(gclk));
	jdff dff_B_wLCrObGZ6_2(.din(w_dff_B_tfumFg1C3_2),.dout(w_dff_B_wLCrObGZ6_2),.clk(gclk));
	jdff dff_B_VVLKQ5Q39_2(.din(w_dff_B_wLCrObGZ6_2),.dout(w_dff_B_VVLKQ5Q39_2),.clk(gclk));
	jdff dff_B_ezfXU9GF3_2(.din(w_dff_B_VVLKQ5Q39_2),.dout(w_dff_B_ezfXU9GF3_2),.clk(gclk));
	jdff dff_B_cdb9Mvoj9_2(.din(w_dff_B_ezfXU9GF3_2),.dout(w_dff_B_cdb9Mvoj9_2),.clk(gclk));
	jdff dff_B_lLLZcuUT7_2(.din(w_dff_B_cdb9Mvoj9_2),.dout(w_dff_B_lLLZcuUT7_2),.clk(gclk));
	jdff dff_B_6O5EvuP08_2(.din(w_dff_B_lLLZcuUT7_2),.dout(w_dff_B_6O5EvuP08_2),.clk(gclk));
	jdff dff_B_Ooj3M8kE1_2(.din(w_dff_B_6O5EvuP08_2),.dout(w_dff_B_Ooj3M8kE1_2),.clk(gclk));
	jdff dff_B_MKSnQWk41_2(.din(w_dff_B_Ooj3M8kE1_2),.dout(w_dff_B_MKSnQWk41_2),.clk(gclk));
	jdff dff_B_oLOudchR1_2(.din(w_dff_B_MKSnQWk41_2),.dout(w_dff_B_oLOudchR1_2),.clk(gclk));
	jdff dff_B_zLTCYzRl5_2(.din(w_dff_B_oLOudchR1_2),.dout(w_dff_B_zLTCYzRl5_2),.clk(gclk));
	jdff dff_B_16exLBNQ7_2(.din(w_dff_B_zLTCYzRl5_2),.dout(w_dff_B_16exLBNQ7_2),.clk(gclk));
	jdff dff_B_EdcHSJMl5_2(.din(w_dff_B_16exLBNQ7_2),.dout(w_dff_B_EdcHSJMl5_2),.clk(gclk));
	jdff dff_B_shG9GEvp3_2(.din(w_dff_B_EdcHSJMl5_2),.dout(w_dff_B_shG9GEvp3_2),.clk(gclk));
	jdff dff_B_27VPICdG5_2(.din(w_dff_B_shG9GEvp3_2),.dout(w_dff_B_27VPICdG5_2),.clk(gclk));
	jdff dff_B_S6AkPJPj3_2(.din(w_dff_B_27VPICdG5_2),.dout(w_dff_B_S6AkPJPj3_2),.clk(gclk));
	jdff dff_B_YJTAuJ945_2(.din(n1444),.dout(w_dff_B_YJTAuJ945_2),.clk(gclk));
	jdff dff_B_vokYGC0b9_1(.din(n1406),.dout(w_dff_B_vokYGC0b9_1),.clk(gclk));
	jdff dff_B_Rs2hwzpB6_2(.din(n1327),.dout(w_dff_B_Rs2hwzpB6_2),.clk(gclk));
	jdff dff_B_aasmsvVd2_2(.din(w_dff_B_Rs2hwzpB6_2),.dout(w_dff_B_aasmsvVd2_2),.clk(gclk));
	jdff dff_B_4LFEAv2j1_2(.din(w_dff_B_aasmsvVd2_2),.dout(w_dff_B_4LFEAv2j1_2),.clk(gclk));
	jdff dff_B_eaDDy6O16_2(.din(w_dff_B_4LFEAv2j1_2),.dout(w_dff_B_eaDDy6O16_2),.clk(gclk));
	jdff dff_B_OcaGUfCW3_2(.din(w_dff_B_eaDDy6O16_2),.dout(w_dff_B_OcaGUfCW3_2),.clk(gclk));
	jdff dff_B_PNv8s8b13_2(.din(w_dff_B_OcaGUfCW3_2),.dout(w_dff_B_PNv8s8b13_2),.clk(gclk));
	jdff dff_B_vBZLomtJ0_2(.din(w_dff_B_PNv8s8b13_2),.dout(w_dff_B_vBZLomtJ0_2),.clk(gclk));
	jdff dff_B_pFNvnAe62_2(.din(w_dff_B_vBZLomtJ0_2),.dout(w_dff_B_pFNvnAe62_2),.clk(gclk));
	jdff dff_B_JH47gPyU9_2(.din(w_dff_B_pFNvnAe62_2),.dout(w_dff_B_JH47gPyU9_2),.clk(gclk));
	jdff dff_B_rV3xResR9_2(.din(w_dff_B_JH47gPyU9_2),.dout(w_dff_B_rV3xResR9_2),.clk(gclk));
	jdff dff_B_63Ip9KMa2_2(.din(w_dff_B_rV3xResR9_2),.dout(w_dff_B_63Ip9KMa2_2),.clk(gclk));
	jdff dff_B_6M2EC8Sh4_2(.din(w_dff_B_63Ip9KMa2_2),.dout(w_dff_B_6M2EC8Sh4_2),.clk(gclk));
	jdff dff_B_bcnpDTA37_2(.din(w_dff_B_6M2EC8Sh4_2),.dout(w_dff_B_bcnpDTA37_2),.clk(gclk));
	jdff dff_B_CZEdGSg04_2(.din(w_dff_B_bcnpDTA37_2),.dout(w_dff_B_CZEdGSg04_2),.clk(gclk));
	jdff dff_B_mm5R5TOt7_2(.din(w_dff_B_CZEdGSg04_2),.dout(w_dff_B_mm5R5TOt7_2),.clk(gclk));
	jdff dff_B_60Pm7ex72_2(.din(w_dff_B_mm5R5TOt7_2),.dout(w_dff_B_60Pm7ex72_2),.clk(gclk));
	jdff dff_B_PblsyD8d8_2(.din(w_dff_B_60Pm7ex72_2),.dout(w_dff_B_PblsyD8d8_2),.clk(gclk));
	jdff dff_B_RwT1Wr1B0_2(.din(w_dff_B_PblsyD8d8_2),.dout(w_dff_B_RwT1Wr1B0_2),.clk(gclk));
	jdff dff_B_vzNWISLk7_2(.din(w_dff_B_RwT1Wr1B0_2),.dout(w_dff_B_vzNWISLk7_2),.clk(gclk));
	jdff dff_B_3Kovejb60_2(.din(w_dff_B_vzNWISLk7_2),.dout(w_dff_B_3Kovejb60_2),.clk(gclk));
	jdff dff_B_fYZ8xuDg6_2(.din(w_dff_B_3Kovejb60_2),.dout(w_dff_B_fYZ8xuDg6_2),.clk(gclk));
	jdff dff_B_chM9taEi2_2(.din(w_dff_B_fYZ8xuDg6_2),.dout(w_dff_B_chM9taEi2_2),.clk(gclk));
	jdff dff_B_74WmtdW34_2(.din(w_dff_B_chM9taEi2_2),.dout(w_dff_B_74WmtdW34_2),.clk(gclk));
	jdff dff_B_j07Wur1H8_2(.din(w_dff_B_74WmtdW34_2),.dout(w_dff_B_j07Wur1H8_2),.clk(gclk));
	jdff dff_B_oqLzKfjo0_2(.din(w_dff_B_j07Wur1H8_2),.dout(w_dff_B_oqLzKfjo0_2),.clk(gclk));
	jdff dff_B_AcLahKgS3_2(.din(w_dff_B_oqLzKfjo0_2),.dout(w_dff_B_AcLahKgS3_2),.clk(gclk));
	jdff dff_B_t5uMJZv03_2(.din(w_dff_B_AcLahKgS3_2),.dout(w_dff_B_t5uMJZv03_2),.clk(gclk));
	jdff dff_B_3hXUBDKd9_2(.din(w_dff_B_t5uMJZv03_2),.dout(w_dff_B_3hXUBDKd9_2),.clk(gclk));
	jdff dff_B_V6ganN2S2_2(.din(w_dff_B_3hXUBDKd9_2),.dout(w_dff_B_V6ganN2S2_2),.clk(gclk));
	jdff dff_B_ZnWklMm30_2(.din(w_dff_B_V6ganN2S2_2),.dout(w_dff_B_ZnWklMm30_2),.clk(gclk));
	jdff dff_B_HPrd3aYp5_2(.din(w_dff_B_ZnWklMm30_2),.dout(w_dff_B_HPrd3aYp5_2),.clk(gclk));
	jdff dff_B_FQxKZDL89_2(.din(w_dff_B_HPrd3aYp5_2),.dout(w_dff_B_FQxKZDL89_2),.clk(gclk));
	jdff dff_B_Iax4cSnN7_2(.din(n1366),.dout(w_dff_B_Iax4cSnN7_2),.clk(gclk));
	jdff dff_B_UmQpK0rO6_1(.din(n1328),.dout(w_dff_B_UmQpK0rO6_1),.clk(gclk));
	jdff dff_B_FsbPAJqs4_2(.din(n1242),.dout(w_dff_B_FsbPAJqs4_2),.clk(gclk));
	jdff dff_B_hr2bwteo6_2(.din(w_dff_B_FsbPAJqs4_2),.dout(w_dff_B_hr2bwteo6_2),.clk(gclk));
	jdff dff_B_SPLLnP7V4_2(.din(w_dff_B_hr2bwteo6_2),.dout(w_dff_B_SPLLnP7V4_2),.clk(gclk));
	jdff dff_B_ZQK7VYsx0_2(.din(w_dff_B_SPLLnP7V4_2),.dout(w_dff_B_ZQK7VYsx0_2),.clk(gclk));
	jdff dff_B_eP6flCHu8_2(.din(w_dff_B_ZQK7VYsx0_2),.dout(w_dff_B_eP6flCHu8_2),.clk(gclk));
	jdff dff_B_brZIFypa5_2(.din(w_dff_B_eP6flCHu8_2),.dout(w_dff_B_brZIFypa5_2),.clk(gclk));
	jdff dff_B_pqV4ZWSR7_2(.din(w_dff_B_brZIFypa5_2),.dout(w_dff_B_pqV4ZWSR7_2),.clk(gclk));
	jdff dff_B_UYsBVN7x8_2(.din(w_dff_B_pqV4ZWSR7_2),.dout(w_dff_B_UYsBVN7x8_2),.clk(gclk));
	jdff dff_B_tBOkJJb40_2(.din(w_dff_B_UYsBVN7x8_2),.dout(w_dff_B_tBOkJJb40_2),.clk(gclk));
	jdff dff_B_nsVhCZI74_2(.din(w_dff_B_tBOkJJb40_2),.dout(w_dff_B_nsVhCZI74_2),.clk(gclk));
	jdff dff_B_cuijBt0D2_2(.din(w_dff_B_nsVhCZI74_2),.dout(w_dff_B_cuijBt0D2_2),.clk(gclk));
	jdff dff_B_9wj8SFYG0_2(.din(w_dff_B_cuijBt0D2_2),.dout(w_dff_B_9wj8SFYG0_2),.clk(gclk));
	jdff dff_B_tsTS65vP0_2(.din(w_dff_B_9wj8SFYG0_2),.dout(w_dff_B_tsTS65vP0_2),.clk(gclk));
	jdff dff_B_9Kcyb6XJ9_2(.din(w_dff_B_tsTS65vP0_2),.dout(w_dff_B_9Kcyb6XJ9_2),.clk(gclk));
	jdff dff_B_9PupgfsD7_2(.din(w_dff_B_9Kcyb6XJ9_2),.dout(w_dff_B_9PupgfsD7_2),.clk(gclk));
	jdff dff_B_6XqStstz9_2(.din(w_dff_B_9PupgfsD7_2),.dout(w_dff_B_6XqStstz9_2),.clk(gclk));
	jdff dff_B_6eOq1zfV8_2(.din(w_dff_B_6XqStstz9_2),.dout(w_dff_B_6eOq1zfV8_2),.clk(gclk));
	jdff dff_B_ILwT88TU8_2(.din(w_dff_B_6eOq1zfV8_2),.dout(w_dff_B_ILwT88TU8_2),.clk(gclk));
	jdff dff_B_BUWLskyo8_2(.din(w_dff_B_ILwT88TU8_2),.dout(w_dff_B_BUWLskyo8_2),.clk(gclk));
	jdff dff_B_N4sZZfxb6_2(.din(w_dff_B_BUWLskyo8_2),.dout(w_dff_B_N4sZZfxb6_2),.clk(gclk));
	jdff dff_B_eqDd9iGy1_2(.din(w_dff_B_N4sZZfxb6_2),.dout(w_dff_B_eqDd9iGy1_2),.clk(gclk));
	jdff dff_B_wpPzMh8I8_2(.din(w_dff_B_eqDd9iGy1_2),.dout(w_dff_B_wpPzMh8I8_2),.clk(gclk));
	jdff dff_B_c7gFdwpw1_2(.din(w_dff_B_wpPzMh8I8_2),.dout(w_dff_B_c7gFdwpw1_2),.clk(gclk));
	jdff dff_B_cIlPVjOn5_2(.din(w_dff_B_c7gFdwpw1_2),.dout(w_dff_B_cIlPVjOn5_2),.clk(gclk));
	jdff dff_B_NqV9IsLF5_2(.din(w_dff_B_cIlPVjOn5_2),.dout(w_dff_B_NqV9IsLF5_2),.clk(gclk));
	jdff dff_B_Rb0pOu6w7_2(.din(w_dff_B_NqV9IsLF5_2),.dout(w_dff_B_Rb0pOu6w7_2),.clk(gclk));
	jdff dff_B_662tQZJI7_2(.din(w_dff_B_Rb0pOu6w7_2),.dout(w_dff_B_662tQZJI7_2),.clk(gclk));
	jdff dff_B_kSVCW75S1_2(.din(w_dff_B_662tQZJI7_2),.dout(w_dff_B_kSVCW75S1_2),.clk(gclk));
	jdff dff_B_BJnENFj11_2(.din(w_dff_B_kSVCW75S1_2),.dout(w_dff_B_BJnENFj11_2),.clk(gclk));
	jdff dff_B_iPNammup2_2(.din(n1281),.dout(w_dff_B_iPNammup2_2),.clk(gclk));
	jdff dff_B_kV5BDMjF1_1(.din(n1243),.dout(w_dff_B_kV5BDMjF1_1),.clk(gclk));
	jdff dff_B_XhDtq3AJ2_2(.din(n1151),.dout(w_dff_B_XhDtq3AJ2_2),.clk(gclk));
	jdff dff_B_OtLSsN8s5_2(.din(w_dff_B_XhDtq3AJ2_2),.dout(w_dff_B_OtLSsN8s5_2),.clk(gclk));
	jdff dff_B_bnGijKmp3_2(.din(w_dff_B_OtLSsN8s5_2),.dout(w_dff_B_bnGijKmp3_2),.clk(gclk));
	jdff dff_B_hG63Xueq7_2(.din(w_dff_B_bnGijKmp3_2),.dout(w_dff_B_hG63Xueq7_2),.clk(gclk));
	jdff dff_B_n7O1Vi9l0_2(.din(w_dff_B_hG63Xueq7_2),.dout(w_dff_B_n7O1Vi9l0_2),.clk(gclk));
	jdff dff_B_EFcVe6XA3_2(.din(w_dff_B_n7O1Vi9l0_2),.dout(w_dff_B_EFcVe6XA3_2),.clk(gclk));
	jdff dff_B_gUOyplqD7_2(.din(w_dff_B_EFcVe6XA3_2),.dout(w_dff_B_gUOyplqD7_2),.clk(gclk));
	jdff dff_B_fOUSJ79E6_2(.din(w_dff_B_gUOyplqD7_2),.dout(w_dff_B_fOUSJ79E6_2),.clk(gclk));
	jdff dff_B_C8o3RLos2_2(.din(w_dff_B_fOUSJ79E6_2),.dout(w_dff_B_C8o3RLos2_2),.clk(gclk));
	jdff dff_B_pFQjw1tg7_2(.din(w_dff_B_C8o3RLos2_2),.dout(w_dff_B_pFQjw1tg7_2),.clk(gclk));
	jdff dff_B_FI3zd4kB1_2(.din(w_dff_B_pFQjw1tg7_2),.dout(w_dff_B_FI3zd4kB1_2),.clk(gclk));
	jdff dff_B_2OInZIqZ2_2(.din(w_dff_B_FI3zd4kB1_2),.dout(w_dff_B_2OInZIqZ2_2),.clk(gclk));
	jdff dff_B_UZfuMZFs9_2(.din(w_dff_B_2OInZIqZ2_2),.dout(w_dff_B_UZfuMZFs9_2),.clk(gclk));
	jdff dff_B_7JcPBHQe5_2(.din(w_dff_B_UZfuMZFs9_2),.dout(w_dff_B_7JcPBHQe5_2),.clk(gclk));
	jdff dff_B_ndH0dVsQ9_2(.din(w_dff_B_7JcPBHQe5_2),.dout(w_dff_B_ndH0dVsQ9_2),.clk(gclk));
	jdff dff_B_pkbBsHLO6_2(.din(w_dff_B_ndH0dVsQ9_2),.dout(w_dff_B_pkbBsHLO6_2),.clk(gclk));
	jdff dff_B_NnntY5257_2(.din(w_dff_B_pkbBsHLO6_2),.dout(w_dff_B_NnntY5257_2),.clk(gclk));
	jdff dff_B_iOERsrR15_2(.din(w_dff_B_NnntY5257_2),.dout(w_dff_B_iOERsrR15_2),.clk(gclk));
	jdff dff_B_XxpYyPVq8_2(.din(w_dff_B_iOERsrR15_2),.dout(w_dff_B_XxpYyPVq8_2),.clk(gclk));
	jdff dff_B_Q5tekKKe3_2(.din(w_dff_B_XxpYyPVq8_2),.dout(w_dff_B_Q5tekKKe3_2),.clk(gclk));
	jdff dff_B_vLguwKsV5_2(.din(w_dff_B_Q5tekKKe3_2),.dout(w_dff_B_vLguwKsV5_2),.clk(gclk));
	jdff dff_B_0dbO5Wv47_2(.din(w_dff_B_vLguwKsV5_2),.dout(w_dff_B_0dbO5Wv47_2),.clk(gclk));
	jdff dff_B_OtmVuPkN3_2(.din(w_dff_B_0dbO5Wv47_2),.dout(w_dff_B_OtmVuPkN3_2),.clk(gclk));
	jdff dff_B_zByO5G0a4_2(.din(w_dff_B_OtmVuPkN3_2),.dout(w_dff_B_zByO5G0a4_2),.clk(gclk));
	jdff dff_B_7Pig3tyK4_2(.din(w_dff_B_zByO5G0a4_2),.dout(w_dff_B_7Pig3tyK4_2),.clk(gclk));
	jdff dff_B_JryGpri68_2(.din(w_dff_B_7Pig3tyK4_2),.dout(w_dff_B_JryGpri68_2),.clk(gclk));
	jdff dff_B_Plxwei5y9_2(.din(n1190),.dout(w_dff_B_Plxwei5y9_2),.clk(gclk));
	jdff dff_B_OjcRlY2h2_1(.din(n1152),.dout(w_dff_B_OjcRlY2h2_1),.clk(gclk));
	jdff dff_B_HPLnmYZ77_2(.din(n1053),.dout(w_dff_B_HPLnmYZ77_2),.clk(gclk));
	jdff dff_B_LbOgLdUB8_2(.din(w_dff_B_HPLnmYZ77_2),.dout(w_dff_B_LbOgLdUB8_2),.clk(gclk));
	jdff dff_B_8NvYTmhn2_2(.din(w_dff_B_LbOgLdUB8_2),.dout(w_dff_B_8NvYTmhn2_2),.clk(gclk));
	jdff dff_B_MEBeBxjM5_2(.din(w_dff_B_8NvYTmhn2_2),.dout(w_dff_B_MEBeBxjM5_2),.clk(gclk));
	jdff dff_B_IGindAYx2_2(.din(w_dff_B_MEBeBxjM5_2),.dout(w_dff_B_IGindAYx2_2),.clk(gclk));
	jdff dff_B_ZQPs9dvB0_2(.din(w_dff_B_IGindAYx2_2),.dout(w_dff_B_ZQPs9dvB0_2),.clk(gclk));
	jdff dff_B_ZCpSSidV1_2(.din(w_dff_B_ZQPs9dvB0_2),.dout(w_dff_B_ZCpSSidV1_2),.clk(gclk));
	jdff dff_B_jXxu9ANi9_2(.din(w_dff_B_ZCpSSidV1_2),.dout(w_dff_B_jXxu9ANi9_2),.clk(gclk));
	jdff dff_B_tu67hxLv5_2(.din(w_dff_B_jXxu9ANi9_2),.dout(w_dff_B_tu67hxLv5_2),.clk(gclk));
	jdff dff_B_0blAYzrs3_2(.din(w_dff_B_tu67hxLv5_2),.dout(w_dff_B_0blAYzrs3_2),.clk(gclk));
	jdff dff_B_TbBUV0R14_2(.din(w_dff_B_0blAYzrs3_2),.dout(w_dff_B_TbBUV0R14_2),.clk(gclk));
	jdff dff_B_JDREr97s5_2(.din(w_dff_B_TbBUV0R14_2),.dout(w_dff_B_JDREr97s5_2),.clk(gclk));
	jdff dff_B_yb7PB9Q66_2(.din(w_dff_B_JDREr97s5_2),.dout(w_dff_B_yb7PB9Q66_2),.clk(gclk));
	jdff dff_B_nb3SKiOT1_2(.din(w_dff_B_yb7PB9Q66_2),.dout(w_dff_B_nb3SKiOT1_2),.clk(gclk));
	jdff dff_B_WWQgLknE4_2(.din(w_dff_B_nb3SKiOT1_2),.dout(w_dff_B_WWQgLknE4_2),.clk(gclk));
	jdff dff_B_3O4752CT8_2(.din(w_dff_B_WWQgLknE4_2),.dout(w_dff_B_3O4752CT8_2),.clk(gclk));
	jdff dff_B_vQ44mGwc6_2(.din(w_dff_B_3O4752CT8_2),.dout(w_dff_B_vQ44mGwc6_2),.clk(gclk));
	jdff dff_B_raAU1QSt2_2(.din(w_dff_B_vQ44mGwc6_2),.dout(w_dff_B_raAU1QSt2_2),.clk(gclk));
	jdff dff_B_mvcsrnVc6_2(.din(w_dff_B_raAU1QSt2_2),.dout(w_dff_B_mvcsrnVc6_2),.clk(gclk));
	jdff dff_B_TNAedXlp4_2(.din(w_dff_B_mvcsrnVc6_2),.dout(w_dff_B_TNAedXlp4_2),.clk(gclk));
	jdff dff_B_UNstYPRl4_2(.din(w_dff_B_TNAedXlp4_2),.dout(w_dff_B_UNstYPRl4_2),.clk(gclk));
	jdff dff_B_86jlqXc21_2(.din(w_dff_B_UNstYPRl4_2),.dout(w_dff_B_86jlqXc21_2),.clk(gclk));
	jdff dff_B_tSTxillR3_2(.din(w_dff_B_86jlqXc21_2),.dout(w_dff_B_tSTxillR3_2),.clk(gclk));
	jdff dff_B_hTlA5sbm7_2(.din(n1091),.dout(w_dff_B_hTlA5sbm7_2),.clk(gclk));
	jdff dff_B_4uKjXcCu3_1(.din(n1054),.dout(w_dff_B_4uKjXcCu3_1),.clk(gclk));
	jdff dff_B_fQlxMl3S2_2(.din(n954),.dout(w_dff_B_fQlxMl3S2_2),.clk(gclk));
	jdff dff_B_vOfmXFxe6_2(.din(w_dff_B_fQlxMl3S2_2),.dout(w_dff_B_vOfmXFxe6_2),.clk(gclk));
	jdff dff_B_Dnm3OYAp9_2(.din(w_dff_B_vOfmXFxe6_2),.dout(w_dff_B_Dnm3OYAp9_2),.clk(gclk));
	jdff dff_B_6BoHQNdw7_2(.din(w_dff_B_Dnm3OYAp9_2),.dout(w_dff_B_6BoHQNdw7_2),.clk(gclk));
	jdff dff_B_8skwEj4r5_2(.din(w_dff_B_6BoHQNdw7_2),.dout(w_dff_B_8skwEj4r5_2),.clk(gclk));
	jdff dff_B_SDPVJy5z0_2(.din(w_dff_B_8skwEj4r5_2),.dout(w_dff_B_SDPVJy5z0_2),.clk(gclk));
	jdff dff_B_1eEa4Tww7_2(.din(w_dff_B_SDPVJy5z0_2),.dout(w_dff_B_1eEa4Tww7_2),.clk(gclk));
	jdff dff_B_5oxYSuVg4_2(.din(w_dff_B_1eEa4Tww7_2),.dout(w_dff_B_5oxYSuVg4_2),.clk(gclk));
	jdff dff_B_qVWTOqfh8_2(.din(w_dff_B_5oxYSuVg4_2),.dout(w_dff_B_qVWTOqfh8_2),.clk(gclk));
	jdff dff_B_ebnHM4xV7_2(.din(w_dff_B_qVWTOqfh8_2),.dout(w_dff_B_ebnHM4xV7_2),.clk(gclk));
	jdff dff_B_NnQfzU9z1_2(.din(w_dff_B_ebnHM4xV7_2),.dout(w_dff_B_NnQfzU9z1_2),.clk(gclk));
	jdff dff_B_IozRSbbz6_2(.din(w_dff_B_NnQfzU9z1_2),.dout(w_dff_B_IozRSbbz6_2),.clk(gclk));
	jdff dff_B_vM7YJ0Xz1_2(.din(w_dff_B_IozRSbbz6_2),.dout(w_dff_B_vM7YJ0Xz1_2),.clk(gclk));
	jdff dff_B_qD9Fs3SU4_2(.din(w_dff_B_vM7YJ0Xz1_2),.dout(w_dff_B_qD9Fs3SU4_2),.clk(gclk));
	jdff dff_B_xmQi2xox5_2(.din(w_dff_B_qD9Fs3SU4_2),.dout(w_dff_B_xmQi2xox5_2),.clk(gclk));
	jdff dff_B_jBhYpXq06_2(.din(w_dff_B_xmQi2xox5_2),.dout(w_dff_B_jBhYpXq06_2),.clk(gclk));
	jdff dff_B_CAA55B1Q4_2(.din(w_dff_B_jBhYpXq06_2),.dout(w_dff_B_CAA55B1Q4_2),.clk(gclk));
	jdff dff_B_abYapm3v1_2(.din(w_dff_B_CAA55B1Q4_2),.dout(w_dff_B_abYapm3v1_2),.clk(gclk));
	jdff dff_B_x7NgL6XT6_2(.din(w_dff_B_abYapm3v1_2),.dout(w_dff_B_x7NgL6XT6_2),.clk(gclk));
	jdff dff_B_f5N2DkNH4_2(.din(w_dff_B_x7NgL6XT6_2),.dout(w_dff_B_f5N2DkNH4_2),.clk(gclk));
	jdff dff_B_D286X2Hh9_2(.din(n992),.dout(w_dff_B_D286X2Hh9_2),.clk(gclk));
	jdff dff_B_UxsF3NTc2_1(.din(n955),.dout(w_dff_B_UxsF3NTc2_1),.clk(gclk));
	jdff dff_B_hX83ipm33_2(.din(n852),.dout(w_dff_B_hX83ipm33_2),.clk(gclk));
	jdff dff_B_zHvMk9Xz7_2(.din(w_dff_B_hX83ipm33_2),.dout(w_dff_B_zHvMk9Xz7_2),.clk(gclk));
	jdff dff_B_HWcn8jjT1_2(.din(w_dff_B_zHvMk9Xz7_2),.dout(w_dff_B_HWcn8jjT1_2),.clk(gclk));
	jdff dff_B_mGgKSy1w6_2(.din(w_dff_B_HWcn8jjT1_2),.dout(w_dff_B_mGgKSy1w6_2),.clk(gclk));
	jdff dff_B_LkwT9Bz25_2(.din(w_dff_B_mGgKSy1w6_2),.dout(w_dff_B_LkwT9Bz25_2),.clk(gclk));
	jdff dff_B_UygJsp3C1_2(.din(w_dff_B_LkwT9Bz25_2),.dout(w_dff_B_UygJsp3C1_2),.clk(gclk));
	jdff dff_B_Fj9SQ95y6_2(.din(w_dff_B_UygJsp3C1_2),.dout(w_dff_B_Fj9SQ95y6_2),.clk(gclk));
	jdff dff_B_OOIce2499_2(.din(w_dff_B_Fj9SQ95y6_2),.dout(w_dff_B_OOIce2499_2),.clk(gclk));
	jdff dff_B_fCJYw80P6_2(.din(w_dff_B_OOIce2499_2),.dout(w_dff_B_fCJYw80P6_2),.clk(gclk));
	jdff dff_B_3bHjyah09_2(.din(w_dff_B_fCJYw80P6_2),.dout(w_dff_B_3bHjyah09_2),.clk(gclk));
	jdff dff_B_Bz4Qlem84_2(.din(w_dff_B_3bHjyah09_2),.dout(w_dff_B_Bz4Qlem84_2),.clk(gclk));
	jdff dff_B_5G53VeFP1_2(.din(w_dff_B_Bz4Qlem84_2),.dout(w_dff_B_5G53VeFP1_2),.clk(gclk));
	jdff dff_B_ydf0zOwQ6_2(.din(w_dff_B_5G53VeFP1_2),.dout(w_dff_B_ydf0zOwQ6_2),.clk(gclk));
	jdff dff_B_Mr9PeNBM7_2(.din(w_dff_B_ydf0zOwQ6_2),.dout(w_dff_B_Mr9PeNBM7_2),.clk(gclk));
	jdff dff_B_mijPNv5Q7_2(.din(w_dff_B_Mr9PeNBM7_2),.dout(w_dff_B_mijPNv5Q7_2),.clk(gclk));
	jdff dff_B_EfAza7EV0_2(.din(w_dff_B_mijPNv5Q7_2),.dout(w_dff_B_EfAza7EV0_2),.clk(gclk));
	jdff dff_B_QFBFxzKh3_2(.din(w_dff_B_EfAza7EV0_2),.dout(w_dff_B_QFBFxzKh3_2),.clk(gclk));
	jdff dff_B_FYrpa1pl8_2(.din(n886),.dout(w_dff_B_FYrpa1pl8_2),.clk(gclk));
	jdff dff_B_0SQLVANx9_1(.din(n853),.dout(w_dff_B_0SQLVANx9_1),.clk(gclk));
	jdff dff_B_JMyW1ypF9_2(.din(n754),.dout(w_dff_B_JMyW1ypF9_2),.clk(gclk));
	jdff dff_B_ZabHqtev9_2(.din(w_dff_B_JMyW1ypF9_2),.dout(w_dff_B_ZabHqtev9_2),.clk(gclk));
	jdff dff_B_IgmttBZF3_2(.din(w_dff_B_ZabHqtev9_2),.dout(w_dff_B_IgmttBZF3_2),.clk(gclk));
	jdff dff_B_kxWji1ZO6_2(.din(w_dff_B_IgmttBZF3_2),.dout(w_dff_B_kxWji1ZO6_2),.clk(gclk));
	jdff dff_B_d0AN3yjj9_2(.din(w_dff_B_kxWji1ZO6_2),.dout(w_dff_B_d0AN3yjj9_2),.clk(gclk));
	jdff dff_B_Yyo1N9A11_2(.din(w_dff_B_d0AN3yjj9_2),.dout(w_dff_B_Yyo1N9A11_2),.clk(gclk));
	jdff dff_B_vNMxwU1F8_2(.din(w_dff_B_Yyo1N9A11_2),.dout(w_dff_B_vNMxwU1F8_2),.clk(gclk));
	jdff dff_B_WhY8Jqys4_2(.din(w_dff_B_vNMxwU1F8_2),.dout(w_dff_B_WhY8Jqys4_2),.clk(gclk));
	jdff dff_B_E0b8Qx8l9_2(.din(w_dff_B_WhY8Jqys4_2),.dout(w_dff_B_E0b8Qx8l9_2),.clk(gclk));
	jdff dff_B_FGUSWCTU2_2(.din(w_dff_B_E0b8Qx8l9_2),.dout(w_dff_B_FGUSWCTU2_2),.clk(gclk));
	jdff dff_B_wZjoefnz4_2(.din(w_dff_B_FGUSWCTU2_2),.dout(w_dff_B_wZjoefnz4_2),.clk(gclk));
	jdff dff_B_DLMpgKeL7_2(.din(w_dff_B_wZjoefnz4_2),.dout(w_dff_B_DLMpgKeL7_2),.clk(gclk));
	jdff dff_B_KgWTyaJP3_2(.din(w_dff_B_DLMpgKeL7_2),.dout(w_dff_B_KgWTyaJP3_2),.clk(gclk));
	jdff dff_B_VRnjLZMF3_2(.din(w_dff_B_KgWTyaJP3_2),.dout(w_dff_B_VRnjLZMF3_2),.clk(gclk));
	jdff dff_B_1GKvZS0y0_2(.din(n783),.dout(w_dff_B_1GKvZS0y0_2),.clk(gclk));
	jdff dff_B_L9dAiNeY6_1(.din(n755),.dout(w_dff_B_L9dAiNeY6_1),.clk(gclk));
	jdff dff_B_2hQyrjfp5_2(.din(n662),.dout(w_dff_B_2hQyrjfp5_2),.clk(gclk));
	jdff dff_B_BOZk9Qht4_2(.din(w_dff_B_2hQyrjfp5_2),.dout(w_dff_B_BOZk9Qht4_2),.clk(gclk));
	jdff dff_B_r1xfYZN53_2(.din(w_dff_B_BOZk9Qht4_2),.dout(w_dff_B_r1xfYZN53_2),.clk(gclk));
	jdff dff_B_EPQRGGMb7_2(.din(w_dff_B_r1xfYZN53_2),.dout(w_dff_B_EPQRGGMb7_2),.clk(gclk));
	jdff dff_B_iIKiHArP0_2(.din(w_dff_B_EPQRGGMb7_2),.dout(w_dff_B_iIKiHArP0_2),.clk(gclk));
	jdff dff_B_Eu9Ud1cb9_2(.din(w_dff_B_iIKiHArP0_2),.dout(w_dff_B_Eu9Ud1cb9_2),.clk(gclk));
	jdff dff_B_kH1awpSJ2_2(.din(w_dff_B_Eu9Ud1cb9_2),.dout(w_dff_B_kH1awpSJ2_2),.clk(gclk));
	jdff dff_B_epbDVz3U0_2(.din(w_dff_B_kH1awpSJ2_2),.dout(w_dff_B_epbDVz3U0_2),.clk(gclk));
	jdff dff_B_KZTDu68j0_2(.din(w_dff_B_epbDVz3U0_2),.dout(w_dff_B_KZTDu68j0_2),.clk(gclk));
	jdff dff_B_v20WeeIt3_2(.din(w_dff_B_KZTDu68j0_2),.dout(w_dff_B_v20WeeIt3_2),.clk(gclk));
	jdff dff_B_RmOrkIc96_2(.din(w_dff_B_v20WeeIt3_2),.dout(w_dff_B_RmOrkIc96_2),.clk(gclk));
	jdff dff_B_6vOacekQ0_2(.din(n684),.dout(w_dff_B_6vOacekQ0_2),.clk(gclk));
	jdff dff_B_fhsB5pI32_1(.din(n663),.dout(w_dff_B_fhsB5pI32_1),.clk(gclk));
	jdff dff_B_j6r1Pr0z6_2(.din(n577),.dout(w_dff_B_j6r1Pr0z6_2),.clk(gclk));
	jdff dff_B_RyfUBfVm0_2(.din(w_dff_B_j6r1Pr0z6_2),.dout(w_dff_B_RyfUBfVm0_2),.clk(gclk));
	jdff dff_B_ZW9y5cSy0_2(.din(w_dff_B_RyfUBfVm0_2),.dout(w_dff_B_ZW9y5cSy0_2),.clk(gclk));
	jdff dff_B_zvjJeL4G4_2(.din(w_dff_B_ZW9y5cSy0_2),.dout(w_dff_B_zvjJeL4G4_2),.clk(gclk));
	jdff dff_B_oPHvr82C4_2(.din(w_dff_B_zvjJeL4G4_2),.dout(w_dff_B_oPHvr82C4_2),.clk(gclk));
	jdff dff_B_Gng1ttnp6_2(.din(w_dff_B_oPHvr82C4_2),.dout(w_dff_B_Gng1ttnp6_2),.clk(gclk));
	jdff dff_B_IDqVQHuX0_2(.din(w_dff_B_Gng1ttnp6_2),.dout(w_dff_B_IDqVQHuX0_2),.clk(gclk));
	jdff dff_B_SF8nTlbT9_2(.din(w_dff_B_IDqVQHuX0_2),.dout(w_dff_B_SF8nTlbT9_2),.clk(gclk));
	jdff dff_B_1peuGQj02_2(.din(n592),.dout(w_dff_B_1peuGQj02_2),.clk(gclk));
	jdff dff_B_ioxh8fVC2_2(.din(w_dff_B_1peuGQj02_2),.dout(w_dff_B_ioxh8fVC2_2),.clk(gclk));
	jdff dff_B_7qNLUpmv4_2(.din(w_dff_B_ioxh8fVC2_2),.dout(w_dff_B_7qNLUpmv4_2),.clk(gclk));
	jdff dff_B_4LAuJUSU0_1(.din(n578),.dout(w_dff_B_4LAuJUSU0_1),.clk(gclk));
	jdff dff_B_Zdg8hQQA3_1(.din(w_dff_B_4LAuJUSU0_1),.dout(w_dff_B_Zdg8hQQA3_1),.clk(gclk));
	jdff dff_B_ESJgNDMp1_2(.din(n501),.dout(w_dff_B_ESJgNDMp1_2),.clk(gclk));
	jdff dff_B_L6eWh6e09_2(.din(w_dff_B_ESJgNDMp1_2),.dout(w_dff_B_L6eWh6e09_2),.clk(gclk));
	jdff dff_B_7ZZLxOsm6_2(.din(w_dff_B_L6eWh6e09_2),.dout(w_dff_B_7ZZLxOsm6_2),.clk(gclk));
	jdff dff_B_pZTOoJE89_0(.din(n506),.dout(w_dff_B_pZTOoJE89_0),.clk(gclk));
	jdff dff_A_5Se624DU4_0(.dout(w_n427_0[0]),.din(w_dff_A_5Se624DU4_0),.clk(gclk));
	jdff dff_A_tI7GeNyK3_0(.dout(w_dff_A_5Se624DU4_0),.din(w_dff_A_tI7GeNyK3_0),.clk(gclk));
	jdff dff_A_ZWzEZO8B7_1(.dout(w_n427_0[1]),.din(w_dff_A_ZWzEZO8B7_1),.clk(gclk));
	jdff dff_A_4MM8phz66_1(.dout(w_dff_A_ZWzEZO8B7_1),.din(w_dff_A_4MM8phz66_1),.clk(gclk));
	jdff dff_B_GwYof2122_1(.din(n1729),.dout(w_dff_B_GwYof2122_1),.clk(gclk));
	jdff dff_A_SwQ6ri8m3_1(.dout(w_n1697_0[1]),.din(w_dff_A_SwQ6ri8m3_1),.clk(gclk));
	jdff dff_B_2BO5H3Fh3_1(.din(n1695),.dout(w_dff_B_2BO5H3Fh3_1),.clk(gclk));
	jdff dff_B_RcXJoA6M0_2(.din(n1653),.dout(w_dff_B_RcXJoA6M0_2),.clk(gclk));
	jdff dff_B_Y2oKoKr14_2(.din(w_dff_B_RcXJoA6M0_2),.dout(w_dff_B_Y2oKoKr14_2),.clk(gclk));
	jdff dff_B_AqPVFHW88_2(.din(w_dff_B_Y2oKoKr14_2),.dout(w_dff_B_AqPVFHW88_2),.clk(gclk));
	jdff dff_B_LXSgQJGn9_2(.din(w_dff_B_AqPVFHW88_2),.dout(w_dff_B_LXSgQJGn9_2),.clk(gclk));
	jdff dff_B_tnyuM3JP5_2(.din(w_dff_B_LXSgQJGn9_2),.dout(w_dff_B_tnyuM3JP5_2),.clk(gclk));
	jdff dff_B_EsATly1H6_2(.din(w_dff_B_tnyuM3JP5_2),.dout(w_dff_B_EsATly1H6_2),.clk(gclk));
	jdff dff_B_drNmJrFC1_2(.din(w_dff_B_EsATly1H6_2),.dout(w_dff_B_drNmJrFC1_2),.clk(gclk));
	jdff dff_B_IZfbzlGw3_2(.din(w_dff_B_drNmJrFC1_2),.dout(w_dff_B_IZfbzlGw3_2),.clk(gclk));
	jdff dff_B_kwFoYC738_2(.din(w_dff_B_IZfbzlGw3_2),.dout(w_dff_B_kwFoYC738_2),.clk(gclk));
	jdff dff_B_48rGiQOT0_2(.din(w_dff_B_kwFoYC738_2),.dout(w_dff_B_48rGiQOT0_2),.clk(gclk));
	jdff dff_B_SJPeioDR3_2(.din(w_dff_B_48rGiQOT0_2),.dout(w_dff_B_SJPeioDR3_2),.clk(gclk));
	jdff dff_B_lFPka0Mg0_2(.din(w_dff_B_SJPeioDR3_2),.dout(w_dff_B_lFPka0Mg0_2),.clk(gclk));
	jdff dff_B_q4jIGpo08_2(.din(w_dff_B_lFPka0Mg0_2),.dout(w_dff_B_q4jIGpo08_2),.clk(gclk));
	jdff dff_B_6I0723fN9_2(.din(w_dff_B_q4jIGpo08_2),.dout(w_dff_B_6I0723fN9_2),.clk(gclk));
	jdff dff_B_4Rmj2au51_2(.din(w_dff_B_6I0723fN9_2),.dout(w_dff_B_4Rmj2au51_2),.clk(gclk));
	jdff dff_B_QsbgupvY5_2(.din(w_dff_B_4Rmj2au51_2),.dout(w_dff_B_QsbgupvY5_2),.clk(gclk));
	jdff dff_B_gR31hLuU8_2(.din(w_dff_B_QsbgupvY5_2),.dout(w_dff_B_gR31hLuU8_2),.clk(gclk));
	jdff dff_B_ayIruosr3_2(.din(w_dff_B_gR31hLuU8_2),.dout(w_dff_B_ayIruosr3_2),.clk(gclk));
	jdff dff_B_FR4NXnEc2_2(.din(w_dff_B_ayIruosr3_2),.dout(w_dff_B_FR4NXnEc2_2),.clk(gclk));
	jdff dff_B_U8P0ZI8H6_2(.din(w_dff_B_FR4NXnEc2_2),.dout(w_dff_B_U8P0ZI8H6_2),.clk(gclk));
	jdff dff_B_3uuSu37e9_2(.din(w_dff_B_U8P0ZI8H6_2),.dout(w_dff_B_3uuSu37e9_2),.clk(gclk));
	jdff dff_B_pJgnBA9L0_2(.din(w_dff_B_3uuSu37e9_2),.dout(w_dff_B_pJgnBA9L0_2),.clk(gclk));
	jdff dff_B_oMVFEaJZ8_2(.din(w_dff_B_pJgnBA9L0_2),.dout(w_dff_B_oMVFEaJZ8_2),.clk(gclk));
	jdff dff_B_SNcH6jEJ1_2(.din(w_dff_B_oMVFEaJZ8_2),.dout(w_dff_B_SNcH6jEJ1_2),.clk(gclk));
	jdff dff_B_Y9glgvmM9_2(.din(w_dff_B_SNcH6jEJ1_2),.dout(w_dff_B_Y9glgvmM9_2),.clk(gclk));
	jdff dff_B_FSEjjpyd0_2(.din(w_dff_B_Y9glgvmM9_2),.dout(w_dff_B_FSEjjpyd0_2),.clk(gclk));
	jdff dff_B_1crG85sG9_2(.din(w_dff_B_FSEjjpyd0_2),.dout(w_dff_B_1crG85sG9_2),.clk(gclk));
	jdff dff_B_vTiA19Pk2_2(.din(w_dff_B_1crG85sG9_2),.dout(w_dff_B_vTiA19Pk2_2),.clk(gclk));
	jdff dff_B_Lyc5LJAo0_2(.din(w_dff_B_vTiA19Pk2_2),.dout(w_dff_B_Lyc5LJAo0_2),.clk(gclk));
	jdff dff_B_bGXVEpuy0_2(.din(w_dff_B_Lyc5LJAo0_2),.dout(w_dff_B_bGXVEpuy0_2),.clk(gclk));
	jdff dff_B_mSs1jPUu0_2(.din(w_dff_B_bGXVEpuy0_2),.dout(w_dff_B_mSs1jPUu0_2),.clk(gclk));
	jdff dff_B_Pku4wRHZ5_2(.din(w_dff_B_mSs1jPUu0_2),.dout(w_dff_B_Pku4wRHZ5_2),.clk(gclk));
	jdff dff_B_B7nL4GdN8_2(.din(w_dff_B_Pku4wRHZ5_2),.dout(w_dff_B_B7nL4GdN8_2),.clk(gclk));
	jdff dff_B_KGXfH1jC9_2(.din(w_dff_B_B7nL4GdN8_2),.dout(w_dff_B_KGXfH1jC9_2),.clk(gclk));
	jdff dff_B_J2KmmILp8_2(.din(w_dff_B_KGXfH1jC9_2),.dout(w_dff_B_J2KmmILp8_2),.clk(gclk));
	jdff dff_B_OJ7Z7NdO4_2(.din(w_dff_B_J2KmmILp8_2),.dout(w_dff_B_OJ7Z7NdO4_2),.clk(gclk));
	jdff dff_B_4gXtPzDy4_2(.din(w_dff_B_OJ7Z7NdO4_2),.dout(w_dff_B_4gXtPzDy4_2),.clk(gclk));
	jdff dff_B_JGdoBNXQ8_2(.din(w_dff_B_4gXtPzDy4_2),.dout(w_dff_B_JGdoBNXQ8_2),.clk(gclk));
	jdff dff_B_VD9mQd8f7_2(.din(w_dff_B_JGdoBNXQ8_2),.dout(w_dff_B_VD9mQd8f7_2),.clk(gclk));
	jdff dff_B_Ch4NS9AK4_2(.din(w_dff_B_VD9mQd8f7_2),.dout(w_dff_B_Ch4NS9AK4_2),.clk(gclk));
	jdff dff_B_J1tycnE23_2(.din(w_dff_B_Ch4NS9AK4_2),.dout(w_dff_B_J1tycnE23_2),.clk(gclk));
	jdff dff_B_aVyGAD361_2(.din(w_dff_B_J1tycnE23_2),.dout(w_dff_B_aVyGAD361_2),.clk(gclk));
	jdff dff_B_7v498nzy0_2(.din(w_dff_B_aVyGAD361_2),.dout(w_dff_B_7v498nzy0_2),.clk(gclk));
	jdff dff_B_JaHyIaEv7_2(.din(w_dff_B_7v498nzy0_2),.dout(w_dff_B_JaHyIaEv7_2),.clk(gclk));
	jdff dff_B_0Z2jdXNz8_2(.din(w_dff_B_JaHyIaEv7_2),.dout(w_dff_B_0Z2jdXNz8_2),.clk(gclk));
	jdff dff_B_nBxfy3Zo3_2(.din(w_dff_B_0Z2jdXNz8_2),.dout(w_dff_B_nBxfy3Zo3_2),.clk(gclk));
	jdff dff_B_toABSUla3_2(.din(n1656),.dout(w_dff_B_toABSUla3_2),.clk(gclk));
	jdff dff_B_fL374ioq5_1(.din(n1654),.dout(w_dff_B_fL374ioq5_1),.clk(gclk));
	jdff dff_B_srz84Pgv4_2(.din(n1602),.dout(w_dff_B_srz84Pgv4_2),.clk(gclk));
	jdff dff_B_sUGcgf2X2_2(.din(w_dff_B_srz84Pgv4_2),.dout(w_dff_B_sUGcgf2X2_2),.clk(gclk));
	jdff dff_B_RUO0MwKQ6_2(.din(w_dff_B_sUGcgf2X2_2),.dout(w_dff_B_RUO0MwKQ6_2),.clk(gclk));
	jdff dff_B_5CxXe5pG9_2(.din(w_dff_B_RUO0MwKQ6_2),.dout(w_dff_B_5CxXe5pG9_2),.clk(gclk));
	jdff dff_B_50FqWL0Y6_2(.din(w_dff_B_5CxXe5pG9_2),.dout(w_dff_B_50FqWL0Y6_2),.clk(gclk));
	jdff dff_B_ArT0Qvck4_2(.din(w_dff_B_50FqWL0Y6_2),.dout(w_dff_B_ArT0Qvck4_2),.clk(gclk));
	jdff dff_B_QYaoqqG31_2(.din(w_dff_B_ArT0Qvck4_2),.dout(w_dff_B_QYaoqqG31_2),.clk(gclk));
	jdff dff_B_bRblvbew7_2(.din(w_dff_B_QYaoqqG31_2),.dout(w_dff_B_bRblvbew7_2),.clk(gclk));
	jdff dff_B_WLVMwxOw3_2(.din(w_dff_B_bRblvbew7_2),.dout(w_dff_B_WLVMwxOw3_2),.clk(gclk));
	jdff dff_B_vqFZ7Nlo6_2(.din(w_dff_B_WLVMwxOw3_2),.dout(w_dff_B_vqFZ7Nlo6_2),.clk(gclk));
	jdff dff_B_azEYAeet3_2(.din(w_dff_B_vqFZ7Nlo6_2),.dout(w_dff_B_azEYAeet3_2),.clk(gclk));
	jdff dff_B_6GDNLp3L0_2(.din(w_dff_B_azEYAeet3_2),.dout(w_dff_B_6GDNLp3L0_2),.clk(gclk));
	jdff dff_B_GR1mAU6h5_2(.din(w_dff_B_6GDNLp3L0_2),.dout(w_dff_B_GR1mAU6h5_2),.clk(gclk));
	jdff dff_B_iG84c0cQ4_2(.din(w_dff_B_GR1mAU6h5_2),.dout(w_dff_B_iG84c0cQ4_2),.clk(gclk));
	jdff dff_B_c0IoGkQP4_2(.din(w_dff_B_iG84c0cQ4_2),.dout(w_dff_B_c0IoGkQP4_2),.clk(gclk));
	jdff dff_B_gmBvsdYM9_2(.din(w_dff_B_c0IoGkQP4_2),.dout(w_dff_B_gmBvsdYM9_2),.clk(gclk));
	jdff dff_B_NrddrdD48_2(.din(w_dff_B_gmBvsdYM9_2),.dout(w_dff_B_NrddrdD48_2),.clk(gclk));
	jdff dff_B_qbGeRZxD1_2(.din(w_dff_B_NrddrdD48_2),.dout(w_dff_B_qbGeRZxD1_2),.clk(gclk));
	jdff dff_B_2ser7ZdF1_2(.din(w_dff_B_qbGeRZxD1_2),.dout(w_dff_B_2ser7ZdF1_2),.clk(gclk));
	jdff dff_B_47goirtf3_2(.din(w_dff_B_2ser7ZdF1_2),.dout(w_dff_B_47goirtf3_2),.clk(gclk));
	jdff dff_B_D7XGDyVJ9_2(.din(w_dff_B_47goirtf3_2),.dout(w_dff_B_D7XGDyVJ9_2),.clk(gclk));
	jdff dff_B_sHbW1fKC7_2(.din(w_dff_B_D7XGDyVJ9_2),.dout(w_dff_B_sHbW1fKC7_2),.clk(gclk));
	jdff dff_B_0Vhg79P96_2(.din(w_dff_B_sHbW1fKC7_2),.dout(w_dff_B_0Vhg79P96_2),.clk(gclk));
	jdff dff_B_hvuTvXpA6_2(.din(w_dff_B_0Vhg79P96_2),.dout(w_dff_B_hvuTvXpA6_2),.clk(gclk));
	jdff dff_B_5xX9sl2J5_2(.din(w_dff_B_hvuTvXpA6_2),.dout(w_dff_B_5xX9sl2J5_2),.clk(gclk));
	jdff dff_B_NQN0w1Pi1_2(.din(w_dff_B_5xX9sl2J5_2),.dout(w_dff_B_NQN0w1Pi1_2),.clk(gclk));
	jdff dff_B_Ch0jz0Lk7_2(.din(w_dff_B_NQN0w1Pi1_2),.dout(w_dff_B_Ch0jz0Lk7_2),.clk(gclk));
	jdff dff_B_6RVLTVQF5_2(.din(w_dff_B_Ch0jz0Lk7_2),.dout(w_dff_B_6RVLTVQF5_2),.clk(gclk));
	jdff dff_B_VKIDSFkq0_2(.din(w_dff_B_6RVLTVQF5_2),.dout(w_dff_B_VKIDSFkq0_2),.clk(gclk));
	jdff dff_B_6WOtqA6l9_2(.din(w_dff_B_VKIDSFkq0_2),.dout(w_dff_B_6WOtqA6l9_2),.clk(gclk));
	jdff dff_B_EUwzOq7b3_2(.din(w_dff_B_6WOtqA6l9_2),.dout(w_dff_B_EUwzOq7b3_2),.clk(gclk));
	jdff dff_B_YLDpHNXV0_2(.din(w_dff_B_EUwzOq7b3_2),.dout(w_dff_B_YLDpHNXV0_2),.clk(gclk));
	jdff dff_B_36NqWeYd2_2(.din(w_dff_B_YLDpHNXV0_2),.dout(w_dff_B_36NqWeYd2_2),.clk(gclk));
	jdff dff_B_2brQbtMX9_2(.din(w_dff_B_36NqWeYd2_2),.dout(w_dff_B_2brQbtMX9_2),.clk(gclk));
	jdff dff_B_DqxQL4XO5_2(.din(w_dff_B_2brQbtMX9_2),.dout(w_dff_B_DqxQL4XO5_2),.clk(gclk));
	jdff dff_B_NniZN1Ep7_2(.din(w_dff_B_DqxQL4XO5_2),.dout(w_dff_B_NniZN1Ep7_2),.clk(gclk));
	jdff dff_B_mgg01KfN9_2(.din(w_dff_B_NniZN1Ep7_2),.dout(w_dff_B_mgg01KfN9_2),.clk(gclk));
	jdff dff_B_O9TiFwU31_2(.din(w_dff_B_mgg01KfN9_2),.dout(w_dff_B_O9TiFwU31_2),.clk(gclk));
	jdff dff_B_KzSalANb9_2(.din(w_dff_B_O9TiFwU31_2),.dout(w_dff_B_KzSalANb9_2),.clk(gclk));
	jdff dff_B_Z8fkM5Ii2_2(.din(w_dff_B_KzSalANb9_2),.dout(w_dff_B_Z8fkM5Ii2_2),.clk(gclk));
	jdff dff_B_IPbenLDB9_2(.din(w_dff_B_Z8fkM5Ii2_2),.dout(w_dff_B_IPbenLDB9_2),.clk(gclk));
	jdff dff_B_7sCSoUGO2_2(.din(w_dff_B_IPbenLDB9_2),.dout(w_dff_B_7sCSoUGO2_2),.clk(gclk));
	jdff dff_B_JeVevLGF2_2(.din(n1605),.dout(w_dff_B_JeVevLGF2_2),.clk(gclk));
	jdff dff_B_72FCd2WI3_1(.din(n1603),.dout(w_dff_B_72FCd2WI3_1),.clk(gclk));
	jdff dff_B_0Vkd3RTi3_2(.din(n1545),.dout(w_dff_B_0Vkd3RTi3_2),.clk(gclk));
	jdff dff_B_viszoCbb1_2(.din(w_dff_B_0Vkd3RTi3_2),.dout(w_dff_B_viszoCbb1_2),.clk(gclk));
	jdff dff_B_HKpayDrq0_2(.din(w_dff_B_viszoCbb1_2),.dout(w_dff_B_HKpayDrq0_2),.clk(gclk));
	jdff dff_B_E9oVdWO76_2(.din(w_dff_B_HKpayDrq0_2),.dout(w_dff_B_E9oVdWO76_2),.clk(gclk));
	jdff dff_B_jhOmsjKU5_2(.din(w_dff_B_E9oVdWO76_2),.dout(w_dff_B_jhOmsjKU5_2),.clk(gclk));
	jdff dff_B_xtnw1jPq3_2(.din(w_dff_B_jhOmsjKU5_2),.dout(w_dff_B_xtnw1jPq3_2),.clk(gclk));
	jdff dff_B_vMVUCDk53_2(.din(w_dff_B_xtnw1jPq3_2),.dout(w_dff_B_vMVUCDk53_2),.clk(gclk));
	jdff dff_B_LLlFAXGO4_2(.din(w_dff_B_vMVUCDk53_2),.dout(w_dff_B_LLlFAXGO4_2),.clk(gclk));
	jdff dff_B_WSTci83g3_2(.din(w_dff_B_LLlFAXGO4_2),.dout(w_dff_B_WSTci83g3_2),.clk(gclk));
	jdff dff_B_Sy19B0WV3_2(.din(w_dff_B_WSTci83g3_2),.dout(w_dff_B_Sy19B0WV3_2),.clk(gclk));
	jdff dff_B_hSeXNY4M3_2(.din(w_dff_B_Sy19B0WV3_2),.dout(w_dff_B_hSeXNY4M3_2),.clk(gclk));
	jdff dff_B_knrWhgjB0_2(.din(w_dff_B_hSeXNY4M3_2),.dout(w_dff_B_knrWhgjB0_2),.clk(gclk));
	jdff dff_B_AlE2HCrZ7_2(.din(w_dff_B_knrWhgjB0_2),.dout(w_dff_B_AlE2HCrZ7_2),.clk(gclk));
	jdff dff_B_pUKBjtUL4_2(.din(w_dff_B_AlE2HCrZ7_2),.dout(w_dff_B_pUKBjtUL4_2),.clk(gclk));
	jdff dff_B_x9Vc4eVj3_2(.din(w_dff_B_pUKBjtUL4_2),.dout(w_dff_B_x9Vc4eVj3_2),.clk(gclk));
	jdff dff_B_YlLyWT2v8_2(.din(w_dff_B_x9Vc4eVj3_2),.dout(w_dff_B_YlLyWT2v8_2),.clk(gclk));
	jdff dff_B_hE1A2bxz0_2(.din(w_dff_B_YlLyWT2v8_2),.dout(w_dff_B_hE1A2bxz0_2),.clk(gclk));
	jdff dff_B_RViGyZXN7_2(.din(w_dff_B_hE1A2bxz0_2),.dout(w_dff_B_RViGyZXN7_2),.clk(gclk));
	jdff dff_B_js2biHo04_2(.din(w_dff_B_RViGyZXN7_2),.dout(w_dff_B_js2biHo04_2),.clk(gclk));
	jdff dff_B_WXYXMVMO7_2(.din(w_dff_B_js2biHo04_2),.dout(w_dff_B_WXYXMVMO7_2),.clk(gclk));
	jdff dff_B_P71syNyq0_2(.din(w_dff_B_WXYXMVMO7_2),.dout(w_dff_B_P71syNyq0_2),.clk(gclk));
	jdff dff_B_3ubAaHD18_2(.din(w_dff_B_P71syNyq0_2),.dout(w_dff_B_3ubAaHD18_2),.clk(gclk));
	jdff dff_B_ZKTx0qP55_2(.din(w_dff_B_3ubAaHD18_2),.dout(w_dff_B_ZKTx0qP55_2),.clk(gclk));
	jdff dff_B_NRRn0mRd2_2(.din(w_dff_B_ZKTx0qP55_2),.dout(w_dff_B_NRRn0mRd2_2),.clk(gclk));
	jdff dff_B_qGaMJt2o9_2(.din(w_dff_B_NRRn0mRd2_2),.dout(w_dff_B_qGaMJt2o9_2),.clk(gclk));
	jdff dff_B_UOKfX48y1_2(.din(w_dff_B_qGaMJt2o9_2),.dout(w_dff_B_UOKfX48y1_2),.clk(gclk));
	jdff dff_B_UAhTtrPE9_2(.din(w_dff_B_UOKfX48y1_2),.dout(w_dff_B_UAhTtrPE9_2),.clk(gclk));
	jdff dff_B_qp6leGgL9_2(.din(w_dff_B_UAhTtrPE9_2),.dout(w_dff_B_qp6leGgL9_2),.clk(gclk));
	jdff dff_B_Fun1EjNk6_2(.din(w_dff_B_qp6leGgL9_2),.dout(w_dff_B_Fun1EjNk6_2),.clk(gclk));
	jdff dff_B_9F7rfMuK1_2(.din(w_dff_B_Fun1EjNk6_2),.dout(w_dff_B_9F7rfMuK1_2),.clk(gclk));
	jdff dff_B_N588Bo4B8_2(.din(w_dff_B_9F7rfMuK1_2),.dout(w_dff_B_N588Bo4B8_2),.clk(gclk));
	jdff dff_B_jIJU7zvh7_2(.din(w_dff_B_N588Bo4B8_2),.dout(w_dff_B_jIJU7zvh7_2),.clk(gclk));
	jdff dff_B_ywrMII1O9_2(.din(w_dff_B_jIJU7zvh7_2),.dout(w_dff_B_ywrMII1O9_2),.clk(gclk));
	jdff dff_B_HHFWSoPB6_2(.din(w_dff_B_ywrMII1O9_2),.dout(w_dff_B_HHFWSoPB6_2),.clk(gclk));
	jdff dff_B_FCpTu1Oa8_2(.din(w_dff_B_HHFWSoPB6_2),.dout(w_dff_B_FCpTu1Oa8_2),.clk(gclk));
	jdff dff_B_Xjo0NHRN6_2(.din(w_dff_B_FCpTu1Oa8_2),.dout(w_dff_B_Xjo0NHRN6_2),.clk(gclk));
	jdff dff_B_6gaVyu1c2_2(.din(w_dff_B_Xjo0NHRN6_2),.dout(w_dff_B_6gaVyu1c2_2),.clk(gclk));
	jdff dff_B_T9xSZq4u2_2(.din(w_dff_B_6gaVyu1c2_2),.dout(w_dff_B_T9xSZq4u2_2),.clk(gclk));
	jdff dff_B_rtoEWXzK4_1(.din(n1546),.dout(w_dff_B_rtoEWXzK4_1),.clk(gclk));
	jdff dff_B_gnbereKi1_2(.din(n1481),.dout(w_dff_B_gnbereKi1_2),.clk(gclk));
	jdff dff_B_4sCXKAMt1_2(.din(w_dff_B_gnbereKi1_2),.dout(w_dff_B_4sCXKAMt1_2),.clk(gclk));
	jdff dff_B_6isl9lQp4_2(.din(w_dff_B_4sCXKAMt1_2),.dout(w_dff_B_6isl9lQp4_2),.clk(gclk));
	jdff dff_B_Hdl40UF99_2(.din(w_dff_B_6isl9lQp4_2),.dout(w_dff_B_Hdl40UF99_2),.clk(gclk));
	jdff dff_B_k3FqWsEE3_2(.din(w_dff_B_Hdl40UF99_2),.dout(w_dff_B_k3FqWsEE3_2),.clk(gclk));
	jdff dff_B_iWKtQyWh8_2(.din(w_dff_B_k3FqWsEE3_2),.dout(w_dff_B_iWKtQyWh8_2),.clk(gclk));
	jdff dff_B_nvr54PpG3_2(.din(w_dff_B_iWKtQyWh8_2),.dout(w_dff_B_nvr54PpG3_2),.clk(gclk));
	jdff dff_B_AK8tEOvm0_2(.din(w_dff_B_nvr54PpG3_2),.dout(w_dff_B_AK8tEOvm0_2),.clk(gclk));
	jdff dff_B_1R9eaqrL3_2(.din(w_dff_B_AK8tEOvm0_2),.dout(w_dff_B_1R9eaqrL3_2),.clk(gclk));
	jdff dff_B_AtGAz6sJ3_2(.din(w_dff_B_1R9eaqrL3_2),.dout(w_dff_B_AtGAz6sJ3_2),.clk(gclk));
	jdff dff_B_bxWflXCE9_2(.din(w_dff_B_AtGAz6sJ3_2),.dout(w_dff_B_bxWflXCE9_2),.clk(gclk));
	jdff dff_B_SIXSQ67O1_2(.din(w_dff_B_bxWflXCE9_2),.dout(w_dff_B_SIXSQ67O1_2),.clk(gclk));
	jdff dff_B_7fkhM7wJ7_2(.din(w_dff_B_SIXSQ67O1_2),.dout(w_dff_B_7fkhM7wJ7_2),.clk(gclk));
	jdff dff_B_zYeiN5JJ3_2(.din(w_dff_B_7fkhM7wJ7_2),.dout(w_dff_B_zYeiN5JJ3_2),.clk(gclk));
	jdff dff_B_JMkfEVJD1_2(.din(w_dff_B_zYeiN5JJ3_2),.dout(w_dff_B_JMkfEVJD1_2),.clk(gclk));
	jdff dff_B_Tzx18ChG4_2(.din(w_dff_B_JMkfEVJD1_2),.dout(w_dff_B_Tzx18ChG4_2),.clk(gclk));
	jdff dff_B_yVYF2ret0_2(.din(w_dff_B_Tzx18ChG4_2),.dout(w_dff_B_yVYF2ret0_2),.clk(gclk));
	jdff dff_B_VbsMSVfW1_2(.din(w_dff_B_yVYF2ret0_2),.dout(w_dff_B_VbsMSVfW1_2),.clk(gclk));
	jdff dff_B_GRIBojrQ9_2(.din(w_dff_B_VbsMSVfW1_2),.dout(w_dff_B_GRIBojrQ9_2),.clk(gclk));
	jdff dff_B_ufNGh5Nz9_2(.din(w_dff_B_GRIBojrQ9_2),.dout(w_dff_B_ufNGh5Nz9_2),.clk(gclk));
	jdff dff_B_DDVDSGGr2_2(.din(w_dff_B_ufNGh5Nz9_2),.dout(w_dff_B_DDVDSGGr2_2),.clk(gclk));
	jdff dff_B_mNTMWGwj0_2(.din(w_dff_B_DDVDSGGr2_2),.dout(w_dff_B_mNTMWGwj0_2),.clk(gclk));
	jdff dff_B_VTye8jUV5_2(.din(w_dff_B_mNTMWGwj0_2),.dout(w_dff_B_VTye8jUV5_2),.clk(gclk));
	jdff dff_B_UOQW4Sx61_2(.din(w_dff_B_VTye8jUV5_2),.dout(w_dff_B_UOQW4Sx61_2),.clk(gclk));
	jdff dff_B_AXAewekX7_2(.din(w_dff_B_UOQW4Sx61_2),.dout(w_dff_B_AXAewekX7_2),.clk(gclk));
	jdff dff_B_I64BCFFe1_2(.din(w_dff_B_AXAewekX7_2),.dout(w_dff_B_I64BCFFe1_2),.clk(gclk));
	jdff dff_B_GV3oyR2n5_2(.din(w_dff_B_I64BCFFe1_2),.dout(w_dff_B_GV3oyR2n5_2),.clk(gclk));
	jdff dff_B_mjDJMCsb6_2(.din(w_dff_B_GV3oyR2n5_2),.dout(w_dff_B_mjDJMCsb6_2),.clk(gclk));
	jdff dff_B_8bAUqhY71_2(.din(w_dff_B_mjDJMCsb6_2),.dout(w_dff_B_8bAUqhY71_2),.clk(gclk));
	jdff dff_B_WnYZ6jln3_2(.din(w_dff_B_8bAUqhY71_2),.dout(w_dff_B_WnYZ6jln3_2),.clk(gclk));
	jdff dff_B_5mHy322U6_2(.din(w_dff_B_WnYZ6jln3_2),.dout(w_dff_B_5mHy322U6_2),.clk(gclk));
	jdff dff_B_w2IKrN7g5_2(.din(w_dff_B_5mHy322U6_2),.dout(w_dff_B_w2IKrN7g5_2),.clk(gclk));
	jdff dff_B_Qx7mxZdT6_2(.din(w_dff_B_w2IKrN7g5_2),.dout(w_dff_B_Qx7mxZdT6_2),.clk(gclk));
	jdff dff_B_V8sIV8sd4_2(.din(w_dff_B_Qx7mxZdT6_2),.dout(w_dff_B_V8sIV8sd4_2),.clk(gclk));
	jdff dff_B_YklFauZj3_2(.din(w_dff_B_V8sIV8sd4_2),.dout(w_dff_B_YklFauZj3_2),.clk(gclk));
	jdff dff_B_p7AWjSaB0_2(.din(n1513),.dout(w_dff_B_p7AWjSaB0_2),.clk(gclk));
	jdff dff_B_ISJUd31I5_1(.din(n1482),.dout(w_dff_B_ISJUd31I5_1),.clk(gclk));
	jdff dff_B_ojx5wQ788_2(.din(n1410),.dout(w_dff_B_ojx5wQ788_2),.clk(gclk));
	jdff dff_B_QrGb6vKY1_2(.din(w_dff_B_ojx5wQ788_2),.dout(w_dff_B_QrGb6vKY1_2),.clk(gclk));
	jdff dff_B_XmWNjiDD2_2(.din(w_dff_B_QrGb6vKY1_2),.dout(w_dff_B_XmWNjiDD2_2),.clk(gclk));
	jdff dff_B_U0fFuZLV2_2(.din(w_dff_B_XmWNjiDD2_2),.dout(w_dff_B_U0fFuZLV2_2),.clk(gclk));
	jdff dff_B_OcXYIF8E9_2(.din(w_dff_B_U0fFuZLV2_2),.dout(w_dff_B_OcXYIF8E9_2),.clk(gclk));
	jdff dff_B_gsfkJpD56_2(.din(w_dff_B_OcXYIF8E9_2),.dout(w_dff_B_gsfkJpD56_2),.clk(gclk));
	jdff dff_B_lX7IsoW62_2(.din(w_dff_B_gsfkJpD56_2),.dout(w_dff_B_lX7IsoW62_2),.clk(gclk));
	jdff dff_B_R6nnz4UU4_2(.din(w_dff_B_lX7IsoW62_2),.dout(w_dff_B_R6nnz4UU4_2),.clk(gclk));
	jdff dff_B_iseOWATe5_2(.din(w_dff_B_R6nnz4UU4_2),.dout(w_dff_B_iseOWATe5_2),.clk(gclk));
	jdff dff_B_ekQc6uMI0_2(.din(w_dff_B_iseOWATe5_2),.dout(w_dff_B_ekQc6uMI0_2),.clk(gclk));
	jdff dff_B_Tg2ton5F5_2(.din(w_dff_B_ekQc6uMI0_2),.dout(w_dff_B_Tg2ton5F5_2),.clk(gclk));
	jdff dff_B_NC6bMZWi2_2(.din(w_dff_B_Tg2ton5F5_2),.dout(w_dff_B_NC6bMZWi2_2),.clk(gclk));
	jdff dff_B_OV4Ev9ke2_2(.din(w_dff_B_NC6bMZWi2_2),.dout(w_dff_B_OV4Ev9ke2_2),.clk(gclk));
	jdff dff_B_is4k58l98_2(.din(w_dff_B_OV4Ev9ke2_2),.dout(w_dff_B_is4k58l98_2),.clk(gclk));
	jdff dff_B_lyz9BWDG1_2(.din(w_dff_B_is4k58l98_2),.dout(w_dff_B_lyz9BWDG1_2),.clk(gclk));
	jdff dff_B_guYPLWXn1_2(.din(w_dff_B_lyz9BWDG1_2),.dout(w_dff_B_guYPLWXn1_2),.clk(gclk));
	jdff dff_B_mCemIItI9_2(.din(w_dff_B_guYPLWXn1_2),.dout(w_dff_B_mCemIItI9_2),.clk(gclk));
	jdff dff_B_TqwFgypW8_2(.din(w_dff_B_mCemIItI9_2),.dout(w_dff_B_TqwFgypW8_2),.clk(gclk));
	jdff dff_B_xYAQw4AV9_2(.din(w_dff_B_TqwFgypW8_2),.dout(w_dff_B_xYAQw4AV9_2),.clk(gclk));
	jdff dff_B_EdqLmb3R3_2(.din(w_dff_B_xYAQw4AV9_2),.dout(w_dff_B_EdqLmb3R3_2),.clk(gclk));
	jdff dff_B_wCYtV0fA5_2(.din(w_dff_B_EdqLmb3R3_2),.dout(w_dff_B_wCYtV0fA5_2),.clk(gclk));
	jdff dff_B_C2u7cuHN4_2(.din(w_dff_B_wCYtV0fA5_2),.dout(w_dff_B_C2u7cuHN4_2),.clk(gclk));
	jdff dff_B_57zDsbaF2_2(.din(w_dff_B_C2u7cuHN4_2),.dout(w_dff_B_57zDsbaF2_2),.clk(gclk));
	jdff dff_B_jHyEaw602_2(.din(w_dff_B_57zDsbaF2_2),.dout(w_dff_B_jHyEaw602_2),.clk(gclk));
	jdff dff_B_EGWOWf9O9_2(.din(w_dff_B_jHyEaw602_2),.dout(w_dff_B_EGWOWf9O9_2),.clk(gclk));
	jdff dff_B_3Q829Jkz3_2(.din(w_dff_B_EGWOWf9O9_2),.dout(w_dff_B_3Q829Jkz3_2),.clk(gclk));
	jdff dff_B_sJTrjs2W8_2(.din(w_dff_B_3Q829Jkz3_2),.dout(w_dff_B_sJTrjs2W8_2),.clk(gclk));
	jdff dff_B_tCRWd8Nn7_2(.din(w_dff_B_sJTrjs2W8_2),.dout(w_dff_B_tCRWd8Nn7_2),.clk(gclk));
	jdff dff_B_lgAIjsaz4_2(.din(w_dff_B_tCRWd8Nn7_2),.dout(w_dff_B_lgAIjsaz4_2),.clk(gclk));
	jdff dff_B_gFPDvHSl5_2(.din(w_dff_B_lgAIjsaz4_2),.dout(w_dff_B_gFPDvHSl5_2),.clk(gclk));
	jdff dff_B_XWMtnGVA1_2(.din(w_dff_B_gFPDvHSl5_2),.dout(w_dff_B_XWMtnGVA1_2),.clk(gclk));
	jdff dff_B_b6jgOv2c9_2(.din(w_dff_B_XWMtnGVA1_2),.dout(w_dff_B_b6jgOv2c9_2),.clk(gclk));
	jdff dff_B_OMXvXjla2_2(.din(n1442),.dout(w_dff_B_OMXvXjla2_2),.clk(gclk));
	jdff dff_B_Np1v8xsj0_1(.din(n1411),.dout(w_dff_B_Np1v8xsj0_1),.clk(gclk));
	jdff dff_B_r9gpkzOX2_2(.din(n1332),.dout(w_dff_B_r9gpkzOX2_2),.clk(gclk));
	jdff dff_B_Q5FUyK8T8_2(.din(w_dff_B_r9gpkzOX2_2),.dout(w_dff_B_Q5FUyK8T8_2),.clk(gclk));
	jdff dff_B_WR9kmS2X1_2(.din(w_dff_B_Q5FUyK8T8_2),.dout(w_dff_B_WR9kmS2X1_2),.clk(gclk));
	jdff dff_B_1DoWVFXC1_2(.din(w_dff_B_WR9kmS2X1_2),.dout(w_dff_B_1DoWVFXC1_2),.clk(gclk));
	jdff dff_B_ZAbB7ElF1_2(.din(w_dff_B_1DoWVFXC1_2),.dout(w_dff_B_ZAbB7ElF1_2),.clk(gclk));
	jdff dff_B_DPWgG65B2_2(.din(w_dff_B_ZAbB7ElF1_2),.dout(w_dff_B_DPWgG65B2_2),.clk(gclk));
	jdff dff_B_d4tDt8xY2_2(.din(w_dff_B_DPWgG65B2_2),.dout(w_dff_B_d4tDt8xY2_2),.clk(gclk));
	jdff dff_B_SE9M4N407_2(.din(w_dff_B_d4tDt8xY2_2),.dout(w_dff_B_SE9M4N407_2),.clk(gclk));
	jdff dff_B_4KpCWajW6_2(.din(w_dff_B_SE9M4N407_2),.dout(w_dff_B_4KpCWajW6_2),.clk(gclk));
	jdff dff_B_7rAnPWkD7_2(.din(w_dff_B_4KpCWajW6_2),.dout(w_dff_B_7rAnPWkD7_2),.clk(gclk));
	jdff dff_B_OAgzgMeN7_2(.din(w_dff_B_7rAnPWkD7_2),.dout(w_dff_B_OAgzgMeN7_2),.clk(gclk));
	jdff dff_B_f3bO6ym16_2(.din(w_dff_B_OAgzgMeN7_2),.dout(w_dff_B_f3bO6ym16_2),.clk(gclk));
	jdff dff_B_HesHG1wa0_2(.din(w_dff_B_f3bO6ym16_2),.dout(w_dff_B_HesHG1wa0_2),.clk(gclk));
	jdff dff_B_n536rLtD1_2(.din(w_dff_B_HesHG1wa0_2),.dout(w_dff_B_n536rLtD1_2),.clk(gclk));
	jdff dff_B_6lxU23xG7_2(.din(w_dff_B_n536rLtD1_2),.dout(w_dff_B_6lxU23xG7_2),.clk(gclk));
	jdff dff_B_oK34vapg7_2(.din(w_dff_B_6lxU23xG7_2),.dout(w_dff_B_oK34vapg7_2),.clk(gclk));
	jdff dff_B_RIE4rCTD5_2(.din(w_dff_B_oK34vapg7_2),.dout(w_dff_B_RIE4rCTD5_2),.clk(gclk));
	jdff dff_B_tP5Jx9bR0_2(.din(w_dff_B_RIE4rCTD5_2),.dout(w_dff_B_tP5Jx9bR0_2),.clk(gclk));
	jdff dff_B_jY14pEFG1_2(.din(w_dff_B_tP5Jx9bR0_2),.dout(w_dff_B_jY14pEFG1_2),.clk(gclk));
	jdff dff_B_MnnwXFB70_2(.din(w_dff_B_jY14pEFG1_2),.dout(w_dff_B_MnnwXFB70_2),.clk(gclk));
	jdff dff_B_3EnhQxlt8_2(.din(w_dff_B_MnnwXFB70_2),.dout(w_dff_B_3EnhQxlt8_2),.clk(gclk));
	jdff dff_B_exRvzMEK2_2(.din(w_dff_B_3EnhQxlt8_2),.dout(w_dff_B_exRvzMEK2_2),.clk(gclk));
	jdff dff_B_yAKnvj3u6_2(.din(w_dff_B_exRvzMEK2_2),.dout(w_dff_B_yAKnvj3u6_2),.clk(gclk));
	jdff dff_B_j4vFqJ064_2(.din(w_dff_B_yAKnvj3u6_2),.dout(w_dff_B_j4vFqJ064_2),.clk(gclk));
	jdff dff_B_yJX6VZx83_2(.din(w_dff_B_j4vFqJ064_2),.dout(w_dff_B_yJX6VZx83_2),.clk(gclk));
	jdff dff_B_GWUwXBzq6_2(.din(w_dff_B_yJX6VZx83_2),.dout(w_dff_B_GWUwXBzq6_2),.clk(gclk));
	jdff dff_B_YFRCnf3a8_2(.din(w_dff_B_GWUwXBzq6_2),.dout(w_dff_B_YFRCnf3a8_2),.clk(gclk));
	jdff dff_B_8IqsvRsL8_2(.din(w_dff_B_YFRCnf3a8_2),.dout(w_dff_B_8IqsvRsL8_2),.clk(gclk));
	jdff dff_B_FIqkKil95_2(.din(w_dff_B_8IqsvRsL8_2),.dout(w_dff_B_FIqkKil95_2),.clk(gclk));
	jdff dff_B_QCqWFUuj5_2(.din(n1364),.dout(w_dff_B_QCqWFUuj5_2),.clk(gclk));
	jdff dff_B_sVmjXq6O1_1(.din(n1333),.dout(w_dff_B_sVmjXq6O1_1),.clk(gclk));
	jdff dff_B_EEabGscb2_2(.din(n1247),.dout(w_dff_B_EEabGscb2_2),.clk(gclk));
	jdff dff_B_C5w2kazg8_2(.din(w_dff_B_EEabGscb2_2),.dout(w_dff_B_C5w2kazg8_2),.clk(gclk));
	jdff dff_B_r9Sv5kHl7_2(.din(w_dff_B_C5w2kazg8_2),.dout(w_dff_B_r9Sv5kHl7_2),.clk(gclk));
	jdff dff_B_uGOE5r0T1_2(.din(w_dff_B_r9Sv5kHl7_2),.dout(w_dff_B_uGOE5r0T1_2),.clk(gclk));
	jdff dff_B_9TwJOURK2_2(.din(w_dff_B_uGOE5r0T1_2),.dout(w_dff_B_9TwJOURK2_2),.clk(gclk));
	jdff dff_B_TfOF2y5w2_2(.din(w_dff_B_9TwJOURK2_2),.dout(w_dff_B_TfOF2y5w2_2),.clk(gclk));
	jdff dff_B_6IR98p932_2(.din(w_dff_B_TfOF2y5w2_2),.dout(w_dff_B_6IR98p932_2),.clk(gclk));
	jdff dff_B_btSoseQP4_2(.din(w_dff_B_6IR98p932_2),.dout(w_dff_B_btSoseQP4_2),.clk(gclk));
	jdff dff_B_fS0yraMI8_2(.din(w_dff_B_btSoseQP4_2),.dout(w_dff_B_fS0yraMI8_2),.clk(gclk));
	jdff dff_B_scyRMOS63_2(.din(w_dff_B_fS0yraMI8_2),.dout(w_dff_B_scyRMOS63_2),.clk(gclk));
	jdff dff_B_pVniVI5P7_2(.din(w_dff_B_scyRMOS63_2),.dout(w_dff_B_pVniVI5P7_2),.clk(gclk));
	jdff dff_B_9uNclzfI9_2(.din(w_dff_B_pVniVI5P7_2),.dout(w_dff_B_9uNclzfI9_2),.clk(gclk));
	jdff dff_B_c3VBUoBz3_2(.din(w_dff_B_9uNclzfI9_2),.dout(w_dff_B_c3VBUoBz3_2),.clk(gclk));
	jdff dff_B_4ifoD7h11_2(.din(w_dff_B_c3VBUoBz3_2),.dout(w_dff_B_4ifoD7h11_2),.clk(gclk));
	jdff dff_B_hlolFbYN3_2(.din(w_dff_B_4ifoD7h11_2),.dout(w_dff_B_hlolFbYN3_2),.clk(gclk));
	jdff dff_B_GcVyUEG90_2(.din(w_dff_B_hlolFbYN3_2),.dout(w_dff_B_GcVyUEG90_2),.clk(gclk));
	jdff dff_B_IVrARRAJ7_2(.din(w_dff_B_GcVyUEG90_2),.dout(w_dff_B_IVrARRAJ7_2),.clk(gclk));
	jdff dff_B_7JJpx3z64_2(.din(w_dff_B_IVrARRAJ7_2),.dout(w_dff_B_7JJpx3z64_2),.clk(gclk));
	jdff dff_B_Jewm9tFG1_2(.din(w_dff_B_7JJpx3z64_2),.dout(w_dff_B_Jewm9tFG1_2),.clk(gclk));
	jdff dff_B_p9A0L6m08_2(.din(w_dff_B_Jewm9tFG1_2),.dout(w_dff_B_p9A0L6m08_2),.clk(gclk));
	jdff dff_B_lHK1nEr31_2(.din(w_dff_B_p9A0L6m08_2),.dout(w_dff_B_lHK1nEr31_2),.clk(gclk));
	jdff dff_B_xgDKfvmL6_2(.din(w_dff_B_lHK1nEr31_2),.dout(w_dff_B_xgDKfvmL6_2),.clk(gclk));
	jdff dff_B_9SBAGRw60_2(.din(w_dff_B_xgDKfvmL6_2),.dout(w_dff_B_9SBAGRw60_2),.clk(gclk));
	jdff dff_B_77LkU9Lp6_2(.din(w_dff_B_9SBAGRw60_2),.dout(w_dff_B_77LkU9Lp6_2),.clk(gclk));
	jdff dff_B_oo3hJmBa6_2(.din(w_dff_B_77LkU9Lp6_2),.dout(w_dff_B_oo3hJmBa6_2),.clk(gclk));
	jdff dff_B_lI9bCXDS3_2(.din(w_dff_B_oo3hJmBa6_2),.dout(w_dff_B_lI9bCXDS3_2),.clk(gclk));
	jdff dff_B_vcCq38sD8_2(.din(n1279),.dout(w_dff_B_vcCq38sD8_2),.clk(gclk));
	jdff dff_B_D0MLO62s7_1(.din(n1248),.dout(w_dff_B_D0MLO62s7_1),.clk(gclk));
	jdff dff_B_lDD5EwiP7_2(.din(n1156),.dout(w_dff_B_lDD5EwiP7_2),.clk(gclk));
	jdff dff_B_Hdwz1ovf6_2(.din(w_dff_B_lDD5EwiP7_2),.dout(w_dff_B_Hdwz1ovf6_2),.clk(gclk));
	jdff dff_B_jqabLlTY0_2(.din(w_dff_B_Hdwz1ovf6_2),.dout(w_dff_B_jqabLlTY0_2),.clk(gclk));
	jdff dff_B_uKePzSI57_2(.din(w_dff_B_jqabLlTY0_2),.dout(w_dff_B_uKePzSI57_2),.clk(gclk));
	jdff dff_B_gaOYESsH8_2(.din(w_dff_B_uKePzSI57_2),.dout(w_dff_B_gaOYESsH8_2),.clk(gclk));
	jdff dff_B_CniT0wFX8_2(.din(w_dff_B_gaOYESsH8_2),.dout(w_dff_B_CniT0wFX8_2),.clk(gclk));
	jdff dff_B_dHg9dOE06_2(.din(w_dff_B_CniT0wFX8_2),.dout(w_dff_B_dHg9dOE06_2),.clk(gclk));
	jdff dff_B_NIVvBHeG0_2(.din(w_dff_B_dHg9dOE06_2),.dout(w_dff_B_NIVvBHeG0_2),.clk(gclk));
	jdff dff_B_VzNCio8K6_2(.din(w_dff_B_NIVvBHeG0_2),.dout(w_dff_B_VzNCio8K6_2),.clk(gclk));
	jdff dff_B_8w6j5v7y6_2(.din(w_dff_B_VzNCio8K6_2),.dout(w_dff_B_8w6j5v7y6_2),.clk(gclk));
	jdff dff_B_pcyUuP953_2(.din(w_dff_B_8w6j5v7y6_2),.dout(w_dff_B_pcyUuP953_2),.clk(gclk));
	jdff dff_B_0Hiugs2T1_2(.din(w_dff_B_pcyUuP953_2),.dout(w_dff_B_0Hiugs2T1_2),.clk(gclk));
	jdff dff_B_BAdALqCA6_2(.din(w_dff_B_0Hiugs2T1_2),.dout(w_dff_B_BAdALqCA6_2),.clk(gclk));
	jdff dff_B_mSwIxkXj7_2(.din(w_dff_B_BAdALqCA6_2),.dout(w_dff_B_mSwIxkXj7_2),.clk(gclk));
	jdff dff_B_T0QRnaFX5_2(.din(w_dff_B_mSwIxkXj7_2),.dout(w_dff_B_T0QRnaFX5_2),.clk(gclk));
	jdff dff_B_GNuTaNYm0_2(.din(w_dff_B_T0QRnaFX5_2),.dout(w_dff_B_GNuTaNYm0_2),.clk(gclk));
	jdff dff_B_Dy29BoGg8_2(.din(w_dff_B_GNuTaNYm0_2),.dout(w_dff_B_Dy29BoGg8_2),.clk(gclk));
	jdff dff_B_tSwhzLp33_2(.din(w_dff_B_Dy29BoGg8_2),.dout(w_dff_B_tSwhzLp33_2),.clk(gclk));
	jdff dff_B_gGSt85UG0_2(.din(w_dff_B_tSwhzLp33_2),.dout(w_dff_B_gGSt85UG0_2),.clk(gclk));
	jdff dff_B_YYxGgZYu9_2(.din(w_dff_B_gGSt85UG0_2),.dout(w_dff_B_YYxGgZYu9_2),.clk(gclk));
	jdff dff_B_d5I3Ey5t8_2(.din(w_dff_B_YYxGgZYu9_2),.dout(w_dff_B_d5I3Ey5t8_2),.clk(gclk));
	jdff dff_B_QuqzS3fK1_2(.din(w_dff_B_d5I3Ey5t8_2),.dout(w_dff_B_QuqzS3fK1_2),.clk(gclk));
	jdff dff_B_mNza9tcW4_2(.din(w_dff_B_QuqzS3fK1_2),.dout(w_dff_B_mNza9tcW4_2),.clk(gclk));
	jdff dff_B_WUYVu1hl2_2(.din(n1188),.dout(w_dff_B_WUYVu1hl2_2),.clk(gclk));
	jdff dff_B_QMF8uRl06_1(.din(n1157),.dout(w_dff_B_QMF8uRl06_1),.clk(gclk));
	jdff dff_B_GWeOCnPO4_2(.din(n1058),.dout(w_dff_B_GWeOCnPO4_2),.clk(gclk));
	jdff dff_B_dp9fFCs86_2(.din(w_dff_B_GWeOCnPO4_2),.dout(w_dff_B_dp9fFCs86_2),.clk(gclk));
	jdff dff_B_VCj82tDn3_2(.din(w_dff_B_dp9fFCs86_2),.dout(w_dff_B_VCj82tDn3_2),.clk(gclk));
	jdff dff_B_vR181oxi7_2(.din(w_dff_B_VCj82tDn3_2),.dout(w_dff_B_vR181oxi7_2),.clk(gclk));
	jdff dff_B_IxfaIcaT8_2(.din(w_dff_B_vR181oxi7_2),.dout(w_dff_B_IxfaIcaT8_2),.clk(gclk));
	jdff dff_B_IztkZPXG7_2(.din(w_dff_B_IxfaIcaT8_2),.dout(w_dff_B_IztkZPXG7_2),.clk(gclk));
	jdff dff_B_hrt4Mc5x8_2(.din(w_dff_B_IztkZPXG7_2),.dout(w_dff_B_hrt4Mc5x8_2),.clk(gclk));
	jdff dff_B_8G0zxng01_2(.din(w_dff_B_hrt4Mc5x8_2),.dout(w_dff_B_8G0zxng01_2),.clk(gclk));
	jdff dff_B_iSS9SgOM1_2(.din(w_dff_B_8G0zxng01_2),.dout(w_dff_B_iSS9SgOM1_2),.clk(gclk));
	jdff dff_B_61yb0ejX0_2(.din(w_dff_B_iSS9SgOM1_2),.dout(w_dff_B_61yb0ejX0_2),.clk(gclk));
	jdff dff_B_DyhUzHgK1_2(.din(w_dff_B_61yb0ejX0_2),.dout(w_dff_B_DyhUzHgK1_2),.clk(gclk));
	jdff dff_B_Q1Z70QoM6_2(.din(w_dff_B_DyhUzHgK1_2),.dout(w_dff_B_Q1Z70QoM6_2),.clk(gclk));
	jdff dff_B_rKgbTX9Z3_2(.din(w_dff_B_Q1Z70QoM6_2),.dout(w_dff_B_rKgbTX9Z3_2),.clk(gclk));
	jdff dff_B_ZyRBvNaZ5_2(.din(w_dff_B_rKgbTX9Z3_2),.dout(w_dff_B_ZyRBvNaZ5_2),.clk(gclk));
	jdff dff_B_JiEXtOrC9_2(.din(w_dff_B_ZyRBvNaZ5_2),.dout(w_dff_B_JiEXtOrC9_2),.clk(gclk));
	jdff dff_B_Ac5JdQf82_2(.din(w_dff_B_JiEXtOrC9_2),.dout(w_dff_B_Ac5JdQf82_2),.clk(gclk));
	jdff dff_B_QPIfgRm07_2(.din(w_dff_B_Ac5JdQf82_2),.dout(w_dff_B_QPIfgRm07_2),.clk(gclk));
	jdff dff_B_dvVVJkmv8_2(.din(w_dff_B_QPIfgRm07_2),.dout(w_dff_B_dvVVJkmv8_2),.clk(gclk));
	jdff dff_B_9c7T0okH9_2(.din(w_dff_B_dvVVJkmv8_2),.dout(w_dff_B_9c7T0okH9_2),.clk(gclk));
	jdff dff_B_652yf0Nx1_2(.din(w_dff_B_9c7T0okH9_2),.dout(w_dff_B_652yf0Nx1_2),.clk(gclk));
	jdff dff_B_NeEOwLOI0_2(.din(n1089),.dout(w_dff_B_NeEOwLOI0_2),.clk(gclk));
	jdff dff_B_Fipv8Gnp4_1(.din(n1059),.dout(w_dff_B_Fipv8Gnp4_1),.clk(gclk));
	jdff dff_B_D7jdRNo73_2(.din(n959),.dout(w_dff_B_D7jdRNo73_2),.clk(gclk));
	jdff dff_B_BtA0HKAD4_2(.din(w_dff_B_D7jdRNo73_2),.dout(w_dff_B_BtA0HKAD4_2),.clk(gclk));
	jdff dff_B_AhycjzWL7_2(.din(w_dff_B_BtA0HKAD4_2),.dout(w_dff_B_AhycjzWL7_2),.clk(gclk));
	jdff dff_B_3xKiqqXz9_2(.din(w_dff_B_AhycjzWL7_2),.dout(w_dff_B_3xKiqqXz9_2),.clk(gclk));
	jdff dff_B_T7FWyf9u6_2(.din(w_dff_B_3xKiqqXz9_2),.dout(w_dff_B_T7FWyf9u6_2),.clk(gclk));
	jdff dff_B_OU22KPS90_2(.din(w_dff_B_T7FWyf9u6_2),.dout(w_dff_B_OU22KPS90_2),.clk(gclk));
	jdff dff_B_RjM9ejhg4_2(.din(w_dff_B_OU22KPS90_2),.dout(w_dff_B_RjM9ejhg4_2),.clk(gclk));
	jdff dff_B_gab97HyR4_2(.din(w_dff_B_RjM9ejhg4_2),.dout(w_dff_B_gab97HyR4_2),.clk(gclk));
	jdff dff_B_rMKqRuTO1_2(.din(w_dff_B_gab97HyR4_2),.dout(w_dff_B_rMKqRuTO1_2),.clk(gclk));
	jdff dff_B_dSkZkfJE4_2(.din(w_dff_B_rMKqRuTO1_2),.dout(w_dff_B_dSkZkfJE4_2),.clk(gclk));
	jdff dff_B_sN3aDqCS2_2(.din(w_dff_B_dSkZkfJE4_2),.dout(w_dff_B_sN3aDqCS2_2),.clk(gclk));
	jdff dff_B_ncNNF4w89_2(.din(w_dff_B_sN3aDqCS2_2),.dout(w_dff_B_ncNNF4w89_2),.clk(gclk));
	jdff dff_B_mNnMG2Nw2_2(.din(w_dff_B_ncNNF4w89_2),.dout(w_dff_B_mNnMG2Nw2_2),.clk(gclk));
	jdff dff_B_Nu24rtER5_2(.din(w_dff_B_mNnMG2Nw2_2),.dout(w_dff_B_Nu24rtER5_2),.clk(gclk));
	jdff dff_B_EH87Q9Ja2_2(.din(w_dff_B_Nu24rtER5_2),.dout(w_dff_B_EH87Q9Ja2_2),.clk(gclk));
	jdff dff_B_v7n9ZdN78_2(.din(w_dff_B_EH87Q9Ja2_2),.dout(w_dff_B_v7n9ZdN78_2),.clk(gclk));
	jdff dff_B_vel3G9qh4_2(.din(w_dff_B_v7n9ZdN78_2),.dout(w_dff_B_vel3G9qh4_2),.clk(gclk));
	jdff dff_B_BygthE7M4_2(.din(n990),.dout(w_dff_B_BygthE7M4_2),.clk(gclk));
	jdff dff_B_8eTRNjEg9_1(.din(n960),.dout(w_dff_B_8eTRNjEg9_1),.clk(gclk));
	jdff dff_B_dSdzBKzL6_2(.din(n857),.dout(w_dff_B_dSdzBKzL6_2),.clk(gclk));
	jdff dff_B_kRD1cGHm0_2(.din(w_dff_B_dSdzBKzL6_2),.dout(w_dff_B_kRD1cGHm0_2),.clk(gclk));
	jdff dff_B_XSB0ImkT2_2(.din(w_dff_B_kRD1cGHm0_2),.dout(w_dff_B_XSB0ImkT2_2),.clk(gclk));
	jdff dff_B_XFmF0o247_2(.din(w_dff_B_XSB0ImkT2_2),.dout(w_dff_B_XFmF0o247_2),.clk(gclk));
	jdff dff_B_PD1NDFcd8_2(.din(w_dff_B_XFmF0o247_2),.dout(w_dff_B_PD1NDFcd8_2),.clk(gclk));
	jdff dff_B_NB5zcMHp8_2(.din(w_dff_B_PD1NDFcd8_2),.dout(w_dff_B_NB5zcMHp8_2),.clk(gclk));
	jdff dff_B_LoTM9iGp8_2(.din(w_dff_B_NB5zcMHp8_2),.dout(w_dff_B_LoTM9iGp8_2),.clk(gclk));
	jdff dff_B_vh1z7EQf4_2(.din(w_dff_B_LoTM9iGp8_2),.dout(w_dff_B_vh1z7EQf4_2),.clk(gclk));
	jdff dff_B_zQxCkmZz4_2(.din(w_dff_B_vh1z7EQf4_2),.dout(w_dff_B_zQxCkmZz4_2),.clk(gclk));
	jdff dff_B_f8lY0Vet6_2(.din(w_dff_B_zQxCkmZz4_2),.dout(w_dff_B_f8lY0Vet6_2),.clk(gclk));
	jdff dff_B_dx4pguYu7_2(.din(w_dff_B_f8lY0Vet6_2),.dout(w_dff_B_dx4pguYu7_2),.clk(gclk));
	jdff dff_B_QmuKa4eK6_2(.din(w_dff_B_dx4pguYu7_2),.dout(w_dff_B_QmuKa4eK6_2),.clk(gclk));
	jdff dff_B_7X7O8SjT0_2(.din(w_dff_B_QmuKa4eK6_2),.dout(w_dff_B_7X7O8SjT0_2),.clk(gclk));
	jdff dff_B_y521lsx49_2(.din(w_dff_B_7X7O8SjT0_2),.dout(w_dff_B_y521lsx49_2),.clk(gclk));
	jdff dff_B_nNHk4TPi9_2(.din(n884),.dout(w_dff_B_nNHk4TPi9_2),.clk(gclk));
	jdff dff_B_ls7eEVDF7_1(.din(n858),.dout(w_dff_B_ls7eEVDF7_1),.clk(gclk));
	jdff dff_B_zKkPmLf05_2(.din(n759),.dout(w_dff_B_zKkPmLf05_2),.clk(gclk));
	jdff dff_B_TqMtYgbm1_2(.din(w_dff_B_zKkPmLf05_2),.dout(w_dff_B_TqMtYgbm1_2),.clk(gclk));
	jdff dff_B_jE18dZpw0_2(.din(w_dff_B_TqMtYgbm1_2),.dout(w_dff_B_jE18dZpw0_2),.clk(gclk));
	jdff dff_B_DJpvfd7x3_2(.din(w_dff_B_jE18dZpw0_2),.dout(w_dff_B_DJpvfd7x3_2),.clk(gclk));
	jdff dff_B_RhTWUUQC2_2(.din(w_dff_B_DJpvfd7x3_2),.dout(w_dff_B_RhTWUUQC2_2),.clk(gclk));
	jdff dff_B_lUQaqNA31_2(.din(w_dff_B_RhTWUUQC2_2),.dout(w_dff_B_lUQaqNA31_2),.clk(gclk));
	jdff dff_B_jhO1V4YD3_2(.din(w_dff_B_lUQaqNA31_2),.dout(w_dff_B_jhO1V4YD3_2),.clk(gclk));
	jdff dff_B_OmTWrffi8_2(.din(w_dff_B_jhO1V4YD3_2),.dout(w_dff_B_OmTWrffi8_2),.clk(gclk));
	jdff dff_B_6XF6CHzP5_2(.din(w_dff_B_OmTWrffi8_2),.dout(w_dff_B_6XF6CHzP5_2),.clk(gclk));
	jdff dff_B_AZbtr5c57_2(.din(w_dff_B_6XF6CHzP5_2),.dout(w_dff_B_AZbtr5c57_2),.clk(gclk));
	jdff dff_B_L4nzzlCr2_2(.din(w_dff_B_AZbtr5c57_2),.dout(w_dff_B_L4nzzlCr2_2),.clk(gclk));
	jdff dff_B_t4bNrN1L3_2(.din(n781),.dout(w_dff_B_t4bNrN1L3_2),.clk(gclk));
	jdff dff_B_MeaEWRaU7_1(.din(n760),.dout(w_dff_B_MeaEWRaU7_1),.clk(gclk));
	jdff dff_B_BHp6WDKG1_2(.din(n667),.dout(w_dff_B_BHp6WDKG1_2),.clk(gclk));
	jdff dff_B_DSmInTRM0_2(.din(w_dff_B_BHp6WDKG1_2),.dout(w_dff_B_DSmInTRM0_2),.clk(gclk));
	jdff dff_B_3QYMA24v9_2(.din(w_dff_B_DSmInTRM0_2),.dout(w_dff_B_3QYMA24v9_2),.clk(gclk));
	jdff dff_B_SFGCOXC16_2(.din(w_dff_B_3QYMA24v9_2),.dout(w_dff_B_SFGCOXC16_2),.clk(gclk));
	jdff dff_B_PjFtCOgg4_2(.din(w_dff_B_SFGCOXC16_2),.dout(w_dff_B_PjFtCOgg4_2),.clk(gclk));
	jdff dff_B_gWzcO45F1_2(.din(w_dff_B_PjFtCOgg4_2),.dout(w_dff_B_gWzcO45F1_2),.clk(gclk));
	jdff dff_B_e3dMIBCj6_2(.din(w_dff_B_gWzcO45F1_2),.dout(w_dff_B_e3dMIBCj6_2),.clk(gclk));
	jdff dff_B_KiS2yLUk1_2(.din(w_dff_B_e3dMIBCj6_2),.dout(w_dff_B_KiS2yLUk1_2),.clk(gclk));
	jdff dff_B_5fbQ0Tdx8_2(.din(n682),.dout(w_dff_B_5fbQ0Tdx8_2),.clk(gclk));
	jdff dff_B_FXkMh77Y8_2(.din(w_dff_B_5fbQ0Tdx8_2),.dout(w_dff_B_FXkMh77Y8_2),.clk(gclk));
	jdff dff_B_BJLQn1AZ7_2(.din(w_dff_B_FXkMh77Y8_2),.dout(w_dff_B_BJLQn1AZ7_2),.clk(gclk));
	jdff dff_B_HdovCmk45_1(.din(n668),.dout(w_dff_B_HdovCmk45_1),.clk(gclk));
	jdff dff_B_Q8Jhx20V3_1(.din(w_dff_B_HdovCmk45_1),.dout(w_dff_B_Q8Jhx20V3_1),.clk(gclk));
	jdff dff_B_uImFXF9W3_2(.din(n584),.dout(w_dff_B_uImFXF9W3_2),.clk(gclk));
	jdff dff_B_Mzhg2ssD0_2(.din(w_dff_B_uImFXF9W3_2),.dout(w_dff_B_Mzhg2ssD0_2),.clk(gclk));
	jdff dff_B_ts3WuSzZ2_2(.din(w_dff_B_Mzhg2ssD0_2),.dout(w_dff_B_ts3WuSzZ2_2),.clk(gclk));
	jdff dff_B_vPj7a03l5_0(.din(n589),.dout(w_dff_B_vPj7a03l5_0),.clk(gclk));
	jdff dff_A_KX7Rd5572_0(.dout(w_n503_0[0]),.din(w_dff_A_KX7Rd5572_0),.clk(gclk));
	jdff dff_A_rWc83jMO0_0(.dout(w_dff_A_KX7Rd5572_0),.din(w_dff_A_rWc83jMO0_0),.clk(gclk));
	jdff dff_A_gy46G8l43_1(.dout(w_n503_0[1]),.din(w_dff_A_gy46G8l43_1),.clk(gclk));
	jdff dff_A_mOLit72c0_1(.dout(w_dff_A_gy46G8l43_1),.din(w_dff_A_mOLit72c0_1),.clk(gclk));
	jdff dff_B_s9lPq6nu2_1(.din(n1762),.dout(w_dff_B_s9lPq6nu2_1),.clk(gclk));
	jdff dff_A_xWpozIyr6_1(.dout(w_n1737_0[1]),.din(w_dff_A_xWpozIyr6_1),.clk(gclk));
	jdff dff_B_iOR8SBie2_1(.din(n1735),.dout(w_dff_B_iOR8SBie2_1),.clk(gclk));
	jdff dff_B_xvidG6BS0_2(.din(n1699),.dout(w_dff_B_xvidG6BS0_2),.clk(gclk));
	jdff dff_B_H2JOajln6_2(.din(w_dff_B_xvidG6BS0_2),.dout(w_dff_B_H2JOajln6_2),.clk(gclk));
	jdff dff_B_Ycn68z6x2_2(.din(w_dff_B_H2JOajln6_2),.dout(w_dff_B_Ycn68z6x2_2),.clk(gclk));
	jdff dff_B_Qkicp0Nj0_2(.din(w_dff_B_Ycn68z6x2_2),.dout(w_dff_B_Qkicp0Nj0_2),.clk(gclk));
	jdff dff_B_zlxqnU5T9_2(.din(w_dff_B_Qkicp0Nj0_2),.dout(w_dff_B_zlxqnU5T9_2),.clk(gclk));
	jdff dff_B_mSDuYZpA9_2(.din(w_dff_B_zlxqnU5T9_2),.dout(w_dff_B_mSDuYZpA9_2),.clk(gclk));
	jdff dff_B_vmDLUHHK1_2(.din(w_dff_B_mSDuYZpA9_2),.dout(w_dff_B_vmDLUHHK1_2),.clk(gclk));
	jdff dff_B_eHd2FTqC3_2(.din(w_dff_B_vmDLUHHK1_2),.dout(w_dff_B_eHd2FTqC3_2),.clk(gclk));
	jdff dff_B_uBOGlqrS6_2(.din(w_dff_B_eHd2FTqC3_2),.dout(w_dff_B_uBOGlqrS6_2),.clk(gclk));
	jdff dff_B_gyLmnItY4_2(.din(w_dff_B_uBOGlqrS6_2),.dout(w_dff_B_gyLmnItY4_2),.clk(gclk));
	jdff dff_B_A0NbFXRA3_2(.din(w_dff_B_gyLmnItY4_2),.dout(w_dff_B_A0NbFXRA3_2),.clk(gclk));
	jdff dff_B_KZ3Pl0a95_2(.din(w_dff_B_A0NbFXRA3_2),.dout(w_dff_B_KZ3Pl0a95_2),.clk(gclk));
	jdff dff_B_68pFLTaF9_2(.din(w_dff_B_KZ3Pl0a95_2),.dout(w_dff_B_68pFLTaF9_2),.clk(gclk));
	jdff dff_B_Nblkd6oV4_2(.din(w_dff_B_68pFLTaF9_2),.dout(w_dff_B_Nblkd6oV4_2),.clk(gclk));
	jdff dff_B_msA6pmMP5_2(.din(w_dff_B_Nblkd6oV4_2),.dout(w_dff_B_msA6pmMP5_2),.clk(gclk));
	jdff dff_B_OTPIfpTj9_2(.din(w_dff_B_msA6pmMP5_2),.dout(w_dff_B_OTPIfpTj9_2),.clk(gclk));
	jdff dff_B_ThheJh362_2(.din(w_dff_B_OTPIfpTj9_2),.dout(w_dff_B_ThheJh362_2),.clk(gclk));
	jdff dff_B_78wLyOoW3_2(.din(w_dff_B_ThheJh362_2),.dout(w_dff_B_78wLyOoW3_2),.clk(gclk));
	jdff dff_B_K1WphjVx7_2(.din(w_dff_B_78wLyOoW3_2),.dout(w_dff_B_K1WphjVx7_2),.clk(gclk));
	jdff dff_B_y3jsG4hi1_2(.din(w_dff_B_K1WphjVx7_2),.dout(w_dff_B_y3jsG4hi1_2),.clk(gclk));
	jdff dff_B_wBCu0QuX0_2(.din(w_dff_B_y3jsG4hi1_2),.dout(w_dff_B_wBCu0QuX0_2),.clk(gclk));
	jdff dff_B_k9OXH5N45_2(.din(w_dff_B_wBCu0QuX0_2),.dout(w_dff_B_k9OXH5N45_2),.clk(gclk));
	jdff dff_B_mcAs9FME2_2(.din(w_dff_B_k9OXH5N45_2),.dout(w_dff_B_mcAs9FME2_2),.clk(gclk));
	jdff dff_B_xzlCFREP8_2(.din(w_dff_B_mcAs9FME2_2),.dout(w_dff_B_xzlCFREP8_2),.clk(gclk));
	jdff dff_B_EFUzlIud0_2(.din(w_dff_B_xzlCFREP8_2),.dout(w_dff_B_EFUzlIud0_2),.clk(gclk));
	jdff dff_B_0yo6G0Im4_2(.din(w_dff_B_EFUzlIud0_2),.dout(w_dff_B_0yo6G0Im4_2),.clk(gclk));
	jdff dff_B_KIwlVoas2_2(.din(w_dff_B_0yo6G0Im4_2),.dout(w_dff_B_KIwlVoas2_2),.clk(gclk));
	jdff dff_B_usAQ4Qhc7_2(.din(w_dff_B_KIwlVoas2_2),.dout(w_dff_B_usAQ4Qhc7_2),.clk(gclk));
	jdff dff_B_QKoOKo823_2(.din(w_dff_B_usAQ4Qhc7_2),.dout(w_dff_B_QKoOKo823_2),.clk(gclk));
	jdff dff_B_D7HvH2q07_2(.din(w_dff_B_QKoOKo823_2),.dout(w_dff_B_D7HvH2q07_2),.clk(gclk));
	jdff dff_B_iZ8Cg2jB2_2(.din(w_dff_B_D7HvH2q07_2),.dout(w_dff_B_iZ8Cg2jB2_2),.clk(gclk));
	jdff dff_B_XrxrqQa70_2(.din(w_dff_B_iZ8Cg2jB2_2),.dout(w_dff_B_XrxrqQa70_2),.clk(gclk));
	jdff dff_B_AimAZ4rY5_2(.din(w_dff_B_XrxrqQa70_2),.dout(w_dff_B_AimAZ4rY5_2),.clk(gclk));
	jdff dff_B_0mGKjRwK7_2(.din(w_dff_B_AimAZ4rY5_2),.dout(w_dff_B_0mGKjRwK7_2),.clk(gclk));
	jdff dff_B_SLqgLeUz6_2(.din(w_dff_B_0mGKjRwK7_2),.dout(w_dff_B_SLqgLeUz6_2),.clk(gclk));
	jdff dff_B_0Notq8cF1_2(.din(w_dff_B_SLqgLeUz6_2),.dout(w_dff_B_0Notq8cF1_2),.clk(gclk));
	jdff dff_B_cmmxr5wm9_2(.din(w_dff_B_0Notq8cF1_2),.dout(w_dff_B_cmmxr5wm9_2),.clk(gclk));
	jdff dff_B_HsDwihJM1_2(.din(w_dff_B_cmmxr5wm9_2),.dout(w_dff_B_HsDwihJM1_2),.clk(gclk));
	jdff dff_B_kU29M0Bi9_2(.din(w_dff_B_HsDwihJM1_2),.dout(w_dff_B_kU29M0Bi9_2),.clk(gclk));
	jdff dff_B_OO6lC5Ma8_2(.din(w_dff_B_kU29M0Bi9_2),.dout(w_dff_B_OO6lC5Ma8_2),.clk(gclk));
	jdff dff_B_u8os5wxt0_2(.din(w_dff_B_OO6lC5Ma8_2),.dout(w_dff_B_u8os5wxt0_2),.clk(gclk));
	jdff dff_B_9aw1YUF01_2(.din(w_dff_B_u8os5wxt0_2),.dout(w_dff_B_9aw1YUF01_2),.clk(gclk));
	jdff dff_B_H41Oumqr2_2(.din(w_dff_B_9aw1YUF01_2),.dout(w_dff_B_H41Oumqr2_2),.clk(gclk));
	jdff dff_B_MLozTtSE3_2(.din(w_dff_B_H41Oumqr2_2),.dout(w_dff_B_MLozTtSE3_2),.clk(gclk));
	jdff dff_B_u2iNC7Yd9_2(.din(w_dff_B_MLozTtSE3_2),.dout(w_dff_B_u2iNC7Yd9_2),.clk(gclk));
	jdff dff_B_lFhYoAov1_2(.din(w_dff_B_u2iNC7Yd9_2),.dout(w_dff_B_lFhYoAov1_2),.clk(gclk));
	jdff dff_B_FFxwMcAg2_2(.din(w_dff_B_lFhYoAov1_2),.dout(w_dff_B_FFxwMcAg2_2),.clk(gclk));
	jdff dff_B_4Kjf9Xzu5_2(.din(w_dff_B_FFxwMcAg2_2),.dout(w_dff_B_4Kjf9Xzu5_2),.clk(gclk));
	jdff dff_B_AUJVVuZs7_2(.din(n1702),.dout(w_dff_B_AUJVVuZs7_2),.clk(gclk));
	jdff dff_B_rhnCP9QY2_1(.din(n1700),.dout(w_dff_B_rhnCP9QY2_1),.clk(gclk));
	jdff dff_B_C7LHpqBI3_2(.din(n1658),.dout(w_dff_B_C7LHpqBI3_2),.clk(gclk));
	jdff dff_B_UeWfbcrz7_2(.din(w_dff_B_C7LHpqBI3_2),.dout(w_dff_B_UeWfbcrz7_2),.clk(gclk));
	jdff dff_B_n4tpqdkJ5_2(.din(w_dff_B_UeWfbcrz7_2),.dout(w_dff_B_n4tpqdkJ5_2),.clk(gclk));
	jdff dff_B_G7YogIVE9_2(.din(w_dff_B_n4tpqdkJ5_2),.dout(w_dff_B_G7YogIVE9_2),.clk(gclk));
	jdff dff_B_J8LjVr9Z2_2(.din(w_dff_B_G7YogIVE9_2),.dout(w_dff_B_J8LjVr9Z2_2),.clk(gclk));
	jdff dff_B_Y0KJbX4N0_2(.din(w_dff_B_J8LjVr9Z2_2),.dout(w_dff_B_Y0KJbX4N0_2),.clk(gclk));
	jdff dff_B_4qNiEXOt8_2(.din(w_dff_B_Y0KJbX4N0_2),.dout(w_dff_B_4qNiEXOt8_2),.clk(gclk));
	jdff dff_B_9kFeaxVf5_2(.din(w_dff_B_4qNiEXOt8_2),.dout(w_dff_B_9kFeaxVf5_2),.clk(gclk));
	jdff dff_B_HsptdJyG0_2(.din(w_dff_B_9kFeaxVf5_2),.dout(w_dff_B_HsptdJyG0_2),.clk(gclk));
	jdff dff_B_TKzAi6Gl3_2(.din(w_dff_B_HsptdJyG0_2),.dout(w_dff_B_TKzAi6Gl3_2),.clk(gclk));
	jdff dff_B_6ynsMQ2l0_2(.din(w_dff_B_TKzAi6Gl3_2),.dout(w_dff_B_6ynsMQ2l0_2),.clk(gclk));
	jdff dff_B_bhnIZjwp3_2(.din(w_dff_B_6ynsMQ2l0_2),.dout(w_dff_B_bhnIZjwp3_2),.clk(gclk));
	jdff dff_B_tXVk6FcT9_2(.din(w_dff_B_bhnIZjwp3_2),.dout(w_dff_B_tXVk6FcT9_2),.clk(gclk));
	jdff dff_B_58LdgK666_2(.din(w_dff_B_tXVk6FcT9_2),.dout(w_dff_B_58LdgK666_2),.clk(gclk));
	jdff dff_B_gzIk7S020_2(.din(w_dff_B_58LdgK666_2),.dout(w_dff_B_gzIk7S020_2),.clk(gclk));
	jdff dff_B_szxKorJG7_2(.din(w_dff_B_gzIk7S020_2),.dout(w_dff_B_szxKorJG7_2),.clk(gclk));
	jdff dff_B_f5OiTOd96_2(.din(w_dff_B_szxKorJG7_2),.dout(w_dff_B_f5OiTOd96_2),.clk(gclk));
	jdff dff_B_e6WLPQm50_2(.din(w_dff_B_f5OiTOd96_2),.dout(w_dff_B_e6WLPQm50_2),.clk(gclk));
	jdff dff_B_2F000M8A6_2(.din(w_dff_B_e6WLPQm50_2),.dout(w_dff_B_2F000M8A6_2),.clk(gclk));
	jdff dff_B_IFocsjVe8_2(.din(w_dff_B_2F000M8A6_2),.dout(w_dff_B_IFocsjVe8_2),.clk(gclk));
	jdff dff_B_1Y0NbcHw4_2(.din(w_dff_B_IFocsjVe8_2),.dout(w_dff_B_1Y0NbcHw4_2),.clk(gclk));
	jdff dff_B_8w1rBpYa0_2(.din(w_dff_B_1Y0NbcHw4_2),.dout(w_dff_B_8w1rBpYa0_2),.clk(gclk));
	jdff dff_B_eGCw48JR6_2(.din(w_dff_B_8w1rBpYa0_2),.dout(w_dff_B_eGCw48JR6_2),.clk(gclk));
	jdff dff_B_Ym96BF5n5_2(.din(w_dff_B_eGCw48JR6_2),.dout(w_dff_B_Ym96BF5n5_2),.clk(gclk));
	jdff dff_B_7GNR9CiQ1_2(.din(w_dff_B_Ym96BF5n5_2),.dout(w_dff_B_7GNR9CiQ1_2),.clk(gclk));
	jdff dff_B_jydhBZkv3_2(.din(w_dff_B_7GNR9CiQ1_2),.dout(w_dff_B_jydhBZkv3_2),.clk(gclk));
	jdff dff_B_XwbwARax8_2(.din(w_dff_B_jydhBZkv3_2),.dout(w_dff_B_XwbwARax8_2),.clk(gclk));
	jdff dff_B_XUXLl9PZ6_2(.din(w_dff_B_XwbwARax8_2),.dout(w_dff_B_XUXLl9PZ6_2),.clk(gclk));
	jdff dff_B_9s5BgiKq1_2(.din(w_dff_B_XUXLl9PZ6_2),.dout(w_dff_B_9s5BgiKq1_2),.clk(gclk));
	jdff dff_B_cbhmIanl0_2(.din(w_dff_B_9s5BgiKq1_2),.dout(w_dff_B_cbhmIanl0_2),.clk(gclk));
	jdff dff_B_53C2nhS84_2(.din(w_dff_B_cbhmIanl0_2),.dout(w_dff_B_53C2nhS84_2),.clk(gclk));
	jdff dff_B_UbLtddzG5_2(.din(w_dff_B_53C2nhS84_2),.dout(w_dff_B_UbLtddzG5_2),.clk(gclk));
	jdff dff_B_KsXZ429F1_2(.din(w_dff_B_UbLtddzG5_2),.dout(w_dff_B_KsXZ429F1_2),.clk(gclk));
	jdff dff_B_rrGJcutx6_2(.din(w_dff_B_KsXZ429F1_2),.dout(w_dff_B_rrGJcutx6_2),.clk(gclk));
	jdff dff_B_mdjShcxc7_2(.din(w_dff_B_rrGJcutx6_2),.dout(w_dff_B_mdjShcxc7_2),.clk(gclk));
	jdff dff_B_6MPxDqRq9_2(.din(w_dff_B_mdjShcxc7_2),.dout(w_dff_B_6MPxDqRq9_2),.clk(gclk));
	jdff dff_B_Uj77CKxn5_2(.din(w_dff_B_6MPxDqRq9_2),.dout(w_dff_B_Uj77CKxn5_2),.clk(gclk));
	jdff dff_B_VDZ8DIOG4_2(.din(w_dff_B_Uj77CKxn5_2),.dout(w_dff_B_VDZ8DIOG4_2),.clk(gclk));
	jdff dff_B_lS3yPT7e4_2(.din(w_dff_B_VDZ8DIOG4_2),.dout(w_dff_B_lS3yPT7e4_2),.clk(gclk));
	jdff dff_B_8uBAOWGH5_2(.din(w_dff_B_lS3yPT7e4_2),.dout(w_dff_B_8uBAOWGH5_2),.clk(gclk));
	jdff dff_B_26cPxGU03_2(.din(w_dff_B_8uBAOWGH5_2),.dout(w_dff_B_26cPxGU03_2),.clk(gclk));
	jdff dff_B_LrqcIO5M8_2(.din(w_dff_B_26cPxGU03_2),.dout(w_dff_B_LrqcIO5M8_2),.clk(gclk));
	jdff dff_B_aE2A8Mk01_2(.din(w_dff_B_LrqcIO5M8_2),.dout(w_dff_B_aE2A8Mk01_2),.clk(gclk));
	jdff dff_B_x0b2LiBp2_2(.din(w_dff_B_aE2A8Mk01_2),.dout(w_dff_B_x0b2LiBp2_2),.clk(gclk));
	jdff dff_B_oh5mULbq1_2(.din(n1661),.dout(w_dff_B_oh5mULbq1_2),.clk(gclk));
	jdff dff_B_eWtrvpIs8_1(.din(n1659),.dout(w_dff_B_eWtrvpIs8_1),.clk(gclk));
	jdff dff_B_SEXWdAiT6_2(.din(n1607),.dout(w_dff_B_SEXWdAiT6_2),.clk(gclk));
	jdff dff_B_mNob9bnb3_2(.din(w_dff_B_SEXWdAiT6_2),.dout(w_dff_B_mNob9bnb3_2),.clk(gclk));
	jdff dff_B_Rq2NlqbI9_2(.din(w_dff_B_mNob9bnb3_2),.dout(w_dff_B_Rq2NlqbI9_2),.clk(gclk));
	jdff dff_B_Mx0VVGVZ5_2(.din(w_dff_B_Rq2NlqbI9_2),.dout(w_dff_B_Mx0VVGVZ5_2),.clk(gclk));
	jdff dff_B_dViLjMkg3_2(.din(w_dff_B_Mx0VVGVZ5_2),.dout(w_dff_B_dViLjMkg3_2),.clk(gclk));
	jdff dff_B_2ZNy9ijD6_2(.din(w_dff_B_dViLjMkg3_2),.dout(w_dff_B_2ZNy9ijD6_2),.clk(gclk));
	jdff dff_B_zYGaFDGy4_2(.din(w_dff_B_2ZNy9ijD6_2),.dout(w_dff_B_zYGaFDGy4_2),.clk(gclk));
	jdff dff_B_tEeN3z9T5_2(.din(w_dff_B_zYGaFDGy4_2),.dout(w_dff_B_tEeN3z9T5_2),.clk(gclk));
	jdff dff_B_AxSFZzne9_2(.din(w_dff_B_tEeN3z9T5_2),.dout(w_dff_B_AxSFZzne9_2),.clk(gclk));
	jdff dff_B_tWQnD0L75_2(.din(w_dff_B_AxSFZzne9_2),.dout(w_dff_B_tWQnD0L75_2),.clk(gclk));
	jdff dff_B_sDYprePW0_2(.din(w_dff_B_tWQnD0L75_2),.dout(w_dff_B_sDYprePW0_2),.clk(gclk));
	jdff dff_B_WQqs7YsP8_2(.din(w_dff_B_sDYprePW0_2),.dout(w_dff_B_WQqs7YsP8_2),.clk(gclk));
	jdff dff_B_OG5ng1w95_2(.din(w_dff_B_WQqs7YsP8_2),.dout(w_dff_B_OG5ng1w95_2),.clk(gclk));
	jdff dff_B_MiR8bfbQ0_2(.din(w_dff_B_OG5ng1w95_2),.dout(w_dff_B_MiR8bfbQ0_2),.clk(gclk));
	jdff dff_B_YZLiTGSk0_2(.din(w_dff_B_MiR8bfbQ0_2),.dout(w_dff_B_YZLiTGSk0_2),.clk(gclk));
	jdff dff_B_EnkYOP629_2(.din(w_dff_B_YZLiTGSk0_2),.dout(w_dff_B_EnkYOP629_2),.clk(gclk));
	jdff dff_B_Mr0QJ2Rl2_2(.din(w_dff_B_EnkYOP629_2),.dout(w_dff_B_Mr0QJ2Rl2_2),.clk(gclk));
	jdff dff_B_7Sbwzsal4_2(.din(w_dff_B_Mr0QJ2Rl2_2),.dout(w_dff_B_7Sbwzsal4_2),.clk(gclk));
	jdff dff_B_ZBxEJg4i8_2(.din(w_dff_B_7Sbwzsal4_2),.dout(w_dff_B_ZBxEJg4i8_2),.clk(gclk));
	jdff dff_B_D6LTuJuE5_2(.din(w_dff_B_ZBxEJg4i8_2),.dout(w_dff_B_D6LTuJuE5_2),.clk(gclk));
	jdff dff_B_saW3zqss9_2(.din(w_dff_B_D6LTuJuE5_2),.dout(w_dff_B_saW3zqss9_2),.clk(gclk));
	jdff dff_B_KcjWQJfm3_2(.din(w_dff_B_saW3zqss9_2),.dout(w_dff_B_KcjWQJfm3_2),.clk(gclk));
	jdff dff_B_i9E5E1I67_2(.din(w_dff_B_KcjWQJfm3_2),.dout(w_dff_B_i9E5E1I67_2),.clk(gclk));
	jdff dff_B_JW1bkQxN0_2(.din(w_dff_B_i9E5E1I67_2),.dout(w_dff_B_JW1bkQxN0_2),.clk(gclk));
	jdff dff_B_e2OkxWGi5_2(.din(w_dff_B_JW1bkQxN0_2),.dout(w_dff_B_e2OkxWGi5_2),.clk(gclk));
	jdff dff_B_xJhJw2nF1_2(.din(w_dff_B_e2OkxWGi5_2),.dout(w_dff_B_xJhJw2nF1_2),.clk(gclk));
	jdff dff_B_wXwwq99M3_2(.din(w_dff_B_xJhJw2nF1_2),.dout(w_dff_B_wXwwq99M3_2),.clk(gclk));
	jdff dff_B_GbvRjd4Z4_2(.din(w_dff_B_wXwwq99M3_2),.dout(w_dff_B_GbvRjd4Z4_2),.clk(gclk));
	jdff dff_B_wEKKARbf3_2(.din(w_dff_B_GbvRjd4Z4_2),.dout(w_dff_B_wEKKARbf3_2),.clk(gclk));
	jdff dff_B_Apw4MyEK7_2(.din(w_dff_B_wEKKARbf3_2),.dout(w_dff_B_Apw4MyEK7_2),.clk(gclk));
	jdff dff_B_vVS5O0Tl3_2(.din(w_dff_B_Apw4MyEK7_2),.dout(w_dff_B_vVS5O0Tl3_2),.clk(gclk));
	jdff dff_B_bhfZ3va88_2(.din(w_dff_B_vVS5O0Tl3_2),.dout(w_dff_B_bhfZ3va88_2),.clk(gclk));
	jdff dff_B_P4om3MHF6_2(.din(w_dff_B_bhfZ3va88_2),.dout(w_dff_B_P4om3MHF6_2),.clk(gclk));
	jdff dff_B_ulKX7iad3_2(.din(w_dff_B_P4om3MHF6_2),.dout(w_dff_B_ulKX7iad3_2),.clk(gclk));
	jdff dff_B_7qJFgdvK6_2(.din(w_dff_B_ulKX7iad3_2),.dout(w_dff_B_7qJFgdvK6_2),.clk(gclk));
	jdff dff_B_1c96IQu83_2(.din(w_dff_B_7qJFgdvK6_2),.dout(w_dff_B_1c96IQu83_2),.clk(gclk));
	jdff dff_B_9Dh0EJpF6_2(.din(w_dff_B_1c96IQu83_2),.dout(w_dff_B_9Dh0EJpF6_2),.clk(gclk));
	jdff dff_B_wYij6kNY8_2(.din(w_dff_B_9Dh0EJpF6_2),.dout(w_dff_B_wYij6kNY8_2),.clk(gclk));
	jdff dff_B_4GVMkThx5_2(.din(w_dff_B_wYij6kNY8_2),.dout(w_dff_B_4GVMkThx5_2),.clk(gclk));
	jdff dff_B_KFTi04Gr6_2(.din(w_dff_B_4GVMkThx5_2),.dout(w_dff_B_KFTi04Gr6_2),.clk(gclk));
	jdff dff_B_lTDcgB0E7_2(.din(n1610),.dout(w_dff_B_lTDcgB0E7_2),.clk(gclk));
	jdff dff_B_EBXg5wWk4_1(.din(n1608),.dout(w_dff_B_EBXg5wWk4_1),.clk(gclk));
	jdff dff_B_CS0Eygq89_2(.din(n1550),.dout(w_dff_B_CS0Eygq89_2),.clk(gclk));
	jdff dff_B_tZDpSqCR3_2(.din(w_dff_B_CS0Eygq89_2),.dout(w_dff_B_tZDpSqCR3_2),.clk(gclk));
	jdff dff_B_KbDKyaV90_2(.din(w_dff_B_tZDpSqCR3_2),.dout(w_dff_B_KbDKyaV90_2),.clk(gclk));
	jdff dff_B_aNfeVkdx7_2(.din(w_dff_B_KbDKyaV90_2),.dout(w_dff_B_aNfeVkdx7_2),.clk(gclk));
	jdff dff_B_HjDldspW8_2(.din(w_dff_B_aNfeVkdx7_2),.dout(w_dff_B_HjDldspW8_2),.clk(gclk));
	jdff dff_B_vsXKsXhd8_2(.din(w_dff_B_HjDldspW8_2),.dout(w_dff_B_vsXKsXhd8_2),.clk(gclk));
	jdff dff_B_mworufgv5_2(.din(w_dff_B_vsXKsXhd8_2),.dout(w_dff_B_mworufgv5_2),.clk(gclk));
	jdff dff_B_EAgftY1d4_2(.din(w_dff_B_mworufgv5_2),.dout(w_dff_B_EAgftY1d4_2),.clk(gclk));
	jdff dff_B_5mH1526m9_2(.din(w_dff_B_EAgftY1d4_2),.dout(w_dff_B_5mH1526m9_2),.clk(gclk));
	jdff dff_B_MGMWnnIC6_2(.din(w_dff_B_5mH1526m9_2),.dout(w_dff_B_MGMWnnIC6_2),.clk(gclk));
	jdff dff_B_gsLYPoQi5_2(.din(w_dff_B_MGMWnnIC6_2),.dout(w_dff_B_gsLYPoQi5_2),.clk(gclk));
	jdff dff_B_EznCGRIn1_2(.din(w_dff_B_gsLYPoQi5_2),.dout(w_dff_B_EznCGRIn1_2),.clk(gclk));
	jdff dff_B_CHsZoZUY8_2(.din(w_dff_B_EznCGRIn1_2),.dout(w_dff_B_CHsZoZUY8_2),.clk(gclk));
	jdff dff_B_JsWHldx16_2(.din(w_dff_B_CHsZoZUY8_2),.dout(w_dff_B_JsWHldx16_2),.clk(gclk));
	jdff dff_B_LYm6CVXr4_2(.din(w_dff_B_JsWHldx16_2),.dout(w_dff_B_LYm6CVXr4_2),.clk(gclk));
	jdff dff_B_jWypSJo20_2(.din(w_dff_B_LYm6CVXr4_2),.dout(w_dff_B_jWypSJo20_2),.clk(gclk));
	jdff dff_B_Sqw4sEgo6_2(.din(w_dff_B_jWypSJo20_2),.dout(w_dff_B_Sqw4sEgo6_2),.clk(gclk));
	jdff dff_B_kVl59ngq4_2(.din(w_dff_B_Sqw4sEgo6_2),.dout(w_dff_B_kVl59ngq4_2),.clk(gclk));
	jdff dff_B_k48YUVn62_2(.din(w_dff_B_kVl59ngq4_2),.dout(w_dff_B_k48YUVn62_2),.clk(gclk));
	jdff dff_B_JXehVPJs1_2(.din(w_dff_B_k48YUVn62_2),.dout(w_dff_B_JXehVPJs1_2),.clk(gclk));
	jdff dff_B_d9IGH2WH9_2(.din(w_dff_B_JXehVPJs1_2),.dout(w_dff_B_d9IGH2WH9_2),.clk(gclk));
	jdff dff_B_EFMcX0Bi4_2(.din(w_dff_B_d9IGH2WH9_2),.dout(w_dff_B_EFMcX0Bi4_2),.clk(gclk));
	jdff dff_B_pBk6d6VG7_2(.din(w_dff_B_EFMcX0Bi4_2),.dout(w_dff_B_pBk6d6VG7_2),.clk(gclk));
	jdff dff_B_B7dy0SCz9_2(.din(w_dff_B_pBk6d6VG7_2),.dout(w_dff_B_B7dy0SCz9_2),.clk(gclk));
	jdff dff_B_wV1OtUmf9_2(.din(w_dff_B_B7dy0SCz9_2),.dout(w_dff_B_wV1OtUmf9_2),.clk(gclk));
	jdff dff_B_0fkp3bTY3_2(.din(w_dff_B_wV1OtUmf9_2),.dout(w_dff_B_0fkp3bTY3_2),.clk(gclk));
	jdff dff_B_Jug4uxFi6_2(.din(w_dff_B_0fkp3bTY3_2),.dout(w_dff_B_Jug4uxFi6_2),.clk(gclk));
	jdff dff_B_dHAEEWK13_2(.din(w_dff_B_Jug4uxFi6_2),.dout(w_dff_B_dHAEEWK13_2),.clk(gclk));
	jdff dff_B_fQPqUJfB7_2(.din(w_dff_B_dHAEEWK13_2),.dout(w_dff_B_fQPqUJfB7_2),.clk(gclk));
	jdff dff_B_dsG3ScMA0_2(.din(w_dff_B_fQPqUJfB7_2),.dout(w_dff_B_dsG3ScMA0_2),.clk(gclk));
	jdff dff_B_xXtdYtIG7_2(.din(w_dff_B_dsG3ScMA0_2),.dout(w_dff_B_xXtdYtIG7_2),.clk(gclk));
	jdff dff_B_MJMUtV6s6_2(.din(w_dff_B_xXtdYtIG7_2),.dout(w_dff_B_MJMUtV6s6_2),.clk(gclk));
	jdff dff_B_JAChyVXO1_2(.din(w_dff_B_MJMUtV6s6_2),.dout(w_dff_B_JAChyVXO1_2),.clk(gclk));
	jdff dff_B_cC53jNmb5_2(.din(w_dff_B_JAChyVXO1_2),.dout(w_dff_B_cC53jNmb5_2),.clk(gclk));
	jdff dff_B_Ypjycl5A1_2(.din(w_dff_B_cC53jNmb5_2),.dout(w_dff_B_Ypjycl5A1_2),.clk(gclk));
	jdff dff_B_Qs83rpz59_2(.din(w_dff_B_Ypjycl5A1_2),.dout(w_dff_B_Qs83rpz59_2),.clk(gclk));
	jdff dff_B_g95BrBah1_2(.din(n1553),.dout(w_dff_B_g95BrBah1_2),.clk(gclk));
	jdff dff_B_kTo0wJwr9_1(.din(n1551),.dout(w_dff_B_kTo0wJwr9_1),.clk(gclk));
	jdff dff_B_xXfvTIEd0_2(.din(n1486),.dout(w_dff_B_xXfvTIEd0_2),.clk(gclk));
	jdff dff_B_ctNTb8Vz8_2(.din(w_dff_B_xXfvTIEd0_2),.dout(w_dff_B_ctNTb8Vz8_2),.clk(gclk));
	jdff dff_B_OYTBoBDN5_2(.din(w_dff_B_ctNTb8Vz8_2),.dout(w_dff_B_OYTBoBDN5_2),.clk(gclk));
	jdff dff_B_sxvJC70M6_2(.din(w_dff_B_OYTBoBDN5_2),.dout(w_dff_B_sxvJC70M6_2),.clk(gclk));
	jdff dff_B_x7kPA3hh2_2(.din(w_dff_B_sxvJC70M6_2),.dout(w_dff_B_x7kPA3hh2_2),.clk(gclk));
	jdff dff_B_A0qOBcfU0_2(.din(w_dff_B_x7kPA3hh2_2),.dout(w_dff_B_A0qOBcfU0_2),.clk(gclk));
	jdff dff_B_dNMv3fYf8_2(.din(w_dff_B_A0qOBcfU0_2),.dout(w_dff_B_dNMv3fYf8_2),.clk(gclk));
	jdff dff_B_MLygmdTh6_2(.din(w_dff_B_dNMv3fYf8_2),.dout(w_dff_B_MLygmdTh6_2),.clk(gclk));
	jdff dff_B_qHf0FhW84_2(.din(w_dff_B_MLygmdTh6_2),.dout(w_dff_B_qHf0FhW84_2),.clk(gclk));
	jdff dff_B_hG1YzoXd2_2(.din(w_dff_B_qHf0FhW84_2),.dout(w_dff_B_hG1YzoXd2_2),.clk(gclk));
	jdff dff_B_EyEr9Flw2_2(.din(w_dff_B_hG1YzoXd2_2),.dout(w_dff_B_EyEr9Flw2_2),.clk(gclk));
	jdff dff_B_Yq8VIdSQ8_2(.din(w_dff_B_EyEr9Flw2_2),.dout(w_dff_B_Yq8VIdSQ8_2),.clk(gclk));
	jdff dff_B_Gku1QtqH0_2(.din(w_dff_B_Yq8VIdSQ8_2),.dout(w_dff_B_Gku1QtqH0_2),.clk(gclk));
	jdff dff_B_RNxEJiZe6_2(.din(w_dff_B_Gku1QtqH0_2),.dout(w_dff_B_RNxEJiZe6_2),.clk(gclk));
	jdff dff_B_m2PhG3Yg5_2(.din(w_dff_B_RNxEJiZe6_2),.dout(w_dff_B_m2PhG3Yg5_2),.clk(gclk));
	jdff dff_B_LxhWNwgI0_2(.din(w_dff_B_m2PhG3Yg5_2),.dout(w_dff_B_LxhWNwgI0_2),.clk(gclk));
	jdff dff_B_l56bxpkC6_2(.din(w_dff_B_LxhWNwgI0_2),.dout(w_dff_B_l56bxpkC6_2),.clk(gclk));
	jdff dff_B_YpCP5Imj6_2(.din(w_dff_B_l56bxpkC6_2),.dout(w_dff_B_YpCP5Imj6_2),.clk(gclk));
	jdff dff_B_Bf7M6seD1_2(.din(w_dff_B_YpCP5Imj6_2),.dout(w_dff_B_Bf7M6seD1_2),.clk(gclk));
	jdff dff_B_MmXmCIyY0_2(.din(w_dff_B_Bf7M6seD1_2),.dout(w_dff_B_MmXmCIyY0_2),.clk(gclk));
	jdff dff_B_Spc6bhKa1_2(.din(w_dff_B_MmXmCIyY0_2),.dout(w_dff_B_Spc6bhKa1_2),.clk(gclk));
	jdff dff_B_r5cNsBke1_2(.din(w_dff_B_Spc6bhKa1_2),.dout(w_dff_B_r5cNsBke1_2),.clk(gclk));
	jdff dff_B_nHrTzs1x6_2(.din(w_dff_B_r5cNsBke1_2),.dout(w_dff_B_nHrTzs1x6_2),.clk(gclk));
	jdff dff_B_z8BuF0Ov7_2(.din(w_dff_B_nHrTzs1x6_2),.dout(w_dff_B_z8BuF0Ov7_2),.clk(gclk));
	jdff dff_B_Qy6Ze7tF0_2(.din(w_dff_B_z8BuF0Ov7_2),.dout(w_dff_B_Qy6Ze7tF0_2),.clk(gclk));
	jdff dff_B_g8XNXJmE1_2(.din(w_dff_B_Qy6Ze7tF0_2),.dout(w_dff_B_g8XNXJmE1_2),.clk(gclk));
	jdff dff_B_YcrhXcAJ0_2(.din(w_dff_B_g8XNXJmE1_2),.dout(w_dff_B_YcrhXcAJ0_2),.clk(gclk));
	jdff dff_B_DyvprqCN1_2(.din(w_dff_B_YcrhXcAJ0_2),.dout(w_dff_B_DyvprqCN1_2),.clk(gclk));
	jdff dff_B_iVPqHczQ2_2(.din(w_dff_B_DyvprqCN1_2),.dout(w_dff_B_iVPqHczQ2_2),.clk(gclk));
	jdff dff_B_Ui4cwZhr5_2(.din(w_dff_B_iVPqHczQ2_2),.dout(w_dff_B_Ui4cwZhr5_2),.clk(gclk));
	jdff dff_B_ugUEf2eZ9_2(.din(w_dff_B_Ui4cwZhr5_2),.dout(w_dff_B_ugUEf2eZ9_2),.clk(gclk));
	jdff dff_B_6ZFVxRWY6_2(.din(w_dff_B_ugUEf2eZ9_2),.dout(w_dff_B_6ZFVxRWY6_2),.clk(gclk));
	jdff dff_B_IFTw00kJ0_1(.din(n1487),.dout(w_dff_B_IFTw00kJ0_1),.clk(gclk));
	jdff dff_B_RdtKvNYk3_2(.din(n1415),.dout(w_dff_B_RdtKvNYk3_2),.clk(gclk));
	jdff dff_B_PYP44jYz2_2(.din(w_dff_B_RdtKvNYk3_2),.dout(w_dff_B_PYP44jYz2_2),.clk(gclk));
	jdff dff_B_VC9rdrPe5_2(.din(w_dff_B_PYP44jYz2_2),.dout(w_dff_B_VC9rdrPe5_2),.clk(gclk));
	jdff dff_B_683VvSZM6_2(.din(w_dff_B_VC9rdrPe5_2),.dout(w_dff_B_683VvSZM6_2),.clk(gclk));
	jdff dff_B_HDIY0YNw2_2(.din(w_dff_B_683VvSZM6_2),.dout(w_dff_B_HDIY0YNw2_2),.clk(gclk));
	jdff dff_B_alUXG5IP2_2(.din(w_dff_B_HDIY0YNw2_2),.dout(w_dff_B_alUXG5IP2_2),.clk(gclk));
	jdff dff_B_SH10VcSh0_2(.din(w_dff_B_alUXG5IP2_2),.dout(w_dff_B_SH10VcSh0_2),.clk(gclk));
	jdff dff_B_7aTyqGo02_2(.din(w_dff_B_SH10VcSh0_2),.dout(w_dff_B_7aTyqGo02_2),.clk(gclk));
	jdff dff_B_plSKXuKT6_2(.din(w_dff_B_7aTyqGo02_2),.dout(w_dff_B_plSKXuKT6_2),.clk(gclk));
	jdff dff_B_EPFTNTCF3_2(.din(w_dff_B_plSKXuKT6_2),.dout(w_dff_B_EPFTNTCF3_2),.clk(gclk));
	jdff dff_B_Aqhfj5nR5_2(.din(w_dff_B_EPFTNTCF3_2),.dout(w_dff_B_Aqhfj5nR5_2),.clk(gclk));
	jdff dff_B_YfFf0rx90_2(.din(w_dff_B_Aqhfj5nR5_2),.dout(w_dff_B_YfFf0rx90_2),.clk(gclk));
	jdff dff_B_59uJ2E770_2(.din(w_dff_B_YfFf0rx90_2),.dout(w_dff_B_59uJ2E770_2),.clk(gclk));
	jdff dff_B_NU8mHIPF2_2(.din(w_dff_B_59uJ2E770_2),.dout(w_dff_B_NU8mHIPF2_2),.clk(gclk));
	jdff dff_B_Nh5cQURV0_2(.din(w_dff_B_NU8mHIPF2_2),.dout(w_dff_B_Nh5cQURV0_2),.clk(gclk));
	jdff dff_B_Qwg1tJgI4_2(.din(w_dff_B_Nh5cQURV0_2),.dout(w_dff_B_Qwg1tJgI4_2),.clk(gclk));
	jdff dff_B_oBTCs1Ic9_2(.din(w_dff_B_Qwg1tJgI4_2),.dout(w_dff_B_oBTCs1Ic9_2),.clk(gclk));
	jdff dff_B_XklLRYk78_2(.din(w_dff_B_oBTCs1Ic9_2),.dout(w_dff_B_XklLRYk78_2),.clk(gclk));
	jdff dff_B_GPxNX4dw3_2(.din(w_dff_B_XklLRYk78_2),.dout(w_dff_B_GPxNX4dw3_2),.clk(gclk));
	jdff dff_B_jDbtH2FR7_2(.din(w_dff_B_GPxNX4dw3_2),.dout(w_dff_B_jDbtH2FR7_2),.clk(gclk));
	jdff dff_B_7ezMDUGa6_2(.din(w_dff_B_jDbtH2FR7_2),.dout(w_dff_B_7ezMDUGa6_2),.clk(gclk));
	jdff dff_B_ieCxqmrM1_2(.din(w_dff_B_7ezMDUGa6_2),.dout(w_dff_B_ieCxqmrM1_2),.clk(gclk));
	jdff dff_B_58kcIXwr5_2(.din(w_dff_B_ieCxqmrM1_2),.dout(w_dff_B_58kcIXwr5_2),.clk(gclk));
	jdff dff_B_jgVScGte7_2(.din(w_dff_B_58kcIXwr5_2),.dout(w_dff_B_jgVScGte7_2),.clk(gclk));
	jdff dff_B_kVei2QwS4_2(.din(w_dff_B_jgVScGte7_2),.dout(w_dff_B_kVei2QwS4_2),.clk(gclk));
	jdff dff_B_G6KMSaKk6_2(.din(w_dff_B_kVei2QwS4_2),.dout(w_dff_B_G6KMSaKk6_2),.clk(gclk));
	jdff dff_B_0MYWOVCF2_2(.din(w_dff_B_G6KMSaKk6_2),.dout(w_dff_B_0MYWOVCF2_2),.clk(gclk));
	jdff dff_B_RqFGWpq18_2(.din(w_dff_B_0MYWOVCF2_2),.dout(w_dff_B_RqFGWpq18_2),.clk(gclk));
	jdff dff_B_SaWBszGf8_2(.din(w_dff_B_RqFGWpq18_2),.dout(w_dff_B_SaWBszGf8_2),.clk(gclk));
	jdff dff_B_DMjZiILv3_2(.din(n1440),.dout(w_dff_B_DMjZiILv3_2),.clk(gclk));
	jdff dff_B_P7pV3xtN2_1(.din(n1416),.dout(w_dff_B_P7pV3xtN2_1),.clk(gclk));
	jdff dff_B_cAv5JQXD4_2(.din(n1337),.dout(w_dff_B_cAv5JQXD4_2),.clk(gclk));
	jdff dff_B_Ci97n3TX3_2(.din(w_dff_B_cAv5JQXD4_2),.dout(w_dff_B_Ci97n3TX3_2),.clk(gclk));
	jdff dff_B_QUZc3E899_2(.din(w_dff_B_Ci97n3TX3_2),.dout(w_dff_B_QUZc3E899_2),.clk(gclk));
	jdff dff_B_OXQttdKS8_2(.din(w_dff_B_QUZc3E899_2),.dout(w_dff_B_OXQttdKS8_2),.clk(gclk));
	jdff dff_B_MrVLvbVi6_2(.din(w_dff_B_OXQttdKS8_2),.dout(w_dff_B_MrVLvbVi6_2),.clk(gclk));
	jdff dff_B_2r5jHqnC5_2(.din(w_dff_B_MrVLvbVi6_2),.dout(w_dff_B_2r5jHqnC5_2),.clk(gclk));
	jdff dff_B_yNIcBTNp0_2(.din(w_dff_B_2r5jHqnC5_2),.dout(w_dff_B_yNIcBTNp0_2),.clk(gclk));
	jdff dff_B_uLGDsaIN0_2(.din(w_dff_B_yNIcBTNp0_2),.dout(w_dff_B_uLGDsaIN0_2),.clk(gclk));
	jdff dff_B_y1WSSNpM2_2(.din(w_dff_B_uLGDsaIN0_2),.dout(w_dff_B_y1WSSNpM2_2),.clk(gclk));
	jdff dff_B_YtGwdiAQ3_2(.din(w_dff_B_y1WSSNpM2_2),.dout(w_dff_B_YtGwdiAQ3_2),.clk(gclk));
	jdff dff_B_qe8iiywU7_2(.din(w_dff_B_YtGwdiAQ3_2),.dout(w_dff_B_qe8iiywU7_2),.clk(gclk));
	jdff dff_B_6l0Wpm4N9_2(.din(w_dff_B_qe8iiywU7_2),.dout(w_dff_B_6l0Wpm4N9_2),.clk(gclk));
	jdff dff_B_VZVm6zFy0_2(.din(w_dff_B_6l0Wpm4N9_2),.dout(w_dff_B_VZVm6zFy0_2),.clk(gclk));
	jdff dff_B_q2C1g8q56_2(.din(w_dff_B_VZVm6zFy0_2),.dout(w_dff_B_q2C1g8q56_2),.clk(gclk));
	jdff dff_B_boap64Cn4_2(.din(w_dff_B_q2C1g8q56_2),.dout(w_dff_B_boap64Cn4_2),.clk(gclk));
	jdff dff_B_oxSfq6k95_2(.din(w_dff_B_boap64Cn4_2),.dout(w_dff_B_oxSfq6k95_2),.clk(gclk));
	jdff dff_B_WVnCnoJi5_2(.din(w_dff_B_oxSfq6k95_2),.dout(w_dff_B_WVnCnoJi5_2),.clk(gclk));
	jdff dff_B_Q0dkQHni8_2(.din(w_dff_B_WVnCnoJi5_2),.dout(w_dff_B_Q0dkQHni8_2),.clk(gclk));
	jdff dff_B_xlSSTIkI9_2(.din(w_dff_B_Q0dkQHni8_2),.dout(w_dff_B_xlSSTIkI9_2),.clk(gclk));
	jdff dff_B_rUa4M8Eg4_2(.din(w_dff_B_xlSSTIkI9_2),.dout(w_dff_B_rUa4M8Eg4_2),.clk(gclk));
	jdff dff_B_OTarkhj05_2(.din(w_dff_B_rUa4M8Eg4_2),.dout(w_dff_B_OTarkhj05_2),.clk(gclk));
	jdff dff_B_Xh3xVpyD0_2(.din(w_dff_B_OTarkhj05_2),.dout(w_dff_B_Xh3xVpyD0_2),.clk(gclk));
	jdff dff_B_7AhYg2xx1_2(.din(w_dff_B_Xh3xVpyD0_2),.dout(w_dff_B_7AhYg2xx1_2),.clk(gclk));
	jdff dff_B_IDndbqFh3_2(.din(w_dff_B_7AhYg2xx1_2),.dout(w_dff_B_IDndbqFh3_2),.clk(gclk));
	jdff dff_B_MbvSBqjA3_2(.din(w_dff_B_IDndbqFh3_2),.dout(w_dff_B_MbvSBqjA3_2),.clk(gclk));
	jdff dff_B_59Rap77Z8_2(.din(w_dff_B_MbvSBqjA3_2),.dout(w_dff_B_59Rap77Z8_2),.clk(gclk));
	jdff dff_B_8SaeRHr09_2(.din(n1362),.dout(w_dff_B_8SaeRHr09_2),.clk(gclk));
	jdff dff_B_fvBuavZm2_1(.din(n1338),.dout(w_dff_B_fvBuavZm2_1),.clk(gclk));
	jdff dff_B_rikRDUoQ1_2(.din(n1252),.dout(w_dff_B_rikRDUoQ1_2),.clk(gclk));
	jdff dff_B_ODqYfBd60_2(.din(w_dff_B_rikRDUoQ1_2),.dout(w_dff_B_ODqYfBd60_2),.clk(gclk));
	jdff dff_B_stjmCUix9_2(.din(w_dff_B_ODqYfBd60_2),.dout(w_dff_B_stjmCUix9_2),.clk(gclk));
	jdff dff_B_W1CnToUL2_2(.din(w_dff_B_stjmCUix9_2),.dout(w_dff_B_W1CnToUL2_2),.clk(gclk));
	jdff dff_B_nQibsh9b1_2(.din(w_dff_B_W1CnToUL2_2),.dout(w_dff_B_nQibsh9b1_2),.clk(gclk));
	jdff dff_B_kKp3HgM66_2(.din(w_dff_B_nQibsh9b1_2),.dout(w_dff_B_kKp3HgM66_2),.clk(gclk));
	jdff dff_B_umLtDdPn9_2(.din(w_dff_B_kKp3HgM66_2),.dout(w_dff_B_umLtDdPn9_2),.clk(gclk));
	jdff dff_B_BPR8izXS1_2(.din(w_dff_B_umLtDdPn9_2),.dout(w_dff_B_BPR8izXS1_2),.clk(gclk));
	jdff dff_B_qkOfTQAf0_2(.din(w_dff_B_BPR8izXS1_2),.dout(w_dff_B_qkOfTQAf0_2),.clk(gclk));
	jdff dff_B_WLXmD37M5_2(.din(w_dff_B_qkOfTQAf0_2),.dout(w_dff_B_WLXmD37M5_2),.clk(gclk));
	jdff dff_B_1jGcuY3J0_2(.din(w_dff_B_WLXmD37M5_2),.dout(w_dff_B_1jGcuY3J0_2),.clk(gclk));
	jdff dff_B_MssQaZhz4_2(.din(w_dff_B_1jGcuY3J0_2),.dout(w_dff_B_MssQaZhz4_2),.clk(gclk));
	jdff dff_B_4Y6TmLK67_2(.din(w_dff_B_MssQaZhz4_2),.dout(w_dff_B_4Y6TmLK67_2),.clk(gclk));
	jdff dff_B_aI1Fc56f5_2(.din(w_dff_B_4Y6TmLK67_2),.dout(w_dff_B_aI1Fc56f5_2),.clk(gclk));
	jdff dff_B_3pmW3EdN4_2(.din(w_dff_B_aI1Fc56f5_2),.dout(w_dff_B_3pmW3EdN4_2),.clk(gclk));
	jdff dff_B_72SL8DNq3_2(.din(w_dff_B_3pmW3EdN4_2),.dout(w_dff_B_72SL8DNq3_2),.clk(gclk));
	jdff dff_B_LGk9zbWS5_2(.din(w_dff_B_72SL8DNq3_2),.dout(w_dff_B_LGk9zbWS5_2),.clk(gclk));
	jdff dff_B_O5NBdmpQ8_2(.din(w_dff_B_LGk9zbWS5_2),.dout(w_dff_B_O5NBdmpQ8_2),.clk(gclk));
	jdff dff_B_2AiuQ0aa5_2(.din(w_dff_B_O5NBdmpQ8_2),.dout(w_dff_B_2AiuQ0aa5_2),.clk(gclk));
	jdff dff_B_R4gBO1sg1_2(.din(w_dff_B_2AiuQ0aa5_2),.dout(w_dff_B_R4gBO1sg1_2),.clk(gclk));
	jdff dff_B_6S7DUVKu4_2(.din(w_dff_B_R4gBO1sg1_2),.dout(w_dff_B_6S7DUVKu4_2),.clk(gclk));
	jdff dff_B_s3V2nT0A2_2(.din(w_dff_B_6S7DUVKu4_2),.dout(w_dff_B_s3V2nT0A2_2),.clk(gclk));
	jdff dff_B_mIQobraJ3_2(.din(w_dff_B_s3V2nT0A2_2),.dout(w_dff_B_mIQobraJ3_2),.clk(gclk));
	jdff dff_B_FU4KmCfZ3_2(.din(n1277),.dout(w_dff_B_FU4KmCfZ3_2),.clk(gclk));
	jdff dff_B_8eTcrcM07_1(.din(n1253),.dout(w_dff_B_8eTcrcM07_1),.clk(gclk));
	jdff dff_B_BpDJCnWy6_2(.din(n1161),.dout(w_dff_B_BpDJCnWy6_2),.clk(gclk));
	jdff dff_B_c4Ac7gBD1_2(.din(w_dff_B_BpDJCnWy6_2),.dout(w_dff_B_c4Ac7gBD1_2),.clk(gclk));
	jdff dff_B_q5sa0PWj0_2(.din(w_dff_B_c4Ac7gBD1_2),.dout(w_dff_B_q5sa0PWj0_2),.clk(gclk));
	jdff dff_B_embPnHVU0_2(.din(w_dff_B_q5sa0PWj0_2),.dout(w_dff_B_embPnHVU0_2),.clk(gclk));
	jdff dff_B_VdXsQq5V5_2(.din(w_dff_B_embPnHVU0_2),.dout(w_dff_B_VdXsQq5V5_2),.clk(gclk));
	jdff dff_B_ClWm7J4h1_2(.din(w_dff_B_VdXsQq5V5_2),.dout(w_dff_B_ClWm7J4h1_2),.clk(gclk));
	jdff dff_B_96uQTumw9_2(.din(w_dff_B_ClWm7J4h1_2),.dout(w_dff_B_96uQTumw9_2),.clk(gclk));
	jdff dff_B_ZlA23hll0_2(.din(w_dff_B_96uQTumw9_2),.dout(w_dff_B_ZlA23hll0_2),.clk(gclk));
	jdff dff_B_8DPtsfbq1_2(.din(w_dff_B_ZlA23hll0_2),.dout(w_dff_B_8DPtsfbq1_2),.clk(gclk));
	jdff dff_B_1qKzQJJP8_2(.din(w_dff_B_8DPtsfbq1_2),.dout(w_dff_B_1qKzQJJP8_2),.clk(gclk));
	jdff dff_B_M0w7T2lc0_2(.din(w_dff_B_1qKzQJJP8_2),.dout(w_dff_B_M0w7T2lc0_2),.clk(gclk));
	jdff dff_B_mBifnvAS7_2(.din(w_dff_B_M0w7T2lc0_2),.dout(w_dff_B_mBifnvAS7_2),.clk(gclk));
	jdff dff_B_8JcM7pM71_2(.din(w_dff_B_mBifnvAS7_2),.dout(w_dff_B_8JcM7pM71_2),.clk(gclk));
	jdff dff_B_EwOgen9I2_2(.din(w_dff_B_8JcM7pM71_2),.dout(w_dff_B_EwOgen9I2_2),.clk(gclk));
	jdff dff_B_Vcf7JBKS5_2(.din(w_dff_B_EwOgen9I2_2),.dout(w_dff_B_Vcf7JBKS5_2),.clk(gclk));
	jdff dff_B_e7VYbVbi1_2(.din(w_dff_B_Vcf7JBKS5_2),.dout(w_dff_B_e7VYbVbi1_2),.clk(gclk));
	jdff dff_B_9pHvuOoV7_2(.din(w_dff_B_e7VYbVbi1_2),.dout(w_dff_B_9pHvuOoV7_2),.clk(gclk));
	jdff dff_B_83EA3s7T5_2(.din(w_dff_B_9pHvuOoV7_2),.dout(w_dff_B_83EA3s7T5_2),.clk(gclk));
	jdff dff_B_V6q3kUu22_2(.din(w_dff_B_83EA3s7T5_2),.dout(w_dff_B_V6q3kUu22_2),.clk(gclk));
	jdff dff_B_sx23HeQZ2_2(.din(w_dff_B_V6q3kUu22_2),.dout(w_dff_B_sx23HeQZ2_2),.clk(gclk));
	jdff dff_B_aZm2xLBW4_2(.din(n1186),.dout(w_dff_B_aZm2xLBW4_2),.clk(gclk));
	jdff dff_B_S4B5uJt66_1(.din(n1162),.dout(w_dff_B_S4B5uJt66_1),.clk(gclk));
	jdff dff_B_WJNUuhNB8_2(.din(n1063),.dout(w_dff_B_WJNUuhNB8_2),.clk(gclk));
	jdff dff_B_ErLCSPMA9_2(.din(w_dff_B_WJNUuhNB8_2),.dout(w_dff_B_ErLCSPMA9_2),.clk(gclk));
	jdff dff_B_3U4Xjlvm5_2(.din(w_dff_B_ErLCSPMA9_2),.dout(w_dff_B_3U4Xjlvm5_2),.clk(gclk));
	jdff dff_B_7nm19qju8_2(.din(w_dff_B_3U4Xjlvm5_2),.dout(w_dff_B_7nm19qju8_2),.clk(gclk));
	jdff dff_B_3fJvhWbh9_2(.din(w_dff_B_7nm19qju8_2),.dout(w_dff_B_3fJvhWbh9_2),.clk(gclk));
	jdff dff_B_oSfWurtQ4_2(.din(w_dff_B_3fJvhWbh9_2),.dout(w_dff_B_oSfWurtQ4_2),.clk(gclk));
	jdff dff_B_f4WRCaVE0_2(.din(w_dff_B_oSfWurtQ4_2),.dout(w_dff_B_f4WRCaVE0_2),.clk(gclk));
	jdff dff_B_2Mtrg2IV3_2(.din(w_dff_B_f4WRCaVE0_2),.dout(w_dff_B_2Mtrg2IV3_2),.clk(gclk));
	jdff dff_B_1F4gxY6Q7_2(.din(w_dff_B_2Mtrg2IV3_2),.dout(w_dff_B_1F4gxY6Q7_2),.clk(gclk));
	jdff dff_B_NuWwU2qs6_2(.din(w_dff_B_1F4gxY6Q7_2),.dout(w_dff_B_NuWwU2qs6_2),.clk(gclk));
	jdff dff_B_MIncjyIH1_2(.din(w_dff_B_NuWwU2qs6_2),.dout(w_dff_B_MIncjyIH1_2),.clk(gclk));
	jdff dff_B_ZgAoVJIJ3_2(.din(w_dff_B_MIncjyIH1_2),.dout(w_dff_B_ZgAoVJIJ3_2),.clk(gclk));
	jdff dff_B_efVkfXK28_2(.din(w_dff_B_ZgAoVJIJ3_2),.dout(w_dff_B_efVkfXK28_2),.clk(gclk));
	jdff dff_B_kFYl820U7_2(.din(w_dff_B_efVkfXK28_2),.dout(w_dff_B_kFYl820U7_2),.clk(gclk));
	jdff dff_B_M8n77AtN2_2(.din(w_dff_B_kFYl820U7_2),.dout(w_dff_B_M8n77AtN2_2),.clk(gclk));
	jdff dff_B_qFN8LtCW0_2(.din(w_dff_B_M8n77AtN2_2),.dout(w_dff_B_qFN8LtCW0_2),.clk(gclk));
	jdff dff_B_7weLBBiR8_2(.din(w_dff_B_qFN8LtCW0_2),.dout(w_dff_B_7weLBBiR8_2),.clk(gclk));
	jdff dff_B_3TVnsZem2_2(.din(n1087),.dout(w_dff_B_3TVnsZem2_2),.clk(gclk));
	jdff dff_B_tEIsuwSY6_1(.din(n1064),.dout(w_dff_B_tEIsuwSY6_1),.clk(gclk));
	jdff dff_B_7D12UUX70_2(.din(n964),.dout(w_dff_B_7D12UUX70_2),.clk(gclk));
	jdff dff_B_eHnnMSzG1_2(.din(w_dff_B_7D12UUX70_2),.dout(w_dff_B_eHnnMSzG1_2),.clk(gclk));
	jdff dff_B_S24SvMsw7_2(.din(w_dff_B_eHnnMSzG1_2),.dout(w_dff_B_S24SvMsw7_2),.clk(gclk));
	jdff dff_B_345aMDvI1_2(.din(w_dff_B_S24SvMsw7_2),.dout(w_dff_B_345aMDvI1_2),.clk(gclk));
	jdff dff_B_oLj4Ws795_2(.din(w_dff_B_345aMDvI1_2),.dout(w_dff_B_oLj4Ws795_2),.clk(gclk));
	jdff dff_B_bq8Tivif7_2(.din(w_dff_B_oLj4Ws795_2),.dout(w_dff_B_bq8Tivif7_2),.clk(gclk));
	jdff dff_B_PKtjp3DY0_2(.din(w_dff_B_bq8Tivif7_2),.dout(w_dff_B_PKtjp3DY0_2),.clk(gclk));
	jdff dff_B_D8Aa3MQq6_2(.din(w_dff_B_PKtjp3DY0_2),.dout(w_dff_B_D8Aa3MQq6_2),.clk(gclk));
	jdff dff_B_kwYhMsJa9_2(.din(w_dff_B_D8Aa3MQq6_2),.dout(w_dff_B_kwYhMsJa9_2),.clk(gclk));
	jdff dff_B_ShhZK4Dh8_2(.din(w_dff_B_kwYhMsJa9_2),.dout(w_dff_B_ShhZK4Dh8_2),.clk(gclk));
	jdff dff_B_BrJCwibb1_2(.din(w_dff_B_ShhZK4Dh8_2),.dout(w_dff_B_BrJCwibb1_2),.clk(gclk));
	jdff dff_B_R3ndHCbo9_2(.din(w_dff_B_BrJCwibb1_2),.dout(w_dff_B_R3ndHCbo9_2),.clk(gclk));
	jdff dff_B_YR6wcwMd9_2(.din(w_dff_B_R3ndHCbo9_2),.dout(w_dff_B_YR6wcwMd9_2),.clk(gclk));
	jdff dff_B_0qnDpiRu7_2(.din(w_dff_B_YR6wcwMd9_2),.dout(w_dff_B_0qnDpiRu7_2),.clk(gclk));
	jdff dff_B_8aMSco662_2(.din(n988),.dout(w_dff_B_8aMSco662_2),.clk(gclk));
	jdff dff_B_dvYDu3121_1(.din(n965),.dout(w_dff_B_dvYDu3121_1),.clk(gclk));
	jdff dff_B_sGKYpW7A1_2(.din(n862),.dout(w_dff_B_sGKYpW7A1_2),.clk(gclk));
	jdff dff_B_bfIW92sH1_2(.din(w_dff_B_sGKYpW7A1_2),.dout(w_dff_B_bfIW92sH1_2),.clk(gclk));
	jdff dff_B_Fsgw87Dp9_2(.din(w_dff_B_bfIW92sH1_2),.dout(w_dff_B_Fsgw87Dp9_2),.clk(gclk));
	jdff dff_B_9T1ypWOQ6_2(.din(w_dff_B_Fsgw87Dp9_2),.dout(w_dff_B_9T1ypWOQ6_2),.clk(gclk));
	jdff dff_B_OcvriUyv4_2(.din(w_dff_B_9T1ypWOQ6_2),.dout(w_dff_B_OcvriUyv4_2),.clk(gclk));
	jdff dff_B_1L2foCBo2_2(.din(w_dff_B_OcvriUyv4_2),.dout(w_dff_B_1L2foCBo2_2),.clk(gclk));
	jdff dff_B_dbicMcUa1_2(.din(w_dff_B_1L2foCBo2_2),.dout(w_dff_B_dbicMcUa1_2),.clk(gclk));
	jdff dff_B_2INhwtRo7_2(.din(w_dff_B_dbicMcUa1_2),.dout(w_dff_B_2INhwtRo7_2),.clk(gclk));
	jdff dff_B_WjTeDR5t1_2(.din(w_dff_B_2INhwtRo7_2),.dout(w_dff_B_WjTeDR5t1_2),.clk(gclk));
	jdff dff_B_lhZez3Wi3_2(.din(w_dff_B_WjTeDR5t1_2),.dout(w_dff_B_lhZez3Wi3_2),.clk(gclk));
	jdff dff_B_lEt3Fjqo3_2(.din(w_dff_B_lhZez3Wi3_2),.dout(w_dff_B_lEt3Fjqo3_2),.clk(gclk));
	jdff dff_B_Vd6fMmaD0_2(.din(n882),.dout(w_dff_B_Vd6fMmaD0_2),.clk(gclk));
	jdff dff_B_rX2M1cWh8_1(.din(n863),.dout(w_dff_B_rX2M1cWh8_1),.clk(gclk));
	jdff dff_B_c50el4ku7_2(.din(n764),.dout(w_dff_B_c50el4ku7_2),.clk(gclk));
	jdff dff_B_c98Z24RB0_2(.din(w_dff_B_c50el4ku7_2),.dout(w_dff_B_c98Z24RB0_2),.clk(gclk));
	jdff dff_B_h0AshvrR1_2(.din(w_dff_B_c98Z24RB0_2),.dout(w_dff_B_h0AshvrR1_2),.clk(gclk));
	jdff dff_B_Cl50itll5_2(.din(w_dff_B_h0AshvrR1_2),.dout(w_dff_B_Cl50itll5_2),.clk(gclk));
	jdff dff_B_lq4ZSHCx9_2(.din(w_dff_B_Cl50itll5_2),.dout(w_dff_B_lq4ZSHCx9_2),.clk(gclk));
	jdff dff_B_I93lvMkg4_2(.din(w_dff_B_lq4ZSHCx9_2),.dout(w_dff_B_I93lvMkg4_2),.clk(gclk));
	jdff dff_B_oe9DYwCn9_2(.din(w_dff_B_I93lvMkg4_2),.dout(w_dff_B_oe9DYwCn9_2),.clk(gclk));
	jdff dff_B_GURg5o5w9_2(.din(w_dff_B_oe9DYwCn9_2),.dout(w_dff_B_GURg5o5w9_2),.clk(gclk));
	jdff dff_B_VI1NDn6o2_2(.din(n779),.dout(w_dff_B_VI1NDn6o2_2),.clk(gclk));
	jdff dff_B_ifZxfT5A3_2(.din(w_dff_B_VI1NDn6o2_2),.dout(w_dff_B_ifZxfT5A3_2),.clk(gclk));
	jdff dff_B_9WGQxfkY6_2(.din(w_dff_B_ifZxfT5A3_2),.dout(w_dff_B_9WGQxfkY6_2),.clk(gclk));
	jdff dff_B_kuP3yNXd4_1(.din(n765),.dout(w_dff_B_kuP3yNXd4_1),.clk(gclk));
	jdff dff_B_6JvFeimc6_1(.din(w_dff_B_kuP3yNXd4_1),.dout(w_dff_B_6JvFeimc6_1),.clk(gclk));
	jdff dff_B_j4e8ueRL0_2(.din(n674),.dout(w_dff_B_j4e8ueRL0_2),.clk(gclk));
	jdff dff_B_bJXOhhWn9_2(.din(w_dff_B_j4e8ueRL0_2),.dout(w_dff_B_bJXOhhWn9_2),.clk(gclk));
	jdff dff_B_3QPnI6HQ7_2(.din(w_dff_B_bJXOhhWn9_2),.dout(w_dff_B_3QPnI6HQ7_2),.clk(gclk));
	jdff dff_B_P53qelmo0_0(.din(n679),.dout(w_dff_B_P53qelmo0_0),.clk(gclk));
	jdff dff_A_46UlZCZ00_0(.dout(w_n586_0[0]),.din(w_dff_A_46UlZCZ00_0),.clk(gclk));
	jdff dff_A_Y85roqRL0_0(.dout(w_dff_A_46UlZCZ00_0),.din(w_dff_A_Y85roqRL0_0),.clk(gclk));
	jdff dff_A_c6VNpxpW0_1(.dout(w_n586_0[1]),.din(w_dff_A_c6VNpxpW0_1),.clk(gclk));
	jdff dff_A_as2XVWPH6_1(.dout(w_dff_A_c6VNpxpW0_1),.din(w_dff_A_as2XVWPH6_1),.clk(gclk));
	jdff dff_B_IuxRMeHR7_1(.din(n1788),.dout(w_dff_B_IuxRMeHR7_1),.clk(gclk));
	jdff dff_A_XICyd0S42_1(.dout(w_n1770_0[1]),.din(w_dff_A_XICyd0S42_1),.clk(gclk));
	jdff dff_B_cNIx8qef4_1(.din(n1768),.dout(w_dff_B_cNIx8qef4_1),.clk(gclk));
	jdff dff_B_5VH3S5KC4_2(.din(n1739),.dout(w_dff_B_5VH3S5KC4_2),.clk(gclk));
	jdff dff_B_eonfFV8u8_2(.din(w_dff_B_5VH3S5KC4_2),.dout(w_dff_B_eonfFV8u8_2),.clk(gclk));
	jdff dff_B_56vQnV2A8_2(.din(w_dff_B_eonfFV8u8_2),.dout(w_dff_B_56vQnV2A8_2),.clk(gclk));
	jdff dff_B_eO0lWiz65_2(.din(w_dff_B_56vQnV2A8_2),.dout(w_dff_B_eO0lWiz65_2),.clk(gclk));
	jdff dff_B_oC8nM5Yi5_2(.din(w_dff_B_eO0lWiz65_2),.dout(w_dff_B_oC8nM5Yi5_2),.clk(gclk));
	jdff dff_B_vwgx5DcS3_2(.din(w_dff_B_oC8nM5Yi5_2),.dout(w_dff_B_vwgx5DcS3_2),.clk(gclk));
	jdff dff_B_fFVJZIG67_2(.din(w_dff_B_vwgx5DcS3_2),.dout(w_dff_B_fFVJZIG67_2),.clk(gclk));
	jdff dff_B_d4FGOjfo9_2(.din(w_dff_B_fFVJZIG67_2),.dout(w_dff_B_d4FGOjfo9_2),.clk(gclk));
	jdff dff_B_UILQIAy54_2(.din(w_dff_B_d4FGOjfo9_2),.dout(w_dff_B_UILQIAy54_2),.clk(gclk));
	jdff dff_B_KoF4gMht1_2(.din(w_dff_B_UILQIAy54_2),.dout(w_dff_B_KoF4gMht1_2),.clk(gclk));
	jdff dff_B_Wn5ugI7L7_2(.din(w_dff_B_KoF4gMht1_2),.dout(w_dff_B_Wn5ugI7L7_2),.clk(gclk));
	jdff dff_B_rjqHnoJX9_2(.din(w_dff_B_Wn5ugI7L7_2),.dout(w_dff_B_rjqHnoJX9_2),.clk(gclk));
	jdff dff_B_n6GBJcvL2_2(.din(w_dff_B_rjqHnoJX9_2),.dout(w_dff_B_n6GBJcvL2_2),.clk(gclk));
	jdff dff_B_Dt4sJqKx5_2(.din(w_dff_B_n6GBJcvL2_2),.dout(w_dff_B_Dt4sJqKx5_2),.clk(gclk));
	jdff dff_B_BJI9yP0M9_2(.din(w_dff_B_Dt4sJqKx5_2),.dout(w_dff_B_BJI9yP0M9_2),.clk(gclk));
	jdff dff_B_vrLlW9cl6_2(.din(w_dff_B_BJI9yP0M9_2),.dout(w_dff_B_vrLlW9cl6_2),.clk(gclk));
	jdff dff_B_3LRHKtQS9_2(.din(w_dff_B_vrLlW9cl6_2),.dout(w_dff_B_3LRHKtQS9_2),.clk(gclk));
	jdff dff_B_aCKGDVyq4_2(.din(w_dff_B_3LRHKtQS9_2),.dout(w_dff_B_aCKGDVyq4_2),.clk(gclk));
	jdff dff_B_ORugJqgg6_2(.din(w_dff_B_aCKGDVyq4_2),.dout(w_dff_B_ORugJqgg6_2),.clk(gclk));
	jdff dff_B_5efZ3p6X7_2(.din(w_dff_B_ORugJqgg6_2),.dout(w_dff_B_5efZ3p6X7_2),.clk(gclk));
	jdff dff_B_UwK4YVAB1_2(.din(w_dff_B_5efZ3p6X7_2),.dout(w_dff_B_UwK4YVAB1_2),.clk(gclk));
	jdff dff_B_euxLNvD36_2(.din(w_dff_B_UwK4YVAB1_2),.dout(w_dff_B_euxLNvD36_2),.clk(gclk));
	jdff dff_B_Dd2Sk7f24_2(.din(w_dff_B_euxLNvD36_2),.dout(w_dff_B_Dd2Sk7f24_2),.clk(gclk));
	jdff dff_B_LVENd3dJ2_2(.din(w_dff_B_Dd2Sk7f24_2),.dout(w_dff_B_LVENd3dJ2_2),.clk(gclk));
	jdff dff_B_73vxsRqY7_2(.din(w_dff_B_LVENd3dJ2_2),.dout(w_dff_B_73vxsRqY7_2),.clk(gclk));
	jdff dff_B_lwlF5osT4_2(.din(w_dff_B_73vxsRqY7_2),.dout(w_dff_B_lwlF5osT4_2),.clk(gclk));
	jdff dff_B_E2oGo5wO3_2(.din(w_dff_B_lwlF5osT4_2),.dout(w_dff_B_E2oGo5wO3_2),.clk(gclk));
	jdff dff_B_0ECbxJA31_2(.din(w_dff_B_E2oGo5wO3_2),.dout(w_dff_B_0ECbxJA31_2),.clk(gclk));
	jdff dff_B_X4oyjOEb6_2(.din(w_dff_B_0ECbxJA31_2),.dout(w_dff_B_X4oyjOEb6_2),.clk(gclk));
	jdff dff_B_mhVll2lE1_2(.din(w_dff_B_X4oyjOEb6_2),.dout(w_dff_B_mhVll2lE1_2),.clk(gclk));
	jdff dff_B_f6oVvfJU1_2(.din(w_dff_B_mhVll2lE1_2),.dout(w_dff_B_f6oVvfJU1_2),.clk(gclk));
	jdff dff_B_kyuORWib9_2(.din(w_dff_B_f6oVvfJU1_2),.dout(w_dff_B_kyuORWib9_2),.clk(gclk));
	jdff dff_B_xPcuBZK88_2(.din(w_dff_B_kyuORWib9_2),.dout(w_dff_B_xPcuBZK88_2),.clk(gclk));
	jdff dff_B_5PC7VOl03_2(.din(w_dff_B_xPcuBZK88_2),.dout(w_dff_B_5PC7VOl03_2),.clk(gclk));
	jdff dff_B_u6CBGsXu3_2(.din(w_dff_B_5PC7VOl03_2),.dout(w_dff_B_u6CBGsXu3_2),.clk(gclk));
	jdff dff_B_Jd60A3Jd8_2(.din(w_dff_B_u6CBGsXu3_2),.dout(w_dff_B_Jd60A3Jd8_2),.clk(gclk));
	jdff dff_B_4ugWdidr7_2(.din(w_dff_B_Jd60A3Jd8_2),.dout(w_dff_B_4ugWdidr7_2),.clk(gclk));
	jdff dff_B_Wv25tivg8_2(.din(w_dff_B_4ugWdidr7_2),.dout(w_dff_B_Wv25tivg8_2),.clk(gclk));
	jdff dff_B_Fcmq35nS5_2(.din(w_dff_B_Wv25tivg8_2),.dout(w_dff_B_Fcmq35nS5_2),.clk(gclk));
	jdff dff_B_6bRSeZ6Y0_2(.din(w_dff_B_Fcmq35nS5_2),.dout(w_dff_B_6bRSeZ6Y0_2),.clk(gclk));
	jdff dff_B_k9zFCfFa8_2(.din(w_dff_B_6bRSeZ6Y0_2),.dout(w_dff_B_k9zFCfFa8_2),.clk(gclk));
	jdff dff_B_UIxhGLUA5_2(.din(w_dff_B_k9zFCfFa8_2),.dout(w_dff_B_UIxhGLUA5_2),.clk(gclk));
	jdff dff_B_eTtUuq7z1_2(.din(w_dff_B_UIxhGLUA5_2),.dout(w_dff_B_eTtUuq7z1_2),.clk(gclk));
	jdff dff_B_eG0Dg59U6_2(.din(w_dff_B_eTtUuq7z1_2),.dout(w_dff_B_eG0Dg59U6_2),.clk(gclk));
	jdff dff_B_QtGIqCeq3_2(.din(w_dff_B_eG0Dg59U6_2),.dout(w_dff_B_QtGIqCeq3_2),.clk(gclk));
	jdff dff_B_Vd1YzWeS3_2(.din(w_dff_B_QtGIqCeq3_2),.dout(w_dff_B_Vd1YzWeS3_2),.clk(gclk));
	jdff dff_B_Eq8KXynb3_2(.din(w_dff_B_Vd1YzWeS3_2),.dout(w_dff_B_Eq8KXynb3_2),.clk(gclk));
	jdff dff_B_42Kb9K9Y3_2(.din(w_dff_B_Eq8KXynb3_2),.dout(w_dff_B_42Kb9K9Y3_2),.clk(gclk));
	jdff dff_B_wOQWxcFM9_2(.din(w_dff_B_42Kb9K9Y3_2),.dout(w_dff_B_wOQWxcFM9_2),.clk(gclk));
	jdff dff_B_kZfnxLQn1_2(.din(w_dff_B_wOQWxcFM9_2),.dout(w_dff_B_kZfnxLQn1_2),.clk(gclk));
	jdff dff_B_XI9aL1kA6_2(.din(n1742),.dout(w_dff_B_XI9aL1kA6_2),.clk(gclk));
	jdff dff_B_YZ2J9A3L8_1(.din(n1740),.dout(w_dff_B_YZ2J9A3L8_1),.clk(gclk));
	jdff dff_B_qmakESc91_2(.din(n1704),.dout(w_dff_B_qmakESc91_2),.clk(gclk));
	jdff dff_B_eu2GnKC27_2(.din(w_dff_B_qmakESc91_2),.dout(w_dff_B_eu2GnKC27_2),.clk(gclk));
	jdff dff_B_PwLcmGNU4_2(.din(w_dff_B_eu2GnKC27_2),.dout(w_dff_B_PwLcmGNU4_2),.clk(gclk));
	jdff dff_B_WAsqVksa8_2(.din(w_dff_B_PwLcmGNU4_2),.dout(w_dff_B_WAsqVksa8_2),.clk(gclk));
	jdff dff_B_6WIRJcBQ2_2(.din(w_dff_B_WAsqVksa8_2),.dout(w_dff_B_6WIRJcBQ2_2),.clk(gclk));
	jdff dff_B_BhEidsID0_2(.din(w_dff_B_6WIRJcBQ2_2),.dout(w_dff_B_BhEidsID0_2),.clk(gclk));
	jdff dff_B_GbCx0CF75_2(.din(w_dff_B_BhEidsID0_2),.dout(w_dff_B_GbCx0CF75_2),.clk(gclk));
	jdff dff_B_PLhHUix31_2(.din(w_dff_B_GbCx0CF75_2),.dout(w_dff_B_PLhHUix31_2),.clk(gclk));
	jdff dff_B_Gu0HUX2A1_2(.din(w_dff_B_PLhHUix31_2),.dout(w_dff_B_Gu0HUX2A1_2),.clk(gclk));
	jdff dff_B_Sn5Vhz4B5_2(.din(w_dff_B_Gu0HUX2A1_2),.dout(w_dff_B_Sn5Vhz4B5_2),.clk(gclk));
	jdff dff_B_FuwVTXdU6_2(.din(w_dff_B_Sn5Vhz4B5_2),.dout(w_dff_B_FuwVTXdU6_2),.clk(gclk));
	jdff dff_B_1rVF39iu2_2(.din(w_dff_B_FuwVTXdU6_2),.dout(w_dff_B_1rVF39iu2_2),.clk(gclk));
	jdff dff_B_KsixzHA04_2(.din(w_dff_B_1rVF39iu2_2),.dout(w_dff_B_KsixzHA04_2),.clk(gclk));
	jdff dff_B_fYltOazL9_2(.din(w_dff_B_KsixzHA04_2),.dout(w_dff_B_fYltOazL9_2),.clk(gclk));
	jdff dff_B_GK1aQCcu0_2(.din(w_dff_B_fYltOazL9_2),.dout(w_dff_B_GK1aQCcu0_2),.clk(gclk));
	jdff dff_B_eMqGJ8F13_2(.din(w_dff_B_GK1aQCcu0_2),.dout(w_dff_B_eMqGJ8F13_2),.clk(gclk));
	jdff dff_B_3zEYds2h1_2(.din(w_dff_B_eMqGJ8F13_2),.dout(w_dff_B_3zEYds2h1_2),.clk(gclk));
	jdff dff_B_gcFnD3vg5_2(.din(w_dff_B_3zEYds2h1_2),.dout(w_dff_B_gcFnD3vg5_2),.clk(gclk));
	jdff dff_B_rgjRzDTl7_2(.din(w_dff_B_gcFnD3vg5_2),.dout(w_dff_B_rgjRzDTl7_2),.clk(gclk));
	jdff dff_B_FGUL7rSd9_2(.din(w_dff_B_rgjRzDTl7_2),.dout(w_dff_B_FGUL7rSd9_2),.clk(gclk));
	jdff dff_B_AE4XgTMc7_2(.din(w_dff_B_FGUL7rSd9_2),.dout(w_dff_B_AE4XgTMc7_2),.clk(gclk));
	jdff dff_B_OpgnOYYm3_2(.din(w_dff_B_AE4XgTMc7_2),.dout(w_dff_B_OpgnOYYm3_2),.clk(gclk));
	jdff dff_B_GLwLq8Om5_2(.din(w_dff_B_OpgnOYYm3_2),.dout(w_dff_B_GLwLq8Om5_2),.clk(gclk));
	jdff dff_B_8IGFw4n75_2(.din(w_dff_B_GLwLq8Om5_2),.dout(w_dff_B_8IGFw4n75_2),.clk(gclk));
	jdff dff_B_o3nhPfho0_2(.din(w_dff_B_8IGFw4n75_2),.dout(w_dff_B_o3nhPfho0_2),.clk(gclk));
	jdff dff_B_aBT5OuNh7_2(.din(w_dff_B_o3nhPfho0_2),.dout(w_dff_B_aBT5OuNh7_2),.clk(gclk));
	jdff dff_B_NS0kfxfQ2_2(.din(w_dff_B_aBT5OuNh7_2),.dout(w_dff_B_NS0kfxfQ2_2),.clk(gclk));
	jdff dff_B_emF6X8te7_2(.din(w_dff_B_NS0kfxfQ2_2),.dout(w_dff_B_emF6X8te7_2),.clk(gclk));
	jdff dff_B_s1XKdGf11_2(.din(w_dff_B_emF6X8te7_2),.dout(w_dff_B_s1XKdGf11_2),.clk(gclk));
	jdff dff_B_t5twnAwt4_2(.din(w_dff_B_s1XKdGf11_2),.dout(w_dff_B_t5twnAwt4_2),.clk(gclk));
	jdff dff_B_RWA8z1rd4_2(.din(w_dff_B_t5twnAwt4_2),.dout(w_dff_B_RWA8z1rd4_2),.clk(gclk));
	jdff dff_B_tGQ1HdrO5_2(.din(w_dff_B_RWA8z1rd4_2),.dout(w_dff_B_tGQ1HdrO5_2),.clk(gclk));
	jdff dff_B_cnVcqDy19_2(.din(w_dff_B_tGQ1HdrO5_2),.dout(w_dff_B_cnVcqDy19_2),.clk(gclk));
	jdff dff_B_YcoEt3Rc4_2(.din(w_dff_B_cnVcqDy19_2),.dout(w_dff_B_YcoEt3Rc4_2),.clk(gclk));
	jdff dff_B_Ke7e9Ui86_2(.din(w_dff_B_YcoEt3Rc4_2),.dout(w_dff_B_Ke7e9Ui86_2),.clk(gclk));
	jdff dff_B_8OtDWy1P2_2(.din(w_dff_B_Ke7e9Ui86_2),.dout(w_dff_B_8OtDWy1P2_2),.clk(gclk));
	jdff dff_B_sG4f9neP9_2(.din(w_dff_B_8OtDWy1P2_2),.dout(w_dff_B_sG4f9neP9_2),.clk(gclk));
	jdff dff_B_JRXAlELz5_2(.din(w_dff_B_sG4f9neP9_2),.dout(w_dff_B_JRXAlELz5_2),.clk(gclk));
	jdff dff_B_XoZAkpvS4_2(.din(w_dff_B_JRXAlELz5_2),.dout(w_dff_B_XoZAkpvS4_2),.clk(gclk));
	jdff dff_B_LWMAvW8f8_2(.din(w_dff_B_XoZAkpvS4_2),.dout(w_dff_B_LWMAvW8f8_2),.clk(gclk));
	jdff dff_B_32XNziaG7_2(.din(w_dff_B_LWMAvW8f8_2),.dout(w_dff_B_32XNziaG7_2),.clk(gclk));
	jdff dff_B_zULAgVPI8_2(.din(w_dff_B_32XNziaG7_2),.dout(w_dff_B_zULAgVPI8_2),.clk(gclk));
	jdff dff_B_Dc2eUq571_2(.din(w_dff_B_zULAgVPI8_2),.dout(w_dff_B_Dc2eUq571_2),.clk(gclk));
	jdff dff_B_9yEx8lTI4_2(.din(w_dff_B_Dc2eUq571_2),.dout(w_dff_B_9yEx8lTI4_2),.clk(gclk));
	jdff dff_B_7wcgc0jE1_2(.din(w_dff_B_9yEx8lTI4_2),.dout(w_dff_B_7wcgc0jE1_2),.clk(gclk));
	jdff dff_B_R2b2iea10_2(.din(w_dff_B_7wcgc0jE1_2),.dout(w_dff_B_R2b2iea10_2),.clk(gclk));
	jdff dff_B_9JNkZehn3_2(.din(n1707),.dout(w_dff_B_9JNkZehn3_2),.clk(gclk));
	jdff dff_B_qIxe3vd75_1(.din(n1705),.dout(w_dff_B_qIxe3vd75_1),.clk(gclk));
	jdff dff_B_NVfbZG8w5_2(.din(n1663),.dout(w_dff_B_NVfbZG8w5_2),.clk(gclk));
	jdff dff_B_q31nTGiS3_2(.din(w_dff_B_NVfbZG8w5_2),.dout(w_dff_B_q31nTGiS3_2),.clk(gclk));
	jdff dff_B_yj1Oysll0_2(.din(w_dff_B_q31nTGiS3_2),.dout(w_dff_B_yj1Oysll0_2),.clk(gclk));
	jdff dff_B_NNh7bi0w6_2(.din(w_dff_B_yj1Oysll0_2),.dout(w_dff_B_NNh7bi0w6_2),.clk(gclk));
	jdff dff_B_OMaqo4Ru2_2(.din(w_dff_B_NNh7bi0w6_2),.dout(w_dff_B_OMaqo4Ru2_2),.clk(gclk));
	jdff dff_B_XHID7XCf1_2(.din(w_dff_B_OMaqo4Ru2_2),.dout(w_dff_B_XHID7XCf1_2),.clk(gclk));
	jdff dff_B_MOkMZ7Md9_2(.din(w_dff_B_XHID7XCf1_2),.dout(w_dff_B_MOkMZ7Md9_2),.clk(gclk));
	jdff dff_B_s9qYIOlf6_2(.din(w_dff_B_MOkMZ7Md9_2),.dout(w_dff_B_s9qYIOlf6_2),.clk(gclk));
	jdff dff_B_9wN18sTM0_2(.din(w_dff_B_s9qYIOlf6_2),.dout(w_dff_B_9wN18sTM0_2),.clk(gclk));
	jdff dff_B_nAWgq8vi1_2(.din(w_dff_B_9wN18sTM0_2),.dout(w_dff_B_nAWgq8vi1_2),.clk(gclk));
	jdff dff_B_ZGYvdwqG6_2(.din(w_dff_B_nAWgq8vi1_2),.dout(w_dff_B_ZGYvdwqG6_2),.clk(gclk));
	jdff dff_B_BwM7BUln4_2(.din(w_dff_B_ZGYvdwqG6_2),.dout(w_dff_B_BwM7BUln4_2),.clk(gclk));
	jdff dff_B_3DYt0mkP2_2(.din(w_dff_B_BwM7BUln4_2),.dout(w_dff_B_3DYt0mkP2_2),.clk(gclk));
	jdff dff_B_TjitmiLP6_2(.din(w_dff_B_3DYt0mkP2_2),.dout(w_dff_B_TjitmiLP6_2),.clk(gclk));
	jdff dff_B_B6KatWc69_2(.din(w_dff_B_TjitmiLP6_2),.dout(w_dff_B_B6KatWc69_2),.clk(gclk));
	jdff dff_B_jJyY4cTE7_2(.din(w_dff_B_B6KatWc69_2),.dout(w_dff_B_jJyY4cTE7_2),.clk(gclk));
	jdff dff_B_ZDJN93Bu5_2(.din(w_dff_B_jJyY4cTE7_2),.dout(w_dff_B_ZDJN93Bu5_2),.clk(gclk));
	jdff dff_B_4ybuubSP4_2(.din(w_dff_B_ZDJN93Bu5_2),.dout(w_dff_B_4ybuubSP4_2),.clk(gclk));
	jdff dff_B_qYAC7WbY1_2(.din(w_dff_B_4ybuubSP4_2),.dout(w_dff_B_qYAC7WbY1_2),.clk(gclk));
	jdff dff_B_HYOiJHHU0_2(.din(w_dff_B_qYAC7WbY1_2),.dout(w_dff_B_HYOiJHHU0_2),.clk(gclk));
	jdff dff_B_slKoBVAO3_2(.din(w_dff_B_HYOiJHHU0_2),.dout(w_dff_B_slKoBVAO3_2),.clk(gclk));
	jdff dff_B_v73g2qe33_2(.din(w_dff_B_slKoBVAO3_2),.dout(w_dff_B_v73g2qe33_2),.clk(gclk));
	jdff dff_B_RRwZcDg88_2(.din(w_dff_B_v73g2qe33_2),.dout(w_dff_B_RRwZcDg88_2),.clk(gclk));
	jdff dff_B_v7PMVfU24_2(.din(w_dff_B_RRwZcDg88_2),.dout(w_dff_B_v7PMVfU24_2),.clk(gclk));
	jdff dff_B_Ig3GQaC66_2(.din(w_dff_B_v7PMVfU24_2),.dout(w_dff_B_Ig3GQaC66_2),.clk(gclk));
	jdff dff_B_UH5SJ1ty1_2(.din(w_dff_B_Ig3GQaC66_2),.dout(w_dff_B_UH5SJ1ty1_2),.clk(gclk));
	jdff dff_B_gbY1j1Mp7_2(.din(w_dff_B_UH5SJ1ty1_2),.dout(w_dff_B_gbY1j1Mp7_2),.clk(gclk));
	jdff dff_B_Nan30Hjt2_2(.din(w_dff_B_gbY1j1Mp7_2),.dout(w_dff_B_Nan30Hjt2_2),.clk(gclk));
	jdff dff_B_9PByZS5W8_2(.din(w_dff_B_Nan30Hjt2_2),.dout(w_dff_B_9PByZS5W8_2),.clk(gclk));
	jdff dff_B_qwSj470X6_2(.din(w_dff_B_9PByZS5W8_2),.dout(w_dff_B_qwSj470X6_2),.clk(gclk));
	jdff dff_B_9MKSPDSP3_2(.din(w_dff_B_qwSj470X6_2),.dout(w_dff_B_9MKSPDSP3_2),.clk(gclk));
	jdff dff_B_u8vTxEML2_2(.din(w_dff_B_9MKSPDSP3_2),.dout(w_dff_B_u8vTxEML2_2),.clk(gclk));
	jdff dff_B_YXpqEmOj2_2(.din(w_dff_B_u8vTxEML2_2),.dout(w_dff_B_YXpqEmOj2_2),.clk(gclk));
	jdff dff_B_9j7eYWqM0_2(.din(w_dff_B_YXpqEmOj2_2),.dout(w_dff_B_9j7eYWqM0_2),.clk(gclk));
	jdff dff_B_I7XImHNI4_2(.din(w_dff_B_9j7eYWqM0_2),.dout(w_dff_B_I7XImHNI4_2),.clk(gclk));
	jdff dff_B_z9Rgkd8u4_2(.din(w_dff_B_I7XImHNI4_2),.dout(w_dff_B_z9Rgkd8u4_2),.clk(gclk));
	jdff dff_B_0pDl5VBX2_2(.din(w_dff_B_z9Rgkd8u4_2),.dout(w_dff_B_0pDl5VBX2_2),.clk(gclk));
	jdff dff_B_ZkHN4mcn7_2(.din(w_dff_B_0pDl5VBX2_2),.dout(w_dff_B_ZkHN4mcn7_2),.clk(gclk));
	jdff dff_B_JfmcWgGP3_2(.din(w_dff_B_ZkHN4mcn7_2),.dout(w_dff_B_JfmcWgGP3_2),.clk(gclk));
	jdff dff_B_R82lrEbb0_2(.din(w_dff_B_JfmcWgGP3_2),.dout(w_dff_B_R82lrEbb0_2),.clk(gclk));
	jdff dff_B_VDz2SiDw3_2(.din(w_dff_B_R82lrEbb0_2),.dout(w_dff_B_VDz2SiDw3_2),.clk(gclk));
	jdff dff_B_QBDy5FYn6_2(.din(w_dff_B_VDz2SiDw3_2),.dout(w_dff_B_QBDy5FYn6_2),.clk(gclk));
	jdff dff_B_uQ6Ji3YS2_2(.din(n1666),.dout(w_dff_B_uQ6Ji3YS2_2),.clk(gclk));
	jdff dff_B_2UH6Sju27_1(.din(n1664),.dout(w_dff_B_2UH6Sju27_1),.clk(gclk));
	jdff dff_B_KPqezL1z7_2(.din(n1612),.dout(w_dff_B_KPqezL1z7_2),.clk(gclk));
	jdff dff_B_LKVCHkt39_2(.din(w_dff_B_KPqezL1z7_2),.dout(w_dff_B_LKVCHkt39_2),.clk(gclk));
	jdff dff_B_Kub1RPoA5_2(.din(w_dff_B_LKVCHkt39_2),.dout(w_dff_B_Kub1RPoA5_2),.clk(gclk));
	jdff dff_B_KxCVWRow4_2(.din(w_dff_B_Kub1RPoA5_2),.dout(w_dff_B_KxCVWRow4_2),.clk(gclk));
	jdff dff_B_CCr9oJcR6_2(.din(w_dff_B_KxCVWRow4_2),.dout(w_dff_B_CCr9oJcR6_2),.clk(gclk));
	jdff dff_B_BgfVez5E5_2(.din(w_dff_B_CCr9oJcR6_2),.dout(w_dff_B_BgfVez5E5_2),.clk(gclk));
	jdff dff_B_JvFE5xG48_2(.din(w_dff_B_BgfVez5E5_2),.dout(w_dff_B_JvFE5xG48_2),.clk(gclk));
	jdff dff_B_wAeifTfD6_2(.din(w_dff_B_JvFE5xG48_2),.dout(w_dff_B_wAeifTfD6_2),.clk(gclk));
	jdff dff_B_r7SEr9GN3_2(.din(w_dff_B_wAeifTfD6_2),.dout(w_dff_B_r7SEr9GN3_2),.clk(gclk));
	jdff dff_B_iWc8oDqp6_2(.din(w_dff_B_r7SEr9GN3_2),.dout(w_dff_B_iWc8oDqp6_2),.clk(gclk));
	jdff dff_B_PjOst9vO6_2(.din(w_dff_B_iWc8oDqp6_2),.dout(w_dff_B_PjOst9vO6_2),.clk(gclk));
	jdff dff_B_KFSz1UYg8_2(.din(w_dff_B_PjOst9vO6_2),.dout(w_dff_B_KFSz1UYg8_2),.clk(gclk));
	jdff dff_B_stk4p4U24_2(.din(w_dff_B_KFSz1UYg8_2),.dout(w_dff_B_stk4p4U24_2),.clk(gclk));
	jdff dff_B_LzvV4MbZ0_2(.din(w_dff_B_stk4p4U24_2),.dout(w_dff_B_LzvV4MbZ0_2),.clk(gclk));
	jdff dff_B_SZIE7ewA0_2(.din(w_dff_B_LzvV4MbZ0_2),.dout(w_dff_B_SZIE7ewA0_2),.clk(gclk));
	jdff dff_B_PSpzbNGq7_2(.din(w_dff_B_SZIE7ewA0_2),.dout(w_dff_B_PSpzbNGq7_2),.clk(gclk));
	jdff dff_B_6wEnHQ3O8_2(.din(w_dff_B_PSpzbNGq7_2),.dout(w_dff_B_6wEnHQ3O8_2),.clk(gclk));
	jdff dff_B_9rBjxFsq1_2(.din(w_dff_B_6wEnHQ3O8_2),.dout(w_dff_B_9rBjxFsq1_2),.clk(gclk));
	jdff dff_B_3QJIp8YZ9_2(.din(w_dff_B_9rBjxFsq1_2),.dout(w_dff_B_3QJIp8YZ9_2),.clk(gclk));
	jdff dff_B_Yjt6tcos6_2(.din(w_dff_B_3QJIp8YZ9_2),.dout(w_dff_B_Yjt6tcos6_2),.clk(gclk));
	jdff dff_B_nc5pdmiF8_2(.din(w_dff_B_Yjt6tcos6_2),.dout(w_dff_B_nc5pdmiF8_2),.clk(gclk));
	jdff dff_B_QDHaZHBr1_2(.din(w_dff_B_nc5pdmiF8_2),.dout(w_dff_B_QDHaZHBr1_2),.clk(gclk));
	jdff dff_B_g9QSn8kA9_2(.din(w_dff_B_QDHaZHBr1_2),.dout(w_dff_B_g9QSn8kA9_2),.clk(gclk));
	jdff dff_B_zzJ2wYow2_2(.din(w_dff_B_g9QSn8kA9_2),.dout(w_dff_B_zzJ2wYow2_2),.clk(gclk));
	jdff dff_B_xJW8AOW98_2(.din(w_dff_B_zzJ2wYow2_2),.dout(w_dff_B_xJW8AOW98_2),.clk(gclk));
	jdff dff_B_YLOkRTk84_2(.din(w_dff_B_xJW8AOW98_2),.dout(w_dff_B_YLOkRTk84_2),.clk(gclk));
	jdff dff_B_c8afeDPF4_2(.din(w_dff_B_YLOkRTk84_2),.dout(w_dff_B_c8afeDPF4_2),.clk(gclk));
	jdff dff_B_6qhEYN629_2(.din(w_dff_B_c8afeDPF4_2),.dout(w_dff_B_6qhEYN629_2),.clk(gclk));
	jdff dff_B_8L7B1R8z3_2(.din(w_dff_B_6qhEYN629_2),.dout(w_dff_B_8L7B1R8z3_2),.clk(gclk));
	jdff dff_B_MvYxJbrD3_2(.din(w_dff_B_8L7B1R8z3_2),.dout(w_dff_B_MvYxJbrD3_2),.clk(gclk));
	jdff dff_B_0hN6HVNw3_2(.din(w_dff_B_MvYxJbrD3_2),.dout(w_dff_B_0hN6HVNw3_2),.clk(gclk));
	jdff dff_B_MjmfVJrZ1_2(.din(w_dff_B_0hN6HVNw3_2),.dout(w_dff_B_MjmfVJrZ1_2),.clk(gclk));
	jdff dff_B_ybvTQLDj6_2(.din(w_dff_B_MjmfVJrZ1_2),.dout(w_dff_B_ybvTQLDj6_2),.clk(gclk));
	jdff dff_B_NBui3msE9_2(.din(w_dff_B_ybvTQLDj6_2),.dout(w_dff_B_NBui3msE9_2),.clk(gclk));
	jdff dff_B_b7o55a3V5_2(.din(w_dff_B_NBui3msE9_2),.dout(w_dff_B_b7o55a3V5_2),.clk(gclk));
	jdff dff_B_bYHH4Yfc8_2(.din(w_dff_B_b7o55a3V5_2),.dout(w_dff_B_bYHH4Yfc8_2),.clk(gclk));
	jdff dff_B_N9AL9DrK6_2(.din(w_dff_B_bYHH4Yfc8_2),.dout(w_dff_B_N9AL9DrK6_2),.clk(gclk));
	jdff dff_B_g4sqGszj0_2(.din(w_dff_B_N9AL9DrK6_2),.dout(w_dff_B_g4sqGszj0_2),.clk(gclk));
	jdff dff_B_YuhbQnDV1_2(.din(n1615),.dout(w_dff_B_YuhbQnDV1_2),.clk(gclk));
	jdff dff_B_QaZA6LOD3_1(.din(n1613),.dout(w_dff_B_QaZA6LOD3_1),.clk(gclk));
	jdff dff_B_RzWB5iSg2_2(.din(n1555),.dout(w_dff_B_RzWB5iSg2_2),.clk(gclk));
	jdff dff_B_NdfeGn7z7_2(.din(w_dff_B_RzWB5iSg2_2),.dout(w_dff_B_NdfeGn7z7_2),.clk(gclk));
	jdff dff_B_I4ubmTIl0_2(.din(w_dff_B_NdfeGn7z7_2),.dout(w_dff_B_I4ubmTIl0_2),.clk(gclk));
	jdff dff_B_iWz0g9oD4_2(.din(w_dff_B_I4ubmTIl0_2),.dout(w_dff_B_iWz0g9oD4_2),.clk(gclk));
	jdff dff_B_CjGinJYp1_2(.din(w_dff_B_iWz0g9oD4_2),.dout(w_dff_B_CjGinJYp1_2),.clk(gclk));
	jdff dff_B_BLnkTZ9F0_2(.din(w_dff_B_CjGinJYp1_2),.dout(w_dff_B_BLnkTZ9F0_2),.clk(gclk));
	jdff dff_B_V1dW6LMn0_2(.din(w_dff_B_BLnkTZ9F0_2),.dout(w_dff_B_V1dW6LMn0_2),.clk(gclk));
	jdff dff_B_UlYrC57j3_2(.din(w_dff_B_V1dW6LMn0_2),.dout(w_dff_B_UlYrC57j3_2),.clk(gclk));
	jdff dff_B_oKIsmv7I1_2(.din(w_dff_B_UlYrC57j3_2),.dout(w_dff_B_oKIsmv7I1_2),.clk(gclk));
	jdff dff_B_s0T3wLst3_2(.din(w_dff_B_oKIsmv7I1_2),.dout(w_dff_B_s0T3wLst3_2),.clk(gclk));
	jdff dff_B_DsevGJRv5_2(.din(w_dff_B_s0T3wLst3_2),.dout(w_dff_B_DsevGJRv5_2),.clk(gclk));
	jdff dff_B_3HG2h4uj7_2(.din(w_dff_B_DsevGJRv5_2),.dout(w_dff_B_3HG2h4uj7_2),.clk(gclk));
	jdff dff_B_bl2F6YaM6_2(.din(w_dff_B_3HG2h4uj7_2),.dout(w_dff_B_bl2F6YaM6_2),.clk(gclk));
	jdff dff_B_jW8y2dBd1_2(.din(w_dff_B_bl2F6YaM6_2),.dout(w_dff_B_jW8y2dBd1_2),.clk(gclk));
	jdff dff_B_XHAP7rNe0_2(.din(w_dff_B_jW8y2dBd1_2),.dout(w_dff_B_XHAP7rNe0_2),.clk(gclk));
	jdff dff_B_j5ZlGhP52_2(.din(w_dff_B_XHAP7rNe0_2),.dout(w_dff_B_j5ZlGhP52_2),.clk(gclk));
	jdff dff_B_7Nc3XTFA8_2(.din(w_dff_B_j5ZlGhP52_2),.dout(w_dff_B_7Nc3XTFA8_2),.clk(gclk));
	jdff dff_B_5TvAHopH4_2(.din(w_dff_B_7Nc3XTFA8_2),.dout(w_dff_B_5TvAHopH4_2),.clk(gclk));
	jdff dff_B_uJ0AlV0R0_2(.din(w_dff_B_5TvAHopH4_2),.dout(w_dff_B_uJ0AlV0R0_2),.clk(gclk));
	jdff dff_B_c1mHGTGw3_2(.din(w_dff_B_uJ0AlV0R0_2),.dout(w_dff_B_c1mHGTGw3_2),.clk(gclk));
	jdff dff_B_P2x1g1VB8_2(.din(w_dff_B_c1mHGTGw3_2),.dout(w_dff_B_P2x1g1VB8_2),.clk(gclk));
	jdff dff_B_T6aPQNht1_2(.din(w_dff_B_P2x1g1VB8_2),.dout(w_dff_B_T6aPQNht1_2),.clk(gclk));
	jdff dff_B_70n6rwZV7_2(.din(w_dff_B_T6aPQNht1_2),.dout(w_dff_B_70n6rwZV7_2),.clk(gclk));
	jdff dff_B_YNZMNGWQ8_2(.din(w_dff_B_70n6rwZV7_2),.dout(w_dff_B_YNZMNGWQ8_2),.clk(gclk));
	jdff dff_B_dDnYqVIC0_2(.din(w_dff_B_YNZMNGWQ8_2),.dout(w_dff_B_dDnYqVIC0_2),.clk(gclk));
	jdff dff_B_LCP5en5G1_2(.din(w_dff_B_dDnYqVIC0_2),.dout(w_dff_B_LCP5en5G1_2),.clk(gclk));
	jdff dff_B_UDmQUMAb0_2(.din(w_dff_B_LCP5en5G1_2),.dout(w_dff_B_UDmQUMAb0_2),.clk(gclk));
	jdff dff_B_1Rf4n2bq3_2(.din(w_dff_B_UDmQUMAb0_2),.dout(w_dff_B_1Rf4n2bq3_2),.clk(gclk));
	jdff dff_B_KQuy6tPL7_2(.din(w_dff_B_1Rf4n2bq3_2),.dout(w_dff_B_KQuy6tPL7_2),.clk(gclk));
	jdff dff_B_2SX8haRQ9_2(.din(w_dff_B_KQuy6tPL7_2),.dout(w_dff_B_2SX8haRQ9_2),.clk(gclk));
	jdff dff_B_kZx66CwO6_2(.din(w_dff_B_2SX8haRQ9_2),.dout(w_dff_B_kZx66CwO6_2),.clk(gclk));
	jdff dff_B_5ix9SUyF4_2(.din(w_dff_B_kZx66CwO6_2),.dout(w_dff_B_5ix9SUyF4_2),.clk(gclk));
	jdff dff_B_g8O4kjua5_2(.din(w_dff_B_5ix9SUyF4_2),.dout(w_dff_B_g8O4kjua5_2),.clk(gclk));
	jdff dff_B_8XvW1uyN8_2(.din(w_dff_B_g8O4kjua5_2),.dout(w_dff_B_8XvW1uyN8_2),.clk(gclk));
	jdff dff_B_mKfxyogV8_2(.din(n1558),.dout(w_dff_B_mKfxyogV8_2),.clk(gclk));
	jdff dff_B_iQ0mUJQH6_1(.din(n1556),.dout(w_dff_B_iQ0mUJQH6_1),.clk(gclk));
	jdff dff_B_dQdqVN723_2(.din(n1491),.dout(w_dff_B_dQdqVN723_2),.clk(gclk));
	jdff dff_B_NTPd2rSh2_2(.din(w_dff_B_dQdqVN723_2),.dout(w_dff_B_NTPd2rSh2_2),.clk(gclk));
	jdff dff_B_zqV67sBM5_2(.din(w_dff_B_NTPd2rSh2_2),.dout(w_dff_B_zqV67sBM5_2),.clk(gclk));
	jdff dff_B_n099u9Pv0_2(.din(w_dff_B_zqV67sBM5_2),.dout(w_dff_B_n099u9Pv0_2),.clk(gclk));
	jdff dff_B_6Sab7Gvb9_2(.din(w_dff_B_n099u9Pv0_2),.dout(w_dff_B_6Sab7Gvb9_2),.clk(gclk));
	jdff dff_B_gLeGkFh78_2(.din(w_dff_B_6Sab7Gvb9_2),.dout(w_dff_B_gLeGkFh78_2),.clk(gclk));
	jdff dff_B_ddkL6cTG5_2(.din(w_dff_B_gLeGkFh78_2),.dout(w_dff_B_ddkL6cTG5_2),.clk(gclk));
	jdff dff_B_XCUWzEbc6_2(.din(w_dff_B_ddkL6cTG5_2),.dout(w_dff_B_XCUWzEbc6_2),.clk(gclk));
	jdff dff_B_UrPrCatm2_2(.din(w_dff_B_XCUWzEbc6_2),.dout(w_dff_B_UrPrCatm2_2),.clk(gclk));
	jdff dff_B_eu3o8Ibq0_2(.din(w_dff_B_UrPrCatm2_2),.dout(w_dff_B_eu3o8Ibq0_2),.clk(gclk));
	jdff dff_B_hzY9z3lZ4_2(.din(w_dff_B_eu3o8Ibq0_2),.dout(w_dff_B_hzY9z3lZ4_2),.clk(gclk));
	jdff dff_B_n2NpeEVV3_2(.din(w_dff_B_hzY9z3lZ4_2),.dout(w_dff_B_n2NpeEVV3_2),.clk(gclk));
	jdff dff_B_mNy4Cxjq4_2(.din(w_dff_B_n2NpeEVV3_2),.dout(w_dff_B_mNy4Cxjq4_2),.clk(gclk));
	jdff dff_B_xZQFpAmx4_2(.din(w_dff_B_mNy4Cxjq4_2),.dout(w_dff_B_xZQFpAmx4_2),.clk(gclk));
	jdff dff_B_HsqbjUEV3_2(.din(w_dff_B_xZQFpAmx4_2),.dout(w_dff_B_HsqbjUEV3_2),.clk(gclk));
	jdff dff_B_wCzqPmun3_2(.din(w_dff_B_HsqbjUEV3_2),.dout(w_dff_B_wCzqPmun3_2),.clk(gclk));
	jdff dff_B_u0zIWOXM2_2(.din(w_dff_B_wCzqPmun3_2),.dout(w_dff_B_u0zIWOXM2_2),.clk(gclk));
	jdff dff_B_UEzWtuxx1_2(.din(w_dff_B_u0zIWOXM2_2),.dout(w_dff_B_UEzWtuxx1_2),.clk(gclk));
	jdff dff_B_O71PxFAS5_2(.din(w_dff_B_UEzWtuxx1_2),.dout(w_dff_B_O71PxFAS5_2),.clk(gclk));
	jdff dff_B_wIaZn0DU1_2(.din(w_dff_B_O71PxFAS5_2),.dout(w_dff_B_wIaZn0DU1_2),.clk(gclk));
	jdff dff_B_s7c5mmix7_2(.din(w_dff_B_wIaZn0DU1_2),.dout(w_dff_B_s7c5mmix7_2),.clk(gclk));
	jdff dff_B_G4522sUc5_2(.din(w_dff_B_s7c5mmix7_2),.dout(w_dff_B_G4522sUc5_2),.clk(gclk));
	jdff dff_B_9Q1p4yba0_2(.din(w_dff_B_G4522sUc5_2),.dout(w_dff_B_9Q1p4yba0_2),.clk(gclk));
	jdff dff_B_jhCC9DdC0_2(.din(w_dff_B_9Q1p4yba0_2),.dout(w_dff_B_jhCC9DdC0_2),.clk(gclk));
	jdff dff_B_c6yzg8PN3_2(.din(w_dff_B_jhCC9DdC0_2),.dout(w_dff_B_c6yzg8PN3_2),.clk(gclk));
	jdff dff_B_LCNauuFj0_2(.din(w_dff_B_c6yzg8PN3_2),.dout(w_dff_B_LCNauuFj0_2),.clk(gclk));
	jdff dff_B_xLJgt0sl3_2(.din(w_dff_B_LCNauuFj0_2),.dout(w_dff_B_xLJgt0sl3_2),.clk(gclk));
	jdff dff_B_jx55aJCp5_2(.din(w_dff_B_xLJgt0sl3_2),.dout(w_dff_B_jx55aJCp5_2),.clk(gclk));
	jdff dff_B_84X8Q3Iq5_2(.din(w_dff_B_jx55aJCp5_2),.dout(w_dff_B_84X8Q3Iq5_2),.clk(gclk));
	jdff dff_B_qrmTfwrb9_2(.din(w_dff_B_84X8Q3Iq5_2),.dout(w_dff_B_qrmTfwrb9_2),.clk(gclk));
	jdff dff_B_KkbJhSEQ3_2(.din(n1494),.dout(w_dff_B_KkbJhSEQ3_2),.clk(gclk));
	jdff dff_B_ho8lWHFt5_1(.din(n1492),.dout(w_dff_B_ho8lWHFt5_1),.clk(gclk));
	jdff dff_B_S58oYmMa0_2(.din(n1420),.dout(w_dff_B_S58oYmMa0_2),.clk(gclk));
	jdff dff_B_IKGTS3zP1_2(.din(w_dff_B_S58oYmMa0_2),.dout(w_dff_B_IKGTS3zP1_2),.clk(gclk));
	jdff dff_B_DUCn5t4Q7_2(.din(w_dff_B_IKGTS3zP1_2),.dout(w_dff_B_DUCn5t4Q7_2),.clk(gclk));
	jdff dff_B_1MiFA5151_2(.din(w_dff_B_DUCn5t4Q7_2),.dout(w_dff_B_1MiFA5151_2),.clk(gclk));
	jdff dff_B_C6Zyxbbl3_2(.din(w_dff_B_1MiFA5151_2),.dout(w_dff_B_C6Zyxbbl3_2),.clk(gclk));
	jdff dff_B_ZGPI2EY02_2(.din(w_dff_B_C6Zyxbbl3_2),.dout(w_dff_B_ZGPI2EY02_2),.clk(gclk));
	jdff dff_B_DkH4Sp0K4_2(.din(w_dff_B_ZGPI2EY02_2),.dout(w_dff_B_DkH4Sp0K4_2),.clk(gclk));
	jdff dff_B_BciaIpX67_2(.din(w_dff_B_DkH4Sp0K4_2),.dout(w_dff_B_BciaIpX67_2),.clk(gclk));
	jdff dff_B_hPADyZlN8_2(.din(w_dff_B_BciaIpX67_2),.dout(w_dff_B_hPADyZlN8_2),.clk(gclk));
	jdff dff_B_uN7n0fjF1_2(.din(w_dff_B_hPADyZlN8_2),.dout(w_dff_B_uN7n0fjF1_2),.clk(gclk));
	jdff dff_B_LEEUnOa70_2(.din(w_dff_B_uN7n0fjF1_2),.dout(w_dff_B_LEEUnOa70_2),.clk(gclk));
	jdff dff_B_KhVTjsAB2_2(.din(w_dff_B_LEEUnOa70_2),.dout(w_dff_B_KhVTjsAB2_2),.clk(gclk));
	jdff dff_B_GcII21Rg3_2(.din(w_dff_B_KhVTjsAB2_2),.dout(w_dff_B_GcII21Rg3_2),.clk(gclk));
	jdff dff_B_U71n6pbz7_2(.din(w_dff_B_GcII21Rg3_2),.dout(w_dff_B_U71n6pbz7_2),.clk(gclk));
	jdff dff_B_XulHHwSR3_2(.din(w_dff_B_U71n6pbz7_2),.dout(w_dff_B_XulHHwSR3_2),.clk(gclk));
	jdff dff_B_KpREJOeS1_2(.din(w_dff_B_XulHHwSR3_2),.dout(w_dff_B_KpREJOeS1_2),.clk(gclk));
	jdff dff_B_jTA3M3jC7_2(.din(w_dff_B_KpREJOeS1_2),.dout(w_dff_B_jTA3M3jC7_2),.clk(gclk));
	jdff dff_B_vyF548bN1_2(.din(w_dff_B_jTA3M3jC7_2),.dout(w_dff_B_vyF548bN1_2),.clk(gclk));
	jdff dff_B_OMv3a6iv1_2(.din(w_dff_B_vyF548bN1_2),.dout(w_dff_B_OMv3a6iv1_2),.clk(gclk));
	jdff dff_B_Z8u58FAa3_2(.din(w_dff_B_OMv3a6iv1_2),.dout(w_dff_B_Z8u58FAa3_2),.clk(gclk));
	jdff dff_B_5p5T4rIz2_2(.din(w_dff_B_Z8u58FAa3_2),.dout(w_dff_B_5p5T4rIz2_2),.clk(gclk));
	jdff dff_B_vtpdGxVm4_2(.din(w_dff_B_5p5T4rIz2_2),.dout(w_dff_B_vtpdGxVm4_2),.clk(gclk));
	jdff dff_B_KMI7p34y5_2(.din(w_dff_B_vtpdGxVm4_2),.dout(w_dff_B_KMI7p34y5_2),.clk(gclk));
	jdff dff_B_QH1yS4HV2_2(.din(w_dff_B_KMI7p34y5_2),.dout(w_dff_B_QH1yS4HV2_2),.clk(gclk));
	jdff dff_B_AHxknJIR7_2(.din(w_dff_B_QH1yS4HV2_2),.dout(w_dff_B_AHxknJIR7_2),.clk(gclk));
	jdff dff_B_1BL8Ahqj1_2(.din(w_dff_B_AHxknJIR7_2),.dout(w_dff_B_1BL8Ahqj1_2),.clk(gclk));
	jdff dff_B_XCPKuwD08_1(.din(n1421),.dout(w_dff_B_XCPKuwD08_1),.clk(gclk));
	jdff dff_B_8fWD4FDZ5_2(.din(n1342),.dout(w_dff_B_8fWD4FDZ5_2),.clk(gclk));
	jdff dff_B_0bmhFsBP2_2(.din(w_dff_B_8fWD4FDZ5_2),.dout(w_dff_B_0bmhFsBP2_2),.clk(gclk));
	jdff dff_B_L8tmRKeS6_2(.din(w_dff_B_0bmhFsBP2_2),.dout(w_dff_B_L8tmRKeS6_2),.clk(gclk));
	jdff dff_B_Zq0PgvtI0_2(.din(w_dff_B_L8tmRKeS6_2),.dout(w_dff_B_Zq0PgvtI0_2),.clk(gclk));
	jdff dff_B_bh9e0hKE9_2(.din(w_dff_B_Zq0PgvtI0_2),.dout(w_dff_B_bh9e0hKE9_2),.clk(gclk));
	jdff dff_B_gvCo8ja90_2(.din(w_dff_B_bh9e0hKE9_2),.dout(w_dff_B_gvCo8ja90_2),.clk(gclk));
	jdff dff_B_vPabyj2N4_2(.din(w_dff_B_gvCo8ja90_2),.dout(w_dff_B_vPabyj2N4_2),.clk(gclk));
	jdff dff_B_C4KObj3N2_2(.din(w_dff_B_vPabyj2N4_2),.dout(w_dff_B_C4KObj3N2_2),.clk(gclk));
	jdff dff_B_6tM6Bikm2_2(.din(w_dff_B_C4KObj3N2_2),.dout(w_dff_B_6tM6Bikm2_2),.clk(gclk));
	jdff dff_B_Fxh8FrRE8_2(.din(w_dff_B_6tM6Bikm2_2),.dout(w_dff_B_Fxh8FrRE8_2),.clk(gclk));
	jdff dff_B_1eMWfmE62_2(.din(w_dff_B_Fxh8FrRE8_2),.dout(w_dff_B_1eMWfmE62_2),.clk(gclk));
	jdff dff_B_iLlOrbvU8_2(.din(w_dff_B_1eMWfmE62_2),.dout(w_dff_B_iLlOrbvU8_2),.clk(gclk));
	jdff dff_B_LoGDqp0X6_2(.din(w_dff_B_iLlOrbvU8_2),.dout(w_dff_B_LoGDqp0X6_2),.clk(gclk));
	jdff dff_B_24k2RjLd8_2(.din(w_dff_B_LoGDqp0X6_2),.dout(w_dff_B_24k2RjLd8_2),.clk(gclk));
	jdff dff_B_2fR7Wl904_2(.din(w_dff_B_24k2RjLd8_2),.dout(w_dff_B_2fR7Wl904_2),.clk(gclk));
	jdff dff_B_k1RGTAP00_2(.din(w_dff_B_2fR7Wl904_2),.dout(w_dff_B_k1RGTAP00_2),.clk(gclk));
	jdff dff_B_ccpovmWP2_2(.din(w_dff_B_k1RGTAP00_2),.dout(w_dff_B_ccpovmWP2_2),.clk(gclk));
	jdff dff_B_fyHA7Bdf4_2(.din(w_dff_B_ccpovmWP2_2),.dout(w_dff_B_fyHA7Bdf4_2),.clk(gclk));
	jdff dff_B_fu7MWsCY7_2(.din(w_dff_B_fyHA7Bdf4_2),.dout(w_dff_B_fu7MWsCY7_2),.clk(gclk));
	jdff dff_B_i43YjZIH4_2(.din(w_dff_B_fu7MWsCY7_2),.dout(w_dff_B_i43YjZIH4_2),.clk(gclk));
	jdff dff_B_Wv5N0oYO3_2(.din(w_dff_B_i43YjZIH4_2),.dout(w_dff_B_Wv5N0oYO3_2),.clk(gclk));
	jdff dff_B_cb5H1mkX6_2(.din(w_dff_B_Wv5N0oYO3_2),.dout(w_dff_B_cb5H1mkX6_2),.clk(gclk));
	jdff dff_B_QDSLTbY30_2(.din(w_dff_B_cb5H1mkX6_2),.dout(w_dff_B_QDSLTbY30_2),.clk(gclk));
	jdff dff_B_HCQgwVJi0_2(.din(n1360),.dout(w_dff_B_HCQgwVJi0_2),.clk(gclk));
	jdff dff_B_JqAWgDf77_1(.din(n1343),.dout(w_dff_B_JqAWgDf77_1),.clk(gclk));
	jdff dff_B_cjg5O9F09_2(.din(n1257),.dout(w_dff_B_cjg5O9F09_2),.clk(gclk));
	jdff dff_B_eD6PzqY11_2(.din(w_dff_B_cjg5O9F09_2),.dout(w_dff_B_eD6PzqY11_2),.clk(gclk));
	jdff dff_B_0mU4iFnm1_2(.din(w_dff_B_eD6PzqY11_2),.dout(w_dff_B_0mU4iFnm1_2),.clk(gclk));
	jdff dff_B_sXGLcywk4_2(.din(w_dff_B_0mU4iFnm1_2),.dout(w_dff_B_sXGLcywk4_2),.clk(gclk));
	jdff dff_B_83KL4U2s0_2(.din(w_dff_B_sXGLcywk4_2),.dout(w_dff_B_83KL4U2s0_2),.clk(gclk));
	jdff dff_B_qnPe1rC34_2(.din(w_dff_B_83KL4U2s0_2),.dout(w_dff_B_qnPe1rC34_2),.clk(gclk));
	jdff dff_B_FjH128Yc7_2(.din(w_dff_B_qnPe1rC34_2),.dout(w_dff_B_FjH128Yc7_2),.clk(gclk));
	jdff dff_B_3MVQSV9i7_2(.din(w_dff_B_FjH128Yc7_2),.dout(w_dff_B_3MVQSV9i7_2),.clk(gclk));
	jdff dff_B_7RFmhv6M5_2(.din(w_dff_B_3MVQSV9i7_2),.dout(w_dff_B_7RFmhv6M5_2),.clk(gclk));
	jdff dff_B_9bqj45Az9_2(.din(w_dff_B_7RFmhv6M5_2),.dout(w_dff_B_9bqj45Az9_2),.clk(gclk));
	jdff dff_B_jcI5yAf75_2(.din(w_dff_B_9bqj45Az9_2),.dout(w_dff_B_jcI5yAf75_2),.clk(gclk));
	jdff dff_B_e3mmbSYq6_2(.din(w_dff_B_jcI5yAf75_2),.dout(w_dff_B_e3mmbSYq6_2),.clk(gclk));
	jdff dff_B_jtjhHmXu3_2(.din(w_dff_B_e3mmbSYq6_2),.dout(w_dff_B_jtjhHmXu3_2),.clk(gclk));
	jdff dff_B_BQSGshNK2_2(.din(w_dff_B_jtjhHmXu3_2),.dout(w_dff_B_BQSGshNK2_2),.clk(gclk));
	jdff dff_B_hiE1BAur6_2(.din(w_dff_B_BQSGshNK2_2),.dout(w_dff_B_hiE1BAur6_2),.clk(gclk));
	jdff dff_B_PBJpxvx89_2(.din(w_dff_B_hiE1BAur6_2),.dout(w_dff_B_PBJpxvx89_2),.clk(gclk));
	jdff dff_B_2sugV3bU7_2(.din(w_dff_B_PBJpxvx89_2),.dout(w_dff_B_2sugV3bU7_2),.clk(gclk));
	jdff dff_B_xIxdlzct2_2(.din(w_dff_B_2sugV3bU7_2),.dout(w_dff_B_xIxdlzct2_2),.clk(gclk));
	jdff dff_B_swwuuHOT8_2(.din(w_dff_B_xIxdlzct2_2),.dout(w_dff_B_swwuuHOT8_2),.clk(gclk));
	jdff dff_B_f1fCDRhk4_2(.din(w_dff_B_swwuuHOT8_2),.dout(w_dff_B_f1fCDRhk4_2),.clk(gclk));
	jdff dff_B_Xe6He2ej0_2(.din(n1275),.dout(w_dff_B_Xe6He2ej0_2),.clk(gclk));
	jdff dff_B_bVIrtuqp5_1(.din(n1258),.dout(w_dff_B_bVIrtuqp5_1),.clk(gclk));
	jdff dff_B_6m1xM35V8_2(.din(n1166),.dout(w_dff_B_6m1xM35V8_2),.clk(gclk));
	jdff dff_B_Cg7d4s2f6_2(.din(w_dff_B_6m1xM35V8_2),.dout(w_dff_B_Cg7d4s2f6_2),.clk(gclk));
	jdff dff_B_WXTTm8Gk6_2(.din(w_dff_B_Cg7d4s2f6_2),.dout(w_dff_B_WXTTm8Gk6_2),.clk(gclk));
	jdff dff_B_QmjzsAcW2_2(.din(w_dff_B_WXTTm8Gk6_2),.dout(w_dff_B_QmjzsAcW2_2),.clk(gclk));
	jdff dff_B_LtJR30tu6_2(.din(w_dff_B_QmjzsAcW2_2),.dout(w_dff_B_LtJR30tu6_2),.clk(gclk));
	jdff dff_B_Nsc63dWk3_2(.din(w_dff_B_LtJR30tu6_2),.dout(w_dff_B_Nsc63dWk3_2),.clk(gclk));
	jdff dff_B_DompU1Mn5_2(.din(w_dff_B_Nsc63dWk3_2),.dout(w_dff_B_DompU1Mn5_2),.clk(gclk));
	jdff dff_B_qNgr9wnv7_2(.din(w_dff_B_DompU1Mn5_2),.dout(w_dff_B_qNgr9wnv7_2),.clk(gclk));
	jdff dff_B_7qLpwFRF7_2(.din(w_dff_B_qNgr9wnv7_2),.dout(w_dff_B_7qLpwFRF7_2),.clk(gclk));
	jdff dff_B_FMwohWg13_2(.din(w_dff_B_7qLpwFRF7_2),.dout(w_dff_B_FMwohWg13_2),.clk(gclk));
	jdff dff_B_sm3ZAiPd7_2(.din(w_dff_B_FMwohWg13_2),.dout(w_dff_B_sm3ZAiPd7_2),.clk(gclk));
	jdff dff_B_PGvRhzpx8_2(.din(w_dff_B_sm3ZAiPd7_2),.dout(w_dff_B_PGvRhzpx8_2),.clk(gclk));
	jdff dff_B_Ff6loTOH1_2(.din(w_dff_B_PGvRhzpx8_2),.dout(w_dff_B_Ff6loTOH1_2),.clk(gclk));
	jdff dff_B_JGntCBvc0_2(.din(w_dff_B_Ff6loTOH1_2),.dout(w_dff_B_JGntCBvc0_2),.clk(gclk));
	jdff dff_B_tgJVvPhR1_2(.din(w_dff_B_JGntCBvc0_2),.dout(w_dff_B_tgJVvPhR1_2),.clk(gclk));
	jdff dff_B_fYzdwXKl8_2(.din(w_dff_B_tgJVvPhR1_2),.dout(w_dff_B_fYzdwXKl8_2),.clk(gclk));
	jdff dff_B_n2dKzKE83_2(.din(w_dff_B_fYzdwXKl8_2),.dout(w_dff_B_n2dKzKE83_2),.clk(gclk));
	jdff dff_B_I90VvDvk6_2(.din(n1184),.dout(w_dff_B_I90VvDvk6_2),.clk(gclk));
	jdff dff_B_RyEVqxOx9_1(.din(n1167),.dout(w_dff_B_RyEVqxOx9_1),.clk(gclk));
	jdff dff_B_5y5m7if40_2(.din(n1068),.dout(w_dff_B_5y5m7if40_2),.clk(gclk));
	jdff dff_B_C7NOqQmo0_2(.din(w_dff_B_5y5m7if40_2),.dout(w_dff_B_C7NOqQmo0_2),.clk(gclk));
	jdff dff_B_nOiyILY67_2(.din(w_dff_B_C7NOqQmo0_2),.dout(w_dff_B_nOiyILY67_2),.clk(gclk));
	jdff dff_B_Nr3nNIHK5_2(.din(w_dff_B_nOiyILY67_2),.dout(w_dff_B_Nr3nNIHK5_2),.clk(gclk));
	jdff dff_B_Sldwm07Z4_2(.din(w_dff_B_Nr3nNIHK5_2),.dout(w_dff_B_Sldwm07Z4_2),.clk(gclk));
	jdff dff_B_696ONaBT7_2(.din(w_dff_B_Sldwm07Z4_2),.dout(w_dff_B_696ONaBT7_2),.clk(gclk));
	jdff dff_B_5WJOaiIf6_2(.din(w_dff_B_696ONaBT7_2),.dout(w_dff_B_5WJOaiIf6_2),.clk(gclk));
	jdff dff_B_owGEMTNz7_2(.din(w_dff_B_5WJOaiIf6_2),.dout(w_dff_B_owGEMTNz7_2),.clk(gclk));
	jdff dff_B_MTvfbLHM2_2(.din(w_dff_B_owGEMTNz7_2),.dout(w_dff_B_MTvfbLHM2_2),.clk(gclk));
	jdff dff_B_QejiHL5P1_2(.din(w_dff_B_MTvfbLHM2_2),.dout(w_dff_B_QejiHL5P1_2),.clk(gclk));
	jdff dff_B_blyeLdE39_2(.din(w_dff_B_QejiHL5P1_2),.dout(w_dff_B_blyeLdE39_2),.clk(gclk));
	jdff dff_B_ftThUZDC8_2(.din(w_dff_B_blyeLdE39_2),.dout(w_dff_B_ftThUZDC8_2),.clk(gclk));
	jdff dff_B_1OYb2m226_2(.din(w_dff_B_ftThUZDC8_2),.dout(w_dff_B_1OYb2m226_2),.clk(gclk));
	jdff dff_B_Ci9wtgQJ5_2(.din(w_dff_B_1OYb2m226_2),.dout(w_dff_B_Ci9wtgQJ5_2),.clk(gclk));
	jdff dff_B_smVEtmv42_2(.din(n1085),.dout(w_dff_B_smVEtmv42_2),.clk(gclk));
	jdff dff_B_zrwX1Wfj8_1(.din(n1069),.dout(w_dff_B_zrwX1Wfj8_1),.clk(gclk));
	jdff dff_B_Vyrvde2k7_2(.din(n969),.dout(w_dff_B_Vyrvde2k7_2),.clk(gclk));
	jdff dff_B_7dHNVaiX3_2(.din(w_dff_B_Vyrvde2k7_2),.dout(w_dff_B_7dHNVaiX3_2),.clk(gclk));
	jdff dff_B_Z07SO9pK4_2(.din(w_dff_B_7dHNVaiX3_2),.dout(w_dff_B_Z07SO9pK4_2),.clk(gclk));
	jdff dff_B_CU3VdFFs7_2(.din(w_dff_B_Z07SO9pK4_2),.dout(w_dff_B_CU3VdFFs7_2),.clk(gclk));
	jdff dff_B_1pRFknuG1_2(.din(w_dff_B_CU3VdFFs7_2),.dout(w_dff_B_1pRFknuG1_2),.clk(gclk));
	jdff dff_B_pDyPHFbo8_2(.din(w_dff_B_1pRFknuG1_2),.dout(w_dff_B_pDyPHFbo8_2),.clk(gclk));
	jdff dff_B_hW581FkD7_2(.din(w_dff_B_pDyPHFbo8_2),.dout(w_dff_B_hW581FkD7_2),.clk(gclk));
	jdff dff_B_ax2HaJUt4_2(.din(w_dff_B_hW581FkD7_2),.dout(w_dff_B_ax2HaJUt4_2),.clk(gclk));
	jdff dff_B_XyB4ET0e1_2(.din(w_dff_B_ax2HaJUt4_2),.dout(w_dff_B_XyB4ET0e1_2),.clk(gclk));
	jdff dff_B_7FkRkUes7_2(.din(w_dff_B_XyB4ET0e1_2),.dout(w_dff_B_7FkRkUes7_2),.clk(gclk));
	jdff dff_B_imKGIIwC7_2(.din(w_dff_B_7FkRkUes7_2),.dout(w_dff_B_imKGIIwC7_2),.clk(gclk));
	jdff dff_B_NGWTcjpH5_2(.din(n986),.dout(w_dff_B_NGWTcjpH5_2),.clk(gclk));
	jdff dff_B_4oC1homs9_1(.din(n970),.dout(w_dff_B_4oC1homs9_1),.clk(gclk));
	jdff dff_B_aWKR5lhH0_2(.din(n867),.dout(w_dff_B_aWKR5lhH0_2),.clk(gclk));
	jdff dff_B_AciXEQ3X1_2(.din(w_dff_B_aWKR5lhH0_2),.dout(w_dff_B_AciXEQ3X1_2),.clk(gclk));
	jdff dff_B_RC2f9G3l3_2(.din(w_dff_B_AciXEQ3X1_2),.dout(w_dff_B_RC2f9G3l3_2),.clk(gclk));
	jdff dff_B_EuFkQLMU9_2(.din(w_dff_B_RC2f9G3l3_2),.dout(w_dff_B_EuFkQLMU9_2),.clk(gclk));
	jdff dff_B_d7qrxhmy8_2(.din(w_dff_B_EuFkQLMU9_2),.dout(w_dff_B_d7qrxhmy8_2),.clk(gclk));
	jdff dff_B_lKZInh7R6_2(.din(w_dff_B_d7qrxhmy8_2),.dout(w_dff_B_lKZInh7R6_2),.clk(gclk));
	jdff dff_B_lvn5e4YR2_2(.din(w_dff_B_lKZInh7R6_2),.dout(w_dff_B_lvn5e4YR2_2),.clk(gclk));
	jdff dff_B_wSpih1Qt8_2(.din(w_dff_B_lvn5e4YR2_2),.dout(w_dff_B_wSpih1Qt8_2),.clk(gclk));
	jdff dff_B_9x4o2KCf7_2(.din(n880),.dout(w_dff_B_9x4o2KCf7_2),.clk(gclk));
	jdff dff_B_OzCmzcbf7_2(.din(w_dff_B_9x4o2KCf7_2),.dout(w_dff_B_OzCmzcbf7_2),.clk(gclk));
	jdff dff_B_aL4m3DRC6_2(.din(w_dff_B_OzCmzcbf7_2),.dout(w_dff_B_aL4m3DRC6_2),.clk(gclk));
	jdff dff_B_9hdXcse39_1(.din(n868),.dout(w_dff_B_9hdXcse39_1),.clk(gclk));
	jdff dff_B_IPyqcC861_1(.din(w_dff_B_9hdXcse39_1),.dout(w_dff_B_IPyqcC861_1),.clk(gclk));
	jdff dff_B_U4bDjFzh5_2(.din(n771),.dout(w_dff_B_U4bDjFzh5_2),.clk(gclk));
	jdff dff_B_LYiWz5wH8_2(.din(w_dff_B_U4bDjFzh5_2),.dout(w_dff_B_LYiWz5wH8_2),.clk(gclk));
	jdff dff_B_BUBibZu93_2(.din(w_dff_B_LYiWz5wH8_2),.dout(w_dff_B_BUBibZu93_2),.clk(gclk));
	jdff dff_B_A0THsbh72_0(.din(n776),.dout(w_dff_B_A0THsbh72_0),.clk(gclk));
	jdff dff_A_sRUxz9k22_0(.dout(w_n676_0[0]),.din(w_dff_A_sRUxz9k22_0),.clk(gclk));
	jdff dff_A_sb8ifWuf6_0(.dout(w_dff_A_sRUxz9k22_0),.din(w_dff_A_sb8ifWuf6_0),.clk(gclk));
	jdff dff_A_v5IQem1f2_1(.dout(w_n676_0[1]),.din(w_dff_A_v5IQem1f2_1),.clk(gclk));
	jdff dff_A_YptSCDAG8_1(.dout(w_dff_A_v5IQem1f2_1),.din(w_dff_A_YptSCDAG8_1),.clk(gclk));
	jdff dff_B_3khtPMZW2_1(.din(n1812),.dout(w_dff_B_3khtPMZW2_1),.clk(gclk));
	jdff dff_B_9DLV4WV10_1(.din(n1799),.dout(w_dff_B_9DLV4WV10_1),.clk(gclk));
	jdff dff_B_faZ3ZuPl5_1(.din(w_dff_B_9DLV4WV10_1),.dout(w_dff_B_faZ3ZuPl5_1),.clk(gclk));
	jdff dff_B_MfPpxzJJ9_2(.din(n1798),.dout(w_dff_B_MfPpxzJJ9_2),.clk(gclk));
	jdff dff_B_wqld1sS99_2(.din(w_dff_B_MfPpxzJJ9_2),.dout(w_dff_B_wqld1sS99_2),.clk(gclk));
	jdff dff_B_TFMUueFe3_2(.din(w_dff_B_wqld1sS99_2),.dout(w_dff_B_TFMUueFe3_2),.clk(gclk));
	jdff dff_B_meT1L5XU9_2(.din(w_dff_B_TFMUueFe3_2),.dout(w_dff_B_meT1L5XU9_2),.clk(gclk));
	jdff dff_B_eIGPAlFf5_2(.din(w_dff_B_meT1L5XU9_2),.dout(w_dff_B_eIGPAlFf5_2),.clk(gclk));
	jdff dff_B_GYFatfmk0_2(.din(w_dff_B_eIGPAlFf5_2),.dout(w_dff_B_GYFatfmk0_2),.clk(gclk));
	jdff dff_B_UFZSArsj2_2(.din(w_dff_B_GYFatfmk0_2),.dout(w_dff_B_UFZSArsj2_2),.clk(gclk));
	jdff dff_B_brlA7cSV0_2(.din(w_dff_B_UFZSArsj2_2),.dout(w_dff_B_brlA7cSV0_2),.clk(gclk));
	jdff dff_B_m91rymN61_2(.din(w_dff_B_brlA7cSV0_2),.dout(w_dff_B_m91rymN61_2),.clk(gclk));
	jdff dff_B_bZPLzYsL4_2(.din(w_dff_B_m91rymN61_2),.dout(w_dff_B_bZPLzYsL4_2),.clk(gclk));
	jdff dff_B_g3fF2vhK7_2(.din(w_dff_B_bZPLzYsL4_2),.dout(w_dff_B_g3fF2vhK7_2),.clk(gclk));
	jdff dff_B_NSDCk7Dd7_2(.din(w_dff_B_g3fF2vhK7_2),.dout(w_dff_B_NSDCk7Dd7_2),.clk(gclk));
	jdff dff_B_GX258PLG1_2(.din(w_dff_B_NSDCk7Dd7_2),.dout(w_dff_B_GX258PLG1_2),.clk(gclk));
	jdff dff_B_GlgEY3dY5_2(.din(w_dff_B_GX258PLG1_2),.dout(w_dff_B_GlgEY3dY5_2),.clk(gclk));
	jdff dff_B_w9khd0Be5_2(.din(w_dff_B_GlgEY3dY5_2),.dout(w_dff_B_w9khd0Be5_2),.clk(gclk));
	jdff dff_B_2lfrzC9f1_2(.din(w_dff_B_w9khd0Be5_2),.dout(w_dff_B_2lfrzC9f1_2),.clk(gclk));
	jdff dff_B_9PLjGxQl9_2(.din(w_dff_B_2lfrzC9f1_2),.dout(w_dff_B_9PLjGxQl9_2),.clk(gclk));
	jdff dff_B_LiCwUIuV8_2(.din(w_dff_B_9PLjGxQl9_2),.dout(w_dff_B_LiCwUIuV8_2),.clk(gclk));
	jdff dff_B_hYnWIWjr6_2(.din(w_dff_B_LiCwUIuV8_2),.dout(w_dff_B_hYnWIWjr6_2),.clk(gclk));
	jdff dff_B_Xmzl4cMp4_2(.din(w_dff_B_hYnWIWjr6_2),.dout(w_dff_B_Xmzl4cMp4_2),.clk(gclk));
	jdff dff_B_NoZ2XuEd6_2(.din(w_dff_B_Xmzl4cMp4_2),.dout(w_dff_B_NoZ2XuEd6_2),.clk(gclk));
	jdff dff_B_uHW3695z4_2(.din(w_dff_B_NoZ2XuEd6_2),.dout(w_dff_B_uHW3695z4_2),.clk(gclk));
	jdff dff_B_YYFN2Zed4_2(.din(w_dff_B_uHW3695z4_2),.dout(w_dff_B_YYFN2Zed4_2),.clk(gclk));
	jdff dff_B_yYEalvjV5_2(.din(w_dff_B_YYFN2Zed4_2),.dout(w_dff_B_yYEalvjV5_2),.clk(gclk));
	jdff dff_B_NvM6fDmN8_2(.din(w_dff_B_yYEalvjV5_2),.dout(w_dff_B_NvM6fDmN8_2),.clk(gclk));
	jdff dff_B_BuhkKyiz1_2(.din(w_dff_B_NvM6fDmN8_2),.dout(w_dff_B_BuhkKyiz1_2),.clk(gclk));
	jdff dff_B_USWE1dzW0_2(.din(w_dff_B_BuhkKyiz1_2),.dout(w_dff_B_USWE1dzW0_2),.clk(gclk));
	jdff dff_B_HpAjlrzA1_2(.din(w_dff_B_USWE1dzW0_2),.dout(w_dff_B_HpAjlrzA1_2),.clk(gclk));
	jdff dff_B_vYBqpBVu4_2(.din(w_dff_B_HpAjlrzA1_2),.dout(w_dff_B_vYBqpBVu4_2),.clk(gclk));
	jdff dff_B_UJbJAONb9_2(.din(w_dff_B_vYBqpBVu4_2),.dout(w_dff_B_UJbJAONb9_2),.clk(gclk));
	jdff dff_B_PHo3CXyP2_2(.din(w_dff_B_UJbJAONb9_2),.dout(w_dff_B_PHo3CXyP2_2),.clk(gclk));
	jdff dff_B_mcM7JGJ51_2(.din(w_dff_B_PHo3CXyP2_2),.dout(w_dff_B_mcM7JGJ51_2),.clk(gclk));
	jdff dff_B_fdrUX4wB3_2(.din(w_dff_B_mcM7JGJ51_2),.dout(w_dff_B_fdrUX4wB3_2),.clk(gclk));
	jdff dff_B_s1gwsI996_2(.din(w_dff_B_fdrUX4wB3_2),.dout(w_dff_B_s1gwsI996_2),.clk(gclk));
	jdff dff_B_FQBwSGez0_2(.din(w_dff_B_s1gwsI996_2),.dout(w_dff_B_FQBwSGez0_2),.clk(gclk));
	jdff dff_B_sHeUz6nC6_2(.din(w_dff_B_FQBwSGez0_2),.dout(w_dff_B_sHeUz6nC6_2),.clk(gclk));
	jdff dff_B_cOsl4YVb1_2(.din(w_dff_B_sHeUz6nC6_2),.dout(w_dff_B_cOsl4YVb1_2),.clk(gclk));
	jdff dff_B_fTwFTflT5_2(.din(w_dff_B_cOsl4YVb1_2),.dout(w_dff_B_fTwFTflT5_2),.clk(gclk));
	jdff dff_B_H5yL1yby8_2(.din(w_dff_B_fTwFTflT5_2),.dout(w_dff_B_H5yL1yby8_2),.clk(gclk));
	jdff dff_B_a8SEDwBz6_2(.din(w_dff_B_H5yL1yby8_2),.dout(w_dff_B_a8SEDwBz6_2),.clk(gclk));
	jdff dff_B_TwxTjr6m7_2(.din(w_dff_B_a8SEDwBz6_2),.dout(w_dff_B_TwxTjr6m7_2),.clk(gclk));
	jdff dff_B_Yxnipmd05_2(.din(w_dff_B_TwxTjr6m7_2),.dout(w_dff_B_Yxnipmd05_2),.clk(gclk));
	jdff dff_B_0gvTZBI68_2(.din(w_dff_B_Yxnipmd05_2),.dout(w_dff_B_0gvTZBI68_2),.clk(gclk));
	jdff dff_B_PB7KWXqT8_2(.din(w_dff_B_0gvTZBI68_2),.dout(w_dff_B_PB7KWXqT8_2),.clk(gclk));
	jdff dff_B_Lko5MVvg3_2(.din(w_dff_B_PB7KWXqT8_2),.dout(w_dff_B_Lko5MVvg3_2),.clk(gclk));
	jdff dff_B_HSCpKC7y0_2(.din(w_dff_B_Lko5MVvg3_2),.dout(w_dff_B_HSCpKC7y0_2),.clk(gclk));
	jdff dff_B_OrMGwLI38_2(.din(w_dff_B_HSCpKC7y0_2),.dout(w_dff_B_OrMGwLI38_2),.clk(gclk));
	jdff dff_B_uTO94k8z0_2(.din(w_dff_B_OrMGwLI38_2),.dout(w_dff_B_uTO94k8z0_2),.clk(gclk));
	jdff dff_B_Jj1COXCJ9_2(.din(w_dff_B_uTO94k8z0_2),.dout(w_dff_B_Jj1COXCJ9_2),.clk(gclk));
	jdff dff_B_Ar2B9dB93_2(.din(w_dff_B_Jj1COXCJ9_2),.dout(w_dff_B_Ar2B9dB93_2),.clk(gclk));
	jdff dff_B_fkpKJ1nu2_2(.din(w_dff_B_Ar2B9dB93_2),.dout(w_dff_B_fkpKJ1nu2_2),.clk(gclk));
	jdff dff_B_77zVpOrb5_2(.din(w_dff_B_fkpKJ1nu2_2),.dout(w_dff_B_77zVpOrb5_2),.clk(gclk));
	jdff dff_B_6aixUHpW2_2(.din(w_dff_B_77zVpOrb5_2),.dout(w_dff_B_6aixUHpW2_2),.clk(gclk));
	jdff dff_B_IGeMV9ib9_2(.din(n1797),.dout(w_dff_B_IGeMV9ib9_2),.clk(gclk));
	jdff dff_B_1hXPoMWS8_2(.din(w_dff_B_IGeMV9ib9_2),.dout(w_dff_B_1hXPoMWS8_2),.clk(gclk));
	jdff dff_B_hTm9IOLP4_2(.din(w_dff_B_1hXPoMWS8_2),.dout(w_dff_B_hTm9IOLP4_2),.clk(gclk));
	jdff dff_B_lUSdTHp65_2(.din(w_dff_B_hTm9IOLP4_2),.dout(w_dff_B_lUSdTHp65_2),.clk(gclk));
	jdff dff_B_nkhFoypa0_2(.din(w_dff_B_lUSdTHp65_2),.dout(w_dff_B_nkhFoypa0_2),.clk(gclk));
	jdff dff_B_hFKUTLDw7_2(.din(w_dff_B_nkhFoypa0_2),.dout(w_dff_B_hFKUTLDw7_2),.clk(gclk));
	jdff dff_B_OlSnPDNG8_2(.din(w_dff_B_hFKUTLDw7_2),.dout(w_dff_B_OlSnPDNG8_2),.clk(gclk));
	jdff dff_B_MJVdG18b0_2(.din(w_dff_B_OlSnPDNG8_2),.dout(w_dff_B_MJVdG18b0_2),.clk(gclk));
	jdff dff_B_uHrKPwcu2_2(.din(w_dff_B_MJVdG18b0_2),.dout(w_dff_B_uHrKPwcu2_2),.clk(gclk));
	jdff dff_B_ARfFCk4c8_2(.din(w_dff_B_uHrKPwcu2_2),.dout(w_dff_B_ARfFCk4c8_2),.clk(gclk));
	jdff dff_B_0uOtnRUs4_2(.din(w_dff_B_ARfFCk4c8_2),.dout(w_dff_B_0uOtnRUs4_2),.clk(gclk));
	jdff dff_B_GgziSO107_2(.din(w_dff_B_0uOtnRUs4_2),.dout(w_dff_B_GgziSO107_2),.clk(gclk));
	jdff dff_B_f2H1AQPX8_2(.din(w_dff_B_GgziSO107_2),.dout(w_dff_B_f2H1AQPX8_2),.clk(gclk));
	jdff dff_B_Wbda1GtI8_2(.din(w_dff_B_f2H1AQPX8_2),.dout(w_dff_B_Wbda1GtI8_2),.clk(gclk));
	jdff dff_B_YzgAQTqb6_2(.din(w_dff_B_Wbda1GtI8_2),.dout(w_dff_B_YzgAQTqb6_2),.clk(gclk));
	jdff dff_B_5a1WIX7l3_2(.din(w_dff_B_YzgAQTqb6_2),.dout(w_dff_B_5a1WIX7l3_2),.clk(gclk));
	jdff dff_B_DGGBXSaQ6_2(.din(w_dff_B_5a1WIX7l3_2),.dout(w_dff_B_DGGBXSaQ6_2),.clk(gclk));
	jdff dff_B_zKSRgERY3_2(.din(w_dff_B_DGGBXSaQ6_2),.dout(w_dff_B_zKSRgERY3_2),.clk(gclk));
	jdff dff_B_ZH41LcwF6_2(.din(w_dff_B_zKSRgERY3_2),.dout(w_dff_B_ZH41LcwF6_2),.clk(gclk));
	jdff dff_B_JxGqPK4N2_2(.din(w_dff_B_ZH41LcwF6_2),.dout(w_dff_B_JxGqPK4N2_2),.clk(gclk));
	jdff dff_B_vdOInZ5o7_2(.din(w_dff_B_JxGqPK4N2_2),.dout(w_dff_B_vdOInZ5o7_2),.clk(gclk));
	jdff dff_B_wq5U4Wf54_2(.din(w_dff_B_vdOInZ5o7_2),.dout(w_dff_B_wq5U4Wf54_2),.clk(gclk));
	jdff dff_B_8DNgGRHO6_2(.din(w_dff_B_wq5U4Wf54_2),.dout(w_dff_B_8DNgGRHO6_2),.clk(gclk));
	jdff dff_B_hBdRicXW5_2(.din(w_dff_B_8DNgGRHO6_2),.dout(w_dff_B_hBdRicXW5_2),.clk(gclk));
	jdff dff_B_y05gS8lc0_2(.din(w_dff_B_hBdRicXW5_2),.dout(w_dff_B_y05gS8lc0_2),.clk(gclk));
	jdff dff_B_CKs8n0Ga0_2(.din(w_dff_B_y05gS8lc0_2),.dout(w_dff_B_CKs8n0Ga0_2),.clk(gclk));
	jdff dff_B_QSqeWaxf5_2(.din(w_dff_B_CKs8n0Ga0_2),.dout(w_dff_B_QSqeWaxf5_2),.clk(gclk));
	jdff dff_B_vkXyBreC2_2(.din(w_dff_B_QSqeWaxf5_2),.dout(w_dff_B_vkXyBreC2_2),.clk(gclk));
	jdff dff_B_RH3bIGlB7_2(.din(w_dff_B_vkXyBreC2_2),.dout(w_dff_B_RH3bIGlB7_2),.clk(gclk));
	jdff dff_B_nkG0x9KF5_2(.din(w_dff_B_RH3bIGlB7_2),.dout(w_dff_B_nkG0x9KF5_2),.clk(gclk));
	jdff dff_B_99JDZfRv1_2(.din(w_dff_B_nkG0x9KF5_2),.dout(w_dff_B_99JDZfRv1_2),.clk(gclk));
	jdff dff_B_gC5WPp5f2_2(.din(w_dff_B_99JDZfRv1_2),.dout(w_dff_B_gC5WPp5f2_2),.clk(gclk));
	jdff dff_B_9gwnppzM2_2(.din(w_dff_B_gC5WPp5f2_2),.dout(w_dff_B_9gwnppzM2_2),.clk(gclk));
	jdff dff_B_UGPfeOys5_2(.din(w_dff_B_9gwnppzM2_2),.dout(w_dff_B_UGPfeOys5_2),.clk(gclk));
	jdff dff_B_1p3qAfnr3_2(.din(w_dff_B_UGPfeOys5_2),.dout(w_dff_B_1p3qAfnr3_2),.clk(gclk));
	jdff dff_B_nzqDpM5g9_2(.din(w_dff_B_1p3qAfnr3_2),.dout(w_dff_B_nzqDpM5g9_2),.clk(gclk));
	jdff dff_B_j2gRuAmv6_2(.din(w_dff_B_nzqDpM5g9_2),.dout(w_dff_B_j2gRuAmv6_2),.clk(gclk));
	jdff dff_B_qjyyVmx96_2(.din(w_dff_B_j2gRuAmv6_2),.dout(w_dff_B_qjyyVmx96_2),.clk(gclk));
	jdff dff_B_MOd2wavx1_2(.din(w_dff_B_qjyyVmx96_2),.dout(w_dff_B_MOd2wavx1_2),.clk(gclk));
	jdff dff_B_edEKACBM9_2(.din(w_dff_B_MOd2wavx1_2),.dout(w_dff_B_edEKACBM9_2),.clk(gclk));
	jdff dff_B_iMCb9WWC1_2(.din(w_dff_B_edEKACBM9_2),.dout(w_dff_B_iMCb9WWC1_2),.clk(gclk));
	jdff dff_B_2EolgRcV6_2(.din(w_dff_B_iMCb9WWC1_2),.dout(w_dff_B_2EolgRcV6_2),.clk(gclk));
	jdff dff_B_eQikfSyF9_2(.din(w_dff_B_2EolgRcV6_2),.dout(w_dff_B_eQikfSyF9_2),.clk(gclk));
	jdff dff_B_zZP6iBpU1_2(.din(w_dff_B_eQikfSyF9_2),.dout(w_dff_B_zZP6iBpU1_2),.clk(gclk));
	jdff dff_B_sxPkbQoA5_2(.din(w_dff_B_zZP6iBpU1_2),.dout(w_dff_B_sxPkbQoA5_2),.clk(gclk));
	jdff dff_B_UVizJ9OA6_2(.din(w_dff_B_sxPkbQoA5_2),.dout(w_dff_B_UVizJ9OA6_2),.clk(gclk));
	jdff dff_B_Qmo4U34Y5_2(.din(w_dff_B_UVizJ9OA6_2),.dout(w_dff_B_Qmo4U34Y5_2),.clk(gclk));
	jdff dff_B_PxKGak9c1_2(.din(w_dff_B_Qmo4U34Y5_2),.dout(w_dff_B_PxKGak9c1_2),.clk(gclk));
	jdff dff_B_bZvZbHM05_2(.din(w_dff_B_PxKGak9c1_2),.dout(w_dff_B_bZvZbHM05_2),.clk(gclk));
	jdff dff_B_BTIdkmGU8_2(.din(w_dff_B_bZvZbHM05_2),.dout(w_dff_B_BTIdkmGU8_2),.clk(gclk));
	jdff dff_B_LjShF65B1_2(.din(w_dff_B_BTIdkmGU8_2),.dout(w_dff_B_LjShF65B1_2),.clk(gclk));
	jdff dff_B_Sx5j2Lhm8_2(.din(w_dff_B_LjShF65B1_2),.dout(w_dff_B_Sx5j2Lhm8_2),.clk(gclk));
	jdff dff_B_wGYfX4iD3_2(.din(w_dff_B_Sx5j2Lhm8_2),.dout(w_dff_B_wGYfX4iD3_2),.clk(gclk));
	jdff dff_B_77mgntCa2_2(.din(w_dff_B_wGYfX4iD3_2),.dout(w_dff_B_77mgntCa2_2),.clk(gclk));
	jdff dff_B_JTBAVYp00_2(.din(w_dff_B_77mgntCa2_2),.dout(w_dff_B_JTBAVYp00_2),.clk(gclk));
	jdff dff_A_kIMEJZuV4_1(.dout(w_n1796_0[1]),.din(w_dff_A_kIMEJZuV4_1),.clk(gclk));
	jdff dff_B_kLCCYxg90_1(.din(n1794),.dout(w_dff_B_kLCCYxg90_1),.clk(gclk));
	jdff dff_B_6WvChU4n7_2(.din(n1772),.dout(w_dff_B_6WvChU4n7_2),.clk(gclk));
	jdff dff_B_VeE8k1Js9_2(.din(w_dff_B_6WvChU4n7_2),.dout(w_dff_B_VeE8k1Js9_2),.clk(gclk));
	jdff dff_B_b0ffJJZ37_2(.din(w_dff_B_VeE8k1Js9_2),.dout(w_dff_B_b0ffJJZ37_2),.clk(gclk));
	jdff dff_B_qUAGjAFZ7_2(.din(w_dff_B_b0ffJJZ37_2),.dout(w_dff_B_qUAGjAFZ7_2),.clk(gclk));
	jdff dff_B_HbUZ7giP6_2(.din(w_dff_B_qUAGjAFZ7_2),.dout(w_dff_B_HbUZ7giP6_2),.clk(gclk));
	jdff dff_B_225T9Tfg2_2(.din(w_dff_B_HbUZ7giP6_2),.dout(w_dff_B_225T9Tfg2_2),.clk(gclk));
	jdff dff_B_2Ebq5G2f8_2(.din(w_dff_B_225T9Tfg2_2),.dout(w_dff_B_2Ebq5G2f8_2),.clk(gclk));
	jdff dff_B_qLonYJt09_2(.din(w_dff_B_2Ebq5G2f8_2),.dout(w_dff_B_qLonYJt09_2),.clk(gclk));
	jdff dff_B_rW4he9le3_2(.din(w_dff_B_qLonYJt09_2),.dout(w_dff_B_rW4he9le3_2),.clk(gclk));
	jdff dff_B_WltqSuis1_2(.din(w_dff_B_rW4he9le3_2),.dout(w_dff_B_WltqSuis1_2),.clk(gclk));
	jdff dff_B_WH1ZPVG68_2(.din(w_dff_B_WltqSuis1_2),.dout(w_dff_B_WH1ZPVG68_2),.clk(gclk));
	jdff dff_B_JxdmMQdi8_2(.din(w_dff_B_WH1ZPVG68_2),.dout(w_dff_B_JxdmMQdi8_2),.clk(gclk));
	jdff dff_B_YtQ5t4BL2_2(.din(w_dff_B_JxdmMQdi8_2),.dout(w_dff_B_YtQ5t4BL2_2),.clk(gclk));
	jdff dff_B_9cMtjPah8_2(.din(w_dff_B_YtQ5t4BL2_2),.dout(w_dff_B_9cMtjPah8_2),.clk(gclk));
	jdff dff_B_T714fXWc2_2(.din(w_dff_B_9cMtjPah8_2),.dout(w_dff_B_T714fXWc2_2),.clk(gclk));
	jdff dff_B_5ehTGXKN0_2(.din(w_dff_B_T714fXWc2_2),.dout(w_dff_B_5ehTGXKN0_2),.clk(gclk));
	jdff dff_B_U3HENvgj9_2(.din(w_dff_B_5ehTGXKN0_2),.dout(w_dff_B_U3HENvgj9_2),.clk(gclk));
	jdff dff_B_sale1tLe9_2(.din(w_dff_B_U3HENvgj9_2),.dout(w_dff_B_sale1tLe9_2),.clk(gclk));
	jdff dff_B_uG6YmGoK2_2(.din(w_dff_B_sale1tLe9_2),.dout(w_dff_B_uG6YmGoK2_2),.clk(gclk));
	jdff dff_B_ucI4AD7R8_2(.din(w_dff_B_uG6YmGoK2_2),.dout(w_dff_B_ucI4AD7R8_2),.clk(gclk));
	jdff dff_B_2AtVjVru3_2(.din(w_dff_B_ucI4AD7R8_2),.dout(w_dff_B_2AtVjVru3_2),.clk(gclk));
	jdff dff_B_wi2x7uf67_2(.din(w_dff_B_2AtVjVru3_2),.dout(w_dff_B_wi2x7uf67_2),.clk(gclk));
	jdff dff_B_oWb3rbPn0_2(.din(w_dff_B_wi2x7uf67_2),.dout(w_dff_B_oWb3rbPn0_2),.clk(gclk));
	jdff dff_B_GAs5Apbm0_2(.din(w_dff_B_oWb3rbPn0_2),.dout(w_dff_B_GAs5Apbm0_2),.clk(gclk));
	jdff dff_B_89P7xuT70_2(.din(w_dff_B_GAs5Apbm0_2),.dout(w_dff_B_89P7xuT70_2),.clk(gclk));
	jdff dff_B_UzxMRUuo1_2(.din(w_dff_B_89P7xuT70_2),.dout(w_dff_B_UzxMRUuo1_2),.clk(gclk));
	jdff dff_B_UtvfWYMs8_2(.din(w_dff_B_UzxMRUuo1_2),.dout(w_dff_B_UtvfWYMs8_2),.clk(gclk));
	jdff dff_B_vTVOUeVN0_2(.din(w_dff_B_UtvfWYMs8_2),.dout(w_dff_B_vTVOUeVN0_2),.clk(gclk));
	jdff dff_B_tnw1i2EO3_2(.din(w_dff_B_vTVOUeVN0_2),.dout(w_dff_B_tnw1i2EO3_2),.clk(gclk));
	jdff dff_B_utnlB5gF5_2(.din(w_dff_B_tnw1i2EO3_2),.dout(w_dff_B_utnlB5gF5_2),.clk(gclk));
	jdff dff_B_0jtgF9Pa2_2(.din(w_dff_B_utnlB5gF5_2),.dout(w_dff_B_0jtgF9Pa2_2),.clk(gclk));
	jdff dff_B_ToWwYuCP9_2(.din(w_dff_B_0jtgF9Pa2_2),.dout(w_dff_B_ToWwYuCP9_2),.clk(gclk));
	jdff dff_B_3ElCogYp8_2(.din(w_dff_B_ToWwYuCP9_2),.dout(w_dff_B_3ElCogYp8_2),.clk(gclk));
	jdff dff_B_da2by9p20_2(.din(w_dff_B_3ElCogYp8_2),.dout(w_dff_B_da2by9p20_2),.clk(gclk));
	jdff dff_B_XiqeBoTE8_2(.din(w_dff_B_da2by9p20_2),.dout(w_dff_B_XiqeBoTE8_2),.clk(gclk));
	jdff dff_B_7PW0mHnc6_2(.din(w_dff_B_XiqeBoTE8_2),.dout(w_dff_B_7PW0mHnc6_2),.clk(gclk));
	jdff dff_B_LvrPfIdk7_2(.din(w_dff_B_7PW0mHnc6_2),.dout(w_dff_B_LvrPfIdk7_2),.clk(gclk));
	jdff dff_B_DFZ8lVSh3_2(.din(w_dff_B_LvrPfIdk7_2),.dout(w_dff_B_DFZ8lVSh3_2),.clk(gclk));
	jdff dff_B_pXOmb06k6_2(.din(w_dff_B_DFZ8lVSh3_2),.dout(w_dff_B_pXOmb06k6_2),.clk(gclk));
	jdff dff_B_FrGaBkqP7_2(.din(w_dff_B_pXOmb06k6_2),.dout(w_dff_B_FrGaBkqP7_2),.clk(gclk));
	jdff dff_B_DRKSCwm95_2(.din(w_dff_B_FrGaBkqP7_2),.dout(w_dff_B_DRKSCwm95_2),.clk(gclk));
	jdff dff_B_CfL2HHFE9_2(.din(w_dff_B_DRKSCwm95_2),.dout(w_dff_B_CfL2HHFE9_2),.clk(gclk));
	jdff dff_B_R1wbpUy81_2(.din(w_dff_B_CfL2HHFE9_2),.dout(w_dff_B_R1wbpUy81_2),.clk(gclk));
	jdff dff_B_u2A0zG2l8_2(.din(w_dff_B_R1wbpUy81_2),.dout(w_dff_B_u2A0zG2l8_2),.clk(gclk));
	jdff dff_B_bGYF4gsT3_2(.din(w_dff_B_u2A0zG2l8_2),.dout(w_dff_B_bGYF4gsT3_2),.clk(gclk));
	jdff dff_B_5DYZp9407_2(.din(w_dff_B_bGYF4gsT3_2),.dout(w_dff_B_5DYZp9407_2),.clk(gclk));
	jdff dff_B_n49NGnNO7_2(.din(w_dff_B_5DYZp9407_2),.dout(w_dff_B_n49NGnNO7_2),.clk(gclk));
	jdff dff_B_0p1ewIGR8_2(.din(w_dff_B_n49NGnNO7_2),.dout(w_dff_B_0p1ewIGR8_2),.clk(gclk));
	jdff dff_B_pee5vlDs6_2(.din(w_dff_B_0p1ewIGR8_2),.dout(w_dff_B_pee5vlDs6_2),.clk(gclk));
	jdff dff_B_Nu1GZGt17_2(.din(w_dff_B_pee5vlDs6_2),.dout(w_dff_B_Nu1GZGt17_2),.clk(gclk));
	jdff dff_B_04UzHpm74_2(.din(w_dff_B_Nu1GZGt17_2),.dout(w_dff_B_04UzHpm74_2),.clk(gclk));
	jdff dff_B_vc5rPiNp8_2(.din(w_dff_B_04UzHpm74_2),.dout(w_dff_B_vc5rPiNp8_2),.clk(gclk));
	jdff dff_B_IIrK9S8e4_1(.din(n1778),.dout(w_dff_B_IIrK9S8e4_1),.clk(gclk));
	jdff dff_B_KInWw2Ze8_1(.din(w_dff_B_IIrK9S8e4_1),.dout(w_dff_B_KInWw2Ze8_1),.clk(gclk));
	jdff dff_B_NvrZTT2W4_2(.din(n1777),.dout(w_dff_B_NvrZTT2W4_2),.clk(gclk));
	jdff dff_B_De0raXHb8_2(.din(w_dff_B_NvrZTT2W4_2),.dout(w_dff_B_De0raXHb8_2),.clk(gclk));
	jdff dff_B_8ufEoUho1_2(.din(w_dff_B_De0raXHb8_2),.dout(w_dff_B_8ufEoUho1_2),.clk(gclk));
	jdff dff_B_WfiKk9ED1_2(.din(w_dff_B_8ufEoUho1_2),.dout(w_dff_B_WfiKk9ED1_2),.clk(gclk));
	jdff dff_B_RR8CyNt29_2(.din(w_dff_B_WfiKk9ED1_2),.dout(w_dff_B_RR8CyNt29_2),.clk(gclk));
	jdff dff_B_fwbLCIO69_2(.din(w_dff_B_RR8CyNt29_2),.dout(w_dff_B_fwbLCIO69_2),.clk(gclk));
	jdff dff_B_bIZv65pX6_2(.din(w_dff_B_fwbLCIO69_2),.dout(w_dff_B_bIZv65pX6_2),.clk(gclk));
	jdff dff_B_WlTNzLHA3_2(.din(w_dff_B_bIZv65pX6_2),.dout(w_dff_B_WlTNzLHA3_2),.clk(gclk));
	jdff dff_B_bZc4q3YB1_2(.din(w_dff_B_WlTNzLHA3_2),.dout(w_dff_B_bZc4q3YB1_2),.clk(gclk));
	jdff dff_B_IhhxcOd89_2(.din(w_dff_B_bZc4q3YB1_2),.dout(w_dff_B_IhhxcOd89_2),.clk(gclk));
	jdff dff_B_bvdpctnm3_2(.din(w_dff_B_IhhxcOd89_2),.dout(w_dff_B_bvdpctnm3_2),.clk(gclk));
	jdff dff_B_GHdlnLmj6_2(.din(w_dff_B_bvdpctnm3_2),.dout(w_dff_B_GHdlnLmj6_2),.clk(gclk));
	jdff dff_B_mtzGz4AY3_2(.din(w_dff_B_GHdlnLmj6_2),.dout(w_dff_B_mtzGz4AY3_2),.clk(gclk));
	jdff dff_B_QGx8HGMa5_2(.din(w_dff_B_mtzGz4AY3_2),.dout(w_dff_B_QGx8HGMa5_2),.clk(gclk));
	jdff dff_B_L91D3la25_2(.din(w_dff_B_QGx8HGMa5_2),.dout(w_dff_B_L91D3la25_2),.clk(gclk));
	jdff dff_B_CZ8Y5NwY2_2(.din(w_dff_B_L91D3la25_2),.dout(w_dff_B_CZ8Y5NwY2_2),.clk(gclk));
	jdff dff_B_tpEbFM308_2(.din(w_dff_B_CZ8Y5NwY2_2),.dout(w_dff_B_tpEbFM308_2),.clk(gclk));
	jdff dff_B_9NpQc4t86_2(.din(w_dff_B_tpEbFM308_2),.dout(w_dff_B_9NpQc4t86_2),.clk(gclk));
	jdff dff_B_YCFMKMzF9_2(.din(w_dff_B_9NpQc4t86_2),.dout(w_dff_B_YCFMKMzF9_2),.clk(gclk));
	jdff dff_B_B3EHuTda0_2(.din(w_dff_B_YCFMKMzF9_2),.dout(w_dff_B_B3EHuTda0_2),.clk(gclk));
	jdff dff_B_JhLcc2yb1_2(.din(w_dff_B_B3EHuTda0_2),.dout(w_dff_B_JhLcc2yb1_2),.clk(gclk));
	jdff dff_B_mquBrRvZ8_2(.din(w_dff_B_JhLcc2yb1_2),.dout(w_dff_B_mquBrRvZ8_2),.clk(gclk));
	jdff dff_B_QaQo3S3Q2_2(.din(w_dff_B_mquBrRvZ8_2),.dout(w_dff_B_QaQo3S3Q2_2),.clk(gclk));
	jdff dff_B_3VG0ynRn9_2(.din(w_dff_B_QaQo3S3Q2_2),.dout(w_dff_B_3VG0ynRn9_2),.clk(gclk));
	jdff dff_B_t2D9BH491_2(.din(w_dff_B_3VG0ynRn9_2),.dout(w_dff_B_t2D9BH491_2),.clk(gclk));
	jdff dff_B_wZwMO1n63_2(.din(w_dff_B_t2D9BH491_2),.dout(w_dff_B_wZwMO1n63_2),.clk(gclk));
	jdff dff_B_CSEUDD1e1_2(.din(w_dff_B_wZwMO1n63_2),.dout(w_dff_B_CSEUDD1e1_2),.clk(gclk));
	jdff dff_B_saawBkeW2_2(.din(w_dff_B_CSEUDD1e1_2),.dout(w_dff_B_saawBkeW2_2),.clk(gclk));
	jdff dff_B_UemBGa1j1_2(.din(w_dff_B_saawBkeW2_2),.dout(w_dff_B_UemBGa1j1_2),.clk(gclk));
	jdff dff_B_98nErRHJ8_2(.din(w_dff_B_UemBGa1j1_2),.dout(w_dff_B_98nErRHJ8_2),.clk(gclk));
	jdff dff_B_11LC3EgX4_2(.din(w_dff_B_98nErRHJ8_2),.dout(w_dff_B_11LC3EgX4_2),.clk(gclk));
	jdff dff_B_MjhrhxhZ0_2(.din(w_dff_B_11LC3EgX4_2),.dout(w_dff_B_MjhrhxhZ0_2),.clk(gclk));
	jdff dff_B_EZjFtKMT9_2(.din(w_dff_B_MjhrhxhZ0_2),.dout(w_dff_B_EZjFtKMT9_2),.clk(gclk));
	jdff dff_B_jdkNWGqi4_2(.din(w_dff_B_EZjFtKMT9_2),.dout(w_dff_B_jdkNWGqi4_2),.clk(gclk));
	jdff dff_B_BQuO9eMB8_2(.din(w_dff_B_jdkNWGqi4_2),.dout(w_dff_B_BQuO9eMB8_2),.clk(gclk));
	jdff dff_B_qwHNU55a6_2(.din(w_dff_B_BQuO9eMB8_2),.dout(w_dff_B_qwHNU55a6_2),.clk(gclk));
	jdff dff_B_iciNOIY51_2(.din(w_dff_B_qwHNU55a6_2),.dout(w_dff_B_iciNOIY51_2),.clk(gclk));
	jdff dff_B_S48muyIX0_2(.din(w_dff_B_iciNOIY51_2),.dout(w_dff_B_S48muyIX0_2),.clk(gclk));
	jdff dff_B_K7cPHnl28_2(.din(w_dff_B_S48muyIX0_2),.dout(w_dff_B_K7cPHnl28_2),.clk(gclk));
	jdff dff_B_f6nEfctv1_2(.din(w_dff_B_K7cPHnl28_2),.dout(w_dff_B_f6nEfctv1_2),.clk(gclk));
	jdff dff_B_IDk7U9bE4_2(.din(w_dff_B_f6nEfctv1_2),.dout(w_dff_B_IDk7U9bE4_2),.clk(gclk));
	jdff dff_B_e6LfYu1o8_2(.din(w_dff_B_IDk7U9bE4_2),.dout(w_dff_B_e6LfYu1o8_2),.clk(gclk));
	jdff dff_B_NxnBI4752_2(.din(w_dff_B_e6LfYu1o8_2),.dout(w_dff_B_NxnBI4752_2),.clk(gclk));
	jdff dff_B_ExZacyRm6_2(.din(w_dff_B_NxnBI4752_2),.dout(w_dff_B_ExZacyRm6_2),.clk(gclk));
	jdff dff_B_x5WR6gah7_2(.din(w_dff_B_ExZacyRm6_2),.dout(w_dff_B_x5WR6gah7_2),.clk(gclk));
	jdff dff_B_PaHaOLhD0_2(.din(w_dff_B_x5WR6gah7_2),.dout(w_dff_B_PaHaOLhD0_2),.clk(gclk));
	jdff dff_B_0IALB7UA1_2(.din(w_dff_B_PaHaOLhD0_2),.dout(w_dff_B_0IALB7UA1_2),.clk(gclk));
	jdff dff_B_NBVbAG3x8_2(.din(w_dff_B_0IALB7UA1_2),.dout(w_dff_B_NBVbAG3x8_2),.clk(gclk));
	jdff dff_B_PIWEmWL32_2(.din(w_dff_B_NBVbAG3x8_2),.dout(w_dff_B_PIWEmWL32_2),.clk(gclk));
	jdff dff_B_iImEmESC3_2(.din(n1776),.dout(w_dff_B_iImEmESC3_2),.clk(gclk));
	jdff dff_B_ioW0lsdf2_2(.din(w_dff_B_iImEmESC3_2),.dout(w_dff_B_ioW0lsdf2_2),.clk(gclk));
	jdff dff_B_b8avPETQ4_2(.din(w_dff_B_ioW0lsdf2_2),.dout(w_dff_B_b8avPETQ4_2),.clk(gclk));
	jdff dff_B_Gl93NYTU5_2(.din(w_dff_B_b8avPETQ4_2),.dout(w_dff_B_Gl93NYTU5_2),.clk(gclk));
	jdff dff_B_Bv4Iw56G1_2(.din(w_dff_B_Gl93NYTU5_2),.dout(w_dff_B_Bv4Iw56G1_2),.clk(gclk));
	jdff dff_B_NFDbYbnJ8_2(.din(w_dff_B_Bv4Iw56G1_2),.dout(w_dff_B_NFDbYbnJ8_2),.clk(gclk));
	jdff dff_B_ZHjLGGQq6_2(.din(w_dff_B_NFDbYbnJ8_2),.dout(w_dff_B_ZHjLGGQq6_2),.clk(gclk));
	jdff dff_B_vHlc8EKC4_2(.din(w_dff_B_ZHjLGGQq6_2),.dout(w_dff_B_vHlc8EKC4_2),.clk(gclk));
	jdff dff_B_aN7Pusvh5_2(.din(w_dff_B_vHlc8EKC4_2),.dout(w_dff_B_aN7Pusvh5_2),.clk(gclk));
	jdff dff_B_ZJeEpx7f1_2(.din(w_dff_B_aN7Pusvh5_2),.dout(w_dff_B_ZJeEpx7f1_2),.clk(gclk));
	jdff dff_B_hNeWZUh13_2(.din(w_dff_B_ZJeEpx7f1_2),.dout(w_dff_B_hNeWZUh13_2),.clk(gclk));
	jdff dff_B_Wv0oDHv37_2(.din(w_dff_B_hNeWZUh13_2),.dout(w_dff_B_Wv0oDHv37_2),.clk(gclk));
	jdff dff_B_DY2AlFEn3_2(.din(w_dff_B_Wv0oDHv37_2),.dout(w_dff_B_DY2AlFEn3_2),.clk(gclk));
	jdff dff_B_AxjmYavE4_2(.din(w_dff_B_DY2AlFEn3_2),.dout(w_dff_B_AxjmYavE4_2),.clk(gclk));
	jdff dff_B_OFJpi7aV4_2(.din(w_dff_B_AxjmYavE4_2),.dout(w_dff_B_OFJpi7aV4_2),.clk(gclk));
	jdff dff_B_viHaDg3n8_2(.din(w_dff_B_OFJpi7aV4_2),.dout(w_dff_B_viHaDg3n8_2),.clk(gclk));
	jdff dff_B_6KAxKkF52_2(.din(w_dff_B_viHaDg3n8_2),.dout(w_dff_B_6KAxKkF52_2),.clk(gclk));
	jdff dff_B_WvUy9Xgj7_2(.din(w_dff_B_6KAxKkF52_2),.dout(w_dff_B_WvUy9Xgj7_2),.clk(gclk));
	jdff dff_B_yjPwEgj65_2(.din(w_dff_B_WvUy9Xgj7_2),.dout(w_dff_B_yjPwEgj65_2),.clk(gclk));
	jdff dff_B_ceBBZEjj7_2(.din(w_dff_B_yjPwEgj65_2),.dout(w_dff_B_ceBBZEjj7_2),.clk(gclk));
	jdff dff_B_xn6GsXHo8_2(.din(w_dff_B_ceBBZEjj7_2),.dout(w_dff_B_xn6GsXHo8_2),.clk(gclk));
	jdff dff_B_cGsJNLJ77_2(.din(w_dff_B_xn6GsXHo8_2),.dout(w_dff_B_cGsJNLJ77_2),.clk(gclk));
	jdff dff_B_dibxXs7f9_2(.din(w_dff_B_cGsJNLJ77_2),.dout(w_dff_B_dibxXs7f9_2),.clk(gclk));
	jdff dff_B_BVXcjW8O3_2(.din(w_dff_B_dibxXs7f9_2),.dout(w_dff_B_BVXcjW8O3_2),.clk(gclk));
	jdff dff_B_WHKlnkAW0_2(.din(w_dff_B_BVXcjW8O3_2),.dout(w_dff_B_WHKlnkAW0_2),.clk(gclk));
	jdff dff_B_JS1aW1tV3_2(.din(w_dff_B_WHKlnkAW0_2),.dout(w_dff_B_JS1aW1tV3_2),.clk(gclk));
	jdff dff_B_TOrT2Hal9_2(.din(w_dff_B_JS1aW1tV3_2),.dout(w_dff_B_TOrT2Hal9_2),.clk(gclk));
	jdff dff_B_edlU4s8A5_2(.din(w_dff_B_TOrT2Hal9_2),.dout(w_dff_B_edlU4s8A5_2),.clk(gclk));
	jdff dff_B_N2b6l1Lb9_2(.din(w_dff_B_edlU4s8A5_2),.dout(w_dff_B_N2b6l1Lb9_2),.clk(gclk));
	jdff dff_B_1Q8PyZCg0_2(.din(w_dff_B_N2b6l1Lb9_2),.dout(w_dff_B_1Q8PyZCg0_2),.clk(gclk));
	jdff dff_B_Ryb6VMY08_2(.din(w_dff_B_1Q8PyZCg0_2),.dout(w_dff_B_Ryb6VMY08_2),.clk(gclk));
	jdff dff_B_mL8KOsxt8_2(.din(w_dff_B_Ryb6VMY08_2),.dout(w_dff_B_mL8KOsxt8_2),.clk(gclk));
	jdff dff_B_Lqpb9cmN6_2(.din(w_dff_B_mL8KOsxt8_2),.dout(w_dff_B_Lqpb9cmN6_2),.clk(gclk));
	jdff dff_B_we1dICRd6_2(.din(w_dff_B_Lqpb9cmN6_2),.dout(w_dff_B_we1dICRd6_2),.clk(gclk));
	jdff dff_B_hlQ9slZK8_2(.din(w_dff_B_we1dICRd6_2),.dout(w_dff_B_hlQ9slZK8_2),.clk(gclk));
	jdff dff_B_OTAyjO1U2_2(.din(w_dff_B_hlQ9slZK8_2),.dout(w_dff_B_OTAyjO1U2_2),.clk(gclk));
	jdff dff_B_0t2RPjdF7_2(.din(w_dff_B_OTAyjO1U2_2),.dout(w_dff_B_0t2RPjdF7_2),.clk(gclk));
	jdff dff_B_VNckG46C8_2(.din(w_dff_B_0t2RPjdF7_2),.dout(w_dff_B_VNckG46C8_2),.clk(gclk));
	jdff dff_B_5AnD0mq88_2(.din(w_dff_B_VNckG46C8_2),.dout(w_dff_B_5AnD0mq88_2),.clk(gclk));
	jdff dff_B_64R7jRtM0_2(.din(w_dff_B_5AnD0mq88_2),.dout(w_dff_B_64R7jRtM0_2),.clk(gclk));
	jdff dff_B_yZFX5zYs1_2(.din(w_dff_B_64R7jRtM0_2),.dout(w_dff_B_yZFX5zYs1_2),.clk(gclk));
	jdff dff_B_rat0vrnm5_2(.din(w_dff_B_yZFX5zYs1_2),.dout(w_dff_B_rat0vrnm5_2),.clk(gclk));
	jdff dff_B_cjrXDAJm2_2(.din(w_dff_B_rat0vrnm5_2),.dout(w_dff_B_cjrXDAJm2_2),.clk(gclk));
	jdff dff_B_SX2lUEYc6_2(.din(w_dff_B_cjrXDAJm2_2),.dout(w_dff_B_SX2lUEYc6_2),.clk(gclk));
	jdff dff_B_fP9B9w7o9_2(.din(w_dff_B_SX2lUEYc6_2),.dout(w_dff_B_fP9B9w7o9_2),.clk(gclk));
	jdff dff_B_YdQuE3et0_2(.din(w_dff_B_fP9B9w7o9_2),.dout(w_dff_B_YdQuE3et0_2),.clk(gclk));
	jdff dff_B_mDd0gWwf2_2(.din(w_dff_B_YdQuE3et0_2),.dout(w_dff_B_mDd0gWwf2_2),.clk(gclk));
	jdff dff_B_hEINZUw46_2(.din(w_dff_B_mDd0gWwf2_2),.dout(w_dff_B_hEINZUw46_2),.clk(gclk));
	jdff dff_B_4S6Z5FUH4_2(.din(w_dff_B_hEINZUw46_2),.dout(w_dff_B_4S6Z5FUH4_2),.clk(gclk));
	jdff dff_B_GAvzG52H4_2(.din(w_dff_B_4S6Z5FUH4_2),.dout(w_dff_B_GAvzG52H4_2),.clk(gclk));
	jdff dff_B_Lam9kCm25_2(.din(w_dff_B_GAvzG52H4_2),.dout(w_dff_B_Lam9kCm25_2),.clk(gclk));
	jdff dff_B_962kAxAN4_2(.din(n1775),.dout(w_dff_B_962kAxAN4_2),.clk(gclk));
	jdff dff_B_w3zmnl6r0_1(.din(n1773),.dout(w_dff_B_w3zmnl6r0_1),.clk(gclk));
	jdff dff_B_doL0YCC16_2(.din(n1744),.dout(w_dff_B_doL0YCC16_2),.clk(gclk));
	jdff dff_B_PO80Hljs3_2(.din(w_dff_B_doL0YCC16_2),.dout(w_dff_B_PO80Hljs3_2),.clk(gclk));
	jdff dff_B_tAoJnxxI7_2(.din(w_dff_B_PO80Hljs3_2),.dout(w_dff_B_tAoJnxxI7_2),.clk(gclk));
	jdff dff_B_I9tNYdXt6_2(.din(w_dff_B_tAoJnxxI7_2),.dout(w_dff_B_I9tNYdXt6_2),.clk(gclk));
	jdff dff_B_xVYa1lsO8_2(.din(w_dff_B_I9tNYdXt6_2),.dout(w_dff_B_xVYa1lsO8_2),.clk(gclk));
	jdff dff_B_eGZKkaC31_2(.din(w_dff_B_xVYa1lsO8_2),.dout(w_dff_B_eGZKkaC31_2),.clk(gclk));
	jdff dff_B_ag97yKCq3_2(.din(w_dff_B_eGZKkaC31_2),.dout(w_dff_B_ag97yKCq3_2),.clk(gclk));
	jdff dff_B_r5LZPEN60_2(.din(w_dff_B_ag97yKCq3_2),.dout(w_dff_B_r5LZPEN60_2),.clk(gclk));
	jdff dff_B_8GMA7ssn8_2(.din(w_dff_B_r5LZPEN60_2),.dout(w_dff_B_8GMA7ssn8_2),.clk(gclk));
	jdff dff_B_HZSYmuGw2_2(.din(w_dff_B_8GMA7ssn8_2),.dout(w_dff_B_HZSYmuGw2_2),.clk(gclk));
	jdff dff_B_zpNYHYiv5_2(.din(w_dff_B_HZSYmuGw2_2),.dout(w_dff_B_zpNYHYiv5_2),.clk(gclk));
	jdff dff_B_GK7qFWiW3_2(.din(w_dff_B_zpNYHYiv5_2),.dout(w_dff_B_GK7qFWiW3_2),.clk(gclk));
	jdff dff_B_Tv4ccQm50_2(.din(w_dff_B_GK7qFWiW3_2),.dout(w_dff_B_Tv4ccQm50_2),.clk(gclk));
	jdff dff_B_lx9X790e1_2(.din(w_dff_B_Tv4ccQm50_2),.dout(w_dff_B_lx9X790e1_2),.clk(gclk));
	jdff dff_B_69GtdHYW0_2(.din(w_dff_B_lx9X790e1_2),.dout(w_dff_B_69GtdHYW0_2),.clk(gclk));
	jdff dff_B_H8BvjoBO4_2(.din(w_dff_B_69GtdHYW0_2),.dout(w_dff_B_H8BvjoBO4_2),.clk(gclk));
	jdff dff_B_U0rRh0O24_2(.din(w_dff_B_H8BvjoBO4_2),.dout(w_dff_B_U0rRh0O24_2),.clk(gclk));
	jdff dff_B_Yft8nIWx2_2(.din(w_dff_B_U0rRh0O24_2),.dout(w_dff_B_Yft8nIWx2_2),.clk(gclk));
	jdff dff_B_TULcQlcD6_2(.din(w_dff_B_Yft8nIWx2_2),.dout(w_dff_B_TULcQlcD6_2),.clk(gclk));
	jdff dff_B_I6nnn3an5_2(.din(w_dff_B_TULcQlcD6_2),.dout(w_dff_B_I6nnn3an5_2),.clk(gclk));
	jdff dff_B_4UavkAXR7_2(.din(w_dff_B_I6nnn3an5_2),.dout(w_dff_B_4UavkAXR7_2),.clk(gclk));
	jdff dff_B_meDrfdmn5_2(.din(w_dff_B_4UavkAXR7_2),.dout(w_dff_B_meDrfdmn5_2),.clk(gclk));
	jdff dff_B_mZmAkMTK6_2(.din(w_dff_B_meDrfdmn5_2),.dout(w_dff_B_mZmAkMTK6_2),.clk(gclk));
	jdff dff_B_DWy7vFSZ3_2(.din(w_dff_B_mZmAkMTK6_2),.dout(w_dff_B_DWy7vFSZ3_2),.clk(gclk));
	jdff dff_B_u9cOpx384_2(.din(w_dff_B_DWy7vFSZ3_2),.dout(w_dff_B_u9cOpx384_2),.clk(gclk));
	jdff dff_B_PrUIrbZJ0_2(.din(w_dff_B_u9cOpx384_2),.dout(w_dff_B_PrUIrbZJ0_2),.clk(gclk));
	jdff dff_B_d0RyFGEL1_2(.din(w_dff_B_PrUIrbZJ0_2),.dout(w_dff_B_d0RyFGEL1_2),.clk(gclk));
	jdff dff_B_w4FEVQiI4_2(.din(w_dff_B_d0RyFGEL1_2),.dout(w_dff_B_w4FEVQiI4_2),.clk(gclk));
	jdff dff_B_2V7g2ufw7_2(.din(w_dff_B_w4FEVQiI4_2),.dout(w_dff_B_2V7g2ufw7_2),.clk(gclk));
	jdff dff_B_qmcX0Slb6_2(.din(w_dff_B_2V7g2ufw7_2),.dout(w_dff_B_qmcX0Slb6_2),.clk(gclk));
	jdff dff_B_bi3efb5G8_2(.din(w_dff_B_qmcX0Slb6_2),.dout(w_dff_B_bi3efb5G8_2),.clk(gclk));
	jdff dff_B_GGyeunjO4_2(.din(w_dff_B_bi3efb5G8_2),.dout(w_dff_B_GGyeunjO4_2),.clk(gclk));
	jdff dff_B_YYY4kqJg7_2(.din(w_dff_B_GGyeunjO4_2),.dout(w_dff_B_YYY4kqJg7_2),.clk(gclk));
	jdff dff_B_c2rmAP3l6_2(.din(w_dff_B_YYY4kqJg7_2),.dout(w_dff_B_c2rmAP3l6_2),.clk(gclk));
	jdff dff_B_usUNnHza6_2(.din(w_dff_B_c2rmAP3l6_2),.dout(w_dff_B_usUNnHza6_2),.clk(gclk));
	jdff dff_B_P4zJadhL9_2(.din(w_dff_B_usUNnHza6_2),.dout(w_dff_B_P4zJadhL9_2),.clk(gclk));
	jdff dff_B_cc8eC8nn5_2(.din(w_dff_B_P4zJadhL9_2),.dout(w_dff_B_cc8eC8nn5_2),.clk(gclk));
	jdff dff_B_A6n8MjoI5_2(.din(w_dff_B_cc8eC8nn5_2),.dout(w_dff_B_A6n8MjoI5_2),.clk(gclk));
	jdff dff_B_meZHDjPW6_2(.din(w_dff_B_A6n8MjoI5_2),.dout(w_dff_B_meZHDjPW6_2),.clk(gclk));
	jdff dff_B_hYYQqhYG9_2(.din(w_dff_B_meZHDjPW6_2),.dout(w_dff_B_hYYQqhYG9_2),.clk(gclk));
	jdff dff_B_h5C3FUQk0_2(.din(w_dff_B_hYYQqhYG9_2),.dout(w_dff_B_h5C3FUQk0_2),.clk(gclk));
	jdff dff_B_hgpcHUij2_2(.din(w_dff_B_h5C3FUQk0_2),.dout(w_dff_B_hgpcHUij2_2),.clk(gclk));
	jdff dff_B_waOVNIE37_2(.din(w_dff_B_hgpcHUij2_2),.dout(w_dff_B_waOVNIE37_2),.clk(gclk));
	jdff dff_B_xnqK7Byh6_2(.din(w_dff_B_waOVNIE37_2),.dout(w_dff_B_xnqK7Byh6_2),.clk(gclk));
	jdff dff_B_p7B7sbbP7_2(.din(w_dff_B_xnqK7Byh6_2),.dout(w_dff_B_p7B7sbbP7_2),.clk(gclk));
	jdff dff_B_DcLUZTiI2_2(.din(w_dff_B_p7B7sbbP7_2),.dout(w_dff_B_DcLUZTiI2_2),.clk(gclk));
	jdff dff_B_G20dCVcg1_2(.din(w_dff_B_DcLUZTiI2_2),.dout(w_dff_B_G20dCVcg1_2),.clk(gclk));
	jdff dff_B_Gqhqk55Q6_2(.din(w_dff_B_G20dCVcg1_2),.dout(w_dff_B_Gqhqk55Q6_2),.clk(gclk));
	jdff dff_B_KSBx9hgd8_1(.din(n1750),.dout(w_dff_B_KSBx9hgd8_1),.clk(gclk));
	jdff dff_B_HuYfgTST5_1(.din(w_dff_B_KSBx9hgd8_1),.dout(w_dff_B_HuYfgTST5_1),.clk(gclk));
	jdff dff_B_NRarIm481_2(.din(n1749),.dout(w_dff_B_NRarIm481_2),.clk(gclk));
	jdff dff_B_bNkLPfhj3_2(.din(w_dff_B_NRarIm481_2),.dout(w_dff_B_bNkLPfhj3_2),.clk(gclk));
	jdff dff_B_HsTrgkDH7_2(.din(w_dff_B_bNkLPfhj3_2),.dout(w_dff_B_HsTrgkDH7_2),.clk(gclk));
	jdff dff_B_WJ1K3ROM2_2(.din(w_dff_B_HsTrgkDH7_2),.dout(w_dff_B_WJ1K3ROM2_2),.clk(gclk));
	jdff dff_B_Sy2gkp6g9_2(.din(w_dff_B_WJ1K3ROM2_2),.dout(w_dff_B_Sy2gkp6g9_2),.clk(gclk));
	jdff dff_B_vQw3N8xP1_2(.din(w_dff_B_Sy2gkp6g9_2),.dout(w_dff_B_vQw3N8xP1_2),.clk(gclk));
	jdff dff_B_hu3d0up95_2(.din(w_dff_B_vQw3N8xP1_2),.dout(w_dff_B_hu3d0up95_2),.clk(gclk));
	jdff dff_B_bwTsxGle8_2(.din(w_dff_B_hu3d0up95_2),.dout(w_dff_B_bwTsxGle8_2),.clk(gclk));
	jdff dff_B_ZVHMzRyU3_2(.din(w_dff_B_bwTsxGle8_2),.dout(w_dff_B_ZVHMzRyU3_2),.clk(gclk));
	jdff dff_B_Aa3Ruav88_2(.din(w_dff_B_ZVHMzRyU3_2),.dout(w_dff_B_Aa3Ruav88_2),.clk(gclk));
	jdff dff_B_1hOm2KMg3_2(.din(w_dff_B_Aa3Ruav88_2),.dout(w_dff_B_1hOm2KMg3_2),.clk(gclk));
	jdff dff_B_PstwEAOL5_2(.din(w_dff_B_1hOm2KMg3_2),.dout(w_dff_B_PstwEAOL5_2),.clk(gclk));
	jdff dff_B_SBC3Jut87_2(.din(w_dff_B_PstwEAOL5_2),.dout(w_dff_B_SBC3Jut87_2),.clk(gclk));
	jdff dff_B_1x4BOWQm9_2(.din(w_dff_B_SBC3Jut87_2),.dout(w_dff_B_1x4BOWQm9_2),.clk(gclk));
	jdff dff_B_FPk5bM1R3_2(.din(w_dff_B_1x4BOWQm9_2),.dout(w_dff_B_FPk5bM1R3_2),.clk(gclk));
	jdff dff_B_AZNJ5v4x4_2(.din(w_dff_B_FPk5bM1R3_2),.dout(w_dff_B_AZNJ5v4x4_2),.clk(gclk));
	jdff dff_B_TCdxf6yk6_2(.din(w_dff_B_AZNJ5v4x4_2),.dout(w_dff_B_TCdxf6yk6_2),.clk(gclk));
	jdff dff_B_13eA2AlI8_2(.din(w_dff_B_TCdxf6yk6_2),.dout(w_dff_B_13eA2AlI8_2),.clk(gclk));
	jdff dff_B_BneWj0V76_2(.din(w_dff_B_13eA2AlI8_2),.dout(w_dff_B_BneWj0V76_2),.clk(gclk));
	jdff dff_B_4GUV5hjH8_2(.din(w_dff_B_BneWj0V76_2),.dout(w_dff_B_4GUV5hjH8_2),.clk(gclk));
	jdff dff_B_GytnC5GA3_2(.din(w_dff_B_4GUV5hjH8_2),.dout(w_dff_B_GytnC5GA3_2),.clk(gclk));
	jdff dff_B_vgouNKQR2_2(.din(w_dff_B_GytnC5GA3_2),.dout(w_dff_B_vgouNKQR2_2),.clk(gclk));
	jdff dff_B_ARMT9Ao40_2(.din(w_dff_B_vgouNKQR2_2),.dout(w_dff_B_ARMT9Ao40_2),.clk(gclk));
	jdff dff_B_KyBIYozU9_2(.din(w_dff_B_ARMT9Ao40_2),.dout(w_dff_B_KyBIYozU9_2),.clk(gclk));
	jdff dff_B_EnifDq9L0_2(.din(w_dff_B_KyBIYozU9_2),.dout(w_dff_B_EnifDq9L0_2),.clk(gclk));
	jdff dff_B_6uVhiURb5_2(.din(w_dff_B_EnifDq9L0_2),.dout(w_dff_B_6uVhiURb5_2),.clk(gclk));
	jdff dff_B_doFOBq3C3_2(.din(w_dff_B_6uVhiURb5_2),.dout(w_dff_B_doFOBq3C3_2),.clk(gclk));
	jdff dff_B_PiALsGyr0_2(.din(w_dff_B_doFOBq3C3_2),.dout(w_dff_B_PiALsGyr0_2),.clk(gclk));
	jdff dff_B_edLLhkFo3_2(.din(w_dff_B_PiALsGyr0_2),.dout(w_dff_B_edLLhkFo3_2),.clk(gclk));
	jdff dff_B_SCokj42K4_2(.din(w_dff_B_edLLhkFo3_2),.dout(w_dff_B_SCokj42K4_2),.clk(gclk));
	jdff dff_B_1UDNjSQa5_2(.din(w_dff_B_SCokj42K4_2),.dout(w_dff_B_1UDNjSQa5_2),.clk(gclk));
	jdff dff_B_RcZVIRtI1_2(.din(w_dff_B_1UDNjSQa5_2),.dout(w_dff_B_RcZVIRtI1_2),.clk(gclk));
	jdff dff_B_l14ZrkSU1_2(.din(w_dff_B_RcZVIRtI1_2),.dout(w_dff_B_l14ZrkSU1_2),.clk(gclk));
	jdff dff_B_nsUfkMOK9_2(.din(w_dff_B_l14ZrkSU1_2),.dout(w_dff_B_nsUfkMOK9_2),.clk(gclk));
	jdff dff_B_iYkn4oJr6_2(.din(w_dff_B_nsUfkMOK9_2),.dout(w_dff_B_iYkn4oJr6_2),.clk(gclk));
	jdff dff_B_qY0Midl32_2(.din(w_dff_B_iYkn4oJr6_2),.dout(w_dff_B_qY0Midl32_2),.clk(gclk));
	jdff dff_B_YrCBHve83_2(.din(w_dff_B_qY0Midl32_2),.dout(w_dff_B_YrCBHve83_2),.clk(gclk));
	jdff dff_B_RzP8ufSE6_2(.din(w_dff_B_YrCBHve83_2),.dout(w_dff_B_RzP8ufSE6_2),.clk(gclk));
	jdff dff_B_3OaYdXdL7_2(.din(w_dff_B_RzP8ufSE6_2),.dout(w_dff_B_3OaYdXdL7_2),.clk(gclk));
	jdff dff_B_sIdjzXAe4_2(.din(w_dff_B_3OaYdXdL7_2),.dout(w_dff_B_sIdjzXAe4_2),.clk(gclk));
	jdff dff_B_iNTIn2dh8_2(.din(w_dff_B_sIdjzXAe4_2),.dout(w_dff_B_iNTIn2dh8_2),.clk(gclk));
	jdff dff_B_eJivWHm39_2(.din(w_dff_B_iNTIn2dh8_2),.dout(w_dff_B_eJivWHm39_2),.clk(gclk));
	jdff dff_B_OsKF9fUF4_2(.din(w_dff_B_eJivWHm39_2),.dout(w_dff_B_OsKF9fUF4_2),.clk(gclk));
	jdff dff_B_7atpzyXC7_2(.din(w_dff_B_OsKF9fUF4_2),.dout(w_dff_B_7atpzyXC7_2),.clk(gclk));
	jdff dff_B_f45WlC394_2(.din(w_dff_B_7atpzyXC7_2),.dout(w_dff_B_f45WlC394_2),.clk(gclk));
	jdff dff_B_hbLmOOlo1_2(.din(n1748),.dout(w_dff_B_hbLmOOlo1_2),.clk(gclk));
	jdff dff_B_YjCazqQQ3_2(.din(w_dff_B_hbLmOOlo1_2),.dout(w_dff_B_YjCazqQQ3_2),.clk(gclk));
	jdff dff_B_t1xsbvDJ0_2(.din(w_dff_B_YjCazqQQ3_2),.dout(w_dff_B_t1xsbvDJ0_2),.clk(gclk));
	jdff dff_B_ZgDqR1Pc8_2(.din(w_dff_B_t1xsbvDJ0_2),.dout(w_dff_B_ZgDqR1Pc8_2),.clk(gclk));
	jdff dff_B_jC8a5Z0i6_2(.din(w_dff_B_ZgDqR1Pc8_2),.dout(w_dff_B_jC8a5Z0i6_2),.clk(gclk));
	jdff dff_B_CtOC030R1_2(.din(w_dff_B_jC8a5Z0i6_2),.dout(w_dff_B_CtOC030R1_2),.clk(gclk));
	jdff dff_B_KvAkGQWQ1_2(.din(w_dff_B_CtOC030R1_2),.dout(w_dff_B_KvAkGQWQ1_2),.clk(gclk));
	jdff dff_B_GxhBTZam8_2(.din(w_dff_B_KvAkGQWQ1_2),.dout(w_dff_B_GxhBTZam8_2),.clk(gclk));
	jdff dff_B_hmvdfGcC1_2(.din(w_dff_B_GxhBTZam8_2),.dout(w_dff_B_hmvdfGcC1_2),.clk(gclk));
	jdff dff_B_WofEt4Ay7_2(.din(w_dff_B_hmvdfGcC1_2),.dout(w_dff_B_WofEt4Ay7_2),.clk(gclk));
	jdff dff_B_Dq5naBde3_2(.din(w_dff_B_WofEt4Ay7_2),.dout(w_dff_B_Dq5naBde3_2),.clk(gclk));
	jdff dff_B_tM7YFD2G3_2(.din(w_dff_B_Dq5naBde3_2),.dout(w_dff_B_tM7YFD2G3_2),.clk(gclk));
	jdff dff_B_ES7BqhXo1_2(.din(w_dff_B_tM7YFD2G3_2),.dout(w_dff_B_ES7BqhXo1_2),.clk(gclk));
	jdff dff_B_04aS6UYb8_2(.din(w_dff_B_ES7BqhXo1_2),.dout(w_dff_B_04aS6UYb8_2),.clk(gclk));
	jdff dff_B_bdSMKOBd5_2(.din(w_dff_B_04aS6UYb8_2),.dout(w_dff_B_bdSMKOBd5_2),.clk(gclk));
	jdff dff_B_mF38fRtk7_2(.din(w_dff_B_bdSMKOBd5_2),.dout(w_dff_B_mF38fRtk7_2),.clk(gclk));
	jdff dff_B_CutgmOio5_2(.din(w_dff_B_mF38fRtk7_2),.dout(w_dff_B_CutgmOio5_2),.clk(gclk));
	jdff dff_B_SjFGFVOn6_2(.din(w_dff_B_CutgmOio5_2),.dout(w_dff_B_SjFGFVOn6_2),.clk(gclk));
	jdff dff_B_L0kR6tUv3_2(.din(w_dff_B_SjFGFVOn6_2),.dout(w_dff_B_L0kR6tUv3_2),.clk(gclk));
	jdff dff_B_KI5fYqMu0_2(.din(w_dff_B_L0kR6tUv3_2),.dout(w_dff_B_KI5fYqMu0_2),.clk(gclk));
	jdff dff_B_iX5CW8J70_2(.din(w_dff_B_KI5fYqMu0_2),.dout(w_dff_B_iX5CW8J70_2),.clk(gclk));
	jdff dff_B_YDENOHEJ1_2(.din(w_dff_B_iX5CW8J70_2),.dout(w_dff_B_YDENOHEJ1_2),.clk(gclk));
	jdff dff_B_0aMEzOUL1_2(.din(w_dff_B_YDENOHEJ1_2),.dout(w_dff_B_0aMEzOUL1_2),.clk(gclk));
	jdff dff_B_xbVwIZ758_2(.din(w_dff_B_0aMEzOUL1_2),.dout(w_dff_B_xbVwIZ758_2),.clk(gclk));
	jdff dff_B_uCaqHB5Y1_2(.din(w_dff_B_xbVwIZ758_2),.dout(w_dff_B_uCaqHB5Y1_2),.clk(gclk));
	jdff dff_B_lnPNylQo6_2(.din(w_dff_B_uCaqHB5Y1_2),.dout(w_dff_B_lnPNylQo6_2),.clk(gclk));
	jdff dff_B_0edCn8cW7_2(.din(w_dff_B_lnPNylQo6_2),.dout(w_dff_B_0edCn8cW7_2),.clk(gclk));
	jdff dff_B_tlPVmLpa7_2(.din(w_dff_B_0edCn8cW7_2),.dout(w_dff_B_tlPVmLpa7_2),.clk(gclk));
	jdff dff_B_CrNf6jlH1_2(.din(w_dff_B_tlPVmLpa7_2),.dout(w_dff_B_CrNf6jlH1_2),.clk(gclk));
	jdff dff_B_5uTOTLMr7_2(.din(w_dff_B_CrNf6jlH1_2),.dout(w_dff_B_5uTOTLMr7_2),.clk(gclk));
	jdff dff_B_ayMTJqjq5_2(.din(w_dff_B_5uTOTLMr7_2),.dout(w_dff_B_ayMTJqjq5_2),.clk(gclk));
	jdff dff_B_ZJSE5A6u8_2(.din(w_dff_B_ayMTJqjq5_2),.dout(w_dff_B_ZJSE5A6u8_2),.clk(gclk));
	jdff dff_B_JOaVQVlj1_2(.din(w_dff_B_ZJSE5A6u8_2),.dout(w_dff_B_JOaVQVlj1_2),.clk(gclk));
	jdff dff_B_87GpAEat4_2(.din(w_dff_B_JOaVQVlj1_2),.dout(w_dff_B_87GpAEat4_2),.clk(gclk));
	jdff dff_B_R4e1XHKk7_2(.din(w_dff_B_87GpAEat4_2),.dout(w_dff_B_R4e1XHKk7_2),.clk(gclk));
	jdff dff_B_acDlqHo75_2(.din(w_dff_B_R4e1XHKk7_2),.dout(w_dff_B_acDlqHo75_2),.clk(gclk));
	jdff dff_B_tzmShRyT4_2(.din(w_dff_B_acDlqHo75_2),.dout(w_dff_B_tzmShRyT4_2),.clk(gclk));
	jdff dff_B_5gTMTT226_2(.din(w_dff_B_tzmShRyT4_2),.dout(w_dff_B_5gTMTT226_2),.clk(gclk));
	jdff dff_B_qf7enKqJ3_2(.din(w_dff_B_5gTMTT226_2),.dout(w_dff_B_qf7enKqJ3_2),.clk(gclk));
	jdff dff_B_SjS9F0V23_2(.din(w_dff_B_qf7enKqJ3_2),.dout(w_dff_B_SjS9F0V23_2),.clk(gclk));
	jdff dff_B_81SDYdzI1_2(.din(w_dff_B_SjS9F0V23_2),.dout(w_dff_B_81SDYdzI1_2),.clk(gclk));
	jdff dff_B_r6NlxRvS2_2(.din(w_dff_B_81SDYdzI1_2),.dout(w_dff_B_r6NlxRvS2_2),.clk(gclk));
	jdff dff_B_honvnWC47_2(.din(w_dff_B_r6NlxRvS2_2),.dout(w_dff_B_honvnWC47_2),.clk(gclk));
	jdff dff_B_Pm4lz2TE6_2(.din(w_dff_B_honvnWC47_2),.dout(w_dff_B_Pm4lz2TE6_2),.clk(gclk));
	jdff dff_B_qNm5DonE1_2(.din(w_dff_B_Pm4lz2TE6_2),.dout(w_dff_B_qNm5DonE1_2),.clk(gclk));
	jdff dff_B_SV2kvBoR0_2(.din(w_dff_B_qNm5DonE1_2),.dout(w_dff_B_SV2kvBoR0_2),.clk(gclk));
	jdff dff_B_EBIpuuQR8_2(.din(w_dff_B_SV2kvBoR0_2),.dout(w_dff_B_EBIpuuQR8_2),.clk(gclk));
	jdff dff_B_WeM40RcL6_2(.din(n1747),.dout(w_dff_B_WeM40RcL6_2),.clk(gclk));
	jdff dff_B_ntpkS7Lg8_1(.din(n1745),.dout(w_dff_B_ntpkS7Lg8_1),.clk(gclk));
	jdff dff_B_lG7B0dfC4_2(.din(n1709),.dout(w_dff_B_lG7B0dfC4_2),.clk(gclk));
	jdff dff_B_KJecEGLT1_2(.din(w_dff_B_lG7B0dfC4_2),.dout(w_dff_B_KJecEGLT1_2),.clk(gclk));
	jdff dff_B_5mxEd2ES5_2(.din(w_dff_B_KJecEGLT1_2),.dout(w_dff_B_5mxEd2ES5_2),.clk(gclk));
	jdff dff_B_p5mWZGv34_2(.din(w_dff_B_5mxEd2ES5_2),.dout(w_dff_B_p5mWZGv34_2),.clk(gclk));
	jdff dff_B_ojpNVx150_2(.din(w_dff_B_p5mWZGv34_2),.dout(w_dff_B_ojpNVx150_2),.clk(gclk));
	jdff dff_B_si9fCXoa2_2(.din(w_dff_B_ojpNVx150_2),.dout(w_dff_B_si9fCXoa2_2),.clk(gclk));
	jdff dff_B_OCgk9N5P9_2(.din(w_dff_B_si9fCXoa2_2),.dout(w_dff_B_OCgk9N5P9_2),.clk(gclk));
	jdff dff_B_WnmibGQH6_2(.din(w_dff_B_OCgk9N5P9_2),.dout(w_dff_B_WnmibGQH6_2),.clk(gclk));
	jdff dff_B_ph9dCYgJ7_2(.din(w_dff_B_WnmibGQH6_2),.dout(w_dff_B_ph9dCYgJ7_2),.clk(gclk));
	jdff dff_B_5VGsv4e43_2(.din(w_dff_B_ph9dCYgJ7_2),.dout(w_dff_B_5VGsv4e43_2),.clk(gclk));
	jdff dff_B_XZbLP5Lf1_2(.din(w_dff_B_5VGsv4e43_2),.dout(w_dff_B_XZbLP5Lf1_2),.clk(gclk));
	jdff dff_B_MNC0GTuQ2_2(.din(w_dff_B_XZbLP5Lf1_2),.dout(w_dff_B_MNC0GTuQ2_2),.clk(gclk));
	jdff dff_B_JbaTNY7h6_2(.din(w_dff_B_MNC0GTuQ2_2),.dout(w_dff_B_JbaTNY7h6_2),.clk(gclk));
	jdff dff_B_HQyyC0Ks2_2(.din(w_dff_B_JbaTNY7h6_2),.dout(w_dff_B_HQyyC0Ks2_2),.clk(gclk));
	jdff dff_B_vY6PerlF7_2(.din(w_dff_B_HQyyC0Ks2_2),.dout(w_dff_B_vY6PerlF7_2),.clk(gclk));
	jdff dff_B_1hAp9e208_2(.din(w_dff_B_vY6PerlF7_2),.dout(w_dff_B_1hAp9e208_2),.clk(gclk));
	jdff dff_B_XlhxLxdf4_2(.din(w_dff_B_1hAp9e208_2),.dout(w_dff_B_XlhxLxdf4_2),.clk(gclk));
	jdff dff_B_ya1aadhD8_2(.din(w_dff_B_XlhxLxdf4_2),.dout(w_dff_B_ya1aadhD8_2),.clk(gclk));
	jdff dff_B_6b2jPVpP9_2(.din(w_dff_B_ya1aadhD8_2),.dout(w_dff_B_6b2jPVpP9_2),.clk(gclk));
	jdff dff_B_ls1Z6PYf3_2(.din(w_dff_B_6b2jPVpP9_2),.dout(w_dff_B_ls1Z6PYf3_2),.clk(gclk));
	jdff dff_B_Q32PWZgJ5_2(.din(w_dff_B_ls1Z6PYf3_2),.dout(w_dff_B_Q32PWZgJ5_2),.clk(gclk));
	jdff dff_B_nOu8jI8L3_2(.din(w_dff_B_Q32PWZgJ5_2),.dout(w_dff_B_nOu8jI8L3_2),.clk(gclk));
	jdff dff_B_ThscDitp7_2(.din(w_dff_B_nOu8jI8L3_2),.dout(w_dff_B_ThscDitp7_2),.clk(gclk));
	jdff dff_B_RJkYcvaE6_2(.din(w_dff_B_ThscDitp7_2),.dout(w_dff_B_RJkYcvaE6_2),.clk(gclk));
	jdff dff_B_XxLkv4WB8_2(.din(w_dff_B_RJkYcvaE6_2),.dout(w_dff_B_XxLkv4WB8_2),.clk(gclk));
	jdff dff_B_4a0Znj3O4_2(.din(w_dff_B_XxLkv4WB8_2),.dout(w_dff_B_4a0Znj3O4_2),.clk(gclk));
	jdff dff_B_j9tULFLz3_2(.din(w_dff_B_4a0Znj3O4_2),.dout(w_dff_B_j9tULFLz3_2),.clk(gclk));
	jdff dff_B_n8hs05Cd5_2(.din(w_dff_B_j9tULFLz3_2),.dout(w_dff_B_n8hs05Cd5_2),.clk(gclk));
	jdff dff_B_LPoWhfUl3_2(.din(w_dff_B_n8hs05Cd5_2),.dout(w_dff_B_LPoWhfUl3_2),.clk(gclk));
	jdff dff_B_j1zwFrvm4_2(.din(w_dff_B_LPoWhfUl3_2),.dout(w_dff_B_j1zwFrvm4_2),.clk(gclk));
	jdff dff_B_xtrKM9KJ5_2(.din(w_dff_B_j1zwFrvm4_2),.dout(w_dff_B_xtrKM9KJ5_2),.clk(gclk));
	jdff dff_B_gStlqySk1_2(.din(w_dff_B_xtrKM9KJ5_2),.dout(w_dff_B_gStlqySk1_2),.clk(gclk));
	jdff dff_B_m1XEFau04_2(.din(w_dff_B_gStlqySk1_2),.dout(w_dff_B_m1XEFau04_2),.clk(gclk));
	jdff dff_B_rgFpqpQt5_2(.din(w_dff_B_m1XEFau04_2),.dout(w_dff_B_rgFpqpQt5_2),.clk(gclk));
	jdff dff_B_pJTzBIea4_2(.din(w_dff_B_rgFpqpQt5_2),.dout(w_dff_B_pJTzBIea4_2),.clk(gclk));
	jdff dff_B_VmGD0QdK1_2(.din(w_dff_B_pJTzBIea4_2),.dout(w_dff_B_VmGD0QdK1_2),.clk(gclk));
	jdff dff_B_tL8n37lo1_2(.din(w_dff_B_VmGD0QdK1_2),.dout(w_dff_B_tL8n37lo1_2),.clk(gclk));
	jdff dff_B_1EEhgPRe6_2(.din(w_dff_B_tL8n37lo1_2),.dout(w_dff_B_1EEhgPRe6_2),.clk(gclk));
	jdff dff_B_W2gLu4uP4_2(.din(w_dff_B_1EEhgPRe6_2),.dout(w_dff_B_W2gLu4uP4_2),.clk(gclk));
	jdff dff_B_zrvBGAS09_2(.din(w_dff_B_W2gLu4uP4_2),.dout(w_dff_B_zrvBGAS09_2),.clk(gclk));
	jdff dff_B_k9bITiLT4_2(.din(w_dff_B_zrvBGAS09_2),.dout(w_dff_B_k9bITiLT4_2),.clk(gclk));
	jdff dff_B_BamoOFI32_2(.din(w_dff_B_k9bITiLT4_2),.dout(w_dff_B_BamoOFI32_2),.clk(gclk));
	jdff dff_B_kY5qNx0X4_2(.din(w_dff_B_BamoOFI32_2),.dout(w_dff_B_kY5qNx0X4_2),.clk(gclk));
	jdff dff_B_hc8D6Meq7_2(.din(w_dff_B_kY5qNx0X4_2),.dout(w_dff_B_hc8D6Meq7_2),.clk(gclk));
	jdff dff_B_WENRyFSp3_1(.din(n1715),.dout(w_dff_B_WENRyFSp3_1),.clk(gclk));
	jdff dff_B_dofnAvnv2_1(.din(w_dff_B_WENRyFSp3_1),.dout(w_dff_B_dofnAvnv2_1),.clk(gclk));
	jdff dff_B_pSBUtnzf2_2(.din(n1714),.dout(w_dff_B_pSBUtnzf2_2),.clk(gclk));
	jdff dff_B_O3wxnIq12_2(.din(w_dff_B_pSBUtnzf2_2),.dout(w_dff_B_O3wxnIq12_2),.clk(gclk));
	jdff dff_B_14OyNwMz8_2(.din(w_dff_B_O3wxnIq12_2),.dout(w_dff_B_14OyNwMz8_2),.clk(gclk));
	jdff dff_B_R2UkBLZN6_2(.din(w_dff_B_14OyNwMz8_2),.dout(w_dff_B_R2UkBLZN6_2),.clk(gclk));
	jdff dff_B_Ir5t8v328_2(.din(w_dff_B_R2UkBLZN6_2),.dout(w_dff_B_Ir5t8v328_2),.clk(gclk));
	jdff dff_B_vvhWlZZ94_2(.din(w_dff_B_Ir5t8v328_2),.dout(w_dff_B_vvhWlZZ94_2),.clk(gclk));
	jdff dff_B_p3wJfSXo4_2(.din(w_dff_B_vvhWlZZ94_2),.dout(w_dff_B_p3wJfSXo4_2),.clk(gclk));
	jdff dff_B_FI3lRxcy8_2(.din(w_dff_B_p3wJfSXo4_2),.dout(w_dff_B_FI3lRxcy8_2),.clk(gclk));
	jdff dff_B_hUfJYE093_2(.din(w_dff_B_FI3lRxcy8_2),.dout(w_dff_B_hUfJYE093_2),.clk(gclk));
	jdff dff_B_GnXh7Pqn2_2(.din(w_dff_B_hUfJYE093_2),.dout(w_dff_B_GnXh7Pqn2_2),.clk(gclk));
	jdff dff_B_98zCHcyQ2_2(.din(w_dff_B_GnXh7Pqn2_2),.dout(w_dff_B_98zCHcyQ2_2),.clk(gclk));
	jdff dff_B_e1qiWSwR7_2(.din(w_dff_B_98zCHcyQ2_2),.dout(w_dff_B_e1qiWSwR7_2),.clk(gclk));
	jdff dff_B_SOnsn3GE9_2(.din(w_dff_B_e1qiWSwR7_2),.dout(w_dff_B_SOnsn3GE9_2),.clk(gclk));
	jdff dff_B_S6xX9IMr5_2(.din(w_dff_B_SOnsn3GE9_2),.dout(w_dff_B_S6xX9IMr5_2),.clk(gclk));
	jdff dff_B_U2PTNmWC1_2(.din(w_dff_B_S6xX9IMr5_2),.dout(w_dff_B_U2PTNmWC1_2),.clk(gclk));
	jdff dff_B_HhKI1uqI6_2(.din(w_dff_B_U2PTNmWC1_2),.dout(w_dff_B_HhKI1uqI6_2),.clk(gclk));
	jdff dff_B_AuJP7aRH3_2(.din(w_dff_B_HhKI1uqI6_2),.dout(w_dff_B_AuJP7aRH3_2),.clk(gclk));
	jdff dff_B_E4oFzWpb5_2(.din(w_dff_B_AuJP7aRH3_2),.dout(w_dff_B_E4oFzWpb5_2),.clk(gclk));
	jdff dff_B_hR4v2NY77_2(.din(w_dff_B_E4oFzWpb5_2),.dout(w_dff_B_hR4v2NY77_2),.clk(gclk));
	jdff dff_B_vFwUmgL80_2(.din(w_dff_B_hR4v2NY77_2),.dout(w_dff_B_vFwUmgL80_2),.clk(gclk));
	jdff dff_B_CUYVvrqS3_2(.din(w_dff_B_vFwUmgL80_2),.dout(w_dff_B_CUYVvrqS3_2),.clk(gclk));
	jdff dff_B_C5fZiopT0_2(.din(w_dff_B_CUYVvrqS3_2),.dout(w_dff_B_C5fZiopT0_2),.clk(gclk));
	jdff dff_B_QuAmi1I34_2(.din(w_dff_B_C5fZiopT0_2),.dout(w_dff_B_QuAmi1I34_2),.clk(gclk));
	jdff dff_B_vr3iXH2W2_2(.din(w_dff_B_QuAmi1I34_2),.dout(w_dff_B_vr3iXH2W2_2),.clk(gclk));
	jdff dff_B_HotQv0NS4_2(.din(w_dff_B_vr3iXH2W2_2),.dout(w_dff_B_HotQv0NS4_2),.clk(gclk));
	jdff dff_B_HCGhOKUu4_2(.din(w_dff_B_HotQv0NS4_2),.dout(w_dff_B_HCGhOKUu4_2),.clk(gclk));
	jdff dff_B_1MuYgIjq2_2(.din(w_dff_B_HCGhOKUu4_2),.dout(w_dff_B_1MuYgIjq2_2),.clk(gclk));
	jdff dff_B_MB9s2mwy8_2(.din(w_dff_B_1MuYgIjq2_2),.dout(w_dff_B_MB9s2mwy8_2),.clk(gclk));
	jdff dff_B_g3DZWlK20_2(.din(w_dff_B_MB9s2mwy8_2),.dout(w_dff_B_g3DZWlK20_2),.clk(gclk));
	jdff dff_B_Q1XIJ01N1_2(.din(w_dff_B_g3DZWlK20_2),.dout(w_dff_B_Q1XIJ01N1_2),.clk(gclk));
	jdff dff_B_pl1VKKq94_2(.din(w_dff_B_Q1XIJ01N1_2),.dout(w_dff_B_pl1VKKq94_2),.clk(gclk));
	jdff dff_B_6M08i3Rs0_2(.din(w_dff_B_pl1VKKq94_2),.dout(w_dff_B_6M08i3Rs0_2),.clk(gclk));
	jdff dff_B_ueYOJYnk6_2(.din(w_dff_B_6M08i3Rs0_2),.dout(w_dff_B_ueYOJYnk6_2),.clk(gclk));
	jdff dff_B_RMmkhvFz7_2(.din(w_dff_B_ueYOJYnk6_2),.dout(w_dff_B_RMmkhvFz7_2),.clk(gclk));
	jdff dff_B_m1BpQfr49_2(.din(w_dff_B_RMmkhvFz7_2),.dout(w_dff_B_m1BpQfr49_2),.clk(gclk));
	jdff dff_B_ScpP36Ta3_2(.din(w_dff_B_m1BpQfr49_2),.dout(w_dff_B_ScpP36Ta3_2),.clk(gclk));
	jdff dff_B_y7uob3vh7_2(.din(w_dff_B_ScpP36Ta3_2),.dout(w_dff_B_y7uob3vh7_2),.clk(gclk));
	jdff dff_B_cSZHN7Iz6_2(.din(w_dff_B_y7uob3vh7_2),.dout(w_dff_B_cSZHN7Iz6_2),.clk(gclk));
	jdff dff_B_T0aF33hJ2_2(.din(w_dff_B_cSZHN7Iz6_2),.dout(w_dff_B_T0aF33hJ2_2),.clk(gclk));
	jdff dff_B_8V6d5mBP2_2(.din(w_dff_B_T0aF33hJ2_2),.dout(w_dff_B_8V6d5mBP2_2),.clk(gclk));
	jdff dff_B_qvorlkVc9_2(.din(w_dff_B_8V6d5mBP2_2),.dout(w_dff_B_qvorlkVc9_2),.clk(gclk));
	jdff dff_B_ORVskRRL0_2(.din(n1713),.dout(w_dff_B_ORVskRRL0_2),.clk(gclk));
	jdff dff_B_uFLbA16n0_2(.din(w_dff_B_ORVskRRL0_2),.dout(w_dff_B_uFLbA16n0_2),.clk(gclk));
	jdff dff_B_hPPU42YS7_2(.din(w_dff_B_uFLbA16n0_2),.dout(w_dff_B_hPPU42YS7_2),.clk(gclk));
	jdff dff_B_zSHorKoy5_2(.din(w_dff_B_hPPU42YS7_2),.dout(w_dff_B_zSHorKoy5_2),.clk(gclk));
	jdff dff_B_Dsq5ntar3_2(.din(w_dff_B_zSHorKoy5_2),.dout(w_dff_B_Dsq5ntar3_2),.clk(gclk));
	jdff dff_B_hkowsfGn2_2(.din(w_dff_B_Dsq5ntar3_2),.dout(w_dff_B_hkowsfGn2_2),.clk(gclk));
	jdff dff_B_zzUlKvej9_2(.din(w_dff_B_hkowsfGn2_2),.dout(w_dff_B_zzUlKvej9_2),.clk(gclk));
	jdff dff_B_nlG2aPkr8_2(.din(w_dff_B_zzUlKvej9_2),.dout(w_dff_B_nlG2aPkr8_2),.clk(gclk));
	jdff dff_B_hpD5bY4P9_2(.din(w_dff_B_nlG2aPkr8_2),.dout(w_dff_B_hpD5bY4P9_2),.clk(gclk));
	jdff dff_B_lwvS4Zqz8_2(.din(w_dff_B_hpD5bY4P9_2),.dout(w_dff_B_lwvS4Zqz8_2),.clk(gclk));
	jdff dff_B_h47sk5SR6_2(.din(w_dff_B_lwvS4Zqz8_2),.dout(w_dff_B_h47sk5SR6_2),.clk(gclk));
	jdff dff_B_z07UA75T7_2(.din(w_dff_B_h47sk5SR6_2),.dout(w_dff_B_z07UA75T7_2),.clk(gclk));
	jdff dff_B_hoiRqGj51_2(.din(w_dff_B_z07UA75T7_2),.dout(w_dff_B_hoiRqGj51_2),.clk(gclk));
	jdff dff_B_BU8PtD0b4_2(.din(w_dff_B_hoiRqGj51_2),.dout(w_dff_B_BU8PtD0b4_2),.clk(gclk));
	jdff dff_B_ruquY5fG5_2(.din(w_dff_B_BU8PtD0b4_2),.dout(w_dff_B_ruquY5fG5_2),.clk(gclk));
	jdff dff_B_ZoTcBwNy0_2(.din(w_dff_B_ruquY5fG5_2),.dout(w_dff_B_ZoTcBwNy0_2),.clk(gclk));
	jdff dff_B_zHr4kXGj1_2(.din(w_dff_B_ZoTcBwNy0_2),.dout(w_dff_B_zHr4kXGj1_2),.clk(gclk));
	jdff dff_B_ACzXzg0L4_2(.din(w_dff_B_zHr4kXGj1_2),.dout(w_dff_B_ACzXzg0L4_2),.clk(gclk));
	jdff dff_B_rP9G3l960_2(.din(w_dff_B_ACzXzg0L4_2),.dout(w_dff_B_rP9G3l960_2),.clk(gclk));
	jdff dff_B_Rp6DzqGG0_2(.din(w_dff_B_rP9G3l960_2),.dout(w_dff_B_Rp6DzqGG0_2),.clk(gclk));
	jdff dff_B_GBP0cfjm9_2(.din(w_dff_B_Rp6DzqGG0_2),.dout(w_dff_B_GBP0cfjm9_2),.clk(gclk));
	jdff dff_B_MVtfaO6K0_2(.din(w_dff_B_GBP0cfjm9_2),.dout(w_dff_B_MVtfaO6K0_2),.clk(gclk));
	jdff dff_B_QXqo12Wh5_2(.din(w_dff_B_MVtfaO6K0_2),.dout(w_dff_B_QXqo12Wh5_2),.clk(gclk));
	jdff dff_B_X11AiJN49_2(.din(w_dff_B_QXqo12Wh5_2),.dout(w_dff_B_X11AiJN49_2),.clk(gclk));
	jdff dff_B_rSkWizs21_2(.din(w_dff_B_X11AiJN49_2),.dout(w_dff_B_rSkWizs21_2),.clk(gclk));
	jdff dff_B_GbEMdghI6_2(.din(w_dff_B_rSkWizs21_2),.dout(w_dff_B_GbEMdghI6_2),.clk(gclk));
	jdff dff_B_CghXusbL2_2(.din(w_dff_B_GbEMdghI6_2),.dout(w_dff_B_CghXusbL2_2),.clk(gclk));
	jdff dff_B_AHRYWI4h6_2(.din(w_dff_B_CghXusbL2_2),.dout(w_dff_B_AHRYWI4h6_2),.clk(gclk));
	jdff dff_B_b10RUB805_2(.din(w_dff_B_AHRYWI4h6_2),.dout(w_dff_B_b10RUB805_2),.clk(gclk));
	jdff dff_B_E0DuHRWX5_2(.din(w_dff_B_b10RUB805_2),.dout(w_dff_B_E0DuHRWX5_2),.clk(gclk));
	jdff dff_B_DQki4TfN8_2(.din(w_dff_B_E0DuHRWX5_2),.dout(w_dff_B_DQki4TfN8_2),.clk(gclk));
	jdff dff_B_BJxRN4Rq8_2(.din(w_dff_B_DQki4TfN8_2),.dout(w_dff_B_BJxRN4Rq8_2),.clk(gclk));
	jdff dff_B_gUA60vJn9_2(.din(w_dff_B_BJxRN4Rq8_2),.dout(w_dff_B_gUA60vJn9_2),.clk(gclk));
	jdff dff_B_NKbBbhAo5_2(.din(w_dff_B_gUA60vJn9_2),.dout(w_dff_B_NKbBbhAo5_2),.clk(gclk));
	jdff dff_B_OY1yIeMD6_2(.din(w_dff_B_NKbBbhAo5_2),.dout(w_dff_B_OY1yIeMD6_2),.clk(gclk));
	jdff dff_B_1AsiLKXu0_2(.din(w_dff_B_OY1yIeMD6_2),.dout(w_dff_B_1AsiLKXu0_2),.clk(gclk));
	jdff dff_B_YOk2K5Xj7_2(.din(w_dff_B_1AsiLKXu0_2),.dout(w_dff_B_YOk2K5Xj7_2),.clk(gclk));
	jdff dff_B_5QgVmLnI6_2(.din(w_dff_B_YOk2K5Xj7_2),.dout(w_dff_B_5QgVmLnI6_2),.clk(gclk));
	jdff dff_B_6Qk5svwe4_2(.din(w_dff_B_5QgVmLnI6_2),.dout(w_dff_B_6Qk5svwe4_2),.clk(gclk));
	jdff dff_B_V6ItlT3I2_2(.din(w_dff_B_6Qk5svwe4_2),.dout(w_dff_B_V6ItlT3I2_2),.clk(gclk));
	jdff dff_B_82aBdxM65_2(.din(w_dff_B_V6ItlT3I2_2),.dout(w_dff_B_82aBdxM65_2),.clk(gclk));
	jdff dff_B_GZT2zF813_2(.din(w_dff_B_82aBdxM65_2),.dout(w_dff_B_GZT2zF813_2),.clk(gclk));
	jdff dff_B_Iwu0JBoY1_2(.din(w_dff_B_GZT2zF813_2),.dout(w_dff_B_Iwu0JBoY1_2),.clk(gclk));
	jdff dff_B_fSAmthdF5_2(.din(n1712),.dout(w_dff_B_fSAmthdF5_2),.clk(gclk));
	jdff dff_B_so3bvXCA9_1(.din(n1710),.dout(w_dff_B_so3bvXCA9_1),.clk(gclk));
	jdff dff_B_vtEi4Kpz3_2(.din(n1668),.dout(w_dff_B_vtEi4Kpz3_2),.clk(gclk));
	jdff dff_B_rMh5kDWf4_2(.din(w_dff_B_vtEi4Kpz3_2),.dout(w_dff_B_rMh5kDWf4_2),.clk(gclk));
	jdff dff_B_W3huiePw8_2(.din(w_dff_B_rMh5kDWf4_2),.dout(w_dff_B_W3huiePw8_2),.clk(gclk));
	jdff dff_B_GmeMhhA71_2(.din(w_dff_B_W3huiePw8_2),.dout(w_dff_B_GmeMhhA71_2),.clk(gclk));
	jdff dff_B_C7QERlP91_2(.din(w_dff_B_GmeMhhA71_2),.dout(w_dff_B_C7QERlP91_2),.clk(gclk));
	jdff dff_B_84s5c5Nz2_2(.din(w_dff_B_C7QERlP91_2),.dout(w_dff_B_84s5c5Nz2_2),.clk(gclk));
	jdff dff_B_7ZW0x3g02_2(.din(w_dff_B_84s5c5Nz2_2),.dout(w_dff_B_7ZW0x3g02_2),.clk(gclk));
	jdff dff_B_aPDhGeFP9_2(.din(w_dff_B_7ZW0x3g02_2),.dout(w_dff_B_aPDhGeFP9_2),.clk(gclk));
	jdff dff_B_KaUutlwy9_2(.din(w_dff_B_aPDhGeFP9_2),.dout(w_dff_B_KaUutlwy9_2),.clk(gclk));
	jdff dff_B_bySvzJn36_2(.din(w_dff_B_KaUutlwy9_2),.dout(w_dff_B_bySvzJn36_2),.clk(gclk));
	jdff dff_B_O66wpek53_2(.din(w_dff_B_bySvzJn36_2),.dout(w_dff_B_O66wpek53_2),.clk(gclk));
	jdff dff_B_aizqsT1X0_2(.din(w_dff_B_O66wpek53_2),.dout(w_dff_B_aizqsT1X0_2),.clk(gclk));
	jdff dff_B_aiutfzTc1_2(.din(w_dff_B_aizqsT1X0_2),.dout(w_dff_B_aiutfzTc1_2),.clk(gclk));
	jdff dff_B_12oASWHn1_2(.din(w_dff_B_aiutfzTc1_2),.dout(w_dff_B_12oASWHn1_2),.clk(gclk));
	jdff dff_B_alXqnom34_2(.din(w_dff_B_12oASWHn1_2),.dout(w_dff_B_alXqnom34_2),.clk(gclk));
	jdff dff_B_ONerYRmf7_2(.din(w_dff_B_alXqnom34_2),.dout(w_dff_B_ONerYRmf7_2),.clk(gclk));
	jdff dff_B_Rrpl6yNC2_2(.din(w_dff_B_ONerYRmf7_2),.dout(w_dff_B_Rrpl6yNC2_2),.clk(gclk));
	jdff dff_B_ix0Gi1mB1_2(.din(w_dff_B_Rrpl6yNC2_2),.dout(w_dff_B_ix0Gi1mB1_2),.clk(gclk));
	jdff dff_B_zNqUTJr67_2(.din(w_dff_B_ix0Gi1mB1_2),.dout(w_dff_B_zNqUTJr67_2),.clk(gclk));
	jdff dff_B_EmUI2uyv6_2(.din(w_dff_B_zNqUTJr67_2),.dout(w_dff_B_EmUI2uyv6_2),.clk(gclk));
	jdff dff_B_x5jrItde3_2(.din(w_dff_B_EmUI2uyv6_2),.dout(w_dff_B_x5jrItde3_2),.clk(gclk));
	jdff dff_B_PvovAB4y7_2(.din(w_dff_B_x5jrItde3_2),.dout(w_dff_B_PvovAB4y7_2),.clk(gclk));
	jdff dff_B_Bh9Ch4t81_2(.din(w_dff_B_PvovAB4y7_2),.dout(w_dff_B_Bh9Ch4t81_2),.clk(gclk));
	jdff dff_B_i92uPmxT6_2(.din(w_dff_B_Bh9Ch4t81_2),.dout(w_dff_B_i92uPmxT6_2),.clk(gclk));
	jdff dff_B_raTTTJJC9_2(.din(w_dff_B_i92uPmxT6_2),.dout(w_dff_B_raTTTJJC9_2),.clk(gclk));
	jdff dff_B_niThLe7M3_2(.din(w_dff_B_raTTTJJC9_2),.dout(w_dff_B_niThLe7M3_2),.clk(gclk));
	jdff dff_B_JuaK0qrj5_2(.din(w_dff_B_niThLe7M3_2),.dout(w_dff_B_JuaK0qrj5_2),.clk(gclk));
	jdff dff_B_NBcwkllt8_2(.din(w_dff_B_JuaK0qrj5_2),.dout(w_dff_B_NBcwkllt8_2),.clk(gclk));
	jdff dff_B_aYlYT9TL0_2(.din(w_dff_B_NBcwkllt8_2),.dout(w_dff_B_aYlYT9TL0_2),.clk(gclk));
	jdff dff_B_0rHLpv2Q3_2(.din(w_dff_B_aYlYT9TL0_2),.dout(w_dff_B_0rHLpv2Q3_2),.clk(gclk));
	jdff dff_B_aspizn5w9_2(.din(w_dff_B_0rHLpv2Q3_2),.dout(w_dff_B_aspizn5w9_2),.clk(gclk));
	jdff dff_B_Lh31jnUz8_2(.din(w_dff_B_aspizn5w9_2),.dout(w_dff_B_Lh31jnUz8_2),.clk(gclk));
	jdff dff_B_tQKoUhBA2_2(.din(w_dff_B_Lh31jnUz8_2),.dout(w_dff_B_tQKoUhBA2_2),.clk(gclk));
	jdff dff_B_BaVR6MCD1_2(.din(w_dff_B_tQKoUhBA2_2),.dout(w_dff_B_BaVR6MCD1_2),.clk(gclk));
	jdff dff_B_Eq2yXbdA5_2(.din(w_dff_B_BaVR6MCD1_2),.dout(w_dff_B_Eq2yXbdA5_2),.clk(gclk));
	jdff dff_B_EW9AYF2q3_2(.din(w_dff_B_Eq2yXbdA5_2),.dout(w_dff_B_EW9AYF2q3_2),.clk(gclk));
	jdff dff_B_rjDBiP412_2(.din(w_dff_B_EW9AYF2q3_2),.dout(w_dff_B_rjDBiP412_2),.clk(gclk));
	jdff dff_B_VlbZDsvX9_2(.din(w_dff_B_rjDBiP412_2),.dout(w_dff_B_VlbZDsvX9_2),.clk(gclk));
	jdff dff_B_EZofrVWs8_2(.din(w_dff_B_VlbZDsvX9_2),.dout(w_dff_B_EZofrVWs8_2),.clk(gclk));
	jdff dff_B_YSlYmL2F6_2(.din(w_dff_B_EZofrVWs8_2),.dout(w_dff_B_YSlYmL2F6_2),.clk(gclk));
	jdff dff_B_Jfqm8b2C2_1(.din(n1674),.dout(w_dff_B_Jfqm8b2C2_1),.clk(gclk));
	jdff dff_B_XGro1DDU8_1(.din(w_dff_B_Jfqm8b2C2_1),.dout(w_dff_B_XGro1DDU8_1),.clk(gclk));
	jdff dff_B_DCt7W3KY5_2(.din(n1673),.dout(w_dff_B_DCt7W3KY5_2),.clk(gclk));
	jdff dff_B_Ze1Gbbtc4_2(.din(w_dff_B_DCt7W3KY5_2),.dout(w_dff_B_Ze1Gbbtc4_2),.clk(gclk));
	jdff dff_B_afN3qDdr6_2(.din(w_dff_B_Ze1Gbbtc4_2),.dout(w_dff_B_afN3qDdr6_2),.clk(gclk));
	jdff dff_B_zNipOtPz0_2(.din(w_dff_B_afN3qDdr6_2),.dout(w_dff_B_zNipOtPz0_2),.clk(gclk));
	jdff dff_B_T48beAEl9_2(.din(w_dff_B_zNipOtPz0_2),.dout(w_dff_B_T48beAEl9_2),.clk(gclk));
	jdff dff_B_zanLY2pj5_2(.din(w_dff_B_T48beAEl9_2),.dout(w_dff_B_zanLY2pj5_2),.clk(gclk));
	jdff dff_B_o3WkWxfY1_2(.din(w_dff_B_zanLY2pj5_2),.dout(w_dff_B_o3WkWxfY1_2),.clk(gclk));
	jdff dff_B_4ODzqni49_2(.din(w_dff_B_o3WkWxfY1_2),.dout(w_dff_B_4ODzqni49_2),.clk(gclk));
	jdff dff_B_Nd0ab4CN2_2(.din(w_dff_B_4ODzqni49_2),.dout(w_dff_B_Nd0ab4CN2_2),.clk(gclk));
	jdff dff_B_ZQLpiDU95_2(.din(w_dff_B_Nd0ab4CN2_2),.dout(w_dff_B_ZQLpiDU95_2),.clk(gclk));
	jdff dff_B_mGISbn4m9_2(.din(w_dff_B_ZQLpiDU95_2),.dout(w_dff_B_mGISbn4m9_2),.clk(gclk));
	jdff dff_B_lSaa4y9E0_2(.din(w_dff_B_mGISbn4m9_2),.dout(w_dff_B_lSaa4y9E0_2),.clk(gclk));
	jdff dff_B_bMaQ7bwB8_2(.din(w_dff_B_lSaa4y9E0_2),.dout(w_dff_B_bMaQ7bwB8_2),.clk(gclk));
	jdff dff_B_V7dQB2OC2_2(.din(w_dff_B_bMaQ7bwB8_2),.dout(w_dff_B_V7dQB2OC2_2),.clk(gclk));
	jdff dff_B_cyHswZPc6_2(.din(w_dff_B_V7dQB2OC2_2),.dout(w_dff_B_cyHswZPc6_2),.clk(gclk));
	jdff dff_B_24iqTy5j5_2(.din(w_dff_B_cyHswZPc6_2),.dout(w_dff_B_24iqTy5j5_2),.clk(gclk));
	jdff dff_B_8xclsG7e0_2(.din(w_dff_B_24iqTy5j5_2),.dout(w_dff_B_8xclsG7e0_2),.clk(gclk));
	jdff dff_B_wOx0yO1d7_2(.din(w_dff_B_8xclsG7e0_2),.dout(w_dff_B_wOx0yO1d7_2),.clk(gclk));
	jdff dff_B_HnLvbag86_2(.din(w_dff_B_wOx0yO1d7_2),.dout(w_dff_B_HnLvbag86_2),.clk(gclk));
	jdff dff_B_1dpNgc582_2(.din(w_dff_B_HnLvbag86_2),.dout(w_dff_B_1dpNgc582_2),.clk(gclk));
	jdff dff_B_inlD8xDw3_2(.din(w_dff_B_1dpNgc582_2),.dout(w_dff_B_inlD8xDw3_2),.clk(gclk));
	jdff dff_B_rpjd2GH41_2(.din(w_dff_B_inlD8xDw3_2),.dout(w_dff_B_rpjd2GH41_2),.clk(gclk));
	jdff dff_B_DjxsCOey1_2(.din(w_dff_B_rpjd2GH41_2),.dout(w_dff_B_DjxsCOey1_2),.clk(gclk));
	jdff dff_B_EF4Ictk27_2(.din(w_dff_B_DjxsCOey1_2),.dout(w_dff_B_EF4Ictk27_2),.clk(gclk));
	jdff dff_B_Mbcn8u8I1_2(.din(w_dff_B_EF4Ictk27_2),.dout(w_dff_B_Mbcn8u8I1_2),.clk(gclk));
	jdff dff_B_KZy9Wzyl2_2(.din(w_dff_B_Mbcn8u8I1_2),.dout(w_dff_B_KZy9Wzyl2_2),.clk(gclk));
	jdff dff_B_oTyIkkL54_2(.din(w_dff_B_KZy9Wzyl2_2),.dout(w_dff_B_oTyIkkL54_2),.clk(gclk));
	jdff dff_B_2Eqq8dfa6_2(.din(w_dff_B_oTyIkkL54_2),.dout(w_dff_B_2Eqq8dfa6_2),.clk(gclk));
	jdff dff_B_RplELcYv5_2(.din(w_dff_B_2Eqq8dfa6_2),.dout(w_dff_B_RplELcYv5_2),.clk(gclk));
	jdff dff_B_Mpd7KjoO9_2(.din(w_dff_B_RplELcYv5_2),.dout(w_dff_B_Mpd7KjoO9_2),.clk(gclk));
	jdff dff_B_6ZIO1vSb3_2(.din(w_dff_B_Mpd7KjoO9_2),.dout(w_dff_B_6ZIO1vSb3_2),.clk(gclk));
	jdff dff_B_r1Iwv30N4_2(.din(w_dff_B_6ZIO1vSb3_2),.dout(w_dff_B_r1Iwv30N4_2),.clk(gclk));
	jdff dff_B_7LBpGpU68_2(.din(w_dff_B_r1Iwv30N4_2),.dout(w_dff_B_7LBpGpU68_2),.clk(gclk));
	jdff dff_B_jrTO1hzs4_2(.din(w_dff_B_7LBpGpU68_2),.dout(w_dff_B_jrTO1hzs4_2),.clk(gclk));
	jdff dff_B_0dPZOt1m0_2(.din(w_dff_B_jrTO1hzs4_2),.dout(w_dff_B_0dPZOt1m0_2),.clk(gclk));
	jdff dff_B_Xqy7mTJH3_2(.din(w_dff_B_0dPZOt1m0_2),.dout(w_dff_B_Xqy7mTJH3_2),.clk(gclk));
	jdff dff_B_nLDF5s0E1_2(.din(w_dff_B_Xqy7mTJH3_2),.dout(w_dff_B_nLDF5s0E1_2),.clk(gclk));
	jdff dff_B_Gn5z5N8B7_2(.din(n1672),.dout(w_dff_B_Gn5z5N8B7_2),.clk(gclk));
	jdff dff_B_oxrMN8Kh5_2(.din(w_dff_B_Gn5z5N8B7_2),.dout(w_dff_B_oxrMN8Kh5_2),.clk(gclk));
	jdff dff_B_4Na5e2Ve2_2(.din(w_dff_B_oxrMN8Kh5_2),.dout(w_dff_B_4Na5e2Ve2_2),.clk(gclk));
	jdff dff_B_mqT7sGcI9_2(.din(w_dff_B_4Na5e2Ve2_2),.dout(w_dff_B_mqT7sGcI9_2),.clk(gclk));
	jdff dff_B_I0wq4VfE7_2(.din(w_dff_B_mqT7sGcI9_2),.dout(w_dff_B_I0wq4VfE7_2),.clk(gclk));
	jdff dff_B_4p7ifI9w6_2(.din(w_dff_B_I0wq4VfE7_2),.dout(w_dff_B_4p7ifI9w6_2),.clk(gclk));
	jdff dff_B_8KitNCqB3_2(.din(w_dff_B_4p7ifI9w6_2),.dout(w_dff_B_8KitNCqB3_2),.clk(gclk));
	jdff dff_B_E8h5qvUD1_2(.din(w_dff_B_8KitNCqB3_2),.dout(w_dff_B_E8h5qvUD1_2),.clk(gclk));
	jdff dff_B_wDljcrXF6_2(.din(w_dff_B_E8h5qvUD1_2),.dout(w_dff_B_wDljcrXF6_2),.clk(gclk));
	jdff dff_B_FGQZMneQ8_2(.din(w_dff_B_wDljcrXF6_2),.dout(w_dff_B_FGQZMneQ8_2),.clk(gclk));
	jdff dff_B_S4IAZWVB1_2(.din(w_dff_B_FGQZMneQ8_2),.dout(w_dff_B_S4IAZWVB1_2),.clk(gclk));
	jdff dff_B_2Kh34KYl0_2(.din(w_dff_B_S4IAZWVB1_2),.dout(w_dff_B_2Kh34KYl0_2),.clk(gclk));
	jdff dff_B_ZPGuMP478_2(.din(w_dff_B_2Kh34KYl0_2),.dout(w_dff_B_ZPGuMP478_2),.clk(gclk));
	jdff dff_B_xxvAtJO13_2(.din(w_dff_B_ZPGuMP478_2),.dout(w_dff_B_xxvAtJO13_2),.clk(gclk));
	jdff dff_B_w8vxuQ7V0_2(.din(w_dff_B_xxvAtJO13_2),.dout(w_dff_B_w8vxuQ7V0_2),.clk(gclk));
	jdff dff_B_IG7nORry1_2(.din(w_dff_B_w8vxuQ7V0_2),.dout(w_dff_B_IG7nORry1_2),.clk(gclk));
	jdff dff_B_PSJ3wbRG5_2(.din(w_dff_B_IG7nORry1_2),.dout(w_dff_B_PSJ3wbRG5_2),.clk(gclk));
	jdff dff_B_IwR4VEJz9_2(.din(w_dff_B_PSJ3wbRG5_2),.dout(w_dff_B_IwR4VEJz9_2),.clk(gclk));
	jdff dff_B_0AN5FYnj7_2(.din(w_dff_B_IwR4VEJz9_2),.dout(w_dff_B_0AN5FYnj7_2),.clk(gclk));
	jdff dff_B_rUYiWd898_2(.din(w_dff_B_0AN5FYnj7_2),.dout(w_dff_B_rUYiWd898_2),.clk(gclk));
	jdff dff_B_YAml3ti30_2(.din(w_dff_B_rUYiWd898_2),.dout(w_dff_B_YAml3ti30_2),.clk(gclk));
	jdff dff_B_KXMdH0Dv1_2(.din(w_dff_B_YAml3ti30_2),.dout(w_dff_B_KXMdH0Dv1_2),.clk(gclk));
	jdff dff_B_GoOFHact8_2(.din(w_dff_B_KXMdH0Dv1_2),.dout(w_dff_B_GoOFHact8_2),.clk(gclk));
	jdff dff_B_y1NWIWDG0_2(.din(w_dff_B_GoOFHact8_2),.dout(w_dff_B_y1NWIWDG0_2),.clk(gclk));
	jdff dff_B_2PNBIXAu4_2(.din(w_dff_B_y1NWIWDG0_2),.dout(w_dff_B_2PNBIXAu4_2),.clk(gclk));
	jdff dff_B_rqmfBGFq8_2(.din(w_dff_B_2PNBIXAu4_2),.dout(w_dff_B_rqmfBGFq8_2),.clk(gclk));
	jdff dff_B_LlQ4oQ0Q5_2(.din(w_dff_B_rqmfBGFq8_2),.dout(w_dff_B_LlQ4oQ0Q5_2),.clk(gclk));
	jdff dff_B_zXddmIFX4_2(.din(w_dff_B_LlQ4oQ0Q5_2),.dout(w_dff_B_zXddmIFX4_2),.clk(gclk));
	jdff dff_B_VMphltbY0_2(.din(w_dff_B_zXddmIFX4_2),.dout(w_dff_B_VMphltbY0_2),.clk(gclk));
	jdff dff_B_mcgQLaqK0_2(.din(w_dff_B_VMphltbY0_2),.dout(w_dff_B_mcgQLaqK0_2),.clk(gclk));
	jdff dff_B_islzgUuV1_2(.din(w_dff_B_mcgQLaqK0_2),.dout(w_dff_B_islzgUuV1_2),.clk(gclk));
	jdff dff_B_HzXEvtSl7_2(.din(w_dff_B_islzgUuV1_2),.dout(w_dff_B_HzXEvtSl7_2),.clk(gclk));
	jdff dff_B_90Nz1PCK0_2(.din(w_dff_B_HzXEvtSl7_2),.dout(w_dff_B_90Nz1PCK0_2),.clk(gclk));
	jdff dff_B_QcZsuWx58_2(.din(w_dff_B_90Nz1PCK0_2),.dout(w_dff_B_QcZsuWx58_2),.clk(gclk));
	jdff dff_B_qpxyykvy9_2(.din(w_dff_B_QcZsuWx58_2),.dout(w_dff_B_qpxyykvy9_2),.clk(gclk));
	jdff dff_B_tjsDtm5i5_2(.din(w_dff_B_qpxyykvy9_2),.dout(w_dff_B_tjsDtm5i5_2),.clk(gclk));
	jdff dff_B_PwJXIweD9_2(.din(w_dff_B_tjsDtm5i5_2),.dout(w_dff_B_PwJXIweD9_2),.clk(gclk));
	jdff dff_B_f2N7aWOk5_2(.din(w_dff_B_PwJXIweD9_2),.dout(w_dff_B_f2N7aWOk5_2),.clk(gclk));
	jdff dff_B_SKoI0v3m4_2(.din(w_dff_B_f2N7aWOk5_2),.dout(w_dff_B_SKoI0v3m4_2),.clk(gclk));
	jdff dff_B_GhTEZuUV2_2(.din(n1671),.dout(w_dff_B_GhTEZuUV2_2),.clk(gclk));
	jdff dff_B_egK88UFU6_1(.din(n1669),.dout(w_dff_B_egK88UFU6_1),.clk(gclk));
	jdff dff_B_nuPRXyN19_2(.din(n1617),.dout(w_dff_B_nuPRXyN19_2),.clk(gclk));
	jdff dff_B_OV3k2TzR9_2(.din(w_dff_B_nuPRXyN19_2),.dout(w_dff_B_OV3k2TzR9_2),.clk(gclk));
	jdff dff_B_AkPfrcEy4_2(.din(w_dff_B_OV3k2TzR9_2),.dout(w_dff_B_AkPfrcEy4_2),.clk(gclk));
	jdff dff_B_B9JU5BK58_2(.din(w_dff_B_AkPfrcEy4_2),.dout(w_dff_B_B9JU5BK58_2),.clk(gclk));
	jdff dff_B_95thr4gk8_2(.din(w_dff_B_B9JU5BK58_2),.dout(w_dff_B_95thr4gk8_2),.clk(gclk));
	jdff dff_B_3Qn4gqZ09_2(.din(w_dff_B_95thr4gk8_2),.dout(w_dff_B_3Qn4gqZ09_2),.clk(gclk));
	jdff dff_B_5GvkDcz38_2(.din(w_dff_B_3Qn4gqZ09_2),.dout(w_dff_B_5GvkDcz38_2),.clk(gclk));
	jdff dff_B_EPcGO0WF1_2(.din(w_dff_B_5GvkDcz38_2),.dout(w_dff_B_EPcGO0WF1_2),.clk(gclk));
	jdff dff_B_bnL5c9sb2_2(.din(w_dff_B_EPcGO0WF1_2),.dout(w_dff_B_bnL5c9sb2_2),.clk(gclk));
	jdff dff_B_T8XW9peQ7_2(.din(w_dff_B_bnL5c9sb2_2),.dout(w_dff_B_T8XW9peQ7_2),.clk(gclk));
	jdff dff_B_9Yad3EFy0_2(.din(w_dff_B_T8XW9peQ7_2),.dout(w_dff_B_9Yad3EFy0_2),.clk(gclk));
	jdff dff_B_zn8z2mBb6_2(.din(w_dff_B_9Yad3EFy0_2),.dout(w_dff_B_zn8z2mBb6_2),.clk(gclk));
	jdff dff_B_h4DXpltR5_2(.din(w_dff_B_zn8z2mBb6_2),.dout(w_dff_B_h4DXpltR5_2),.clk(gclk));
	jdff dff_B_lKBVVANg4_2(.din(w_dff_B_h4DXpltR5_2),.dout(w_dff_B_lKBVVANg4_2),.clk(gclk));
	jdff dff_B_ENot0orb1_2(.din(w_dff_B_lKBVVANg4_2),.dout(w_dff_B_ENot0orb1_2),.clk(gclk));
	jdff dff_B_D09HICv27_2(.din(w_dff_B_ENot0orb1_2),.dout(w_dff_B_D09HICv27_2),.clk(gclk));
	jdff dff_B_OAfFfalN6_2(.din(w_dff_B_D09HICv27_2),.dout(w_dff_B_OAfFfalN6_2),.clk(gclk));
	jdff dff_B_nMq9dOsC3_2(.din(w_dff_B_OAfFfalN6_2),.dout(w_dff_B_nMq9dOsC3_2),.clk(gclk));
	jdff dff_B_K0ZaFbJq8_2(.din(w_dff_B_nMq9dOsC3_2),.dout(w_dff_B_K0ZaFbJq8_2),.clk(gclk));
	jdff dff_B_uvcL2WJG4_2(.din(w_dff_B_K0ZaFbJq8_2),.dout(w_dff_B_uvcL2WJG4_2),.clk(gclk));
	jdff dff_B_CZZznmh27_2(.din(w_dff_B_uvcL2WJG4_2),.dout(w_dff_B_CZZznmh27_2),.clk(gclk));
	jdff dff_B_OhNPlfJw6_2(.din(w_dff_B_CZZznmh27_2),.dout(w_dff_B_OhNPlfJw6_2),.clk(gclk));
	jdff dff_B_kW2INgSM3_2(.din(w_dff_B_OhNPlfJw6_2),.dout(w_dff_B_kW2INgSM3_2),.clk(gclk));
	jdff dff_B_9bj1JdwC4_2(.din(w_dff_B_kW2INgSM3_2),.dout(w_dff_B_9bj1JdwC4_2),.clk(gclk));
	jdff dff_B_KpoYko7H8_2(.din(w_dff_B_9bj1JdwC4_2),.dout(w_dff_B_KpoYko7H8_2),.clk(gclk));
	jdff dff_B_x6RjqWcj0_2(.din(w_dff_B_KpoYko7H8_2),.dout(w_dff_B_x6RjqWcj0_2),.clk(gclk));
	jdff dff_B_HKZYHUZX9_2(.din(w_dff_B_x6RjqWcj0_2),.dout(w_dff_B_HKZYHUZX9_2),.clk(gclk));
	jdff dff_B_nGncQTUi1_2(.din(w_dff_B_HKZYHUZX9_2),.dout(w_dff_B_nGncQTUi1_2),.clk(gclk));
	jdff dff_B_rwrnzylx8_2(.din(w_dff_B_nGncQTUi1_2),.dout(w_dff_B_rwrnzylx8_2),.clk(gclk));
	jdff dff_B_5rPQpd1L3_2(.din(w_dff_B_rwrnzylx8_2),.dout(w_dff_B_5rPQpd1L3_2),.clk(gclk));
	jdff dff_B_bExroYum5_2(.din(w_dff_B_5rPQpd1L3_2),.dout(w_dff_B_bExroYum5_2),.clk(gclk));
	jdff dff_B_yxQpWcGX6_2(.din(w_dff_B_bExroYum5_2),.dout(w_dff_B_yxQpWcGX6_2),.clk(gclk));
	jdff dff_B_higTDy5o0_2(.din(w_dff_B_yxQpWcGX6_2),.dout(w_dff_B_higTDy5o0_2),.clk(gclk));
	jdff dff_B_lL1HJHi17_2(.din(w_dff_B_higTDy5o0_2),.dout(w_dff_B_lL1HJHi17_2),.clk(gclk));
	jdff dff_B_uqQT0TR96_2(.din(w_dff_B_lL1HJHi17_2),.dout(w_dff_B_uqQT0TR96_2),.clk(gclk));
	jdff dff_B_MoL9CwpP0_2(.din(w_dff_B_uqQT0TR96_2),.dout(w_dff_B_MoL9CwpP0_2),.clk(gclk));
	jdff dff_B_N4JfSr7n1_1(.din(n1623),.dout(w_dff_B_N4JfSr7n1_1),.clk(gclk));
	jdff dff_B_5qq234Sr4_1(.din(w_dff_B_N4JfSr7n1_1),.dout(w_dff_B_5qq234Sr4_1),.clk(gclk));
	jdff dff_B_K68rkaQn9_2(.din(n1622),.dout(w_dff_B_K68rkaQn9_2),.clk(gclk));
	jdff dff_B_CiM7q6Xq9_2(.din(w_dff_B_K68rkaQn9_2),.dout(w_dff_B_CiM7q6Xq9_2),.clk(gclk));
	jdff dff_B_dkzLxwFq0_2(.din(w_dff_B_CiM7q6Xq9_2),.dout(w_dff_B_dkzLxwFq0_2),.clk(gclk));
	jdff dff_B_uDDFTSOm6_2(.din(w_dff_B_dkzLxwFq0_2),.dout(w_dff_B_uDDFTSOm6_2),.clk(gclk));
	jdff dff_B_mgJMzQa61_2(.din(w_dff_B_uDDFTSOm6_2),.dout(w_dff_B_mgJMzQa61_2),.clk(gclk));
	jdff dff_B_VrpVDPnN9_2(.din(w_dff_B_mgJMzQa61_2),.dout(w_dff_B_VrpVDPnN9_2),.clk(gclk));
	jdff dff_B_G4RSUY8j0_2(.din(w_dff_B_VrpVDPnN9_2),.dout(w_dff_B_G4RSUY8j0_2),.clk(gclk));
	jdff dff_B_4cME2GAL0_2(.din(w_dff_B_G4RSUY8j0_2),.dout(w_dff_B_4cME2GAL0_2),.clk(gclk));
	jdff dff_B_ez5PiuDK8_2(.din(w_dff_B_4cME2GAL0_2),.dout(w_dff_B_ez5PiuDK8_2),.clk(gclk));
	jdff dff_B_LLI0imW92_2(.din(w_dff_B_ez5PiuDK8_2),.dout(w_dff_B_LLI0imW92_2),.clk(gclk));
	jdff dff_B_QmHDANHS5_2(.din(w_dff_B_LLI0imW92_2),.dout(w_dff_B_QmHDANHS5_2),.clk(gclk));
	jdff dff_B_kI9ytiqq9_2(.din(w_dff_B_QmHDANHS5_2),.dout(w_dff_B_kI9ytiqq9_2),.clk(gclk));
	jdff dff_B_rjTU1pez0_2(.din(w_dff_B_kI9ytiqq9_2),.dout(w_dff_B_rjTU1pez0_2),.clk(gclk));
	jdff dff_B_lpMXW1jg1_2(.din(w_dff_B_rjTU1pez0_2),.dout(w_dff_B_lpMXW1jg1_2),.clk(gclk));
	jdff dff_B_hoUfVHa60_2(.din(w_dff_B_lpMXW1jg1_2),.dout(w_dff_B_hoUfVHa60_2),.clk(gclk));
	jdff dff_B_j0iP1Hub7_2(.din(w_dff_B_hoUfVHa60_2),.dout(w_dff_B_j0iP1Hub7_2),.clk(gclk));
	jdff dff_B_aLBmGYDK6_2(.din(w_dff_B_j0iP1Hub7_2),.dout(w_dff_B_aLBmGYDK6_2),.clk(gclk));
	jdff dff_B_fzDOd8fJ1_2(.din(w_dff_B_aLBmGYDK6_2),.dout(w_dff_B_fzDOd8fJ1_2),.clk(gclk));
	jdff dff_B_TpOVAHZl7_2(.din(w_dff_B_fzDOd8fJ1_2),.dout(w_dff_B_TpOVAHZl7_2),.clk(gclk));
	jdff dff_B_NKzhgmlF2_2(.din(w_dff_B_TpOVAHZl7_2),.dout(w_dff_B_NKzhgmlF2_2),.clk(gclk));
	jdff dff_B_bncAS4Pf5_2(.din(w_dff_B_NKzhgmlF2_2),.dout(w_dff_B_bncAS4Pf5_2),.clk(gclk));
	jdff dff_B_LlbdaGVx6_2(.din(w_dff_B_bncAS4Pf5_2),.dout(w_dff_B_LlbdaGVx6_2),.clk(gclk));
	jdff dff_B_u1oLIKQV6_2(.din(w_dff_B_LlbdaGVx6_2),.dout(w_dff_B_u1oLIKQV6_2),.clk(gclk));
	jdff dff_B_uq7RaOV39_2(.din(w_dff_B_u1oLIKQV6_2),.dout(w_dff_B_uq7RaOV39_2),.clk(gclk));
	jdff dff_B_auCKxZI85_2(.din(w_dff_B_uq7RaOV39_2),.dout(w_dff_B_auCKxZI85_2),.clk(gclk));
	jdff dff_B_X5V6IUaz7_2(.din(w_dff_B_auCKxZI85_2),.dout(w_dff_B_X5V6IUaz7_2),.clk(gclk));
	jdff dff_B_eiviAIJK3_2(.din(w_dff_B_X5V6IUaz7_2),.dout(w_dff_B_eiviAIJK3_2),.clk(gclk));
	jdff dff_B_BGC8ItBU0_2(.din(w_dff_B_eiviAIJK3_2),.dout(w_dff_B_BGC8ItBU0_2),.clk(gclk));
	jdff dff_B_K35cnsZx0_2(.din(w_dff_B_BGC8ItBU0_2),.dout(w_dff_B_K35cnsZx0_2),.clk(gclk));
	jdff dff_B_WaZa6cDR7_2(.din(w_dff_B_K35cnsZx0_2),.dout(w_dff_B_WaZa6cDR7_2),.clk(gclk));
	jdff dff_B_hvBdxNAh1_2(.din(w_dff_B_WaZa6cDR7_2),.dout(w_dff_B_hvBdxNAh1_2),.clk(gclk));
	jdff dff_B_1Bs6bCOl1_2(.din(w_dff_B_hvBdxNAh1_2),.dout(w_dff_B_1Bs6bCOl1_2),.clk(gclk));
	jdff dff_B_3fu1YQq02_2(.din(w_dff_B_1Bs6bCOl1_2),.dout(w_dff_B_3fu1YQq02_2),.clk(gclk));
	jdff dff_B_R9BpI6KK7_2(.din(n1621),.dout(w_dff_B_R9BpI6KK7_2),.clk(gclk));
	jdff dff_B_rgqCiTNK7_2(.din(w_dff_B_R9BpI6KK7_2),.dout(w_dff_B_rgqCiTNK7_2),.clk(gclk));
	jdff dff_B_pW0QKm1x8_2(.din(w_dff_B_rgqCiTNK7_2),.dout(w_dff_B_pW0QKm1x8_2),.clk(gclk));
	jdff dff_B_xg1axJwk5_2(.din(w_dff_B_pW0QKm1x8_2),.dout(w_dff_B_xg1axJwk5_2),.clk(gclk));
	jdff dff_B_z8qdQBbT6_2(.din(w_dff_B_xg1axJwk5_2),.dout(w_dff_B_z8qdQBbT6_2),.clk(gclk));
	jdff dff_B_xn1SH1mG0_2(.din(w_dff_B_z8qdQBbT6_2),.dout(w_dff_B_xn1SH1mG0_2),.clk(gclk));
	jdff dff_B_0A83RMKG1_2(.din(w_dff_B_xn1SH1mG0_2),.dout(w_dff_B_0A83RMKG1_2),.clk(gclk));
	jdff dff_B_rb4pol9V8_2(.din(w_dff_B_0A83RMKG1_2),.dout(w_dff_B_rb4pol9V8_2),.clk(gclk));
	jdff dff_B_Ih7bEQca3_2(.din(w_dff_B_rb4pol9V8_2),.dout(w_dff_B_Ih7bEQca3_2),.clk(gclk));
	jdff dff_B_CXOJ9m5j8_2(.din(w_dff_B_Ih7bEQca3_2),.dout(w_dff_B_CXOJ9m5j8_2),.clk(gclk));
	jdff dff_B_AKdxi1Rf0_2(.din(w_dff_B_CXOJ9m5j8_2),.dout(w_dff_B_AKdxi1Rf0_2),.clk(gclk));
	jdff dff_B_dHN7jQjp8_2(.din(w_dff_B_AKdxi1Rf0_2),.dout(w_dff_B_dHN7jQjp8_2),.clk(gclk));
	jdff dff_B_mcPNcui82_2(.din(w_dff_B_dHN7jQjp8_2),.dout(w_dff_B_mcPNcui82_2),.clk(gclk));
	jdff dff_B_rzKFESw93_2(.din(w_dff_B_mcPNcui82_2),.dout(w_dff_B_rzKFESw93_2),.clk(gclk));
	jdff dff_B_UhrocrFL1_2(.din(w_dff_B_rzKFESw93_2),.dout(w_dff_B_UhrocrFL1_2),.clk(gclk));
	jdff dff_B_RU89xR409_2(.din(w_dff_B_UhrocrFL1_2),.dout(w_dff_B_RU89xR409_2),.clk(gclk));
	jdff dff_B_fHbRt2Nq6_2(.din(w_dff_B_RU89xR409_2),.dout(w_dff_B_fHbRt2Nq6_2),.clk(gclk));
	jdff dff_B_QJgFrR4p9_2(.din(w_dff_B_fHbRt2Nq6_2),.dout(w_dff_B_QJgFrR4p9_2),.clk(gclk));
	jdff dff_B_Sxvk3fOd2_2(.din(w_dff_B_QJgFrR4p9_2),.dout(w_dff_B_Sxvk3fOd2_2),.clk(gclk));
	jdff dff_B_pMUf683H6_2(.din(w_dff_B_Sxvk3fOd2_2),.dout(w_dff_B_pMUf683H6_2),.clk(gclk));
	jdff dff_B_2pLBPppL5_2(.din(w_dff_B_pMUf683H6_2),.dout(w_dff_B_2pLBPppL5_2),.clk(gclk));
	jdff dff_B_jsv79wMI0_2(.din(w_dff_B_2pLBPppL5_2),.dout(w_dff_B_jsv79wMI0_2),.clk(gclk));
	jdff dff_B_8vTgenk18_2(.din(w_dff_B_jsv79wMI0_2),.dout(w_dff_B_8vTgenk18_2),.clk(gclk));
	jdff dff_B_V1SX7UNt0_2(.din(w_dff_B_8vTgenk18_2),.dout(w_dff_B_V1SX7UNt0_2),.clk(gclk));
	jdff dff_B_31X9wV946_2(.din(w_dff_B_V1SX7UNt0_2),.dout(w_dff_B_31X9wV946_2),.clk(gclk));
	jdff dff_B_3NQYAGCw8_2(.din(w_dff_B_31X9wV946_2),.dout(w_dff_B_3NQYAGCw8_2),.clk(gclk));
	jdff dff_B_zSEpyaj96_2(.din(w_dff_B_3NQYAGCw8_2),.dout(w_dff_B_zSEpyaj96_2),.clk(gclk));
	jdff dff_B_HKUMPwgn9_2(.din(w_dff_B_zSEpyaj96_2),.dout(w_dff_B_HKUMPwgn9_2),.clk(gclk));
	jdff dff_B_o7bljNKx1_2(.din(w_dff_B_HKUMPwgn9_2),.dout(w_dff_B_o7bljNKx1_2),.clk(gclk));
	jdff dff_B_vBkPOOmw4_2(.din(w_dff_B_o7bljNKx1_2),.dout(w_dff_B_vBkPOOmw4_2),.clk(gclk));
	jdff dff_B_QtazNloG8_2(.din(w_dff_B_vBkPOOmw4_2),.dout(w_dff_B_QtazNloG8_2),.clk(gclk));
	jdff dff_B_rRJOtmUo5_2(.din(w_dff_B_QtazNloG8_2),.dout(w_dff_B_rRJOtmUo5_2),.clk(gclk));
	jdff dff_B_tid6EDcB4_2(.din(w_dff_B_rRJOtmUo5_2),.dout(w_dff_B_tid6EDcB4_2),.clk(gclk));
	jdff dff_B_ThuaIvl45_2(.din(w_dff_B_tid6EDcB4_2),.dout(w_dff_B_ThuaIvl45_2),.clk(gclk));
	jdff dff_B_UxFdy8pr2_2(.din(w_dff_B_ThuaIvl45_2),.dout(w_dff_B_UxFdy8pr2_2),.clk(gclk));
	jdff dff_B_S9b9GWiV5_2(.din(n1620),.dout(w_dff_B_S9b9GWiV5_2),.clk(gclk));
	jdff dff_B_HJZteJoN3_1(.din(n1618),.dout(w_dff_B_HJZteJoN3_1),.clk(gclk));
	jdff dff_B_OmvMAqTT0_2(.din(n1560),.dout(w_dff_B_OmvMAqTT0_2),.clk(gclk));
	jdff dff_B_pvsZFsx15_2(.din(w_dff_B_OmvMAqTT0_2),.dout(w_dff_B_pvsZFsx15_2),.clk(gclk));
	jdff dff_B_AXr4O4ty0_2(.din(w_dff_B_pvsZFsx15_2),.dout(w_dff_B_AXr4O4ty0_2),.clk(gclk));
	jdff dff_B_862N7lLh1_2(.din(w_dff_B_AXr4O4ty0_2),.dout(w_dff_B_862N7lLh1_2),.clk(gclk));
	jdff dff_B_P7AhAO7I5_2(.din(w_dff_B_862N7lLh1_2),.dout(w_dff_B_P7AhAO7I5_2),.clk(gclk));
	jdff dff_B_x1kZzuYt4_2(.din(w_dff_B_P7AhAO7I5_2),.dout(w_dff_B_x1kZzuYt4_2),.clk(gclk));
	jdff dff_B_XKApxCph2_2(.din(w_dff_B_x1kZzuYt4_2),.dout(w_dff_B_XKApxCph2_2),.clk(gclk));
	jdff dff_B_JaHfiVvu5_2(.din(w_dff_B_XKApxCph2_2),.dout(w_dff_B_JaHfiVvu5_2),.clk(gclk));
	jdff dff_B_yvXraZ4b0_2(.din(w_dff_B_JaHfiVvu5_2),.dout(w_dff_B_yvXraZ4b0_2),.clk(gclk));
	jdff dff_B_osxJEzY77_2(.din(w_dff_B_yvXraZ4b0_2),.dout(w_dff_B_osxJEzY77_2),.clk(gclk));
	jdff dff_B_gtYJYOf66_2(.din(w_dff_B_osxJEzY77_2),.dout(w_dff_B_gtYJYOf66_2),.clk(gclk));
	jdff dff_B_XqkQqxjt0_2(.din(w_dff_B_gtYJYOf66_2),.dout(w_dff_B_XqkQqxjt0_2),.clk(gclk));
	jdff dff_B_Oh9Z1gqE0_2(.din(w_dff_B_XqkQqxjt0_2),.dout(w_dff_B_Oh9Z1gqE0_2),.clk(gclk));
	jdff dff_B_sJ956VoH2_2(.din(w_dff_B_Oh9Z1gqE0_2),.dout(w_dff_B_sJ956VoH2_2),.clk(gclk));
	jdff dff_B_NFSfL3w03_2(.din(w_dff_B_sJ956VoH2_2),.dout(w_dff_B_NFSfL3w03_2),.clk(gclk));
	jdff dff_B_bhMsQ0N37_2(.din(w_dff_B_NFSfL3w03_2),.dout(w_dff_B_bhMsQ0N37_2),.clk(gclk));
	jdff dff_B_dWoWhe207_2(.din(w_dff_B_bhMsQ0N37_2),.dout(w_dff_B_dWoWhe207_2),.clk(gclk));
	jdff dff_B_7FrM7QSE4_2(.din(w_dff_B_dWoWhe207_2),.dout(w_dff_B_7FrM7QSE4_2),.clk(gclk));
	jdff dff_B_jp38REXl8_2(.din(w_dff_B_7FrM7QSE4_2),.dout(w_dff_B_jp38REXl8_2),.clk(gclk));
	jdff dff_B_JVrL0fzG6_2(.din(w_dff_B_jp38REXl8_2),.dout(w_dff_B_JVrL0fzG6_2),.clk(gclk));
	jdff dff_B_rgx8hFa92_2(.din(w_dff_B_JVrL0fzG6_2),.dout(w_dff_B_rgx8hFa92_2),.clk(gclk));
	jdff dff_B_mqpK7Xad6_2(.din(w_dff_B_rgx8hFa92_2),.dout(w_dff_B_mqpK7Xad6_2),.clk(gclk));
	jdff dff_B_zeToHgRv0_2(.din(w_dff_B_mqpK7Xad6_2),.dout(w_dff_B_zeToHgRv0_2),.clk(gclk));
	jdff dff_B_EbJNOq1D7_2(.din(w_dff_B_zeToHgRv0_2),.dout(w_dff_B_EbJNOq1D7_2),.clk(gclk));
	jdff dff_B_ZIMh5qSI7_2(.din(w_dff_B_EbJNOq1D7_2),.dout(w_dff_B_ZIMh5qSI7_2),.clk(gclk));
	jdff dff_B_Ln9EsESf0_2(.din(w_dff_B_ZIMh5qSI7_2),.dout(w_dff_B_Ln9EsESf0_2),.clk(gclk));
	jdff dff_B_trsadETY7_2(.din(w_dff_B_Ln9EsESf0_2),.dout(w_dff_B_trsadETY7_2),.clk(gclk));
	jdff dff_B_xqcF2OXE4_2(.din(w_dff_B_trsadETY7_2),.dout(w_dff_B_xqcF2OXE4_2),.clk(gclk));
	jdff dff_B_LCJfPLE72_2(.din(w_dff_B_xqcF2OXE4_2),.dout(w_dff_B_LCJfPLE72_2),.clk(gclk));
	jdff dff_B_snsH9h506_2(.din(w_dff_B_LCJfPLE72_2),.dout(w_dff_B_snsH9h506_2),.clk(gclk));
	jdff dff_B_If3bHUL46_2(.din(w_dff_B_snsH9h506_2),.dout(w_dff_B_If3bHUL46_2),.clk(gclk));
	jdff dff_B_vCWHOO814_2(.din(w_dff_B_If3bHUL46_2),.dout(w_dff_B_vCWHOO814_2),.clk(gclk));
	jdff dff_B_lyZCPGs11_1(.din(n1566),.dout(w_dff_B_lyZCPGs11_1),.clk(gclk));
	jdff dff_B_R8uxWo708_1(.din(w_dff_B_lyZCPGs11_1),.dout(w_dff_B_R8uxWo708_1),.clk(gclk));
	jdff dff_B_46WPqBBn2_2(.din(n1565),.dout(w_dff_B_46WPqBBn2_2),.clk(gclk));
	jdff dff_B_1XWtqaD66_2(.din(w_dff_B_46WPqBBn2_2),.dout(w_dff_B_1XWtqaD66_2),.clk(gclk));
	jdff dff_B_knW16qmU7_2(.din(w_dff_B_1XWtqaD66_2),.dout(w_dff_B_knW16qmU7_2),.clk(gclk));
	jdff dff_B_4GCSMxTt4_2(.din(w_dff_B_knW16qmU7_2),.dout(w_dff_B_4GCSMxTt4_2),.clk(gclk));
	jdff dff_B_bcXDzk9i8_2(.din(w_dff_B_4GCSMxTt4_2),.dout(w_dff_B_bcXDzk9i8_2),.clk(gclk));
	jdff dff_B_ssevscCk1_2(.din(w_dff_B_bcXDzk9i8_2),.dout(w_dff_B_ssevscCk1_2),.clk(gclk));
	jdff dff_B_t9CUpARs6_2(.din(w_dff_B_ssevscCk1_2),.dout(w_dff_B_t9CUpARs6_2),.clk(gclk));
	jdff dff_B_PKkvjSv16_2(.din(w_dff_B_t9CUpARs6_2),.dout(w_dff_B_PKkvjSv16_2),.clk(gclk));
	jdff dff_B_1tQLeOoh5_2(.din(w_dff_B_PKkvjSv16_2),.dout(w_dff_B_1tQLeOoh5_2),.clk(gclk));
	jdff dff_B_iQ0u0b7B8_2(.din(w_dff_B_1tQLeOoh5_2),.dout(w_dff_B_iQ0u0b7B8_2),.clk(gclk));
	jdff dff_B_2HVBPVYn0_2(.din(w_dff_B_iQ0u0b7B8_2),.dout(w_dff_B_2HVBPVYn0_2),.clk(gclk));
	jdff dff_B_Tmz9uCix5_2(.din(w_dff_B_2HVBPVYn0_2),.dout(w_dff_B_Tmz9uCix5_2),.clk(gclk));
	jdff dff_B_1a7KvG528_2(.din(w_dff_B_Tmz9uCix5_2),.dout(w_dff_B_1a7KvG528_2),.clk(gclk));
	jdff dff_B_Y5s6eiW44_2(.din(w_dff_B_1a7KvG528_2),.dout(w_dff_B_Y5s6eiW44_2),.clk(gclk));
	jdff dff_B_kqvOaVKo7_2(.din(w_dff_B_Y5s6eiW44_2),.dout(w_dff_B_kqvOaVKo7_2),.clk(gclk));
	jdff dff_B_r9B0GuIM5_2(.din(w_dff_B_kqvOaVKo7_2),.dout(w_dff_B_r9B0GuIM5_2),.clk(gclk));
	jdff dff_B_ostB113k4_2(.din(w_dff_B_r9B0GuIM5_2),.dout(w_dff_B_ostB113k4_2),.clk(gclk));
	jdff dff_B_ivdue0726_2(.din(w_dff_B_ostB113k4_2),.dout(w_dff_B_ivdue0726_2),.clk(gclk));
	jdff dff_B_SbTmByqZ9_2(.din(w_dff_B_ivdue0726_2),.dout(w_dff_B_SbTmByqZ9_2),.clk(gclk));
	jdff dff_B_UpzIo9X63_2(.din(w_dff_B_SbTmByqZ9_2),.dout(w_dff_B_UpzIo9X63_2),.clk(gclk));
	jdff dff_B_9M1mJqd92_2(.din(w_dff_B_UpzIo9X63_2),.dout(w_dff_B_9M1mJqd92_2),.clk(gclk));
	jdff dff_B_1jWpo7Xj0_2(.din(w_dff_B_9M1mJqd92_2),.dout(w_dff_B_1jWpo7Xj0_2),.clk(gclk));
	jdff dff_B_AGK4g5ti1_2(.din(w_dff_B_1jWpo7Xj0_2),.dout(w_dff_B_AGK4g5ti1_2),.clk(gclk));
	jdff dff_B_vcJ09U567_2(.din(w_dff_B_AGK4g5ti1_2),.dout(w_dff_B_vcJ09U567_2),.clk(gclk));
	jdff dff_B_uhJs6o5p9_2(.din(w_dff_B_vcJ09U567_2),.dout(w_dff_B_uhJs6o5p9_2),.clk(gclk));
	jdff dff_B_ZgdaOcBh9_2(.din(w_dff_B_uhJs6o5p9_2),.dout(w_dff_B_ZgdaOcBh9_2),.clk(gclk));
	jdff dff_B_N5MWngKd2_2(.din(w_dff_B_ZgdaOcBh9_2),.dout(w_dff_B_N5MWngKd2_2),.clk(gclk));
	jdff dff_B_BtMKTer00_2(.din(w_dff_B_N5MWngKd2_2),.dout(w_dff_B_BtMKTer00_2),.clk(gclk));
	jdff dff_B_00H811zv5_2(.din(w_dff_B_BtMKTer00_2),.dout(w_dff_B_00H811zv5_2),.clk(gclk));
	jdff dff_B_XI8wn8Uu3_2(.din(n1564),.dout(w_dff_B_XI8wn8Uu3_2),.clk(gclk));
	jdff dff_B_7BwIwi7Z2_2(.din(w_dff_B_XI8wn8Uu3_2),.dout(w_dff_B_7BwIwi7Z2_2),.clk(gclk));
	jdff dff_B_K3tdjOh04_2(.din(w_dff_B_7BwIwi7Z2_2),.dout(w_dff_B_K3tdjOh04_2),.clk(gclk));
	jdff dff_B_nluhx48n8_2(.din(w_dff_B_K3tdjOh04_2),.dout(w_dff_B_nluhx48n8_2),.clk(gclk));
	jdff dff_B_NZIDjwhe7_2(.din(w_dff_B_nluhx48n8_2),.dout(w_dff_B_NZIDjwhe7_2),.clk(gclk));
	jdff dff_B_Zffxkm2s6_2(.din(w_dff_B_NZIDjwhe7_2),.dout(w_dff_B_Zffxkm2s6_2),.clk(gclk));
	jdff dff_B_1phQhY8Q9_2(.din(w_dff_B_Zffxkm2s6_2),.dout(w_dff_B_1phQhY8Q9_2),.clk(gclk));
	jdff dff_B_xKjVvZqP4_2(.din(w_dff_B_1phQhY8Q9_2),.dout(w_dff_B_xKjVvZqP4_2),.clk(gclk));
	jdff dff_B_l0ZUqaLf9_2(.din(w_dff_B_xKjVvZqP4_2),.dout(w_dff_B_l0ZUqaLf9_2),.clk(gclk));
	jdff dff_B_MWaep3iz6_2(.din(w_dff_B_l0ZUqaLf9_2),.dout(w_dff_B_MWaep3iz6_2),.clk(gclk));
	jdff dff_B_hU9AkzUJ6_2(.din(w_dff_B_MWaep3iz6_2),.dout(w_dff_B_hU9AkzUJ6_2),.clk(gclk));
	jdff dff_B_AjQpZnQL2_2(.din(w_dff_B_hU9AkzUJ6_2),.dout(w_dff_B_AjQpZnQL2_2),.clk(gclk));
	jdff dff_B_JC37OW3r9_2(.din(w_dff_B_AjQpZnQL2_2),.dout(w_dff_B_JC37OW3r9_2),.clk(gclk));
	jdff dff_B_hXM82lQv5_2(.din(w_dff_B_JC37OW3r9_2),.dout(w_dff_B_hXM82lQv5_2),.clk(gclk));
	jdff dff_B_TVfRBuFz0_2(.din(w_dff_B_hXM82lQv5_2),.dout(w_dff_B_TVfRBuFz0_2),.clk(gclk));
	jdff dff_B_4bp5GJi99_2(.din(w_dff_B_TVfRBuFz0_2),.dout(w_dff_B_4bp5GJi99_2),.clk(gclk));
	jdff dff_B_a1Q1jioX6_2(.din(w_dff_B_4bp5GJi99_2),.dout(w_dff_B_a1Q1jioX6_2),.clk(gclk));
	jdff dff_B_lUUGNdUr8_2(.din(w_dff_B_a1Q1jioX6_2),.dout(w_dff_B_lUUGNdUr8_2),.clk(gclk));
	jdff dff_B_fLdWDGxq5_2(.din(w_dff_B_lUUGNdUr8_2),.dout(w_dff_B_fLdWDGxq5_2),.clk(gclk));
	jdff dff_B_2m5bpYii5_2(.din(w_dff_B_fLdWDGxq5_2),.dout(w_dff_B_2m5bpYii5_2),.clk(gclk));
	jdff dff_B_NTT9AYFE1_2(.din(w_dff_B_2m5bpYii5_2),.dout(w_dff_B_NTT9AYFE1_2),.clk(gclk));
	jdff dff_B_g3vSHVBW2_2(.din(w_dff_B_NTT9AYFE1_2),.dout(w_dff_B_g3vSHVBW2_2),.clk(gclk));
	jdff dff_B_f1BJmZyr2_2(.din(w_dff_B_g3vSHVBW2_2),.dout(w_dff_B_f1BJmZyr2_2),.clk(gclk));
	jdff dff_B_ZJaPvM3o5_2(.din(w_dff_B_f1BJmZyr2_2),.dout(w_dff_B_ZJaPvM3o5_2),.clk(gclk));
	jdff dff_B_KDPqWNWF0_2(.din(w_dff_B_ZJaPvM3o5_2),.dout(w_dff_B_KDPqWNWF0_2),.clk(gclk));
	jdff dff_B_kTuf7nG95_2(.din(w_dff_B_KDPqWNWF0_2),.dout(w_dff_B_kTuf7nG95_2),.clk(gclk));
	jdff dff_B_lCJyOdvc2_2(.din(w_dff_B_kTuf7nG95_2),.dout(w_dff_B_lCJyOdvc2_2),.clk(gclk));
	jdff dff_B_IH3DPNQ59_2(.din(w_dff_B_lCJyOdvc2_2),.dout(w_dff_B_IH3DPNQ59_2),.clk(gclk));
	jdff dff_B_dymqQGsn2_2(.din(w_dff_B_IH3DPNQ59_2),.dout(w_dff_B_dymqQGsn2_2),.clk(gclk));
	jdff dff_B_6ELLYYeu3_2(.din(w_dff_B_dymqQGsn2_2),.dout(w_dff_B_6ELLYYeu3_2),.clk(gclk));
	jdff dff_B_VtqpH4MQ5_2(.din(w_dff_B_6ELLYYeu3_2),.dout(w_dff_B_VtqpH4MQ5_2),.clk(gclk));
	jdff dff_B_ipKRWSpy6_2(.din(n1563),.dout(w_dff_B_ipKRWSpy6_2),.clk(gclk));
	jdff dff_B_plcpmFsX2_1(.din(n1561),.dout(w_dff_B_plcpmFsX2_1),.clk(gclk));
	jdff dff_B_Av03ybjv7_2(.din(n1496),.dout(w_dff_B_Av03ybjv7_2),.clk(gclk));
	jdff dff_B_TOXOZ8v72_2(.din(w_dff_B_Av03ybjv7_2),.dout(w_dff_B_TOXOZ8v72_2),.clk(gclk));
	jdff dff_B_8NNliQ6X1_2(.din(w_dff_B_TOXOZ8v72_2),.dout(w_dff_B_8NNliQ6X1_2),.clk(gclk));
	jdff dff_B_zKqFceEj0_2(.din(w_dff_B_8NNliQ6X1_2),.dout(w_dff_B_zKqFceEj0_2),.clk(gclk));
	jdff dff_B_u8HlRG636_2(.din(w_dff_B_zKqFceEj0_2),.dout(w_dff_B_u8HlRG636_2),.clk(gclk));
	jdff dff_B_1CTfZ9rO2_2(.din(w_dff_B_u8HlRG636_2),.dout(w_dff_B_1CTfZ9rO2_2),.clk(gclk));
	jdff dff_B_NFOgvyNk0_2(.din(w_dff_B_1CTfZ9rO2_2),.dout(w_dff_B_NFOgvyNk0_2),.clk(gclk));
	jdff dff_B_l4BH1Z9j0_2(.din(w_dff_B_NFOgvyNk0_2),.dout(w_dff_B_l4BH1Z9j0_2),.clk(gclk));
	jdff dff_B_ps38PL8f9_2(.din(w_dff_B_l4BH1Z9j0_2),.dout(w_dff_B_ps38PL8f9_2),.clk(gclk));
	jdff dff_B_3yStKIJO4_2(.din(w_dff_B_ps38PL8f9_2),.dout(w_dff_B_3yStKIJO4_2),.clk(gclk));
	jdff dff_B_vekcYn1c4_2(.din(w_dff_B_3yStKIJO4_2),.dout(w_dff_B_vekcYn1c4_2),.clk(gclk));
	jdff dff_B_rUxGzJKf2_2(.din(w_dff_B_vekcYn1c4_2),.dout(w_dff_B_rUxGzJKf2_2),.clk(gclk));
	jdff dff_B_0GKuh1zB5_2(.din(w_dff_B_rUxGzJKf2_2),.dout(w_dff_B_0GKuh1zB5_2),.clk(gclk));
	jdff dff_B_8JPsKB0k2_2(.din(w_dff_B_0GKuh1zB5_2),.dout(w_dff_B_8JPsKB0k2_2),.clk(gclk));
	jdff dff_B_dx6bcf6z5_2(.din(w_dff_B_8JPsKB0k2_2),.dout(w_dff_B_dx6bcf6z5_2),.clk(gclk));
	jdff dff_B_O1DiOXmJ6_2(.din(w_dff_B_dx6bcf6z5_2),.dout(w_dff_B_O1DiOXmJ6_2),.clk(gclk));
	jdff dff_B_vkte66X21_2(.din(w_dff_B_O1DiOXmJ6_2),.dout(w_dff_B_vkte66X21_2),.clk(gclk));
	jdff dff_B_aDINbv7V1_2(.din(w_dff_B_vkte66X21_2),.dout(w_dff_B_aDINbv7V1_2),.clk(gclk));
	jdff dff_B_WzghUl385_2(.din(w_dff_B_aDINbv7V1_2),.dout(w_dff_B_WzghUl385_2),.clk(gclk));
	jdff dff_B_z03Ap8BX4_2(.din(w_dff_B_WzghUl385_2),.dout(w_dff_B_z03Ap8BX4_2),.clk(gclk));
	jdff dff_B_WwKReFR89_2(.din(w_dff_B_z03Ap8BX4_2),.dout(w_dff_B_WwKReFR89_2),.clk(gclk));
	jdff dff_B_0huAPqU41_2(.din(w_dff_B_WwKReFR89_2),.dout(w_dff_B_0huAPqU41_2),.clk(gclk));
	jdff dff_B_ucANHPEB7_2(.din(w_dff_B_0huAPqU41_2),.dout(w_dff_B_ucANHPEB7_2),.clk(gclk));
	jdff dff_B_ULZfgP8H2_2(.din(w_dff_B_ucANHPEB7_2),.dout(w_dff_B_ULZfgP8H2_2),.clk(gclk));
	jdff dff_B_hsgHv1xE6_2(.din(w_dff_B_ULZfgP8H2_2),.dout(w_dff_B_hsgHv1xE6_2),.clk(gclk));
	jdff dff_B_aIIDjXAm4_2(.din(w_dff_B_hsgHv1xE6_2),.dout(w_dff_B_aIIDjXAm4_2),.clk(gclk));
	jdff dff_B_9CVhahh19_2(.din(w_dff_B_aIIDjXAm4_2),.dout(w_dff_B_9CVhahh19_2),.clk(gclk));
	jdff dff_B_B2JJaT8Y1_2(.din(w_dff_B_9CVhahh19_2),.dout(w_dff_B_B2JJaT8Y1_2),.clk(gclk));
	jdff dff_B_YFMKMXf99_1(.din(n1502),.dout(w_dff_B_YFMKMXf99_1),.clk(gclk));
	jdff dff_B_zBIB7LIv3_1(.din(w_dff_B_YFMKMXf99_1),.dout(w_dff_B_zBIB7LIv3_1),.clk(gclk));
	jdff dff_B_2lupi1eT7_2(.din(n1501),.dout(w_dff_B_2lupi1eT7_2),.clk(gclk));
	jdff dff_B_lDeJkaEL8_2(.din(w_dff_B_2lupi1eT7_2),.dout(w_dff_B_lDeJkaEL8_2),.clk(gclk));
	jdff dff_B_m2ps2aC25_2(.din(w_dff_B_lDeJkaEL8_2),.dout(w_dff_B_m2ps2aC25_2),.clk(gclk));
	jdff dff_B_QmTK3o6b0_2(.din(w_dff_B_m2ps2aC25_2),.dout(w_dff_B_QmTK3o6b0_2),.clk(gclk));
	jdff dff_B_Z0VOmMi61_2(.din(w_dff_B_QmTK3o6b0_2),.dout(w_dff_B_Z0VOmMi61_2),.clk(gclk));
	jdff dff_B_XLWiyqa95_2(.din(w_dff_B_Z0VOmMi61_2),.dout(w_dff_B_XLWiyqa95_2),.clk(gclk));
	jdff dff_B_EA0yKMqT5_2(.din(w_dff_B_XLWiyqa95_2),.dout(w_dff_B_EA0yKMqT5_2),.clk(gclk));
	jdff dff_B_uYntsCLe6_2(.din(w_dff_B_EA0yKMqT5_2),.dout(w_dff_B_uYntsCLe6_2),.clk(gclk));
	jdff dff_B_W7xGSPqc6_2(.din(w_dff_B_uYntsCLe6_2),.dout(w_dff_B_W7xGSPqc6_2),.clk(gclk));
	jdff dff_B_8BqnZydY8_2(.din(w_dff_B_W7xGSPqc6_2),.dout(w_dff_B_8BqnZydY8_2),.clk(gclk));
	jdff dff_B_KTe0YBW91_2(.din(w_dff_B_8BqnZydY8_2),.dout(w_dff_B_KTe0YBW91_2),.clk(gclk));
	jdff dff_B_TDNCuHUh6_2(.din(w_dff_B_KTe0YBW91_2),.dout(w_dff_B_TDNCuHUh6_2),.clk(gclk));
	jdff dff_B_F7zplMgm0_2(.din(w_dff_B_TDNCuHUh6_2),.dout(w_dff_B_F7zplMgm0_2),.clk(gclk));
	jdff dff_B_7ziRD5KS4_2(.din(w_dff_B_F7zplMgm0_2),.dout(w_dff_B_7ziRD5KS4_2),.clk(gclk));
	jdff dff_B_Zhr77VUE0_2(.din(w_dff_B_7ziRD5KS4_2),.dout(w_dff_B_Zhr77VUE0_2),.clk(gclk));
	jdff dff_B_HvIRCMU08_2(.din(w_dff_B_Zhr77VUE0_2),.dout(w_dff_B_HvIRCMU08_2),.clk(gclk));
	jdff dff_B_Pak5dTBC9_2(.din(w_dff_B_HvIRCMU08_2),.dout(w_dff_B_Pak5dTBC9_2),.clk(gclk));
	jdff dff_B_s7w1pX6x4_2(.din(w_dff_B_Pak5dTBC9_2),.dout(w_dff_B_s7w1pX6x4_2),.clk(gclk));
	jdff dff_B_rlNnwseh7_2(.din(w_dff_B_s7w1pX6x4_2),.dout(w_dff_B_rlNnwseh7_2),.clk(gclk));
	jdff dff_B_0GkVLFEq5_2(.din(w_dff_B_rlNnwseh7_2),.dout(w_dff_B_0GkVLFEq5_2),.clk(gclk));
	jdff dff_B_I4XY41NH0_2(.din(w_dff_B_0GkVLFEq5_2),.dout(w_dff_B_I4XY41NH0_2),.clk(gclk));
	jdff dff_B_8NyDsdmn2_2(.din(w_dff_B_I4XY41NH0_2),.dout(w_dff_B_8NyDsdmn2_2),.clk(gclk));
	jdff dff_B_8Ql4FxcU6_2(.din(w_dff_B_8NyDsdmn2_2),.dout(w_dff_B_8Ql4FxcU6_2),.clk(gclk));
	jdff dff_B_l6HYqmoc5_2(.din(w_dff_B_8Ql4FxcU6_2),.dout(w_dff_B_l6HYqmoc5_2),.clk(gclk));
	jdff dff_B_7pxHhch97_2(.din(w_dff_B_l6HYqmoc5_2),.dout(w_dff_B_7pxHhch97_2),.clk(gclk));
	jdff dff_B_A2NDWBwO0_2(.din(n1500),.dout(w_dff_B_A2NDWBwO0_2),.clk(gclk));
	jdff dff_B_YNYkrfAJ7_2(.din(w_dff_B_A2NDWBwO0_2),.dout(w_dff_B_YNYkrfAJ7_2),.clk(gclk));
	jdff dff_B_bN5RRWSv1_2(.din(w_dff_B_YNYkrfAJ7_2),.dout(w_dff_B_bN5RRWSv1_2),.clk(gclk));
	jdff dff_B_QlHe1He51_2(.din(w_dff_B_bN5RRWSv1_2),.dout(w_dff_B_QlHe1He51_2),.clk(gclk));
	jdff dff_B_g9NgCkTW4_2(.din(w_dff_B_QlHe1He51_2),.dout(w_dff_B_g9NgCkTW4_2),.clk(gclk));
	jdff dff_B_A4GuylTi0_2(.din(w_dff_B_g9NgCkTW4_2),.dout(w_dff_B_A4GuylTi0_2),.clk(gclk));
	jdff dff_B_U0GPJpZ77_2(.din(w_dff_B_A4GuylTi0_2),.dout(w_dff_B_U0GPJpZ77_2),.clk(gclk));
	jdff dff_B_fZoFfEII8_2(.din(w_dff_B_U0GPJpZ77_2),.dout(w_dff_B_fZoFfEII8_2),.clk(gclk));
	jdff dff_B_HUKTMELg4_2(.din(w_dff_B_fZoFfEII8_2),.dout(w_dff_B_HUKTMELg4_2),.clk(gclk));
	jdff dff_B_jqEcdhi14_2(.din(w_dff_B_HUKTMELg4_2),.dout(w_dff_B_jqEcdhi14_2),.clk(gclk));
	jdff dff_B_z3aWz5gU4_2(.din(w_dff_B_jqEcdhi14_2),.dout(w_dff_B_z3aWz5gU4_2),.clk(gclk));
	jdff dff_B_GoEvd0vC6_2(.din(w_dff_B_z3aWz5gU4_2),.dout(w_dff_B_GoEvd0vC6_2),.clk(gclk));
	jdff dff_B_AYPZjyLs3_2(.din(w_dff_B_GoEvd0vC6_2),.dout(w_dff_B_AYPZjyLs3_2),.clk(gclk));
	jdff dff_B_YE4EL8mj1_2(.din(w_dff_B_AYPZjyLs3_2),.dout(w_dff_B_YE4EL8mj1_2),.clk(gclk));
	jdff dff_B_WzOT6QaG6_2(.din(w_dff_B_YE4EL8mj1_2),.dout(w_dff_B_WzOT6QaG6_2),.clk(gclk));
	jdff dff_B_efoCT5ku6_2(.din(w_dff_B_WzOT6QaG6_2),.dout(w_dff_B_efoCT5ku6_2),.clk(gclk));
	jdff dff_B_jD55L0qG7_2(.din(w_dff_B_efoCT5ku6_2),.dout(w_dff_B_jD55L0qG7_2),.clk(gclk));
	jdff dff_B_QFmHvdPf5_2(.din(w_dff_B_jD55L0qG7_2),.dout(w_dff_B_QFmHvdPf5_2),.clk(gclk));
	jdff dff_B_VOFMawPP0_2(.din(w_dff_B_QFmHvdPf5_2),.dout(w_dff_B_VOFMawPP0_2),.clk(gclk));
	jdff dff_B_iiUpzoe22_2(.din(w_dff_B_VOFMawPP0_2),.dout(w_dff_B_iiUpzoe22_2),.clk(gclk));
	jdff dff_B_Y30VZ7cH5_2(.din(w_dff_B_iiUpzoe22_2),.dout(w_dff_B_Y30VZ7cH5_2),.clk(gclk));
	jdff dff_B_wgDX7S5p8_2(.din(w_dff_B_Y30VZ7cH5_2),.dout(w_dff_B_wgDX7S5p8_2),.clk(gclk));
	jdff dff_B_uOzOINEo1_2(.din(w_dff_B_wgDX7S5p8_2),.dout(w_dff_B_uOzOINEo1_2),.clk(gclk));
	jdff dff_B_pmP1MQka3_2(.din(w_dff_B_uOzOINEo1_2),.dout(w_dff_B_pmP1MQka3_2),.clk(gclk));
	jdff dff_B_lCFVNw2c2_2(.din(w_dff_B_pmP1MQka3_2),.dout(w_dff_B_lCFVNw2c2_2),.clk(gclk));
	jdff dff_B_Jm9w6RiA2_2(.din(w_dff_B_lCFVNw2c2_2),.dout(w_dff_B_Jm9w6RiA2_2),.clk(gclk));
	jdff dff_B_2BeACS201_2(.din(w_dff_B_Jm9w6RiA2_2),.dout(w_dff_B_2BeACS201_2),.clk(gclk));
	jdff dff_B_8HqNMCiP7_2(.din(n1499),.dout(w_dff_B_8HqNMCiP7_2),.clk(gclk));
	jdff dff_B_S026EZg56_1(.din(n1497),.dout(w_dff_B_S026EZg56_1),.clk(gclk));
	jdff dff_B_II4gFpzY7_2(.din(n1425),.dout(w_dff_B_II4gFpzY7_2),.clk(gclk));
	jdff dff_B_p6KibwD58_2(.din(w_dff_B_II4gFpzY7_2),.dout(w_dff_B_p6KibwD58_2),.clk(gclk));
	jdff dff_B_0NSAln6R0_2(.din(w_dff_B_p6KibwD58_2),.dout(w_dff_B_0NSAln6R0_2),.clk(gclk));
	jdff dff_B_6GJH66ZJ3_2(.din(w_dff_B_0NSAln6R0_2),.dout(w_dff_B_6GJH66ZJ3_2),.clk(gclk));
	jdff dff_B_arL3XSj35_2(.din(w_dff_B_6GJH66ZJ3_2),.dout(w_dff_B_arL3XSj35_2),.clk(gclk));
	jdff dff_B_uXKY5agJ5_2(.din(w_dff_B_arL3XSj35_2),.dout(w_dff_B_uXKY5agJ5_2),.clk(gclk));
	jdff dff_B_C1ODHJfy8_2(.din(w_dff_B_uXKY5agJ5_2),.dout(w_dff_B_C1ODHJfy8_2),.clk(gclk));
	jdff dff_B_YPbSpx0w3_2(.din(w_dff_B_C1ODHJfy8_2),.dout(w_dff_B_YPbSpx0w3_2),.clk(gclk));
	jdff dff_B_GS2BtMHa6_2(.din(w_dff_B_YPbSpx0w3_2),.dout(w_dff_B_GS2BtMHa6_2),.clk(gclk));
	jdff dff_B_3S7Xee543_2(.din(w_dff_B_GS2BtMHa6_2),.dout(w_dff_B_3S7Xee543_2),.clk(gclk));
	jdff dff_B_YIlu3IVC2_2(.din(w_dff_B_3S7Xee543_2),.dout(w_dff_B_YIlu3IVC2_2),.clk(gclk));
	jdff dff_B_mJEY2d3L8_2(.din(w_dff_B_YIlu3IVC2_2),.dout(w_dff_B_mJEY2d3L8_2),.clk(gclk));
	jdff dff_B_BBMuspAo1_2(.din(w_dff_B_mJEY2d3L8_2),.dout(w_dff_B_BBMuspAo1_2),.clk(gclk));
	jdff dff_B_FUoJSM8P2_2(.din(w_dff_B_BBMuspAo1_2),.dout(w_dff_B_FUoJSM8P2_2),.clk(gclk));
	jdff dff_B_FarZG3x59_2(.din(w_dff_B_FUoJSM8P2_2),.dout(w_dff_B_FarZG3x59_2),.clk(gclk));
	jdff dff_B_D1blQciI4_2(.din(w_dff_B_FarZG3x59_2),.dout(w_dff_B_D1blQciI4_2),.clk(gclk));
	jdff dff_B_PSLsGNfR4_2(.din(w_dff_B_D1blQciI4_2),.dout(w_dff_B_PSLsGNfR4_2),.clk(gclk));
	jdff dff_B_GkV0GfZV3_2(.din(w_dff_B_PSLsGNfR4_2),.dout(w_dff_B_GkV0GfZV3_2),.clk(gclk));
	jdff dff_B_e2573Xix1_2(.din(w_dff_B_GkV0GfZV3_2),.dout(w_dff_B_e2573Xix1_2),.clk(gclk));
	jdff dff_B_S29BS6Mz3_2(.din(w_dff_B_e2573Xix1_2),.dout(w_dff_B_S29BS6Mz3_2),.clk(gclk));
	jdff dff_B_SLJeWLzc9_2(.din(w_dff_B_S29BS6Mz3_2),.dout(w_dff_B_SLJeWLzc9_2),.clk(gclk));
	jdff dff_B_6IidSZij5_2(.din(w_dff_B_SLJeWLzc9_2),.dout(w_dff_B_6IidSZij5_2),.clk(gclk));
	jdff dff_B_Yun8i6zT6_2(.din(w_dff_B_6IidSZij5_2),.dout(w_dff_B_Yun8i6zT6_2),.clk(gclk));
	jdff dff_B_uNJ5Rqbx3_2(.din(w_dff_B_Yun8i6zT6_2),.dout(w_dff_B_uNJ5Rqbx3_2),.clk(gclk));
	jdff dff_B_dfts3IKL9_1(.din(n1431),.dout(w_dff_B_dfts3IKL9_1),.clk(gclk));
	jdff dff_B_L7a03A1l4_1(.din(w_dff_B_dfts3IKL9_1),.dout(w_dff_B_L7a03A1l4_1),.clk(gclk));
	jdff dff_B_t5tatHDx5_2(.din(n1430),.dout(w_dff_B_t5tatHDx5_2),.clk(gclk));
	jdff dff_B_R4NCvGAC8_2(.din(w_dff_B_t5tatHDx5_2),.dout(w_dff_B_R4NCvGAC8_2),.clk(gclk));
	jdff dff_B_iXGGVD222_2(.din(w_dff_B_R4NCvGAC8_2),.dout(w_dff_B_iXGGVD222_2),.clk(gclk));
	jdff dff_B_VcZm2RMr9_2(.din(w_dff_B_iXGGVD222_2),.dout(w_dff_B_VcZm2RMr9_2),.clk(gclk));
	jdff dff_B_7DCWxgRP0_2(.din(w_dff_B_VcZm2RMr9_2),.dout(w_dff_B_7DCWxgRP0_2),.clk(gclk));
	jdff dff_B_FfpEEnUS0_2(.din(w_dff_B_7DCWxgRP0_2),.dout(w_dff_B_FfpEEnUS0_2),.clk(gclk));
	jdff dff_B_bFwnEhbF0_2(.din(w_dff_B_FfpEEnUS0_2),.dout(w_dff_B_bFwnEhbF0_2),.clk(gclk));
	jdff dff_B_xAT24ykD2_2(.din(w_dff_B_bFwnEhbF0_2),.dout(w_dff_B_xAT24ykD2_2),.clk(gclk));
	jdff dff_B_l9Ht3rWf6_2(.din(w_dff_B_xAT24ykD2_2),.dout(w_dff_B_l9Ht3rWf6_2),.clk(gclk));
	jdff dff_B_OhHNcRaJ6_2(.din(w_dff_B_l9Ht3rWf6_2),.dout(w_dff_B_OhHNcRaJ6_2),.clk(gclk));
	jdff dff_B_w8ltom5m9_2(.din(w_dff_B_OhHNcRaJ6_2),.dout(w_dff_B_w8ltom5m9_2),.clk(gclk));
	jdff dff_B_KRVmArpG9_2(.din(w_dff_B_w8ltom5m9_2),.dout(w_dff_B_KRVmArpG9_2),.clk(gclk));
	jdff dff_B_icWNlMFz9_2(.din(w_dff_B_KRVmArpG9_2),.dout(w_dff_B_icWNlMFz9_2),.clk(gclk));
	jdff dff_B_y7zRgHsx7_2(.din(w_dff_B_icWNlMFz9_2),.dout(w_dff_B_y7zRgHsx7_2),.clk(gclk));
	jdff dff_B_292f23vW9_2(.din(w_dff_B_y7zRgHsx7_2),.dout(w_dff_B_292f23vW9_2),.clk(gclk));
	jdff dff_B_lMtldrk21_2(.din(w_dff_B_292f23vW9_2),.dout(w_dff_B_lMtldrk21_2),.clk(gclk));
	jdff dff_B_V0PjiF4E6_2(.din(w_dff_B_lMtldrk21_2),.dout(w_dff_B_V0PjiF4E6_2),.clk(gclk));
	jdff dff_B_JCtWA6Zp9_2(.din(w_dff_B_V0PjiF4E6_2),.dout(w_dff_B_JCtWA6Zp9_2),.clk(gclk));
	jdff dff_B_6Kx7oBwQ2_2(.din(w_dff_B_JCtWA6Zp9_2),.dout(w_dff_B_6Kx7oBwQ2_2),.clk(gclk));
	jdff dff_B_AjSzTbXd6_2(.din(w_dff_B_6Kx7oBwQ2_2),.dout(w_dff_B_AjSzTbXd6_2),.clk(gclk));
	jdff dff_B_KO8C55j57_2(.din(w_dff_B_AjSzTbXd6_2),.dout(w_dff_B_KO8C55j57_2),.clk(gclk));
	jdff dff_B_iHBpOj256_2(.din(n1429),.dout(w_dff_B_iHBpOj256_2),.clk(gclk));
	jdff dff_B_aHWJISxO2_2(.din(w_dff_B_iHBpOj256_2),.dout(w_dff_B_aHWJISxO2_2),.clk(gclk));
	jdff dff_B_figRRYyU9_2(.din(w_dff_B_aHWJISxO2_2),.dout(w_dff_B_figRRYyU9_2),.clk(gclk));
	jdff dff_B_3ALz3QFj1_2(.din(w_dff_B_figRRYyU9_2),.dout(w_dff_B_3ALz3QFj1_2),.clk(gclk));
	jdff dff_B_ylZUh7nx1_2(.din(w_dff_B_3ALz3QFj1_2),.dout(w_dff_B_ylZUh7nx1_2),.clk(gclk));
	jdff dff_B_uJHYtz8k2_2(.din(w_dff_B_ylZUh7nx1_2),.dout(w_dff_B_uJHYtz8k2_2),.clk(gclk));
	jdff dff_B_RA6k6S0C9_2(.din(w_dff_B_uJHYtz8k2_2),.dout(w_dff_B_RA6k6S0C9_2),.clk(gclk));
	jdff dff_B_lllBzQUj4_2(.din(w_dff_B_RA6k6S0C9_2),.dout(w_dff_B_lllBzQUj4_2),.clk(gclk));
	jdff dff_B_o1bQoWKX9_2(.din(w_dff_B_lllBzQUj4_2),.dout(w_dff_B_o1bQoWKX9_2),.clk(gclk));
	jdff dff_B_qxNWYZJC9_2(.din(w_dff_B_o1bQoWKX9_2),.dout(w_dff_B_qxNWYZJC9_2),.clk(gclk));
	jdff dff_B_R9FC6olV1_2(.din(w_dff_B_qxNWYZJC9_2),.dout(w_dff_B_R9FC6olV1_2),.clk(gclk));
	jdff dff_B_NUWo2WtU2_2(.din(w_dff_B_R9FC6olV1_2),.dout(w_dff_B_NUWo2WtU2_2),.clk(gclk));
	jdff dff_B_IXZKlPZk1_2(.din(w_dff_B_NUWo2WtU2_2),.dout(w_dff_B_IXZKlPZk1_2),.clk(gclk));
	jdff dff_B_28AxlOWV2_2(.din(w_dff_B_IXZKlPZk1_2),.dout(w_dff_B_28AxlOWV2_2),.clk(gclk));
	jdff dff_B_gvtEs4qI3_2(.din(w_dff_B_28AxlOWV2_2),.dout(w_dff_B_gvtEs4qI3_2),.clk(gclk));
	jdff dff_B_n0tCGg293_2(.din(w_dff_B_gvtEs4qI3_2),.dout(w_dff_B_n0tCGg293_2),.clk(gclk));
	jdff dff_B_dfRpefxj8_2(.din(w_dff_B_n0tCGg293_2),.dout(w_dff_B_dfRpefxj8_2),.clk(gclk));
	jdff dff_B_HKAXMSIQ3_2(.din(w_dff_B_dfRpefxj8_2),.dout(w_dff_B_HKAXMSIQ3_2),.clk(gclk));
	jdff dff_B_4lF1Wtn35_2(.din(w_dff_B_HKAXMSIQ3_2),.dout(w_dff_B_4lF1Wtn35_2),.clk(gclk));
	jdff dff_B_Ywg0Cgk01_2(.din(w_dff_B_4lF1Wtn35_2),.dout(w_dff_B_Ywg0Cgk01_2),.clk(gclk));
	jdff dff_B_qDAYAYTz6_2(.din(w_dff_B_Ywg0Cgk01_2),.dout(w_dff_B_qDAYAYTz6_2),.clk(gclk));
	jdff dff_B_V6JVcxgo2_2(.din(w_dff_B_qDAYAYTz6_2),.dout(w_dff_B_V6JVcxgo2_2),.clk(gclk));
	jdff dff_B_oHPukJZ31_2(.din(w_dff_B_V6JVcxgo2_2),.dout(w_dff_B_oHPukJZ31_2),.clk(gclk));
	jdff dff_B_q8jcn1tp2_2(.din(n1428),.dout(w_dff_B_q8jcn1tp2_2),.clk(gclk));
	jdff dff_B_Ep9cpCXH0_1(.din(n1426),.dout(w_dff_B_Ep9cpCXH0_1),.clk(gclk));
	jdff dff_B_3ltbbv398_2(.din(n1347),.dout(w_dff_B_3ltbbv398_2),.clk(gclk));
	jdff dff_B_bocfXfef2_2(.din(w_dff_B_3ltbbv398_2),.dout(w_dff_B_bocfXfef2_2),.clk(gclk));
	jdff dff_B_GaYdGWsG5_2(.din(w_dff_B_bocfXfef2_2),.dout(w_dff_B_GaYdGWsG5_2),.clk(gclk));
	jdff dff_B_q9gaTcDu3_2(.din(w_dff_B_GaYdGWsG5_2),.dout(w_dff_B_q9gaTcDu3_2),.clk(gclk));
	jdff dff_B_0QW5N3qY0_2(.din(w_dff_B_q9gaTcDu3_2),.dout(w_dff_B_0QW5N3qY0_2),.clk(gclk));
	jdff dff_B_Aowu6DMd5_2(.din(w_dff_B_0QW5N3qY0_2),.dout(w_dff_B_Aowu6DMd5_2),.clk(gclk));
	jdff dff_B_GvFDmbse0_2(.din(w_dff_B_Aowu6DMd5_2),.dout(w_dff_B_GvFDmbse0_2),.clk(gclk));
	jdff dff_B_HdTcVjcR1_2(.din(w_dff_B_GvFDmbse0_2),.dout(w_dff_B_HdTcVjcR1_2),.clk(gclk));
	jdff dff_B_0JOnG4MU9_2(.din(w_dff_B_HdTcVjcR1_2),.dout(w_dff_B_0JOnG4MU9_2),.clk(gclk));
	jdff dff_B_yVQYx5ct9_2(.din(w_dff_B_0JOnG4MU9_2),.dout(w_dff_B_yVQYx5ct9_2),.clk(gclk));
	jdff dff_B_pMrb1zjr9_2(.din(w_dff_B_yVQYx5ct9_2),.dout(w_dff_B_pMrb1zjr9_2),.clk(gclk));
	jdff dff_B_w9qkHa0X9_2(.din(w_dff_B_pMrb1zjr9_2),.dout(w_dff_B_w9qkHa0X9_2),.clk(gclk));
	jdff dff_B_0wIZXfFx6_2(.din(w_dff_B_w9qkHa0X9_2),.dout(w_dff_B_0wIZXfFx6_2),.clk(gclk));
	jdff dff_B_htGTtLG31_2(.din(w_dff_B_0wIZXfFx6_2),.dout(w_dff_B_htGTtLG31_2),.clk(gclk));
	jdff dff_B_SMleNtAW7_2(.din(w_dff_B_htGTtLG31_2),.dout(w_dff_B_SMleNtAW7_2),.clk(gclk));
	jdff dff_B_E2neHheu8_2(.din(w_dff_B_SMleNtAW7_2),.dout(w_dff_B_E2neHheu8_2),.clk(gclk));
	jdff dff_B_Rmk0nzYJ5_2(.din(w_dff_B_E2neHheu8_2),.dout(w_dff_B_Rmk0nzYJ5_2),.clk(gclk));
	jdff dff_B_4zsRuMEd9_2(.din(w_dff_B_Rmk0nzYJ5_2),.dout(w_dff_B_4zsRuMEd9_2),.clk(gclk));
	jdff dff_B_qy0GjkrA5_2(.din(w_dff_B_4zsRuMEd9_2),.dout(w_dff_B_qy0GjkrA5_2),.clk(gclk));
	jdff dff_B_9qLTKO0M8_2(.din(w_dff_B_qy0GjkrA5_2),.dout(w_dff_B_9qLTKO0M8_2),.clk(gclk));
	jdff dff_B_c8bSl9KV5_1(.din(n1353),.dout(w_dff_B_c8bSl9KV5_1),.clk(gclk));
	jdff dff_B_niqKiDNW8_1(.din(w_dff_B_c8bSl9KV5_1),.dout(w_dff_B_niqKiDNW8_1),.clk(gclk));
	jdff dff_B_p0P3BqH15_2(.din(n1352),.dout(w_dff_B_p0P3BqH15_2),.clk(gclk));
	jdff dff_B_I62c8JQI2_2(.din(w_dff_B_p0P3BqH15_2),.dout(w_dff_B_I62c8JQI2_2),.clk(gclk));
	jdff dff_B_28qhwm4P8_2(.din(w_dff_B_I62c8JQI2_2),.dout(w_dff_B_28qhwm4P8_2),.clk(gclk));
	jdff dff_B_D3dcFmjD0_2(.din(w_dff_B_28qhwm4P8_2),.dout(w_dff_B_D3dcFmjD0_2),.clk(gclk));
	jdff dff_B_C1Fw9SYq6_2(.din(w_dff_B_D3dcFmjD0_2),.dout(w_dff_B_C1Fw9SYq6_2),.clk(gclk));
	jdff dff_B_CEKibw6u6_2(.din(w_dff_B_C1Fw9SYq6_2),.dout(w_dff_B_CEKibw6u6_2),.clk(gclk));
	jdff dff_B_36SM1F5p9_2(.din(w_dff_B_CEKibw6u6_2),.dout(w_dff_B_36SM1F5p9_2),.clk(gclk));
	jdff dff_B_UVad4XiN1_2(.din(w_dff_B_36SM1F5p9_2),.dout(w_dff_B_UVad4XiN1_2),.clk(gclk));
	jdff dff_B_pX10OgSl7_2(.din(w_dff_B_UVad4XiN1_2),.dout(w_dff_B_pX10OgSl7_2),.clk(gclk));
	jdff dff_B_7Ffryffh8_2(.din(w_dff_B_pX10OgSl7_2),.dout(w_dff_B_7Ffryffh8_2),.clk(gclk));
	jdff dff_B_f6WdYUHc7_2(.din(w_dff_B_7Ffryffh8_2),.dout(w_dff_B_f6WdYUHc7_2),.clk(gclk));
	jdff dff_B_P76XU3xn8_2(.din(w_dff_B_f6WdYUHc7_2),.dout(w_dff_B_P76XU3xn8_2),.clk(gclk));
	jdff dff_B_WGSPOU760_2(.din(w_dff_B_P76XU3xn8_2),.dout(w_dff_B_WGSPOU760_2),.clk(gclk));
	jdff dff_B_Nbcylzl11_2(.din(w_dff_B_WGSPOU760_2),.dout(w_dff_B_Nbcylzl11_2),.clk(gclk));
	jdff dff_B_nI0JwNwB0_2(.din(w_dff_B_Nbcylzl11_2),.dout(w_dff_B_nI0JwNwB0_2),.clk(gclk));
	jdff dff_B_NAIdpmZ68_2(.din(w_dff_B_nI0JwNwB0_2),.dout(w_dff_B_NAIdpmZ68_2),.clk(gclk));
	jdff dff_B_6BAj7eS14_2(.din(w_dff_B_NAIdpmZ68_2),.dout(w_dff_B_6BAj7eS14_2),.clk(gclk));
	jdff dff_B_YNZ0gsHV9_2(.din(n1351),.dout(w_dff_B_YNZ0gsHV9_2),.clk(gclk));
	jdff dff_B_C5oaDWd87_2(.din(w_dff_B_YNZ0gsHV9_2),.dout(w_dff_B_C5oaDWd87_2),.clk(gclk));
	jdff dff_B_sTy8tjPG0_2(.din(w_dff_B_C5oaDWd87_2),.dout(w_dff_B_sTy8tjPG0_2),.clk(gclk));
	jdff dff_B_oGCyOuvB8_2(.din(w_dff_B_sTy8tjPG0_2),.dout(w_dff_B_oGCyOuvB8_2),.clk(gclk));
	jdff dff_B_dWMT7Lpx4_2(.din(w_dff_B_oGCyOuvB8_2),.dout(w_dff_B_dWMT7Lpx4_2),.clk(gclk));
	jdff dff_B_EfmG8clW0_2(.din(w_dff_B_dWMT7Lpx4_2),.dout(w_dff_B_EfmG8clW0_2),.clk(gclk));
	jdff dff_B_qAGUZoC20_2(.din(w_dff_B_EfmG8clW0_2),.dout(w_dff_B_qAGUZoC20_2),.clk(gclk));
	jdff dff_B_M8j8a8cD8_2(.din(w_dff_B_qAGUZoC20_2),.dout(w_dff_B_M8j8a8cD8_2),.clk(gclk));
	jdff dff_B_6vxfeEe18_2(.din(w_dff_B_M8j8a8cD8_2),.dout(w_dff_B_6vxfeEe18_2),.clk(gclk));
	jdff dff_B_HnYbGdPz3_2(.din(w_dff_B_6vxfeEe18_2),.dout(w_dff_B_HnYbGdPz3_2),.clk(gclk));
	jdff dff_B_rMASGJuo7_2(.din(w_dff_B_HnYbGdPz3_2),.dout(w_dff_B_rMASGJuo7_2),.clk(gclk));
	jdff dff_B_qFvWF0m06_2(.din(w_dff_B_rMASGJuo7_2),.dout(w_dff_B_qFvWF0m06_2),.clk(gclk));
	jdff dff_B_Y2SThVqk4_2(.din(w_dff_B_qFvWF0m06_2),.dout(w_dff_B_Y2SThVqk4_2),.clk(gclk));
	jdff dff_B_xGwlfjck2_2(.din(w_dff_B_Y2SThVqk4_2),.dout(w_dff_B_xGwlfjck2_2),.clk(gclk));
	jdff dff_B_QP6s4kkk8_2(.din(w_dff_B_xGwlfjck2_2),.dout(w_dff_B_QP6s4kkk8_2),.clk(gclk));
	jdff dff_B_5g7jLAsm7_2(.din(w_dff_B_QP6s4kkk8_2),.dout(w_dff_B_5g7jLAsm7_2),.clk(gclk));
	jdff dff_B_djCIo45C6_2(.din(w_dff_B_5g7jLAsm7_2),.dout(w_dff_B_djCIo45C6_2),.clk(gclk));
	jdff dff_B_EiNPJyiw2_2(.din(w_dff_B_djCIo45C6_2),.dout(w_dff_B_EiNPJyiw2_2),.clk(gclk));
	jdff dff_B_5rhA6zGm7_2(.din(w_dff_B_EiNPJyiw2_2),.dout(w_dff_B_5rhA6zGm7_2),.clk(gclk));
	jdff dff_B_AqizxOau4_1(.din(n1348),.dout(w_dff_B_AqizxOau4_1),.clk(gclk));
	jdff dff_B_nz9DrSU60_2(.din(n1262),.dout(w_dff_B_nz9DrSU60_2),.clk(gclk));
	jdff dff_B_ntXv2OJM3_2(.din(w_dff_B_nz9DrSU60_2),.dout(w_dff_B_ntXv2OJM3_2),.clk(gclk));
	jdff dff_B_PG7YBjra7_2(.din(w_dff_B_ntXv2OJM3_2),.dout(w_dff_B_PG7YBjra7_2),.clk(gclk));
	jdff dff_B_5aRFOs3S3_2(.din(w_dff_B_PG7YBjra7_2),.dout(w_dff_B_5aRFOs3S3_2),.clk(gclk));
	jdff dff_B_VoPP6YrR0_2(.din(w_dff_B_5aRFOs3S3_2),.dout(w_dff_B_VoPP6YrR0_2),.clk(gclk));
	jdff dff_B_vEotDmyG3_2(.din(w_dff_B_VoPP6YrR0_2),.dout(w_dff_B_vEotDmyG3_2),.clk(gclk));
	jdff dff_B_Yq6fbw8A8_2(.din(w_dff_B_vEotDmyG3_2),.dout(w_dff_B_Yq6fbw8A8_2),.clk(gclk));
	jdff dff_B_LZG5QkFe4_2(.din(w_dff_B_Yq6fbw8A8_2),.dout(w_dff_B_LZG5QkFe4_2),.clk(gclk));
	jdff dff_B_YLNYEWHh0_2(.din(w_dff_B_LZG5QkFe4_2),.dout(w_dff_B_YLNYEWHh0_2),.clk(gclk));
	jdff dff_B_6ywo4OgW3_2(.din(w_dff_B_YLNYEWHh0_2),.dout(w_dff_B_6ywo4OgW3_2),.clk(gclk));
	jdff dff_B_wsuBI3Td1_2(.din(w_dff_B_6ywo4OgW3_2),.dout(w_dff_B_wsuBI3Td1_2),.clk(gclk));
	jdff dff_B_jt55LJ7J9_2(.din(w_dff_B_wsuBI3Td1_2),.dout(w_dff_B_jt55LJ7J9_2),.clk(gclk));
	jdff dff_B_1vZzD2DW9_2(.din(w_dff_B_jt55LJ7J9_2),.dout(w_dff_B_1vZzD2DW9_2),.clk(gclk));
	jdff dff_B_wxBL12NL9_2(.din(w_dff_B_1vZzD2DW9_2),.dout(w_dff_B_wxBL12NL9_2),.clk(gclk));
	jdff dff_B_Hw4blZWM1_2(.din(w_dff_B_wxBL12NL9_2),.dout(w_dff_B_Hw4blZWM1_2),.clk(gclk));
	jdff dff_B_dS6gl4Jj2_2(.din(w_dff_B_Hw4blZWM1_2),.dout(w_dff_B_dS6gl4Jj2_2),.clk(gclk));
	jdff dff_B_YDaxvvi08_2(.din(w_dff_B_dS6gl4Jj2_2),.dout(w_dff_B_YDaxvvi08_2),.clk(gclk));
	jdff dff_B_PgfjzkDW5_2(.din(n1273),.dout(w_dff_B_PgfjzkDW5_2),.clk(gclk));
	jdff dff_B_w3UW7JaH0_1(.din(n1268),.dout(w_dff_B_w3UW7JaH0_1),.clk(gclk));
	jdff dff_B_DIHpMLGD7_1(.din(w_dff_B_w3UW7JaH0_1),.dout(w_dff_B_DIHpMLGD7_1),.clk(gclk));
	jdff dff_B_S7miAAlE2_2(.din(n1267),.dout(w_dff_B_S7miAAlE2_2),.clk(gclk));
	jdff dff_B_IUVelolb2_2(.din(w_dff_B_S7miAAlE2_2),.dout(w_dff_B_IUVelolb2_2),.clk(gclk));
	jdff dff_B_BtC00bdT3_2(.din(w_dff_B_IUVelolb2_2),.dout(w_dff_B_BtC00bdT3_2),.clk(gclk));
	jdff dff_B_EZgn3QZ04_2(.din(w_dff_B_BtC00bdT3_2),.dout(w_dff_B_EZgn3QZ04_2),.clk(gclk));
	jdff dff_B_eLLo6tPw3_2(.din(w_dff_B_EZgn3QZ04_2),.dout(w_dff_B_eLLo6tPw3_2),.clk(gclk));
	jdff dff_B_24l28blo8_2(.din(w_dff_B_eLLo6tPw3_2),.dout(w_dff_B_24l28blo8_2),.clk(gclk));
	jdff dff_B_nbQo6sYz5_2(.din(w_dff_B_24l28blo8_2),.dout(w_dff_B_nbQo6sYz5_2),.clk(gclk));
	jdff dff_B_vAaQu0rq1_2(.din(w_dff_B_nbQo6sYz5_2),.dout(w_dff_B_vAaQu0rq1_2),.clk(gclk));
	jdff dff_B_ZRGZ9G752_2(.din(w_dff_B_vAaQu0rq1_2),.dout(w_dff_B_ZRGZ9G752_2),.clk(gclk));
	jdff dff_B_siqKQiPV5_2(.din(w_dff_B_ZRGZ9G752_2),.dout(w_dff_B_siqKQiPV5_2),.clk(gclk));
	jdff dff_B_jOZ1XtX40_2(.din(w_dff_B_siqKQiPV5_2),.dout(w_dff_B_jOZ1XtX40_2),.clk(gclk));
	jdff dff_B_kHxt7nel9_2(.din(w_dff_B_jOZ1XtX40_2),.dout(w_dff_B_kHxt7nel9_2),.clk(gclk));
	jdff dff_B_HYsBGq0B0_2(.din(w_dff_B_kHxt7nel9_2),.dout(w_dff_B_HYsBGq0B0_2),.clk(gclk));
	jdff dff_B_tkPmTYjn8_2(.din(n1266),.dout(w_dff_B_tkPmTYjn8_2),.clk(gclk));
	jdff dff_B_BxPtfmVg5_2(.din(w_dff_B_tkPmTYjn8_2),.dout(w_dff_B_BxPtfmVg5_2),.clk(gclk));
	jdff dff_B_XquK6lfj3_2(.din(w_dff_B_BxPtfmVg5_2),.dout(w_dff_B_XquK6lfj3_2),.clk(gclk));
	jdff dff_B_pgm5CIOg2_2(.din(w_dff_B_XquK6lfj3_2),.dout(w_dff_B_pgm5CIOg2_2),.clk(gclk));
	jdff dff_B_q5f0g6KW4_2(.din(w_dff_B_pgm5CIOg2_2),.dout(w_dff_B_q5f0g6KW4_2),.clk(gclk));
	jdff dff_B_JlVxxxPi2_2(.din(w_dff_B_q5f0g6KW4_2),.dout(w_dff_B_JlVxxxPi2_2),.clk(gclk));
	jdff dff_B_GJtcJ5q20_2(.din(w_dff_B_JlVxxxPi2_2),.dout(w_dff_B_GJtcJ5q20_2),.clk(gclk));
	jdff dff_B_BNAFJrX09_2(.din(w_dff_B_GJtcJ5q20_2),.dout(w_dff_B_BNAFJrX09_2),.clk(gclk));
	jdff dff_B_Zaa1qRCy2_2(.din(w_dff_B_BNAFJrX09_2),.dout(w_dff_B_Zaa1qRCy2_2),.clk(gclk));
	jdff dff_B_rpMtXSaV3_2(.din(w_dff_B_Zaa1qRCy2_2),.dout(w_dff_B_rpMtXSaV3_2),.clk(gclk));
	jdff dff_B_GHJChAcJ6_2(.din(w_dff_B_rpMtXSaV3_2),.dout(w_dff_B_GHJChAcJ6_2),.clk(gclk));
	jdff dff_B_WpxNynRH4_2(.din(w_dff_B_GHJChAcJ6_2),.dout(w_dff_B_WpxNynRH4_2),.clk(gclk));
	jdff dff_B_tYLlUs1z0_2(.din(w_dff_B_WpxNynRH4_2),.dout(w_dff_B_tYLlUs1z0_2),.clk(gclk));
	jdff dff_B_Iu5vrsMQ1_2(.din(w_dff_B_tYLlUs1z0_2),.dout(w_dff_B_Iu5vrsMQ1_2),.clk(gclk));
	jdff dff_B_BP1LWsrF9_2(.din(w_dff_B_Iu5vrsMQ1_2),.dout(w_dff_B_BP1LWsrF9_2),.clk(gclk));
	jdff dff_B_aeNosS844_1(.din(n1263),.dout(w_dff_B_aeNosS844_1),.clk(gclk));
	jdff dff_B_gz4ugIcs0_2(.din(n1171),.dout(w_dff_B_gz4ugIcs0_2),.clk(gclk));
	jdff dff_B_0ZlW6rUd3_2(.din(w_dff_B_gz4ugIcs0_2),.dout(w_dff_B_0ZlW6rUd3_2),.clk(gclk));
	jdff dff_B_iij9tUrU4_2(.din(w_dff_B_0ZlW6rUd3_2),.dout(w_dff_B_iij9tUrU4_2),.clk(gclk));
	jdff dff_B_4vgmQj8H5_2(.din(w_dff_B_iij9tUrU4_2),.dout(w_dff_B_4vgmQj8H5_2),.clk(gclk));
	jdff dff_B_zejx364E6_2(.din(w_dff_B_4vgmQj8H5_2),.dout(w_dff_B_zejx364E6_2),.clk(gclk));
	jdff dff_B_mLmBGkIA4_2(.din(w_dff_B_zejx364E6_2),.dout(w_dff_B_mLmBGkIA4_2),.clk(gclk));
	jdff dff_B_oY9Nxm7D8_2(.din(w_dff_B_mLmBGkIA4_2),.dout(w_dff_B_oY9Nxm7D8_2),.clk(gclk));
	jdff dff_B_gK4EYb8k8_2(.din(w_dff_B_oY9Nxm7D8_2),.dout(w_dff_B_gK4EYb8k8_2),.clk(gclk));
	jdff dff_B_vpbQY6bd2_2(.din(w_dff_B_gK4EYb8k8_2),.dout(w_dff_B_vpbQY6bd2_2),.clk(gclk));
	jdff dff_B_ruSHOu9E3_2(.din(w_dff_B_vpbQY6bd2_2),.dout(w_dff_B_ruSHOu9E3_2),.clk(gclk));
	jdff dff_B_PMHAVfwd9_2(.din(w_dff_B_ruSHOu9E3_2),.dout(w_dff_B_PMHAVfwd9_2),.clk(gclk));
	jdff dff_B_LU2xYyHE0_2(.din(w_dff_B_PMHAVfwd9_2),.dout(w_dff_B_LU2xYyHE0_2),.clk(gclk));
	jdff dff_B_u6FExlep8_2(.din(w_dff_B_LU2xYyHE0_2),.dout(w_dff_B_u6FExlep8_2),.clk(gclk));
	jdff dff_B_DnRcI9J06_2(.din(w_dff_B_u6FExlep8_2),.dout(w_dff_B_DnRcI9J06_2),.clk(gclk));
	jdff dff_B_vLBFI7kX2_2(.din(n1182),.dout(w_dff_B_vLBFI7kX2_2),.clk(gclk));
	jdff dff_B_OJa5jAA83_2(.din(w_dff_B_vLBFI7kX2_2),.dout(w_dff_B_OJa5jAA83_2),.clk(gclk));
	jdff dff_B_OFzGlZfO7_1(.din(n1177),.dout(w_dff_B_OFzGlZfO7_1),.clk(gclk));
	jdff dff_B_SD9sF0Cs1_1(.din(w_dff_B_OFzGlZfO7_1),.dout(w_dff_B_SD9sF0Cs1_1),.clk(gclk));
	jdff dff_B_QaLurC0e0_2(.din(n1176),.dout(w_dff_B_QaLurC0e0_2),.clk(gclk));
	jdff dff_B_bpSmEV1q8_2(.din(w_dff_B_QaLurC0e0_2),.dout(w_dff_B_bpSmEV1q8_2),.clk(gclk));
	jdff dff_B_J7EFGDsQ1_2(.din(w_dff_B_bpSmEV1q8_2),.dout(w_dff_B_J7EFGDsQ1_2),.clk(gclk));
	jdff dff_B_OX3vOu7t7_2(.din(w_dff_B_J7EFGDsQ1_2),.dout(w_dff_B_OX3vOu7t7_2),.clk(gclk));
	jdff dff_B_7bXp8v1W7_2(.din(w_dff_B_OX3vOu7t7_2),.dout(w_dff_B_7bXp8v1W7_2),.clk(gclk));
	jdff dff_B_37Ba0chz7_2(.din(w_dff_B_7bXp8v1W7_2),.dout(w_dff_B_37Ba0chz7_2),.clk(gclk));
	jdff dff_B_2KlZSCcS2_2(.din(w_dff_B_37Ba0chz7_2),.dout(w_dff_B_2KlZSCcS2_2),.clk(gclk));
	jdff dff_B_TbL9iLmj7_2(.din(w_dff_B_2KlZSCcS2_2),.dout(w_dff_B_TbL9iLmj7_2),.clk(gclk));
	jdff dff_B_0k8pGfeg4_2(.din(w_dff_B_TbL9iLmj7_2),.dout(w_dff_B_0k8pGfeg4_2),.clk(gclk));
	jdff dff_B_mPD3MaaR6_2(.din(n1175),.dout(w_dff_B_mPD3MaaR6_2),.clk(gclk));
	jdff dff_B_HvS5g1lJ0_2(.din(w_dff_B_mPD3MaaR6_2),.dout(w_dff_B_HvS5g1lJ0_2),.clk(gclk));
	jdff dff_B_7IvXLYJf4_2(.din(w_dff_B_HvS5g1lJ0_2),.dout(w_dff_B_7IvXLYJf4_2),.clk(gclk));
	jdff dff_B_APs3vc0s8_2(.din(w_dff_B_7IvXLYJf4_2),.dout(w_dff_B_APs3vc0s8_2),.clk(gclk));
	jdff dff_B_CIjp0FNg9_2(.din(w_dff_B_APs3vc0s8_2),.dout(w_dff_B_CIjp0FNg9_2),.clk(gclk));
	jdff dff_B_yr5QtQdn2_2(.din(w_dff_B_CIjp0FNg9_2),.dout(w_dff_B_yr5QtQdn2_2),.clk(gclk));
	jdff dff_B_ucHTXldm6_2(.din(w_dff_B_yr5QtQdn2_2),.dout(w_dff_B_ucHTXldm6_2),.clk(gclk));
	jdff dff_B_R6DVXZaE2_2(.din(w_dff_B_ucHTXldm6_2),.dout(w_dff_B_R6DVXZaE2_2),.clk(gclk));
	jdff dff_B_qGvxvP9i8_2(.din(w_dff_B_R6DVXZaE2_2),.dout(w_dff_B_qGvxvP9i8_2),.clk(gclk));
	jdff dff_B_QVDCbL2V2_2(.din(w_dff_B_qGvxvP9i8_2),.dout(w_dff_B_QVDCbL2V2_2),.clk(gclk));
	jdff dff_B_VjTNHORE0_2(.din(w_dff_B_QVDCbL2V2_2),.dout(w_dff_B_VjTNHORE0_2),.clk(gclk));
	jdff dff_B_5fzawKms6_1(.din(n1172),.dout(w_dff_B_5fzawKms6_1),.clk(gclk));
	jdff dff_B_wsTcT6Du0_2(.din(n1073),.dout(w_dff_B_wsTcT6Du0_2),.clk(gclk));
	jdff dff_B_7r0mPeHX4_2(.din(w_dff_B_wsTcT6Du0_2),.dout(w_dff_B_7r0mPeHX4_2),.clk(gclk));
	jdff dff_B_N2I7r5sW2_2(.din(w_dff_B_7r0mPeHX4_2),.dout(w_dff_B_N2I7r5sW2_2),.clk(gclk));
	jdff dff_B_UF2C35uT0_2(.din(w_dff_B_N2I7r5sW2_2),.dout(w_dff_B_UF2C35uT0_2),.clk(gclk));
	jdff dff_B_aCqy50DP1_2(.din(w_dff_B_UF2C35uT0_2),.dout(w_dff_B_aCqy50DP1_2),.clk(gclk));
	jdff dff_B_JOJvbckc7_2(.din(w_dff_B_aCqy50DP1_2),.dout(w_dff_B_JOJvbckc7_2),.clk(gclk));
	jdff dff_B_pdwwQ1TC8_2(.din(w_dff_B_JOJvbckc7_2),.dout(w_dff_B_pdwwQ1TC8_2),.clk(gclk));
	jdff dff_B_gN1PgTyV2_2(.din(w_dff_B_pdwwQ1TC8_2),.dout(w_dff_B_gN1PgTyV2_2),.clk(gclk));
	jdff dff_B_LoTTiBbr1_2(.din(w_dff_B_gN1PgTyV2_2),.dout(w_dff_B_LoTTiBbr1_2),.clk(gclk));
	jdff dff_B_lBt4bscN8_2(.din(w_dff_B_LoTTiBbr1_2),.dout(w_dff_B_lBt4bscN8_2),.clk(gclk));
	jdff dff_B_dsSb6e5W5_2(.din(w_dff_B_lBt4bscN8_2),.dout(w_dff_B_dsSb6e5W5_2),.clk(gclk));
	jdff dff_B_1KLaqIJr5_2(.din(n1083),.dout(w_dff_B_1KLaqIJr5_2),.clk(gclk));
	jdff dff_B_RbHQ6WDG5_2(.din(w_dff_B_1KLaqIJr5_2),.dout(w_dff_B_RbHQ6WDG5_2),.clk(gclk));
	jdff dff_B_gbsWdu792_2(.din(w_dff_B_RbHQ6WDG5_2),.dout(w_dff_B_gbsWdu792_2),.clk(gclk));
	jdff dff_B_xBcfH5Hk6_2(.din(n1078),.dout(w_dff_B_xBcfH5Hk6_2),.clk(gclk));
	jdff dff_B_SmC5t9hb1_2(.din(w_dff_B_xBcfH5Hk6_2),.dout(w_dff_B_SmC5t9hb1_2),.clk(gclk));
	jdff dff_B_VHvBBpfl8_2(.din(w_dff_B_SmC5t9hb1_2),.dout(w_dff_B_VHvBBpfl8_2),.clk(gclk));
	jdff dff_B_k7SHEqls8_2(.din(w_dff_B_VHvBBpfl8_2),.dout(w_dff_B_k7SHEqls8_2),.clk(gclk));
	jdff dff_B_PJgaHfRU1_2(.din(w_dff_B_k7SHEqls8_2),.dout(w_dff_B_PJgaHfRU1_2),.clk(gclk));
	jdff dff_B_NO34ytKQ1_2(.din(n1077),.dout(w_dff_B_NO34ytKQ1_2),.clk(gclk));
	jdff dff_B_UIoTEzfY3_2(.din(w_dff_B_NO34ytKQ1_2),.dout(w_dff_B_UIoTEzfY3_2),.clk(gclk));
	jdff dff_B_Hs3Qj9xI6_2(.din(w_dff_B_UIoTEzfY3_2),.dout(w_dff_B_Hs3Qj9xI6_2),.clk(gclk));
	jdff dff_B_dj0bbnkz3_2(.din(w_dff_B_Hs3Qj9xI6_2),.dout(w_dff_B_dj0bbnkz3_2),.clk(gclk));
	jdff dff_B_w1LqP5Ba0_2(.din(w_dff_B_dj0bbnkz3_2),.dout(w_dff_B_w1LqP5Ba0_2),.clk(gclk));
	jdff dff_B_9AOZzDh31_2(.din(w_dff_B_w1LqP5Ba0_2),.dout(w_dff_B_9AOZzDh31_2),.clk(gclk));
	jdff dff_B_nWASdzTi0_2(.din(w_dff_B_9AOZzDh31_2),.dout(w_dff_B_nWASdzTi0_2),.clk(gclk));
	jdff dff_B_Kvu2NZ8E1_1(.din(n1074),.dout(w_dff_B_Kvu2NZ8E1_1),.clk(gclk));
	jdff dff_B_b7VkWaVq0_2(.din(n974),.dout(w_dff_B_b7VkWaVq0_2),.clk(gclk));
	jdff dff_B_mkivJK7r1_2(.din(w_dff_B_b7VkWaVq0_2),.dout(w_dff_B_mkivJK7r1_2),.clk(gclk));
	jdff dff_B_VUMyWcSP6_2(.din(w_dff_B_mkivJK7r1_2),.dout(w_dff_B_VUMyWcSP6_2),.clk(gclk));
	jdff dff_B_5JAcsR253_2(.din(w_dff_B_VUMyWcSP6_2),.dout(w_dff_B_5JAcsR253_2),.clk(gclk));
	jdff dff_B_jomUdwLt9_2(.din(w_dff_B_5JAcsR253_2),.dout(w_dff_B_jomUdwLt9_2),.clk(gclk));
	jdff dff_B_XFWsS37N1_2(.din(w_dff_B_jomUdwLt9_2),.dout(w_dff_B_XFWsS37N1_2),.clk(gclk));
	jdff dff_B_WfJUC5Th7_2(.din(w_dff_B_XFWsS37N1_2),.dout(w_dff_B_WfJUC5Th7_2),.clk(gclk));
	jdff dff_B_rHluWfOf0_2(.din(w_dff_B_WfJUC5Th7_2),.dout(w_dff_B_rHluWfOf0_2),.clk(gclk));
	jdff dff_B_PuzwdCvi4_2(.din(n984),.dout(w_dff_B_PuzwdCvi4_2),.clk(gclk));
	jdff dff_B_pUoWxrfk5_2(.din(w_dff_B_PuzwdCvi4_2),.dout(w_dff_B_pUoWxrfk5_2),.clk(gclk));
	jdff dff_B_P1VSDqeu3_2(.din(w_dff_B_pUoWxrfk5_2),.dout(w_dff_B_P1VSDqeu3_2),.clk(gclk));
	jdff dff_B_uSkMMjTT2_2(.din(w_dff_B_P1VSDqeu3_2),.dout(w_dff_B_uSkMMjTT2_2),.clk(gclk));
	jdff dff_B_zSwb67hh5_2(.din(n983),.dout(w_dff_B_zSwb67hh5_2),.clk(gclk));
	jdff dff_B_4QMQO2HH8_2(.din(w_dff_B_zSwb67hh5_2),.dout(w_dff_B_4QMQO2HH8_2),.clk(gclk));
	jdff dff_B_lQTeKuBM6_2(.din(w_dff_B_4QMQO2HH8_2),.dout(w_dff_B_lQTeKuBM6_2),.clk(gclk));
	jdff dff_A_FudOx7h20_0(.dout(w_n980_0[0]),.din(w_dff_A_FudOx7h20_0),.clk(gclk));
	jdff dff_A_4HSIEWTC5_0(.dout(w_dff_A_FudOx7h20_0),.din(w_dff_A_4HSIEWTC5_0),.clk(gclk));
	jdff dff_A_CQ0L2kB03_0(.dout(w_dff_A_4HSIEWTC5_0),.din(w_dff_A_CQ0L2kB03_0),.clk(gclk));
	jdff dff_B_pWjCZ7xu6_2(.din(n980),.dout(w_dff_B_pWjCZ7xu6_2),.clk(gclk));
	jdff dff_A_UzGkmPuH7_0(.dout(w_n877_0[0]),.din(w_dff_A_UzGkmPuH7_0),.clk(gclk));
	jdff dff_A_MSQpi08P7_0(.dout(w_dff_A_UzGkmPuH7_0),.din(w_dff_A_MSQpi08P7_0),.clk(gclk));
	jdff dff_A_kM3WLGk62_0(.dout(w_dff_A_MSQpi08P7_0),.din(w_dff_A_kM3WLGk62_0),.clk(gclk));
	jdff dff_B_4DEEQ4gN5_2(.din(n877),.dout(w_dff_B_4DEEQ4gN5_2),.clk(gclk));
	jdff dff_A_cIGZ47B76_0(.dout(w_n875_0[0]),.din(w_dff_A_cIGZ47B76_0),.clk(gclk));
	jdff dff_A_ZGZ8rWrU5_0(.dout(w_dff_A_cIGZ47B76_0),.din(w_dff_A_ZGZ8rWrU5_0),.clk(gclk));
	jdff dff_B_rJjPETkF3_2(.din(n874),.dout(w_dff_B_rJjPETkF3_2),.clk(gclk));
	jdff dff_B_iwILiT0Z8_2(.din(w_dff_B_rJjPETkF3_2),.dout(w_dff_B_iwILiT0Z8_2),.clk(gclk));
	jdff dff_B_6xdhJ48v5_2(.din(w_dff_B_iwILiT0Z8_2),.dout(w_dff_B_6xdhJ48v5_2),.clk(gclk));
	jdff dff_A_SBHDbXIx1_1(.dout(w_dff_A_4gQ9ZUKu3_0),.din(w_dff_A_SBHDbXIx1_1),.clk(gclk));
	jdff dff_A_4gQ9ZUKu3_0(.dout(w_dff_A_pPQigq9M5_0),.din(w_dff_A_4gQ9ZUKu3_0),.clk(gclk));
	jdff dff_A_pPQigq9M5_0(.dout(w_dff_A_eI17mUKL4_0),.din(w_dff_A_pPQigq9M5_0),.clk(gclk));
	jdff dff_A_eI17mUKL4_0(.dout(w_dff_A_PdpyK4ry0_0),.din(w_dff_A_eI17mUKL4_0),.clk(gclk));
	jdff dff_A_PdpyK4ry0_0(.dout(w_dff_A_LljHSyni0_0),.din(w_dff_A_PdpyK4ry0_0),.clk(gclk));
	jdff dff_A_LljHSyni0_0(.dout(w_dff_A_YeHL9aIy8_0),.din(w_dff_A_LljHSyni0_0),.clk(gclk));
	jdff dff_A_YeHL9aIy8_0(.dout(w_dff_A_7Y8JO7ZJ2_0),.din(w_dff_A_YeHL9aIy8_0),.clk(gclk));
	jdff dff_A_7Y8JO7ZJ2_0(.dout(w_dff_A_iPlPA2Ip5_0),.din(w_dff_A_7Y8JO7ZJ2_0),.clk(gclk));
	jdff dff_A_iPlPA2Ip5_0(.dout(w_dff_A_zo0549vH2_0),.din(w_dff_A_iPlPA2Ip5_0),.clk(gclk));
	jdff dff_A_zo0549vH2_0(.dout(w_dff_A_QYQci1fk0_0),.din(w_dff_A_zo0549vH2_0),.clk(gclk));
	jdff dff_A_QYQci1fk0_0(.dout(w_dff_A_OiAZEN2v0_0),.din(w_dff_A_QYQci1fk0_0),.clk(gclk));
	jdff dff_A_OiAZEN2v0_0(.dout(w_dff_A_vDxG6o7n8_0),.din(w_dff_A_OiAZEN2v0_0),.clk(gclk));
	jdff dff_A_vDxG6o7n8_0(.dout(w_dff_A_kBEVpuim4_0),.din(w_dff_A_vDxG6o7n8_0),.clk(gclk));
	jdff dff_A_kBEVpuim4_0(.dout(w_dff_A_nhrO4Cok2_0),.din(w_dff_A_kBEVpuim4_0),.clk(gclk));
	jdff dff_A_nhrO4Cok2_0(.dout(w_dff_A_IcvCZ8672_0),.din(w_dff_A_nhrO4Cok2_0),.clk(gclk));
	jdff dff_A_IcvCZ8672_0(.dout(w_dff_A_tltlAlJX5_0),.din(w_dff_A_IcvCZ8672_0),.clk(gclk));
	jdff dff_A_tltlAlJX5_0(.dout(w_dff_A_8G0ZVXKd4_0),.din(w_dff_A_tltlAlJX5_0),.clk(gclk));
	jdff dff_A_8G0ZVXKd4_0(.dout(w_dff_A_vb3okClZ5_0),.din(w_dff_A_8G0ZVXKd4_0),.clk(gclk));
	jdff dff_A_vb3okClZ5_0(.dout(w_dff_A_vQku3r5r0_0),.din(w_dff_A_vb3okClZ5_0),.clk(gclk));
	jdff dff_A_vQku3r5r0_0(.dout(w_dff_A_8rg70ohz8_0),.din(w_dff_A_vQku3r5r0_0),.clk(gclk));
	jdff dff_A_8rg70ohz8_0(.dout(w_dff_A_3n7Q4p9d4_0),.din(w_dff_A_8rg70ohz8_0),.clk(gclk));
	jdff dff_A_3n7Q4p9d4_0(.dout(w_dff_A_y7Vu8jfj0_0),.din(w_dff_A_3n7Q4p9d4_0),.clk(gclk));
	jdff dff_A_y7Vu8jfj0_0(.dout(w_dff_A_9Eor3Hjo5_0),.din(w_dff_A_y7Vu8jfj0_0),.clk(gclk));
	jdff dff_A_9Eor3Hjo5_0(.dout(w_dff_A_1otuXqZt4_0),.din(w_dff_A_9Eor3Hjo5_0),.clk(gclk));
	jdff dff_A_1otuXqZt4_0(.dout(w_dff_A_6VIoMdNo0_0),.din(w_dff_A_1otuXqZt4_0),.clk(gclk));
	jdff dff_A_6VIoMdNo0_0(.dout(w_dff_A_xhkOA6d50_0),.din(w_dff_A_6VIoMdNo0_0),.clk(gclk));
	jdff dff_A_xhkOA6d50_0(.dout(w_dff_A_OlotAoqD8_0),.din(w_dff_A_xhkOA6d50_0),.clk(gclk));
	jdff dff_A_OlotAoqD8_0(.dout(w_dff_A_Fj4mPkYJ5_0),.din(w_dff_A_OlotAoqD8_0),.clk(gclk));
	jdff dff_A_Fj4mPkYJ5_0(.dout(w_dff_A_dd4IHaLo4_0),.din(w_dff_A_Fj4mPkYJ5_0),.clk(gclk));
	jdff dff_A_dd4IHaLo4_0(.dout(w_dff_A_vttlEuDG3_0),.din(w_dff_A_dd4IHaLo4_0),.clk(gclk));
	jdff dff_A_vttlEuDG3_0(.dout(w_dff_A_XFPGfoyo9_0),.din(w_dff_A_vttlEuDG3_0),.clk(gclk));
	jdff dff_A_XFPGfoyo9_0(.dout(w_dff_A_0GuCBN7h6_0),.din(w_dff_A_XFPGfoyo9_0),.clk(gclk));
	jdff dff_A_0GuCBN7h6_0(.dout(w_dff_A_fzMSTGnW4_0),.din(w_dff_A_0GuCBN7h6_0),.clk(gclk));
	jdff dff_A_fzMSTGnW4_0(.dout(w_dff_A_Lq5pI89p4_0),.din(w_dff_A_fzMSTGnW4_0),.clk(gclk));
	jdff dff_A_Lq5pI89p4_0(.dout(w_dff_A_3aywD2BY3_0),.din(w_dff_A_Lq5pI89p4_0),.clk(gclk));
	jdff dff_A_3aywD2BY3_0(.dout(w_dff_A_BvpnkpUv4_0),.din(w_dff_A_3aywD2BY3_0),.clk(gclk));
	jdff dff_A_BvpnkpUv4_0(.dout(w_dff_A_p8qqB4hC7_0),.din(w_dff_A_BvpnkpUv4_0),.clk(gclk));
	jdff dff_A_p8qqB4hC7_0(.dout(w_dff_A_MWZThVTg6_0),.din(w_dff_A_p8qqB4hC7_0),.clk(gclk));
	jdff dff_A_MWZThVTg6_0(.dout(w_dff_A_OW6khchs0_0),.din(w_dff_A_MWZThVTg6_0),.clk(gclk));
	jdff dff_A_OW6khchs0_0(.dout(w_dff_A_LD4LPZq52_0),.din(w_dff_A_OW6khchs0_0),.clk(gclk));
	jdff dff_A_LD4LPZq52_0(.dout(w_dff_A_u9QVAb9v2_0),.din(w_dff_A_LD4LPZq52_0),.clk(gclk));
	jdff dff_A_u9QVAb9v2_0(.dout(w_dff_A_JoN3L7Ym8_0),.din(w_dff_A_u9QVAb9v2_0),.clk(gclk));
	jdff dff_A_JoN3L7Ym8_0(.dout(w_dff_A_wn67Koel0_0),.din(w_dff_A_JoN3L7Ym8_0),.clk(gclk));
	jdff dff_A_wn67Koel0_0(.dout(w_dff_A_80IDQ1SK6_0),.din(w_dff_A_wn67Koel0_0),.clk(gclk));
	jdff dff_A_80IDQ1SK6_0(.dout(w_dff_A_lJavKu555_0),.din(w_dff_A_80IDQ1SK6_0),.clk(gclk));
	jdff dff_A_lJavKu555_0(.dout(w_dff_A_IhD23cpZ7_0),.din(w_dff_A_lJavKu555_0),.clk(gclk));
	jdff dff_A_IhD23cpZ7_0(.dout(w_dff_A_GkZLiVdJ6_0),.din(w_dff_A_IhD23cpZ7_0),.clk(gclk));
	jdff dff_A_GkZLiVdJ6_0(.dout(w_dff_A_PJj3rKIH7_0),.din(w_dff_A_GkZLiVdJ6_0),.clk(gclk));
	jdff dff_A_PJj3rKIH7_0(.dout(w_dff_A_0vxVuywM2_0),.din(w_dff_A_PJj3rKIH7_0),.clk(gclk));
	jdff dff_A_0vxVuywM2_0(.dout(w_dff_A_IsojOi9V4_0),.din(w_dff_A_0vxVuywM2_0),.clk(gclk));
	jdff dff_A_IsojOi9V4_0(.dout(w_dff_A_RBtRBIYw7_0),.din(w_dff_A_IsojOi9V4_0),.clk(gclk));
	jdff dff_A_RBtRBIYw7_0(.dout(w_dff_A_DxGRfkrQ7_0),.din(w_dff_A_RBtRBIYw7_0),.clk(gclk));
	jdff dff_A_DxGRfkrQ7_0(.dout(w_dff_A_er8aXkTg5_0),.din(w_dff_A_DxGRfkrQ7_0),.clk(gclk));
	jdff dff_A_er8aXkTg5_0(.dout(w_dff_A_6ntCjEA50_0),.din(w_dff_A_er8aXkTg5_0),.clk(gclk));
	jdff dff_A_6ntCjEA50_0(.dout(w_dff_A_WxxUDhz89_0),.din(w_dff_A_6ntCjEA50_0),.clk(gclk));
	jdff dff_A_WxxUDhz89_0(.dout(w_dff_A_AsbJXWKL8_0),.din(w_dff_A_WxxUDhz89_0),.clk(gclk));
	jdff dff_A_AsbJXWKL8_0(.dout(w_dff_A_xIqktCFN7_0),.din(w_dff_A_AsbJXWKL8_0),.clk(gclk));
	jdff dff_A_xIqktCFN7_0(.dout(w_dff_A_MKLHHGtO8_0),.din(w_dff_A_xIqktCFN7_0),.clk(gclk));
	jdff dff_A_MKLHHGtO8_0(.dout(w_dff_A_15MuG5kP2_0),.din(w_dff_A_MKLHHGtO8_0),.clk(gclk));
	jdff dff_A_15MuG5kP2_0(.dout(w_dff_A_oOvTVNbi6_0),.din(w_dff_A_15MuG5kP2_0),.clk(gclk));
	jdff dff_A_oOvTVNbi6_0(.dout(w_dff_A_y0Lfbng75_0),.din(w_dff_A_oOvTVNbi6_0),.clk(gclk));
	jdff dff_A_y0Lfbng75_0(.dout(w_dff_A_pw8NBRHb1_0),.din(w_dff_A_y0Lfbng75_0),.clk(gclk));
	jdff dff_A_pw8NBRHb1_0(.dout(w_dff_A_h5p1L6Im0_0),.din(w_dff_A_pw8NBRHb1_0),.clk(gclk));
	jdff dff_A_h5p1L6Im0_0(.dout(w_dff_A_SXdZkzCK8_0),.din(w_dff_A_h5p1L6Im0_0),.clk(gclk));
	jdff dff_A_SXdZkzCK8_0(.dout(w_dff_A_WHkIXC9S7_0),.din(w_dff_A_SXdZkzCK8_0),.clk(gclk));
	jdff dff_A_WHkIXC9S7_0(.dout(w_dff_A_PRlghX754_0),.din(w_dff_A_WHkIXC9S7_0),.clk(gclk));
	jdff dff_A_PRlghX754_0(.dout(w_dff_A_890P4iKA2_0),.din(w_dff_A_PRlghX754_0),.clk(gclk));
	jdff dff_A_890P4iKA2_0(.dout(w_dff_A_rDYz4CU07_0),.din(w_dff_A_890P4iKA2_0),.clk(gclk));
	jdff dff_A_rDYz4CU07_0(.dout(w_dff_A_5GQGx5pO5_0),.din(w_dff_A_rDYz4CU07_0),.clk(gclk));
	jdff dff_A_5GQGx5pO5_0(.dout(w_dff_A_ooBTxhM42_0),.din(w_dff_A_5GQGx5pO5_0),.clk(gclk));
	jdff dff_A_ooBTxhM42_0(.dout(w_dff_A_ohbgeCYa9_0),.din(w_dff_A_ooBTxhM42_0),.clk(gclk));
	jdff dff_A_ohbgeCYa9_0(.dout(w_dff_A_JVsAVccg2_0),.din(w_dff_A_ohbgeCYa9_0),.clk(gclk));
	jdff dff_A_JVsAVccg2_0(.dout(w_dff_A_tJS67BLc6_0),.din(w_dff_A_JVsAVccg2_0),.clk(gclk));
	jdff dff_A_tJS67BLc6_0(.dout(G545gat),.din(w_dff_A_tJS67BLc6_0),.clk(gclk));
	jdff dff_A_TXpAQk9U3_2(.dout(w_dff_A_vRJlwoKH4_0),.din(w_dff_A_TXpAQk9U3_2),.clk(gclk));
	jdff dff_A_vRJlwoKH4_0(.dout(w_dff_A_C73LlL5J4_0),.din(w_dff_A_vRJlwoKH4_0),.clk(gclk));
	jdff dff_A_C73LlL5J4_0(.dout(w_dff_A_yFw1wAaJ8_0),.din(w_dff_A_C73LlL5J4_0),.clk(gclk));
	jdff dff_A_yFw1wAaJ8_0(.dout(w_dff_A_rw9zDxdR1_0),.din(w_dff_A_yFw1wAaJ8_0),.clk(gclk));
	jdff dff_A_rw9zDxdR1_0(.dout(w_dff_A_6hyZpext7_0),.din(w_dff_A_rw9zDxdR1_0),.clk(gclk));
	jdff dff_A_6hyZpext7_0(.dout(w_dff_A_Sbe3YF118_0),.din(w_dff_A_6hyZpext7_0),.clk(gclk));
	jdff dff_A_Sbe3YF118_0(.dout(w_dff_A_KQCOlCla5_0),.din(w_dff_A_Sbe3YF118_0),.clk(gclk));
	jdff dff_A_KQCOlCla5_0(.dout(w_dff_A_2TrdDXiy6_0),.din(w_dff_A_KQCOlCla5_0),.clk(gclk));
	jdff dff_A_2TrdDXiy6_0(.dout(w_dff_A_NWvETIUF0_0),.din(w_dff_A_2TrdDXiy6_0),.clk(gclk));
	jdff dff_A_NWvETIUF0_0(.dout(w_dff_A_T1wKX3wU2_0),.din(w_dff_A_NWvETIUF0_0),.clk(gclk));
	jdff dff_A_T1wKX3wU2_0(.dout(w_dff_A_NAQK3TVa0_0),.din(w_dff_A_T1wKX3wU2_0),.clk(gclk));
	jdff dff_A_NAQK3TVa0_0(.dout(w_dff_A_cszTkADn4_0),.din(w_dff_A_NAQK3TVa0_0),.clk(gclk));
	jdff dff_A_cszTkADn4_0(.dout(w_dff_A_unkegTzu8_0),.din(w_dff_A_cszTkADn4_0),.clk(gclk));
	jdff dff_A_unkegTzu8_0(.dout(w_dff_A_jSaQJkPg7_0),.din(w_dff_A_unkegTzu8_0),.clk(gclk));
	jdff dff_A_jSaQJkPg7_0(.dout(w_dff_A_tew7kQNq2_0),.din(w_dff_A_jSaQJkPg7_0),.clk(gclk));
	jdff dff_A_tew7kQNq2_0(.dout(w_dff_A_7HqJiyOl4_0),.din(w_dff_A_tew7kQNq2_0),.clk(gclk));
	jdff dff_A_7HqJiyOl4_0(.dout(w_dff_A_ZwjQEB1m5_0),.din(w_dff_A_7HqJiyOl4_0),.clk(gclk));
	jdff dff_A_ZwjQEB1m5_0(.dout(w_dff_A_ke1r9i094_0),.din(w_dff_A_ZwjQEB1m5_0),.clk(gclk));
	jdff dff_A_ke1r9i094_0(.dout(w_dff_A_csbgERdT2_0),.din(w_dff_A_ke1r9i094_0),.clk(gclk));
	jdff dff_A_csbgERdT2_0(.dout(w_dff_A_Evb8SzQx3_0),.din(w_dff_A_csbgERdT2_0),.clk(gclk));
	jdff dff_A_Evb8SzQx3_0(.dout(w_dff_A_F6cmjWKV8_0),.din(w_dff_A_Evb8SzQx3_0),.clk(gclk));
	jdff dff_A_F6cmjWKV8_0(.dout(w_dff_A_AiXJQjp85_0),.din(w_dff_A_F6cmjWKV8_0),.clk(gclk));
	jdff dff_A_AiXJQjp85_0(.dout(w_dff_A_tuzudz8Y8_0),.din(w_dff_A_AiXJQjp85_0),.clk(gclk));
	jdff dff_A_tuzudz8Y8_0(.dout(w_dff_A_0ExLSiUF7_0),.din(w_dff_A_tuzudz8Y8_0),.clk(gclk));
	jdff dff_A_0ExLSiUF7_0(.dout(w_dff_A_P4W3ewrv5_0),.din(w_dff_A_0ExLSiUF7_0),.clk(gclk));
	jdff dff_A_P4W3ewrv5_0(.dout(w_dff_A_HJyifzUq5_0),.din(w_dff_A_P4W3ewrv5_0),.clk(gclk));
	jdff dff_A_HJyifzUq5_0(.dout(w_dff_A_GtoYfMj76_0),.din(w_dff_A_HJyifzUq5_0),.clk(gclk));
	jdff dff_A_GtoYfMj76_0(.dout(w_dff_A_V3EB6ZcX4_0),.din(w_dff_A_GtoYfMj76_0),.clk(gclk));
	jdff dff_A_V3EB6ZcX4_0(.dout(w_dff_A_W1dEsIh73_0),.din(w_dff_A_V3EB6ZcX4_0),.clk(gclk));
	jdff dff_A_W1dEsIh73_0(.dout(w_dff_A_CkV3fprj9_0),.din(w_dff_A_W1dEsIh73_0),.clk(gclk));
	jdff dff_A_CkV3fprj9_0(.dout(w_dff_A_20HUvyKL2_0),.din(w_dff_A_CkV3fprj9_0),.clk(gclk));
	jdff dff_A_20HUvyKL2_0(.dout(w_dff_A_htP9gWyX3_0),.din(w_dff_A_20HUvyKL2_0),.clk(gclk));
	jdff dff_A_htP9gWyX3_0(.dout(w_dff_A_PhEvehmV8_0),.din(w_dff_A_htP9gWyX3_0),.clk(gclk));
	jdff dff_A_PhEvehmV8_0(.dout(w_dff_A_sMZeNh7a9_0),.din(w_dff_A_PhEvehmV8_0),.clk(gclk));
	jdff dff_A_sMZeNh7a9_0(.dout(w_dff_A_Fv68ae0f3_0),.din(w_dff_A_sMZeNh7a9_0),.clk(gclk));
	jdff dff_A_Fv68ae0f3_0(.dout(w_dff_A_D6UvXoZM2_0),.din(w_dff_A_Fv68ae0f3_0),.clk(gclk));
	jdff dff_A_D6UvXoZM2_0(.dout(w_dff_A_1EVHpBAP4_0),.din(w_dff_A_D6UvXoZM2_0),.clk(gclk));
	jdff dff_A_1EVHpBAP4_0(.dout(w_dff_A_mniHZ3B98_0),.din(w_dff_A_1EVHpBAP4_0),.clk(gclk));
	jdff dff_A_mniHZ3B98_0(.dout(w_dff_A_Eb114fix2_0),.din(w_dff_A_mniHZ3B98_0),.clk(gclk));
	jdff dff_A_Eb114fix2_0(.dout(w_dff_A_K5RERxYj4_0),.din(w_dff_A_Eb114fix2_0),.clk(gclk));
	jdff dff_A_K5RERxYj4_0(.dout(w_dff_A_KUtIuPcF4_0),.din(w_dff_A_K5RERxYj4_0),.clk(gclk));
	jdff dff_A_KUtIuPcF4_0(.dout(w_dff_A_RS0rcUYA9_0),.din(w_dff_A_KUtIuPcF4_0),.clk(gclk));
	jdff dff_A_RS0rcUYA9_0(.dout(w_dff_A_lAIycoQE7_0),.din(w_dff_A_RS0rcUYA9_0),.clk(gclk));
	jdff dff_A_lAIycoQE7_0(.dout(w_dff_A_7gBGe5ps6_0),.din(w_dff_A_lAIycoQE7_0),.clk(gclk));
	jdff dff_A_7gBGe5ps6_0(.dout(w_dff_A_BdaQd5Rb9_0),.din(w_dff_A_7gBGe5ps6_0),.clk(gclk));
	jdff dff_A_BdaQd5Rb9_0(.dout(w_dff_A_dbATNVWm6_0),.din(w_dff_A_BdaQd5Rb9_0),.clk(gclk));
	jdff dff_A_dbATNVWm6_0(.dout(w_dff_A_tBVi5mJQ8_0),.din(w_dff_A_dbATNVWm6_0),.clk(gclk));
	jdff dff_A_tBVi5mJQ8_0(.dout(w_dff_A_INDGoFkg3_0),.din(w_dff_A_tBVi5mJQ8_0),.clk(gclk));
	jdff dff_A_INDGoFkg3_0(.dout(w_dff_A_2tnSaPAX0_0),.din(w_dff_A_INDGoFkg3_0),.clk(gclk));
	jdff dff_A_2tnSaPAX0_0(.dout(w_dff_A_epFCYmGl7_0),.din(w_dff_A_2tnSaPAX0_0),.clk(gclk));
	jdff dff_A_epFCYmGl7_0(.dout(w_dff_A_EsqYMR8O7_0),.din(w_dff_A_epFCYmGl7_0),.clk(gclk));
	jdff dff_A_EsqYMR8O7_0(.dout(w_dff_A_zs9xhk1c1_0),.din(w_dff_A_EsqYMR8O7_0),.clk(gclk));
	jdff dff_A_zs9xhk1c1_0(.dout(w_dff_A_SShDmPL80_0),.din(w_dff_A_zs9xhk1c1_0),.clk(gclk));
	jdff dff_A_SShDmPL80_0(.dout(w_dff_A_UXcMNORi3_0),.din(w_dff_A_SShDmPL80_0),.clk(gclk));
	jdff dff_A_UXcMNORi3_0(.dout(w_dff_A_T0mmnZeG6_0),.din(w_dff_A_UXcMNORi3_0),.clk(gclk));
	jdff dff_A_T0mmnZeG6_0(.dout(w_dff_A_EEkZZj2h4_0),.din(w_dff_A_T0mmnZeG6_0),.clk(gclk));
	jdff dff_A_EEkZZj2h4_0(.dout(w_dff_A_rOD5n1Y23_0),.din(w_dff_A_EEkZZj2h4_0),.clk(gclk));
	jdff dff_A_rOD5n1Y23_0(.dout(w_dff_A_VBddhrBH2_0),.din(w_dff_A_rOD5n1Y23_0),.clk(gclk));
	jdff dff_A_VBddhrBH2_0(.dout(w_dff_A_rOO9VspZ6_0),.din(w_dff_A_VBddhrBH2_0),.clk(gclk));
	jdff dff_A_rOO9VspZ6_0(.dout(w_dff_A_CPjkiGVQ2_0),.din(w_dff_A_rOO9VspZ6_0),.clk(gclk));
	jdff dff_A_CPjkiGVQ2_0(.dout(w_dff_A_AL20DwRz2_0),.din(w_dff_A_CPjkiGVQ2_0),.clk(gclk));
	jdff dff_A_AL20DwRz2_0(.dout(w_dff_A_vwszhUu81_0),.din(w_dff_A_AL20DwRz2_0),.clk(gclk));
	jdff dff_A_vwszhUu81_0(.dout(w_dff_A_81v8lyms0_0),.din(w_dff_A_vwszhUu81_0),.clk(gclk));
	jdff dff_A_81v8lyms0_0(.dout(w_dff_A_WLCOgiXJ7_0),.din(w_dff_A_81v8lyms0_0),.clk(gclk));
	jdff dff_A_WLCOgiXJ7_0(.dout(w_dff_A_0Lq0JNAS8_0),.din(w_dff_A_WLCOgiXJ7_0),.clk(gclk));
	jdff dff_A_0Lq0JNAS8_0(.dout(w_dff_A_vRK7OhD86_0),.din(w_dff_A_0Lq0JNAS8_0),.clk(gclk));
	jdff dff_A_vRK7OhD86_0(.dout(w_dff_A_q6O0bSP29_0),.din(w_dff_A_vRK7OhD86_0),.clk(gclk));
	jdff dff_A_q6O0bSP29_0(.dout(w_dff_A_lamaJPT51_0),.din(w_dff_A_q6O0bSP29_0),.clk(gclk));
	jdff dff_A_lamaJPT51_0(.dout(w_dff_A_blGfFtq53_0),.din(w_dff_A_lamaJPT51_0),.clk(gclk));
	jdff dff_A_blGfFtq53_0(.dout(G1581gat),.din(w_dff_A_blGfFtq53_0),.clk(gclk));
	jdff dff_A_buo4FdL10_2(.dout(w_dff_A_TXQDmXQu9_0),.din(w_dff_A_buo4FdL10_2),.clk(gclk));
	jdff dff_A_TXQDmXQu9_0(.dout(w_dff_A_poLHy51T9_0),.din(w_dff_A_TXQDmXQu9_0),.clk(gclk));
	jdff dff_A_poLHy51T9_0(.dout(w_dff_A_G7Yi1Tj75_0),.din(w_dff_A_poLHy51T9_0),.clk(gclk));
	jdff dff_A_G7Yi1Tj75_0(.dout(w_dff_A_JBM5vqQf6_0),.din(w_dff_A_G7Yi1Tj75_0),.clk(gclk));
	jdff dff_A_JBM5vqQf6_0(.dout(w_dff_A_WaoXTjPl0_0),.din(w_dff_A_JBM5vqQf6_0),.clk(gclk));
	jdff dff_A_WaoXTjPl0_0(.dout(w_dff_A_WOiBWxin6_0),.din(w_dff_A_WaoXTjPl0_0),.clk(gclk));
	jdff dff_A_WOiBWxin6_0(.dout(w_dff_A_X7s0jOUv1_0),.din(w_dff_A_WOiBWxin6_0),.clk(gclk));
	jdff dff_A_X7s0jOUv1_0(.dout(w_dff_A_NBJwJOM78_0),.din(w_dff_A_X7s0jOUv1_0),.clk(gclk));
	jdff dff_A_NBJwJOM78_0(.dout(w_dff_A_7Q7l75KR3_0),.din(w_dff_A_NBJwJOM78_0),.clk(gclk));
	jdff dff_A_7Q7l75KR3_0(.dout(w_dff_A_95RTOtd64_0),.din(w_dff_A_7Q7l75KR3_0),.clk(gclk));
	jdff dff_A_95RTOtd64_0(.dout(w_dff_A_smRvgRlM3_0),.din(w_dff_A_95RTOtd64_0),.clk(gclk));
	jdff dff_A_smRvgRlM3_0(.dout(w_dff_A_IScTT8RI7_0),.din(w_dff_A_smRvgRlM3_0),.clk(gclk));
	jdff dff_A_IScTT8RI7_0(.dout(w_dff_A_kwZ2gT2t5_0),.din(w_dff_A_IScTT8RI7_0),.clk(gclk));
	jdff dff_A_kwZ2gT2t5_0(.dout(w_dff_A_zbTTgX4P1_0),.din(w_dff_A_kwZ2gT2t5_0),.clk(gclk));
	jdff dff_A_zbTTgX4P1_0(.dout(w_dff_A_WijUF9467_0),.din(w_dff_A_zbTTgX4P1_0),.clk(gclk));
	jdff dff_A_WijUF9467_0(.dout(w_dff_A_g0eAg3Co1_0),.din(w_dff_A_WijUF9467_0),.clk(gclk));
	jdff dff_A_g0eAg3Co1_0(.dout(w_dff_A_57ZLz1p54_0),.din(w_dff_A_g0eAg3Co1_0),.clk(gclk));
	jdff dff_A_57ZLz1p54_0(.dout(w_dff_A_Ie2YxNOe9_0),.din(w_dff_A_57ZLz1p54_0),.clk(gclk));
	jdff dff_A_Ie2YxNOe9_0(.dout(w_dff_A_rmuaJVc84_0),.din(w_dff_A_Ie2YxNOe9_0),.clk(gclk));
	jdff dff_A_rmuaJVc84_0(.dout(w_dff_A_kW8m9Uc21_0),.din(w_dff_A_rmuaJVc84_0),.clk(gclk));
	jdff dff_A_kW8m9Uc21_0(.dout(w_dff_A_7hQEarXC6_0),.din(w_dff_A_kW8m9Uc21_0),.clk(gclk));
	jdff dff_A_7hQEarXC6_0(.dout(w_dff_A_NsfJuRvx0_0),.din(w_dff_A_7hQEarXC6_0),.clk(gclk));
	jdff dff_A_NsfJuRvx0_0(.dout(w_dff_A_lySbVBV65_0),.din(w_dff_A_NsfJuRvx0_0),.clk(gclk));
	jdff dff_A_lySbVBV65_0(.dout(w_dff_A_AhkEpVkb3_0),.din(w_dff_A_lySbVBV65_0),.clk(gclk));
	jdff dff_A_AhkEpVkb3_0(.dout(w_dff_A_AARyv2OZ4_0),.din(w_dff_A_AhkEpVkb3_0),.clk(gclk));
	jdff dff_A_AARyv2OZ4_0(.dout(w_dff_A_nv6ZFavq7_0),.din(w_dff_A_AARyv2OZ4_0),.clk(gclk));
	jdff dff_A_nv6ZFavq7_0(.dout(w_dff_A_fIYMeOPI7_0),.din(w_dff_A_nv6ZFavq7_0),.clk(gclk));
	jdff dff_A_fIYMeOPI7_0(.dout(w_dff_A_FMlrkncn3_0),.din(w_dff_A_fIYMeOPI7_0),.clk(gclk));
	jdff dff_A_FMlrkncn3_0(.dout(w_dff_A_seEZ09Bf8_0),.din(w_dff_A_FMlrkncn3_0),.clk(gclk));
	jdff dff_A_seEZ09Bf8_0(.dout(w_dff_A_XvhIP3zA9_0),.din(w_dff_A_seEZ09Bf8_0),.clk(gclk));
	jdff dff_A_XvhIP3zA9_0(.dout(w_dff_A_CqixKKVX0_0),.din(w_dff_A_XvhIP3zA9_0),.clk(gclk));
	jdff dff_A_CqixKKVX0_0(.dout(w_dff_A_gz1GsxHp5_0),.din(w_dff_A_CqixKKVX0_0),.clk(gclk));
	jdff dff_A_gz1GsxHp5_0(.dout(w_dff_A_Tyj5oO2W9_0),.din(w_dff_A_gz1GsxHp5_0),.clk(gclk));
	jdff dff_A_Tyj5oO2W9_0(.dout(w_dff_A_R7C45UMu6_0),.din(w_dff_A_Tyj5oO2W9_0),.clk(gclk));
	jdff dff_A_R7C45UMu6_0(.dout(w_dff_A_kyvCI4jS6_0),.din(w_dff_A_R7C45UMu6_0),.clk(gclk));
	jdff dff_A_kyvCI4jS6_0(.dout(w_dff_A_hdGFVPii0_0),.din(w_dff_A_kyvCI4jS6_0),.clk(gclk));
	jdff dff_A_hdGFVPii0_0(.dout(w_dff_A_mAfEbpZI0_0),.din(w_dff_A_hdGFVPii0_0),.clk(gclk));
	jdff dff_A_mAfEbpZI0_0(.dout(w_dff_A_CoeC1kwg1_0),.din(w_dff_A_mAfEbpZI0_0),.clk(gclk));
	jdff dff_A_CoeC1kwg1_0(.dout(w_dff_A_IGxYFOR93_0),.din(w_dff_A_CoeC1kwg1_0),.clk(gclk));
	jdff dff_A_IGxYFOR93_0(.dout(w_dff_A_Vw5fECnz2_0),.din(w_dff_A_IGxYFOR93_0),.clk(gclk));
	jdff dff_A_Vw5fECnz2_0(.dout(w_dff_A_WpnxNDUE8_0),.din(w_dff_A_Vw5fECnz2_0),.clk(gclk));
	jdff dff_A_WpnxNDUE8_0(.dout(w_dff_A_1YDCgfkD9_0),.din(w_dff_A_WpnxNDUE8_0),.clk(gclk));
	jdff dff_A_1YDCgfkD9_0(.dout(w_dff_A_OLAfH0io7_0),.din(w_dff_A_1YDCgfkD9_0),.clk(gclk));
	jdff dff_A_OLAfH0io7_0(.dout(w_dff_A_jBE172ew3_0),.din(w_dff_A_OLAfH0io7_0),.clk(gclk));
	jdff dff_A_jBE172ew3_0(.dout(w_dff_A_LmlYMnMJ8_0),.din(w_dff_A_jBE172ew3_0),.clk(gclk));
	jdff dff_A_LmlYMnMJ8_0(.dout(w_dff_A_Gr02eWPc5_0),.din(w_dff_A_LmlYMnMJ8_0),.clk(gclk));
	jdff dff_A_Gr02eWPc5_0(.dout(w_dff_A_l8jeQ4254_0),.din(w_dff_A_Gr02eWPc5_0),.clk(gclk));
	jdff dff_A_l8jeQ4254_0(.dout(w_dff_A_JBUAY8Fw0_0),.din(w_dff_A_l8jeQ4254_0),.clk(gclk));
	jdff dff_A_JBUAY8Fw0_0(.dout(w_dff_A_6zutFgaU6_0),.din(w_dff_A_JBUAY8Fw0_0),.clk(gclk));
	jdff dff_A_6zutFgaU6_0(.dout(w_dff_A_rp2XgVWh3_0),.din(w_dff_A_6zutFgaU6_0),.clk(gclk));
	jdff dff_A_rp2XgVWh3_0(.dout(w_dff_A_6wZbilJl2_0),.din(w_dff_A_rp2XgVWh3_0),.clk(gclk));
	jdff dff_A_6wZbilJl2_0(.dout(w_dff_A_GnMpStnz1_0),.din(w_dff_A_6wZbilJl2_0),.clk(gclk));
	jdff dff_A_GnMpStnz1_0(.dout(w_dff_A_cMcUBohz8_0),.din(w_dff_A_GnMpStnz1_0),.clk(gclk));
	jdff dff_A_cMcUBohz8_0(.dout(w_dff_A_UI1R9Le08_0),.din(w_dff_A_cMcUBohz8_0),.clk(gclk));
	jdff dff_A_UI1R9Le08_0(.dout(w_dff_A_w8sKohNk5_0),.din(w_dff_A_UI1R9Le08_0),.clk(gclk));
	jdff dff_A_w8sKohNk5_0(.dout(w_dff_A_zlcWMyib6_0),.din(w_dff_A_w8sKohNk5_0),.clk(gclk));
	jdff dff_A_zlcWMyib6_0(.dout(w_dff_A_O0SO8ROF3_0),.din(w_dff_A_zlcWMyib6_0),.clk(gclk));
	jdff dff_A_O0SO8ROF3_0(.dout(w_dff_A_MdHWVO2B3_0),.din(w_dff_A_O0SO8ROF3_0),.clk(gclk));
	jdff dff_A_MdHWVO2B3_0(.dout(w_dff_A_paKgfGkd1_0),.din(w_dff_A_MdHWVO2B3_0),.clk(gclk));
	jdff dff_A_paKgfGkd1_0(.dout(w_dff_A_c4TVz89o2_0),.din(w_dff_A_paKgfGkd1_0),.clk(gclk));
	jdff dff_A_c4TVz89o2_0(.dout(w_dff_A_wGpiu0r74_0),.din(w_dff_A_c4TVz89o2_0),.clk(gclk));
	jdff dff_A_wGpiu0r74_0(.dout(w_dff_A_U6lDBDTs0_0),.din(w_dff_A_wGpiu0r74_0),.clk(gclk));
	jdff dff_A_U6lDBDTs0_0(.dout(w_dff_A_ZI9Vowwm3_0),.din(w_dff_A_U6lDBDTs0_0),.clk(gclk));
	jdff dff_A_ZI9Vowwm3_0(.dout(w_dff_A_DHpCUB6Q1_0),.din(w_dff_A_ZI9Vowwm3_0),.clk(gclk));
	jdff dff_A_DHpCUB6Q1_0(.dout(w_dff_A_yKS96IHA5_0),.din(w_dff_A_DHpCUB6Q1_0),.clk(gclk));
	jdff dff_A_yKS96IHA5_0(.dout(w_dff_A_yyGiPMnY0_0),.din(w_dff_A_yKS96IHA5_0),.clk(gclk));
	jdff dff_A_yyGiPMnY0_0(.dout(w_dff_A_vUbw6a1X3_0),.din(w_dff_A_yyGiPMnY0_0),.clk(gclk));
	jdff dff_A_vUbw6a1X3_0(.dout(w_dff_A_5QNzbAT64_0),.din(w_dff_A_vUbw6a1X3_0),.clk(gclk));
	jdff dff_A_5QNzbAT64_0(.dout(G1901gat),.din(w_dff_A_5QNzbAT64_0),.clk(gclk));
	jdff dff_A_dMBLpPmk9_2(.dout(w_dff_A_w7Qg4Ogm6_0),.din(w_dff_A_dMBLpPmk9_2),.clk(gclk));
	jdff dff_A_w7Qg4Ogm6_0(.dout(w_dff_A_aAxv4qMc1_0),.din(w_dff_A_w7Qg4Ogm6_0),.clk(gclk));
	jdff dff_A_aAxv4qMc1_0(.dout(w_dff_A_ItSyCivU4_0),.din(w_dff_A_aAxv4qMc1_0),.clk(gclk));
	jdff dff_A_ItSyCivU4_0(.dout(w_dff_A_KceAzcYC0_0),.din(w_dff_A_ItSyCivU4_0),.clk(gclk));
	jdff dff_A_KceAzcYC0_0(.dout(w_dff_A_DJaz2nfu9_0),.din(w_dff_A_KceAzcYC0_0),.clk(gclk));
	jdff dff_A_DJaz2nfu9_0(.dout(w_dff_A_DL4jujl76_0),.din(w_dff_A_DJaz2nfu9_0),.clk(gclk));
	jdff dff_A_DL4jujl76_0(.dout(w_dff_A_M7REda1w2_0),.din(w_dff_A_DL4jujl76_0),.clk(gclk));
	jdff dff_A_M7REda1w2_0(.dout(w_dff_A_T7K3CaY87_0),.din(w_dff_A_M7REda1w2_0),.clk(gclk));
	jdff dff_A_T7K3CaY87_0(.dout(w_dff_A_hmRtgyuR3_0),.din(w_dff_A_T7K3CaY87_0),.clk(gclk));
	jdff dff_A_hmRtgyuR3_0(.dout(w_dff_A_0sdC5CQt8_0),.din(w_dff_A_hmRtgyuR3_0),.clk(gclk));
	jdff dff_A_0sdC5CQt8_0(.dout(w_dff_A_3ho92WB04_0),.din(w_dff_A_0sdC5CQt8_0),.clk(gclk));
	jdff dff_A_3ho92WB04_0(.dout(w_dff_A_Ytp4l8vM7_0),.din(w_dff_A_3ho92WB04_0),.clk(gclk));
	jdff dff_A_Ytp4l8vM7_0(.dout(w_dff_A_mEgezkWX4_0),.din(w_dff_A_Ytp4l8vM7_0),.clk(gclk));
	jdff dff_A_mEgezkWX4_0(.dout(w_dff_A_n0dU0Hwf3_0),.din(w_dff_A_mEgezkWX4_0),.clk(gclk));
	jdff dff_A_n0dU0Hwf3_0(.dout(w_dff_A_sANRdrOi4_0),.din(w_dff_A_n0dU0Hwf3_0),.clk(gclk));
	jdff dff_A_sANRdrOi4_0(.dout(w_dff_A_VoeJeHDR0_0),.din(w_dff_A_sANRdrOi4_0),.clk(gclk));
	jdff dff_A_VoeJeHDR0_0(.dout(w_dff_A_R5d8JNCG8_0),.din(w_dff_A_VoeJeHDR0_0),.clk(gclk));
	jdff dff_A_R5d8JNCG8_0(.dout(w_dff_A_LkTXmiTN2_0),.din(w_dff_A_R5d8JNCG8_0),.clk(gclk));
	jdff dff_A_LkTXmiTN2_0(.dout(w_dff_A_44b5Za3q0_0),.din(w_dff_A_LkTXmiTN2_0),.clk(gclk));
	jdff dff_A_44b5Za3q0_0(.dout(w_dff_A_65S7st0f9_0),.din(w_dff_A_44b5Za3q0_0),.clk(gclk));
	jdff dff_A_65S7st0f9_0(.dout(w_dff_A_qez06FdT3_0),.din(w_dff_A_65S7st0f9_0),.clk(gclk));
	jdff dff_A_qez06FdT3_0(.dout(w_dff_A_jIfjbs3p4_0),.din(w_dff_A_qez06FdT3_0),.clk(gclk));
	jdff dff_A_jIfjbs3p4_0(.dout(w_dff_A_Lp23YidW0_0),.din(w_dff_A_jIfjbs3p4_0),.clk(gclk));
	jdff dff_A_Lp23YidW0_0(.dout(w_dff_A_liEFXoqg6_0),.din(w_dff_A_Lp23YidW0_0),.clk(gclk));
	jdff dff_A_liEFXoqg6_0(.dout(w_dff_A_iSUWP2vl4_0),.din(w_dff_A_liEFXoqg6_0),.clk(gclk));
	jdff dff_A_iSUWP2vl4_0(.dout(w_dff_A_0VBGkh5x9_0),.din(w_dff_A_iSUWP2vl4_0),.clk(gclk));
	jdff dff_A_0VBGkh5x9_0(.dout(w_dff_A_shQg4kMP0_0),.din(w_dff_A_0VBGkh5x9_0),.clk(gclk));
	jdff dff_A_shQg4kMP0_0(.dout(w_dff_A_i74p85CP1_0),.din(w_dff_A_shQg4kMP0_0),.clk(gclk));
	jdff dff_A_i74p85CP1_0(.dout(w_dff_A_htM5lZks8_0),.din(w_dff_A_i74p85CP1_0),.clk(gclk));
	jdff dff_A_htM5lZks8_0(.dout(w_dff_A_6VIPgpEI3_0),.din(w_dff_A_htM5lZks8_0),.clk(gclk));
	jdff dff_A_6VIPgpEI3_0(.dout(w_dff_A_mpJjQPkg4_0),.din(w_dff_A_6VIPgpEI3_0),.clk(gclk));
	jdff dff_A_mpJjQPkg4_0(.dout(w_dff_A_OO8pCVS49_0),.din(w_dff_A_mpJjQPkg4_0),.clk(gclk));
	jdff dff_A_OO8pCVS49_0(.dout(w_dff_A_mSmIWK7j9_0),.din(w_dff_A_OO8pCVS49_0),.clk(gclk));
	jdff dff_A_mSmIWK7j9_0(.dout(w_dff_A_u0gJUiq52_0),.din(w_dff_A_mSmIWK7j9_0),.clk(gclk));
	jdff dff_A_u0gJUiq52_0(.dout(w_dff_A_y9xN8TYu4_0),.din(w_dff_A_u0gJUiq52_0),.clk(gclk));
	jdff dff_A_y9xN8TYu4_0(.dout(w_dff_A_Sr626VtM9_0),.din(w_dff_A_y9xN8TYu4_0),.clk(gclk));
	jdff dff_A_Sr626VtM9_0(.dout(w_dff_A_adCT9SwV1_0),.din(w_dff_A_Sr626VtM9_0),.clk(gclk));
	jdff dff_A_adCT9SwV1_0(.dout(w_dff_A_79qyOkIc4_0),.din(w_dff_A_adCT9SwV1_0),.clk(gclk));
	jdff dff_A_79qyOkIc4_0(.dout(w_dff_A_yWsc2FG58_0),.din(w_dff_A_79qyOkIc4_0),.clk(gclk));
	jdff dff_A_yWsc2FG58_0(.dout(w_dff_A_XvVgFn9P0_0),.din(w_dff_A_yWsc2FG58_0),.clk(gclk));
	jdff dff_A_XvVgFn9P0_0(.dout(w_dff_A_pBRyccUm1_0),.din(w_dff_A_XvVgFn9P0_0),.clk(gclk));
	jdff dff_A_pBRyccUm1_0(.dout(w_dff_A_urcuM0of9_0),.din(w_dff_A_pBRyccUm1_0),.clk(gclk));
	jdff dff_A_urcuM0of9_0(.dout(w_dff_A_YsSHIPp28_0),.din(w_dff_A_urcuM0of9_0),.clk(gclk));
	jdff dff_A_YsSHIPp28_0(.dout(w_dff_A_vL4YCkmB6_0),.din(w_dff_A_YsSHIPp28_0),.clk(gclk));
	jdff dff_A_vL4YCkmB6_0(.dout(w_dff_A_7ao35V7m9_0),.din(w_dff_A_vL4YCkmB6_0),.clk(gclk));
	jdff dff_A_7ao35V7m9_0(.dout(w_dff_A_KPVd0E3G7_0),.din(w_dff_A_7ao35V7m9_0),.clk(gclk));
	jdff dff_A_KPVd0E3G7_0(.dout(w_dff_A_C84v9WI28_0),.din(w_dff_A_KPVd0E3G7_0),.clk(gclk));
	jdff dff_A_C84v9WI28_0(.dout(w_dff_A_merpgjMT5_0),.din(w_dff_A_C84v9WI28_0),.clk(gclk));
	jdff dff_A_merpgjMT5_0(.dout(w_dff_A_i29UEyo96_0),.din(w_dff_A_merpgjMT5_0),.clk(gclk));
	jdff dff_A_i29UEyo96_0(.dout(w_dff_A_6Ljx9aGY4_0),.din(w_dff_A_i29UEyo96_0),.clk(gclk));
	jdff dff_A_6Ljx9aGY4_0(.dout(w_dff_A_8WYA2Jd19_0),.din(w_dff_A_6Ljx9aGY4_0),.clk(gclk));
	jdff dff_A_8WYA2Jd19_0(.dout(w_dff_A_waG2YfAb8_0),.din(w_dff_A_8WYA2Jd19_0),.clk(gclk));
	jdff dff_A_waG2YfAb8_0(.dout(w_dff_A_MZG1aCZA7_0),.din(w_dff_A_waG2YfAb8_0),.clk(gclk));
	jdff dff_A_MZG1aCZA7_0(.dout(w_dff_A_sqbHbFPC4_0),.din(w_dff_A_MZG1aCZA7_0),.clk(gclk));
	jdff dff_A_sqbHbFPC4_0(.dout(w_dff_A_LS7bFTju7_0),.din(w_dff_A_sqbHbFPC4_0),.clk(gclk));
	jdff dff_A_LS7bFTju7_0(.dout(w_dff_A_RZtG7oBe2_0),.din(w_dff_A_LS7bFTju7_0),.clk(gclk));
	jdff dff_A_RZtG7oBe2_0(.dout(w_dff_A_Lo4r26GP1_0),.din(w_dff_A_RZtG7oBe2_0),.clk(gclk));
	jdff dff_A_Lo4r26GP1_0(.dout(w_dff_A_XNimF5mI3_0),.din(w_dff_A_Lo4r26GP1_0),.clk(gclk));
	jdff dff_A_XNimF5mI3_0(.dout(w_dff_A_48zxiKJh3_0),.din(w_dff_A_XNimF5mI3_0),.clk(gclk));
	jdff dff_A_48zxiKJh3_0(.dout(w_dff_A_HXAkp2Hr2_0),.din(w_dff_A_48zxiKJh3_0),.clk(gclk));
	jdff dff_A_HXAkp2Hr2_0(.dout(w_dff_A_D98vrOpP9_0),.din(w_dff_A_HXAkp2Hr2_0),.clk(gclk));
	jdff dff_A_D98vrOpP9_0(.dout(w_dff_A_SbpdLbA98_0),.din(w_dff_A_D98vrOpP9_0),.clk(gclk));
	jdff dff_A_SbpdLbA98_0(.dout(w_dff_A_vjiFzC1H3_0),.din(w_dff_A_SbpdLbA98_0),.clk(gclk));
	jdff dff_A_vjiFzC1H3_0(.dout(w_dff_A_O6hg4Dry9_0),.din(w_dff_A_vjiFzC1H3_0),.clk(gclk));
	jdff dff_A_O6hg4Dry9_0(.dout(w_dff_A_7yE0NEGK3_0),.din(w_dff_A_O6hg4Dry9_0),.clk(gclk));
	jdff dff_A_7yE0NEGK3_0(.dout(G2223gat),.din(w_dff_A_7yE0NEGK3_0),.clk(gclk));
	jdff dff_A_gefk1wav5_2(.dout(w_dff_A_DWMixp4U9_0),.din(w_dff_A_gefk1wav5_2),.clk(gclk));
	jdff dff_A_DWMixp4U9_0(.dout(w_dff_A_yy540UXo8_0),.din(w_dff_A_DWMixp4U9_0),.clk(gclk));
	jdff dff_A_yy540UXo8_0(.dout(w_dff_A_qRfJJhsW8_0),.din(w_dff_A_yy540UXo8_0),.clk(gclk));
	jdff dff_A_qRfJJhsW8_0(.dout(w_dff_A_oTtkERGX3_0),.din(w_dff_A_qRfJJhsW8_0),.clk(gclk));
	jdff dff_A_oTtkERGX3_0(.dout(w_dff_A_5waJCCo93_0),.din(w_dff_A_oTtkERGX3_0),.clk(gclk));
	jdff dff_A_5waJCCo93_0(.dout(w_dff_A_9QY3BGhr5_0),.din(w_dff_A_5waJCCo93_0),.clk(gclk));
	jdff dff_A_9QY3BGhr5_0(.dout(w_dff_A_U5OLYsr97_0),.din(w_dff_A_9QY3BGhr5_0),.clk(gclk));
	jdff dff_A_U5OLYsr97_0(.dout(w_dff_A_pRcNIFEJ4_0),.din(w_dff_A_U5OLYsr97_0),.clk(gclk));
	jdff dff_A_pRcNIFEJ4_0(.dout(w_dff_A_ABzoDVs39_0),.din(w_dff_A_pRcNIFEJ4_0),.clk(gclk));
	jdff dff_A_ABzoDVs39_0(.dout(w_dff_A_pFZUHEKQ7_0),.din(w_dff_A_ABzoDVs39_0),.clk(gclk));
	jdff dff_A_pFZUHEKQ7_0(.dout(w_dff_A_w4Aj6XlB2_0),.din(w_dff_A_pFZUHEKQ7_0),.clk(gclk));
	jdff dff_A_w4Aj6XlB2_0(.dout(w_dff_A_yIzZqKfb5_0),.din(w_dff_A_w4Aj6XlB2_0),.clk(gclk));
	jdff dff_A_yIzZqKfb5_0(.dout(w_dff_A_kTaoyh0S4_0),.din(w_dff_A_yIzZqKfb5_0),.clk(gclk));
	jdff dff_A_kTaoyh0S4_0(.dout(w_dff_A_BHdxHAt01_0),.din(w_dff_A_kTaoyh0S4_0),.clk(gclk));
	jdff dff_A_BHdxHAt01_0(.dout(w_dff_A_EErckhbs1_0),.din(w_dff_A_BHdxHAt01_0),.clk(gclk));
	jdff dff_A_EErckhbs1_0(.dout(w_dff_A_5n9ZpK7C5_0),.din(w_dff_A_EErckhbs1_0),.clk(gclk));
	jdff dff_A_5n9ZpK7C5_0(.dout(w_dff_A_vDpKBRS55_0),.din(w_dff_A_5n9ZpK7C5_0),.clk(gclk));
	jdff dff_A_vDpKBRS55_0(.dout(w_dff_A_xY2YEdT17_0),.din(w_dff_A_vDpKBRS55_0),.clk(gclk));
	jdff dff_A_xY2YEdT17_0(.dout(w_dff_A_O1FQhSMu2_0),.din(w_dff_A_xY2YEdT17_0),.clk(gclk));
	jdff dff_A_O1FQhSMu2_0(.dout(w_dff_A_KwVgtCfR3_0),.din(w_dff_A_O1FQhSMu2_0),.clk(gclk));
	jdff dff_A_KwVgtCfR3_0(.dout(w_dff_A_X8hL8fkt7_0),.din(w_dff_A_KwVgtCfR3_0),.clk(gclk));
	jdff dff_A_X8hL8fkt7_0(.dout(w_dff_A_UJpwuqi06_0),.din(w_dff_A_X8hL8fkt7_0),.clk(gclk));
	jdff dff_A_UJpwuqi06_0(.dout(w_dff_A_KPqNtckk9_0),.din(w_dff_A_UJpwuqi06_0),.clk(gclk));
	jdff dff_A_KPqNtckk9_0(.dout(w_dff_A_Zuq8soWV9_0),.din(w_dff_A_KPqNtckk9_0),.clk(gclk));
	jdff dff_A_Zuq8soWV9_0(.dout(w_dff_A_aVzL60u73_0),.din(w_dff_A_Zuq8soWV9_0),.clk(gclk));
	jdff dff_A_aVzL60u73_0(.dout(w_dff_A_2XcVAt7h1_0),.din(w_dff_A_aVzL60u73_0),.clk(gclk));
	jdff dff_A_2XcVAt7h1_0(.dout(w_dff_A_vi7yjqHw6_0),.din(w_dff_A_2XcVAt7h1_0),.clk(gclk));
	jdff dff_A_vi7yjqHw6_0(.dout(w_dff_A_IOKbtvmm5_0),.din(w_dff_A_vi7yjqHw6_0),.clk(gclk));
	jdff dff_A_IOKbtvmm5_0(.dout(w_dff_A_nValV1yi1_0),.din(w_dff_A_IOKbtvmm5_0),.clk(gclk));
	jdff dff_A_nValV1yi1_0(.dout(w_dff_A_cYohB2Ig3_0),.din(w_dff_A_nValV1yi1_0),.clk(gclk));
	jdff dff_A_cYohB2Ig3_0(.dout(w_dff_A_fcy7mX9L5_0),.din(w_dff_A_cYohB2Ig3_0),.clk(gclk));
	jdff dff_A_fcy7mX9L5_0(.dout(w_dff_A_rV90dYuF4_0),.din(w_dff_A_fcy7mX9L5_0),.clk(gclk));
	jdff dff_A_rV90dYuF4_0(.dout(w_dff_A_IS1vNVL88_0),.din(w_dff_A_rV90dYuF4_0),.clk(gclk));
	jdff dff_A_IS1vNVL88_0(.dout(w_dff_A_8ObDaeqV8_0),.din(w_dff_A_IS1vNVL88_0),.clk(gclk));
	jdff dff_A_8ObDaeqV8_0(.dout(w_dff_A_NJuuxCSy0_0),.din(w_dff_A_8ObDaeqV8_0),.clk(gclk));
	jdff dff_A_NJuuxCSy0_0(.dout(w_dff_A_tExBP91x7_0),.din(w_dff_A_NJuuxCSy0_0),.clk(gclk));
	jdff dff_A_tExBP91x7_0(.dout(w_dff_A_fK22dD7y6_0),.din(w_dff_A_tExBP91x7_0),.clk(gclk));
	jdff dff_A_fK22dD7y6_0(.dout(w_dff_A_kQuEI4zD7_0),.din(w_dff_A_fK22dD7y6_0),.clk(gclk));
	jdff dff_A_kQuEI4zD7_0(.dout(w_dff_A_WdTMREwU5_0),.din(w_dff_A_kQuEI4zD7_0),.clk(gclk));
	jdff dff_A_WdTMREwU5_0(.dout(w_dff_A_fbPW6fY64_0),.din(w_dff_A_WdTMREwU5_0),.clk(gclk));
	jdff dff_A_fbPW6fY64_0(.dout(w_dff_A_I40QanF71_0),.din(w_dff_A_fbPW6fY64_0),.clk(gclk));
	jdff dff_A_I40QanF71_0(.dout(w_dff_A_KHz6G9TZ1_0),.din(w_dff_A_I40QanF71_0),.clk(gclk));
	jdff dff_A_KHz6G9TZ1_0(.dout(w_dff_A_EDJQ5LCw3_0),.din(w_dff_A_KHz6G9TZ1_0),.clk(gclk));
	jdff dff_A_EDJQ5LCw3_0(.dout(w_dff_A_UaAQEaEB1_0),.din(w_dff_A_EDJQ5LCw3_0),.clk(gclk));
	jdff dff_A_UaAQEaEB1_0(.dout(w_dff_A_cKcQoA330_0),.din(w_dff_A_UaAQEaEB1_0),.clk(gclk));
	jdff dff_A_cKcQoA330_0(.dout(w_dff_A_xLl8ZBKx4_0),.din(w_dff_A_cKcQoA330_0),.clk(gclk));
	jdff dff_A_xLl8ZBKx4_0(.dout(w_dff_A_Hy0Ia5YF8_0),.din(w_dff_A_xLl8ZBKx4_0),.clk(gclk));
	jdff dff_A_Hy0Ia5YF8_0(.dout(w_dff_A_MiTYFQNb2_0),.din(w_dff_A_Hy0Ia5YF8_0),.clk(gclk));
	jdff dff_A_MiTYFQNb2_0(.dout(w_dff_A_ej3NMY796_0),.din(w_dff_A_MiTYFQNb2_0),.clk(gclk));
	jdff dff_A_ej3NMY796_0(.dout(w_dff_A_zQLlC5Jg5_0),.din(w_dff_A_ej3NMY796_0),.clk(gclk));
	jdff dff_A_zQLlC5Jg5_0(.dout(w_dff_A_vGJVRWXF6_0),.din(w_dff_A_zQLlC5Jg5_0),.clk(gclk));
	jdff dff_A_vGJVRWXF6_0(.dout(w_dff_A_dbq52p2K5_0),.din(w_dff_A_vGJVRWXF6_0),.clk(gclk));
	jdff dff_A_dbq52p2K5_0(.dout(w_dff_A_wtIb7jUO1_0),.din(w_dff_A_dbq52p2K5_0),.clk(gclk));
	jdff dff_A_wtIb7jUO1_0(.dout(w_dff_A_aODrlKhT3_0),.din(w_dff_A_wtIb7jUO1_0),.clk(gclk));
	jdff dff_A_aODrlKhT3_0(.dout(w_dff_A_v01lq88z1_0),.din(w_dff_A_aODrlKhT3_0),.clk(gclk));
	jdff dff_A_v01lq88z1_0(.dout(w_dff_A_iVSpAhTK7_0),.din(w_dff_A_v01lq88z1_0),.clk(gclk));
	jdff dff_A_iVSpAhTK7_0(.dout(w_dff_A_7WfemrKq0_0),.din(w_dff_A_iVSpAhTK7_0),.clk(gclk));
	jdff dff_A_7WfemrKq0_0(.dout(w_dff_A_IgrKJTUo6_0),.din(w_dff_A_7WfemrKq0_0),.clk(gclk));
	jdff dff_A_IgrKJTUo6_0(.dout(w_dff_A_8ZFaHYJb2_0),.din(w_dff_A_IgrKJTUo6_0),.clk(gclk));
	jdff dff_A_8ZFaHYJb2_0(.dout(w_dff_A_Z8lnYFP37_0),.din(w_dff_A_8ZFaHYJb2_0),.clk(gclk));
	jdff dff_A_Z8lnYFP37_0(.dout(w_dff_A_x5RKSedm6_0),.din(w_dff_A_Z8lnYFP37_0),.clk(gclk));
	jdff dff_A_x5RKSedm6_0(.dout(w_dff_A_YIn3qLDg7_0),.din(w_dff_A_x5RKSedm6_0),.clk(gclk));
	jdff dff_A_YIn3qLDg7_0(.dout(G2548gat),.din(w_dff_A_YIn3qLDg7_0),.clk(gclk));
	jdff dff_A_4JhpDJQk1_2(.dout(w_dff_A_nscWjhLV4_0),.din(w_dff_A_4JhpDJQk1_2),.clk(gclk));
	jdff dff_A_nscWjhLV4_0(.dout(w_dff_A_QQtvKVR79_0),.din(w_dff_A_nscWjhLV4_0),.clk(gclk));
	jdff dff_A_QQtvKVR79_0(.dout(w_dff_A_zwrkMT7A1_0),.din(w_dff_A_QQtvKVR79_0),.clk(gclk));
	jdff dff_A_zwrkMT7A1_0(.dout(w_dff_A_QwIXjRXM8_0),.din(w_dff_A_zwrkMT7A1_0),.clk(gclk));
	jdff dff_A_QwIXjRXM8_0(.dout(w_dff_A_CQnTGkZN9_0),.din(w_dff_A_QwIXjRXM8_0),.clk(gclk));
	jdff dff_A_CQnTGkZN9_0(.dout(w_dff_A_FF4UYeuX9_0),.din(w_dff_A_CQnTGkZN9_0),.clk(gclk));
	jdff dff_A_FF4UYeuX9_0(.dout(w_dff_A_bo9Idjg63_0),.din(w_dff_A_FF4UYeuX9_0),.clk(gclk));
	jdff dff_A_bo9Idjg63_0(.dout(w_dff_A_alVAfPKn5_0),.din(w_dff_A_bo9Idjg63_0),.clk(gclk));
	jdff dff_A_alVAfPKn5_0(.dout(w_dff_A_0B793M7y4_0),.din(w_dff_A_alVAfPKn5_0),.clk(gclk));
	jdff dff_A_0B793M7y4_0(.dout(w_dff_A_hmCun4bB8_0),.din(w_dff_A_0B793M7y4_0),.clk(gclk));
	jdff dff_A_hmCun4bB8_0(.dout(w_dff_A_05M9lXxp1_0),.din(w_dff_A_hmCun4bB8_0),.clk(gclk));
	jdff dff_A_05M9lXxp1_0(.dout(w_dff_A_CIi0AJt59_0),.din(w_dff_A_05M9lXxp1_0),.clk(gclk));
	jdff dff_A_CIi0AJt59_0(.dout(w_dff_A_7tYKSSNk7_0),.din(w_dff_A_CIi0AJt59_0),.clk(gclk));
	jdff dff_A_7tYKSSNk7_0(.dout(w_dff_A_AH7xB5E76_0),.din(w_dff_A_7tYKSSNk7_0),.clk(gclk));
	jdff dff_A_AH7xB5E76_0(.dout(w_dff_A_K7xAnZbI1_0),.din(w_dff_A_AH7xB5E76_0),.clk(gclk));
	jdff dff_A_K7xAnZbI1_0(.dout(w_dff_A_2MQGX1sc5_0),.din(w_dff_A_K7xAnZbI1_0),.clk(gclk));
	jdff dff_A_2MQGX1sc5_0(.dout(w_dff_A_BXAf8yXK6_0),.din(w_dff_A_2MQGX1sc5_0),.clk(gclk));
	jdff dff_A_BXAf8yXK6_0(.dout(w_dff_A_NSmRaWpA6_0),.din(w_dff_A_BXAf8yXK6_0),.clk(gclk));
	jdff dff_A_NSmRaWpA6_0(.dout(w_dff_A_6S5w8DWx4_0),.din(w_dff_A_NSmRaWpA6_0),.clk(gclk));
	jdff dff_A_6S5w8DWx4_0(.dout(w_dff_A_bLq4l5x63_0),.din(w_dff_A_6S5w8DWx4_0),.clk(gclk));
	jdff dff_A_bLq4l5x63_0(.dout(w_dff_A_15wk6lWG7_0),.din(w_dff_A_bLq4l5x63_0),.clk(gclk));
	jdff dff_A_15wk6lWG7_0(.dout(w_dff_A_npCZH30I8_0),.din(w_dff_A_15wk6lWG7_0),.clk(gclk));
	jdff dff_A_npCZH30I8_0(.dout(w_dff_A_lEqnh4SU5_0),.din(w_dff_A_npCZH30I8_0),.clk(gclk));
	jdff dff_A_lEqnh4SU5_0(.dout(w_dff_A_pqHE9Al20_0),.din(w_dff_A_lEqnh4SU5_0),.clk(gclk));
	jdff dff_A_pqHE9Al20_0(.dout(w_dff_A_xRpkV9632_0),.din(w_dff_A_pqHE9Al20_0),.clk(gclk));
	jdff dff_A_xRpkV9632_0(.dout(w_dff_A_vCbl7ueO9_0),.din(w_dff_A_xRpkV9632_0),.clk(gclk));
	jdff dff_A_vCbl7ueO9_0(.dout(w_dff_A_MDG60FCl4_0),.din(w_dff_A_vCbl7ueO9_0),.clk(gclk));
	jdff dff_A_MDG60FCl4_0(.dout(w_dff_A_3ohWSRwp6_0),.din(w_dff_A_MDG60FCl4_0),.clk(gclk));
	jdff dff_A_3ohWSRwp6_0(.dout(w_dff_A_JpKvjN0Q8_0),.din(w_dff_A_3ohWSRwp6_0),.clk(gclk));
	jdff dff_A_JpKvjN0Q8_0(.dout(w_dff_A_8ctyCZPs9_0),.din(w_dff_A_JpKvjN0Q8_0),.clk(gclk));
	jdff dff_A_8ctyCZPs9_0(.dout(w_dff_A_dQW0Y0CM0_0),.din(w_dff_A_8ctyCZPs9_0),.clk(gclk));
	jdff dff_A_dQW0Y0CM0_0(.dout(w_dff_A_lIMMJ4mF0_0),.din(w_dff_A_dQW0Y0CM0_0),.clk(gclk));
	jdff dff_A_lIMMJ4mF0_0(.dout(w_dff_A_X3aSuwpr7_0),.din(w_dff_A_lIMMJ4mF0_0),.clk(gclk));
	jdff dff_A_X3aSuwpr7_0(.dout(w_dff_A_So9rCyCz4_0),.din(w_dff_A_X3aSuwpr7_0),.clk(gclk));
	jdff dff_A_So9rCyCz4_0(.dout(w_dff_A_0UJhvR7F7_0),.din(w_dff_A_So9rCyCz4_0),.clk(gclk));
	jdff dff_A_0UJhvR7F7_0(.dout(w_dff_A_XMy9xEqY6_0),.din(w_dff_A_0UJhvR7F7_0),.clk(gclk));
	jdff dff_A_XMy9xEqY6_0(.dout(w_dff_A_mKHUZWye9_0),.din(w_dff_A_XMy9xEqY6_0),.clk(gclk));
	jdff dff_A_mKHUZWye9_0(.dout(w_dff_A_wWWm1iD94_0),.din(w_dff_A_mKHUZWye9_0),.clk(gclk));
	jdff dff_A_wWWm1iD94_0(.dout(w_dff_A_lzbFtxis8_0),.din(w_dff_A_wWWm1iD94_0),.clk(gclk));
	jdff dff_A_lzbFtxis8_0(.dout(w_dff_A_LcacxyjB4_0),.din(w_dff_A_lzbFtxis8_0),.clk(gclk));
	jdff dff_A_LcacxyjB4_0(.dout(w_dff_A_pajuTJ4l9_0),.din(w_dff_A_LcacxyjB4_0),.clk(gclk));
	jdff dff_A_pajuTJ4l9_0(.dout(w_dff_A_gajrwyFc3_0),.din(w_dff_A_pajuTJ4l9_0),.clk(gclk));
	jdff dff_A_gajrwyFc3_0(.dout(w_dff_A_UbCLgaYO7_0),.din(w_dff_A_gajrwyFc3_0),.clk(gclk));
	jdff dff_A_UbCLgaYO7_0(.dout(w_dff_A_XSaSblFD4_0),.din(w_dff_A_UbCLgaYO7_0),.clk(gclk));
	jdff dff_A_XSaSblFD4_0(.dout(w_dff_A_q5LOD2tg7_0),.din(w_dff_A_XSaSblFD4_0),.clk(gclk));
	jdff dff_A_q5LOD2tg7_0(.dout(w_dff_A_diZSij045_0),.din(w_dff_A_q5LOD2tg7_0),.clk(gclk));
	jdff dff_A_diZSij045_0(.dout(w_dff_A_Ah9bIosR8_0),.din(w_dff_A_diZSij045_0),.clk(gclk));
	jdff dff_A_Ah9bIosR8_0(.dout(w_dff_A_X2xmfMcN5_0),.din(w_dff_A_Ah9bIosR8_0),.clk(gclk));
	jdff dff_A_X2xmfMcN5_0(.dout(w_dff_A_2stJmJAI3_0),.din(w_dff_A_X2xmfMcN5_0),.clk(gclk));
	jdff dff_A_2stJmJAI3_0(.dout(w_dff_A_C3F1ytOH2_0),.din(w_dff_A_2stJmJAI3_0),.clk(gclk));
	jdff dff_A_C3F1ytOH2_0(.dout(w_dff_A_IRQLmgfl1_0),.din(w_dff_A_C3F1ytOH2_0),.clk(gclk));
	jdff dff_A_IRQLmgfl1_0(.dout(w_dff_A_33pAvLiG4_0),.din(w_dff_A_IRQLmgfl1_0),.clk(gclk));
	jdff dff_A_33pAvLiG4_0(.dout(w_dff_A_VDOZAGKJ3_0),.din(w_dff_A_33pAvLiG4_0),.clk(gclk));
	jdff dff_A_VDOZAGKJ3_0(.dout(w_dff_A_D67H8ryT4_0),.din(w_dff_A_VDOZAGKJ3_0),.clk(gclk));
	jdff dff_A_D67H8ryT4_0(.dout(w_dff_A_ZcD82bRK2_0),.din(w_dff_A_D67H8ryT4_0),.clk(gclk));
	jdff dff_A_ZcD82bRK2_0(.dout(w_dff_A_gffDqlbO2_0),.din(w_dff_A_ZcD82bRK2_0),.clk(gclk));
	jdff dff_A_gffDqlbO2_0(.dout(w_dff_A_jMtAlfG86_0),.din(w_dff_A_gffDqlbO2_0),.clk(gclk));
	jdff dff_A_jMtAlfG86_0(.dout(w_dff_A_PIQxSxvV7_0),.din(w_dff_A_jMtAlfG86_0),.clk(gclk));
	jdff dff_A_PIQxSxvV7_0(.dout(w_dff_A_V5ARinu60_0),.din(w_dff_A_PIQxSxvV7_0),.clk(gclk));
	jdff dff_A_V5ARinu60_0(.dout(G2877gat),.din(w_dff_A_V5ARinu60_0),.clk(gclk));
	jdff dff_A_fzty24Fg7_2(.dout(w_dff_A_6iTRBODh0_0),.din(w_dff_A_fzty24Fg7_2),.clk(gclk));
	jdff dff_A_6iTRBODh0_0(.dout(w_dff_A_m3ufP3LF0_0),.din(w_dff_A_6iTRBODh0_0),.clk(gclk));
	jdff dff_A_m3ufP3LF0_0(.dout(w_dff_A_22qSoX7d0_0),.din(w_dff_A_m3ufP3LF0_0),.clk(gclk));
	jdff dff_A_22qSoX7d0_0(.dout(w_dff_A_ijIFejDa8_0),.din(w_dff_A_22qSoX7d0_0),.clk(gclk));
	jdff dff_A_ijIFejDa8_0(.dout(w_dff_A_RMJAOgWq7_0),.din(w_dff_A_ijIFejDa8_0),.clk(gclk));
	jdff dff_A_RMJAOgWq7_0(.dout(w_dff_A_OOkiQ2DN0_0),.din(w_dff_A_RMJAOgWq7_0),.clk(gclk));
	jdff dff_A_OOkiQ2DN0_0(.dout(w_dff_A_1nyx4VDY1_0),.din(w_dff_A_OOkiQ2DN0_0),.clk(gclk));
	jdff dff_A_1nyx4VDY1_0(.dout(w_dff_A_gKZFgW2Y3_0),.din(w_dff_A_1nyx4VDY1_0),.clk(gclk));
	jdff dff_A_gKZFgW2Y3_0(.dout(w_dff_A_bSzpXqiR9_0),.din(w_dff_A_gKZFgW2Y3_0),.clk(gclk));
	jdff dff_A_bSzpXqiR9_0(.dout(w_dff_A_vxA7COBK1_0),.din(w_dff_A_bSzpXqiR9_0),.clk(gclk));
	jdff dff_A_vxA7COBK1_0(.dout(w_dff_A_AGXvGq6D7_0),.din(w_dff_A_vxA7COBK1_0),.clk(gclk));
	jdff dff_A_AGXvGq6D7_0(.dout(w_dff_A_KINI6req8_0),.din(w_dff_A_AGXvGq6D7_0),.clk(gclk));
	jdff dff_A_KINI6req8_0(.dout(w_dff_A_EAgXLHIO1_0),.din(w_dff_A_KINI6req8_0),.clk(gclk));
	jdff dff_A_EAgXLHIO1_0(.dout(w_dff_A_2KUCl9DI3_0),.din(w_dff_A_EAgXLHIO1_0),.clk(gclk));
	jdff dff_A_2KUCl9DI3_0(.dout(w_dff_A_8NgEBRJE8_0),.din(w_dff_A_2KUCl9DI3_0),.clk(gclk));
	jdff dff_A_8NgEBRJE8_0(.dout(w_dff_A_R16Af9wA2_0),.din(w_dff_A_8NgEBRJE8_0),.clk(gclk));
	jdff dff_A_R16Af9wA2_0(.dout(w_dff_A_dlri9R6W5_0),.din(w_dff_A_R16Af9wA2_0),.clk(gclk));
	jdff dff_A_dlri9R6W5_0(.dout(w_dff_A_uXKjIZUZ8_0),.din(w_dff_A_dlri9R6W5_0),.clk(gclk));
	jdff dff_A_uXKjIZUZ8_0(.dout(w_dff_A_ocPFOu4n9_0),.din(w_dff_A_uXKjIZUZ8_0),.clk(gclk));
	jdff dff_A_ocPFOu4n9_0(.dout(w_dff_A_3GNKu7tj4_0),.din(w_dff_A_ocPFOu4n9_0),.clk(gclk));
	jdff dff_A_3GNKu7tj4_0(.dout(w_dff_A_6Klz3CAM9_0),.din(w_dff_A_3GNKu7tj4_0),.clk(gclk));
	jdff dff_A_6Klz3CAM9_0(.dout(w_dff_A_d9dXtT5D1_0),.din(w_dff_A_6Klz3CAM9_0),.clk(gclk));
	jdff dff_A_d9dXtT5D1_0(.dout(w_dff_A_Y45WbqMa1_0),.din(w_dff_A_d9dXtT5D1_0),.clk(gclk));
	jdff dff_A_Y45WbqMa1_0(.dout(w_dff_A_94PULiMl6_0),.din(w_dff_A_Y45WbqMa1_0),.clk(gclk));
	jdff dff_A_94PULiMl6_0(.dout(w_dff_A_VnGbh9Xj3_0),.din(w_dff_A_94PULiMl6_0),.clk(gclk));
	jdff dff_A_VnGbh9Xj3_0(.dout(w_dff_A_wRWZrKDl9_0),.din(w_dff_A_VnGbh9Xj3_0),.clk(gclk));
	jdff dff_A_wRWZrKDl9_0(.dout(w_dff_A_rTm3ETE66_0),.din(w_dff_A_wRWZrKDl9_0),.clk(gclk));
	jdff dff_A_rTm3ETE66_0(.dout(w_dff_A_cMnCFvqz6_0),.din(w_dff_A_rTm3ETE66_0),.clk(gclk));
	jdff dff_A_cMnCFvqz6_0(.dout(w_dff_A_EqIcwaNl4_0),.din(w_dff_A_cMnCFvqz6_0),.clk(gclk));
	jdff dff_A_EqIcwaNl4_0(.dout(w_dff_A_PYTHsVSV6_0),.din(w_dff_A_EqIcwaNl4_0),.clk(gclk));
	jdff dff_A_PYTHsVSV6_0(.dout(w_dff_A_zW3StyU38_0),.din(w_dff_A_PYTHsVSV6_0),.clk(gclk));
	jdff dff_A_zW3StyU38_0(.dout(w_dff_A_TiiRIfM07_0),.din(w_dff_A_zW3StyU38_0),.clk(gclk));
	jdff dff_A_TiiRIfM07_0(.dout(w_dff_A_Z8m1LNur4_0),.din(w_dff_A_TiiRIfM07_0),.clk(gclk));
	jdff dff_A_Z8m1LNur4_0(.dout(w_dff_A_pDxQtBqK4_0),.din(w_dff_A_Z8m1LNur4_0),.clk(gclk));
	jdff dff_A_pDxQtBqK4_0(.dout(w_dff_A_Xxxmtu9M9_0),.din(w_dff_A_pDxQtBqK4_0),.clk(gclk));
	jdff dff_A_Xxxmtu9M9_0(.dout(w_dff_A_v1i21oW54_0),.din(w_dff_A_Xxxmtu9M9_0),.clk(gclk));
	jdff dff_A_v1i21oW54_0(.dout(w_dff_A_Q3nwZ8B10_0),.din(w_dff_A_v1i21oW54_0),.clk(gclk));
	jdff dff_A_Q3nwZ8B10_0(.dout(w_dff_A_SxpUWssj6_0),.din(w_dff_A_Q3nwZ8B10_0),.clk(gclk));
	jdff dff_A_SxpUWssj6_0(.dout(w_dff_A_8oG1HlPz7_0),.din(w_dff_A_SxpUWssj6_0),.clk(gclk));
	jdff dff_A_8oG1HlPz7_0(.dout(w_dff_A_XuZzfXVF6_0),.din(w_dff_A_8oG1HlPz7_0),.clk(gclk));
	jdff dff_A_XuZzfXVF6_0(.dout(w_dff_A_Pwa9WOzs5_0),.din(w_dff_A_XuZzfXVF6_0),.clk(gclk));
	jdff dff_A_Pwa9WOzs5_0(.dout(w_dff_A_PfzGn3X40_0),.din(w_dff_A_Pwa9WOzs5_0),.clk(gclk));
	jdff dff_A_PfzGn3X40_0(.dout(w_dff_A_BfQIop7N9_0),.din(w_dff_A_PfzGn3X40_0),.clk(gclk));
	jdff dff_A_BfQIop7N9_0(.dout(w_dff_A_3Wp3jCBv0_0),.din(w_dff_A_BfQIop7N9_0),.clk(gclk));
	jdff dff_A_3Wp3jCBv0_0(.dout(w_dff_A_zOl2rtiz9_0),.din(w_dff_A_3Wp3jCBv0_0),.clk(gclk));
	jdff dff_A_zOl2rtiz9_0(.dout(w_dff_A_yjXakVSd2_0),.din(w_dff_A_zOl2rtiz9_0),.clk(gclk));
	jdff dff_A_yjXakVSd2_0(.dout(w_dff_A_uAUxLrQH5_0),.din(w_dff_A_yjXakVSd2_0),.clk(gclk));
	jdff dff_A_uAUxLrQH5_0(.dout(w_dff_A_ySqeQT9u0_0),.din(w_dff_A_uAUxLrQH5_0),.clk(gclk));
	jdff dff_A_ySqeQT9u0_0(.dout(w_dff_A_tTPD9ViQ9_0),.din(w_dff_A_ySqeQT9u0_0),.clk(gclk));
	jdff dff_A_tTPD9ViQ9_0(.dout(w_dff_A_S5aMvSkZ1_0),.din(w_dff_A_tTPD9ViQ9_0),.clk(gclk));
	jdff dff_A_S5aMvSkZ1_0(.dout(w_dff_A_Aj89iEXp0_0),.din(w_dff_A_S5aMvSkZ1_0),.clk(gclk));
	jdff dff_A_Aj89iEXp0_0(.dout(w_dff_A_i15bLFzL8_0),.din(w_dff_A_Aj89iEXp0_0),.clk(gclk));
	jdff dff_A_i15bLFzL8_0(.dout(w_dff_A_r47pQr0d3_0),.din(w_dff_A_i15bLFzL8_0),.clk(gclk));
	jdff dff_A_r47pQr0d3_0(.dout(w_dff_A_DcnzQsiz7_0),.din(w_dff_A_r47pQr0d3_0),.clk(gclk));
	jdff dff_A_DcnzQsiz7_0(.dout(w_dff_A_9mk7is8K3_0),.din(w_dff_A_DcnzQsiz7_0),.clk(gclk));
	jdff dff_A_9mk7is8K3_0(.dout(w_dff_A_68phYQ4d9_0),.din(w_dff_A_9mk7is8K3_0),.clk(gclk));
	jdff dff_A_68phYQ4d9_0(.dout(G3211gat),.din(w_dff_A_68phYQ4d9_0),.clk(gclk));
	jdff dff_A_1S7EK9uC0_2(.dout(w_dff_A_HPUO8x400_0),.din(w_dff_A_1S7EK9uC0_2),.clk(gclk));
	jdff dff_A_HPUO8x400_0(.dout(w_dff_A_WC9m3MTH6_0),.din(w_dff_A_HPUO8x400_0),.clk(gclk));
	jdff dff_A_WC9m3MTH6_0(.dout(w_dff_A_yV6upp311_0),.din(w_dff_A_WC9m3MTH6_0),.clk(gclk));
	jdff dff_A_yV6upp311_0(.dout(w_dff_A_NkTNLiv69_0),.din(w_dff_A_yV6upp311_0),.clk(gclk));
	jdff dff_A_NkTNLiv69_0(.dout(w_dff_A_TEWSREFY8_0),.din(w_dff_A_NkTNLiv69_0),.clk(gclk));
	jdff dff_A_TEWSREFY8_0(.dout(w_dff_A_hahDbAXu3_0),.din(w_dff_A_TEWSREFY8_0),.clk(gclk));
	jdff dff_A_hahDbAXu3_0(.dout(w_dff_A_QqVaIVsn3_0),.din(w_dff_A_hahDbAXu3_0),.clk(gclk));
	jdff dff_A_QqVaIVsn3_0(.dout(w_dff_A_kPlYeg6T3_0),.din(w_dff_A_QqVaIVsn3_0),.clk(gclk));
	jdff dff_A_kPlYeg6T3_0(.dout(w_dff_A_88CXVLny9_0),.din(w_dff_A_kPlYeg6T3_0),.clk(gclk));
	jdff dff_A_88CXVLny9_0(.dout(w_dff_A_pln3Ak7p8_0),.din(w_dff_A_88CXVLny9_0),.clk(gclk));
	jdff dff_A_pln3Ak7p8_0(.dout(w_dff_A_C6QyKAcU4_0),.din(w_dff_A_pln3Ak7p8_0),.clk(gclk));
	jdff dff_A_C6QyKAcU4_0(.dout(w_dff_A_V3wRKQ6T0_0),.din(w_dff_A_C6QyKAcU4_0),.clk(gclk));
	jdff dff_A_V3wRKQ6T0_0(.dout(w_dff_A_vspatCTH4_0),.din(w_dff_A_V3wRKQ6T0_0),.clk(gclk));
	jdff dff_A_vspatCTH4_0(.dout(w_dff_A_ONKKmu3q0_0),.din(w_dff_A_vspatCTH4_0),.clk(gclk));
	jdff dff_A_ONKKmu3q0_0(.dout(w_dff_A_dFA43SZV8_0),.din(w_dff_A_ONKKmu3q0_0),.clk(gclk));
	jdff dff_A_dFA43SZV8_0(.dout(w_dff_A_zgdFauPo1_0),.din(w_dff_A_dFA43SZV8_0),.clk(gclk));
	jdff dff_A_zgdFauPo1_0(.dout(w_dff_A_2gmMJMzL1_0),.din(w_dff_A_zgdFauPo1_0),.clk(gclk));
	jdff dff_A_2gmMJMzL1_0(.dout(w_dff_A_V79hsKxC5_0),.din(w_dff_A_2gmMJMzL1_0),.clk(gclk));
	jdff dff_A_V79hsKxC5_0(.dout(w_dff_A_swYR5ZIm2_0),.din(w_dff_A_V79hsKxC5_0),.clk(gclk));
	jdff dff_A_swYR5ZIm2_0(.dout(w_dff_A_1QJpCATX3_0),.din(w_dff_A_swYR5ZIm2_0),.clk(gclk));
	jdff dff_A_1QJpCATX3_0(.dout(w_dff_A_RN94JaGJ7_0),.din(w_dff_A_1QJpCATX3_0),.clk(gclk));
	jdff dff_A_RN94JaGJ7_0(.dout(w_dff_A_UAPm7bfk6_0),.din(w_dff_A_RN94JaGJ7_0),.clk(gclk));
	jdff dff_A_UAPm7bfk6_0(.dout(w_dff_A_rfc8MkMO1_0),.din(w_dff_A_UAPm7bfk6_0),.clk(gclk));
	jdff dff_A_rfc8MkMO1_0(.dout(w_dff_A_8kmJIDCC6_0),.din(w_dff_A_rfc8MkMO1_0),.clk(gclk));
	jdff dff_A_8kmJIDCC6_0(.dout(w_dff_A_vnxznyvI0_0),.din(w_dff_A_8kmJIDCC6_0),.clk(gclk));
	jdff dff_A_vnxznyvI0_0(.dout(w_dff_A_w36IsMES2_0),.din(w_dff_A_vnxznyvI0_0),.clk(gclk));
	jdff dff_A_w36IsMES2_0(.dout(w_dff_A_J0AoCJDc7_0),.din(w_dff_A_w36IsMES2_0),.clk(gclk));
	jdff dff_A_J0AoCJDc7_0(.dout(w_dff_A_GLZ5Xeui5_0),.din(w_dff_A_J0AoCJDc7_0),.clk(gclk));
	jdff dff_A_GLZ5Xeui5_0(.dout(w_dff_A_Wc3AONrK4_0),.din(w_dff_A_GLZ5Xeui5_0),.clk(gclk));
	jdff dff_A_Wc3AONrK4_0(.dout(w_dff_A_DRa0OLxR4_0),.din(w_dff_A_Wc3AONrK4_0),.clk(gclk));
	jdff dff_A_DRa0OLxR4_0(.dout(w_dff_A_btiNppzx2_0),.din(w_dff_A_DRa0OLxR4_0),.clk(gclk));
	jdff dff_A_btiNppzx2_0(.dout(w_dff_A_DFFZ0xWL5_0),.din(w_dff_A_btiNppzx2_0),.clk(gclk));
	jdff dff_A_DFFZ0xWL5_0(.dout(w_dff_A_5xZ55Ezy0_0),.din(w_dff_A_DFFZ0xWL5_0),.clk(gclk));
	jdff dff_A_5xZ55Ezy0_0(.dout(w_dff_A_ubRN5I0d2_0),.din(w_dff_A_5xZ55Ezy0_0),.clk(gclk));
	jdff dff_A_ubRN5I0d2_0(.dout(w_dff_A_48kgtEq73_0),.din(w_dff_A_ubRN5I0d2_0),.clk(gclk));
	jdff dff_A_48kgtEq73_0(.dout(w_dff_A_Mo7K6gIZ5_0),.din(w_dff_A_48kgtEq73_0),.clk(gclk));
	jdff dff_A_Mo7K6gIZ5_0(.dout(w_dff_A_2EloxUDu8_0),.din(w_dff_A_Mo7K6gIZ5_0),.clk(gclk));
	jdff dff_A_2EloxUDu8_0(.dout(w_dff_A_7gmrsr0L6_0),.din(w_dff_A_2EloxUDu8_0),.clk(gclk));
	jdff dff_A_7gmrsr0L6_0(.dout(w_dff_A_BTqd9MWm2_0),.din(w_dff_A_7gmrsr0L6_0),.clk(gclk));
	jdff dff_A_BTqd9MWm2_0(.dout(w_dff_A_XzN1SUH75_0),.din(w_dff_A_BTqd9MWm2_0),.clk(gclk));
	jdff dff_A_XzN1SUH75_0(.dout(w_dff_A_CI30zncL7_0),.din(w_dff_A_XzN1SUH75_0),.clk(gclk));
	jdff dff_A_CI30zncL7_0(.dout(w_dff_A_cTzWC01n7_0),.din(w_dff_A_CI30zncL7_0),.clk(gclk));
	jdff dff_A_cTzWC01n7_0(.dout(w_dff_A_nCyqUpG01_0),.din(w_dff_A_cTzWC01n7_0),.clk(gclk));
	jdff dff_A_nCyqUpG01_0(.dout(w_dff_A_IAwfR51o0_0),.din(w_dff_A_nCyqUpG01_0),.clk(gclk));
	jdff dff_A_IAwfR51o0_0(.dout(w_dff_A_mhy64e4S5_0),.din(w_dff_A_IAwfR51o0_0),.clk(gclk));
	jdff dff_A_mhy64e4S5_0(.dout(w_dff_A_KJnPgomu6_0),.din(w_dff_A_mhy64e4S5_0),.clk(gclk));
	jdff dff_A_KJnPgomu6_0(.dout(w_dff_A_Xhq0SttG8_0),.din(w_dff_A_KJnPgomu6_0),.clk(gclk));
	jdff dff_A_Xhq0SttG8_0(.dout(w_dff_A_7uhaWb3b0_0),.din(w_dff_A_Xhq0SttG8_0),.clk(gclk));
	jdff dff_A_7uhaWb3b0_0(.dout(w_dff_A_c2T70DH62_0),.din(w_dff_A_7uhaWb3b0_0),.clk(gclk));
	jdff dff_A_c2T70DH62_0(.dout(w_dff_A_0NeDqDHN7_0),.din(w_dff_A_c2T70DH62_0),.clk(gclk));
	jdff dff_A_0NeDqDHN7_0(.dout(w_dff_A_N1CbjniU6_0),.din(w_dff_A_0NeDqDHN7_0),.clk(gclk));
	jdff dff_A_N1CbjniU6_0(.dout(w_dff_A_RaSdH8Ma7_0),.din(w_dff_A_N1CbjniU6_0),.clk(gclk));
	jdff dff_A_RaSdH8Ma7_0(.dout(w_dff_A_uZFEBlv00_0),.din(w_dff_A_RaSdH8Ma7_0),.clk(gclk));
	jdff dff_A_uZFEBlv00_0(.dout(G3552gat),.din(w_dff_A_uZFEBlv00_0),.clk(gclk));
	jdff dff_A_fdK3GZD42_2(.dout(w_dff_A_D1ljxla53_0),.din(w_dff_A_fdK3GZD42_2),.clk(gclk));
	jdff dff_A_D1ljxla53_0(.dout(w_dff_A_tEARLD7D6_0),.din(w_dff_A_D1ljxla53_0),.clk(gclk));
	jdff dff_A_tEARLD7D6_0(.dout(w_dff_A_76c5jxDK0_0),.din(w_dff_A_tEARLD7D6_0),.clk(gclk));
	jdff dff_A_76c5jxDK0_0(.dout(w_dff_A_zBD61QgE5_0),.din(w_dff_A_76c5jxDK0_0),.clk(gclk));
	jdff dff_A_zBD61QgE5_0(.dout(w_dff_A_ztwIVD195_0),.din(w_dff_A_zBD61QgE5_0),.clk(gclk));
	jdff dff_A_ztwIVD195_0(.dout(w_dff_A_46XjdZOD8_0),.din(w_dff_A_ztwIVD195_0),.clk(gclk));
	jdff dff_A_46XjdZOD8_0(.dout(w_dff_A_ubCCc7Ut7_0),.din(w_dff_A_46XjdZOD8_0),.clk(gclk));
	jdff dff_A_ubCCc7Ut7_0(.dout(w_dff_A_19AlYVxb6_0),.din(w_dff_A_ubCCc7Ut7_0),.clk(gclk));
	jdff dff_A_19AlYVxb6_0(.dout(w_dff_A_7nhZJRs75_0),.din(w_dff_A_19AlYVxb6_0),.clk(gclk));
	jdff dff_A_7nhZJRs75_0(.dout(w_dff_A_o7mc7g1c8_0),.din(w_dff_A_7nhZJRs75_0),.clk(gclk));
	jdff dff_A_o7mc7g1c8_0(.dout(w_dff_A_PNytZXnZ6_0),.din(w_dff_A_o7mc7g1c8_0),.clk(gclk));
	jdff dff_A_PNytZXnZ6_0(.dout(w_dff_A_pYQCQtA32_0),.din(w_dff_A_PNytZXnZ6_0),.clk(gclk));
	jdff dff_A_pYQCQtA32_0(.dout(w_dff_A_KD3YEOd65_0),.din(w_dff_A_pYQCQtA32_0),.clk(gclk));
	jdff dff_A_KD3YEOd65_0(.dout(w_dff_A_EGwqlcHe5_0),.din(w_dff_A_KD3YEOd65_0),.clk(gclk));
	jdff dff_A_EGwqlcHe5_0(.dout(w_dff_A_EoZBtHPh3_0),.din(w_dff_A_EGwqlcHe5_0),.clk(gclk));
	jdff dff_A_EoZBtHPh3_0(.dout(w_dff_A_AYNaDx281_0),.din(w_dff_A_EoZBtHPh3_0),.clk(gclk));
	jdff dff_A_AYNaDx281_0(.dout(w_dff_A_UMl2PSNY9_0),.din(w_dff_A_AYNaDx281_0),.clk(gclk));
	jdff dff_A_UMl2PSNY9_0(.dout(w_dff_A_MvOEAy0u1_0),.din(w_dff_A_UMl2PSNY9_0),.clk(gclk));
	jdff dff_A_MvOEAy0u1_0(.dout(w_dff_A_5g1JbNwe1_0),.din(w_dff_A_MvOEAy0u1_0),.clk(gclk));
	jdff dff_A_5g1JbNwe1_0(.dout(w_dff_A_UvrOH25s6_0),.din(w_dff_A_5g1JbNwe1_0),.clk(gclk));
	jdff dff_A_UvrOH25s6_0(.dout(w_dff_A_MQ0iiGvh3_0),.din(w_dff_A_UvrOH25s6_0),.clk(gclk));
	jdff dff_A_MQ0iiGvh3_0(.dout(w_dff_A_EDcfrQLi4_0),.din(w_dff_A_MQ0iiGvh3_0),.clk(gclk));
	jdff dff_A_EDcfrQLi4_0(.dout(w_dff_A_pqKVAr1L2_0),.din(w_dff_A_EDcfrQLi4_0),.clk(gclk));
	jdff dff_A_pqKVAr1L2_0(.dout(w_dff_A_h48HmMfn9_0),.din(w_dff_A_pqKVAr1L2_0),.clk(gclk));
	jdff dff_A_h48HmMfn9_0(.dout(w_dff_A_FciaFmtN9_0),.din(w_dff_A_h48HmMfn9_0),.clk(gclk));
	jdff dff_A_FciaFmtN9_0(.dout(w_dff_A_Q3yKlTyM2_0),.din(w_dff_A_FciaFmtN9_0),.clk(gclk));
	jdff dff_A_Q3yKlTyM2_0(.dout(w_dff_A_jyS6FEhA3_0),.din(w_dff_A_Q3yKlTyM2_0),.clk(gclk));
	jdff dff_A_jyS6FEhA3_0(.dout(w_dff_A_c87I8tIR1_0),.din(w_dff_A_jyS6FEhA3_0),.clk(gclk));
	jdff dff_A_c87I8tIR1_0(.dout(w_dff_A_HcoYOmkU1_0),.din(w_dff_A_c87I8tIR1_0),.clk(gclk));
	jdff dff_A_HcoYOmkU1_0(.dout(w_dff_A_dbNCtryU3_0),.din(w_dff_A_HcoYOmkU1_0),.clk(gclk));
	jdff dff_A_dbNCtryU3_0(.dout(w_dff_A_8aYcfREe7_0),.din(w_dff_A_dbNCtryU3_0),.clk(gclk));
	jdff dff_A_8aYcfREe7_0(.dout(w_dff_A_0W8NKevD2_0),.din(w_dff_A_8aYcfREe7_0),.clk(gclk));
	jdff dff_A_0W8NKevD2_0(.dout(w_dff_A_fvZktCYV2_0),.din(w_dff_A_0W8NKevD2_0),.clk(gclk));
	jdff dff_A_fvZktCYV2_0(.dout(w_dff_A_d4PDu5js1_0),.din(w_dff_A_fvZktCYV2_0),.clk(gclk));
	jdff dff_A_d4PDu5js1_0(.dout(w_dff_A_emgBjAc66_0),.din(w_dff_A_d4PDu5js1_0),.clk(gclk));
	jdff dff_A_emgBjAc66_0(.dout(w_dff_A_IcrTRLzk1_0),.din(w_dff_A_emgBjAc66_0),.clk(gclk));
	jdff dff_A_IcrTRLzk1_0(.dout(w_dff_A_EmEDWUDA7_0),.din(w_dff_A_IcrTRLzk1_0),.clk(gclk));
	jdff dff_A_EmEDWUDA7_0(.dout(w_dff_A_ppQja7TY5_0),.din(w_dff_A_EmEDWUDA7_0),.clk(gclk));
	jdff dff_A_ppQja7TY5_0(.dout(w_dff_A_IBxT8tdI5_0),.din(w_dff_A_ppQja7TY5_0),.clk(gclk));
	jdff dff_A_IBxT8tdI5_0(.dout(w_dff_A_fum6iNeP8_0),.din(w_dff_A_IBxT8tdI5_0),.clk(gclk));
	jdff dff_A_fum6iNeP8_0(.dout(w_dff_A_JaRRQPGI6_0),.din(w_dff_A_fum6iNeP8_0),.clk(gclk));
	jdff dff_A_JaRRQPGI6_0(.dout(w_dff_A_q1dML4Pk2_0),.din(w_dff_A_JaRRQPGI6_0),.clk(gclk));
	jdff dff_A_q1dML4Pk2_0(.dout(w_dff_A_2Jk1u5j47_0),.din(w_dff_A_q1dML4Pk2_0),.clk(gclk));
	jdff dff_A_2Jk1u5j47_0(.dout(w_dff_A_PzDEvjIy5_0),.din(w_dff_A_2Jk1u5j47_0),.clk(gclk));
	jdff dff_A_PzDEvjIy5_0(.dout(w_dff_A_IBHNEwXx5_0),.din(w_dff_A_PzDEvjIy5_0),.clk(gclk));
	jdff dff_A_IBHNEwXx5_0(.dout(w_dff_A_ksiK7KtB0_0),.din(w_dff_A_IBHNEwXx5_0),.clk(gclk));
	jdff dff_A_ksiK7KtB0_0(.dout(w_dff_A_nbbZbNnd3_0),.din(w_dff_A_ksiK7KtB0_0),.clk(gclk));
	jdff dff_A_nbbZbNnd3_0(.dout(w_dff_A_cd5jhFgd7_0),.din(w_dff_A_nbbZbNnd3_0),.clk(gclk));
	jdff dff_A_cd5jhFgd7_0(.dout(w_dff_A_yKbQ2N8Z4_0),.din(w_dff_A_cd5jhFgd7_0),.clk(gclk));
	jdff dff_A_yKbQ2N8Z4_0(.dout(w_dff_A_pWkdBPgJ1_0),.din(w_dff_A_yKbQ2N8Z4_0),.clk(gclk));
	jdff dff_A_pWkdBPgJ1_0(.dout(G3895gat),.din(w_dff_A_pWkdBPgJ1_0),.clk(gclk));
	jdff dff_A_rFD3ruyP8_2(.dout(w_dff_A_wCy1wkOG8_0),.din(w_dff_A_rFD3ruyP8_2),.clk(gclk));
	jdff dff_A_wCy1wkOG8_0(.dout(w_dff_A_f8dCr8qN6_0),.din(w_dff_A_wCy1wkOG8_0),.clk(gclk));
	jdff dff_A_f8dCr8qN6_0(.dout(w_dff_A_kG6bMXmL9_0),.din(w_dff_A_f8dCr8qN6_0),.clk(gclk));
	jdff dff_A_kG6bMXmL9_0(.dout(w_dff_A_nE69rSCD7_0),.din(w_dff_A_kG6bMXmL9_0),.clk(gclk));
	jdff dff_A_nE69rSCD7_0(.dout(w_dff_A_liYaWvap4_0),.din(w_dff_A_nE69rSCD7_0),.clk(gclk));
	jdff dff_A_liYaWvap4_0(.dout(w_dff_A_YZwxnTFa8_0),.din(w_dff_A_liYaWvap4_0),.clk(gclk));
	jdff dff_A_YZwxnTFa8_0(.dout(w_dff_A_HYrZCvr05_0),.din(w_dff_A_YZwxnTFa8_0),.clk(gclk));
	jdff dff_A_HYrZCvr05_0(.dout(w_dff_A_H1MTa1pn2_0),.din(w_dff_A_HYrZCvr05_0),.clk(gclk));
	jdff dff_A_H1MTa1pn2_0(.dout(w_dff_A_WJWPnB9Q8_0),.din(w_dff_A_H1MTa1pn2_0),.clk(gclk));
	jdff dff_A_WJWPnB9Q8_0(.dout(w_dff_A_2eYmAzvl3_0),.din(w_dff_A_WJWPnB9Q8_0),.clk(gclk));
	jdff dff_A_2eYmAzvl3_0(.dout(w_dff_A_Lerj2lpD7_0),.din(w_dff_A_2eYmAzvl3_0),.clk(gclk));
	jdff dff_A_Lerj2lpD7_0(.dout(w_dff_A_p8WJsDxe2_0),.din(w_dff_A_Lerj2lpD7_0),.clk(gclk));
	jdff dff_A_p8WJsDxe2_0(.dout(w_dff_A_BtXZHzpo6_0),.din(w_dff_A_p8WJsDxe2_0),.clk(gclk));
	jdff dff_A_BtXZHzpo6_0(.dout(w_dff_A_T2pNZOI31_0),.din(w_dff_A_BtXZHzpo6_0),.clk(gclk));
	jdff dff_A_T2pNZOI31_0(.dout(w_dff_A_S5XawaYp1_0),.din(w_dff_A_T2pNZOI31_0),.clk(gclk));
	jdff dff_A_S5XawaYp1_0(.dout(w_dff_A_AdmSjIPk7_0),.din(w_dff_A_S5XawaYp1_0),.clk(gclk));
	jdff dff_A_AdmSjIPk7_0(.dout(w_dff_A_Rz9JcqBr3_0),.din(w_dff_A_AdmSjIPk7_0),.clk(gclk));
	jdff dff_A_Rz9JcqBr3_0(.dout(w_dff_A_3R3qCcjJ9_0),.din(w_dff_A_Rz9JcqBr3_0),.clk(gclk));
	jdff dff_A_3R3qCcjJ9_0(.dout(w_dff_A_lTAA7f5n6_0),.din(w_dff_A_3R3qCcjJ9_0),.clk(gclk));
	jdff dff_A_lTAA7f5n6_0(.dout(w_dff_A_sfwro9XK1_0),.din(w_dff_A_lTAA7f5n6_0),.clk(gclk));
	jdff dff_A_sfwro9XK1_0(.dout(w_dff_A_OWnu9flQ8_0),.din(w_dff_A_sfwro9XK1_0),.clk(gclk));
	jdff dff_A_OWnu9flQ8_0(.dout(w_dff_A_ueVP981F2_0),.din(w_dff_A_OWnu9flQ8_0),.clk(gclk));
	jdff dff_A_ueVP981F2_0(.dout(w_dff_A_t339kxfb7_0),.din(w_dff_A_ueVP981F2_0),.clk(gclk));
	jdff dff_A_t339kxfb7_0(.dout(w_dff_A_ZcDslSaE2_0),.din(w_dff_A_t339kxfb7_0),.clk(gclk));
	jdff dff_A_ZcDslSaE2_0(.dout(w_dff_A_kIFd3SPK5_0),.din(w_dff_A_ZcDslSaE2_0),.clk(gclk));
	jdff dff_A_kIFd3SPK5_0(.dout(w_dff_A_HtpdOZjk3_0),.din(w_dff_A_kIFd3SPK5_0),.clk(gclk));
	jdff dff_A_HtpdOZjk3_0(.dout(w_dff_A_ffaHNuvX1_0),.din(w_dff_A_HtpdOZjk3_0),.clk(gclk));
	jdff dff_A_ffaHNuvX1_0(.dout(w_dff_A_el1TYYkf6_0),.din(w_dff_A_ffaHNuvX1_0),.clk(gclk));
	jdff dff_A_el1TYYkf6_0(.dout(w_dff_A_VXlBulOn1_0),.din(w_dff_A_el1TYYkf6_0),.clk(gclk));
	jdff dff_A_VXlBulOn1_0(.dout(w_dff_A_ftGxvHZw6_0),.din(w_dff_A_VXlBulOn1_0),.clk(gclk));
	jdff dff_A_ftGxvHZw6_0(.dout(w_dff_A_jVvIQzwF0_0),.din(w_dff_A_ftGxvHZw6_0),.clk(gclk));
	jdff dff_A_jVvIQzwF0_0(.dout(w_dff_A_fnJRMVzh6_0),.din(w_dff_A_jVvIQzwF0_0),.clk(gclk));
	jdff dff_A_fnJRMVzh6_0(.dout(w_dff_A_fioCgruU3_0),.din(w_dff_A_fnJRMVzh6_0),.clk(gclk));
	jdff dff_A_fioCgruU3_0(.dout(w_dff_A_HcBfl0mh6_0),.din(w_dff_A_fioCgruU3_0),.clk(gclk));
	jdff dff_A_HcBfl0mh6_0(.dout(w_dff_A_hBewRon32_0),.din(w_dff_A_HcBfl0mh6_0),.clk(gclk));
	jdff dff_A_hBewRon32_0(.dout(w_dff_A_46sTgkrF7_0),.din(w_dff_A_hBewRon32_0),.clk(gclk));
	jdff dff_A_46sTgkrF7_0(.dout(w_dff_A_ahm8CCsf0_0),.din(w_dff_A_46sTgkrF7_0),.clk(gclk));
	jdff dff_A_ahm8CCsf0_0(.dout(w_dff_A_SitAz65p3_0),.din(w_dff_A_ahm8CCsf0_0),.clk(gclk));
	jdff dff_A_SitAz65p3_0(.dout(w_dff_A_wuCqWLwH1_0),.din(w_dff_A_SitAz65p3_0),.clk(gclk));
	jdff dff_A_wuCqWLwH1_0(.dout(w_dff_A_1OeTwyEH9_0),.din(w_dff_A_wuCqWLwH1_0),.clk(gclk));
	jdff dff_A_1OeTwyEH9_0(.dout(w_dff_A_jWvUl0xN3_0),.din(w_dff_A_1OeTwyEH9_0),.clk(gclk));
	jdff dff_A_jWvUl0xN3_0(.dout(w_dff_A_v0BdXfzU6_0),.din(w_dff_A_jWvUl0xN3_0),.clk(gclk));
	jdff dff_A_v0BdXfzU6_0(.dout(w_dff_A_yFAQckSv6_0),.din(w_dff_A_v0BdXfzU6_0),.clk(gclk));
	jdff dff_A_yFAQckSv6_0(.dout(w_dff_A_KXkzmyTm3_0),.din(w_dff_A_yFAQckSv6_0),.clk(gclk));
	jdff dff_A_KXkzmyTm3_0(.dout(w_dff_A_LXNOeWHW9_0),.din(w_dff_A_KXkzmyTm3_0),.clk(gclk));
	jdff dff_A_LXNOeWHW9_0(.dout(w_dff_A_YFPYsXl46_0),.din(w_dff_A_LXNOeWHW9_0),.clk(gclk));
	jdff dff_A_YFPYsXl46_0(.dout(w_dff_A_HLXQTx3j8_0),.din(w_dff_A_YFPYsXl46_0),.clk(gclk));
	jdff dff_A_HLXQTx3j8_0(.dout(G4241gat),.din(w_dff_A_HLXQTx3j8_0),.clk(gclk));
	jdff dff_A_xANsDdVz6_2(.dout(w_dff_A_pXTROB3q9_0),.din(w_dff_A_xANsDdVz6_2),.clk(gclk));
	jdff dff_A_pXTROB3q9_0(.dout(w_dff_A_jTOenI3v4_0),.din(w_dff_A_pXTROB3q9_0),.clk(gclk));
	jdff dff_A_jTOenI3v4_0(.dout(w_dff_A_r8okHQLl2_0),.din(w_dff_A_jTOenI3v4_0),.clk(gclk));
	jdff dff_A_r8okHQLl2_0(.dout(w_dff_A_fM681KaE7_0),.din(w_dff_A_r8okHQLl2_0),.clk(gclk));
	jdff dff_A_fM681KaE7_0(.dout(w_dff_A_jHmMc3Ki1_0),.din(w_dff_A_fM681KaE7_0),.clk(gclk));
	jdff dff_A_jHmMc3Ki1_0(.dout(w_dff_A_fLjFoE160_0),.din(w_dff_A_jHmMc3Ki1_0),.clk(gclk));
	jdff dff_A_fLjFoE160_0(.dout(w_dff_A_h0g5HjaA9_0),.din(w_dff_A_fLjFoE160_0),.clk(gclk));
	jdff dff_A_h0g5HjaA9_0(.dout(w_dff_A_aS2bhrfJ1_0),.din(w_dff_A_h0g5HjaA9_0),.clk(gclk));
	jdff dff_A_aS2bhrfJ1_0(.dout(w_dff_A_GL7PML9S7_0),.din(w_dff_A_aS2bhrfJ1_0),.clk(gclk));
	jdff dff_A_GL7PML9S7_0(.dout(w_dff_A_obzNNO2M9_0),.din(w_dff_A_GL7PML9S7_0),.clk(gclk));
	jdff dff_A_obzNNO2M9_0(.dout(w_dff_A_rC9QR0lC5_0),.din(w_dff_A_obzNNO2M9_0),.clk(gclk));
	jdff dff_A_rC9QR0lC5_0(.dout(w_dff_A_G3oFA62V3_0),.din(w_dff_A_rC9QR0lC5_0),.clk(gclk));
	jdff dff_A_G3oFA62V3_0(.dout(w_dff_A_gPMwZevJ4_0),.din(w_dff_A_G3oFA62V3_0),.clk(gclk));
	jdff dff_A_gPMwZevJ4_0(.dout(w_dff_A_Ahq83ELf3_0),.din(w_dff_A_gPMwZevJ4_0),.clk(gclk));
	jdff dff_A_Ahq83ELf3_0(.dout(w_dff_A_3Gxy1OxP4_0),.din(w_dff_A_Ahq83ELf3_0),.clk(gclk));
	jdff dff_A_3Gxy1OxP4_0(.dout(w_dff_A_tsng1w7b9_0),.din(w_dff_A_3Gxy1OxP4_0),.clk(gclk));
	jdff dff_A_tsng1w7b9_0(.dout(w_dff_A_e9OojFyN1_0),.din(w_dff_A_tsng1w7b9_0),.clk(gclk));
	jdff dff_A_e9OojFyN1_0(.dout(w_dff_A_lhRRBONw1_0),.din(w_dff_A_e9OojFyN1_0),.clk(gclk));
	jdff dff_A_lhRRBONw1_0(.dout(w_dff_A_9K9WqwCv8_0),.din(w_dff_A_lhRRBONw1_0),.clk(gclk));
	jdff dff_A_9K9WqwCv8_0(.dout(w_dff_A_JQlLSURC0_0),.din(w_dff_A_9K9WqwCv8_0),.clk(gclk));
	jdff dff_A_JQlLSURC0_0(.dout(w_dff_A_fQm5pxXj3_0),.din(w_dff_A_JQlLSURC0_0),.clk(gclk));
	jdff dff_A_fQm5pxXj3_0(.dout(w_dff_A_jgkdZ4zw3_0),.din(w_dff_A_fQm5pxXj3_0),.clk(gclk));
	jdff dff_A_jgkdZ4zw3_0(.dout(w_dff_A_2UBEBqK12_0),.din(w_dff_A_jgkdZ4zw3_0),.clk(gclk));
	jdff dff_A_2UBEBqK12_0(.dout(w_dff_A_TECjVfwv6_0),.din(w_dff_A_2UBEBqK12_0),.clk(gclk));
	jdff dff_A_TECjVfwv6_0(.dout(w_dff_A_nSqJEH3d4_0),.din(w_dff_A_TECjVfwv6_0),.clk(gclk));
	jdff dff_A_nSqJEH3d4_0(.dout(w_dff_A_SN8bqs2Q8_0),.din(w_dff_A_nSqJEH3d4_0),.clk(gclk));
	jdff dff_A_SN8bqs2Q8_0(.dout(w_dff_A_T5LinO5h6_0),.din(w_dff_A_SN8bqs2Q8_0),.clk(gclk));
	jdff dff_A_T5LinO5h6_0(.dout(w_dff_A_IM87GUaO0_0),.din(w_dff_A_T5LinO5h6_0),.clk(gclk));
	jdff dff_A_IM87GUaO0_0(.dout(w_dff_A_FySOt3Ij6_0),.din(w_dff_A_IM87GUaO0_0),.clk(gclk));
	jdff dff_A_FySOt3Ij6_0(.dout(w_dff_A_Sid51fXI9_0),.din(w_dff_A_FySOt3Ij6_0),.clk(gclk));
	jdff dff_A_Sid51fXI9_0(.dout(w_dff_A_tcKMdUFV7_0),.din(w_dff_A_Sid51fXI9_0),.clk(gclk));
	jdff dff_A_tcKMdUFV7_0(.dout(w_dff_A_Z1MctO2O6_0),.din(w_dff_A_tcKMdUFV7_0),.clk(gclk));
	jdff dff_A_Z1MctO2O6_0(.dout(w_dff_A_RIlCVX171_0),.din(w_dff_A_Z1MctO2O6_0),.clk(gclk));
	jdff dff_A_RIlCVX171_0(.dout(w_dff_A_y0kfxqN95_0),.din(w_dff_A_RIlCVX171_0),.clk(gclk));
	jdff dff_A_y0kfxqN95_0(.dout(w_dff_A_YZlIMUAR2_0),.din(w_dff_A_y0kfxqN95_0),.clk(gclk));
	jdff dff_A_YZlIMUAR2_0(.dout(w_dff_A_uMQoYzc75_0),.din(w_dff_A_YZlIMUAR2_0),.clk(gclk));
	jdff dff_A_uMQoYzc75_0(.dout(w_dff_A_ATFtiSAo6_0),.din(w_dff_A_uMQoYzc75_0),.clk(gclk));
	jdff dff_A_ATFtiSAo6_0(.dout(w_dff_A_9vqiQXsy9_0),.din(w_dff_A_ATFtiSAo6_0),.clk(gclk));
	jdff dff_A_9vqiQXsy9_0(.dout(w_dff_A_B3kiD3K41_0),.din(w_dff_A_9vqiQXsy9_0),.clk(gclk));
	jdff dff_A_B3kiD3K41_0(.dout(w_dff_A_J7KP6UIZ4_0),.din(w_dff_A_B3kiD3K41_0),.clk(gclk));
	jdff dff_A_J7KP6UIZ4_0(.dout(w_dff_A_KlfMuHA29_0),.din(w_dff_A_J7KP6UIZ4_0),.clk(gclk));
	jdff dff_A_KlfMuHA29_0(.dout(w_dff_A_pIiXC78S0_0),.din(w_dff_A_KlfMuHA29_0),.clk(gclk));
	jdff dff_A_pIiXC78S0_0(.dout(w_dff_A_uHFALARi1_0),.din(w_dff_A_pIiXC78S0_0),.clk(gclk));
	jdff dff_A_uHFALARi1_0(.dout(w_dff_A_sCnUazWe3_0),.din(w_dff_A_uHFALARi1_0),.clk(gclk));
	jdff dff_A_sCnUazWe3_0(.dout(G4591gat),.din(w_dff_A_sCnUazWe3_0),.clk(gclk));
	jdff dff_A_k3iKXLIe4_2(.dout(w_dff_A_Aglkn81E6_0),.din(w_dff_A_k3iKXLIe4_2),.clk(gclk));
	jdff dff_A_Aglkn81E6_0(.dout(w_dff_A_XL6evCQi0_0),.din(w_dff_A_Aglkn81E6_0),.clk(gclk));
	jdff dff_A_XL6evCQi0_0(.dout(w_dff_A_u11dQkLr8_0),.din(w_dff_A_XL6evCQi0_0),.clk(gclk));
	jdff dff_A_u11dQkLr8_0(.dout(w_dff_A_XnWeIXQY3_0),.din(w_dff_A_u11dQkLr8_0),.clk(gclk));
	jdff dff_A_XnWeIXQY3_0(.dout(w_dff_A_VZNs2JDX5_0),.din(w_dff_A_XnWeIXQY3_0),.clk(gclk));
	jdff dff_A_VZNs2JDX5_0(.dout(w_dff_A_6aVrzrep2_0),.din(w_dff_A_VZNs2JDX5_0),.clk(gclk));
	jdff dff_A_6aVrzrep2_0(.dout(w_dff_A_ljf05tGS0_0),.din(w_dff_A_6aVrzrep2_0),.clk(gclk));
	jdff dff_A_ljf05tGS0_0(.dout(w_dff_A_UrPv5nGB4_0),.din(w_dff_A_ljf05tGS0_0),.clk(gclk));
	jdff dff_A_UrPv5nGB4_0(.dout(w_dff_A_5VnNimcs2_0),.din(w_dff_A_UrPv5nGB4_0),.clk(gclk));
	jdff dff_A_5VnNimcs2_0(.dout(w_dff_A_Hrg1rnYa5_0),.din(w_dff_A_5VnNimcs2_0),.clk(gclk));
	jdff dff_A_Hrg1rnYa5_0(.dout(w_dff_A_QcnA24mZ2_0),.din(w_dff_A_Hrg1rnYa5_0),.clk(gclk));
	jdff dff_A_QcnA24mZ2_0(.dout(w_dff_A_J2rQYll28_0),.din(w_dff_A_QcnA24mZ2_0),.clk(gclk));
	jdff dff_A_J2rQYll28_0(.dout(w_dff_A_n7I5sYsL8_0),.din(w_dff_A_J2rQYll28_0),.clk(gclk));
	jdff dff_A_n7I5sYsL8_0(.dout(w_dff_A_S9hkccD34_0),.din(w_dff_A_n7I5sYsL8_0),.clk(gclk));
	jdff dff_A_S9hkccD34_0(.dout(w_dff_A_lpelPjES3_0),.din(w_dff_A_S9hkccD34_0),.clk(gclk));
	jdff dff_A_lpelPjES3_0(.dout(w_dff_A_YzZJmEw44_0),.din(w_dff_A_lpelPjES3_0),.clk(gclk));
	jdff dff_A_YzZJmEw44_0(.dout(w_dff_A_9lcWTbCJ1_0),.din(w_dff_A_YzZJmEw44_0),.clk(gclk));
	jdff dff_A_9lcWTbCJ1_0(.dout(w_dff_A_Ov99oSIH4_0),.din(w_dff_A_9lcWTbCJ1_0),.clk(gclk));
	jdff dff_A_Ov99oSIH4_0(.dout(w_dff_A_D0caj4ux5_0),.din(w_dff_A_Ov99oSIH4_0),.clk(gclk));
	jdff dff_A_D0caj4ux5_0(.dout(w_dff_A_bsshSqi58_0),.din(w_dff_A_D0caj4ux5_0),.clk(gclk));
	jdff dff_A_bsshSqi58_0(.dout(w_dff_A_Nda5H63m0_0),.din(w_dff_A_bsshSqi58_0),.clk(gclk));
	jdff dff_A_Nda5H63m0_0(.dout(w_dff_A_buRSM4VA9_0),.din(w_dff_A_Nda5H63m0_0),.clk(gclk));
	jdff dff_A_buRSM4VA9_0(.dout(w_dff_A_HePwnezM4_0),.din(w_dff_A_buRSM4VA9_0),.clk(gclk));
	jdff dff_A_HePwnezM4_0(.dout(w_dff_A_gc1VAXFE5_0),.din(w_dff_A_HePwnezM4_0),.clk(gclk));
	jdff dff_A_gc1VAXFE5_0(.dout(w_dff_A_fgwJtztX6_0),.din(w_dff_A_gc1VAXFE5_0),.clk(gclk));
	jdff dff_A_fgwJtztX6_0(.dout(w_dff_A_l2OkezNQ1_0),.din(w_dff_A_fgwJtztX6_0),.clk(gclk));
	jdff dff_A_l2OkezNQ1_0(.dout(w_dff_A_V4m9BGio9_0),.din(w_dff_A_l2OkezNQ1_0),.clk(gclk));
	jdff dff_A_V4m9BGio9_0(.dout(w_dff_A_WoDYBINQ3_0),.din(w_dff_A_V4m9BGio9_0),.clk(gclk));
	jdff dff_A_WoDYBINQ3_0(.dout(w_dff_A_RwfZcAnT6_0),.din(w_dff_A_WoDYBINQ3_0),.clk(gclk));
	jdff dff_A_RwfZcAnT6_0(.dout(w_dff_A_iervmNT84_0),.din(w_dff_A_RwfZcAnT6_0),.clk(gclk));
	jdff dff_A_iervmNT84_0(.dout(w_dff_A_sbxqpdEo3_0),.din(w_dff_A_iervmNT84_0),.clk(gclk));
	jdff dff_A_sbxqpdEo3_0(.dout(w_dff_A_Lw05cSSz2_0),.din(w_dff_A_sbxqpdEo3_0),.clk(gclk));
	jdff dff_A_Lw05cSSz2_0(.dout(w_dff_A_GmhKQyBS2_0),.din(w_dff_A_Lw05cSSz2_0),.clk(gclk));
	jdff dff_A_GmhKQyBS2_0(.dout(w_dff_A_8zV5OEf07_0),.din(w_dff_A_GmhKQyBS2_0),.clk(gclk));
	jdff dff_A_8zV5OEf07_0(.dout(w_dff_A_77moib451_0),.din(w_dff_A_8zV5OEf07_0),.clk(gclk));
	jdff dff_A_77moib451_0(.dout(w_dff_A_DOBWTF6i9_0),.din(w_dff_A_77moib451_0),.clk(gclk));
	jdff dff_A_DOBWTF6i9_0(.dout(w_dff_A_JODvmQXA8_0),.din(w_dff_A_DOBWTF6i9_0),.clk(gclk));
	jdff dff_A_JODvmQXA8_0(.dout(w_dff_A_J58U6LNq4_0),.din(w_dff_A_JODvmQXA8_0),.clk(gclk));
	jdff dff_A_J58U6LNq4_0(.dout(w_dff_A_0SptStsj3_0),.din(w_dff_A_J58U6LNq4_0),.clk(gclk));
	jdff dff_A_0SptStsj3_0(.dout(w_dff_A_CXuqsHmV8_0),.din(w_dff_A_0SptStsj3_0),.clk(gclk));
	jdff dff_A_CXuqsHmV8_0(.dout(w_dff_A_akbihhF17_0),.din(w_dff_A_CXuqsHmV8_0),.clk(gclk));
	jdff dff_A_akbihhF17_0(.dout(G4946gat),.din(w_dff_A_akbihhF17_0),.clk(gclk));
	jdff dff_A_Whz6y90z4_2(.dout(w_dff_A_HZt5ri3T9_0),.din(w_dff_A_Whz6y90z4_2),.clk(gclk));
	jdff dff_A_HZt5ri3T9_0(.dout(w_dff_A_MjSvTIG88_0),.din(w_dff_A_HZt5ri3T9_0),.clk(gclk));
	jdff dff_A_MjSvTIG88_0(.dout(w_dff_A_JrxqGUmX7_0),.din(w_dff_A_MjSvTIG88_0),.clk(gclk));
	jdff dff_A_JrxqGUmX7_0(.dout(w_dff_A_42z0BhHr9_0),.din(w_dff_A_JrxqGUmX7_0),.clk(gclk));
	jdff dff_A_42z0BhHr9_0(.dout(w_dff_A_WA9QuyfT8_0),.din(w_dff_A_42z0BhHr9_0),.clk(gclk));
	jdff dff_A_WA9QuyfT8_0(.dout(w_dff_A_hV3B999W1_0),.din(w_dff_A_WA9QuyfT8_0),.clk(gclk));
	jdff dff_A_hV3B999W1_0(.dout(w_dff_A_yw5RLx8R4_0),.din(w_dff_A_hV3B999W1_0),.clk(gclk));
	jdff dff_A_yw5RLx8R4_0(.dout(w_dff_A_GlRNSy3p5_0),.din(w_dff_A_yw5RLx8R4_0),.clk(gclk));
	jdff dff_A_GlRNSy3p5_0(.dout(w_dff_A_Ifjcdlbu3_0),.din(w_dff_A_GlRNSy3p5_0),.clk(gclk));
	jdff dff_A_Ifjcdlbu3_0(.dout(w_dff_A_sSoUT4GB2_0),.din(w_dff_A_Ifjcdlbu3_0),.clk(gclk));
	jdff dff_A_sSoUT4GB2_0(.dout(w_dff_A_7z4bE0cu6_0),.din(w_dff_A_sSoUT4GB2_0),.clk(gclk));
	jdff dff_A_7z4bE0cu6_0(.dout(w_dff_A_fBj8Bayd6_0),.din(w_dff_A_7z4bE0cu6_0),.clk(gclk));
	jdff dff_A_fBj8Bayd6_0(.dout(w_dff_A_ARnkUL2z7_0),.din(w_dff_A_fBj8Bayd6_0),.clk(gclk));
	jdff dff_A_ARnkUL2z7_0(.dout(w_dff_A_phchnPF09_0),.din(w_dff_A_ARnkUL2z7_0),.clk(gclk));
	jdff dff_A_phchnPF09_0(.dout(w_dff_A_AbD197dt4_0),.din(w_dff_A_phchnPF09_0),.clk(gclk));
	jdff dff_A_AbD197dt4_0(.dout(w_dff_A_qZU0jvS74_0),.din(w_dff_A_AbD197dt4_0),.clk(gclk));
	jdff dff_A_qZU0jvS74_0(.dout(w_dff_A_AC60Ks0n6_0),.din(w_dff_A_qZU0jvS74_0),.clk(gclk));
	jdff dff_A_AC60Ks0n6_0(.dout(w_dff_A_zowmw9a57_0),.din(w_dff_A_AC60Ks0n6_0),.clk(gclk));
	jdff dff_A_zowmw9a57_0(.dout(w_dff_A_fwwJw1VS2_0),.din(w_dff_A_zowmw9a57_0),.clk(gclk));
	jdff dff_A_fwwJw1VS2_0(.dout(w_dff_A_8Kb0HGMS8_0),.din(w_dff_A_fwwJw1VS2_0),.clk(gclk));
	jdff dff_A_8Kb0HGMS8_0(.dout(w_dff_A_GawTFX1o1_0),.din(w_dff_A_8Kb0HGMS8_0),.clk(gclk));
	jdff dff_A_GawTFX1o1_0(.dout(w_dff_A_1QWCMiNR1_0),.din(w_dff_A_GawTFX1o1_0),.clk(gclk));
	jdff dff_A_1QWCMiNR1_0(.dout(w_dff_A_jCTNTG1a6_0),.din(w_dff_A_1QWCMiNR1_0),.clk(gclk));
	jdff dff_A_jCTNTG1a6_0(.dout(w_dff_A_KI8nbasE7_0),.din(w_dff_A_jCTNTG1a6_0),.clk(gclk));
	jdff dff_A_KI8nbasE7_0(.dout(w_dff_A_wRVKJ3jY9_0),.din(w_dff_A_KI8nbasE7_0),.clk(gclk));
	jdff dff_A_wRVKJ3jY9_0(.dout(w_dff_A_4k8yGm471_0),.din(w_dff_A_wRVKJ3jY9_0),.clk(gclk));
	jdff dff_A_4k8yGm471_0(.dout(w_dff_A_dYamHiU94_0),.din(w_dff_A_4k8yGm471_0),.clk(gclk));
	jdff dff_A_dYamHiU94_0(.dout(w_dff_A_Hb5cXusa5_0),.din(w_dff_A_dYamHiU94_0),.clk(gclk));
	jdff dff_A_Hb5cXusa5_0(.dout(w_dff_A_EGGfkYTS7_0),.din(w_dff_A_Hb5cXusa5_0),.clk(gclk));
	jdff dff_A_EGGfkYTS7_0(.dout(w_dff_A_T5g9g3CF7_0),.din(w_dff_A_EGGfkYTS7_0),.clk(gclk));
	jdff dff_A_T5g9g3CF7_0(.dout(w_dff_A_BPTIuZLw0_0),.din(w_dff_A_T5g9g3CF7_0),.clk(gclk));
	jdff dff_A_BPTIuZLw0_0(.dout(w_dff_A_CYdXihWS8_0),.din(w_dff_A_BPTIuZLw0_0),.clk(gclk));
	jdff dff_A_CYdXihWS8_0(.dout(w_dff_A_JfbYWNPY1_0),.din(w_dff_A_CYdXihWS8_0),.clk(gclk));
	jdff dff_A_JfbYWNPY1_0(.dout(w_dff_A_uYc1LZQA9_0),.din(w_dff_A_JfbYWNPY1_0),.clk(gclk));
	jdff dff_A_uYc1LZQA9_0(.dout(w_dff_A_5JzA5IOY5_0),.din(w_dff_A_uYc1LZQA9_0),.clk(gclk));
	jdff dff_A_5JzA5IOY5_0(.dout(w_dff_A_zlYlzgot0_0),.din(w_dff_A_5JzA5IOY5_0),.clk(gclk));
	jdff dff_A_zlYlzgot0_0(.dout(w_dff_A_J77gEn0R7_0),.din(w_dff_A_zlYlzgot0_0),.clk(gclk));
	jdff dff_A_J77gEn0R7_0(.dout(w_dff_A_IOeZXjCa0_0),.din(w_dff_A_J77gEn0R7_0),.clk(gclk));
	jdff dff_A_IOeZXjCa0_0(.dout(G5308gat),.din(w_dff_A_IOeZXjCa0_0),.clk(gclk));
	jdff dff_A_dSuBmHpc5_2(.dout(w_dff_A_mdoLfKW24_0),.din(w_dff_A_dSuBmHpc5_2),.clk(gclk));
	jdff dff_A_mdoLfKW24_0(.dout(w_dff_A_fdPLxgoC7_0),.din(w_dff_A_mdoLfKW24_0),.clk(gclk));
	jdff dff_A_fdPLxgoC7_0(.dout(w_dff_A_p0IlcEKG9_0),.din(w_dff_A_fdPLxgoC7_0),.clk(gclk));
	jdff dff_A_p0IlcEKG9_0(.dout(w_dff_A_3Pq8IOer9_0),.din(w_dff_A_p0IlcEKG9_0),.clk(gclk));
	jdff dff_A_3Pq8IOer9_0(.dout(w_dff_A_EopLJP5f8_0),.din(w_dff_A_3Pq8IOer9_0),.clk(gclk));
	jdff dff_A_EopLJP5f8_0(.dout(w_dff_A_aZpy6ceA4_0),.din(w_dff_A_EopLJP5f8_0),.clk(gclk));
	jdff dff_A_aZpy6ceA4_0(.dout(w_dff_A_u2yetZ701_0),.din(w_dff_A_aZpy6ceA4_0),.clk(gclk));
	jdff dff_A_u2yetZ701_0(.dout(w_dff_A_XRjeNN6X4_0),.din(w_dff_A_u2yetZ701_0),.clk(gclk));
	jdff dff_A_XRjeNN6X4_0(.dout(w_dff_A_J9I248Jp1_0),.din(w_dff_A_XRjeNN6X4_0),.clk(gclk));
	jdff dff_A_J9I248Jp1_0(.dout(w_dff_A_htZXRUfj3_0),.din(w_dff_A_J9I248Jp1_0),.clk(gclk));
	jdff dff_A_htZXRUfj3_0(.dout(w_dff_A_U4JsR3Uq9_0),.din(w_dff_A_htZXRUfj3_0),.clk(gclk));
	jdff dff_A_U4JsR3Uq9_0(.dout(w_dff_A_p6E1KrtO2_0),.din(w_dff_A_U4JsR3Uq9_0),.clk(gclk));
	jdff dff_A_p6E1KrtO2_0(.dout(w_dff_A_Q1tb5loz6_0),.din(w_dff_A_p6E1KrtO2_0),.clk(gclk));
	jdff dff_A_Q1tb5loz6_0(.dout(w_dff_A_h2AvVCpa7_0),.din(w_dff_A_Q1tb5loz6_0),.clk(gclk));
	jdff dff_A_h2AvVCpa7_0(.dout(w_dff_A_bzvuPIrZ7_0),.din(w_dff_A_h2AvVCpa7_0),.clk(gclk));
	jdff dff_A_bzvuPIrZ7_0(.dout(w_dff_A_yy7jIqcN3_0),.din(w_dff_A_bzvuPIrZ7_0),.clk(gclk));
	jdff dff_A_yy7jIqcN3_0(.dout(w_dff_A_JlQ5wT8n6_0),.din(w_dff_A_yy7jIqcN3_0),.clk(gclk));
	jdff dff_A_JlQ5wT8n6_0(.dout(w_dff_A_yxNV3cxa8_0),.din(w_dff_A_JlQ5wT8n6_0),.clk(gclk));
	jdff dff_A_yxNV3cxa8_0(.dout(w_dff_A_9VucbSb85_0),.din(w_dff_A_yxNV3cxa8_0),.clk(gclk));
	jdff dff_A_9VucbSb85_0(.dout(w_dff_A_s7UaRNx12_0),.din(w_dff_A_9VucbSb85_0),.clk(gclk));
	jdff dff_A_s7UaRNx12_0(.dout(w_dff_A_9shebP5b4_0),.din(w_dff_A_s7UaRNx12_0),.clk(gclk));
	jdff dff_A_9shebP5b4_0(.dout(w_dff_A_BphnsUee2_0),.din(w_dff_A_9shebP5b4_0),.clk(gclk));
	jdff dff_A_BphnsUee2_0(.dout(w_dff_A_7MN3KpQd6_0),.din(w_dff_A_BphnsUee2_0),.clk(gclk));
	jdff dff_A_7MN3KpQd6_0(.dout(w_dff_A_vw1RV2NV0_0),.din(w_dff_A_7MN3KpQd6_0),.clk(gclk));
	jdff dff_A_vw1RV2NV0_0(.dout(w_dff_A_SHwyh0c18_0),.din(w_dff_A_vw1RV2NV0_0),.clk(gclk));
	jdff dff_A_SHwyh0c18_0(.dout(w_dff_A_DDAQjcyZ1_0),.din(w_dff_A_SHwyh0c18_0),.clk(gclk));
	jdff dff_A_DDAQjcyZ1_0(.dout(w_dff_A_Dg9NJat15_0),.din(w_dff_A_DDAQjcyZ1_0),.clk(gclk));
	jdff dff_A_Dg9NJat15_0(.dout(w_dff_A_2CJ6JoJ82_0),.din(w_dff_A_Dg9NJat15_0),.clk(gclk));
	jdff dff_A_2CJ6JoJ82_0(.dout(w_dff_A_cJ2U47NJ9_0),.din(w_dff_A_2CJ6JoJ82_0),.clk(gclk));
	jdff dff_A_cJ2U47NJ9_0(.dout(w_dff_A_w16I4wIA3_0),.din(w_dff_A_cJ2U47NJ9_0),.clk(gclk));
	jdff dff_A_w16I4wIA3_0(.dout(w_dff_A_zwpytITb0_0),.din(w_dff_A_w16I4wIA3_0),.clk(gclk));
	jdff dff_A_zwpytITb0_0(.dout(w_dff_A_EgeqZIwH2_0),.din(w_dff_A_zwpytITb0_0),.clk(gclk));
	jdff dff_A_EgeqZIwH2_0(.dout(w_dff_A_tjFBlMny9_0),.din(w_dff_A_EgeqZIwH2_0),.clk(gclk));
	jdff dff_A_tjFBlMny9_0(.dout(w_dff_A_iKzjfTVX4_0),.din(w_dff_A_tjFBlMny9_0),.clk(gclk));
	jdff dff_A_iKzjfTVX4_0(.dout(w_dff_A_6VkxC2es4_0),.din(w_dff_A_iKzjfTVX4_0),.clk(gclk));
	jdff dff_A_6VkxC2es4_0(.dout(G5672gat),.din(w_dff_A_6VkxC2es4_0),.clk(gclk));
	jdff dff_A_GrvPvRzD1_2(.dout(w_dff_A_pqB8Fko46_0),.din(w_dff_A_GrvPvRzD1_2),.clk(gclk));
	jdff dff_A_pqB8Fko46_0(.dout(w_dff_A_3f80n6Gs2_0),.din(w_dff_A_pqB8Fko46_0),.clk(gclk));
	jdff dff_A_3f80n6Gs2_0(.dout(w_dff_A_Udra6jHd0_0),.din(w_dff_A_3f80n6Gs2_0),.clk(gclk));
	jdff dff_A_Udra6jHd0_0(.dout(w_dff_A_034Fj5gR5_0),.din(w_dff_A_Udra6jHd0_0),.clk(gclk));
	jdff dff_A_034Fj5gR5_0(.dout(w_dff_A_we1nG2fK9_0),.din(w_dff_A_034Fj5gR5_0),.clk(gclk));
	jdff dff_A_we1nG2fK9_0(.dout(w_dff_A_8uBpOEXy0_0),.din(w_dff_A_we1nG2fK9_0),.clk(gclk));
	jdff dff_A_8uBpOEXy0_0(.dout(w_dff_A_AFM0uJ5l6_0),.din(w_dff_A_8uBpOEXy0_0),.clk(gclk));
	jdff dff_A_AFM0uJ5l6_0(.dout(w_dff_A_tqQXvXDU0_0),.din(w_dff_A_AFM0uJ5l6_0),.clk(gclk));
	jdff dff_A_tqQXvXDU0_0(.dout(w_dff_A_w1ApzctC7_0),.din(w_dff_A_tqQXvXDU0_0),.clk(gclk));
	jdff dff_A_w1ApzctC7_0(.dout(w_dff_A_ztgUPg7q4_0),.din(w_dff_A_w1ApzctC7_0),.clk(gclk));
	jdff dff_A_ztgUPg7q4_0(.dout(w_dff_A_XwcQiECs5_0),.din(w_dff_A_ztgUPg7q4_0),.clk(gclk));
	jdff dff_A_XwcQiECs5_0(.dout(w_dff_A_vvzIJkBd2_0),.din(w_dff_A_XwcQiECs5_0),.clk(gclk));
	jdff dff_A_vvzIJkBd2_0(.dout(w_dff_A_ujjTKTyt5_0),.din(w_dff_A_vvzIJkBd2_0),.clk(gclk));
	jdff dff_A_ujjTKTyt5_0(.dout(w_dff_A_0To7aDDQ0_0),.din(w_dff_A_ujjTKTyt5_0),.clk(gclk));
	jdff dff_A_0To7aDDQ0_0(.dout(w_dff_A_PNOJfyzw4_0),.din(w_dff_A_0To7aDDQ0_0),.clk(gclk));
	jdff dff_A_PNOJfyzw4_0(.dout(w_dff_A_fP7OT9lk4_0),.din(w_dff_A_PNOJfyzw4_0),.clk(gclk));
	jdff dff_A_fP7OT9lk4_0(.dout(w_dff_A_v2uaTy926_0),.din(w_dff_A_fP7OT9lk4_0),.clk(gclk));
	jdff dff_A_v2uaTy926_0(.dout(w_dff_A_wfeZErTh7_0),.din(w_dff_A_v2uaTy926_0),.clk(gclk));
	jdff dff_A_wfeZErTh7_0(.dout(w_dff_A_7m7ZrYDo0_0),.din(w_dff_A_wfeZErTh7_0),.clk(gclk));
	jdff dff_A_7m7ZrYDo0_0(.dout(w_dff_A_IIEnOhAI5_0),.din(w_dff_A_7m7ZrYDo0_0),.clk(gclk));
	jdff dff_A_IIEnOhAI5_0(.dout(w_dff_A_BdpJywMH1_0),.din(w_dff_A_IIEnOhAI5_0),.clk(gclk));
	jdff dff_A_BdpJywMH1_0(.dout(w_dff_A_OeX0mVef4_0),.din(w_dff_A_BdpJywMH1_0),.clk(gclk));
	jdff dff_A_OeX0mVef4_0(.dout(w_dff_A_dCOIv1RO8_0),.din(w_dff_A_OeX0mVef4_0),.clk(gclk));
	jdff dff_A_dCOIv1RO8_0(.dout(w_dff_A_gilxwOXP8_0),.din(w_dff_A_dCOIv1RO8_0),.clk(gclk));
	jdff dff_A_gilxwOXP8_0(.dout(w_dff_A_9s0IZ3cU9_0),.din(w_dff_A_gilxwOXP8_0),.clk(gclk));
	jdff dff_A_9s0IZ3cU9_0(.dout(w_dff_A_nd2IUhhm0_0),.din(w_dff_A_9s0IZ3cU9_0),.clk(gclk));
	jdff dff_A_nd2IUhhm0_0(.dout(w_dff_A_B55TaYlr1_0),.din(w_dff_A_nd2IUhhm0_0),.clk(gclk));
	jdff dff_A_B55TaYlr1_0(.dout(w_dff_A_hwYXCZVQ2_0),.din(w_dff_A_B55TaYlr1_0),.clk(gclk));
	jdff dff_A_hwYXCZVQ2_0(.dout(w_dff_A_K83xiXkF9_0),.din(w_dff_A_hwYXCZVQ2_0),.clk(gclk));
	jdff dff_A_K83xiXkF9_0(.dout(w_dff_A_rL6AXHc15_0),.din(w_dff_A_K83xiXkF9_0),.clk(gclk));
	jdff dff_A_rL6AXHc15_0(.dout(w_dff_A_kD19nGPu9_0),.din(w_dff_A_rL6AXHc15_0),.clk(gclk));
	jdff dff_A_kD19nGPu9_0(.dout(w_dff_A_QAAJOoP98_0),.din(w_dff_A_kD19nGPu9_0),.clk(gclk));
	jdff dff_A_QAAJOoP98_0(.dout(G5971gat),.din(w_dff_A_QAAJOoP98_0),.clk(gclk));
	jdff dff_A_b9xSmEOi6_2(.dout(w_dff_A_Xgwsrhnl1_0),.din(w_dff_A_b9xSmEOi6_2),.clk(gclk));
	jdff dff_A_Xgwsrhnl1_0(.dout(w_dff_A_RzkSdMIb4_0),.din(w_dff_A_Xgwsrhnl1_0),.clk(gclk));
	jdff dff_A_RzkSdMIb4_0(.dout(w_dff_A_zaboybat2_0),.din(w_dff_A_RzkSdMIb4_0),.clk(gclk));
	jdff dff_A_zaboybat2_0(.dout(w_dff_A_ZlJw7U003_0),.din(w_dff_A_zaboybat2_0),.clk(gclk));
	jdff dff_A_ZlJw7U003_0(.dout(w_dff_A_ieo9pNzn8_0),.din(w_dff_A_ZlJw7U003_0),.clk(gclk));
	jdff dff_A_ieo9pNzn8_0(.dout(w_dff_A_vrhsss888_0),.din(w_dff_A_ieo9pNzn8_0),.clk(gclk));
	jdff dff_A_vrhsss888_0(.dout(w_dff_A_woTG74pO7_0),.din(w_dff_A_vrhsss888_0),.clk(gclk));
	jdff dff_A_woTG74pO7_0(.dout(w_dff_A_72D0u0by4_0),.din(w_dff_A_woTG74pO7_0),.clk(gclk));
	jdff dff_A_72D0u0by4_0(.dout(w_dff_A_PLOyHNKq5_0),.din(w_dff_A_72D0u0by4_0),.clk(gclk));
	jdff dff_A_PLOyHNKq5_0(.dout(w_dff_A_29S28ue60_0),.din(w_dff_A_PLOyHNKq5_0),.clk(gclk));
	jdff dff_A_29S28ue60_0(.dout(w_dff_A_keZsIW5T0_0),.din(w_dff_A_29S28ue60_0),.clk(gclk));
	jdff dff_A_keZsIW5T0_0(.dout(w_dff_A_Q8l7aJsV0_0),.din(w_dff_A_keZsIW5T0_0),.clk(gclk));
	jdff dff_A_Q8l7aJsV0_0(.dout(w_dff_A_OhTY83Rd8_0),.din(w_dff_A_Q8l7aJsV0_0),.clk(gclk));
	jdff dff_A_OhTY83Rd8_0(.dout(w_dff_A_kM3AliSJ6_0),.din(w_dff_A_OhTY83Rd8_0),.clk(gclk));
	jdff dff_A_kM3AliSJ6_0(.dout(w_dff_A_86whUlow5_0),.din(w_dff_A_kM3AliSJ6_0),.clk(gclk));
	jdff dff_A_86whUlow5_0(.dout(w_dff_A_8UlC83LO4_0),.din(w_dff_A_86whUlow5_0),.clk(gclk));
	jdff dff_A_8UlC83LO4_0(.dout(w_dff_A_iKGDNwfx3_0),.din(w_dff_A_8UlC83LO4_0),.clk(gclk));
	jdff dff_A_iKGDNwfx3_0(.dout(w_dff_A_hN7dwSJE8_0),.din(w_dff_A_iKGDNwfx3_0),.clk(gclk));
	jdff dff_A_hN7dwSJE8_0(.dout(w_dff_A_TnokJ5nQ7_0),.din(w_dff_A_hN7dwSJE8_0),.clk(gclk));
	jdff dff_A_TnokJ5nQ7_0(.dout(w_dff_A_m86Z4tSp8_0),.din(w_dff_A_TnokJ5nQ7_0),.clk(gclk));
	jdff dff_A_m86Z4tSp8_0(.dout(w_dff_A_02Bq87UL8_0),.din(w_dff_A_m86Z4tSp8_0),.clk(gclk));
	jdff dff_A_02Bq87UL8_0(.dout(w_dff_A_WUnYuut38_0),.din(w_dff_A_02Bq87UL8_0),.clk(gclk));
	jdff dff_A_WUnYuut38_0(.dout(w_dff_A_cBWohS1Z9_0),.din(w_dff_A_WUnYuut38_0),.clk(gclk));
	jdff dff_A_cBWohS1Z9_0(.dout(w_dff_A_5sxAXsZZ2_0),.din(w_dff_A_cBWohS1Z9_0),.clk(gclk));
	jdff dff_A_5sxAXsZZ2_0(.dout(w_dff_A_NqQJ7Q9N7_0),.din(w_dff_A_5sxAXsZZ2_0),.clk(gclk));
	jdff dff_A_NqQJ7Q9N7_0(.dout(w_dff_A_edrMVVhI0_0),.din(w_dff_A_NqQJ7Q9N7_0),.clk(gclk));
	jdff dff_A_edrMVVhI0_0(.dout(w_dff_A_mc2ocRHi5_0),.din(w_dff_A_edrMVVhI0_0),.clk(gclk));
	jdff dff_A_mc2ocRHi5_0(.dout(w_dff_A_ClIG4uEj0_0),.din(w_dff_A_mc2ocRHi5_0),.clk(gclk));
	jdff dff_A_ClIG4uEj0_0(.dout(w_dff_A_qTqooJ4g5_0),.din(w_dff_A_ClIG4uEj0_0),.clk(gclk));
	jdff dff_A_qTqooJ4g5_0(.dout(G6123gat),.din(w_dff_A_qTqooJ4g5_0),.clk(gclk));
	jdff dff_A_okMi2w5I6_2(.dout(w_dff_A_mmqCAwQQ0_0),.din(w_dff_A_okMi2w5I6_2),.clk(gclk));
	jdff dff_A_mmqCAwQQ0_0(.dout(w_dff_A_jqnpxvNa9_0),.din(w_dff_A_mmqCAwQQ0_0),.clk(gclk));
	jdff dff_A_jqnpxvNa9_0(.dout(w_dff_A_D4aIypSf1_0),.din(w_dff_A_jqnpxvNa9_0),.clk(gclk));
	jdff dff_A_D4aIypSf1_0(.dout(w_dff_A_9F7A4NHn8_0),.din(w_dff_A_D4aIypSf1_0),.clk(gclk));
	jdff dff_A_9F7A4NHn8_0(.dout(w_dff_A_vSOF2bZ24_0),.din(w_dff_A_9F7A4NHn8_0),.clk(gclk));
	jdff dff_A_vSOF2bZ24_0(.dout(w_dff_A_uNXe2iYU3_0),.din(w_dff_A_vSOF2bZ24_0),.clk(gclk));
	jdff dff_A_uNXe2iYU3_0(.dout(w_dff_A_lRk8e8la5_0),.din(w_dff_A_uNXe2iYU3_0),.clk(gclk));
	jdff dff_A_lRk8e8la5_0(.dout(w_dff_A_cHwFbjZE0_0),.din(w_dff_A_lRk8e8la5_0),.clk(gclk));
	jdff dff_A_cHwFbjZE0_0(.dout(w_dff_A_lgumkYTG3_0),.din(w_dff_A_cHwFbjZE0_0),.clk(gclk));
	jdff dff_A_lgumkYTG3_0(.dout(w_dff_A_eb5JBGlA6_0),.din(w_dff_A_lgumkYTG3_0),.clk(gclk));
	jdff dff_A_eb5JBGlA6_0(.dout(w_dff_A_oic7v7yG5_0),.din(w_dff_A_eb5JBGlA6_0),.clk(gclk));
	jdff dff_A_oic7v7yG5_0(.dout(w_dff_A_FORKC9420_0),.din(w_dff_A_oic7v7yG5_0),.clk(gclk));
	jdff dff_A_FORKC9420_0(.dout(w_dff_A_gfUeqGK95_0),.din(w_dff_A_FORKC9420_0),.clk(gclk));
	jdff dff_A_gfUeqGK95_0(.dout(w_dff_A_Q7M2dmfq1_0),.din(w_dff_A_gfUeqGK95_0),.clk(gclk));
	jdff dff_A_Q7M2dmfq1_0(.dout(w_dff_A_hGO9D4ZK3_0),.din(w_dff_A_Q7M2dmfq1_0),.clk(gclk));
	jdff dff_A_hGO9D4ZK3_0(.dout(w_dff_A_eMN0Lyhf3_0),.din(w_dff_A_hGO9D4ZK3_0),.clk(gclk));
	jdff dff_A_eMN0Lyhf3_0(.dout(w_dff_A_IcRl3GVm5_0),.din(w_dff_A_eMN0Lyhf3_0),.clk(gclk));
	jdff dff_A_IcRl3GVm5_0(.dout(w_dff_A_d4vweEuQ4_0),.din(w_dff_A_IcRl3GVm5_0),.clk(gclk));
	jdff dff_A_d4vweEuQ4_0(.dout(w_dff_A_fhHm3dOI4_0),.din(w_dff_A_d4vweEuQ4_0),.clk(gclk));
	jdff dff_A_fhHm3dOI4_0(.dout(w_dff_A_TjnycSFa1_0),.din(w_dff_A_fhHm3dOI4_0),.clk(gclk));
	jdff dff_A_TjnycSFa1_0(.dout(w_dff_A_XenvYTYa7_0),.din(w_dff_A_TjnycSFa1_0),.clk(gclk));
	jdff dff_A_XenvYTYa7_0(.dout(w_dff_A_3hJ0cqb57_0),.din(w_dff_A_XenvYTYa7_0),.clk(gclk));
	jdff dff_A_3hJ0cqb57_0(.dout(w_dff_A_qvypK3uu5_0),.din(w_dff_A_3hJ0cqb57_0),.clk(gclk));
	jdff dff_A_qvypK3uu5_0(.dout(w_dff_A_TjEhGHcb0_0),.din(w_dff_A_qvypK3uu5_0),.clk(gclk));
	jdff dff_A_TjEhGHcb0_0(.dout(w_dff_A_uQZ1sL6C8_0),.din(w_dff_A_TjEhGHcb0_0),.clk(gclk));
	jdff dff_A_uQZ1sL6C8_0(.dout(w_dff_A_ShKNXAb48_0),.din(w_dff_A_uQZ1sL6C8_0),.clk(gclk));
	jdff dff_A_ShKNXAb48_0(.dout(w_dff_A_hT8zARTA3_0),.din(w_dff_A_ShKNXAb48_0),.clk(gclk));
	jdff dff_A_hT8zARTA3_0(.dout(G6150gat),.din(w_dff_A_hT8zARTA3_0),.clk(gclk));
	jdff dff_A_3iIVPtIy0_2(.dout(w_dff_A_TH0McGuv2_0),.din(w_dff_A_3iIVPtIy0_2),.clk(gclk));
	jdff dff_A_TH0McGuv2_0(.dout(w_dff_A_1tBOBIB03_0),.din(w_dff_A_TH0McGuv2_0),.clk(gclk));
	jdff dff_A_1tBOBIB03_0(.dout(w_dff_A_Qeapd9vl1_0),.din(w_dff_A_1tBOBIB03_0),.clk(gclk));
	jdff dff_A_Qeapd9vl1_0(.dout(w_dff_A_xWsUKLVc5_0),.din(w_dff_A_Qeapd9vl1_0),.clk(gclk));
	jdff dff_A_xWsUKLVc5_0(.dout(w_dff_A_EO82gKr26_0),.din(w_dff_A_xWsUKLVc5_0),.clk(gclk));
	jdff dff_A_EO82gKr26_0(.dout(w_dff_A_cGcdneVv0_0),.din(w_dff_A_EO82gKr26_0),.clk(gclk));
	jdff dff_A_cGcdneVv0_0(.dout(w_dff_A_OXZH8Ev40_0),.din(w_dff_A_cGcdneVv0_0),.clk(gclk));
	jdff dff_A_OXZH8Ev40_0(.dout(w_dff_A_ScY5LJbO9_0),.din(w_dff_A_OXZH8Ev40_0),.clk(gclk));
	jdff dff_A_ScY5LJbO9_0(.dout(w_dff_A_t9AJSCtL8_0),.din(w_dff_A_ScY5LJbO9_0),.clk(gclk));
	jdff dff_A_t9AJSCtL8_0(.dout(w_dff_A_8RJtbIcx6_0),.din(w_dff_A_t9AJSCtL8_0),.clk(gclk));
	jdff dff_A_8RJtbIcx6_0(.dout(w_dff_A_wkmvjhQv7_0),.din(w_dff_A_8RJtbIcx6_0),.clk(gclk));
	jdff dff_A_wkmvjhQv7_0(.dout(w_dff_A_MFUeYaer4_0),.din(w_dff_A_wkmvjhQv7_0),.clk(gclk));
	jdff dff_A_MFUeYaer4_0(.dout(w_dff_A_2r97kzzL1_0),.din(w_dff_A_MFUeYaer4_0),.clk(gclk));
	jdff dff_A_2r97kzzL1_0(.dout(w_dff_A_SZPHObf33_0),.din(w_dff_A_2r97kzzL1_0),.clk(gclk));
	jdff dff_A_SZPHObf33_0(.dout(w_dff_A_m7XT8p5y2_0),.din(w_dff_A_SZPHObf33_0),.clk(gclk));
	jdff dff_A_m7XT8p5y2_0(.dout(w_dff_A_Cqeo3oVs2_0),.din(w_dff_A_m7XT8p5y2_0),.clk(gclk));
	jdff dff_A_Cqeo3oVs2_0(.dout(w_dff_A_yFybcONs6_0),.din(w_dff_A_Cqeo3oVs2_0),.clk(gclk));
	jdff dff_A_yFybcONs6_0(.dout(w_dff_A_Cpf0AO8S8_0),.din(w_dff_A_yFybcONs6_0),.clk(gclk));
	jdff dff_A_Cpf0AO8S8_0(.dout(w_dff_A_mIDikPEU3_0),.din(w_dff_A_Cpf0AO8S8_0),.clk(gclk));
	jdff dff_A_mIDikPEU3_0(.dout(w_dff_A_8CQWHjB58_0),.din(w_dff_A_mIDikPEU3_0),.clk(gclk));
	jdff dff_A_8CQWHjB58_0(.dout(w_dff_A_2kzLPTvc2_0),.din(w_dff_A_8CQWHjB58_0),.clk(gclk));
	jdff dff_A_2kzLPTvc2_0(.dout(w_dff_A_CnQxLwoq5_0),.din(w_dff_A_2kzLPTvc2_0),.clk(gclk));
	jdff dff_A_CnQxLwoq5_0(.dout(w_dff_A_NM6yUNZu4_0),.din(w_dff_A_CnQxLwoq5_0),.clk(gclk));
	jdff dff_A_NM6yUNZu4_0(.dout(w_dff_A_QvzwaO3j7_0),.din(w_dff_A_NM6yUNZu4_0),.clk(gclk));
	jdff dff_A_QvzwaO3j7_0(.dout(w_dff_A_nESaPY9Y1_0),.din(w_dff_A_QvzwaO3j7_0),.clk(gclk));
	jdff dff_A_nESaPY9Y1_0(.dout(G6160gat),.din(w_dff_A_nESaPY9Y1_0),.clk(gclk));
	jdff dff_A_UyaYymEo5_2(.dout(w_dff_A_CLR1cD3l5_0),.din(w_dff_A_UyaYymEo5_2),.clk(gclk));
	jdff dff_A_CLR1cD3l5_0(.dout(w_dff_A_qbNEzUsY4_0),.din(w_dff_A_CLR1cD3l5_0),.clk(gclk));
	jdff dff_A_qbNEzUsY4_0(.dout(w_dff_A_7RC0Upu28_0),.din(w_dff_A_qbNEzUsY4_0),.clk(gclk));
	jdff dff_A_7RC0Upu28_0(.dout(w_dff_A_LZyI69R21_0),.din(w_dff_A_7RC0Upu28_0),.clk(gclk));
	jdff dff_A_LZyI69R21_0(.dout(w_dff_A_NpWq06f96_0),.din(w_dff_A_LZyI69R21_0),.clk(gclk));
	jdff dff_A_NpWq06f96_0(.dout(w_dff_A_jGs2LuPI6_0),.din(w_dff_A_NpWq06f96_0),.clk(gclk));
	jdff dff_A_jGs2LuPI6_0(.dout(w_dff_A_xvfqY82a2_0),.din(w_dff_A_jGs2LuPI6_0),.clk(gclk));
	jdff dff_A_xvfqY82a2_0(.dout(w_dff_A_7wOeM5Yg7_0),.din(w_dff_A_xvfqY82a2_0),.clk(gclk));
	jdff dff_A_7wOeM5Yg7_0(.dout(w_dff_A_a4aepqnD1_0),.din(w_dff_A_7wOeM5Yg7_0),.clk(gclk));
	jdff dff_A_a4aepqnD1_0(.dout(w_dff_A_N30RBU3j1_0),.din(w_dff_A_a4aepqnD1_0),.clk(gclk));
	jdff dff_A_N30RBU3j1_0(.dout(w_dff_A_H0X0Wm9v6_0),.din(w_dff_A_N30RBU3j1_0),.clk(gclk));
	jdff dff_A_H0X0Wm9v6_0(.dout(w_dff_A_c5N44hHk3_0),.din(w_dff_A_H0X0Wm9v6_0),.clk(gclk));
	jdff dff_A_c5N44hHk3_0(.dout(w_dff_A_JkVAFg4G2_0),.din(w_dff_A_c5N44hHk3_0),.clk(gclk));
	jdff dff_A_JkVAFg4G2_0(.dout(w_dff_A_T5wClN0H7_0),.din(w_dff_A_JkVAFg4G2_0),.clk(gclk));
	jdff dff_A_T5wClN0H7_0(.dout(w_dff_A_SE7CBLWH4_0),.din(w_dff_A_T5wClN0H7_0),.clk(gclk));
	jdff dff_A_SE7CBLWH4_0(.dout(w_dff_A_gS5j8tEI6_0),.din(w_dff_A_SE7CBLWH4_0),.clk(gclk));
	jdff dff_A_gS5j8tEI6_0(.dout(w_dff_A_oUED2Fr67_0),.din(w_dff_A_gS5j8tEI6_0),.clk(gclk));
	jdff dff_A_oUED2Fr67_0(.dout(w_dff_A_sQEAefrg6_0),.din(w_dff_A_oUED2Fr67_0),.clk(gclk));
	jdff dff_A_sQEAefrg6_0(.dout(w_dff_A_j1s66bpE5_0),.din(w_dff_A_sQEAefrg6_0),.clk(gclk));
	jdff dff_A_j1s66bpE5_0(.dout(w_dff_A_qXI94FpI0_0),.din(w_dff_A_j1s66bpE5_0),.clk(gclk));
	jdff dff_A_qXI94FpI0_0(.dout(w_dff_A_K7faFUhy4_0),.din(w_dff_A_qXI94FpI0_0),.clk(gclk));
	jdff dff_A_K7faFUhy4_0(.dout(w_dff_A_72L7YKCR9_0),.din(w_dff_A_K7faFUhy4_0),.clk(gclk));
	jdff dff_A_72L7YKCR9_0(.dout(w_dff_A_3MmwWSic9_0),.din(w_dff_A_72L7YKCR9_0),.clk(gclk));
	jdff dff_A_3MmwWSic9_0(.dout(w_dff_A_nCWPNuLc1_0),.din(w_dff_A_3MmwWSic9_0),.clk(gclk));
	jdff dff_A_nCWPNuLc1_0(.dout(G6170gat),.din(w_dff_A_nCWPNuLc1_0),.clk(gclk));
	jdff dff_A_5lkC1ky40_2(.dout(w_dff_A_OISVg6qP5_0),.din(w_dff_A_5lkC1ky40_2),.clk(gclk));
	jdff dff_A_OISVg6qP5_0(.dout(w_dff_A_y9lT7fhQ5_0),.din(w_dff_A_OISVg6qP5_0),.clk(gclk));
	jdff dff_A_y9lT7fhQ5_0(.dout(w_dff_A_2oxaerVo3_0),.din(w_dff_A_y9lT7fhQ5_0),.clk(gclk));
	jdff dff_A_2oxaerVo3_0(.dout(w_dff_A_dk5s9Qxe5_0),.din(w_dff_A_2oxaerVo3_0),.clk(gclk));
	jdff dff_A_dk5s9Qxe5_0(.dout(w_dff_A_LEc3BTSR4_0),.din(w_dff_A_dk5s9Qxe5_0),.clk(gclk));
	jdff dff_A_LEc3BTSR4_0(.dout(w_dff_A_1Jc7roqJ1_0),.din(w_dff_A_LEc3BTSR4_0),.clk(gclk));
	jdff dff_A_1Jc7roqJ1_0(.dout(w_dff_A_3sKt7CUo6_0),.din(w_dff_A_1Jc7roqJ1_0),.clk(gclk));
	jdff dff_A_3sKt7CUo6_0(.dout(w_dff_A_olkl87Jj3_0),.din(w_dff_A_3sKt7CUo6_0),.clk(gclk));
	jdff dff_A_olkl87Jj3_0(.dout(w_dff_A_wsZ5ojC10_0),.din(w_dff_A_olkl87Jj3_0),.clk(gclk));
	jdff dff_A_wsZ5ojC10_0(.dout(w_dff_A_Sb09y2jW7_0),.din(w_dff_A_wsZ5ojC10_0),.clk(gclk));
	jdff dff_A_Sb09y2jW7_0(.dout(w_dff_A_QtSPrnah2_0),.din(w_dff_A_Sb09y2jW7_0),.clk(gclk));
	jdff dff_A_QtSPrnah2_0(.dout(w_dff_A_dV7twkBH2_0),.din(w_dff_A_QtSPrnah2_0),.clk(gclk));
	jdff dff_A_dV7twkBH2_0(.dout(w_dff_A_A4pMx8fq4_0),.din(w_dff_A_dV7twkBH2_0),.clk(gclk));
	jdff dff_A_A4pMx8fq4_0(.dout(w_dff_A_hSmILgKU8_0),.din(w_dff_A_A4pMx8fq4_0),.clk(gclk));
	jdff dff_A_hSmILgKU8_0(.dout(w_dff_A_HIv5fYST7_0),.din(w_dff_A_hSmILgKU8_0),.clk(gclk));
	jdff dff_A_HIv5fYST7_0(.dout(w_dff_A_zWlbSlYz7_0),.din(w_dff_A_HIv5fYST7_0),.clk(gclk));
	jdff dff_A_zWlbSlYz7_0(.dout(w_dff_A_lInS9lwp3_0),.din(w_dff_A_zWlbSlYz7_0),.clk(gclk));
	jdff dff_A_lInS9lwp3_0(.dout(w_dff_A_PKjcF8ZR7_0),.din(w_dff_A_lInS9lwp3_0),.clk(gclk));
	jdff dff_A_PKjcF8ZR7_0(.dout(w_dff_A_sezIkoQa5_0),.din(w_dff_A_PKjcF8ZR7_0),.clk(gclk));
	jdff dff_A_sezIkoQa5_0(.dout(w_dff_A_5hturpCd7_0),.din(w_dff_A_sezIkoQa5_0),.clk(gclk));
	jdff dff_A_5hturpCd7_0(.dout(w_dff_A_HeJUNTxn5_0),.din(w_dff_A_5hturpCd7_0),.clk(gclk));
	jdff dff_A_HeJUNTxn5_0(.dout(w_dff_A_ZzX8KFrT7_0),.din(w_dff_A_HeJUNTxn5_0),.clk(gclk));
	jdff dff_A_ZzX8KFrT7_0(.dout(G6180gat),.din(w_dff_A_ZzX8KFrT7_0),.clk(gclk));
	jdff dff_A_yzVOykgA5_2(.dout(w_dff_A_nYyHfqI36_0),.din(w_dff_A_yzVOykgA5_2),.clk(gclk));
	jdff dff_A_nYyHfqI36_0(.dout(w_dff_A_t3iTvneP3_0),.din(w_dff_A_nYyHfqI36_0),.clk(gclk));
	jdff dff_A_t3iTvneP3_0(.dout(w_dff_A_I70Es19W1_0),.din(w_dff_A_t3iTvneP3_0),.clk(gclk));
	jdff dff_A_I70Es19W1_0(.dout(w_dff_A_V1TQ6Yxg8_0),.din(w_dff_A_I70Es19W1_0),.clk(gclk));
	jdff dff_A_V1TQ6Yxg8_0(.dout(w_dff_A_KJIJFdNi3_0),.din(w_dff_A_V1TQ6Yxg8_0),.clk(gclk));
	jdff dff_A_KJIJFdNi3_0(.dout(w_dff_A_ou10IiEt3_0),.din(w_dff_A_KJIJFdNi3_0),.clk(gclk));
	jdff dff_A_ou10IiEt3_0(.dout(w_dff_A_EuHGMMbj1_0),.din(w_dff_A_ou10IiEt3_0),.clk(gclk));
	jdff dff_A_EuHGMMbj1_0(.dout(w_dff_A_dv9MIYmE0_0),.din(w_dff_A_EuHGMMbj1_0),.clk(gclk));
	jdff dff_A_dv9MIYmE0_0(.dout(w_dff_A_wU7Ypb4D1_0),.din(w_dff_A_dv9MIYmE0_0),.clk(gclk));
	jdff dff_A_wU7Ypb4D1_0(.dout(w_dff_A_y3QdUFRR8_0),.din(w_dff_A_wU7Ypb4D1_0),.clk(gclk));
	jdff dff_A_y3QdUFRR8_0(.dout(w_dff_A_uXi4uYz30_0),.din(w_dff_A_y3QdUFRR8_0),.clk(gclk));
	jdff dff_A_uXi4uYz30_0(.dout(w_dff_A_nmauDiGY8_0),.din(w_dff_A_uXi4uYz30_0),.clk(gclk));
	jdff dff_A_nmauDiGY8_0(.dout(w_dff_A_nvlstr0F3_0),.din(w_dff_A_nmauDiGY8_0),.clk(gclk));
	jdff dff_A_nvlstr0F3_0(.dout(w_dff_A_uK05PgXN7_0),.din(w_dff_A_nvlstr0F3_0),.clk(gclk));
	jdff dff_A_uK05PgXN7_0(.dout(w_dff_A_2gUMQ6Ez8_0),.din(w_dff_A_uK05PgXN7_0),.clk(gclk));
	jdff dff_A_2gUMQ6Ez8_0(.dout(w_dff_A_hz74bhKB2_0),.din(w_dff_A_2gUMQ6Ez8_0),.clk(gclk));
	jdff dff_A_hz74bhKB2_0(.dout(w_dff_A_Fkys4IKG2_0),.din(w_dff_A_hz74bhKB2_0),.clk(gclk));
	jdff dff_A_Fkys4IKG2_0(.dout(w_dff_A_oVAjaGor1_0),.din(w_dff_A_Fkys4IKG2_0),.clk(gclk));
	jdff dff_A_oVAjaGor1_0(.dout(w_dff_A_mMZtzphy0_0),.din(w_dff_A_oVAjaGor1_0),.clk(gclk));
	jdff dff_A_mMZtzphy0_0(.dout(w_dff_A_upFUzfVE3_0),.din(w_dff_A_mMZtzphy0_0),.clk(gclk));
	jdff dff_A_upFUzfVE3_0(.dout(G6190gat),.din(w_dff_A_upFUzfVE3_0),.clk(gclk));
	jdff dff_A_CdP4FEpr4_2(.dout(w_dff_A_YmJQOPXe6_0),.din(w_dff_A_CdP4FEpr4_2),.clk(gclk));
	jdff dff_A_YmJQOPXe6_0(.dout(w_dff_A_dZ5hM3BL9_0),.din(w_dff_A_YmJQOPXe6_0),.clk(gclk));
	jdff dff_A_dZ5hM3BL9_0(.dout(w_dff_A_zMy2P6rC1_0),.din(w_dff_A_dZ5hM3BL9_0),.clk(gclk));
	jdff dff_A_zMy2P6rC1_0(.dout(w_dff_A_GThilhKC2_0),.din(w_dff_A_zMy2P6rC1_0),.clk(gclk));
	jdff dff_A_GThilhKC2_0(.dout(w_dff_A_ZlkLXRqS6_0),.din(w_dff_A_GThilhKC2_0),.clk(gclk));
	jdff dff_A_ZlkLXRqS6_0(.dout(w_dff_A_0gGD8cSC0_0),.din(w_dff_A_ZlkLXRqS6_0),.clk(gclk));
	jdff dff_A_0gGD8cSC0_0(.dout(w_dff_A_z6O5gkmr2_0),.din(w_dff_A_0gGD8cSC0_0),.clk(gclk));
	jdff dff_A_z6O5gkmr2_0(.dout(w_dff_A_KDyyAq3I6_0),.din(w_dff_A_z6O5gkmr2_0),.clk(gclk));
	jdff dff_A_KDyyAq3I6_0(.dout(w_dff_A_ENYoDgN90_0),.din(w_dff_A_KDyyAq3I6_0),.clk(gclk));
	jdff dff_A_ENYoDgN90_0(.dout(w_dff_A_giftbn219_0),.din(w_dff_A_ENYoDgN90_0),.clk(gclk));
	jdff dff_A_giftbn219_0(.dout(w_dff_A_pA2bGjJH7_0),.din(w_dff_A_giftbn219_0),.clk(gclk));
	jdff dff_A_pA2bGjJH7_0(.dout(w_dff_A_hwvQOeus6_0),.din(w_dff_A_pA2bGjJH7_0),.clk(gclk));
	jdff dff_A_hwvQOeus6_0(.dout(w_dff_A_snNeLaxx7_0),.din(w_dff_A_hwvQOeus6_0),.clk(gclk));
	jdff dff_A_snNeLaxx7_0(.dout(w_dff_A_XRf37nWQ7_0),.din(w_dff_A_snNeLaxx7_0),.clk(gclk));
	jdff dff_A_XRf37nWQ7_0(.dout(w_dff_A_oOspxazI5_0),.din(w_dff_A_XRf37nWQ7_0),.clk(gclk));
	jdff dff_A_oOspxazI5_0(.dout(w_dff_A_105n3lWY2_0),.din(w_dff_A_oOspxazI5_0),.clk(gclk));
	jdff dff_A_105n3lWY2_0(.dout(w_dff_A_l2BaYcZ29_0),.din(w_dff_A_105n3lWY2_0),.clk(gclk));
	jdff dff_A_l2BaYcZ29_0(.dout(w_dff_A_euOPKNzS4_0),.din(w_dff_A_l2BaYcZ29_0),.clk(gclk));
	jdff dff_A_euOPKNzS4_0(.dout(G6200gat),.din(w_dff_A_euOPKNzS4_0),.clk(gclk));
	jdff dff_A_HN7yDTv85_2(.dout(w_dff_A_RpX5OA6x2_0),.din(w_dff_A_HN7yDTv85_2),.clk(gclk));
	jdff dff_A_RpX5OA6x2_0(.dout(w_dff_A_jmf8UfBV6_0),.din(w_dff_A_RpX5OA6x2_0),.clk(gclk));
	jdff dff_A_jmf8UfBV6_0(.dout(w_dff_A_6ivIQwPA9_0),.din(w_dff_A_jmf8UfBV6_0),.clk(gclk));
	jdff dff_A_6ivIQwPA9_0(.dout(w_dff_A_JNkMfS620_0),.din(w_dff_A_6ivIQwPA9_0),.clk(gclk));
	jdff dff_A_JNkMfS620_0(.dout(w_dff_A_hkNq3aHH0_0),.din(w_dff_A_JNkMfS620_0),.clk(gclk));
	jdff dff_A_hkNq3aHH0_0(.dout(w_dff_A_kM1wyV0K5_0),.din(w_dff_A_hkNq3aHH0_0),.clk(gclk));
	jdff dff_A_kM1wyV0K5_0(.dout(w_dff_A_RyDYXRC51_0),.din(w_dff_A_kM1wyV0K5_0),.clk(gclk));
	jdff dff_A_RyDYXRC51_0(.dout(w_dff_A_3GSiUFl94_0),.din(w_dff_A_RyDYXRC51_0),.clk(gclk));
	jdff dff_A_3GSiUFl94_0(.dout(w_dff_A_Qm70PGdU8_0),.din(w_dff_A_3GSiUFl94_0),.clk(gclk));
	jdff dff_A_Qm70PGdU8_0(.dout(w_dff_A_EAGjHtSv9_0),.din(w_dff_A_Qm70PGdU8_0),.clk(gclk));
	jdff dff_A_EAGjHtSv9_0(.dout(w_dff_A_kD5VZRvd3_0),.din(w_dff_A_EAGjHtSv9_0),.clk(gclk));
	jdff dff_A_kD5VZRvd3_0(.dout(w_dff_A_HaGpOdSV0_0),.din(w_dff_A_kD5VZRvd3_0),.clk(gclk));
	jdff dff_A_HaGpOdSV0_0(.dout(w_dff_A_MSuQjyhW9_0),.din(w_dff_A_HaGpOdSV0_0),.clk(gclk));
	jdff dff_A_MSuQjyhW9_0(.dout(w_dff_A_QYdJGrRl3_0),.din(w_dff_A_MSuQjyhW9_0),.clk(gclk));
	jdff dff_A_QYdJGrRl3_0(.dout(w_dff_A_WU8237Lx4_0),.din(w_dff_A_QYdJGrRl3_0),.clk(gclk));
	jdff dff_A_WU8237Lx4_0(.dout(w_dff_A_uQFiSjFw0_0),.din(w_dff_A_WU8237Lx4_0),.clk(gclk));
	jdff dff_A_uQFiSjFw0_0(.dout(G6210gat),.din(w_dff_A_uQFiSjFw0_0),.clk(gclk));
	jdff dff_A_5arqhEZw5_2(.dout(w_dff_A_9CKZi3AS6_0),.din(w_dff_A_5arqhEZw5_2),.clk(gclk));
	jdff dff_A_9CKZi3AS6_0(.dout(w_dff_A_8al8690v7_0),.din(w_dff_A_9CKZi3AS6_0),.clk(gclk));
	jdff dff_A_8al8690v7_0(.dout(w_dff_A_CL7wU4204_0),.din(w_dff_A_8al8690v7_0),.clk(gclk));
	jdff dff_A_CL7wU4204_0(.dout(w_dff_A_Bi1nK5XC8_0),.din(w_dff_A_CL7wU4204_0),.clk(gclk));
	jdff dff_A_Bi1nK5XC8_0(.dout(w_dff_A_9sFUi5mS4_0),.din(w_dff_A_Bi1nK5XC8_0),.clk(gclk));
	jdff dff_A_9sFUi5mS4_0(.dout(w_dff_A_cfkZlF4D1_0),.din(w_dff_A_9sFUi5mS4_0),.clk(gclk));
	jdff dff_A_cfkZlF4D1_0(.dout(w_dff_A_vM5byLDi9_0),.din(w_dff_A_cfkZlF4D1_0),.clk(gclk));
	jdff dff_A_vM5byLDi9_0(.dout(w_dff_A_f1KZGQfn5_0),.din(w_dff_A_vM5byLDi9_0),.clk(gclk));
	jdff dff_A_f1KZGQfn5_0(.dout(w_dff_A_MaLPbrWR8_0),.din(w_dff_A_f1KZGQfn5_0),.clk(gclk));
	jdff dff_A_MaLPbrWR8_0(.dout(w_dff_A_EbVELEbw0_0),.din(w_dff_A_MaLPbrWR8_0),.clk(gclk));
	jdff dff_A_EbVELEbw0_0(.dout(w_dff_A_5CXZnEeV2_0),.din(w_dff_A_EbVELEbw0_0),.clk(gclk));
	jdff dff_A_5CXZnEeV2_0(.dout(w_dff_A_ZJxOxn1Z9_0),.din(w_dff_A_5CXZnEeV2_0),.clk(gclk));
	jdff dff_A_ZJxOxn1Z9_0(.dout(w_dff_A_cW4hY6gH8_0),.din(w_dff_A_ZJxOxn1Z9_0),.clk(gclk));
	jdff dff_A_cW4hY6gH8_0(.dout(w_dff_A_VtS6o35P7_0),.din(w_dff_A_cW4hY6gH8_0),.clk(gclk));
	jdff dff_A_VtS6o35P7_0(.dout(G6220gat),.din(w_dff_A_VtS6o35P7_0),.clk(gclk));
	jdff dff_A_OWGNsutV7_2(.dout(w_dff_A_H03cf2lL9_0),.din(w_dff_A_OWGNsutV7_2),.clk(gclk));
	jdff dff_A_H03cf2lL9_0(.dout(w_dff_A_5lHIJwDH5_0),.din(w_dff_A_H03cf2lL9_0),.clk(gclk));
	jdff dff_A_5lHIJwDH5_0(.dout(w_dff_A_j2EuERaM6_0),.din(w_dff_A_5lHIJwDH5_0),.clk(gclk));
	jdff dff_A_j2EuERaM6_0(.dout(w_dff_A_CG92fvNm1_0),.din(w_dff_A_j2EuERaM6_0),.clk(gclk));
	jdff dff_A_CG92fvNm1_0(.dout(w_dff_A_P87da74r3_0),.din(w_dff_A_CG92fvNm1_0),.clk(gclk));
	jdff dff_A_P87da74r3_0(.dout(w_dff_A_XTmRmp8A1_0),.din(w_dff_A_P87da74r3_0),.clk(gclk));
	jdff dff_A_XTmRmp8A1_0(.dout(w_dff_A_GgkbaN2K3_0),.din(w_dff_A_XTmRmp8A1_0),.clk(gclk));
	jdff dff_A_GgkbaN2K3_0(.dout(w_dff_A_DKlpFjiM6_0),.din(w_dff_A_GgkbaN2K3_0),.clk(gclk));
	jdff dff_A_DKlpFjiM6_0(.dout(w_dff_A_Cv8Wk0hu7_0),.din(w_dff_A_DKlpFjiM6_0),.clk(gclk));
	jdff dff_A_Cv8Wk0hu7_0(.dout(w_dff_A_uD06ZPIu0_0),.din(w_dff_A_Cv8Wk0hu7_0),.clk(gclk));
	jdff dff_A_uD06ZPIu0_0(.dout(w_dff_A_PM8G6V623_0),.din(w_dff_A_uD06ZPIu0_0),.clk(gclk));
	jdff dff_A_PM8G6V623_0(.dout(w_dff_A_ldmD4Pg34_0),.din(w_dff_A_PM8G6V623_0),.clk(gclk));
	jdff dff_A_ldmD4Pg34_0(.dout(G6230gat),.din(w_dff_A_ldmD4Pg34_0),.clk(gclk));
	jdff dff_A_FgSjYYdM3_2(.dout(w_dff_A_tJmfc1aX8_0),.din(w_dff_A_FgSjYYdM3_2),.clk(gclk));
	jdff dff_A_tJmfc1aX8_0(.dout(w_dff_A_esA7WomA6_0),.din(w_dff_A_tJmfc1aX8_0),.clk(gclk));
	jdff dff_A_esA7WomA6_0(.dout(w_dff_A_bV8WZ6pc6_0),.din(w_dff_A_esA7WomA6_0),.clk(gclk));
	jdff dff_A_bV8WZ6pc6_0(.dout(w_dff_A_Tyex67UV2_0),.din(w_dff_A_bV8WZ6pc6_0),.clk(gclk));
	jdff dff_A_Tyex67UV2_0(.dout(w_dff_A_tBkbXq5g4_0),.din(w_dff_A_Tyex67UV2_0),.clk(gclk));
	jdff dff_A_tBkbXq5g4_0(.dout(w_dff_A_udNx3lHZ0_0),.din(w_dff_A_tBkbXq5g4_0),.clk(gclk));
	jdff dff_A_udNx3lHZ0_0(.dout(w_dff_A_4PmcjKeH8_0),.din(w_dff_A_udNx3lHZ0_0),.clk(gclk));
	jdff dff_A_4PmcjKeH8_0(.dout(w_dff_A_b1vuRf3a4_0),.din(w_dff_A_4PmcjKeH8_0),.clk(gclk));
	jdff dff_A_b1vuRf3a4_0(.dout(w_dff_A_dua3Bi0M8_0),.din(w_dff_A_b1vuRf3a4_0),.clk(gclk));
	jdff dff_A_dua3Bi0M8_0(.dout(w_dff_A_vcl3bDJl7_0),.din(w_dff_A_dua3Bi0M8_0),.clk(gclk));
	jdff dff_A_vcl3bDJl7_0(.dout(G6240gat),.din(w_dff_A_vcl3bDJl7_0),.clk(gclk));
	jdff dff_A_c6Fm6OCo3_2(.dout(w_dff_A_x8t5Shk49_0),.din(w_dff_A_c6Fm6OCo3_2),.clk(gclk));
	jdff dff_A_x8t5Shk49_0(.dout(w_dff_A_wDfxn7zY6_0),.din(w_dff_A_x8t5Shk49_0),.clk(gclk));
	jdff dff_A_wDfxn7zY6_0(.dout(w_dff_A_AjLI4VpR0_0),.din(w_dff_A_wDfxn7zY6_0),.clk(gclk));
	jdff dff_A_AjLI4VpR0_0(.dout(w_dff_A_r3sMAMPb3_0),.din(w_dff_A_AjLI4VpR0_0),.clk(gclk));
	jdff dff_A_r3sMAMPb3_0(.dout(w_dff_A_WR9E9Aag2_0),.din(w_dff_A_r3sMAMPb3_0),.clk(gclk));
	jdff dff_A_WR9E9Aag2_0(.dout(w_dff_A_kuq4Pi7Z7_0),.din(w_dff_A_WR9E9Aag2_0),.clk(gclk));
	jdff dff_A_kuq4Pi7Z7_0(.dout(w_dff_A_ytZxEyU76_0),.din(w_dff_A_kuq4Pi7Z7_0),.clk(gclk));
	jdff dff_A_ytZxEyU76_0(.dout(w_dff_A_JW9f4wSa2_0),.din(w_dff_A_ytZxEyU76_0),.clk(gclk));
	jdff dff_A_JW9f4wSa2_0(.dout(G6250gat),.din(w_dff_A_JW9f4wSa2_0),.clk(gclk));
	jdff dff_A_cTXjgFSt7_2(.dout(w_dff_A_zgz3aUWA5_0),.din(w_dff_A_cTXjgFSt7_2),.clk(gclk));
	jdff dff_A_zgz3aUWA5_0(.dout(w_dff_A_AvJiQkvT6_0),.din(w_dff_A_zgz3aUWA5_0),.clk(gclk));
	jdff dff_A_AvJiQkvT6_0(.dout(w_dff_A_apui6QwY8_0),.din(w_dff_A_AvJiQkvT6_0),.clk(gclk));
	jdff dff_A_apui6QwY8_0(.dout(w_dff_A_QWaLqLGT0_0),.din(w_dff_A_apui6QwY8_0),.clk(gclk));
	jdff dff_A_QWaLqLGT0_0(.dout(w_dff_A_7HV5KXse8_0),.din(w_dff_A_QWaLqLGT0_0),.clk(gclk));
	jdff dff_A_7HV5KXse8_0(.dout(w_dff_A_OnBH3vUl3_0),.din(w_dff_A_7HV5KXse8_0),.clk(gclk));
	jdff dff_A_OnBH3vUl3_0(.dout(G6260gat),.din(w_dff_A_OnBH3vUl3_0),.clk(gclk));
	jdff dff_A_MtaWg8ib7_2(.dout(w_dff_A_KzyXslny6_0),.din(w_dff_A_MtaWg8ib7_2),.clk(gclk));
	jdff dff_A_KzyXslny6_0(.dout(w_dff_A_wSRmAakt8_0),.din(w_dff_A_KzyXslny6_0),.clk(gclk));
	jdff dff_A_wSRmAakt8_0(.dout(w_dff_A_ZVdSCnXX0_0),.din(w_dff_A_wSRmAakt8_0),.clk(gclk));
	jdff dff_A_ZVdSCnXX0_0(.dout(w_dff_A_j9NUrqag8_0),.din(w_dff_A_ZVdSCnXX0_0),.clk(gclk));
	jdff dff_A_j9NUrqag8_0(.dout(G6270gat),.din(w_dff_A_j9NUrqag8_0),.clk(gclk));
	jdff dff_A_GvGhDXPx3_2(.dout(w_dff_A_PAyX2J2a8_0),.din(w_dff_A_GvGhDXPx3_2),.clk(gclk));
	jdff dff_A_PAyX2J2a8_0(.dout(w_dff_A_N2tTzVE14_0),.din(w_dff_A_PAyX2J2a8_0),.clk(gclk));
	jdff dff_A_N2tTzVE14_0(.dout(G6280gat),.din(w_dff_A_N2tTzVE14_0),.clk(gclk));
	jdff dff_A_l6uLDiYR0_2(.dout(G6288gat),.din(w_dff_A_l6uLDiYR0_2),.clk(gclk));
endmodule

