// Benchmark "top" written by ABC on Thu May 28 22:02:24 2020

module rf_sqrt (a, asqrt);
  input [127:0] a;
  output [63:0] asqrt;
  wire n192, n193, n194, n195, n196, n197, n199, n200, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n258, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n428, n429, n430,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n504, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n593, n594, n595, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n687, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n794, n795, n796, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n910, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1037, n1038, n1039, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1169, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1315, n1316,
    n1317, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1472, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1644, n1645, n1646, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1817, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2008,
    n2009, n2010, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2206, n2208, n2209, n2210, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2423, n2424,
    n2425, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2637,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2873, n2874, n2875, n2877, n2878, n2879, n2880, n2881,
    n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
    n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
    n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
    n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
    n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
    n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3112, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
    n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
    n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3374, n3375, n3376,
    n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
    n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
    n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
    n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
    n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
    n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
    n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
    n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3629,
    n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
    n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
    n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
    n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
    n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3910, n3911, n3912,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
    n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
    n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
    n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
    n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
    n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4190, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
    n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4497, n4498,
    n4499, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
    n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4793, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
    n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
    n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
    n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
    n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
    n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
    n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
    n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
    n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
    n5113, n5114, n5115, n5116, n5119, n5120, n5121, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
    n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
    n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
    n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5440, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
    n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
    n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
    n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
    n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
    n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
    n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
    n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
    n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
    n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
    n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
    n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
    n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
    n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
    n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
    n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
    n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
    n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
    n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
    n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
    n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
    n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
    n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
    n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
    n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
    n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
    n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6128, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
    n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
    n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
    n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
    n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
    n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
    n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
    n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
    n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
    n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
    n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
    n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
    n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
    n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
    n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
    n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
    n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
    n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
    n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
    n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
    n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
    n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
    n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
    n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
    n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
    n6858, n6859, n6860, n6861, n6862, n6865, n6867, n6868, n6869, n6870,
    n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
    n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
    n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
    n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
    n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
    n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
    n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
    n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
    n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
    n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
    n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
    n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
    n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
    n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
    n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
    n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
    n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
    n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
    n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
    n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
    n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
    n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
    n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
    n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
    n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
    n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
    n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
    n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7640, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
    n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
    n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
    n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
    n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
    n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
    n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
    n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
    n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
    n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
    n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
    n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
    n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
    n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
    n8450, n8451, n8454, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
    n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
    n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
    n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
    n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
    n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
    n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
    n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
    n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
    n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
    n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9311, n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
    n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
    n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
    n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
    n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
    n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
    n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
    n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
    n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
    n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
    n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
    n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
    n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
    n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
    n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
    n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
    n9769, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
    n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
    n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
    n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
    n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
    n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
    n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
    n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
    n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
    n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
    n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
    n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
    n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
    n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
    n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
    n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
    n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
    n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
    n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
    n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
    n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
    n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
    n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
    n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
    n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
    n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
    n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
    n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
    n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10212, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
    n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
    n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
    n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
    n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
    n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
    n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
    n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
    n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
    n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
    n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
    n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
    n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
    n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
    n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
    n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
    n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
    n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
    n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
    n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
    n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
    n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
    n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
    n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
    n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
    n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
    n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
    n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
    n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11154, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
    n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
    n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
    n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
    n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
    n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
    n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
    n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
    n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
    n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
    n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
    n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
    n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
    n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
    n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
    n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
    n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
    n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
    n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
    n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
    n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
    n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
    n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
    n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
    n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
    n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
    n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
    n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719, n11721, n11722, n11723,
    n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
    n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
    n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
    n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
    n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
    n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
    n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
    n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
    n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12141, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12673,
    n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
    n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
    n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
    n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733, n12735, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
    n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
    n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
    n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
    n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
    n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
    n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
    n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
    n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
    n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
    n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
    n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
    n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
    n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
    n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
    n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
    n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
    n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
    n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
    n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13170, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
    n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
    n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
    n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
    n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
    n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
    n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
    n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
    n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
    n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
    n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
    n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
    n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
    n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
    n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
    n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
    n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
    n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
    n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
    n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
    n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
    n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
    n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
    n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13782, n13783, n13784, n13785, n13786, n13787,
    n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
    n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
    n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
    n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
    n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
    n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
    n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
    n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
    n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
    n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
    n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
    n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
    n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
    n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
    n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
    n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
    n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
    n14238, n14239, n14242, n14244, n14245, n14246, n14247, n14248, n14249,
    n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
    n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
    n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
    n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
    n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
    n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
    n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
    n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
    n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
    n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
    n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
    n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
    n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
    n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
    n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
    n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
    n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
    n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
    n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
    n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
    n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
    n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
    n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
    n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
    n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
    n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
    n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
    n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
    n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
    n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
    n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
    n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
    n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
    n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
    n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
    n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
    n14873, n14874, n14875, n14876, n14877, n14878, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
    n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
    n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
    n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
    n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
    n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
    n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
    n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
    n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
    n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
    n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
    n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
    n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
    n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
    n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
    n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
    n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
    n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
    n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
    n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
    n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
    n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
    n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
    n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
    n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
    n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
    n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15357, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
    n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
    n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
    n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
    n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
    n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
    n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
    n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
    n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
    n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
    n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
    n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
    n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
    n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
    n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
    n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
    n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
    n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
    n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
    n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
    n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
    n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
    n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
    n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
    n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
    n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
    n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
    n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
    n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
    n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
    n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
    n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
    n15948, n15949, n15950, n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
    n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
    n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
    n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
    n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
    n16013, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
    n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
    n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
    n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
    n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
    n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
    n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
    n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
    n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
    n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
    n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
    n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
    n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
    n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16516, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
    n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
    n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
    n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
    n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
    n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
    n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
    n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
    n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
    n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
    n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
    n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
    n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
    n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
    n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
    n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
    n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
    n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
    n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
    n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
    n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
    n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
    n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
    n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
    n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
    n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
    n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
    n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
    n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
    n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
    n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
    n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
    n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17138, n17139, n17140, n17141, n17142, n17143,
    n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
    n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
    n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
    n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
    n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
    n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
    n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
    n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
    n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
    n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
    n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
    n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
    n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
    n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
    n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
    n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
    n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
    n17712, n17713, n17716, n17718, n17719, n17720, n17721, n17722, n17723,
    n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
    n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
    n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
    n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
    n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
    n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
    n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
    n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
    n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
    n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
    n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
    n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
    n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
    n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
    n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
    n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
    n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
    n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
    n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
    n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
    n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
    n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
    n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
    n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
    n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
    n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
    n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
    n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
    n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
    n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
    n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
    n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
    n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
    n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
    n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
    n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
    n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
    n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
    n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
    n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
    n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
    n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
    n18372, n18373, n18374, n18375, n18376, n18377, n18379, n18380, n18381,
    n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
    n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
    n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
    n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
    n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
    n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
    n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
    n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
    n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
    n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
    n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
    n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
    n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
    n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
    n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
    n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
    n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
    n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
    n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
    n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
    n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
    n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
    n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
    n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
    n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
    n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
    n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
    n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
    n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
    n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
    n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
    n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
    n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
    n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
    n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
    n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
    n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
    n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
    n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
    n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
    n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
    n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
    n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
    n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
    n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
    n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
    n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
    n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
    n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
    n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
    n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
    n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
    n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
    n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
    n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
    n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
    n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
    n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
    n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
    n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
    n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
    n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
    n18949, n18950, n18951, n18952, n18953, n18954, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
    n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
    n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
    n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
    n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
    n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
    n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
    n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
    n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
    n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
    n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
    n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
    n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
    n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
    n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
    n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
    n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
    n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
    n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
    n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
    n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
    n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
    n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
    n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
    n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
    n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
    n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
    n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
    n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
    n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
    n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
    n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
    n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
    n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
    n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
    n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
    n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
    n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
    n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
    n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
    n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
    n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
    n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
    n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
    n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
    n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
    n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19639, n19640, n19641, n19642, n19643,
    n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
    n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
    n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
    n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
    n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
    n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
    n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
    n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
    n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
    n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
    n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
    n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
    n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
    n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
    n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
    n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
    n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
    n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
    n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
    n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
    n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
    n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
    n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
    n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
    n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
    n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
    n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
    n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
    n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
    n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
    n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
    n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
    n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
    n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
    n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
    n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
    n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
    n20229, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
    n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
    n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
    n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
    n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
    n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
    n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
    n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
    n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
    n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
    n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
    n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
    n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
    n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
    n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
    n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
    n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
    n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
    n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
    n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
    n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
    n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
    n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
    n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
    n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
    n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
    n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
    n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
    n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
    n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
    n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
    n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
    n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
    n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
    n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
    n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
    n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
    n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
    n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
    n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
    n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
    n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
    n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
    n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
    n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
    n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
    n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
    n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
    n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
    n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
    n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
    n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
    n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
    n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
    n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
    n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
    n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
    n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
    n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
    n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
    n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
    n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
    n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
    n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
    n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
    n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
    n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
    n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
    n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
    n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
    n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
    n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
    n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
    n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
    n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
    n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
    n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
    n20923, n20924, n20925, n20926, n20928, n20929, n20930, n20931, n20932,
    n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
    n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
    n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
    n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
    n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
    n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
    n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
    n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
    n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
    n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
    n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
    n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
    n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
    n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
    n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
    n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
    n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
    n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
    n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
    n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
    n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
    n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
    n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
    n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
    n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
    n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
    n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
    n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
    n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
    n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
    n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
    n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
    n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
    n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
    n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
    n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
    n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
    n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
    n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
    n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
    n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
    n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
    n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
    n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
    n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
    n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
    n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
    n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
    n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
    n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
    n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
    n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
    n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
    n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
    n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
    n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
    n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
    n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
    n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508;
  jnot g00000(.din(a[126] ), .dout(n192));
  jnot g00001(.din(a[127] ), .dout(n193));
  jand g00002(.dina(n193), .dinb(n192), .dout(n194));
  jand g00003(.dina(a[127] ), .dinb(a[126] ), .dout(n195));
  jor  g00004(.dina(a[125] ), .dinb(a[124] ), .dout(n196));
  jand g00005(.dina(n196), .dinb(n192), .dout(n197));
  jor  g00006(.dina(n197), .dinb(n195), .dout(asqrt[62] ));
  jnot g00007(.din(asqrt[62] ), .dout(n199));
  jnot g00008(.din(a[63] ), .dout(n200));
  jnot g00009(.din(n194), .dout(asqrt[63] ));
  jnot g00010(.din(a[125] ), .dout(n202));
  jnot g00011(.din(a[124] ), .dout(n203));
  jand g00012(.dina(asqrt[62] ), .dinb(n203), .dout(n204));
  jor  g00013(.dina(n204), .dinb(n202), .dout(n205));
  jnot g00014(.din(n196), .dout(n206));
  jand g00015(.dina(n206), .dinb(n195), .dout(n207));
  jnot g00016(.din(n207), .dout(n208));
  jand g00017(.dina(n208), .dinb(n205), .dout(n209));
  jand g00018(.dina(asqrt[62] ), .dinb(a[124] ), .dout(n210));
  jnot g00019(.din(a[122] ), .dout(n211));
  jnot g00020(.din(a[123] ), .dout(n212));
  jand g00021(.dina(n203), .dinb(n212), .dout(n213));
  jand g00022(.dina(n213), .dinb(n211), .dout(n214));
  jor  g00023(.dina(n214), .dinb(n210), .dout(n215));
  jand g00024(.dina(n215), .dinb(n209), .dout(n216));
  jor  g00025(.dina(n216), .dinb(asqrt[63] ), .dout(n217));
  jor  g00026(.dina(n215), .dinb(n209), .dout(n218));
  jand g00027(.dina(n206), .dinb(a[126] ), .dout(n219));
  jor  g00028(.dina(n197), .dinb(n193), .dout(n220));
  jor  g00029(.dina(n220), .dinb(n219), .dout(n221));
  jand g00030(.dina(n221), .dinb(n218), .dout(n222));
  jand g00031(.dina(n222), .dinb(n217), .dout(n223));
  jnot g00032(.din(n223), .dout(asqrt[61] ));
  jor  g00033(.dina(asqrt[61] ), .dinb(n199), .dout(n225));
  jor  g00034(.dina(n223), .dinb(a[122] ), .dout(n226));
  jor  g00035(.dina(n226), .dinb(a[123] ), .dout(n227));
  jand g00036(.dina(n227), .dinb(n225), .dout(n228));
  jxor g00037(.dina(n228), .dinb(n203), .dout(n229));
  jor  g00038(.dina(n223), .dinb(n211), .dout(n230));
  jnot g00039(.din(a[120] ), .dout(n231));
  jnot g00040(.din(a[121] ), .dout(n232));
  jand g00041(.dina(n211), .dinb(n232), .dout(n233));
  jand g00042(.dina(n233), .dinb(n231), .dout(n234));
  jnot g00043(.din(n234), .dout(n235));
  jand g00044(.dina(n235), .dinb(n230), .dout(n236));
  jor  g00045(.dina(n236), .dinb(n199), .dout(n237));
  jand g00046(.dina(n236), .dinb(n199), .dout(n238));
  jxor g00047(.dina(n226), .dinb(n212), .dout(n239));
  jor  g00048(.dina(n239), .dinb(n238), .dout(n240));
  jand g00049(.dina(n240), .dinb(n237), .dout(n241));
  jor  g00050(.dina(n241), .dinb(n229), .dout(n242));
  jnot g00051(.din(n218), .dout(n243));
  jnot g00052(.din(n221), .dout(n244));
  jand g00053(.dina(n244), .dinb(n216), .dout(n245));
  jor  g00054(.dina(n245), .dinb(n243), .dout(n246));
  jor  g00055(.dina(n246), .dinb(n242), .dout(n247));
  jand g00056(.dina(n247), .dinb(n194), .dout(n248));
  jand g00057(.dina(n241), .dinb(n229), .dout(n249));
  jand g00058(.dina(asqrt[61] ), .dinb(n209), .dout(n250));
  jor  g00059(.dina(n250), .dinb(n215), .dout(n251));
  jnot g00060(.din(n216), .dout(n252));
  jand g00061(.dina(n252), .dinb(asqrt[63] ), .dout(n253));
  jand g00062(.dina(n253), .dinb(n251), .dout(n254));
  jor  g00063(.dina(n254), .dinb(n249), .dout(n258));
  jor  g00064(.dina(n258), .dinb(n248), .dout(asqrt[60] ));
  jand g00065(.dina(asqrt[60] ), .dinb(a[120] ), .dout(n260));
  jnot g00066(.din(a[118] ), .dout(n261));
  jnot g00067(.din(a[119] ), .dout(n262));
  jand g00068(.dina(n231), .dinb(n262), .dout(n263));
  jand g00069(.dina(n263), .dinb(n261), .dout(n264));
  jor  g00070(.dina(n264), .dinb(n260), .dout(n265));
  jand g00071(.dina(n265), .dinb(asqrt[61] ), .dout(n266));
  jand g00072(.dina(asqrt[60] ), .dinb(n231), .dout(n267));
  jxor g00073(.dina(n267), .dinb(n232), .dout(n268));
  jor  g00074(.dina(n265), .dinb(asqrt[61] ), .dout(n269));
  jand g00075(.dina(n269), .dinb(n268), .dout(n270));
  jor  g00076(.dina(n270), .dinb(n266), .dout(n271));
  jand g00077(.dina(n271), .dinb(asqrt[62] ), .dout(n272));
  jor  g00078(.dina(n266), .dinb(asqrt[62] ), .dout(n273));
  jor  g00079(.dina(n273), .dinb(n270), .dout(n274));
  jand g00080(.dina(n267), .dinb(n232), .dout(n275));
  jnot g00081(.din(n248), .dout(n276));
  jnot g00082(.din(n249), .dout(n277));
  jnot g00083(.din(n254), .dout(n278));
  jand g00084(.dina(n278), .dinb(asqrt[61] ), .dout(n279));
  jand g00085(.dina(n279), .dinb(n277), .dout(n280));
  jand g00086(.dina(n280), .dinb(n276), .dout(n281));
  jor  g00087(.dina(n281), .dinb(n275), .dout(n282));
  jxor g00088(.dina(n282), .dinb(n211), .dout(n283));
  jand g00089(.dina(n283), .dinb(n274), .dout(n284));
  jor  g00090(.dina(n284), .dinb(n272), .dout(n285));
  jnot g00091(.din(n239), .dout(n286));
  jxor g00092(.dina(n236), .dinb(n199), .dout(n287));
  jand g00093(.dina(n287), .dinb(asqrt[60] ), .dout(n288));
  jxor g00094(.dina(n288), .dinb(n286), .dout(n289));
  jnot g00095(.din(asqrt[60] ), .dout(n290));
  jor  g00096(.dina(n290), .dinb(n242), .dout(n291));
  jand g00097(.dina(n291), .dinb(n277), .dout(n292));
  jand g00098(.dina(n292), .dinb(n289), .dout(n293));
  jand g00099(.dina(n293), .dinb(n285), .dout(n294));
  jor  g00100(.dina(n294), .dinb(asqrt[63] ), .dout(n295));
  jor  g00101(.dina(n289), .dinb(n285), .dout(n296));
  jnot g00102(.din(n229), .dout(n297));
  jand g00103(.dina(n290), .dinb(n297), .dout(n298));
  jand g00104(.dina(n277), .dinb(asqrt[63] ), .dout(n299));
  jand g00105(.dina(n299), .dinb(n242), .dout(n300));
  jor  g00106(.dina(n300), .dinb(n290), .dout(n301));
  jnot g00107(.din(n301), .dout(n302));
  jor  g00108(.dina(n302), .dinb(n298), .dout(n303));
  jand g00109(.dina(n303), .dinb(n296), .dout(n304));
  jand g00110(.dina(n304), .dinb(n295), .dout(n305));
  jnot g00111(.din(n305), .dout(asqrt[59] ));
  jor  g00112(.dina(n305), .dinb(n261), .dout(n307));
  jnot g00113(.din(a[116] ), .dout(n308));
  jnot g00114(.din(a[117] ), .dout(n309));
  jand g00115(.dina(n261), .dinb(n309), .dout(n310));
  jand g00116(.dina(n310), .dinb(n308), .dout(n311));
  jnot g00117(.din(n311), .dout(n312));
  jand g00118(.dina(n312), .dinb(n307), .dout(n313));
  jor  g00119(.dina(n313), .dinb(n290), .dout(n314));
  jor  g00120(.dina(n305), .dinb(a[118] ), .dout(n315));
  jxor g00121(.dina(n315), .dinb(n262), .dout(n316));
  jand g00122(.dina(n313), .dinb(n290), .dout(n317));
  jor  g00123(.dina(n317), .dinb(n316), .dout(n318));
  jand g00124(.dina(n318), .dinb(n314), .dout(n319));
  jor  g00125(.dina(n319), .dinb(n223), .dout(n320));
  jand g00126(.dina(n314), .dinb(n223), .dout(n321));
  jand g00127(.dina(n321), .dinb(n318), .dout(n322));
  jor  g00128(.dina(n315), .dinb(a[119] ), .dout(n323));
  jnot g00129(.din(n295), .dout(n324));
  jnot g00130(.din(n296), .dout(n325));
  jor  g00131(.dina(n301), .dinb(n325), .dout(n326));
  jor  g00132(.dina(n326), .dinb(n324), .dout(n327));
  jand g00133(.dina(n327), .dinb(n323), .dout(n328));
  jxor g00134(.dina(n328), .dinb(n231), .dout(n329));
  jor  g00135(.dina(n329), .dinb(n322), .dout(n330));
  jand g00136(.dina(n330), .dinb(n320), .dout(n331));
  jor  g00137(.dina(n331), .dinb(n199), .dout(n332));
  jand g00138(.dina(n331), .dinb(n199), .dout(n333));
  jxor g00139(.dina(n265), .dinb(n223), .dout(n334));
  jor  g00140(.dina(n334), .dinb(n305), .dout(n335));
  jxor g00141(.dina(n335), .dinb(n268), .dout(n336));
  jor  g00142(.dina(n336), .dinb(n333), .dout(n337));
  jand g00143(.dina(n337), .dinb(n332), .dout(n338));
  jnot g00144(.din(n274), .dout(n339));
  jor  g00145(.dina(n339), .dinb(n272), .dout(n340));
  jor  g00146(.dina(n340), .dinb(n305), .dout(n341));
  jxor g00147(.dina(n341), .dinb(n283), .dout(n342));
  jand g00148(.dina(n289), .dinb(n285), .dout(n343));
  jand g00149(.dina(n343), .dinb(asqrt[59] ), .dout(n344));
  jor  g00150(.dina(n344), .dinb(n325), .dout(n345));
  jor  g00151(.dina(n345), .dinb(n342), .dout(n346));
  jor  g00152(.dina(n346), .dinb(n338), .dout(n347));
  jand g00153(.dina(n347), .dinb(n194), .dout(n348));
  jand g00154(.dina(n342), .dinb(n338), .dout(n349));
  jnot g00155(.din(n289), .dout(n350));
  jnot g00156(.din(n285), .dout(n351));
  jand g00157(.dina(asqrt[59] ), .dinb(n351), .dout(n352));
  jor  g00158(.dina(n352), .dinb(n350), .dout(n353));
  jnot g00159(.din(n353), .dout(n354));
  jand g00160(.dina(n296), .dinb(asqrt[63] ), .dout(n355));
  jnot g00161(.din(n355), .dout(n356));
  jand g00162(.dina(n356), .dinb(asqrt[59] ), .dout(n357));
  jor  g00163(.dina(n357), .dinb(n354), .dout(n358));
  jnot g00164(.din(n358), .dout(n359));
  jor  g00165(.dina(n359), .dinb(n349), .dout(n360));
  jor  g00166(.dina(n360), .dinb(n348), .dout(asqrt[58] ));
  jand g00167(.dina(asqrt[58] ), .dinb(a[116] ), .dout(n362));
  jnot g00168(.din(a[114] ), .dout(n363));
  jnot g00169(.din(a[115] ), .dout(n364));
  jand g00170(.dina(n308), .dinb(n364), .dout(n365));
  jand g00171(.dina(n365), .dinb(n363), .dout(n366));
  jor  g00172(.dina(n366), .dinb(n362), .dout(n367));
  jand g00173(.dina(n367), .dinb(asqrt[59] ), .dout(n368));
  jand g00174(.dina(asqrt[58] ), .dinb(n308), .dout(n369));
  jxor g00175(.dina(n369), .dinb(n309), .dout(n370));
  jor  g00176(.dina(n367), .dinb(asqrt[59] ), .dout(n371));
  jand g00177(.dina(n371), .dinb(n370), .dout(n372));
  jor  g00178(.dina(n372), .dinb(n368), .dout(n373));
  jand g00179(.dina(n373), .dinb(asqrt[60] ), .dout(n374));
  jor  g00180(.dina(n368), .dinb(asqrt[60] ), .dout(n375));
  jor  g00181(.dina(n375), .dinb(n372), .dout(n376));
  jand g00182(.dina(n369), .dinb(n309), .dout(n377));
  jnot g00183(.din(n348), .dout(n378));
  jnot g00184(.din(n349), .dout(n379));
  jand g00185(.dina(n358), .dinb(asqrt[59] ), .dout(n381));
  jand g00186(.dina(n381), .dinb(n379), .dout(n382));
  jand g00187(.dina(n382), .dinb(n378), .dout(n383));
  jor  g00188(.dina(n383), .dinb(n377), .dout(n384));
  jxor g00189(.dina(n384), .dinb(n261), .dout(n385));
  jand g00190(.dina(n385), .dinb(n376), .dout(n386));
  jor  g00191(.dina(n386), .dinb(n374), .dout(n387));
  jand g00192(.dina(n387), .dinb(asqrt[61] ), .dout(n388));
  jor  g00193(.dina(n387), .dinb(asqrt[61] ), .dout(n389));
  jxor g00194(.dina(n313), .dinb(n290), .dout(n390));
  jand g00195(.dina(n390), .dinb(asqrt[58] ), .dout(n391));
  jxor g00196(.dina(n391), .dinb(n316), .dout(n392));
  jnot g00197(.din(n392), .dout(n393));
  jand g00198(.dina(n393), .dinb(n389), .dout(n394));
  jor  g00199(.dina(n394), .dinb(n388), .dout(n395));
  jand g00200(.dina(n395), .dinb(asqrt[62] ), .dout(n396));
  jnot g00201(.din(n322), .dout(n397));
  jand g00202(.dina(n397), .dinb(n320), .dout(n398));
  jand g00203(.dina(n398), .dinb(asqrt[58] ), .dout(n399));
  jxor g00204(.dina(n399), .dinb(n329), .dout(n400));
  jnot g00205(.din(n400), .dout(n401));
  jor  g00206(.dina(n388), .dinb(asqrt[62] ), .dout(n402));
  jor  g00207(.dina(n402), .dinb(n394), .dout(n403));
  jand g00208(.dina(n403), .dinb(n401), .dout(n404));
  jor  g00209(.dina(n404), .dinb(n396), .dout(n405));
  jxor g00210(.dina(n331), .dinb(n199), .dout(n406));
  jand g00211(.dina(n406), .dinb(asqrt[58] ), .dout(n407));
  jxor g00212(.dina(n407), .dinb(n336), .dout(n408));
  jnot g00213(.din(n338), .dout(n409));
  jnot g00214(.din(n342), .dout(n410));
  jand g00215(.dina(asqrt[58] ), .dinb(n410), .dout(n411));
  jand g00216(.dina(n411), .dinb(n409), .dout(n412));
  jor  g00217(.dina(n412), .dinb(n349), .dout(n413));
  jor  g00218(.dina(n413), .dinb(n408), .dout(n414));
  jnot g00219(.din(n414), .dout(n415));
  jand g00220(.dina(n415), .dinb(n405), .dout(n416));
  jor  g00221(.dina(n416), .dinb(asqrt[63] ), .dout(n417));
  jnot g00222(.din(n408), .dout(n418));
  jor  g00223(.dina(n418), .dinb(n405), .dout(n419));
  jor  g00224(.dina(n411), .dinb(n409), .dout(n420));
  jand g00225(.dina(n410), .dinb(n409), .dout(n421));
  jor  g00226(.dina(n421), .dinb(n194), .dout(n422));
  jnot g00227(.din(n422), .dout(n423));
  jand g00228(.dina(n423), .dinb(n420), .dout(n424));
  jnot g00229(.din(asqrt[58] ), .dout(n425));
  jnot g00230(.din(n424), .dout(n428));
  jand g00231(.dina(n428), .dinb(n419), .dout(n429));
  jand g00232(.dina(n429), .dinb(n417), .dout(n430));
  jnot g00233(.din(n430), .dout(asqrt[57] ));
  jor  g00234(.dina(n430), .dinb(n363), .dout(n432));
  jnot g00235(.din(a[112] ), .dout(n433));
  jnot g00236(.din(a[113] ), .dout(n434));
  jand g00237(.dina(n363), .dinb(n434), .dout(n435));
  jand g00238(.dina(n435), .dinb(n433), .dout(n436));
  jnot g00239(.din(n436), .dout(n437));
  jand g00240(.dina(n437), .dinb(n432), .dout(n438));
  jor  g00241(.dina(n438), .dinb(n425), .dout(n439));
  jor  g00242(.dina(n430), .dinb(a[114] ), .dout(n440));
  jxor g00243(.dina(n440), .dinb(n364), .dout(n441));
  jand g00244(.dina(n438), .dinb(n425), .dout(n442));
  jor  g00245(.dina(n442), .dinb(n441), .dout(n443));
  jand g00246(.dina(n443), .dinb(n439), .dout(n444));
  jor  g00247(.dina(n444), .dinb(n305), .dout(n445));
  jand g00248(.dina(n439), .dinb(n305), .dout(n446));
  jand g00249(.dina(n446), .dinb(n443), .dout(n447));
  jor  g00250(.dina(n440), .dinb(a[115] ), .dout(n448));
  jnot g00251(.din(n417), .dout(n449));
  jnot g00252(.din(n419), .dout(n450));
  jor  g00253(.dina(n424), .dinb(n425), .dout(n451));
  jor  g00254(.dina(n451), .dinb(n450), .dout(n452));
  jor  g00255(.dina(n452), .dinb(n449), .dout(n453));
  jand g00256(.dina(n453), .dinb(n448), .dout(n454));
  jxor g00257(.dina(n454), .dinb(n308), .dout(n455));
  jor  g00258(.dina(n455), .dinb(n447), .dout(n456));
  jand g00259(.dina(n456), .dinb(n445), .dout(n457));
  jor  g00260(.dina(n457), .dinb(n290), .dout(n458));
  jand g00261(.dina(n457), .dinb(n290), .dout(n459));
  jxor g00262(.dina(n367), .dinb(n305), .dout(n460));
  jor  g00263(.dina(n460), .dinb(n430), .dout(n461));
  jxor g00264(.dina(n461), .dinb(n370), .dout(n462));
  jor  g00265(.dina(n462), .dinb(n459), .dout(n463));
  jand g00266(.dina(n463), .dinb(n458), .dout(n464));
  jor  g00267(.dina(n464), .dinb(n223), .dout(n465));
  jnot g00268(.din(n376), .dout(n466));
  jor  g00269(.dina(n466), .dinb(n374), .dout(n467));
  jor  g00270(.dina(n467), .dinb(n430), .dout(n468));
  jxor g00271(.dina(n468), .dinb(n385), .dout(n469));
  jand g00272(.dina(n458), .dinb(n223), .dout(n470));
  jand g00273(.dina(n470), .dinb(n463), .dout(n471));
  jor  g00274(.dina(n471), .dinb(n469), .dout(n472));
  jand g00275(.dina(n472), .dinb(n465), .dout(n473));
  jor  g00276(.dina(n473), .dinb(n199), .dout(n474));
  jand g00277(.dina(n473), .dinb(n199), .dout(n475));
  jxor g00278(.dina(n387), .dinb(n223), .dout(n476));
  jor  g00279(.dina(n476), .dinb(n430), .dout(n477));
  jxor g00280(.dina(n477), .dinb(n392), .dout(n478));
  jnot g00281(.din(n478), .dout(n479));
  jor  g00282(.dina(n479), .dinb(n475), .dout(n480));
  jand g00283(.dina(n480), .dinb(n474), .dout(n481));
  jnot g00284(.din(n396), .dout(n482));
  jand g00285(.dina(asqrt[57] ), .dinb(n482), .dout(n483));
  jand g00286(.dina(n483), .dinb(n403), .dout(n484));
  jor  g00287(.dina(n484), .dinb(n401), .dout(n485));
  jand g00288(.dina(n483), .dinb(n404), .dout(n486));
  jnot g00289(.din(n486), .dout(n487));
  jand g00290(.dina(n487), .dinb(n485), .dout(n488));
  jnot g00291(.din(n488), .dout(n489));
  jand g00292(.dina(asqrt[57] ), .dinb(n418), .dout(n490));
  jand g00293(.dina(n490), .dinb(n405), .dout(n491));
  jor  g00294(.dina(n491), .dinb(n450), .dout(n492));
  jor  g00295(.dina(n492), .dinb(n489), .dout(n493));
  jor  g00296(.dina(n493), .dinb(n481), .dout(n494));
  jand g00297(.dina(n494), .dinb(n194), .dout(n495));
  jand g00298(.dina(n489), .dinb(n481), .dout(n496));
  jor  g00299(.dina(n490), .dinb(n405), .dout(n497));
  jand g00300(.dina(n418), .dinb(n405), .dout(n498));
  jor  g00301(.dina(n498), .dinb(n194), .dout(n499));
  jnot g00302(.din(n499), .dout(n500));
  jand g00303(.dina(n500), .dinb(n497), .dout(n501));
  jor  g00304(.dina(n501), .dinb(n496), .dout(n504));
  jor  g00305(.dina(n504), .dinb(n495), .dout(asqrt[56] ));
  jand g00306(.dina(asqrt[56] ), .dinb(a[112] ), .dout(n506));
  jnot g00307(.din(a[110] ), .dout(n507));
  jnot g00308(.din(a[111] ), .dout(n508));
  jand g00309(.dina(n433), .dinb(n508), .dout(n509));
  jand g00310(.dina(n509), .dinb(n507), .dout(n510));
  jor  g00311(.dina(n510), .dinb(n506), .dout(n511));
  jand g00312(.dina(n511), .dinb(asqrt[57] ), .dout(n512));
  jand g00313(.dina(asqrt[56] ), .dinb(n433), .dout(n513));
  jxor g00314(.dina(n513), .dinb(n434), .dout(n514));
  jor  g00315(.dina(n511), .dinb(asqrt[57] ), .dout(n515));
  jand g00316(.dina(n515), .dinb(n514), .dout(n516));
  jor  g00317(.dina(n516), .dinb(n512), .dout(n517));
  jand g00318(.dina(n517), .dinb(asqrt[58] ), .dout(n518));
  jor  g00319(.dina(n512), .dinb(asqrt[58] ), .dout(n519));
  jor  g00320(.dina(n519), .dinb(n516), .dout(n520));
  jand g00321(.dina(n513), .dinb(n434), .dout(n521));
  jnot g00322(.din(n495), .dout(n522));
  jnot g00323(.din(n496), .dout(n523));
  jnot g00324(.din(n501), .dout(n524));
  jand g00325(.dina(n524), .dinb(asqrt[57] ), .dout(n525));
  jand g00326(.dina(n525), .dinb(n523), .dout(n526));
  jand g00327(.dina(n526), .dinb(n522), .dout(n527));
  jor  g00328(.dina(n527), .dinb(n521), .dout(n528));
  jxor g00329(.dina(n528), .dinb(n363), .dout(n529));
  jand g00330(.dina(n529), .dinb(n520), .dout(n530));
  jor  g00331(.dina(n530), .dinb(n518), .dout(n531));
  jand g00332(.dina(n531), .dinb(asqrt[59] ), .dout(n532));
  jor  g00333(.dina(n531), .dinb(asqrt[59] ), .dout(n533));
  jxor g00334(.dina(n438), .dinb(n425), .dout(n534));
  jand g00335(.dina(n534), .dinb(asqrt[56] ), .dout(n535));
  jxor g00336(.dina(n535), .dinb(n441), .dout(n536));
  jnot g00337(.din(n536), .dout(n537));
  jand g00338(.dina(n537), .dinb(n533), .dout(n538));
  jor  g00339(.dina(n538), .dinb(n532), .dout(n539));
  jand g00340(.dina(n539), .dinb(asqrt[60] ), .dout(n540));
  jnot g00341(.din(n447), .dout(n541));
  jand g00342(.dina(n541), .dinb(n445), .dout(n542));
  jand g00343(.dina(n542), .dinb(asqrt[56] ), .dout(n543));
  jxor g00344(.dina(n543), .dinb(n455), .dout(n544));
  jnot g00345(.din(n544), .dout(n545));
  jor  g00346(.dina(n532), .dinb(asqrt[60] ), .dout(n546));
  jor  g00347(.dina(n546), .dinb(n538), .dout(n547));
  jand g00348(.dina(n547), .dinb(n545), .dout(n548));
  jor  g00349(.dina(n548), .dinb(n540), .dout(n549));
  jand g00350(.dina(n549), .dinb(asqrt[61] ), .dout(n550));
  jor  g00351(.dina(n549), .dinb(asqrt[61] ), .dout(n551));
  jnot g00352(.din(n462), .dout(n552));
  jxor g00353(.dina(n457), .dinb(n290), .dout(n553));
  jand g00354(.dina(n553), .dinb(asqrt[56] ), .dout(n554));
  jxor g00355(.dina(n554), .dinb(n552), .dout(n555));
  jand g00356(.dina(n555), .dinb(n551), .dout(n556));
  jor  g00357(.dina(n556), .dinb(n550), .dout(n557));
  jand g00358(.dina(n557), .dinb(asqrt[62] ), .dout(n558));
  jor  g00359(.dina(n550), .dinb(asqrt[62] ), .dout(n559));
  jor  g00360(.dina(n559), .dinb(n556), .dout(n560));
  jnot g00361(.din(n469), .dout(n561));
  jnot g00362(.din(n471), .dout(n562));
  jand g00363(.dina(asqrt[56] ), .dinb(n465), .dout(n563));
  jand g00364(.dina(n563), .dinb(n562), .dout(n564));
  jor  g00365(.dina(n564), .dinb(n561), .dout(n565));
  jnot g00366(.din(n472), .dout(n566));
  jand g00367(.dina(n563), .dinb(n566), .dout(n567));
  jnot g00368(.din(n567), .dout(n568));
  jand g00369(.dina(n568), .dinb(n565), .dout(n569));
  jand g00370(.dina(n569), .dinb(n560), .dout(n570));
  jor  g00371(.dina(n570), .dinb(n558), .dout(n571));
  jxor g00372(.dina(n473), .dinb(n199), .dout(n572));
  jand g00373(.dina(n572), .dinb(asqrt[56] ), .dout(n573));
  jxor g00374(.dina(n573), .dinb(n478), .dout(n574));
  jnot g00375(.din(n574), .dout(n575));
  jnot g00376(.din(n481), .dout(n576));
  jand g00377(.dina(asqrt[56] ), .dinb(n488), .dout(n577));
  jand g00378(.dina(n577), .dinb(n576), .dout(n578));
  jor  g00379(.dina(n578), .dinb(n496), .dout(n579));
  jor  g00380(.dina(n579), .dinb(n575), .dout(n580));
  jnot g00381(.din(n580), .dout(n581));
  jand g00382(.dina(n581), .dinb(n571), .dout(n582));
  jor  g00383(.dina(n582), .dinb(asqrt[63] ), .dout(n583));
  jor  g00384(.dina(n574), .dinb(n571), .dout(n584));
  jor  g00385(.dina(n577), .dinb(n576), .dout(n585));
  jand g00386(.dina(n488), .dinb(n576), .dout(n586));
  jor  g00387(.dina(n586), .dinb(n194), .dout(n587));
  jnot g00388(.din(n587), .dout(n588));
  jand g00389(.dina(n588), .dinb(n585), .dout(n589));
  jnot g00390(.din(asqrt[56] ), .dout(n590));
  jnot g00391(.din(n589), .dout(n593));
  jand g00392(.dina(n593), .dinb(n584), .dout(n594));
  jand g00393(.dina(n594), .dinb(n583), .dout(n595));
  jnot g00394(.din(n595), .dout(asqrt[55] ));
  jor  g00395(.dina(n595), .dinb(n507), .dout(n597));
  jnot g00396(.din(a[108] ), .dout(n598));
  jnot g00397(.din(a[109] ), .dout(n599));
  jand g00398(.dina(n507), .dinb(n599), .dout(n600));
  jand g00399(.dina(n600), .dinb(n598), .dout(n601));
  jnot g00400(.din(n601), .dout(n602));
  jand g00401(.dina(n602), .dinb(n597), .dout(n603));
  jor  g00402(.dina(n603), .dinb(n590), .dout(n604));
  jor  g00403(.dina(n595), .dinb(a[110] ), .dout(n605));
  jxor g00404(.dina(n605), .dinb(n508), .dout(n606));
  jand g00405(.dina(n603), .dinb(n590), .dout(n607));
  jor  g00406(.dina(n607), .dinb(n606), .dout(n608));
  jand g00407(.dina(n608), .dinb(n604), .dout(n609));
  jor  g00408(.dina(n609), .dinb(n430), .dout(n610));
  jand g00409(.dina(n604), .dinb(n430), .dout(n611));
  jand g00410(.dina(n611), .dinb(n608), .dout(n612));
  jor  g00411(.dina(n605), .dinb(a[111] ), .dout(n613));
  jnot g00412(.din(n583), .dout(n614));
  jnot g00413(.din(n584), .dout(n615));
  jor  g00414(.dina(n589), .dinb(n590), .dout(n616));
  jor  g00415(.dina(n616), .dinb(n615), .dout(n617));
  jor  g00416(.dina(n617), .dinb(n614), .dout(n618));
  jand g00417(.dina(n618), .dinb(n613), .dout(n619));
  jxor g00418(.dina(n619), .dinb(n433), .dout(n620));
  jor  g00419(.dina(n620), .dinb(n612), .dout(n621));
  jand g00420(.dina(n621), .dinb(n610), .dout(n622));
  jor  g00421(.dina(n622), .dinb(n425), .dout(n623));
  jand g00422(.dina(n622), .dinb(n425), .dout(n624));
  jxor g00423(.dina(n511), .dinb(n430), .dout(n625));
  jor  g00424(.dina(n625), .dinb(n595), .dout(n626));
  jxor g00425(.dina(n626), .dinb(n514), .dout(n627));
  jor  g00426(.dina(n627), .dinb(n624), .dout(n628));
  jand g00427(.dina(n628), .dinb(n623), .dout(n629));
  jor  g00428(.dina(n629), .dinb(n305), .dout(n630));
  jnot g00429(.din(n520), .dout(n631));
  jor  g00430(.dina(n631), .dinb(n518), .dout(n632));
  jor  g00431(.dina(n632), .dinb(n595), .dout(n633));
  jxor g00432(.dina(n633), .dinb(n529), .dout(n634));
  jand g00433(.dina(n623), .dinb(n305), .dout(n635));
  jand g00434(.dina(n635), .dinb(n628), .dout(n636));
  jor  g00435(.dina(n636), .dinb(n634), .dout(n637));
  jand g00436(.dina(n637), .dinb(n630), .dout(n638));
  jor  g00437(.dina(n638), .dinb(n290), .dout(n639));
  jand g00438(.dina(n638), .dinb(n290), .dout(n640));
  jxor g00439(.dina(n531), .dinb(n305), .dout(n641));
  jor  g00440(.dina(n641), .dinb(n595), .dout(n642));
  jxor g00441(.dina(n642), .dinb(n536), .dout(n643));
  jnot g00442(.din(n643), .dout(n644));
  jor  g00443(.dina(n644), .dinb(n640), .dout(n645));
  jand g00444(.dina(n645), .dinb(n639), .dout(n646));
  jor  g00445(.dina(n646), .dinb(n223), .dout(n647));
  jand g00446(.dina(n639), .dinb(n223), .dout(n648));
  jand g00447(.dina(n648), .dinb(n645), .dout(n649));
  jnot g00448(.din(n540), .dout(n650));
  jand g00449(.dina(asqrt[55] ), .dinb(n650), .dout(n651));
  jand g00450(.dina(n651), .dinb(n547), .dout(n652));
  jor  g00451(.dina(n652), .dinb(n545), .dout(n653));
  jand g00452(.dina(n651), .dinb(n548), .dout(n654));
  jnot g00453(.din(n654), .dout(n655));
  jand g00454(.dina(n655), .dinb(n653), .dout(n656));
  jnot g00455(.din(n656), .dout(n657));
  jor  g00456(.dina(n657), .dinb(n649), .dout(n658));
  jand g00457(.dina(n658), .dinb(n647), .dout(n659));
  jor  g00458(.dina(n659), .dinb(n199), .dout(n660));
  jand g00459(.dina(n659), .dinb(n199), .dout(n661));
  jnot g00460(.din(n555), .dout(n662));
  jxor g00461(.dina(n549), .dinb(n223), .dout(n663));
  jor  g00462(.dina(n663), .dinb(n595), .dout(n664));
  jxor g00463(.dina(n664), .dinb(n662), .dout(n665));
  jnot g00464(.din(n665), .dout(n666));
  jor  g00465(.dina(n666), .dinb(n661), .dout(n667));
  jand g00466(.dina(n667), .dinb(n660), .dout(n668));
  jnot g00467(.din(n560), .dout(n669));
  jor  g00468(.dina(n669), .dinb(n558), .dout(n670));
  jor  g00469(.dina(n670), .dinb(n595), .dout(n671));
  jxor g00470(.dina(n671), .dinb(n569), .dout(n672));
  jand g00471(.dina(asqrt[55] ), .dinb(n574), .dout(n673));
  jand g00472(.dina(n673), .dinb(n571), .dout(n674));
  jor  g00473(.dina(n674), .dinb(n615), .dout(n675));
  jor  g00474(.dina(n675), .dinb(n672), .dout(n676));
  jor  g00475(.dina(n676), .dinb(n668), .dout(n677));
  jand g00476(.dina(n677), .dinb(n194), .dout(n678));
  jand g00477(.dina(n672), .dinb(n668), .dout(n679));
  jor  g00478(.dina(n673), .dinb(n571), .dout(n680));
  jand g00479(.dina(n574), .dinb(n571), .dout(n681));
  jor  g00480(.dina(n681), .dinb(n194), .dout(n682));
  jnot g00481(.din(n682), .dout(n683));
  jand g00482(.dina(n683), .dinb(n680), .dout(n684));
  jor  g00483(.dina(n684), .dinb(n679), .dout(n687));
  jor  g00484(.dina(n687), .dinb(n678), .dout(asqrt[54] ));
  jand g00485(.dina(asqrt[54] ), .dinb(a[108] ), .dout(n689));
  jnot g00486(.din(a[106] ), .dout(n690));
  jnot g00487(.din(a[107] ), .dout(n691));
  jand g00488(.dina(n598), .dinb(n691), .dout(n692));
  jand g00489(.dina(n692), .dinb(n690), .dout(n693));
  jor  g00490(.dina(n693), .dinb(n689), .dout(n694));
  jand g00491(.dina(n694), .dinb(asqrt[55] ), .dout(n695));
  jand g00492(.dina(asqrt[54] ), .dinb(n598), .dout(n696));
  jxor g00493(.dina(n696), .dinb(n599), .dout(n697));
  jor  g00494(.dina(n694), .dinb(asqrt[55] ), .dout(n698));
  jand g00495(.dina(n698), .dinb(n697), .dout(n699));
  jor  g00496(.dina(n699), .dinb(n695), .dout(n700));
  jand g00497(.dina(n700), .dinb(asqrt[56] ), .dout(n701));
  jor  g00498(.dina(n695), .dinb(asqrt[56] ), .dout(n702));
  jor  g00499(.dina(n702), .dinb(n699), .dout(n703));
  jand g00500(.dina(n696), .dinb(n599), .dout(n704));
  jnot g00501(.din(n678), .dout(n705));
  jnot g00502(.din(n679), .dout(n706));
  jnot g00503(.din(n684), .dout(n707));
  jand g00504(.dina(n707), .dinb(asqrt[55] ), .dout(n708));
  jand g00505(.dina(n708), .dinb(n706), .dout(n709));
  jand g00506(.dina(n709), .dinb(n705), .dout(n710));
  jor  g00507(.dina(n710), .dinb(n704), .dout(n711));
  jxor g00508(.dina(n711), .dinb(n507), .dout(n712));
  jand g00509(.dina(n712), .dinb(n703), .dout(n713));
  jor  g00510(.dina(n713), .dinb(n701), .dout(n714));
  jand g00511(.dina(n714), .dinb(asqrt[57] ), .dout(n715));
  jor  g00512(.dina(n714), .dinb(asqrt[57] ), .dout(n716));
  jxor g00513(.dina(n603), .dinb(n590), .dout(n717));
  jand g00514(.dina(n717), .dinb(asqrt[54] ), .dout(n718));
  jxor g00515(.dina(n718), .dinb(n606), .dout(n719));
  jnot g00516(.din(n719), .dout(n720));
  jand g00517(.dina(n720), .dinb(n716), .dout(n721));
  jor  g00518(.dina(n721), .dinb(n715), .dout(n722));
  jand g00519(.dina(n722), .dinb(asqrt[58] ), .dout(n723));
  jnot g00520(.din(n612), .dout(n724));
  jand g00521(.dina(n724), .dinb(n610), .dout(n725));
  jand g00522(.dina(n725), .dinb(asqrt[54] ), .dout(n726));
  jxor g00523(.dina(n726), .dinb(n620), .dout(n727));
  jnot g00524(.din(n727), .dout(n728));
  jor  g00525(.dina(n715), .dinb(asqrt[58] ), .dout(n729));
  jor  g00526(.dina(n729), .dinb(n721), .dout(n730));
  jand g00527(.dina(n730), .dinb(n728), .dout(n731));
  jor  g00528(.dina(n731), .dinb(n723), .dout(n732));
  jand g00529(.dina(n732), .dinb(asqrt[59] ), .dout(n733));
  jor  g00530(.dina(n732), .dinb(asqrt[59] ), .dout(n734));
  jnot g00531(.din(n627), .dout(n735));
  jxor g00532(.dina(n622), .dinb(n425), .dout(n736));
  jand g00533(.dina(n736), .dinb(asqrt[54] ), .dout(n737));
  jxor g00534(.dina(n737), .dinb(n735), .dout(n738));
  jand g00535(.dina(n738), .dinb(n734), .dout(n739));
  jor  g00536(.dina(n739), .dinb(n733), .dout(n740));
  jand g00537(.dina(n740), .dinb(asqrt[60] ), .dout(n741));
  jor  g00538(.dina(n733), .dinb(asqrt[60] ), .dout(n742));
  jor  g00539(.dina(n742), .dinb(n739), .dout(n743));
  jnot g00540(.din(n634), .dout(n744));
  jnot g00541(.din(n636), .dout(n745));
  jand g00542(.dina(asqrt[54] ), .dinb(n630), .dout(n746));
  jand g00543(.dina(n746), .dinb(n745), .dout(n747));
  jor  g00544(.dina(n747), .dinb(n744), .dout(n748));
  jnot g00545(.din(n637), .dout(n749));
  jand g00546(.dina(n746), .dinb(n749), .dout(n750));
  jnot g00547(.din(n750), .dout(n751));
  jand g00548(.dina(n751), .dinb(n748), .dout(n752));
  jand g00549(.dina(n752), .dinb(n743), .dout(n753));
  jor  g00550(.dina(n753), .dinb(n741), .dout(n754));
  jand g00551(.dina(n754), .dinb(asqrt[61] ), .dout(n755));
  jor  g00552(.dina(n754), .dinb(asqrt[61] ), .dout(n756));
  jxor g00553(.dina(n638), .dinb(n290), .dout(n757));
  jand g00554(.dina(n757), .dinb(asqrt[54] ), .dout(n758));
  jxor g00555(.dina(n758), .dinb(n643), .dout(n759));
  jand g00556(.dina(n759), .dinb(n756), .dout(n760));
  jor  g00557(.dina(n760), .dinb(n755), .dout(n761));
  jand g00558(.dina(n761), .dinb(asqrt[62] ), .dout(n762));
  jnot g00559(.din(n649), .dout(n763));
  jand g00560(.dina(n763), .dinb(n647), .dout(n764));
  jand g00561(.dina(n764), .dinb(asqrt[54] ), .dout(n765));
  jxor g00562(.dina(n765), .dinb(n657), .dout(n766));
  jnot g00563(.din(n766), .dout(n767));
  jor  g00564(.dina(n755), .dinb(asqrt[62] ), .dout(n768));
  jor  g00565(.dina(n768), .dinb(n760), .dout(n769));
  jand g00566(.dina(n769), .dinb(n767), .dout(n770));
  jor  g00567(.dina(n770), .dinb(n762), .dout(n771));
  jxor g00568(.dina(n659), .dinb(n199), .dout(n772));
  jand g00569(.dina(n772), .dinb(asqrt[54] ), .dout(n773));
  jxor g00570(.dina(n773), .dinb(n665), .dout(n774));
  jnot g00571(.din(n774), .dout(n775));
  jnot g00572(.din(n668), .dout(n776));
  jnot g00573(.din(n672), .dout(n777));
  jand g00574(.dina(asqrt[54] ), .dinb(n777), .dout(n778));
  jand g00575(.dina(n778), .dinb(n776), .dout(n779));
  jor  g00576(.dina(n779), .dinb(n679), .dout(n780));
  jor  g00577(.dina(n780), .dinb(n775), .dout(n781));
  jnot g00578(.din(n781), .dout(n782));
  jand g00579(.dina(n782), .dinb(n771), .dout(n783));
  jor  g00580(.dina(n783), .dinb(asqrt[63] ), .dout(n784));
  jor  g00581(.dina(n774), .dinb(n771), .dout(n785));
  jor  g00582(.dina(n778), .dinb(n776), .dout(n786));
  jand g00583(.dina(n777), .dinb(n776), .dout(n787));
  jor  g00584(.dina(n787), .dinb(n194), .dout(n788));
  jnot g00585(.din(n788), .dout(n789));
  jand g00586(.dina(n789), .dinb(n786), .dout(n790));
  jnot g00587(.din(asqrt[54] ), .dout(n791));
  jnot g00588(.din(n790), .dout(n794));
  jand g00589(.dina(n794), .dinb(n785), .dout(n795));
  jand g00590(.dina(n795), .dinb(n784), .dout(n796));
  jnot g00591(.din(n796), .dout(asqrt[53] ));
  jor  g00592(.dina(n796), .dinb(n690), .dout(n798));
  jnot g00593(.din(a[104] ), .dout(n799));
  jnot g00594(.din(a[105] ), .dout(n800));
  jand g00595(.dina(n690), .dinb(n800), .dout(n801));
  jand g00596(.dina(n801), .dinb(n799), .dout(n802));
  jnot g00597(.din(n802), .dout(n803));
  jand g00598(.dina(n803), .dinb(n798), .dout(n804));
  jor  g00599(.dina(n804), .dinb(n791), .dout(n805));
  jor  g00600(.dina(n796), .dinb(a[106] ), .dout(n806));
  jxor g00601(.dina(n806), .dinb(n691), .dout(n807));
  jand g00602(.dina(n804), .dinb(n791), .dout(n808));
  jor  g00603(.dina(n808), .dinb(n807), .dout(n809));
  jand g00604(.dina(n809), .dinb(n805), .dout(n810));
  jor  g00605(.dina(n810), .dinb(n595), .dout(n811));
  jand g00606(.dina(n805), .dinb(n595), .dout(n812));
  jand g00607(.dina(n812), .dinb(n809), .dout(n813));
  jor  g00608(.dina(n806), .dinb(a[107] ), .dout(n814));
  jnot g00609(.din(n784), .dout(n815));
  jnot g00610(.din(n785), .dout(n816));
  jor  g00611(.dina(n790), .dinb(n791), .dout(n817));
  jor  g00612(.dina(n817), .dinb(n816), .dout(n818));
  jor  g00613(.dina(n818), .dinb(n815), .dout(n819));
  jand g00614(.dina(n819), .dinb(n814), .dout(n820));
  jxor g00615(.dina(n820), .dinb(n598), .dout(n821));
  jor  g00616(.dina(n821), .dinb(n813), .dout(n822));
  jand g00617(.dina(n822), .dinb(n811), .dout(n823));
  jor  g00618(.dina(n823), .dinb(n590), .dout(n824));
  jand g00619(.dina(n823), .dinb(n590), .dout(n825));
  jxor g00620(.dina(n694), .dinb(n595), .dout(n826));
  jor  g00621(.dina(n826), .dinb(n796), .dout(n827));
  jxor g00622(.dina(n827), .dinb(n697), .dout(n828));
  jor  g00623(.dina(n828), .dinb(n825), .dout(n829));
  jand g00624(.dina(n829), .dinb(n824), .dout(n830));
  jor  g00625(.dina(n830), .dinb(n430), .dout(n831));
  jnot g00626(.din(n703), .dout(n832));
  jor  g00627(.dina(n832), .dinb(n701), .dout(n833));
  jor  g00628(.dina(n833), .dinb(n796), .dout(n834));
  jxor g00629(.dina(n834), .dinb(n712), .dout(n835));
  jand g00630(.dina(n824), .dinb(n430), .dout(n836));
  jand g00631(.dina(n836), .dinb(n829), .dout(n837));
  jor  g00632(.dina(n837), .dinb(n835), .dout(n838));
  jand g00633(.dina(n838), .dinb(n831), .dout(n839));
  jor  g00634(.dina(n839), .dinb(n425), .dout(n840));
  jand g00635(.dina(n839), .dinb(n425), .dout(n841));
  jxor g00636(.dina(n714), .dinb(n430), .dout(n842));
  jor  g00637(.dina(n842), .dinb(n796), .dout(n843));
  jxor g00638(.dina(n843), .dinb(n719), .dout(n844));
  jnot g00639(.din(n844), .dout(n845));
  jor  g00640(.dina(n845), .dinb(n841), .dout(n846));
  jand g00641(.dina(n846), .dinb(n840), .dout(n847));
  jor  g00642(.dina(n847), .dinb(n305), .dout(n848));
  jand g00643(.dina(n840), .dinb(n305), .dout(n849));
  jand g00644(.dina(n849), .dinb(n846), .dout(n850));
  jnot g00645(.din(n723), .dout(n851));
  jand g00646(.dina(asqrt[53] ), .dinb(n851), .dout(n852));
  jand g00647(.dina(n852), .dinb(n730), .dout(n853));
  jor  g00648(.dina(n853), .dinb(n728), .dout(n854));
  jand g00649(.dina(n852), .dinb(n731), .dout(n855));
  jnot g00650(.din(n855), .dout(n856));
  jand g00651(.dina(n856), .dinb(n854), .dout(n857));
  jnot g00652(.din(n857), .dout(n858));
  jor  g00653(.dina(n858), .dinb(n850), .dout(n859));
  jand g00654(.dina(n859), .dinb(n848), .dout(n860));
  jor  g00655(.dina(n860), .dinb(n290), .dout(n861));
  jand g00656(.dina(n860), .dinb(n290), .dout(n862));
  jnot g00657(.din(n738), .dout(n863));
  jxor g00658(.dina(n732), .dinb(n305), .dout(n864));
  jor  g00659(.dina(n864), .dinb(n796), .dout(n865));
  jxor g00660(.dina(n865), .dinb(n863), .dout(n866));
  jnot g00661(.din(n866), .dout(n867));
  jor  g00662(.dina(n867), .dinb(n862), .dout(n868));
  jand g00663(.dina(n868), .dinb(n861), .dout(n869));
  jor  g00664(.dina(n869), .dinb(n223), .dout(n870));
  jnot g00665(.din(n743), .dout(n871));
  jor  g00666(.dina(n871), .dinb(n741), .dout(n872));
  jor  g00667(.dina(n872), .dinb(n796), .dout(n873));
  jxor g00668(.dina(n873), .dinb(n752), .dout(n874));
  jand g00669(.dina(n861), .dinb(n223), .dout(n875));
  jand g00670(.dina(n875), .dinb(n868), .dout(n876));
  jor  g00671(.dina(n876), .dinb(n874), .dout(n877));
  jand g00672(.dina(n877), .dinb(n870), .dout(n878));
  jor  g00673(.dina(n878), .dinb(n199), .dout(n879));
  jand g00674(.dina(n878), .dinb(n199), .dout(n880));
  jnot g00675(.din(n759), .dout(n881));
  jxor g00676(.dina(n754), .dinb(n223), .dout(n882));
  jor  g00677(.dina(n882), .dinb(n796), .dout(n883));
  jxor g00678(.dina(n883), .dinb(n881), .dout(n884));
  jnot g00679(.din(n884), .dout(n885));
  jor  g00680(.dina(n885), .dinb(n880), .dout(n886));
  jand g00681(.dina(n886), .dinb(n879), .dout(n887));
  jnot g00682(.din(n762), .dout(n888));
  jand g00683(.dina(asqrt[53] ), .dinb(n888), .dout(n889));
  jand g00684(.dina(n889), .dinb(n769), .dout(n890));
  jor  g00685(.dina(n890), .dinb(n767), .dout(n891));
  jand g00686(.dina(n889), .dinb(n770), .dout(n892));
  jnot g00687(.din(n892), .dout(n893));
  jand g00688(.dina(n893), .dinb(n891), .dout(n894));
  jnot g00689(.din(n894), .dout(n895));
  jand g00690(.dina(asqrt[53] ), .dinb(n774), .dout(n896));
  jand g00691(.dina(n896), .dinb(n771), .dout(n897));
  jor  g00692(.dina(n897), .dinb(n816), .dout(n898));
  jor  g00693(.dina(n898), .dinb(n895), .dout(n899));
  jor  g00694(.dina(n899), .dinb(n887), .dout(n900));
  jand g00695(.dina(n900), .dinb(n194), .dout(n901));
  jand g00696(.dina(n895), .dinb(n887), .dout(n902));
  jor  g00697(.dina(n896), .dinb(n771), .dout(n903));
  jand g00698(.dina(n774), .dinb(n771), .dout(n904));
  jor  g00699(.dina(n904), .dinb(n194), .dout(n905));
  jnot g00700(.din(n905), .dout(n906));
  jand g00701(.dina(n906), .dinb(n903), .dout(n907));
  jor  g00702(.dina(n907), .dinb(n902), .dout(n910));
  jor  g00703(.dina(n910), .dinb(n901), .dout(asqrt[52] ));
  jand g00704(.dina(asqrt[52] ), .dinb(a[104] ), .dout(n912));
  jnot g00705(.din(a[102] ), .dout(n913));
  jnot g00706(.din(a[103] ), .dout(n914));
  jand g00707(.dina(n799), .dinb(n914), .dout(n915));
  jand g00708(.dina(n915), .dinb(n913), .dout(n916));
  jor  g00709(.dina(n916), .dinb(n912), .dout(n917));
  jand g00710(.dina(n917), .dinb(asqrt[53] ), .dout(n918));
  jand g00711(.dina(asqrt[52] ), .dinb(n799), .dout(n919));
  jxor g00712(.dina(n919), .dinb(n800), .dout(n920));
  jor  g00713(.dina(n917), .dinb(asqrt[53] ), .dout(n921));
  jand g00714(.dina(n921), .dinb(n920), .dout(n922));
  jor  g00715(.dina(n922), .dinb(n918), .dout(n923));
  jand g00716(.dina(n923), .dinb(asqrt[54] ), .dout(n924));
  jor  g00717(.dina(n918), .dinb(asqrt[54] ), .dout(n925));
  jor  g00718(.dina(n925), .dinb(n922), .dout(n926));
  jand g00719(.dina(n919), .dinb(n800), .dout(n927));
  jnot g00720(.din(n901), .dout(n928));
  jnot g00721(.din(n902), .dout(n929));
  jnot g00722(.din(n907), .dout(n930));
  jand g00723(.dina(n930), .dinb(asqrt[53] ), .dout(n931));
  jand g00724(.dina(n931), .dinb(n929), .dout(n932));
  jand g00725(.dina(n932), .dinb(n928), .dout(n933));
  jor  g00726(.dina(n933), .dinb(n927), .dout(n934));
  jxor g00727(.dina(n934), .dinb(n690), .dout(n935));
  jand g00728(.dina(n935), .dinb(n926), .dout(n936));
  jor  g00729(.dina(n936), .dinb(n924), .dout(n937));
  jand g00730(.dina(n937), .dinb(asqrt[55] ), .dout(n938));
  jor  g00731(.dina(n937), .dinb(asqrt[55] ), .dout(n939));
  jxor g00732(.dina(n804), .dinb(n791), .dout(n940));
  jand g00733(.dina(n940), .dinb(asqrt[52] ), .dout(n941));
  jxor g00734(.dina(n941), .dinb(n807), .dout(n942));
  jnot g00735(.din(n942), .dout(n943));
  jand g00736(.dina(n943), .dinb(n939), .dout(n944));
  jor  g00737(.dina(n944), .dinb(n938), .dout(n945));
  jand g00738(.dina(n945), .dinb(asqrt[56] ), .dout(n946));
  jnot g00739(.din(n813), .dout(n947));
  jand g00740(.dina(n947), .dinb(n811), .dout(n948));
  jand g00741(.dina(n948), .dinb(asqrt[52] ), .dout(n949));
  jxor g00742(.dina(n949), .dinb(n821), .dout(n950));
  jnot g00743(.din(n950), .dout(n951));
  jor  g00744(.dina(n938), .dinb(asqrt[56] ), .dout(n952));
  jor  g00745(.dina(n952), .dinb(n944), .dout(n953));
  jand g00746(.dina(n953), .dinb(n951), .dout(n954));
  jor  g00747(.dina(n954), .dinb(n946), .dout(n955));
  jand g00748(.dina(n955), .dinb(asqrt[57] ), .dout(n956));
  jor  g00749(.dina(n955), .dinb(asqrt[57] ), .dout(n957));
  jnot g00750(.din(n828), .dout(n958));
  jxor g00751(.dina(n823), .dinb(n590), .dout(n959));
  jand g00752(.dina(n959), .dinb(asqrt[52] ), .dout(n960));
  jxor g00753(.dina(n960), .dinb(n958), .dout(n961));
  jand g00754(.dina(n961), .dinb(n957), .dout(n962));
  jor  g00755(.dina(n962), .dinb(n956), .dout(n963));
  jand g00756(.dina(n963), .dinb(asqrt[58] ), .dout(n964));
  jor  g00757(.dina(n956), .dinb(asqrt[58] ), .dout(n965));
  jor  g00758(.dina(n965), .dinb(n962), .dout(n966));
  jnot g00759(.din(n835), .dout(n967));
  jnot g00760(.din(n837), .dout(n968));
  jand g00761(.dina(asqrt[52] ), .dinb(n831), .dout(n969));
  jand g00762(.dina(n969), .dinb(n968), .dout(n970));
  jor  g00763(.dina(n970), .dinb(n967), .dout(n971));
  jnot g00764(.din(n838), .dout(n972));
  jand g00765(.dina(n969), .dinb(n972), .dout(n973));
  jnot g00766(.din(n973), .dout(n974));
  jand g00767(.dina(n974), .dinb(n971), .dout(n975));
  jand g00768(.dina(n975), .dinb(n966), .dout(n976));
  jor  g00769(.dina(n976), .dinb(n964), .dout(n977));
  jand g00770(.dina(n977), .dinb(asqrt[59] ), .dout(n978));
  jor  g00771(.dina(n977), .dinb(asqrt[59] ), .dout(n979));
  jxor g00772(.dina(n839), .dinb(n425), .dout(n980));
  jand g00773(.dina(n980), .dinb(asqrt[52] ), .dout(n981));
  jxor g00774(.dina(n981), .dinb(n844), .dout(n982));
  jand g00775(.dina(n982), .dinb(n979), .dout(n983));
  jor  g00776(.dina(n983), .dinb(n978), .dout(n984));
  jand g00777(.dina(n984), .dinb(asqrt[60] ), .dout(n985));
  jnot g00778(.din(n850), .dout(n986));
  jand g00779(.dina(n986), .dinb(n848), .dout(n987));
  jand g00780(.dina(n987), .dinb(asqrt[52] ), .dout(n988));
  jxor g00781(.dina(n988), .dinb(n858), .dout(n989));
  jnot g00782(.din(n989), .dout(n990));
  jor  g00783(.dina(n978), .dinb(asqrt[60] ), .dout(n991));
  jor  g00784(.dina(n991), .dinb(n983), .dout(n992));
  jand g00785(.dina(n992), .dinb(n990), .dout(n993));
  jor  g00786(.dina(n993), .dinb(n985), .dout(n994));
  jand g00787(.dina(n994), .dinb(asqrt[61] ), .dout(n995));
  jor  g00788(.dina(n994), .dinb(asqrt[61] ), .dout(n996));
  jxor g00789(.dina(n860), .dinb(n290), .dout(n997));
  jand g00790(.dina(n997), .dinb(asqrt[52] ), .dout(n998));
  jxor g00791(.dina(n998), .dinb(n866), .dout(n999));
  jand g00792(.dina(n999), .dinb(n996), .dout(n1000));
  jor  g00793(.dina(n1000), .dinb(n995), .dout(n1001));
  jand g00794(.dina(n1001), .dinb(asqrt[62] ), .dout(n1002));
  jor  g00795(.dina(n995), .dinb(asqrt[62] ), .dout(n1003));
  jor  g00796(.dina(n1003), .dinb(n1000), .dout(n1004));
  jnot g00797(.din(n874), .dout(n1005));
  jnot g00798(.din(n876), .dout(n1006));
  jand g00799(.dina(asqrt[52] ), .dinb(n870), .dout(n1007));
  jand g00800(.dina(n1007), .dinb(n1006), .dout(n1008));
  jor  g00801(.dina(n1008), .dinb(n1005), .dout(n1009));
  jnot g00802(.din(n877), .dout(n1010));
  jand g00803(.dina(n1007), .dinb(n1010), .dout(n1011));
  jnot g00804(.din(n1011), .dout(n1012));
  jand g00805(.dina(n1012), .dinb(n1009), .dout(n1013));
  jand g00806(.dina(n1013), .dinb(n1004), .dout(n1014));
  jor  g00807(.dina(n1014), .dinb(n1002), .dout(n1015));
  jxor g00808(.dina(n878), .dinb(n199), .dout(n1016));
  jand g00809(.dina(n1016), .dinb(asqrt[52] ), .dout(n1017));
  jxor g00810(.dina(n1017), .dinb(n885), .dout(n1018));
  jnot g00811(.din(n887), .dout(n1019));
  jand g00812(.dina(asqrt[52] ), .dinb(n894), .dout(n1020));
  jand g00813(.dina(n1020), .dinb(n1019), .dout(n1021));
  jor  g00814(.dina(n1021), .dinb(n902), .dout(n1022));
  jor  g00815(.dina(n1022), .dinb(n1018), .dout(n1023));
  jnot g00816(.din(n1023), .dout(n1024));
  jand g00817(.dina(n1024), .dinb(n1015), .dout(n1025));
  jor  g00818(.dina(n1025), .dinb(asqrt[63] ), .dout(n1026));
  jnot g00819(.din(n1018), .dout(n1027));
  jor  g00820(.dina(n1027), .dinb(n1015), .dout(n1028));
  jor  g00821(.dina(n1020), .dinb(n1019), .dout(n1029));
  jand g00822(.dina(n894), .dinb(n1019), .dout(n1030));
  jor  g00823(.dina(n1030), .dinb(n194), .dout(n1031));
  jnot g00824(.din(n1031), .dout(n1032));
  jand g00825(.dina(n1032), .dinb(n1029), .dout(n1033));
  jnot g00826(.din(asqrt[52] ), .dout(n1034));
  jnot g00827(.din(n1033), .dout(n1037));
  jand g00828(.dina(n1037), .dinb(n1028), .dout(n1038));
  jand g00829(.dina(n1038), .dinb(n1026), .dout(n1039));
  jnot g00830(.din(n1039), .dout(asqrt[51] ));
  jor  g00831(.dina(n1039), .dinb(n913), .dout(n1041));
  jnot g00832(.din(a[100] ), .dout(n1042));
  jnot g00833(.din(a[101] ), .dout(n1043));
  jand g00834(.dina(n913), .dinb(n1043), .dout(n1044));
  jand g00835(.dina(n1044), .dinb(n1042), .dout(n1045));
  jnot g00836(.din(n1045), .dout(n1046));
  jand g00837(.dina(n1046), .dinb(n1041), .dout(n1047));
  jor  g00838(.dina(n1047), .dinb(n1034), .dout(n1048));
  jor  g00839(.dina(n1039), .dinb(a[102] ), .dout(n1049));
  jxor g00840(.dina(n1049), .dinb(n914), .dout(n1050));
  jand g00841(.dina(n1047), .dinb(n1034), .dout(n1051));
  jor  g00842(.dina(n1051), .dinb(n1050), .dout(n1052));
  jand g00843(.dina(n1052), .dinb(n1048), .dout(n1053));
  jor  g00844(.dina(n1053), .dinb(n796), .dout(n1054));
  jand g00845(.dina(n1048), .dinb(n796), .dout(n1055));
  jand g00846(.dina(n1055), .dinb(n1052), .dout(n1056));
  jor  g00847(.dina(n1049), .dinb(a[103] ), .dout(n1057));
  jnot g00848(.din(n1026), .dout(n1058));
  jnot g00849(.din(n1028), .dout(n1059));
  jor  g00850(.dina(n1033), .dinb(n1034), .dout(n1060));
  jor  g00851(.dina(n1060), .dinb(n1059), .dout(n1061));
  jor  g00852(.dina(n1061), .dinb(n1058), .dout(n1062));
  jand g00853(.dina(n1062), .dinb(n1057), .dout(n1063));
  jxor g00854(.dina(n1063), .dinb(n799), .dout(n1064));
  jor  g00855(.dina(n1064), .dinb(n1056), .dout(n1065));
  jand g00856(.dina(n1065), .dinb(n1054), .dout(n1066));
  jor  g00857(.dina(n1066), .dinb(n791), .dout(n1067));
  jand g00858(.dina(n1066), .dinb(n791), .dout(n1068));
  jxor g00859(.dina(n917), .dinb(n796), .dout(n1069));
  jor  g00860(.dina(n1069), .dinb(n1039), .dout(n1070));
  jxor g00861(.dina(n1070), .dinb(n920), .dout(n1071));
  jor  g00862(.dina(n1071), .dinb(n1068), .dout(n1072));
  jand g00863(.dina(n1072), .dinb(n1067), .dout(n1073));
  jor  g00864(.dina(n1073), .dinb(n595), .dout(n1074));
  jnot g00865(.din(n926), .dout(n1075));
  jor  g00866(.dina(n1075), .dinb(n924), .dout(n1076));
  jor  g00867(.dina(n1076), .dinb(n1039), .dout(n1077));
  jxor g00868(.dina(n1077), .dinb(n935), .dout(n1078));
  jand g00869(.dina(n1067), .dinb(n595), .dout(n1079));
  jand g00870(.dina(n1079), .dinb(n1072), .dout(n1080));
  jor  g00871(.dina(n1080), .dinb(n1078), .dout(n1081));
  jand g00872(.dina(n1081), .dinb(n1074), .dout(n1082));
  jor  g00873(.dina(n1082), .dinb(n590), .dout(n1083));
  jand g00874(.dina(n1082), .dinb(n590), .dout(n1084));
  jxor g00875(.dina(n937), .dinb(n595), .dout(n1085));
  jor  g00876(.dina(n1085), .dinb(n1039), .dout(n1086));
  jxor g00877(.dina(n1086), .dinb(n942), .dout(n1087));
  jnot g00878(.din(n1087), .dout(n1088));
  jor  g00879(.dina(n1088), .dinb(n1084), .dout(n1089));
  jand g00880(.dina(n1089), .dinb(n1083), .dout(n1090));
  jor  g00881(.dina(n1090), .dinb(n430), .dout(n1091));
  jand g00882(.dina(n1083), .dinb(n430), .dout(n1092));
  jand g00883(.dina(n1092), .dinb(n1089), .dout(n1093));
  jnot g00884(.din(n946), .dout(n1094));
  jand g00885(.dina(asqrt[51] ), .dinb(n1094), .dout(n1095));
  jand g00886(.dina(n1095), .dinb(n953), .dout(n1096));
  jor  g00887(.dina(n1096), .dinb(n951), .dout(n1097));
  jand g00888(.dina(n1095), .dinb(n954), .dout(n1098));
  jnot g00889(.din(n1098), .dout(n1099));
  jand g00890(.dina(n1099), .dinb(n1097), .dout(n1100));
  jnot g00891(.din(n1100), .dout(n1101));
  jor  g00892(.dina(n1101), .dinb(n1093), .dout(n1102));
  jand g00893(.dina(n1102), .dinb(n1091), .dout(n1103));
  jor  g00894(.dina(n1103), .dinb(n425), .dout(n1104));
  jand g00895(.dina(n1103), .dinb(n425), .dout(n1105));
  jnot g00896(.din(n961), .dout(n1106));
  jxor g00897(.dina(n955), .dinb(n430), .dout(n1107));
  jor  g00898(.dina(n1107), .dinb(n1039), .dout(n1108));
  jxor g00899(.dina(n1108), .dinb(n1106), .dout(n1109));
  jnot g00900(.din(n1109), .dout(n1110));
  jor  g00901(.dina(n1110), .dinb(n1105), .dout(n1111));
  jand g00902(.dina(n1111), .dinb(n1104), .dout(n1112));
  jor  g00903(.dina(n1112), .dinb(n305), .dout(n1113));
  jnot g00904(.din(n966), .dout(n1114));
  jor  g00905(.dina(n1114), .dinb(n964), .dout(n1115));
  jor  g00906(.dina(n1115), .dinb(n1039), .dout(n1116));
  jxor g00907(.dina(n1116), .dinb(n975), .dout(n1117));
  jand g00908(.dina(n1104), .dinb(n305), .dout(n1118));
  jand g00909(.dina(n1118), .dinb(n1111), .dout(n1119));
  jor  g00910(.dina(n1119), .dinb(n1117), .dout(n1120));
  jand g00911(.dina(n1120), .dinb(n1113), .dout(n1121));
  jor  g00912(.dina(n1121), .dinb(n290), .dout(n1122));
  jand g00913(.dina(n1121), .dinb(n290), .dout(n1123));
  jnot g00914(.din(n982), .dout(n1124));
  jxor g00915(.dina(n977), .dinb(n305), .dout(n1125));
  jor  g00916(.dina(n1125), .dinb(n1039), .dout(n1126));
  jxor g00917(.dina(n1126), .dinb(n1124), .dout(n1127));
  jnot g00918(.din(n1127), .dout(n1128));
  jor  g00919(.dina(n1128), .dinb(n1123), .dout(n1129));
  jand g00920(.dina(n1129), .dinb(n1122), .dout(n1130));
  jor  g00921(.dina(n1130), .dinb(n223), .dout(n1131));
  jand g00922(.dina(n1122), .dinb(n223), .dout(n1132));
  jand g00923(.dina(n1132), .dinb(n1129), .dout(n1133));
  jnot g00924(.din(n985), .dout(n1134));
  jand g00925(.dina(asqrt[51] ), .dinb(n1134), .dout(n1135));
  jand g00926(.dina(n1135), .dinb(n992), .dout(n1136));
  jor  g00927(.dina(n1136), .dinb(n990), .dout(n1137));
  jand g00928(.dina(n1135), .dinb(n993), .dout(n1138));
  jnot g00929(.din(n1138), .dout(n1139));
  jand g00930(.dina(n1139), .dinb(n1137), .dout(n1140));
  jnot g00931(.din(n1140), .dout(n1141));
  jor  g00932(.dina(n1141), .dinb(n1133), .dout(n1142));
  jand g00933(.dina(n1142), .dinb(n1131), .dout(n1143));
  jor  g00934(.dina(n1143), .dinb(n199), .dout(n1144));
  jand g00935(.dina(n1143), .dinb(n199), .dout(n1145));
  jxor g00936(.dina(n994), .dinb(n223), .dout(n1146));
  jor  g00937(.dina(n1146), .dinb(n1039), .dout(n1147));
  jxor g00938(.dina(n1147), .dinb(n999), .dout(n1148));
  jor  g00939(.dina(n1148), .dinb(n1145), .dout(n1149));
  jand g00940(.dina(n1149), .dinb(n1144), .dout(n1150));
  jnot g00941(.din(n1004), .dout(n1151));
  jor  g00942(.dina(n1151), .dinb(n1002), .dout(n1152));
  jor  g00943(.dina(n1152), .dinb(n1039), .dout(n1153));
  jxor g00944(.dina(n1153), .dinb(n1013), .dout(n1154));
  jand g00945(.dina(asqrt[51] ), .dinb(n1027), .dout(n1155));
  jand g00946(.dina(n1155), .dinb(n1015), .dout(n1156));
  jor  g00947(.dina(n1156), .dinb(n1059), .dout(n1157));
  jor  g00948(.dina(n1157), .dinb(n1154), .dout(n1158));
  jor  g00949(.dina(n1158), .dinb(n1150), .dout(n1159));
  jand g00950(.dina(n1159), .dinb(n194), .dout(n1160));
  jand g00951(.dina(n1154), .dinb(n1150), .dout(n1161));
  jor  g00952(.dina(n1155), .dinb(n1015), .dout(n1162));
  jand g00953(.dina(n1027), .dinb(n1015), .dout(n1163));
  jor  g00954(.dina(n1163), .dinb(n194), .dout(n1164));
  jnot g00955(.din(n1164), .dout(n1165));
  jand g00956(.dina(n1165), .dinb(n1162), .dout(n1166));
  jor  g00957(.dina(n1166), .dinb(n1161), .dout(n1169));
  jor  g00958(.dina(n1169), .dinb(n1160), .dout(asqrt[50] ));
  jand g00959(.dina(asqrt[50] ), .dinb(a[100] ), .dout(n1171));
  jnot g00960(.din(a[98] ), .dout(n1172));
  jnot g00961(.din(a[99] ), .dout(n1173));
  jand g00962(.dina(n1042), .dinb(n1173), .dout(n1174));
  jand g00963(.dina(n1174), .dinb(n1172), .dout(n1175));
  jor  g00964(.dina(n1175), .dinb(n1171), .dout(n1176));
  jand g00965(.dina(n1176), .dinb(asqrt[51] ), .dout(n1177));
  jand g00966(.dina(asqrt[50] ), .dinb(n1042), .dout(n1178));
  jxor g00967(.dina(n1178), .dinb(n1043), .dout(n1179));
  jor  g00968(.dina(n1176), .dinb(asqrt[51] ), .dout(n1180));
  jand g00969(.dina(n1180), .dinb(n1179), .dout(n1181));
  jor  g00970(.dina(n1181), .dinb(n1177), .dout(n1182));
  jand g00971(.dina(n1182), .dinb(asqrt[52] ), .dout(n1183));
  jor  g00972(.dina(n1177), .dinb(asqrt[52] ), .dout(n1184));
  jor  g00973(.dina(n1184), .dinb(n1181), .dout(n1185));
  jand g00974(.dina(n1178), .dinb(n1043), .dout(n1186));
  jnot g00975(.din(n1160), .dout(n1187));
  jnot g00976(.din(n1161), .dout(n1188));
  jnot g00977(.din(n1166), .dout(n1189));
  jand g00978(.dina(n1189), .dinb(asqrt[51] ), .dout(n1190));
  jand g00979(.dina(n1190), .dinb(n1188), .dout(n1191));
  jand g00980(.dina(n1191), .dinb(n1187), .dout(n1192));
  jor  g00981(.dina(n1192), .dinb(n1186), .dout(n1193));
  jxor g00982(.dina(n1193), .dinb(n913), .dout(n1194));
  jand g00983(.dina(n1194), .dinb(n1185), .dout(n1195));
  jor  g00984(.dina(n1195), .dinb(n1183), .dout(n1196));
  jand g00985(.dina(n1196), .dinb(asqrt[53] ), .dout(n1197));
  jor  g00986(.dina(n1196), .dinb(asqrt[53] ), .dout(n1198));
  jxor g00987(.dina(n1047), .dinb(n1034), .dout(n1199));
  jand g00988(.dina(n1199), .dinb(asqrt[50] ), .dout(n1200));
  jxor g00989(.dina(n1200), .dinb(n1050), .dout(n1201));
  jnot g00990(.din(n1201), .dout(n1202));
  jand g00991(.dina(n1202), .dinb(n1198), .dout(n1203));
  jor  g00992(.dina(n1203), .dinb(n1197), .dout(n1204));
  jand g00993(.dina(n1204), .dinb(asqrt[54] ), .dout(n1205));
  jnot g00994(.din(n1056), .dout(n1206));
  jand g00995(.dina(n1206), .dinb(n1054), .dout(n1207));
  jand g00996(.dina(n1207), .dinb(asqrt[50] ), .dout(n1208));
  jxor g00997(.dina(n1208), .dinb(n1064), .dout(n1209));
  jnot g00998(.din(n1209), .dout(n1210));
  jor  g00999(.dina(n1197), .dinb(asqrt[54] ), .dout(n1211));
  jor  g01000(.dina(n1211), .dinb(n1203), .dout(n1212));
  jand g01001(.dina(n1212), .dinb(n1210), .dout(n1213));
  jor  g01002(.dina(n1213), .dinb(n1205), .dout(n1214));
  jand g01003(.dina(n1214), .dinb(asqrt[55] ), .dout(n1215));
  jor  g01004(.dina(n1214), .dinb(asqrt[55] ), .dout(n1216));
  jnot g01005(.din(n1071), .dout(n1217));
  jxor g01006(.dina(n1066), .dinb(n791), .dout(n1218));
  jand g01007(.dina(n1218), .dinb(asqrt[50] ), .dout(n1219));
  jxor g01008(.dina(n1219), .dinb(n1217), .dout(n1220));
  jand g01009(.dina(n1220), .dinb(n1216), .dout(n1221));
  jor  g01010(.dina(n1221), .dinb(n1215), .dout(n1222));
  jand g01011(.dina(n1222), .dinb(asqrt[56] ), .dout(n1223));
  jor  g01012(.dina(n1215), .dinb(asqrt[56] ), .dout(n1224));
  jor  g01013(.dina(n1224), .dinb(n1221), .dout(n1225));
  jnot g01014(.din(n1078), .dout(n1226));
  jnot g01015(.din(n1080), .dout(n1227));
  jand g01016(.dina(asqrt[50] ), .dinb(n1074), .dout(n1228));
  jand g01017(.dina(n1228), .dinb(n1227), .dout(n1229));
  jor  g01018(.dina(n1229), .dinb(n1226), .dout(n1230));
  jnot g01019(.din(n1081), .dout(n1231));
  jand g01020(.dina(n1228), .dinb(n1231), .dout(n1232));
  jnot g01021(.din(n1232), .dout(n1233));
  jand g01022(.dina(n1233), .dinb(n1230), .dout(n1234));
  jand g01023(.dina(n1234), .dinb(n1225), .dout(n1235));
  jor  g01024(.dina(n1235), .dinb(n1223), .dout(n1236));
  jand g01025(.dina(n1236), .dinb(asqrt[57] ), .dout(n1237));
  jor  g01026(.dina(n1236), .dinb(asqrt[57] ), .dout(n1238));
  jxor g01027(.dina(n1082), .dinb(n590), .dout(n1239));
  jand g01028(.dina(n1239), .dinb(asqrt[50] ), .dout(n1240));
  jxor g01029(.dina(n1240), .dinb(n1087), .dout(n1241));
  jand g01030(.dina(n1241), .dinb(n1238), .dout(n1242));
  jor  g01031(.dina(n1242), .dinb(n1237), .dout(n1243));
  jand g01032(.dina(n1243), .dinb(asqrt[58] ), .dout(n1244));
  jnot g01033(.din(n1093), .dout(n1245));
  jand g01034(.dina(n1245), .dinb(n1091), .dout(n1246));
  jand g01035(.dina(n1246), .dinb(asqrt[50] ), .dout(n1247));
  jxor g01036(.dina(n1247), .dinb(n1101), .dout(n1248));
  jnot g01037(.din(n1248), .dout(n1249));
  jor  g01038(.dina(n1237), .dinb(asqrt[58] ), .dout(n1250));
  jor  g01039(.dina(n1250), .dinb(n1242), .dout(n1251));
  jand g01040(.dina(n1251), .dinb(n1249), .dout(n1252));
  jor  g01041(.dina(n1252), .dinb(n1244), .dout(n1253));
  jand g01042(.dina(n1253), .dinb(asqrt[59] ), .dout(n1254));
  jor  g01043(.dina(n1253), .dinb(asqrt[59] ), .dout(n1255));
  jxor g01044(.dina(n1103), .dinb(n425), .dout(n1256));
  jand g01045(.dina(n1256), .dinb(asqrt[50] ), .dout(n1257));
  jxor g01046(.dina(n1257), .dinb(n1109), .dout(n1258));
  jand g01047(.dina(n1258), .dinb(n1255), .dout(n1259));
  jor  g01048(.dina(n1259), .dinb(n1254), .dout(n1260));
  jand g01049(.dina(n1260), .dinb(asqrt[60] ), .dout(n1261));
  jor  g01050(.dina(n1254), .dinb(asqrt[60] ), .dout(n1262));
  jor  g01051(.dina(n1262), .dinb(n1259), .dout(n1263));
  jnot g01052(.din(n1117), .dout(n1264));
  jnot g01053(.din(n1119), .dout(n1265));
  jand g01054(.dina(asqrt[50] ), .dinb(n1113), .dout(n1266));
  jand g01055(.dina(n1266), .dinb(n1265), .dout(n1267));
  jor  g01056(.dina(n1267), .dinb(n1264), .dout(n1268));
  jnot g01057(.din(n1120), .dout(n1269));
  jand g01058(.dina(n1266), .dinb(n1269), .dout(n1270));
  jnot g01059(.din(n1270), .dout(n1271));
  jand g01060(.dina(n1271), .dinb(n1268), .dout(n1272));
  jand g01061(.dina(n1272), .dinb(n1263), .dout(n1273));
  jor  g01062(.dina(n1273), .dinb(n1261), .dout(n1274));
  jand g01063(.dina(n1274), .dinb(asqrt[61] ), .dout(n1275));
  jxor g01064(.dina(n1121), .dinb(n290), .dout(n1276));
  jand g01065(.dina(n1276), .dinb(asqrt[50] ), .dout(n1277));
  jxor g01066(.dina(n1277), .dinb(n1128), .dout(n1278));
  jnot g01067(.din(n1278), .dout(n1279));
  jor  g01068(.dina(n1274), .dinb(asqrt[61] ), .dout(n1280));
  jand g01069(.dina(n1280), .dinb(n1279), .dout(n1281));
  jor  g01070(.dina(n1281), .dinb(n1275), .dout(n1282));
  jand g01071(.dina(n1282), .dinb(asqrt[62] ), .dout(n1283));
  jnot g01072(.din(n1133), .dout(n1284));
  jand g01073(.dina(n1284), .dinb(n1131), .dout(n1285));
  jand g01074(.dina(n1285), .dinb(asqrt[50] ), .dout(n1286));
  jxor g01075(.dina(n1286), .dinb(n1141), .dout(n1287));
  jnot g01076(.din(n1287), .dout(n1288));
  jor  g01077(.dina(n1275), .dinb(asqrt[62] ), .dout(n1289));
  jor  g01078(.dina(n1289), .dinb(n1281), .dout(n1290));
  jand g01079(.dina(n1290), .dinb(n1288), .dout(n1291));
  jor  g01080(.dina(n1291), .dinb(n1283), .dout(n1292));
  jxor g01081(.dina(n1143), .dinb(n199), .dout(n1293));
  jand g01082(.dina(n1293), .dinb(asqrt[50] ), .dout(n1294));
  jxor g01083(.dina(n1294), .dinb(n1148), .dout(n1295));
  jnot g01084(.din(n1150), .dout(n1296));
  jnot g01085(.din(n1154), .dout(n1297));
  jand g01086(.dina(asqrt[50] ), .dinb(n1297), .dout(n1298));
  jand g01087(.dina(n1298), .dinb(n1296), .dout(n1299));
  jor  g01088(.dina(n1299), .dinb(n1161), .dout(n1300));
  jor  g01089(.dina(n1300), .dinb(n1295), .dout(n1301));
  jnot g01090(.din(n1301), .dout(n1302));
  jand g01091(.dina(n1302), .dinb(n1292), .dout(n1303));
  jor  g01092(.dina(n1303), .dinb(asqrt[63] ), .dout(n1304));
  jnot g01093(.din(n1295), .dout(n1305));
  jor  g01094(.dina(n1305), .dinb(n1292), .dout(n1306));
  jor  g01095(.dina(n1298), .dinb(n1296), .dout(n1307));
  jand g01096(.dina(n1297), .dinb(n1296), .dout(n1308));
  jor  g01097(.dina(n1308), .dinb(n194), .dout(n1309));
  jnot g01098(.din(n1309), .dout(n1310));
  jand g01099(.dina(n1310), .dinb(n1307), .dout(n1311));
  jnot g01100(.din(asqrt[50] ), .dout(n1312));
  jnot g01101(.din(n1311), .dout(n1315));
  jand g01102(.dina(n1315), .dinb(n1306), .dout(n1316));
  jand g01103(.dina(n1316), .dinb(n1304), .dout(n1317));
  jnot g01104(.din(n1317), .dout(asqrt[49] ));
  jor  g01105(.dina(n1317), .dinb(n1172), .dout(n1319));
  jnot g01106(.din(a[96] ), .dout(n1320));
  jnot g01107(.din(a[97] ), .dout(n1321));
  jand g01108(.dina(n1172), .dinb(n1321), .dout(n1322));
  jand g01109(.dina(n1322), .dinb(n1320), .dout(n1323));
  jnot g01110(.din(n1323), .dout(n1324));
  jand g01111(.dina(n1324), .dinb(n1319), .dout(n1325));
  jor  g01112(.dina(n1325), .dinb(n1312), .dout(n1326));
  jor  g01113(.dina(n1317), .dinb(a[98] ), .dout(n1327));
  jxor g01114(.dina(n1327), .dinb(n1173), .dout(n1328));
  jand g01115(.dina(n1325), .dinb(n1312), .dout(n1329));
  jor  g01116(.dina(n1329), .dinb(n1328), .dout(n1330));
  jand g01117(.dina(n1330), .dinb(n1326), .dout(n1331));
  jor  g01118(.dina(n1331), .dinb(n1039), .dout(n1332));
  jand g01119(.dina(n1326), .dinb(n1039), .dout(n1333));
  jand g01120(.dina(n1333), .dinb(n1330), .dout(n1334));
  jor  g01121(.dina(n1327), .dinb(a[99] ), .dout(n1335));
  jnot g01122(.din(n1304), .dout(n1336));
  jnot g01123(.din(n1306), .dout(n1337));
  jor  g01124(.dina(n1311), .dinb(n1312), .dout(n1338));
  jor  g01125(.dina(n1338), .dinb(n1337), .dout(n1339));
  jor  g01126(.dina(n1339), .dinb(n1336), .dout(n1340));
  jand g01127(.dina(n1340), .dinb(n1335), .dout(n1341));
  jxor g01128(.dina(n1341), .dinb(n1042), .dout(n1342));
  jor  g01129(.dina(n1342), .dinb(n1334), .dout(n1343));
  jand g01130(.dina(n1343), .dinb(n1332), .dout(n1344));
  jor  g01131(.dina(n1344), .dinb(n1034), .dout(n1345));
  jand g01132(.dina(n1344), .dinb(n1034), .dout(n1346));
  jxor g01133(.dina(n1176), .dinb(n1039), .dout(n1347));
  jor  g01134(.dina(n1347), .dinb(n1317), .dout(n1348));
  jxor g01135(.dina(n1348), .dinb(n1179), .dout(n1349));
  jor  g01136(.dina(n1349), .dinb(n1346), .dout(n1350));
  jand g01137(.dina(n1350), .dinb(n1345), .dout(n1351));
  jor  g01138(.dina(n1351), .dinb(n796), .dout(n1352));
  jnot g01139(.din(n1185), .dout(n1353));
  jor  g01140(.dina(n1353), .dinb(n1183), .dout(n1354));
  jor  g01141(.dina(n1354), .dinb(n1317), .dout(n1355));
  jxor g01142(.dina(n1355), .dinb(n1194), .dout(n1356));
  jand g01143(.dina(n1345), .dinb(n796), .dout(n1357));
  jand g01144(.dina(n1357), .dinb(n1350), .dout(n1358));
  jor  g01145(.dina(n1358), .dinb(n1356), .dout(n1359));
  jand g01146(.dina(n1359), .dinb(n1352), .dout(n1360));
  jor  g01147(.dina(n1360), .dinb(n791), .dout(n1361));
  jand g01148(.dina(n1360), .dinb(n791), .dout(n1362));
  jxor g01149(.dina(n1196), .dinb(n796), .dout(n1363));
  jor  g01150(.dina(n1363), .dinb(n1317), .dout(n1364));
  jxor g01151(.dina(n1364), .dinb(n1201), .dout(n1365));
  jnot g01152(.din(n1365), .dout(n1366));
  jor  g01153(.dina(n1366), .dinb(n1362), .dout(n1367));
  jand g01154(.dina(n1367), .dinb(n1361), .dout(n1368));
  jor  g01155(.dina(n1368), .dinb(n595), .dout(n1369));
  jand g01156(.dina(n1361), .dinb(n595), .dout(n1370));
  jand g01157(.dina(n1370), .dinb(n1367), .dout(n1371));
  jnot g01158(.din(n1205), .dout(n1372));
  jand g01159(.dina(asqrt[49] ), .dinb(n1372), .dout(n1373));
  jand g01160(.dina(n1373), .dinb(n1212), .dout(n1374));
  jor  g01161(.dina(n1374), .dinb(n1210), .dout(n1375));
  jand g01162(.dina(n1373), .dinb(n1213), .dout(n1376));
  jnot g01163(.din(n1376), .dout(n1377));
  jand g01164(.dina(n1377), .dinb(n1375), .dout(n1378));
  jnot g01165(.din(n1378), .dout(n1379));
  jor  g01166(.dina(n1379), .dinb(n1371), .dout(n1380));
  jand g01167(.dina(n1380), .dinb(n1369), .dout(n1381));
  jor  g01168(.dina(n1381), .dinb(n590), .dout(n1382));
  jand g01169(.dina(n1381), .dinb(n590), .dout(n1383));
  jnot g01170(.din(n1220), .dout(n1384));
  jxor g01171(.dina(n1214), .dinb(n595), .dout(n1385));
  jor  g01172(.dina(n1385), .dinb(n1317), .dout(n1386));
  jxor g01173(.dina(n1386), .dinb(n1384), .dout(n1387));
  jnot g01174(.din(n1387), .dout(n1388));
  jor  g01175(.dina(n1388), .dinb(n1383), .dout(n1389));
  jand g01176(.dina(n1389), .dinb(n1382), .dout(n1390));
  jor  g01177(.dina(n1390), .dinb(n430), .dout(n1391));
  jnot g01178(.din(n1225), .dout(n1392));
  jor  g01179(.dina(n1392), .dinb(n1223), .dout(n1393));
  jor  g01180(.dina(n1393), .dinb(n1317), .dout(n1394));
  jxor g01181(.dina(n1394), .dinb(n1234), .dout(n1395));
  jand g01182(.dina(n1382), .dinb(n430), .dout(n1396));
  jand g01183(.dina(n1396), .dinb(n1389), .dout(n1397));
  jor  g01184(.dina(n1397), .dinb(n1395), .dout(n1398));
  jand g01185(.dina(n1398), .dinb(n1391), .dout(n1399));
  jor  g01186(.dina(n1399), .dinb(n425), .dout(n1400));
  jand g01187(.dina(n1399), .dinb(n425), .dout(n1401));
  jnot g01188(.din(n1241), .dout(n1402));
  jxor g01189(.dina(n1236), .dinb(n430), .dout(n1403));
  jor  g01190(.dina(n1403), .dinb(n1317), .dout(n1404));
  jxor g01191(.dina(n1404), .dinb(n1402), .dout(n1405));
  jnot g01192(.din(n1405), .dout(n1406));
  jor  g01193(.dina(n1406), .dinb(n1401), .dout(n1407));
  jand g01194(.dina(n1407), .dinb(n1400), .dout(n1408));
  jor  g01195(.dina(n1408), .dinb(n305), .dout(n1409));
  jand g01196(.dina(n1400), .dinb(n305), .dout(n1410));
  jand g01197(.dina(n1410), .dinb(n1407), .dout(n1411));
  jnot g01198(.din(n1244), .dout(n1412));
  jand g01199(.dina(asqrt[49] ), .dinb(n1412), .dout(n1413));
  jand g01200(.dina(n1413), .dinb(n1251), .dout(n1414));
  jor  g01201(.dina(n1414), .dinb(n1249), .dout(n1415));
  jand g01202(.dina(n1413), .dinb(n1252), .dout(n1416));
  jnot g01203(.din(n1416), .dout(n1417));
  jand g01204(.dina(n1417), .dinb(n1415), .dout(n1418));
  jnot g01205(.din(n1418), .dout(n1419));
  jor  g01206(.dina(n1419), .dinb(n1411), .dout(n1420));
  jand g01207(.dina(n1420), .dinb(n1409), .dout(n1421));
  jor  g01208(.dina(n1421), .dinb(n290), .dout(n1422));
  jxor g01209(.dina(n1253), .dinb(n305), .dout(n1423));
  jor  g01210(.dina(n1423), .dinb(n1317), .dout(n1424));
  jxor g01211(.dina(n1424), .dinb(n1258), .dout(n1425));
  jand g01212(.dina(n1421), .dinb(n290), .dout(n1426));
  jor  g01213(.dina(n1426), .dinb(n1425), .dout(n1427));
  jand g01214(.dina(n1427), .dinb(n1422), .dout(n1428));
  jor  g01215(.dina(n1428), .dinb(n223), .dout(n1429));
  jnot g01216(.din(n1263), .dout(n1430));
  jor  g01217(.dina(n1430), .dinb(n1261), .dout(n1431));
  jor  g01218(.dina(n1431), .dinb(n1317), .dout(n1432));
  jxor g01219(.dina(n1432), .dinb(n1272), .dout(n1433));
  jand g01220(.dina(n1422), .dinb(n223), .dout(n1434));
  jand g01221(.dina(n1434), .dinb(n1427), .dout(n1435));
  jor  g01222(.dina(n1435), .dinb(n1433), .dout(n1436));
  jand g01223(.dina(n1436), .dinb(n1429), .dout(n1437));
  jor  g01224(.dina(n1437), .dinb(n199), .dout(n1438));
  jand g01225(.dina(n1437), .dinb(n199), .dout(n1439));
  jnot g01226(.din(n1275), .dout(n1440));
  jand g01227(.dina(asqrt[49] ), .dinb(n1440), .dout(n1441));
  jand g01228(.dina(n1441), .dinb(n1280), .dout(n1442));
  jor  g01229(.dina(n1442), .dinb(n1279), .dout(n1443));
  jand g01230(.dina(n1441), .dinb(n1281), .dout(n1444));
  jnot g01231(.din(n1444), .dout(n1445));
  jand g01232(.dina(n1445), .dinb(n1443), .dout(n1446));
  jnot g01233(.din(n1446), .dout(n1447));
  jor  g01234(.dina(n1447), .dinb(n1439), .dout(n1448));
  jand g01235(.dina(n1448), .dinb(n1438), .dout(n1449));
  jnot g01236(.din(n1283), .dout(n1450));
  jand g01237(.dina(asqrt[49] ), .dinb(n1450), .dout(n1451));
  jand g01238(.dina(n1451), .dinb(n1290), .dout(n1452));
  jor  g01239(.dina(n1452), .dinb(n1288), .dout(n1453));
  jand g01240(.dina(n1451), .dinb(n1291), .dout(n1454));
  jnot g01241(.din(n1454), .dout(n1455));
  jand g01242(.dina(n1455), .dinb(n1453), .dout(n1456));
  jnot g01243(.din(n1456), .dout(n1457));
  jand g01244(.dina(asqrt[49] ), .dinb(n1305), .dout(n1458));
  jand g01245(.dina(n1458), .dinb(n1292), .dout(n1459));
  jor  g01246(.dina(n1459), .dinb(n1337), .dout(n1460));
  jor  g01247(.dina(n1460), .dinb(n1457), .dout(n1461));
  jor  g01248(.dina(n1461), .dinb(n1449), .dout(n1462));
  jand g01249(.dina(n1462), .dinb(n194), .dout(n1463));
  jand g01250(.dina(n1457), .dinb(n1449), .dout(n1464));
  jor  g01251(.dina(n1458), .dinb(n1292), .dout(n1465));
  jand g01252(.dina(n1305), .dinb(n1292), .dout(n1466));
  jor  g01253(.dina(n1466), .dinb(n194), .dout(n1467));
  jnot g01254(.din(n1467), .dout(n1468));
  jand g01255(.dina(n1468), .dinb(n1465), .dout(n1469));
  jor  g01256(.dina(n1469), .dinb(n1464), .dout(n1472));
  jor  g01257(.dina(n1472), .dinb(n1463), .dout(asqrt[48] ));
  jand g01258(.dina(asqrt[48] ), .dinb(a[96] ), .dout(n1474));
  jnot g01259(.din(a[94] ), .dout(n1475));
  jnot g01260(.din(a[95] ), .dout(n1476));
  jand g01261(.dina(n1320), .dinb(n1476), .dout(n1477));
  jand g01262(.dina(n1477), .dinb(n1475), .dout(n1478));
  jor  g01263(.dina(n1478), .dinb(n1474), .dout(n1479));
  jand g01264(.dina(n1479), .dinb(asqrt[49] ), .dout(n1480));
  jand g01265(.dina(asqrt[48] ), .dinb(n1320), .dout(n1481));
  jxor g01266(.dina(n1481), .dinb(n1321), .dout(n1482));
  jor  g01267(.dina(n1479), .dinb(asqrt[49] ), .dout(n1483));
  jand g01268(.dina(n1483), .dinb(n1482), .dout(n1484));
  jor  g01269(.dina(n1484), .dinb(n1480), .dout(n1485));
  jand g01270(.dina(n1485), .dinb(asqrt[50] ), .dout(n1486));
  jor  g01271(.dina(n1480), .dinb(asqrt[50] ), .dout(n1487));
  jor  g01272(.dina(n1487), .dinb(n1484), .dout(n1488));
  jand g01273(.dina(n1481), .dinb(n1321), .dout(n1489));
  jnot g01274(.din(n1463), .dout(n1490));
  jnot g01275(.din(n1464), .dout(n1491));
  jnot g01276(.din(n1469), .dout(n1492));
  jand g01277(.dina(n1492), .dinb(asqrt[49] ), .dout(n1493));
  jand g01278(.dina(n1493), .dinb(n1491), .dout(n1494));
  jand g01279(.dina(n1494), .dinb(n1490), .dout(n1495));
  jor  g01280(.dina(n1495), .dinb(n1489), .dout(n1496));
  jxor g01281(.dina(n1496), .dinb(n1172), .dout(n1497));
  jand g01282(.dina(n1497), .dinb(n1488), .dout(n1498));
  jor  g01283(.dina(n1498), .dinb(n1486), .dout(n1499));
  jand g01284(.dina(n1499), .dinb(asqrt[51] ), .dout(n1500));
  jor  g01285(.dina(n1499), .dinb(asqrt[51] ), .dout(n1501));
  jxor g01286(.dina(n1325), .dinb(n1312), .dout(n1502));
  jand g01287(.dina(n1502), .dinb(asqrt[48] ), .dout(n1503));
  jxor g01288(.dina(n1503), .dinb(n1328), .dout(n1504));
  jnot g01289(.din(n1504), .dout(n1505));
  jand g01290(.dina(n1505), .dinb(n1501), .dout(n1506));
  jor  g01291(.dina(n1506), .dinb(n1500), .dout(n1507));
  jand g01292(.dina(n1507), .dinb(asqrt[52] ), .dout(n1508));
  jnot g01293(.din(n1334), .dout(n1509));
  jand g01294(.dina(n1509), .dinb(n1332), .dout(n1510));
  jand g01295(.dina(n1510), .dinb(asqrt[48] ), .dout(n1511));
  jxor g01296(.dina(n1511), .dinb(n1342), .dout(n1512));
  jnot g01297(.din(n1512), .dout(n1513));
  jor  g01298(.dina(n1500), .dinb(asqrt[52] ), .dout(n1514));
  jor  g01299(.dina(n1514), .dinb(n1506), .dout(n1515));
  jand g01300(.dina(n1515), .dinb(n1513), .dout(n1516));
  jor  g01301(.dina(n1516), .dinb(n1508), .dout(n1517));
  jand g01302(.dina(n1517), .dinb(asqrt[53] ), .dout(n1518));
  jor  g01303(.dina(n1517), .dinb(asqrt[53] ), .dout(n1519));
  jnot g01304(.din(n1349), .dout(n1520));
  jxor g01305(.dina(n1344), .dinb(n1034), .dout(n1521));
  jand g01306(.dina(n1521), .dinb(asqrt[48] ), .dout(n1522));
  jxor g01307(.dina(n1522), .dinb(n1520), .dout(n1523));
  jand g01308(.dina(n1523), .dinb(n1519), .dout(n1524));
  jor  g01309(.dina(n1524), .dinb(n1518), .dout(n1525));
  jand g01310(.dina(n1525), .dinb(asqrt[54] ), .dout(n1526));
  jor  g01311(.dina(n1518), .dinb(asqrt[54] ), .dout(n1527));
  jor  g01312(.dina(n1527), .dinb(n1524), .dout(n1528));
  jnot g01313(.din(n1356), .dout(n1529));
  jnot g01314(.din(n1358), .dout(n1530));
  jand g01315(.dina(asqrt[48] ), .dinb(n1352), .dout(n1531));
  jand g01316(.dina(n1531), .dinb(n1530), .dout(n1532));
  jor  g01317(.dina(n1532), .dinb(n1529), .dout(n1533));
  jnot g01318(.din(n1359), .dout(n1534));
  jand g01319(.dina(n1531), .dinb(n1534), .dout(n1535));
  jnot g01320(.din(n1535), .dout(n1536));
  jand g01321(.dina(n1536), .dinb(n1533), .dout(n1537));
  jand g01322(.dina(n1537), .dinb(n1528), .dout(n1538));
  jor  g01323(.dina(n1538), .dinb(n1526), .dout(n1539));
  jand g01324(.dina(n1539), .dinb(asqrt[55] ), .dout(n1540));
  jor  g01325(.dina(n1539), .dinb(asqrt[55] ), .dout(n1541));
  jxor g01326(.dina(n1360), .dinb(n791), .dout(n1542));
  jand g01327(.dina(n1542), .dinb(asqrt[48] ), .dout(n1543));
  jxor g01328(.dina(n1543), .dinb(n1365), .dout(n1544));
  jand g01329(.dina(n1544), .dinb(n1541), .dout(n1545));
  jor  g01330(.dina(n1545), .dinb(n1540), .dout(n1546));
  jand g01331(.dina(n1546), .dinb(asqrt[56] ), .dout(n1547));
  jnot g01332(.din(n1371), .dout(n1548));
  jand g01333(.dina(n1548), .dinb(n1369), .dout(n1549));
  jand g01334(.dina(n1549), .dinb(asqrt[48] ), .dout(n1550));
  jxor g01335(.dina(n1550), .dinb(n1379), .dout(n1551));
  jnot g01336(.din(n1551), .dout(n1552));
  jor  g01337(.dina(n1540), .dinb(asqrt[56] ), .dout(n1553));
  jor  g01338(.dina(n1553), .dinb(n1545), .dout(n1554));
  jand g01339(.dina(n1554), .dinb(n1552), .dout(n1555));
  jor  g01340(.dina(n1555), .dinb(n1547), .dout(n1556));
  jand g01341(.dina(n1556), .dinb(asqrt[57] ), .dout(n1557));
  jor  g01342(.dina(n1556), .dinb(asqrt[57] ), .dout(n1558));
  jxor g01343(.dina(n1381), .dinb(n590), .dout(n1559));
  jand g01344(.dina(n1559), .dinb(asqrt[48] ), .dout(n1560));
  jxor g01345(.dina(n1560), .dinb(n1387), .dout(n1561));
  jand g01346(.dina(n1561), .dinb(n1558), .dout(n1562));
  jor  g01347(.dina(n1562), .dinb(n1557), .dout(n1563));
  jand g01348(.dina(n1563), .dinb(asqrt[58] ), .dout(n1564));
  jor  g01349(.dina(n1557), .dinb(asqrt[58] ), .dout(n1565));
  jor  g01350(.dina(n1565), .dinb(n1562), .dout(n1566));
  jnot g01351(.din(n1395), .dout(n1567));
  jnot g01352(.din(n1397), .dout(n1568));
  jand g01353(.dina(asqrt[48] ), .dinb(n1391), .dout(n1569));
  jand g01354(.dina(n1569), .dinb(n1568), .dout(n1570));
  jor  g01355(.dina(n1570), .dinb(n1567), .dout(n1571));
  jnot g01356(.din(n1398), .dout(n1572));
  jand g01357(.dina(n1569), .dinb(n1572), .dout(n1573));
  jnot g01358(.din(n1573), .dout(n1574));
  jand g01359(.dina(n1574), .dinb(n1571), .dout(n1575));
  jand g01360(.dina(n1575), .dinb(n1566), .dout(n1576));
  jor  g01361(.dina(n1576), .dinb(n1564), .dout(n1577));
  jand g01362(.dina(n1577), .dinb(asqrt[59] ), .dout(n1578));
  jxor g01363(.dina(n1399), .dinb(n425), .dout(n1579));
  jand g01364(.dina(n1579), .dinb(asqrt[48] ), .dout(n1580));
  jxor g01365(.dina(n1580), .dinb(n1406), .dout(n1581));
  jnot g01366(.din(n1581), .dout(n1582));
  jor  g01367(.dina(n1577), .dinb(asqrt[59] ), .dout(n1583));
  jand g01368(.dina(n1583), .dinb(n1582), .dout(n1584));
  jor  g01369(.dina(n1584), .dinb(n1578), .dout(n1585));
  jand g01370(.dina(n1585), .dinb(asqrt[60] ), .dout(n1586));
  jnot g01371(.din(n1411), .dout(n1587));
  jand g01372(.dina(n1587), .dinb(n1409), .dout(n1588));
  jand g01373(.dina(n1588), .dinb(asqrt[48] ), .dout(n1589));
  jxor g01374(.dina(n1589), .dinb(n1419), .dout(n1590));
  jnot g01375(.din(n1590), .dout(n1591));
  jor  g01376(.dina(n1578), .dinb(asqrt[60] ), .dout(n1592));
  jor  g01377(.dina(n1592), .dinb(n1584), .dout(n1593));
  jand g01378(.dina(n1593), .dinb(n1591), .dout(n1594));
  jor  g01379(.dina(n1594), .dinb(n1586), .dout(n1595));
  jand g01380(.dina(n1595), .dinb(asqrt[61] ), .dout(n1596));
  jor  g01381(.dina(n1595), .dinb(asqrt[61] ), .dout(n1597));
  jnot g01382(.din(n1425), .dout(n1598));
  jnot g01383(.din(n1426), .dout(n1599));
  jand g01384(.dina(asqrt[48] ), .dinb(n1422), .dout(n1600));
  jand g01385(.dina(n1600), .dinb(n1599), .dout(n1601));
  jor  g01386(.dina(n1601), .dinb(n1598), .dout(n1602));
  jnot g01387(.din(n1427), .dout(n1603));
  jand g01388(.dina(n1600), .dinb(n1603), .dout(n1604));
  jnot g01389(.din(n1604), .dout(n1605));
  jand g01390(.dina(n1605), .dinb(n1602), .dout(n1606));
  jand g01391(.dina(n1606), .dinb(n1597), .dout(n1607));
  jor  g01392(.dina(n1607), .dinb(n1596), .dout(n1608));
  jand g01393(.dina(n1608), .dinb(asqrt[62] ), .dout(n1609));
  jor  g01394(.dina(n1596), .dinb(asqrt[62] ), .dout(n1610));
  jor  g01395(.dina(n1610), .dinb(n1607), .dout(n1611));
  jnot g01396(.din(n1433), .dout(n1612));
  jnot g01397(.din(n1435), .dout(n1613));
  jand g01398(.dina(asqrt[48] ), .dinb(n1429), .dout(n1614));
  jand g01399(.dina(n1614), .dinb(n1613), .dout(n1615));
  jor  g01400(.dina(n1615), .dinb(n1612), .dout(n1616));
  jnot g01401(.din(n1436), .dout(n1617));
  jand g01402(.dina(n1614), .dinb(n1617), .dout(n1618));
  jnot g01403(.din(n1618), .dout(n1619));
  jand g01404(.dina(n1619), .dinb(n1616), .dout(n1620));
  jand g01405(.dina(n1620), .dinb(n1611), .dout(n1621));
  jor  g01406(.dina(n1621), .dinb(n1609), .dout(n1622));
  jxor g01407(.dina(n1437), .dinb(n199), .dout(n1623));
  jand g01408(.dina(n1623), .dinb(asqrt[48] ), .dout(n1624));
  jxor g01409(.dina(n1624), .dinb(n1447), .dout(n1625));
  jnot g01410(.din(n1449), .dout(n1626));
  jand g01411(.dina(asqrt[48] ), .dinb(n1456), .dout(n1627));
  jand g01412(.dina(n1627), .dinb(n1626), .dout(n1628));
  jor  g01413(.dina(n1628), .dinb(n1464), .dout(n1629));
  jor  g01414(.dina(n1629), .dinb(n1625), .dout(n1630));
  jnot g01415(.din(n1630), .dout(n1631));
  jand g01416(.dina(n1631), .dinb(n1622), .dout(n1632));
  jor  g01417(.dina(n1632), .dinb(asqrt[63] ), .dout(n1633));
  jnot g01418(.din(n1625), .dout(n1634));
  jor  g01419(.dina(n1634), .dinb(n1622), .dout(n1635));
  jor  g01420(.dina(n1627), .dinb(n1626), .dout(n1636));
  jand g01421(.dina(n1456), .dinb(n1626), .dout(n1637));
  jor  g01422(.dina(n1637), .dinb(n194), .dout(n1638));
  jnot g01423(.din(n1638), .dout(n1639));
  jand g01424(.dina(n1639), .dinb(n1636), .dout(n1640));
  jnot g01425(.din(asqrt[48] ), .dout(n1641));
  jnot g01426(.din(n1640), .dout(n1644));
  jand g01427(.dina(n1644), .dinb(n1635), .dout(n1645));
  jand g01428(.dina(n1645), .dinb(n1633), .dout(n1646));
  jnot g01429(.din(n1646), .dout(asqrt[47] ));
  jor  g01430(.dina(n1646), .dinb(n1475), .dout(n1648));
  jnot g01431(.din(a[92] ), .dout(n1649));
  jnot g01432(.din(a[93] ), .dout(n1650));
  jand g01433(.dina(n1475), .dinb(n1650), .dout(n1651));
  jand g01434(.dina(n1651), .dinb(n1649), .dout(n1652));
  jnot g01435(.din(n1652), .dout(n1653));
  jand g01436(.dina(n1653), .dinb(n1648), .dout(n1654));
  jor  g01437(.dina(n1654), .dinb(n1641), .dout(n1655));
  jor  g01438(.dina(n1646), .dinb(a[94] ), .dout(n1656));
  jxor g01439(.dina(n1656), .dinb(n1476), .dout(n1657));
  jand g01440(.dina(n1654), .dinb(n1641), .dout(n1658));
  jor  g01441(.dina(n1658), .dinb(n1657), .dout(n1659));
  jand g01442(.dina(n1659), .dinb(n1655), .dout(n1660));
  jor  g01443(.dina(n1660), .dinb(n1317), .dout(n1661));
  jand g01444(.dina(n1655), .dinb(n1317), .dout(n1662));
  jand g01445(.dina(n1662), .dinb(n1659), .dout(n1663));
  jor  g01446(.dina(n1656), .dinb(a[95] ), .dout(n1664));
  jnot g01447(.din(n1633), .dout(n1665));
  jnot g01448(.din(n1635), .dout(n1666));
  jor  g01449(.dina(n1640), .dinb(n1641), .dout(n1667));
  jor  g01450(.dina(n1667), .dinb(n1666), .dout(n1668));
  jor  g01451(.dina(n1668), .dinb(n1665), .dout(n1669));
  jand g01452(.dina(n1669), .dinb(n1664), .dout(n1670));
  jxor g01453(.dina(n1670), .dinb(n1320), .dout(n1671));
  jor  g01454(.dina(n1671), .dinb(n1663), .dout(n1672));
  jand g01455(.dina(n1672), .dinb(n1661), .dout(n1673));
  jor  g01456(.dina(n1673), .dinb(n1312), .dout(n1674));
  jand g01457(.dina(n1673), .dinb(n1312), .dout(n1675));
  jxor g01458(.dina(n1479), .dinb(n1317), .dout(n1676));
  jor  g01459(.dina(n1676), .dinb(n1646), .dout(n1677));
  jxor g01460(.dina(n1677), .dinb(n1482), .dout(n1678));
  jor  g01461(.dina(n1678), .dinb(n1675), .dout(n1679));
  jand g01462(.dina(n1679), .dinb(n1674), .dout(n1680));
  jor  g01463(.dina(n1680), .dinb(n1039), .dout(n1681));
  jnot g01464(.din(n1488), .dout(n1682));
  jor  g01465(.dina(n1682), .dinb(n1486), .dout(n1683));
  jor  g01466(.dina(n1683), .dinb(n1646), .dout(n1684));
  jxor g01467(.dina(n1684), .dinb(n1497), .dout(n1685));
  jand g01468(.dina(n1674), .dinb(n1039), .dout(n1686));
  jand g01469(.dina(n1686), .dinb(n1679), .dout(n1687));
  jor  g01470(.dina(n1687), .dinb(n1685), .dout(n1688));
  jand g01471(.dina(n1688), .dinb(n1681), .dout(n1689));
  jor  g01472(.dina(n1689), .dinb(n1034), .dout(n1690));
  jand g01473(.dina(n1689), .dinb(n1034), .dout(n1691));
  jxor g01474(.dina(n1499), .dinb(n1039), .dout(n1692));
  jor  g01475(.dina(n1692), .dinb(n1646), .dout(n1693));
  jxor g01476(.dina(n1693), .dinb(n1504), .dout(n1694));
  jnot g01477(.din(n1694), .dout(n1695));
  jor  g01478(.dina(n1695), .dinb(n1691), .dout(n1696));
  jand g01479(.dina(n1696), .dinb(n1690), .dout(n1697));
  jor  g01480(.dina(n1697), .dinb(n796), .dout(n1698));
  jand g01481(.dina(n1690), .dinb(n796), .dout(n1699));
  jand g01482(.dina(n1699), .dinb(n1696), .dout(n1700));
  jnot g01483(.din(n1508), .dout(n1701));
  jand g01484(.dina(asqrt[47] ), .dinb(n1701), .dout(n1702));
  jand g01485(.dina(n1702), .dinb(n1515), .dout(n1703));
  jor  g01486(.dina(n1703), .dinb(n1513), .dout(n1704));
  jand g01487(.dina(n1702), .dinb(n1516), .dout(n1705));
  jnot g01488(.din(n1705), .dout(n1706));
  jand g01489(.dina(n1706), .dinb(n1704), .dout(n1707));
  jnot g01490(.din(n1707), .dout(n1708));
  jor  g01491(.dina(n1708), .dinb(n1700), .dout(n1709));
  jand g01492(.dina(n1709), .dinb(n1698), .dout(n1710));
  jor  g01493(.dina(n1710), .dinb(n791), .dout(n1711));
  jand g01494(.dina(n1710), .dinb(n791), .dout(n1712));
  jnot g01495(.din(n1523), .dout(n1713));
  jxor g01496(.dina(n1517), .dinb(n796), .dout(n1714));
  jor  g01497(.dina(n1714), .dinb(n1646), .dout(n1715));
  jxor g01498(.dina(n1715), .dinb(n1713), .dout(n1716));
  jnot g01499(.din(n1716), .dout(n1717));
  jor  g01500(.dina(n1717), .dinb(n1712), .dout(n1718));
  jand g01501(.dina(n1718), .dinb(n1711), .dout(n1719));
  jor  g01502(.dina(n1719), .dinb(n595), .dout(n1720));
  jnot g01503(.din(n1528), .dout(n1721));
  jor  g01504(.dina(n1721), .dinb(n1526), .dout(n1722));
  jor  g01505(.dina(n1722), .dinb(n1646), .dout(n1723));
  jxor g01506(.dina(n1723), .dinb(n1537), .dout(n1724));
  jand g01507(.dina(n1711), .dinb(n595), .dout(n1725));
  jand g01508(.dina(n1725), .dinb(n1718), .dout(n1726));
  jor  g01509(.dina(n1726), .dinb(n1724), .dout(n1727));
  jand g01510(.dina(n1727), .dinb(n1720), .dout(n1728));
  jor  g01511(.dina(n1728), .dinb(n590), .dout(n1729));
  jand g01512(.dina(n1728), .dinb(n590), .dout(n1730));
  jnot g01513(.din(n1544), .dout(n1731));
  jxor g01514(.dina(n1539), .dinb(n595), .dout(n1732));
  jor  g01515(.dina(n1732), .dinb(n1646), .dout(n1733));
  jxor g01516(.dina(n1733), .dinb(n1731), .dout(n1734));
  jnot g01517(.din(n1734), .dout(n1735));
  jor  g01518(.dina(n1735), .dinb(n1730), .dout(n1736));
  jand g01519(.dina(n1736), .dinb(n1729), .dout(n1737));
  jor  g01520(.dina(n1737), .dinb(n430), .dout(n1738));
  jand g01521(.dina(n1729), .dinb(n430), .dout(n1739));
  jand g01522(.dina(n1739), .dinb(n1736), .dout(n1740));
  jnot g01523(.din(n1547), .dout(n1741));
  jand g01524(.dina(asqrt[47] ), .dinb(n1741), .dout(n1742));
  jand g01525(.dina(n1742), .dinb(n1554), .dout(n1743));
  jor  g01526(.dina(n1743), .dinb(n1552), .dout(n1744));
  jand g01527(.dina(n1742), .dinb(n1555), .dout(n1745));
  jnot g01528(.din(n1745), .dout(n1746));
  jand g01529(.dina(n1746), .dinb(n1744), .dout(n1747));
  jnot g01530(.din(n1747), .dout(n1748));
  jor  g01531(.dina(n1748), .dinb(n1740), .dout(n1749));
  jand g01532(.dina(n1749), .dinb(n1738), .dout(n1750));
  jor  g01533(.dina(n1750), .dinb(n425), .dout(n1751));
  jxor g01534(.dina(n1556), .dinb(n430), .dout(n1752));
  jor  g01535(.dina(n1752), .dinb(n1646), .dout(n1753));
  jxor g01536(.dina(n1753), .dinb(n1561), .dout(n1754));
  jand g01537(.dina(n1750), .dinb(n425), .dout(n1755));
  jor  g01538(.dina(n1755), .dinb(n1754), .dout(n1756));
  jand g01539(.dina(n1756), .dinb(n1751), .dout(n1757));
  jor  g01540(.dina(n1757), .dinb(n305), .dout(n1758));
  jnot g01541(.din(n1566), .dout(n1759));
  jor  g01542(.dina(n1759), .dinb(n1564), .dout(n1760));
  jor  g01543(.dina(n1760), .dinb(n1646), .dout(n1761));
  jxor g01544(.dina(n1761), .dinb(n1575), .dout(n1762));
  jand g01545(.dina(n1751), .dinb(n305), .dout(n1763));
  jand g01546(.dina(n1763), .dinb(n1756), .dout(n1764));
  jor  g01547(.dina(n1764), .dinb(n1762), .dout(n1765));
  jand g01548(.dina(n1765), .dinb(n1758), .dout(n1766));
  jor  g01549(.dina(n1766), .dinb(n290), .dout(n1767));
  jand g01550(.dina(n1766), .dinb(n290), .dout(n1768));
  jnot g01551(.din(n1578), .dout(n1769));
  jand g01552(.dina(asqrt[47] ), .dinb(n1769), .dout(n1770));
  jand g01553(.dina(n1770), .dinb(n1583), .dout(n1771));
  jor  g01554(.dina(n1771), .dinb(n1582), .dout(n1772));
  jand g01555(.dina(n1770), .dinb(n1584), .dout(n1773));
  jnot g01556(.din(n1773), .dout(n1774));
  jand g01557(.dina(n1774), .dinb(n1772), .dout(n1775));
  jnot g01558(.din(n1775), .dout(n1776));
  jor  g01559(.dina(n1776), .dinb(n1768), .dout(n1777));
  jand g01560(.dina(n1777), .dinb(n1767), .dout(n1778));
  jor  g01561(.dina(n1778), .dinb(n223), .dout(n1779));
  jand g01562(.dina(n1767), .dinb(n223), .dout(n1780));
  jand g01563(.dina(n1780), .dinb(n1777), .dout(n1781));
  jnot g01564(.din(n1586), .dout(n1782));
  jand g01565(.dina(asqrt[47] ), .dinb(n1782), .dout(n1783));
  jand g01566(.dina(n1783), .dinb(n1593), .dout(n1784));
  jor  g01567(.dina(n1784), .dinb(n1591), .dout(n1785));
  jand g01568(.dina(n1783), .dinb(n1594), .dout(n1786));
  jnot g01569(.din(n1786), .dout(n1787));
  jand g01570(.dina(n1787), .dinb(n1785), .dout(n1788));
  jnot g01571(.din(n1788), .dout(n1789));
  jor  g01572(.dina(n1789), .dinb(n1781), .dout(n1790));
  jand g01573(.dina(n1790), .dinb(n1779), .dout(n1791));
  jor  g01574(.dina(n1791), .dinb(n199), .dout(n1792));
  jand g01575(.dina(n1791), .dinb(n199), .dout(n1793));
  jxor g01576(.dina(n1595), .dinb(n223), .dout(n1794));
  jor  g01577(.dina(n1794), .dinb(n1646), .dout(n1795));
  jxor g01578(.dina(n1795), .dinb(n1606), .dout(n1796));
  jor  g01579(.dina(n1796), .dinb(n1793), .dout(n1797));
  jand g01580(.dina(n1797), .dinb(n1792), .dout(n1798));
  jnot g01581(.din(n1611), .dout(n1799));
  jor  g01582(.dina(n1799), .dinb(n1609), .dout(n1800));
  jor  g01583(.dina(n1800), .dinb(n1646), .dout(n1801));
  jxor g01584(.dina(n1801), .dinb(n1620), .dout(n1802));
  jand g01585(.dina(asqrt[47] ), .dinb(n1634), .dout(n1803));
  jand g01586(.dina(n1803), .dinb(n1622), .dout(n1804));
  jor  g01587(.dina(n1804), .dinb(n1666), .dout(n1805));
  jor  g01588(.dina(n1805), .dinb(n1802), .dout(n1806));
  jor  g01589(.dina(n1806), .dinb(n1798), .dout(n1807));
  jand g01590(.dina(n1807), .dinb(n194), .dout(n1808));
  jand g01591(.dina(n1802), .dinb(n1798), .dout(n1809));
  jor  g01592(.dina(n1803), .dinb(n1622), .dout(n1810));
  jand g01593(.dina(n1634), .dinb(n1622), .dout(n1811));
  jor  g01594(.dina(n1811), .dinb(n194), .dout(n1812));
  jnot g01595(.din(n1812), .dout(n1813));
  jand g01596(.dina(n1813), .dinb(n1810), .dout(n1814));
  jor  g01597(.dina(n1814), .dinb(n1809), .dout(n1817));
  jor  g01598(.dina(n1817), .dinb(n1808), .dout(asqrt[46] ));
  jand g01599(.dina(asqrt[46] ), .dinb(a[92] ), .dout(n1819));
  jnot g01600(.din(a[90] ), .dout(n1820));
  jnot g01601(.din(a[91] ), .dout(n1821));
  jand g01602(.dina(n1649), .dinb(n1821), .dout(n1822));
  jand g01603(.dina(n1822), .dinb(n1820), .dout(n1823));
  jor  g01604(.dina(n1823), .dinb(n1819), .dout(n1824));
  jand g01605(.dina(n1824), .dinb(asqrt[47] ), .dout(n1825));
  jand g01606(.dina(asqrt[46] ), .dinb(n1649), .dout(n1826));
  jxor g01607(.dina(n1826), .dinb(n1650), .dout(n1827));
  jor  g01608(.dina(n1824), .dinb(asqrt[47] ), .dout(n1828));
  jand g01609(.dina(n1828), .dinb(n1827), .dout(n1829));
  jor  g01610(.dina(n1829), .dinb(n1825), .dout(n1830));
  jand g01611(.dina(n1830), .dinb(asqrt[48] ), .dout(n1831));
  jor  g01612(.dina(n1825), .dinb(asqrt[48] ), .dout(n1832));
  jor  g01613(.dina(n1832), .dinb(n1829), .dout(n1833));
  jand g01614(.dina(n1826), .dinb(n1650), .dout(n1834));
  jnot g01615(.din(n1808), .dout(n1835));
  jnot g01616(.din(n1809), .dout(n1836));
  jnot g01617(.din(n1814), .dout(n1837));
  jand g01618(.dina(n1837), .dinb(asqrt[47] ), .dout(n1838));
  jand g01619(.dina(n1838), .dinb(n1836), .dout(n1839));
  jand g01620(.dina(n1839), .dinb(n1835), .dout(n1840));
  jor  g01621(.dina(n1840), .dinb(n1834), .dout(n1841));
  jxor g01622(.dina(n1841), .dinb(n1475), .dout(n1842));
  jand g01623(.dina(n1842), .dinb(n1833), .dout(n1843));
  jor  g01624(.dina(n1843), .dinb(n1831), .dout(n1844));
  jand g01625(.dina(n1844), .dinb(asqrt[49] ), .dout(n1845));
  jor  g01626(.dina(n1844), .dinb(asqrt[49] ), .dout(n1846));
  jxor g01627(.dina(n1654), .dinb(n1641), .dout(n1847));
  jand g01628(.dina(n1847), .dinb(asqrt[46] ), .dout(n1848));
  jxor g01629(.dina(n1848), .dinb(n1657), .dout(n1849));
  jnot g01630(.din(n1849), .dout(n1850));
  jand g01631(.dina(n1850), .dinb(n1846), .dout(n1851));
  jor  g01632(.dina(n1851), .dinb(n1845), .dout(n1852));
  jand g01633(.dina(n1852), .dinb(asqrt[50] ), .dout(n1853));
  jnot g01634(.din(n1663), .dout(n1854));
  jand g01635(.dina(n1854), .dinb(n1661), .dout(n1855));
  jand g01636(.dina(n1855), .dinb(asqrt[46] ), .dout(n1856));
  jxor g01637(.dina(n1856), .dinb(n1671), .dout(n1857));
  jnot g01638(.din(n1857), .dout(n1858));
  jor  g01639(.dina(n1845), .dinb(asqrt[50] ), .dout(n1859));
  jor  g01640(.dina(n1859), .dinb(n1851), .dout(n1860));
  jand g01641(.dina(n1860), .dinb(n1858), .dout(n1861));
  jor  g01642(.dina(n1861), .dinb(n1853), .dout(n1862));
  jand g01643(.dina(n1862), .dinb(asqrt[51] ), .dout(n1863));
  jor  g01644(.dina(n1862), .dinb(asqrt[51] ), .dout(n1864));
  jnot g01645(.din(n1678), .dout(n1865));
  jxor g01646(.dina(n1673), .dinb(n1312), .dout(n1866));
  jand g01647(.dina(n1866), .dinb(asqrt[46] ), .dout(n1867));
  jxor g01648(.dina(n1867), .dinb(n1865), .dout(n1868));
  jand g01649(.dina(n1868), .dinb(n1864), .dout(n1869));
  jor  g01650(.dina(n1869), .dinb(n1863), .dout(n1870));
  jand g01651(.dina(n1870), .dinb(asqrt[52] ), .dout(n1871));
  jor  g01652(.dina(n1863), .dinb(asqrt[52] ), .dout(n1872));
  jor  g01653(.dina(n1872), .dinb(n1869), .dout(n1873));
  jnot g01654(.din(n1685), .dout(n1874));
  jnot g01655(.din(n1687), .dout(n1875));
  jand g01656(.dina(asqrt[46] ), .dinb(n1681), .dout(n1876));
  jand g01657(.dina(n1876), .dinb(n1875), .dout(n1877));
  jor  g01658(.dina(n1877), .dinb(n1874), .dout(n1878));
  jnot g01659(.din(n1688), .dout(n1879));
  jand g01660(.dina(n1876), .dinb(n1879), .dout(n1880));
  jnot g01661(.din(n1880), .dout(n1881));
  jand g01662(.dina(n1881), .dinb(n1878), .dout(n1882));
  jand g01663(.dina(n1882), .dinb(n1873), .dout(n1883));
  jor  g01664(.dina(n1883), .dinb(n1871), .dout(n1884));
  jand g01665(.dina(n1884), .dinb(asqrt[53] ), .dout(n1885));
  jor  g01666(.dina(n1884), .dinb(asqrt[53] ), .dout(n1886));
  jxor g01667(.dina(n1689), .dinb(n1034), .dout(n1887));
  jand g01668(.dina(n1887), .dinb(asqrt[46] ), .dout(n1888));
  jxor g01669(.dina(n1888), .dinb(n1694), .dout(n1889));
  jand g01670(.dina(n1889), .dinb(n1886), .dout(n1890));
  jor  g01671(.dina(n1890), .dinb(n1885), .dout(n1891));
  jand g01672(.dina(n1891), .dinb(asqrt[54] ), .dout(n1892));
  jnot g01673(.din(n1700), .dout(n1893));
  jand g01674(.dina(n1893), .dinb(n1698), .dout(n1894));
  jand g01675(.dina(n1894), .dinb(asqrt[46] ), .dout(n1895));
  jxor g01676(.dina(n1895), .dinb(n1708), .dout(n1896));
  jnot g01677(.din(n1896), .dout(n1897));
  jor  g01678(.dina(n1885), .dinb(asqrt[54] ), .dout(n1898));
  jor  g01679(.dina(n1898), .dinb(n1890), .dout(n1899));
  jand g01680(.dina(n1899), .dinb(n1897), .dout(n1900));
  jor  g01681(.dina(n1900), .dinb(n1892), .dout(n1901));
  jand g01682(.dina(n1901), .dinb(asqrt[55] ), .dout(n1902));
  jor  g01683(.dina(n1901), .dinb(asqrt[55] ), .dout(n1903));
  jxor g01684(.dina(n1710), .dinb(n791), .dout(n1904));
  jand g01685(.dina(n1904), .dinb(asqrt[46] ), .dout(n1905));
  jxor g01686(.dina(n1905), .dinb(n1716), .dout(n1906));
  jand g01687(.dina(n1906), .dinb(n1903), .dout(n1907));
  jor  g01688(.dina(n1907), .dinb(n1902), .dout(n1908));
  jand g01689(.dina(n1908), .dinb(asqrt[56] ), .dout(n1909));
  jor  g01690(.dina(n1902), .dinb(asqrt[56] ), .dout(n1910));
  jor  g01691(.dina(n1910), .dinb(n1907), .dout(n1911));
  jnot g01692(.din(n1724), .dout(n1912));
  jnot g01693(.din(n1726), .dout(n1913));
  jand g01694(.dina(asqrt[46] ), .dinb(n1720), .dout(n1914));
  jand g01695(.dina(n1914), .dinb(n1913), .dout(n1915));
  jor  g01696(.dina(n1915), .dinb(n1912), .dout(n1916));
  jnot g01697(.din(n1727), .dout(n1917));
  jand g01698(.dina(n1914), .dinb(n1917), .dout(n1918));
  jnot g01699(.din(n1918), .dout(n1919));
  jand g01700(.dina(n1919), .dinb(n1916), .dout(n1920));
  jand g01701(.dina(n1920), .dinb(n1911), .dout(n1921));
  jor  g01702(.dina(n1921), .dinb(n1909), .dout(n1922));
  jand g01703(.dina(n1922), .dinb(asqrt[57] ), .dout(n1923));
  jxor g01704(.dina(n1728), .dinb(n590), .dout(n1924));
  jand g01705(.dina(n1924), .dinb(asqrt[46] ), .dout(n1925));
  jxor g01706(.dina(n1925), .dinb(n1735), .dout(n1926));
  jnot g01707(.din(n1926), .dout(n1927));
  jor  g01708(.dina(n1922), .dinb(asqrt[57] ), .dout(n1928));
  jand g01709(.dina(n1928), .dinb(n1927), .dout(n1929));
  jor  g01710(.dina(n1929), .dinb(n1923), .dout(n1930));
  jand g01711(.dina(n1930), .dinb(asqrt[58] ), .dout(n1931));
  jnot g01712(.din(n1740), .dout(n1932));
  jand g01713(.dina(n1932), .dinb(n1738), .dout(n1933));
  jand g01714(.dina(n1933), .dinb(asqrt[46] ), .dout(n1934));
  jxor g01715(.dina(n1934), .dinb(n1748), .dout(n1935));
  jnot g01716(.din(n1935), .dout(n1936));
  jor  g01717(.dina(n1923), .dinb(asqrt[58] ), .dout(n1937));
  jor  g01718(.dina(n1937), .dinb(n1929), .dout(n1938));
  jand g01719(.dina(n1938), .dinb(n1936), .dout(n1939));
  jor  g01720(.dina(n1939), .dinb(n1931), .dout(n1940));
  jand g01721(.dina(n1940), .dinb(asqrt[59] ), .dout(n1941));
  jor  g01722(.dina(n1940), .dinb(asqrt[59] ), .dout(n1942));
  jnot g01723(.din(n1754), .dout(n1943));
  jnot g01724(.din(n1755), .dout(n1944));
  jand g01725(.dina(asqrt[46] ), .dinb(n1751), .dout(n1945));
  jand g01726(.dina(n1945), .dinb(n1944), .dout(n1946));
  jor  g01727(.dina(n1946), .dinb(n1943), .dout(n1947));
  jnot g01728(.din(n1756), .dout(n1948));
  jand g01729(.dina(n1945), .dinb(n1948), .dout(n1949));
  jnot g01730(.din(n1949), .dout(n1950));
  jand g01731(.dina(n1950), .dinb(n1947), .dout(n1951));
  jand g01732(.dina(n1951), .dinb(n1942), .dout(n1952));
  jor  g01733(.dina(n1952), .dinb(n1941), .dout(n1953));
  jand g01734(.dina(n1953), .dinb(asqrt[60] ), .dout(n1954));
  jor  g01735(.dina(n1941), .dinb(asqrt[60] ), .dout(n1955));
  jor  g01736(.dina(n1955), .dinb(n1952), .dout(n1956));
  jnot g01737(.din(n1762), .dout(n1957));
  jnot g01738(.din(n1764), .dout(n1958));
  jand g01739(.dina(asqrt[46] ), .dinb(n1758), .dout(n1959));
  jand g01740(.dina(n1959), .dinb(n1958), .dout(n1960));
  jor  g01741(.dina(n1960), .dinb(n1957), .dout(n1961));
  jnot g01742(.din(n1765), .dout(n1962));
  jand g01743(.dina(n1959), .dinb(n1962), .dout(n1963));
  jnot g01744(.din(n1963), .dout(n1964));
  jand g01745(.dina(n1964), .dinb(n1961), .dout(n1965));
  jand g01746(.dina(n1965), .dinb(n1956), .dout(n1966));
  jor  g01747(.dina(n1966), .dinb(n1954), .dout(n1967));
  jand g01748(.dina(n1967), .dinb(asqrt[61] ), .dout(n1968));
  jxor g01749(.dina(n1766), .dinb(n290), .dout(n1969));
  jand g01750(.dina(n1969), .dinb(asqrt[46] ), .dout(n1970));
  jxor g01751(.dina(n1970), .dinb(n1776), .dout(n1971));
  jnot g01752(.din(n1971), .dout(n1972));
  jor  g01753(.dina(n1967), .dinb(asqrt[61] ), .dout(n1973));
  jand g01754(.dina(n1973), .dinb(n1972), .dout(n1974));
  jor  g01755(.dina(n1974), .dinb(n1968), .dout(n1975));
  jand g01756(.dina(n1975), .dinb(asqrt[62] ), .dout(n1976));
  jnot g01757(.din(n1781), .dout(n1977));
  jand g01758(.dina(n1977), .dinb(n1779), .dout(n1978));
  jand g01759(.dina(n1978), .dinb(asqrt[46] ), .dout(n1979));
  jxor g01760(.dina(n1979), .dinb(n1789), .dout(n1980));
  jnot g01761(.din(n1980), .dout(n1981));
  jor  g01762(.dina(n1968), .dinb(asqrt[62] ), .dout(n1982));
  jor  g01763(.dina(n1982), .dinb(n1974), .dout(n1983));
  jand g01764(.dina(n1983), .dinb(n1981), .dout(n1984));
  jor  g01765(.dina(n1984), .dinb(n1976), .dout(n1985));
  jxor g01766(.dina(n1791), .dinb(n199), .dout(n1986));
  jand g01767(.dina(n1986), .dinb(asqrt[46] ), .dout(n1987));
  jxor g01768(.dina(n1987), .dinb(n1796), .dout(n1988));
  jnot g01769(.din(n1798), .dout(n1989));
  jnot g01770(.din(n1802), .dout(n1990));
  jand g01771(.dina(asqrt[46] ), .dinb(n1990), .dout(n1991));
  jand g01772(.dina(n1991), .dinb(n1989), .dout(n1992));
  jor  g01773(.dina(n1992), .dinb(n1809), .dout(n1993));
  jor  g01774(.dina(n1993), .dinb(n1988), .dout(n1994));
  jnot g01775(.din(n1994), .dout(n1995));
  jand g01776(.dina(n1995), .dinb(n1985), .dout(n1996));
  jor  g01777(.dina(n1996), .dinb(asqrt[63] ), .dout(n1997));
  jnot g01778(.din(n1988), .dout(n1998));
  jor  g01779(.dina(n1998), .dinb(n1985), .dout(n1999));
  jor  g01780(.dina(n1991), .dinb(n1989), .dout(n2000));
  jand g01781(.dina(n1990), .dinb(n1989), .dout(n2001));
  jor  g01782(.dina(n2001), .dinb(n194), .dout(n2002));
  jnot g01783(.din(n2002), .dout(n2003));
  jand g01784(.dina(n2003), .dinb(n2000), .dout(n2004));
  jnot g01785(.din(asqrt[46] ), .dout(n2005));
  jnot g01786(.din(n2004), .dout(n2008));
  jand g01787(.dina(n2008), .dinb(n1999), .dout(n2009));
  jand g01788(.dina(n2009), .dinb(n1997), .dout(n2010));
  jnot g01789(.din(n2010), .dout(asqrt[45] ));
  jor  g01790(.dina(n2010), .dinb(n1820), .dout(n2012));
  jnot g01791(.din(a[88] ), .dout(n2013));
  jnot g01792(.din(a[89] ), .dout(n2014));
  jand g01793(.dina(n1820), .dinb(n2014), .dout(n2015));
  jand g01794(.dina(n2015), .dinb(n2013), .dout(n2016));
  jnot g01795(.din(n2016), .dout(n2017));
  jand g01796(.dina(n2017), .dinb(n2012), .dout(n2018));
  jor  g01797(.dina(n2018), .dinb(n2005), .dout(n2019));
  jor  g01798(.dina(n2010), .dinb(a[90] ), .dout(n2020));
  jxor g01799(.dina(n2020), .dinb(n1821), .dout(n2021));
  jand g01800(.dina(n2018), .dinb(n2005), .dout(n2022));
  jor  g01801(.dina(n2022), .dinb(n2021), .dout(n2023));
  jand g01802(.dina(n2023), .dinb(n2019), .dout(n2024));
  jor  g01803(.dina(n2024), .dinb(n1646), .dout(n2025));
  jand g01804(.dina(n2019), .dinb(n1646), .dout(n2026));
  jand g01805(.dina(n2026), .dinb(n2023), .dout(n2027));
  jor  g01806(.dina(n2020), .dinb(a[91] ), .dout(n2028));
  jnot g01807(.din(n1997), .dout(n2029));
  jnot g01808(.din(n1999), .dout(n2030));
  jor  g01809(.dina(n2004), .dinb(n2005), .dout(n2031));
  jor  g01810(.dina(n2031), .dinb(n2030), .dout(n2032));
  jor  g01811(.dina(n2032), .dinb(n2029), .dout(n2033));
  jand g01812(.dina(n2033), .dinb(n2028), .dout(n2034));
  jxor g01813(.dina(n2034), .dinb(n1649), .dout(n2035));
  jor  g01814(.dina(n2035), .dinb(n2027), .dout(n2036));
  jand g01815(.dina(n2036), .dinb(n2025), .dout(n2037));
  jor  g01816(.dina(n2037), .dinb(n1641), .dout(n2038));
  jand g01817(.dina(n2037), .dinb(n1641), .dout(n2039));
  jxor g01818(.dina(n1824), .dinb(n1646), .dout(n2040));
  jor  g01819(.dina(n2040), .dinb(n2010), .dout(n2041));
  jxor g01820(.dina(n2041), .dinb(n1827), .dout(n2042));
  jor  g01821(.dina(n2042), .dinb(n2039), .dout(n2043));
  jand g01822(.dina(n2043), .dinb(n2038), .dout(n2044));
  jor  g01823(.dina(n2044), .dinb(n1317), .dout(n2045));
  jnot g01824(.din(n1833), .dout(n2046));
  jor  g01825(.dina(n2046), .dinb(n1831), .dout(n2047));
  jor  g01826(.dina(n2047), .dinb(n2010), .dout(n2048));
  jxor g01827(.dina(n2048), .dinb(n1842), .dout(n2049));
  jand g01828(.dina(n2038), .dinb(n1317), .dout(n2050));
  jand g01829(.dina(n2050), .dinb(n2043), .dout(n2051));
  jor  g01830(.dina(n2051), .dinb(n2049), .dout(n2052));
  jand g01831(.dina(n2052), .dinb(n2045), .dout(n2053));
  jor  g01832(.dina(n2053), .dinb(n1312), .dout(n2054));
  jand g01833(.dina(n2053), .dinb(n1312), .dout(n2055));
  jxor g01834(.dina(n1844), .dinb(n1317), .dout(n2056));
  jor  g01835(.dina(n2056), .dinb(n2010), .dout(n2057));
  jxor g01836(.dina(n2057), .dinb(n1849), .dout(n2058));
  jnot g01837(.din(n2058), .dout(n2059));
  jor  g01838(.dina(n2059), .dinb(n2055), .dout(n2060));
  jand g01839(.dina(n2060), .dinb(n2054), .dout(n2061));
  jor  g01840(.dina(n2061), .dinb(n1039), .dout(n2062));
  jand g01841(.dina(n2054), .dinb(n1039), .dout(n2063));
  jand g01842(.dina(n2063), .dinb(n2060), .dout(n2064));
  jnot g01843(.din(n1853), .dout(n2065));
  jand g01844(.dina(asqrt[45] ), .dinb(n2065), .dout(n2066));
  jand g01845(.dina(n2066), .dinb(n1860), .dout(n2067));
  jor  g01846(.dina(n2067), .dinb(n1858), .dout(n2068));
  jand g01847(.dina(n2066), .dinb(n1861), .dout(n2069));
  jnot g01848(.din(n2069), .dout(n2070));
  jand g01849(.dina(n2070), .dinb(n2068), .dout(n2071));
  jnot g01850(.din(n2071), .dout(n2072));
  jor  g01851(.dina(n2072), .dinb(n2064), .dout(n2073));
  jand g01852(.dina(n2073), .dinb(n2062), .dout(n2074));
  jor  g01853(.dina(n2074), .dinb(n1034), .dout(n2075));
  jand g01854(.dina(n2074), .dinb(n1034), .dout(n2076));
  jnot g01855(.din(n1868), .dout(n2077));
  jxor g01856(.dina(n1862), .dinb(n1039), .dout(n2078));
  jor  g01857(.dina(n2078), .dinb(n2010), .dout(n2079));
  jxor g01858(.dina(n2079), .dinb(n2077), .dout(n2080));
  jnot g01859(.din(n2080), .dout(n2081));
  jor  g01860(.dina(n2081), .dinb(n2076), .dout(n2082));
  jand g01861(.dina(n2082), .dinb(n2075), .dout(n2083));
  jor  g01862(.dina(n2083), .dinb(n796), .dout(n2084));
  jnot g01863(.din(n1873), .dout(n2085));
  jor  g01864(.dina(n2085), .dinb(n1871), .dout(n2086));
  jor  g01865(.dina(n2086), .dinb(n2010), .dout(n2087));
  jxor g01866(.dina(n2087), .dinb(n1882), .dout(n2088));
  jand g01867(.dina(n2075), .dinb(n796), .dout(n2089));
  jand g01868(.dina(n2089), .dinb(n2082), .dout(n2090));
  jor  g01869(.dina(n2090), .dinb(n2088), .dout(n2091));
  jand g01870(.dina(n2091), .dinb(n2084), .dout(n2092));
  jor  g01871(.dina(n2092), .dinb(n791), .dout(n2093));
  jand g01872(.dina(n2092), .dinb(n791), .dout(n2094));
  jnot g01873(.din(n1889), .dout(n2095));
  jxor g01874(.dina(n1884), .dinb(n796), .dout(n2096));
  jor  g01875(.dina(n2096), .dinb(n2010), .dout(n2097));
  jxor g01876(.dina(n2097), .dinb(n2095), .dout(n2098));
  jnot g01877(.din(n2098), .dout(n2099));
  jor  g01878(.dina(n2099), .dinb(n2094), .dout(n2100));
  jand g01879(.dina(n2100), .dinb(n2093), .dout(n2101));
  jor  g01880(.dina(n2101), .dinb(n595), .dout(n2102));
  jand g01881(.dina(n2093), .dinb(n595), .dout(n2103));
  jand g01882(.dina(n2103), .dinb(n2100), .dout(n2104));
  jnot g01883(.din(n1892), .dout(n2105));
  jand g01884(.dina(asqrt[45] ), .dinb(n2105), .dout(n2106));
  jand g01885(.dina(n2106), .dinb(n1899), .dout(n2107));
  jor  g01886(.dina(n2107), .dinb(n1897), .dout(n2108));
  jand g01887(.dina(n2106), .dinb(n1900), .dout(n2109));
  jnot g01888(.din(n2109), .dout(n2110));
  jand g01889(.dina(n2110), .dinb(n2108), .dout(n2111));
  jnot g01890(.din(n2111), .dout(n2112));
  jor  g01891(.dina(n2112), .dinb(n2104), .dout(n2113));
  jand g01892(.dina(n2113), .dinb(n2102), .dout(n2114));
  jor  g01893(.dina(n2114), .dinb(n590), .dout(n2115));
  jxor g01894(.dina(n1901), .dinb(n595), .dout(n2116));
  jor  g01895(.dina(n2116), .dinb(n2010), .dout(n2117));
  jxor g01896(.dina(n2117), .dinb(n1906), .dout(n2118));
  jand g01897(.dina(n2114), .dinb(n590), .dout(n2119));
  jor  g01898(.dina(n2119), .dinb(n2118), .dout(n2120));
  jand g01899(.dina(n2120), .dinb(n2115), .dout(n2121));
  jor  g01900(.dina(n2121), .dinb(n430), .dout(n2122));
  jnot g01901(.din(n1911), .dout(n2123));
  jor  g01902(.dina(n2123), .dinb(n1909), .dout(n2124));
  jor  g01903(.dina(n2124), .dinb(n2010), .dout(n2125));
  jxor g01904(.dina(n2125), .dinb(n1920), .dout(n2126));
  jand g01905(.dina(n2115), .dinb(n430), .dout(n2127));
  jand g01906(.dina(n2127), .dinb(n2120), .dout(n2128));
  jor  g01907(.dina(n2128), .dinb(n2126), .dout(n2129));
  jand g01908(.dina(n2129), .dinb(n2122), .dout(n2130));
  jor  g01909(.dina(n2130), .dinb(n425), .dout(n2131));
  jand g01910(.dina(n2130), .dinb(n425), .dout(n2132));
  jnot g01911(.din(n1923), .dout(n2133));
  jand g01912(.dina(asqrt[45] ), .dinb(n2133), .dout(n2134));
  jand g01913(.dina(n2134), .dinb(n1928), .dout(n2135));
  jor  g01914(.dina(n2135), .dinb(n1927), .dout(n2136));
  jand g01915(.dina(n2134), .dinb(n1929), .dout(n2137));
  jnot g01916(.din(n2137), .dout(n2138));
  jand g01917(.dina(n2138), .dinb(n2136), .dout(n2139));
  jnot g01918(.din(n2139), .dout(n2140));
  jor  g01919(.dina(n2140), .dinb(n2132), .dout(n2141));
  jand g01920(.dina(n2141), .dinb(n2131), .dout(n2142));
  jor  g01921(.dina(n2142), .dinb(n305), .dout(n2143));
  jand g01922(.dina(n2131), .dinb(n305), .dout(n2144));
  jand g01923(.dina(n2144), .dinb(n2141), .dout(n2145));
  jnot g01924(.din(n1931), .dout(n2146));
  jand g01925(.dina(asqrt[45] ), .dinb(n2146), .dout(n2147));
  jand g01926(.dina(n2147), .dinb(n1938), .dout(n2148));
  jor  g01927(.dina(n2148), .dinb(n1936), .dout(n2149));
  jand g01928(.dina(n2147), .dinb(n1939), .dout(n2150));
  jnot g01929(.din(n2150), .dout(n2151));
  jand g01930(.dina(n2151), .dinb(n2149), .dout(n2152));
  jnot g01931(.din(n2152), .dout(n2153));
  jor  g01932(.dina(n2153), .dinb(n2145), .dout(n2154));
  jand g01933(.dina(n2154), .dinb(n2143), .dout(n2155));
  jor  g01934(.dina(n2155), .dinb(n290), .dout(n2156));
  jxor g01935(.dina(n1940), .dinb(n305), .dout(n2157));
  jor  g01936(.dina(n2157), .dinb(n2010), .dout(n2158));
  jxor g01937(.dina(n2158), .dinb(n1951), .dout(n2159));
  jand g01938(.dina(n2155), .dinb(n290), .dout(n2160));
  jor  g01939(.dina(n2160), .dinb(n2159), .dout(n2161));
  jand g01940(.dina(n2161), .dinb(n2156), .dout(n2162));
  jor  g01941(.dina(n2162), .dinb(n223), .dout(n2163));
  jnot g01942(.din(n1956), .dout(n2164));
  jor  g01943(.dina(n2164), .dinb(n1954), .dout(n2165));
  jor  g01944(.dina(n2165), .dinb(n2010), .dout(n2166));
  jxor g01945(.dina(n2166), .dinb(n1965), .dout(n2167));
  jand g01946(.dina(n2156), .dinb(n223), .dout(n2168));
  jand g01947(.dina(n2168), .dinb(n2161), .dout(n2169));
  jor  g01948(.dina(n2169), .dinb(n2167), .dout(n2170));
  jand g01949(.dina(n2170), .dinb(n2163), .dout(n2171));
  jor  g01950(.dina(n2171), .dinb(n199), .dout(n2172));
  jand g01951(.dina(n2171), .dinb(n199), .dout(n2173));
  jnot g01952(.din(n1968), .dout(n2174));
  jand g01953(.dina(asqrt[45] ), .dinb(n2174), .dout(n2175));
  jand g01954(.dina(n2175), .dinb(n1973), .dout(n2176));
  jor  g01955(.dina(n2176), .dinb(n1972), .dout(n2177));
  jand g01956(.dina(n2175), .dinb(n1974), .dout(n2178));
  jnot g01957(.din(n2178), .dout(n2179));
  jand g01958(.dina(n2179), .dinb(n2177), .dout(n2180));
  jnot g01959(.din(n2180), .dout(n2181));
  jor  g01960(.dina(n2181), .dinb(n2173), .dout(n2182));
  jand g01961(.dina(n2182), .dinb(n2172), .dout(n2183));
  jnot g01962(.din(n1976), .dout(n2184));
  jand g01963(.dina(asqrt[45] ), .dinb(n2184), .dout(n2185));
  jand g01964(.dina(n2185), .dinb(n1983), .dout(n2186));
  jor  g01965(.dina(n2186), .dinb(n1981), .dout(n2187));
  jand g01966(.dina(n2185), .dinb(n1984), .dout(n2188));
  jnot g01967(.din(n2188), .dout(n2189));
  jand g01968(.dina(n2189), .dinb(n2187), .dout(n2190));
  jnot g01969(.din(n2190), .dout(n2191));
  jand g01970(.dina(asqrt[45] ), .dinb(n1998), .dout(n2192));
  jand g01971(.dina(n2192), .dinb(n1985), .dout(n2193));
  jor  g01972(.dina(n2193), .dinb(n2030), .dout(n2194));
  jor  g01973(.dina(n2194), .dinb(n2191), .dout(n2195));
  jor  g01974(.dina(n2195), .dinb(n2183), .dout(n2196));
  jand g01975(.dina(n2196), .dinb(n194), .dout(n2197));
  jand g01976(.dina(n2191), .dinb(n2183), .dout(n2198));
  jor  g01977(.dina(n2192), .dinb(n1985), .dout(n2199));
  jand g01978(.dina(n1998), .dinb(n1985), .dout(n2200));
  jor  g01979(.dina(n2200), .dinb(n194), .dout(n2201));
  jnot g01980(.din(n2201), .dout(n2202));
  jand g01981(.dina(n2202), .dinb(n2199), .dout(n2203));
  jor  g01982(.dina(n2203), .dinb(n2198), .dout(n2206));
  jor  g01983(.dina(n2206), .dinb(n2197), .dout(asqrt[44] ));
  jand g01984(.dina(asqrt[44] ), .dinb(a[88] ), .dout(n2208));
  jnot g01985(.din(a[86] ), .dout(n2209));
  jnot g01986(.din(a[87] ), .dout(n2210));
  jand g01987(.dina(n2013), .dinb(n2210), .dout(n2211));
  jand g01988(.dina(n2211), .dinb(n2209), .dout(n2212));
  jor  g01989(.dina(n2212), .dinb(n2208), .dout(n2213));
  jand g01990(.dina(n2213), .dinb(asqrt[45] ), .dout(n2214));
  jand g01991(.dina(asqrt[44] ), .dinb(n2013), .dout(n2215));
  jxor g01992(.dina(n2215), .dinb(n2014), .dout(n2216));
  jor  g01993(.dina(n2213), .dinb(asqrt[45] ), .dout(n2217));
  jand g01994(.dina(n2217), .dinb(n2216), .dout(n2218));
  jor  g01995(.dina(n2218), .dinb(n2214), .dout(n2219));
  jand g01996(.dina(n2219), .dinb(asqrt[46] ), .dout(n2220));
  jor  g01997(.dina(n2214), .dinb(asqrt[46] ), .dout(n2221));
  jor  g01998(.dina(n2221), .dinb(n2218), .dout(n2222));
  jand g01999(.dina(n2215), .dinb(n2014), .dout(n2223));
  jnot g02000(.din(n2197), .dout(n2224));
  jnot g02001(.din(n2198), .dout(n2225));
  jnot g02002(.din(n2203), .dout(n2226));
  jand g02003(.dina(n2226), .dinb(asqrt[45] ), .dout(n2227));
  jand g02004(.dina(n2227), .dinb(n2225), .dout(n2228));
  jand g02005(.dina(n2228), .dinb(n2224), .dout(n2229));
  jor  g02006(.dina(n2229), .dinb(n2223), .dout(n2230));
  jxor g02007(.dina(n2230), .dinb(n1820), .dout(n2231));
  jand g02008(.dina(n2231), .dinb(n2222), .dout(n2232));
  jor  g02009(.dina(n2232), .dinb(n2220), .dout(n2233));
  jand g02010(.dina(n2233), .dinb(asqrt[47] ), .dout(n2234));
  jor  g02011(.dina(n2233), .dinb(asqrt[47] ), .dout(n2235));
  jxor g02012(.dina(n2018), .dinb(n2005), .dout(n2236));
  jand g02013(.dina(n2236), .dinb(asqrt[44] ), .dout(n2237));
  jxor g02014(.dina(n2237), .dinb(n2021), .dout(n2238));
  jnot g02015(.din(n2238), .dout(n2239));
  jand g02016(.dina(n2239), .dinb(n2235), .dout(n2240));
  jor  g02017(.dina(n2240), .dinb(n2234), .dout(n2241));
  jand g02018(.dina(n2241), .dinb(asqrt[48] ), .dout(n2242));
  jnot g02019(.din(n2027), .dout(n2243));
  jand g02020(.dina(n2243), .dinb(n2025), .dout(n2244));
  jand g02021(.dina(n2244), .dinb(asqrt[44] ), .dout(n2245));
  jxor g02022(.dina(n2245), .dinb(n2035), .dout(n2246));
  jnot g02023(.din(n2246), .dout(n2247));
  jor  g02024(.dina(n2234), .dinb(asqrt[48] ), .dout(n2248));
  jor  g02025(.dina(n2248), .dinb(n2240), .dout(n2249));
  jand g02026(.dina(n2249), .dinb(n2247), .dout(n2250));
  jor  g02027(.dina(n2250), .dinb(n2242), .dout(n2251));
  jand g02028(.dina(n2251), .dinb(asqrt[49] ), .dout(n2252));
  jor  g02029(.dina(n2251), .dinb(asqrt[49] ), .dout(n2253));
  jnot g02030(.din(n2042), .dout(n2254));
  jxor g02031(.dina(n2037), .dinb(n1641), .dout(n2255));
  jand g02032(.dina(n2255), .dinb(asqrt[44] ), .dout(n2256));
  jxor g02033(.dina(n2256), .dinb(n2254), .dout(n2257));
  jand g02034(.dina(n2257), .dinb(n2253), .dout(n2258));
  jor  g02035(.dina(n2258), .dinb(n2252), .dout(n2259));
  jand g02036(.dina(n2259), .dinb(asqrt[50] ), .dout(n2260));
  jor  g02037(.dina(n2252), .dinb(asqrt[50] ), .dout(n2261));
  jor  g02038(.dina(n2261), .dinb(n2258), .dout(n2262));
  jnot g02039(.din(n2049), .dout(n2263));
  jnot g02040(.din(n2051), .dout(n2264));
  jand g02041(.dina(asqrt[44] ), .dinb(n2045), .dout(n2265));
  jand g02042(.dina(n2265), .dinb(n2264), .dout(n2266));
  jor  g02043(.dina(n2266), .dinb(n2263), .dout(n2267));
  jnot g02044(.din(n2052), .dout(n2268));
  jand g02045(.dina(n2265), .dinb(n2268), .dout(n2269));
  jnot g02046(.din(n2269), .dout(n2270));
  jand g02047(.dina(n2270), .dinb(n2267), .dout(n2271));
  jand g02048(.dina(n2271), .dinb(n2262), .dout(n2272));
  jor  g02049(.dina(n2272), .dinb(n2260), .dout(n2273));
  jand g02050(.dina(n2273), .dinb(asqrt[51] ), .dout(n2274));
  jor  g02051(.dina(n2273), .dinb(asqrt[51] ), .dout(n2275));
  jxor g02052(.dina(n2053), .dinb(n1312), .dout(n2276));
  jand g02053(.dina(n2276), .dinb(asqrt[44] ), .dout(n2277));
  jxor g02054(.dina(n2277), .dinb(n2058), .dout(n2278));
  jand g02055(.dina(n2278), .dinb(n2275), .dout(n2279));
  jor  g02056(.dina(n2279), .dinb(n2274), .dout(n2280));
  jand g02057(.dina(n2280), .dinb(asqrt[52] ), .dout(n2281));
  jnot g02058(.din(n2064), .dout(n2282));
  jand g02059(.dina(n2282), .dinb(n2062), .dout(n2283));
  jand g02060(.dina(n2283), .dinb(asqrt[44] ), .dout(n2284));
  jxor g02061(.dina(n2284), .dinb(n2072), .dout(n2285));
  jnot g02062(.din(n2285), .dout(n2286));
  jor  g02063(.dina(n2274), .dinb(asqrt[52] ), .dout(n2287));
  jor  g02064(.dina(n2287), .dinb(n2279), .dout(n2288));
  jand g02065(.dina(n2288), .dinb(n2286), .dout(n2289));
  jor  g02066(.dina(n2289), .dinb(n2281), .dout(n2290));
  jand g02067(.dina(n2290), .dinb(asqrt[53] ), .dout(n2291));
  jor  g02068(.dina(n2290), .dinb(asqrt[53] ), .dout(n2292));
  jxor g02069(.dina(n2074), .dinb(n1034), .dout(n2293));
  jand g02070(.dina(n2293), .dinb(asqrt[44] ), .dout(n2294));
  jxor g02071(.dina(n2294), .dinb(n2080), .dout(n2295));
  jand g02072(.dina(n2295), .dinb(n2292), .dout(n2296));
  jor  g02073(.dina(n2296), .dinb(n2291), .dout(n2297));
  jand g02074(.dina(n2297), .dinb(asqrt[54] ), .dout(n2298));
  jor  g02075(.dina(n2291), .dinb(asqrt[54] ), .dout(n2299));
  jor  g02076(.dina(n2299), .dinb(n2296), .dout(n2300));
  jnot g02077(.din(n2088), .dout(n2301));
  jnot g02078(.din(n2090), .dout(n2302));
  jand g02079(.dina(asqrt[44] ), .dinb(n2084), .dout(n2303));
  jand g02080(.dina(n2303), .dinb(n2302), .dout(n2304));
  jor  g02081(.dina(n2304), .dinb(n2301), .dout(n2305));
  jnot g02082(.din(n2091), .dout(n2306));
  jand g02083(.dina(n2303), .dinb(n2306), .dout(n2307));
  jnot g02084(.din(n2307), .dout(n2308));
  jand g02085(.dina(n2308), .dinb(n2305), .dout(n2309));
  jand g02086(.dina(n2309), .dinb(n2300), .dout(n2310));
  jor  g02087(.dina(n2310), .dinb(n2298), .dout(n2311));
  jand g02088(.dina(n2311), .dinb(asqrt[55] ), .dout(n2312));
  jxor g02089(.dina(n2092), .dinb(n791), .dout(n2313));
  jand g02090(.dina(n2313), .dinb(asqrt[44] ), .dout(n2314));
  jxor g02091(.dina(n2314), .dinb(n2099), .dout(n2315));
  jnot g02092(.din(n2315), .dout(n2316));
  jor  g02093(.dina(n2311), .dinb(asqrt[55] ), .dout(n2317));
  jand g02094(.dina(n2317), .dinb(n2316), .dout(n2318));
  jor  g02095(.dina(n2318), .dinb(n2312), .dout(n2319));
  jand g02096(.dina(n2319), .dinb(asqrt[56] ), .dout(n2320));
  jnot g02097(.din(n2104), .dout(n2321));
  jand g02098(.dina(n2321), .dinb(n2102), .dout(n2322));
  jand g02099(.dina(n2322), .dinb(asqrt[44] ), .dout(n2323));
  jxor g02100(.dina(n2323), .dinb(n2112), .dout(n2324));
  jnot g02101(.din(n2324), .dout(n2325));
  jor  g02102(.dina(n2312), .dinb(asqrt[56] ), .dout(n2326));
  jor  g02103(.dina(n2326), .dinb(n2318), .dout(n2327));
  jand g02104(.dina(n2327), .dinb(n2325), .dout(n2328));
  jor  g02105(.dina(n2328), .dinb(n2320), .dout(n2329));
  jand g02106(.dina(n2329), .dinb(asqrt[57] ), .dout(n2330));
  jor  g02107(.dina(n2329), .dinb(asqrt[57] ), .dout(n2331));
  jnot g02108(.din(n2118), .dout(n2332));
  jnot g02109(.din(n2119), .dout(n2333));
  jand g02110(.dina(asqrt[44] ), .dinb(n2115), .dout(n2334));
  jand g02111(.dina(n2334), .dinb(n2333), .dout(n2335));
  jor  g02112(.dina(n2335), .dinb(n2332), .dout(n2336));
  jnot g02113(.din(n2120), .dout(n2337));
  jand g02114(.dina(n2334), .dinb(n2337), .dout(n2338));
  jnot g02115(.din(n2338), .dout(n2339));
  jand g02116(.dina(n2339), .dinb(n2336), .dout(n2340));
  jand g02117(.dina(n2340), .dinb(n2331), .dout(n2341));
  jor  g02118(.dina(n2341), .dinb(n2330), .dout(n2342));
  jand g02119(.dina(n2342), .dinb(asqrt[58] ), .dout(n2343));
  jor  g02120(.dina(n2330), .dinb(asqrt[58] ), .dout(n2344));
  jor  g02121(.dina(n2344), .dinb(n2341), .dout(n2345));
  jnot g02122(.din(n2126), .dout(n2346));
  jnot g02123(.din(n2128), .dout(n2347));
  jand g02124(.dina(asqrt[44] ), .dinb(n2122), .dout(n2348));
  jand g02125(.dina(n2348), .dinb(n2347), .dout(n2349));
  jor  g02126(.dina(n2349), .dinb(n2346), .dout(n2350));
  jnot g02127(.din(n2129), .dout(n2351));
  jand g02128(.dina(n2348), .dinb(n2351), .dout(n2352));
  jnot g02129(.din(n2352), .dout(n2353));
  jand g02130(.dina(n2353), .dinb(n2350), .dout(n2354));
  jand g02131(.dina(n2354), .dinb(n2345), .dout(n2355));
  jor  g02132(.dina(n2355), .dinb(n2343), .dout(n2356));
  jand g02133(.dina(n2356), .dinb(asqrt[59] ), .dout(n2357));
  jxor g02134(.dina(n2130), .dinb(n425), .dout(n2358));
  jand g02135(.dina(n2358), .dinb(asqrt[44] ), .dout(n2359));
  jxor g02136(.dina(n2359), .dinb(n2140), .dout(n2360));
  jnot g02137(.din(n2360), .dout(n2361));
  jor  g02138(.dina(n2356), .dinb(asqrt[59] ), .dout(n2362));
  jand g02139(.dina(n2362), .dinb(n2361), .dout(n2363));
  jor  g02140(.dina(n2363), .dinb(n2357), .dout(n2364));
  jand g02141(.dina(n2364), .dinb(asqrt[60] ), .dout(n2365));
  jnot g02142(.din(n2145), .dout(n2366));
  jand g02143(.dina(n2366), .dinb(n2143), .dout(n2367));
  jand g02144(.dina(n2367), .dinb(asqrt[44] ), .dout(n2368));
  jxor g02145(.dina(n2368), .dinb(n2153), .dout(n2369));
  jnot g02146(.din(n2369), .dout(n2370));
  jor  g02147(.dina(n2357), .dinb(asqrt[60] ), .dout(n2371));
  jor  g02148(.dina(n2371), .dinb(n2363), .dout(n2372));
  jand g02149(.dina(n2372), .dinb(n2370), .dout(n2373));
  jor  g02150(.dina(n2373), .dinb(n2365), .dout(n2374));
  jand g02151(.dina(n2374), .dinb(asqrt[61] ), .dout(n2375));
  jor  g02152(.dina(n2374), .dinb(asqrt[61] ), .dout(n2376));
  jnot g02153(.din(n2159), .dout(n2377));
  jnot g02154(.din(n2160), .dout(n2378));
  jand g02155(.dina(asqrt[44] ), .dinb(n2156), .dout(n2379));
  jand g02156(.dina(n2379), .dinb(n2378), .dout(n2380));
  jor  g02157(.dina(n2380), .dinb(n2377), .dout(n2381));
  jnot g02158(.din(n2161), .dout(n2382));
  jand g02159(.dina(n2379), .dinb(n2382), .dout(n2383));
  jnot g02160(.din(n2383), .dout(n2384));
  jand g02161(.dina(n2384), .dinb(n2381), .dout(n2385));
  jand g02162(.dina(n2385), .dinb(n2376), .dout(n2386));
  jor  g02163(.dina(n2386), .dinb(n2375), .dout(n2387));
  jand g02164(.dina(n2387), .dinb(asqrt[62] ), .dout(n2388));
  jor  g02165(.dina(n2375), .dinb(asqrt[62] ), .dout(n2389));
  jor  g02166(.dina(n2389), .dinb(n2386), .dout(n2390));
  jnot g02167(.din(n2167), .dout(n2391));
  jnot g02168(.din(n2169), .dout(n2392));
  jand g02169(.dina(asqrt[44] ), .dinb(n2163), .dout(n2393));
  jand g02170(.dina(n2393), .dinb(n2392), .dout(n2394));
  jor  g02171(.dina(n2394), .dinb(n2391), .dout(n2395));
  jnot g02172(.din(n2170), .dout(n2396));
  jand g02173(.dina(n2393), .dinb(n2396), .dout(n2397));
  jnot g02174(.din(n2397), .dout(n2398));
  jand g02175(.dina(n2398), .dinb(n2395), .dout(n2399));
  jand g02176(.dina(n2399), .dinb(n2390), .dout(n2400));
  jor  g02177(.dina(n2400), .dinb(n2388), .dout(n2401));
  jxor g02178(.dina(n2171), .dinb(n199), .dout(n2402));
  jand g02179(.dina(n2402), .dinb(asqrt[44] ), .dout(n2403));
  jxor g02180(.dina(n2403), .dinb(n2181), .dout(n2404));
  jnot g02181(.din(n2183), .dout(n2405));
  jand g02182(.dina(asqrt[44] ), .dinb(n2190), .dout(n2406));
  jand g02183(.dina(n2406), .dinb(n2405), .dout(n2407));
  jor  g02184(.dina(n2407), .dinb(n2198), .dout(n2408));
  jor  g02185(.dina(n2408), .dinb(n2404), .dout(n2409));
  jnot g02186(.din(n2409), .dout(n2410));
  jand g02187(.dina(n2410), .dinb(n2401), .dout(n2411));
  jor  g02188(.dina(n2411), .dinb(asqrt[63] ), .dout(n2412));
  jnot g02189(.din(n2404), .dout(n2413));
  jor  g02190(.dina(n2413), .dinb(n2401), .dout(n2414));
  jor  g02191(.dina(n2406), .dinb(n2405), .dout(n2415));
  jand g02192(.dina(n2190), .dinb(n2405), .dout(n2416));
  jor  g02193(.dina(n2416), .dinb(n194), .dout(n2417));
  jnot g02194(.din(n2417), .dout(n2418));
  jand g02195(.dina(n2418), .dinb(n2415), .dout(n2419));
  jnot g02196(.din(asqrt[44] ), .dout(n2420));
  jnot g02197(.din(n2419), .dout(n2423));
  jand g02198(.dina(n2423), .dinb(n2414), .dout(n2424));
  jand g02199(.dina(n2424), .dinb(n2412), .dout(n2425));
  jnot g02200(.din(n2425), .dout(asqrt[43] ));
  jor  g02201(.dina(n2425), .dinb(n2209), .dout(n2427));
  jnot g02202(.din(a[84] ), .dout(n2428));
  jnot g02203(.din(a[85] ), .dout(n2429));
  jand g02204(.dina(n2209), .dinb(n2429), .dout(n2430));
  jand g02205(.dina(n2430), .dinb(n2428), .dout(n2431));
  jnot g02206(.din(n2431), .dout(n2432));
  jand g02207(.dina(n2432), .dinb(n2427), .dout(n2433));
  jor  g02208(.dina(n2433), .dinb(n2420), .dout(n2434));
  jor  g02209(.dina(n2425), .dinb(a[86] ), .dout(n2435));
  jxor g02210(.dina(n2435), .dinb(n2210), .dout(n2436));
  jand g02211(.dina(n2433), .dinb(n2420), .dout(n2437));
  jor  g02212(.dina(n2437), .dinb(n2436), .dout(n2438));
  jand g02213(.dina(n2438), .dinb(n2434), .dout(n2439));
  jor  g02214(.dina(n2439), .dinb(n2010), .dout(n2440));
  jand g02215(.dina(n2434), .dinb(n2010), .dout(n2441));
  jand g02216(.dina(n2441), .dinb(n2438), .dout(n2442));
  jor  g02217(.dina(n2435), .dinb(a[87] ), .dout(n2443));
  jnot g02218(.din(n2412), .dout(n2444));
  jnot g02219(.din(n2414), .dout(n2445));
  jor  g02220(.dina(n2419), .dinb(n2420), .dout(n2446));
  jor  g02221(.dina(n2446), .dinb(n2445), .dout(n2447));
  jor  g02222(.dina(n2447), .dinb(n2444), .dout(n2448));
  jand g02223(.dina(n2448), .dinb(n2443), .dout(n2449));
  jxor g02224(.dina(n2449), .dinb(n2013), .dout(n2450));
  jor  g02225(.dina(n2450), .dinb(n2442), .dout(n2451));
  jand g02226(.dina(n2451), .dinb(n2440), .dout(n2452));
  jor  g02227(.dina(n2452), .dinb(n2005), .dout(n2453));
  jand g02228(.dina(n2452), .dinb(n2005), .dout(n2454));
  jxor g02229(.dina(n2213), .dinb(n2010), .dout(n2455));
  jor  g02230(.dina(n2455), .dinb(n2425), .dout(n2456));
  jxor g02231(.dina(n2456), .dinb(n2216), .dout(n2457));
  jor  g02232(.dina(n2457), .dinb(n2454), .dout(n2458));
  jand g02233(.dina(n2458), .dinb(n2453), .dout(n2459));
  jor  g02234(.dina(n2459), .dinb(n1646), .dout(n2460));
  jnot g02235(.din(n2222), .dout(n2461));
  jor  g02236(.dina(n2461), .dinb(n2220), .dout(n2462));
  jor  g02237(.dina(n2462), .dinb(n2425), .dout(n2463));
  jxor g02238(.dina(n2463), .dinb(n2231), .dout(n2464));
  jand g02239(.dina(n2453), .dinb(n1646), .dout(n2465));
  jand g02240(.dina(n2465), .dinb(n2458), .dout(n2466));
  jor  g02241(.dina(n2466), .dinb(n2464), .dout(n2467));
  jand g02242(.dina(n2467), .dinb(n2460), .dout(n2468));
  jor  g02243(.dina(n2468), .dinb(n1641), .dout(n2469));
  jand g02244(.dina(n2468), .dinb(n1641), .dout(n2470));
  jxor g02245(.dina(n2233), .dinb(n1646), .dout(n2471));
  jor  g02246(.dina(n2471), .dinb(n2425), .dout(n2472));
  jxor g02247(.dina(n2472), .dinb(n2238), .dout(n2473));
  jnot g02248(.din(n2473), .dout(n2474));
  jor  g02249(.dina(n2474), .dinb(n2470), .dout(n2475));
  jand g02250(.dina(n2475), .dinb(n2469), .dout(n2476));
  jor  g02251(.dina(n2476), .dinb(n1317), .dout(n2477));
  jand g02252(.dina(n2469), .dinb(n1317), .dout(n2478));
  jand g02253(.dina(n2478), .dinb(n2475), .dout(n2479));
  jnot g02254(.din(n2242), .dout(n2480));
  jand g02255(.dina(asqrt[43] ), .dinb(n2480), .dout(n2481));
  jand g02256(.dina(n2481), .dinb(n2249), .dout(n2482));
  jor  g02257(.dina(n2482), .dinb(n2247), .dout(n2483));
  jand g02258(.dina(n2481), .dinb(n2250), .dout(n2484));
  jnot g02259(.din(n2484), .dout(n2485));
  jand g02260(.dina(n2485), .dinb(n2483), .dout(n2486));
  jnot g02261(.din(n2486), .dout(n2487));
  jor  g02262(.dina(n2487), .dinb(n2479), .dout(n2488));
  jand g02263(.dina(n2488), .dinb(n2477), .dout(n2489));
  jor  g02264(.dina(n2489), .dinb(n1312), .dout(n2490));
  jand g02265(.dina(n2489), .dinb(n1312), .dout(n2491));
  jnot g02266(.din(n2257), .dout(n2492));
  jxor g02267(.dina(n2251), .dinb(n1317), .dout(n2493));
  jor  g02268(.dina(n2493), .dinb(n2425), .dout(n2494));
  jxor g02269(.dina(n2494), .dinb(n2492), .dout(n2495));
  jnot g02270(.din(n2495), .dout(n2496));
  jor  g02271(.dina(n2496), .dinb(n2491), .dout(n2497));
  jand g02272(.dina(n2497), .dinb(n2490), .dout(n2498));
  jor  g02273(.dina(n2498), .dinb(n1039), .dout(n2499));
  jnot g02274(.din(n2262), .dout(n2500));
  jor  g02275(.dina(n2500), .dinb(n2260), .dout(n2501));
  jor  g02276(.dina(n2501), .dinb(n2425), .dout(n2502));
  jxor g02277(.dina(n2502), .dinb(n2271), .dout(n2503));
  jand g02278(.dina(n2490), .dinb(n1039), .dout(n2504));
  jand g02279(.dina(n2504), .dinb(n2497), .dout(n2505));
  jor  g02280(.dina(n2505), .dinb(n2503), .dout(n2506));
  jand g02281(.dina(n2506), .dinb(n2499), .dout(n2507));
  jor  g02282(.dina(n2507), .dinb(n1034), .dout(n2508));
  jand g02283(.dina(n2507), .dinb(n1034), .dout(n2509));
  jnot g02284(.din(n2278), .dout(n2510));
  jxor g02285(.dina(n2273), .dinb(n1039), .dout(n2511));
  jor  g02286(.dina(n2511), .dinb(n2425), .dout(n2512));
  jxor g02287(.dina(n2512), .dinb(n2510), .dout(n2513));
  jnot g02288(.din(n2513), .dout(n2514));
  jor  g02289(.dina(n2514), .dinb(n2509), .dout(n2515));
  jand g02290(.dina(n2515), .dinb(n2508), .dout(n2516));
  jor  g02291(.dina(n2516), .dinb(n796), .dout(n2517));
  jand g02292(.dina(n2508), .dinb(n796), .dout(n2518));
  jand g02293(.dina(n2518), .dinb(n2515), .dout(n2519));
  jnot g02294(.din(n2281), .dout(n2520));
  jand g02295(.dina(asqrt[43] ), .dinb(n2520), .dout(n2521));
  jand g02296(.dina(n2521), .dinb(n2288), .dout(n2522));
  jor  g02297(.dina(n2522), .dinb(n2286), .dout(n2523));
  jand g02298(.dina(n2521), .dinb(n2289), .dout(n2524));
  jnot g02299(.din(n2524), .dout(n2525));
  jand g02300(.dina(n2525), .dinb(n2523), .dout(n2526));
  jnot g02301(.din(n2526), .dout(n2527));
  jor  g02302(.dina(n2527), .dinb(n2519), .dout(n2528));
  jand g02303(.dina(n2528), .dinb(n2517), .dout(n2529));
  jor  g02304(.dina(n2529), .dinb(n791), .dout(n2530));
  jxor g02305(.dina(n2290), .dinb(n796), .dout(n2531));
  jor  g02306(.dina(n2531), .dinb(n2425), .dout(n2532));
  jxor g02307(.dina(n2532), .dinb(n2295), .dout(n2533));
  jand g02308(.dina(n2529), .dinb(n791), .dout(n2534));
  jor  g02309(.dina(n2534), .dinb(n2533), .dout(n2535));
  jand g02310(.dina(n2535), .dinb(n2530), .dout(n2536));
  jor  g02311(.dina(n2536), .dinb(n595), .dout(n2537));
  jnot g02312(.din(n2300), .dout(n2538));
  jor  g02313(.dina(n2538), .dinb(n2298), .dout(n2539));
  jor  g02314(.dina(n2539), .dinb(n2425), .dout(n2540));
  jxor g02315(.dina(n2540), .dinb(n2309), .dout(n2541));
  jand g02316(.dina(n2530), .dinb(n595), .dout(n2542));
  jand g02317(.dina(n2542), .dinb(n2535), .dout(n2543));
  jor  g02318(.dina(n2543), .dinb(n2541), .dout(n2544));
  jand g02319(.dina(n2544), .dinb(n2537), .dout(n2545));
  jor  g02320(.dina(n2545), .dinb(n590), .dout(n2546));
  jand g02321(.dina(n2545), .dinb(n590), .dout(n2547));
  jnot g02322(.din(n2312), .dout(n2548));
  jand g02323(.dina(asqrt[43] ), .dinb(n2548), .dout(n2549));
  jand g02324(.dina(n2549), .dinb(n2317), .dout(n2550));
  jor  g02325(.dina(n2550), .dinb(n2316), .dout(n2551));
  jand g02326(.dina(n2549), .dinb(n2318), .dout(n2552));
  jnot g02327(.din(n2552), .dout(n2553));
  jand g02328(.dina(n2553), .dinb(n2551), .dout(n2554));
  jnot g02329(.din(n2554), .dout(n2555));
  jor  g02330(.dina(n2555), .dinb(n2547), .dout(n2556));
  jand g02331(.dina(n2556), .dinb(n2546), .dout(n2557));
  jor  g02332(.dina(n2557), .dinb(n430), .dout(n2558));
  jand g02333(.dina(n2546), .dinb(n430), .dout(n2559));
  jand g02334(.dina(n2559), .dinb(n2556), .dout(n2560));
  jnot g02335(.din(n2320), .dout(n2561));
  jand g02336(.dina(asqrt[43] ), .dinb(n2561), .dout(n2562));
  jand g02337(.dina(n2562), .dinb(n2327), .dout(n2563));
  jor  g02338(.dina(n2563), .dinb(n2325), .dout(n2564));
  jand g02339(.dina(n2562), .dinb(n2328), .dout(n2565));
  jnot g02340(.din(n2565), .dout(n2566));
  jand g02341(.dina(n2566), .dinb(n2564), .dout(n2567));
  jnot g02342(.din(n2567), .dout(n2568));
  jor  g02343(.dina(n2568), .dinb(n2560), .dout(n2569));
  jand g02344(.dina(n2569), .dinb(n2558), .dout(n2570));
  jor  g02345(.dina(n2570), .dinb(n425), .dout(n2571));
  jxor g02346(.dina(n2329), .dinb(n430), .dout(n2572));
  jor  g02347(.dina(n2572), .dinb(n2425), .dout(n2573));
  jxor g02348(.dina(n2573), .dinb(n2340), .dout(n2574));
  jand g02349(.dina(n2570), .dinb(n425), .dout(n2575));
  jor  g02350(.dina(n2575), .dinb(n2574), .dout(n2576));
  jand g02351(.dina(n2576), .dinb(n2571), .dout(n2577));
  jor  g02352(.dina(n2577), .dinb(n305), .dout(n2578));
  jnot g02353(.din(n2345), .dout(n2579));
  jor  g02354(.dina(n2579), .dinb(n2343), .dout(n2580));
  jor  g02355(.dina(n2580), .dinb(n2425), .dout(n2581));
  jxor g02356(.dina(n2581), .dinb(n2354), .dout(n2582));
  jand g02357(.dina(n2571), .dinb(n305), .dout(n2583));
  jand g02358(.dina(n2583), .dinb(n2576), .dout(n2584));
  jor  g02359(.dina(n2584), .dinb(n2582), .dout(n2585));
  jand g02360(.dina(n2585), .dinb(n2578), .dout(n2586));
  jor  g02361(.dina(n2586), .dinb(n290), .dout(n2587));
  jand g02362(.dina(n2586), .dinb(n290), .dout(n2588));
  jnot g02363(.din(n2357), .dout(n2589));
  jand g02364(.dina(asqrt[43] ), .dinb(n2589), .dout(n2590));
  jand g02365(.dina(n2590), .dinb(n2362), .dout(n2591));
  jor  g02366(.dina(n2591), .dinb(n2361), .dout(n2592));
  jand g02367(.dina(n2590), .dinb(n2363), .dout(n2593));
  jnot g02368(.din(n2593), .dout(n2594));
  jand g02369(.dina(n2594), .dinb(n2592), .dout(n2595));
  jnot g02370(.din(n2595), .dout(n2596));
  jor  g02371(.dina(n2596), .dinb(n2588), .dout(n2597));
  jand g02372(.dina(n2597), .dinb(n2587), .dout(n2598));
  jor  g02373(.dina(n2598), .dinb(n223), .dout(n2599));
  jand g02374(.dina(n2587), .dinb(n223), .dout(n2600));
  jand g02375(.dina(n2600), .dinb(n2597), .dout(n2601));
  jnot g02376(.din(n2365), .dout(n2602));
  jand g02377(.dina(asqrt[43] ), .dinb(n2602), .dout(n2603));
  jand g02378(.dina(n2603), .dinb(n2372), .dout(n2604));
  jor  g02379(.dina(n2604), .dinb(n2370), .dout(n2605));
  jand g02380(.dina(n2603), .dinb(n2373), .dout(n2606));
  jnot g02381(.din(n2606), .dout(n2607));
  jand g02382(.dina(n2607), .dinb(n2605), .dout(n2608));
  jnot g02383(.din(n2608), .dout(n2609));
  jor  g02384(.dina(n2609), .dinb(n2601), .dout(n2610));
  jand g02385(.dina(n2610), .dinb(n2599), .dout(n2611));
  jor  g02386(.dina(n2611), .dinb(n199), .dout(n2612));
  jand g02387(.dina(n2611), .dinb(n199), .dout(n2613));
  jxor g02388(.dina(n2374), .dinb(n223), .dout(n2614));
  jor  g02389(.dina(n2614), .dinb(n2425), .dout(n2615));
  jxor g02390(.dina(n2615), .dinb(n2385), .dout(n2616));
  jor  g02391(.dina(n2616), .dinb(n2613), .dout(n2617));
  jand g02392(.dina(n2617), .dinb(n2612), .dout(n2618));
  jnot g02393(.din(n2390), .dout(n2619));
  jor  g02394(.dina(n2619), .dinb(n2388), .dout(n2620));
  jor  g02395(.dina(n2620), .dinb(n2425), .dout(n2621));
  jxor g02396(.dina(n2621), .dinb(n2399), .dout(n2622));
  jand g02397(.dina(asqrt[43] ), .dinb(n2413), .dout(n2623));
  jand g02398(.dina(n2623), .dinb(n2401), .dout(n2624));
  jor  g02399(.dina(n2624), .dinb(n2445), .dout(n2625));
  jor  g02400(.dina(n2625), .dinb(n2622), .dout(n2626));
  jor  g02401(.dina(n2626), .dinb(n2618), .dout(n2627));
  jand g02402(.dina(n2627), .dinb(n194), .dout(n2628));
  jand g02403(.dina(n2622), .dinb(n2618), .dout(n2629));
  jor  g02404(.dina(n2623), .dinb(n2401), .dout(n2630));
  jand g02405(.dina(n2413), .dinb(n2401), .dout(n2631));
  jor  g02406(.dina(n2631), .dinb(n194), .dout(n2632));
  jnot g02407(.din(n2632), .dout(n2633));
  jand g02408(.dina(n2633), .dinb(n2630), .dout(n2634));
  jor  g02409(.dina(n2634), .dinb(n2629), .dout(n2637));
  jor  g02410(.dina(n2637), .dinb(n2628), .dout(asqrt[42] ));
  jand g02411(.dina(asqrt[42] ), .dinb(a[84] ), .dout(n2639));
  jnot g02412(.din(a[82] ), .dout(n2640));
  jnot g02413(.din(a[83] ), .dout(n2641));
  jand g02414(.dina(n2428), .dinb(n2641), .dout(n2642));
  jand g02415(.dina(n2642), .dinb(n2640), .dout(n2643));
  jor  g02416(.dina(n2643), .dinb(n2639), .dout(n2644));
  jand g02417(.dina(n2644), .dinb(asqrt[43] ), .dout(n2645));
  jand g02418(.dina(asqrt[42] ), .dinb(n2428), .dout(n2646));
  jxor g02419(.dina(n2646), .dinb(n2429), .dout(n2647));
  jor  g02420(.dina(n2644), .dinb(asqrt[43] ), .dout(n2648));
  jand g02421(.dina(n2648), .dinb(n2647), .dout(n2649));
  jor  g02422(.dina(n2649), .dinb(n2645), .dout(n2650));
  jand g02423(.dina(n2650), .dinb(asqrt[44] ), .dout(n2651));
  jor  g02424(.dina(n2645), .dinb(asqrt[44] ), .dout(n2652));
  jor  g02425(.dina(n2652), .dinb(n2649), .dout(n2653));
  jand g02426(.dina(n2646), .dinb(n2429), .dout(n2654));
  jnot g02427(.din(n2628), .dout(n2655));
  jnot g02428(.din(n2629), .dout(n2656));
  jnot g02429(.din(n2634), .dout(n2657));
  jand g02430(.dina(n2657), .dinb(asqrt[43] ), .dout(n2658));
  jand g02431(.dina(n2658), .dinb(n2656), .dout(n2659));
  jand g02432(.dina(n2659), .dinb(n2655), .dout(n2660));
  jor  g02433(.dina(n2660), .dinb(n2654), .dout(n2661));
  jxor g02434(.dina(n2661), .dinb(n2209), .dout(n2662));
  jand g02435(.dina(n2662), .dinb(n2653), .dout(n2663));
  jor  g02436(.dina(n2663), .dinb(n2651), .dout(n2664));
  jand g02437(.dina(n2664), .dinb(asqrt[45] ), .dout(n2665));
  jor  g02438(.dina(n2664), .dinb(asqrt[45] ), .dout(n2666));
  jxor g02439(.dina(n2433), .dinb(n2420), .dout(n2667));
  jand g02440(.dina(n2667), .dinb(asqrt[42] ), .dout(n2668));
  jxor g02441(.dina(n2668), .dinb(n2436), .dout(n2669));
  jnot g02442(.din(n2669), .dout(n2670));
  jand g02443(.dina(n2670), .dinb(n2666), .dout(n2671));
  jor  g02444(.dina(n2671), .dinb(n2665), .dout(n2672));
  jand g02445(.dina(n2672), .dinb(asqrt[46] ), .dout(n2673));
  jnot g02446(.din(n2442), .dout(n2674));
  jand g02447(.dina(n2674), .dinb(n2440), .dout(n2675));
  jand g02448(.dina(n2675), .dinb(asqrt[42] ), .dout(n2676));
  jxor g02449(.dina(n2676), .dinb(n2450), .dout(n2677));
  jnot g02450(.din(n2677), .dout(n2678));
  jor  g02451(.dina(n2665), .dinb(asqrt[46] ), .dout(n2679));
  jor  g02452(.dina(n2679), .dinb(n2671), .dout(n2680));
  jand g02453(.dina(n2680), .dinb(n2678), .dout(n2681));
  jor  g02454(.dina(n2681), .dinb(n2673), .dout(n2682));
  jand g02455(.dina(n2682), .dinb(asqrt[47] ), .dout(n2683));
  jor  g02456(.dina(n2682), .dinb(asqrt[47] ), .dout(n2684));
  jnot g02457(.din(n2457), .dout(n2685));
  jxor g02458(.dina(n2452), .dinb(n2005), .dout(n2686));
  jand g02459(.dina(n2686), .dinb(asqrt[42] ), .dout(n2687));
  jxor g02460(.dina(n2687), .dinb(n2685), .dout(n2688));
  jand g02461(.dina(n2688), .dinb(n2684), .dout(n2689));
  jor  g02462(.dina(n2689), .dinb(n2683), .dout(n2690));
  jand g02463(.dina(n2690), .dinb(asqrt[48] ), .dout(n2691));
  jor  g02464(.dina(n2683), .dinb(asqrt[48] ), .dout(n2692));
  jor  g02465(.dina(n2692), .dinb(n2689), .dout(n2693));
  jnot g02466(.din(n2464), .dout(n2694));
  jnot g02467(.din(n2466), .dout(n2695));
  jand g02468(.dina(asqrt[42] ), .dinb(n2460), .dout(n2696));
  jand g02469(.dina(n2696), .dinb(n2695), .dout(n2697));
  jor  g02470(.dina(n2697), .dinb(n2694), .dout(n2698));
  jnot g02471(.din(n2467), .dout(n2699));
  jand g02472(.dina(n2696), .dinb(n2699), .dout(n2700));
  jnot g02473(.din(n2700), .dout(n2701));
  jand g02474(.dina(n2701), .dinb(n2698), .dout(n2702));
  jand g02475(.dina(n2702), .dinb(n2693), .dout(n2703));
  jor  g02476(.dina(n2703), .dinb(n2691), .dout(n2704));
  jand g02477(.dina(n2704), .dinb(asqrt[49] ), .dout(n2705));
  jor  g02478(.dina(n2704), .dinb(asqrt[49] ), .dout(n2706));
  jxor g02479(.dina(n2468), .dinb(n1641), .dout(n2707));
  jand g02480(.dina(n2707), .dinb(asqrt[42] ), .dout(n2708));
  jxor g02481(.dina(n2708), .dinb(n2473), .dout(n2709));
  jand g02482(.dina(n2709), .dinb(n2706), .dout(n2710));
  jor  g02483(.dina(n2710), .dinb(n2705), .dout(n2711));
  jand g02484(.dina(n2711), .dinb(asqrt[50] ), .dout(n2712));
  jnot g02485(.din(n2479), .dout(n2713));
  jand g02486(.dina(n2713), .dinb(n2477), .dout(n2714));
  jand g02487(.dina(n2714), .dinb(asqrt[42] ), .dout(n2715));
  jxor g02488(.dina(n2715), .dinb(n2487), .dout(n2716));
  jnot g02489(.din(n2716), .dout(n2717));
  jor  g02490(.dina(n2705), .dinb(asqrt[50] ), .dout(n2718));
  jor  g02491(.dina(n2718), .dinb(n2710), .dout(n2719));
  jand g02492(.dina(n2719), .dinb(n2717), .dout(n2720));
  jor  g02493(.dina(n2720), .dinb(n2712), .dout(n2721));
  jand g02494(.dina(n2721), .dinb(asqrt[51] ), .dout(n2722));
  jor  g02495(.dina(n2721), .dinb(asqrt[51] ), .dout(n2723));
  jxor g02496(.dina(n2489), .dinb(n1312), .dout(n2724));
  jand g02497(.dina(n2724), .dinb(asqrt[42] ), .dout(n2725));
  jxor g02498(.dina(n2725), .dinb(n2495), .dout(n2726));
  jand g02499(.dina(n2726), .dinb(n2723), .dout(n2727));
  jor  g02500(.dina(n2727), .dinb(n2722), .dout(n2728));
  jand g02501(.dina(n2728), .dinb(asqrt[52] ), .dout(n2729));
  jor  g02502(.dina(n2722), .dinb(asqrt[52] ), .dout(n2730));
  jor  g02503(.dina(n2730), .dinb(n2727), .dout(n2731));
  jnot g02504(.din(n2503), .dout(n2732));
  jnot g02505(.din(n2505), .dout(n2733));
  jand g02506(.dina(asqrt[42] ), .dinb(n2499), .dout(n2734));
  jand g02507(.dina(n2734), .dinb(n2733), .dout(n2735));
  jor  g02508(.dina(n2735), .dinb(n2732), .dout(n2736));
  jnot g02509(.din(n2506), .dout(n2737));
  jand g02510(.dina(n2734), .dinb(n2737), .dout(n2738));
  jnot g02511(.din(n2738), .dout(n2739));
  jand g02512(.dina(n2739), .dinb(n2736), .dout(n2740));
  jand g02513(.dina(n2740), .dinb(n2731), .dout(n2741));
  jor  g02514(.dina(n2741), .dinb(n2729), .dout(n2742));
  jand g02515(.dina(n2742), .dinb(asqrt[53] ), .dout(n2743));
  jxor g02516(.dina(n2507), .dinb(n1034), .dout(n2744));
  jand g02517(.dina(n2744), .dinb(asqrt[42] ), .dout(n2745));
  jxor g02518(.dina(n2745), .dinb(n2514), .dout(n2746));
  jnot g02519(.din(n2746), .dout(n2747));
  jor  g02520(.dina(n2742), .dinb(asqrt[53] ), .dout(n2748));
  jand g02521(.dina(n2748), .dinb(n2747), .dout(n2749));
  jor  g02522(.dina(n2749), .dinb(n2743), .dout(n2750));
  jand g02523(.dina(n2750), .dinb(asqrt[54] ), .dout(n2751));
  jnot g02524(.din(n2519), .dout(n2752));
  jand g02525(.dina(n2752), .dinb(n2517), .dout(n2753));
  jand g02526(.dina(n2753), .dinb(asqrt[42] ), .dout(n2754));
  jxor g02527(.dina(n2754), .dinb(n2527), .dout(n2755));
  jnot g02528(.din(n2755), .dout(n2756));
  jor  g02529(.dina(n2743), .dinb(asqrt[54] ), .dout(n2757));
  jor  g02530(.dina(n2757), .dinb(n2749), .dout(n2758));
  jand g02531(.dina(n2758), .dinb(n2756), .dout(n2759));
  jor  g02532(.dina(n2759), .dinb(n2751), .dout(n2760));
  jand g02533(.dina(n2760), .dinb(asqrt[55] ), .dout(n2761));
  jor  g02534(.dina(n2760), .dinb(asqrt[55] ), .dout(n2762));
  jnot g02535(.din(n2533), .dout(n2763));
  jnot g02536(.din(n2534), .dout(n2764));
  jand g02537(.dina(asqrt[42] ), .dinb(n2530), .dout(n2765));
  jand g02538(.dina(n2765), .dinb(n2764), .dout(n2766));
  jor  g02539(.dina(n2766), .dinb(n2763), .dout(n2767));
  jnot g02540(.din(n2535), .dout(n2768));
  jand g02541(.dina(n2765), .dinb(n2768), .dout(n2769));
  jnot g02542(.din(n2769), .dout(n2770));
  jand g02543(.dina(n2770), .dinb(n2767), .dout(n2771));
  jand g02544(.dina(n2771), .dinb(n2762), .dout(n2772));
  jor  g02545(.dina(n2772), .dinb(n2761), .dout(n2773));
  jand g02546(.dina(n2773), .dinb(asqrt[56] ), .dout(n2774));
  jor  g02547(.dina(n2761), .dinb(asqrt[56] ), .dout(n2775));
  jor  g02548(.dina(n2775), .dinb(n2772), .dout(n2776));
  jnot g02549(.din(n2541), .dout(n2777));
  jnot g02550(.din(n2543), .dout(n2778));
  jand g02551(.dina(asqrt[42] ), .dinb(n2537), .dout(n2779));
  jand g02552(.dina(n2779), .dinb(n2778), .dout(n2780));
  jor  g02553(.dina(n2780), .dinb(n2777), .dout(n2781));
  jnot g02554(.din(n2544), .dout(n2782));
  jand g02555(.dina(n2779), .dinb(n2782), .dout(n2783));
  jnot g02556(.din(n2783), .dout(n2784));
  jand g02557(.dina(n2784), .dinb(n2781), .dout(n2785));
  jand g02558(.dina(n2785), .dinb(n2776), .dout(n2786));
  jor  g02559(.dina(n2786), .dinb(n2774), .dout(n2787));
  jand g02560(.dina(n2787), .dinb(asqrt[57] ), .dout(n2788));
  jxor g02561(.dina(n2545), .dinb(n590), .dout(n2789));
  jand g02562(.dina(n2789), .dinb(asqrt[42] ), .dout(n2790));
  jxor g02563(.dina(n2790), .dinb(n2555), .dout(n2791));
  jnot g02564(.din(n2791), .dout(n2792));
  jor  g02565(.dina(n2787), .dinb(asqrt[57] ), .dout(n2793));
  jand g02566(.dina(n2793), .dinb(n2792), .dout(n2794));
  jor  g02567(.dina(n2794), .dinb(n2788), .dout(n2795));
  jand g02568(.dina(n2795), .dinb(asqrt[58] ), .dout(n2796));
  jnot g02569(.din(n2560), .dout(n2797));
  jand g02570(.dina(n2797), .dinb(n2558), .dout(n2798));
  jand g02571(.dina(n2798), .dinb(asqrt[42] ), .dout(n2799));
  jxor g02572(.dina(n2799), .dinb(n2568), .dout(n2800));
  jnot g02573(.din(n2800), .dout(n2801));
  jor  g02574(.dina(n2788), .dinb(asqrt[58] ), .dout(n2802));
  jor  g02575(.dina(n2802), .dinb(n2794), .dout(n2803));
  jand g02576(.dina(n2803), .dinb(n2801), .dout(n2804));
  jor  g02577(.dina(n2804), .dinb(n2796), .dout(n2805));
  jand g02578(.dina(n2805), .dinb(asqrt[59] ), .dout(n2806));
  jor  g02579(.dina(n2805), .dinb(asqrt[59] ), .dout(n2807));
  jnot g02580(.din(n2574), .dout(n2808));
  jnot g02581(.din(n2575), .dout(n2809));
  jand g02582(.dina(asqrt[42] ), .dinb(n2571), .dout(n2810));
  jand g02583(.dina(n2810), .dinb(n2809), .dout(n2811));
  jor  g02584(.dina(n2811), .dinb(n2808), .dout(n2812));
  jnot g02585(.din(n2576), .dout(n2813));
  jand g02586(.dina(n2810), .dinb(n2813), .dout(n2814));
  jnot g02587(.din(n2814), .dout(n2815));
  jand g02588(.dina(n2815), .dinb(n2812), .dout(n2816));
  jand g02589(.dina(n2816), .dinb(n2807), .dout(n2817));
  jor  g02590(.dina(n2817), .dinb(n2806), .dout(n2818));
  jand g02591(.dina(n2818), .dinb(asqrt[60] ), .dout(n2819));
  jor  g02592(.dina(n2806), .dinb(asqrt[60] ), .dout(n2820));
  jor  g02593(.dina(n2820), .dinb(n2817), .dout(n2821));
  jnot g02594(.din(n2582), .dout(n2822));
  jnot g02595(.din(n2584), .dout(n2823));
  jand g02596(.dina(asqrt[42] ), .dinb(n2578), .dout(n2824));
  jand g02597(.dina(n2824), .dinb(n2823), .dout(n2825));
  jor  g02598(.dina(n2825), .dinb(n2822), .dout(n2826));
  jnot g02599(.din(n2585), .dout(n2827));
  jand g02600(.dina(n2824), .dinb(n2827), .dout(n2828));
  jnot g02601(.din(n2828), .dout(n2829));
  jand g02602(.dina(n2829), .dinb(n2826), .dout(n2830));
  jand g02603(.dina(n2830), .dinb(n2821), .dout(n2831));
  jor  g02604(.dina(n2831), .dinb(n2819), .dout(n2832));
  jand g02605(.dina(n2832), .dinb(asqrt[61] ), .dout(n2833));
  jxor g02606(.dina(n2586), .dinb(n290), .dout(n2834));
  jand g02607(.dina(n2834), .dinb(asqrt[42] ), .dout(n2835));
  jxor g02608(.dina(n2835), .dinb(n2596), .dout(n2836));
  jnot g02609(.din(n2836), .dout(n2837));
  jor  g02610(.dina(n2832), .dinb(asqrt[61] ), .dout(n2838));
  jand g02611(.dina(n2838), .dinb(n2837), .dout(n2839));
  jor  g02612(.dina(n2839), .dinb(n2833), .dout(n2840));
  jand g02613(.dina(n2840), .dinb(asqrt[62] ), .dout(n2841));
  jnot g02614(.din(n2601), .dout(n2842));
  jand g02615(.dina(n2842), .dinb(n2599), .dout(n2843));
  jand g02616(.dina(n2843), .dinb(asqrt[42] ), .dout(n2844));
  jxor g02617(.dina(n2844), .dinb(n2609), .dout(n2845));
  jnot g02618(.din(n2845), .dout(n2846));
  jor  g02619(.dina(n2833), .dinb(asqrt[62] ), .dout(n2847));
  jor  g02620(.dina(n2847), .dinb(n2839), .dout(n2848));
  jand g02621(.dina(n2848), .dinb(n2846), .dout(n2849));
  jor  g02622(.dina(n2849), .dinb(n2841), .dout(n2850));
  jxor g02623(.dina(n2611), .dinb(n199), .dout(n2851));
  jand g02624(.dina(n2851), .dinb(asqrt[42] ), .dout(n2852));
  jxor g02625(.dina(n2852), .dinb(n2616), .dout(n2853));
  jnot g02626(.din(n2618), .dout(n2854));
  jnot g02627(.din(n2622), .dout(n2855));
  jand g02628(.dina(asqrt[42] ), .dinb(n2855), .dout(n2856));
  jand g02629(.dina(n2856), .dinb(n2854), .dout(n2857));
  jor  g02630(.dina(n2857), .dinb(n2629), .dout(n2858));
  jor  g02631(.dina(n2858), .dinb(n2853), .dout(n2859));
  jnot g02632(.din(n2859), .dout(n2860));
  jand g02633(.dina(n2860), .dinb(n2850), .dout(n2861));
  jor  g02634(.dina(n2861), .dinb(asqrt[63] ), .dout(n2862));
  jnot g02635(.din(n2853), .dout(n2863));
  jor  g02636(.dina(n2863), .dinb(n2850), .dout(n2864));
  jor  g02637(.dina(n2856), .dinb(n2854), .dout(n2865));
  jand g02638(.dina(n2855), .dinb(n2854), .dout(n2866));
  jor  g02639(.dina(n2866), .dinb(n194), .dout(n2867));
  jnot g02640(.din(n2867), .dout(n2868));
  jand g02641(.dina(n2868), .dinb(n2865), .dout(n2869));
  jnot g02642(.din(asqrt[42] ), .dout(n2870));
  jnot g02643(.din(n2869), .dout(n2873));
  jand g02644(.dina(n2873), .dinb(n2864), .dout(n2874));
  jand g02645(.dina(n2874), .dinb(n2862), .dout(n2875));
  jnot g02646(.din(n2875), .dout(asqrt[41] ));
  jor  g02647(.dina(n2875), .dinb(n2640), .dout(n2877));
  jnot g02648(.din(a[80] ), .dout(n2878));
  jnot g02649(.din(a[81] ), .dout(n2879));
  jand g02650(.dina(n2640), .dinb(n2879), .dout(n2880));
  jand g02651(.dina(n2880), .dinb(n2878), .dout(n2881));
  jnot g02652(.din(n2881), .dout(n2882));
  jand g02653(.dina(n2882), .dinb(n2877), .dout(n2883));
  jor  g02654(.dina(n2883), .dinb(n2870), .dout(n2884));
  jor  g02655(.dina(n2875), .dinb(a[82] ), .dout(n2885));
  jxor g02656(.dina(n2885), .dinb(n2641), .dout(n2886));
  jand g02657(.dina(n2883), .dinb(n2870), .dout(n2887));
  jor  g02658(.dina(n2887), .dinb(n2886), .dout(n2888));
  jand g02659(.dina(n2888), .dinb(n2884), .dout(n2889));
  jor  g02660(.dina(n2889), .dinb(n2425), .dout(n2890));
  jand g02661(.dina(n2884), .dinb(n2425), .dout(n2891));
  jand g02662(.dina(n2891), .dinb(n2888), .dout(n2892));
  jor  g02663(.dina(n2885), .dinb(a[83] ), .dout(n2893));
  jnot g02664(.din(n2862), .dout(n2894));
  jnot g02665(.din(n2864), .dout(n2895));
  jor  g02666(.dina(n2869), .dinb(n2870), .dout(n2896));
  jor  g02667(.dina(n2896), .dinb(n2895), .dout(n2897));
  jor  g02668(.dina(n2897), .dinb(n2894), .dout(n2898));
  jand g02669(.dina(n2898), .dinb(n2893), .dout(n2899));
  jxor g02670(.dina(n2899), .dinb(n2428), .dout(n2900));
  jor  g02671(.dina(n2900), .dinb(n2892), .dout(n2901));
  jand g02672(.dina(n2901), .dinb(n2890), .dout(n2902));
  jor  g02673(.dina(n2902), .dinb(n2420), .dout(n2903));
  jand g02674(.dina(n2902), .dinb(n2420), .dout(n2904));
  jxor g02675(.dina(n2644), .dinb(n2425), .dout(n2905));
  jor  g02676(.dina(n2905), .dinb(n2875), .dout(n2906));
  jxor g02677(.dina(n2906), .dinb(n2647), .dout(n2907));
  jor  g02678(.dina(n2907), .dinb(n2904), .dout(n2908));
  jand g02679(.dina(n2908), .dinb(n2903), .dout(n2909));
  jor  g02680(.dina(n2909), .dinb(n2010), .dout(n2910));
  jnot g02681(.din(n2653), .dout(n2911));
  jor  g02682(.dina(n2911), .dinb(n2651), .dout(n2912));
  jor  g02683(.dina(n2912), .dinb(n2875), .dout(n2913));
  jxor g02684(.dina(n2913), .dinb(n2662), .dout(n2914));
  jand g02685(.dina(n2903), .dinb(n2010), .dout(n2915));
  jand g02686(.dina(n2915), .dinb(n2908), .dout(n2916));
  jor  g02687(.dina(n2916), .dinb(n2914), .dout(n2917));
  jand g02688(.dina(n2917), .dinb(n2910), .dout(n2918));
  jor  g02689(.dina(n2918), .dinb(n2005), .dout(n2919));
  jand g02690(.dina(n2918), .dinb(n2005), .dout(n2920));
  jxor g02691(.dina(n2664), .dinb(n2010), .dout(n2921));
  jor  g02692(.dina(n2921), .dinb(n2875), .dout(n2922));
  jxor g02693(.dina(n2922), .dinb(n2669), .dout(n2923));
  jnot g02694(.din(n2923), .dout(n2924));
  jor  g02695(.dina(n2924), .dinb(n2920), .dout(n2925));
  jand g02696(.dina(n2925), .dinb(n2919), .dout(n2926));
  jor  g02697(.dina(n2926), .dinb(n1646), .dout(n2927));
  jand g02698(.dina(n2919), .dinb(n1646), .dout(n2928));
  jand g02699(.dina(n2928), .dinb(n2925), .dout(n2929));
  jnot g02700(.din(n2673), .dout(n2930));
  jand g02701(.dina(asqrt[41] ), .dinb(n2930), .dout(n2931));
  jand g02702(.dina(n2931), .dinb(n2680), .dout(n2932));
  jor  g02703(.dina(n2932), .dinb(n2678), .dout(n2933));
  jand g02704(.dina(n2931), .dinb(n2681), .dout(n2934));
  jnot g02705(.din(n2934), .dout(n2935));
  jand g02706(.dina(n2935), .dinb(n2933), .dout(n2936));
  jnot g02707(.din(n2936), .dout(n2937));
  jor  g02708(.dina(n2937), .dinb(n2929), .dout(n2938));
  jand g02709(.dina(n2938), .dinb(n2927), .dout(n2939));
  jor  g02710(.dina(n2939), .dinb(n1641), .dout(n2940));
  jand g02711(.dina(n2939), .dinb(n1641), .dout(n2941));
  jnot g02712(.din(n2688), .dout(n2942));
  jxor g02713(.dina(n2682), .dinb(n1646), .dout(n2943));
  jor  g02714(.dina(n2943), .dinb(n2875), .dout(n2944));
  jxor g02715(.dina(n2944), .dinb(n2942), .dout(n2945));
  jnot g02716(.din(n2945), .dout(n2946));
  jor  g02717(.dina(n2946), .dinb(n2941), .dout(n2947));
  jand g02718(.dina(n2947), .dinb(n2940), .dout(n2948));
  jor  g02719(.dina(n2948), .dinb(n1317), .dout(n2949));
  jnot g02720(.din(n2693), .dout(n2950));
  jor  g02721(.dina(n2950), .dinb(n2691), .dout(n2951));
  jor  g02722(.dina(n2951), .dinb(n2875), .dout(n2952));
  jxor g02723(.dina(n2952), .dinb(n2702), .dout(n2953));
  jand g02724(.dina(n2940), .dinb(n1317), .dout(n2954));
  jand g02725(.dina(n2954), .dinb(n2947), .dout(n2955));
  jor  g02726(.dina(n2955), .dinb(n2953), .dout(n2956));
  jand g02727(.dina(n2956), .dinb(n2949), .dout(n2957));
  jor  g02728(.dina(n2957), .dinb(n1312), .dout(n2958));
  jand g02729(.dina(n2957), .dinb(n1312), .dout(n2959));
  jnot g02730(.din(n2709), .dout(n2960));
  jxor g02731(.dina(n2704), .dinb(n1317), .dout(n2961));
  jor  g02732(.dina(n2961), .dinb(n2875), .dout(n2962));
  jxor g02733(.dina(n2962), .dinb(n2960), .dout(n2963));
  jnot g02734(.din(n2963), .dout(n2964));
  jor  g02735(.dina(n2964), .dinb(n2959), .dout(n2965));
  jand g02736(.dina(n2965), .dinb(n2958), .dout(n2966));
  jor  g02737(.dina(n2966), .dinb(n1039), .dout(n2967));
  jand g02738(.dina(n2958), .dinb(n1039), .dout(n2968));
  jand g02739(.dina(n2968), .dinb(n2965), .dout(n2969));
  jnot g02740(.din(n2712), .dout(n2970));
  jand g02741(.dina(asqrt[41] ), .dinb(n2970), .dout(n2971));
  jand g02742(.dina(n2971), .dinb(n2719), .dout(n2972));
  jor  g02743(.dina(n2972), .dinb(n2717), .dout(n2973));
  jand g02744(.dina(n2971), .dinb(n2720), .dout(n2974));
  jnot g02745(.din(n2974), .dout(n2975));
  jand g02746(.dina(n2975), .dinb(n2973), .dout(n2976));
  jnot g02747(.din(n2976), .dout(n2977));
  jor  g02748(.dina(n2977), .dinb(n2969), .dout(n2978));
  jand g02749(.dina(n2978), .dinb(n2967), .dout(n2979));
  jor  g02750(.dina(n2979), .dinb(n1034), .dout(n2980));
  jxor g02751(.dina(n2721), .dinb(n1039), .dout(n2981));
  jor  g02752(.dina(n2981), .dinb(n2875), .dout(n2982));
  jxor g02753(.dina(n2982), .dinb(n2726), .dout(n2983));
  jand g02754(.dina(n2979), .dinb(n1034), .dout(n2984));
  jor  g02755(.dina(n2984), .dinb(n2983), .dout(n2985));
  jand g02756(.dina(n2985), .dinb(n2980), .dout(n2986));
  jor  g02757(.dina(n2986), .dinb(n796), .dout(n2987));
  jnot g02758(.din(n2731), .dout(n2988));
  jor  g02759(.dina(n2988), .dinb(n2729), .dout(n2989));
  jor  g02760(.dina(n2989), .dinb(n2875), .dout(n2990));
  jxor g02761(.dina(n2990), .dinb(n2740), .dout(n2991));
  jand g02762(.dina(n2980), .dinb(n796), .dout(n2992));
  jand g02763(.dina(n2992), .dinb(n2985), .dout(n2993));
  jor  g02764(.dina(n2993), .dinb(n2991), .dout(n2994));
  jand g02765(.dina(n2994), .dinb(n2987), .dout(n2995));
  jor  g02766(.dina(n2995), .dinb(n791), .dout(n2996));
  jand g02767(.dina(n2995), .dinb(n791), .dout(n2997));
  jnot g02768(.din(n2743), .dout(n2998));
  jand g02769(.dina(asqrt[41] ), .dinb(n2998), .dout(n2999));
  jand g02770(.dina(n2999), .dinb(n2748), .dout(n3000));
  jor  g02771(.dina(n3000), .dinb(n2747), .dout(n3001));
  jand g02772(.dina(n2999), .dinb(n2749), .dout(n3002));
  jnot g02773(.din(n3002), .dout(n3003));
  jand g02774(.dina(n3003), .dinb(n3001), .dout(n3004));
  jnot g02775(.din(n3004), .dout(n3005));
  jor  g02776(.dina(n3005), .dinb(n2997), .dout(n3006));
  jand g02777(.dina(n3006), .dinb(n2996), .dout(n3007));
  jor  g02778(.dina(n3007), .dinb(n595), .dout(n3008));
  jand g02779(.dina(n2996), .dinb(n595), .dout(n3009));
  jand g02780(.dina(n3009), .dinb(n3006), .dout(n3010));
  jnot g02781(.din(n2751), .dout(n3011));
  jand g02782(.dina(asqrt[41] ), .dinb(n3011), .dout(n3012));
  jand g02783(.dina(n3012), .dinb(n2758), .dout(n3013));
  jor  g02784(.dina(n3013), .dinb(n2756), .dout(n3014));
  jand g02785(.dina(n3012), .dinb(n2759), .dout(n3015));
  jnot g02786(.din(n3015), .dout(n3016));
  jand g02787(.dina(n3016), .dinb(n3014), .dout(n3017));
  jnot g02788(.din(n3017), .dout(n3018));
  jor  g02789(.dina(n3018), .dinb(n3010), .dout(n3019));
  jand g02790(.dina(n3019), .dinb(n3008), .dout(n3020));
  jor  g02791(.dina(n3020), .dinb(n590), .dout(n3021));
  jxor g02792(.dina(n2760), .dinb(n595), .dout(n3022));
  jor  g02793(.dina(n3022), .dinb(n2875), .dout(n3023));
  jxor g02794(.dina(n3023), .dinb(n2771), .dout(n3024));
  jand g02795(.dina(n3020), .dinb(n590), .dout(n3025));
  jor  g02796(.dina(n3025), .dinb(n3024), .dout(n3026));
  jand g02797(.dina(n3026), .dinb(n3021), .dout(n3027));
  jor  g02798(.dina(n3027), .dinb(n430), .dout(n3028));
  jnot g02799(.din(n2776), .dout(n3029));
  jor  g02800(.dina(n3029), .dinb(n2774), .dout(n3030));
  jor  g02801(.dina(n3030), .dinb(n2875), .dout(n3031));
  jxor g02802(.dina(n3031), .dinb(n2785), .dout(n3032));
  jand g02803(.dina(n3021), .dinb(n430), .dout(n3033));
  jand g02804(.dina(n3033), .dinb(n3026), .dout(n3034));
  jor  g02805(.dina(n3034), .dinb(n3032), .dout(n3035));
  jand g02806(.dina(n3035), .dinb(n3028), .dout(n3036));
  jor  g02807(.dina(n3036), .dinb(n425), .dout(n3037));
  jand g02808(.dina(n3036), .dinb(n425), .dout(n3038));
  jnot g02809(.din(n2788), .dout(n3039));
  jand g02810(.dina(asqrt[41] ), .dinb(n3039), .dout(n3040));
  jand g02811(.dina(n3040), .dinb(n2793), .dout(n3041));
  jor  g02812(.dina(n3041), .dinb(n2792), .dout(n3042));
  jand g02813(.dina(n3040), .dinb(n2794), .dout(n3043));
  jnot g02814(.din(n3043), .dout(n3044));
  jand g02815(.dina(n3044), .dinb(n3042), .dout(n3045));
  jnot g02816(.din(n3045), .dout(n3046));
  jor  g02817(.dina(n3046), .dinb(n3038), .dout(n3047));
  jand g02818(.dina(n3047), .dinb(n3037), .dout(n3048));
  jor  g02819(.dina(n3048), .dinb(n305), .dout(n3049));
  jand g02820(.dina(n3037), .dinb(n305), .dout(n3050));
  jand g02821(.dina(n3050), .dinb(n3047), .dout(n3051));
  jnot g02822(.din(n2796), .dout(n3052));
  jand g02823(.dina(asqrt[41] ), .dinb(n3052), .dout(n3053));
  jand g02824(.dina(n3053), .dinb(n2803), .dout(n3054));
  jor  g02825(.dina(n3054), .dinb(n2801), .dout(n3055));
  jand g02826(.dina(n3053), .dinb(n2804), .dout(n3056));
  jnot g02827(.din(n3056), .dout(n3057));
  jand g02828(.dina(n3057), .dinb(n3055), .dout(n3058));
  jnot g02829(.din(n3058), .dout(n3059));
  jor  g02830(.dina(n3059), .dinb(n3051), .dout(n3060));
  jand g02831(.dina(n3060), .dinb(n3049), .dout(n3061));
  jor  g02832(.dina(n3061), .dinb(n290), .dout(n3062));
  jxor g02833(.dina(n2805), .dinb(n305), .dout(n3063));
  jor  g02834(.dina(n3063), .dinb(n2875), .dout(n3064));
  jxor g02835(.dina(n3064), .dinb(n2816), .dout(n3065));
  jand g02836(.dina(n3061), .dinb(n290), .dout(n3066));
  jor  g02837(.dina(n3066), .dinb(n3065), .dout(n3067));
  jand g02838(.dina(n3067), .dinb(n3062), .dout(n3068));
  jor  g02839(.dina(n3068), .dinb(n223), .dout(n3069));
  jnot g02840(.din(n2821), .dout(n3070));
  jor  g02841(.dina(n3070), .dinb(n2819), .dout(n3071));
  jor  g02842(.dina(n3071), .dinb(n2875), .dout(n3072));
  jxor g02843(.dina(n3072), .dinb(n2830), .dout(n3073));
  jand g02844(.dina(n3062), .dinb(n223), .dout(n3074));
  jand g02845(.dina(n3074), .dinb(n3067), .dout(n3075));
  jor  g02846(.dina(n3075), .dinb(n3073), .dout(n3076));
  jand g02847(.dina(n3076), .dinb(n3069), .dout(n3077));
  jor  g02848(.dina(n3077), .dinb(n199), .dout(n3078));
  jand g02849(.dina(n3077), .dinb(n199), .dout(n3079));
  jnot g02850(.din(n2833), .dout(n3080));
  jand g02851(.dina(asqrt[41] ), .dinb(n3080), .dout(n3081));
  jand g02852(.dina(n3081), .dinb(n2838), .dout(n3082));
  jor  g02853(.dina(n3082), .dinb(n2837), .dout(n3083));
  jand g02854(.dina(n3081), .dinb(n2839), .dout(n3084));
  jnot g02855(.din(n3084), .dout(n3085));
  jand g02856(.dina(n3085), .dinb(n3083), .dout(n3086));
  jnot g02857(.din(n3086), .dout(n3087));
  jor  g02858(.dina(n3087), .dinb(n3079), .dout(n3088));
  jand g02859(.dina(n3088), .dinb(n3078), .dout(n3089));
  jnot g02860(.din(n2841), .dout(n3090));
  jand g02861(.dina(asqrt[41] ), .dinb(n3090), .dout(n3091));
  jand g02862(.dina(n3091), .dinb(n2848), .dout(n3092));
  jor  g02863(.dina(n3092), .dinb(n2846), .dout(n3093));
  jand g02864(.dina(n3091), .dinb(n2849), .dout(n3094));
  jnot g02865(.din(n3094), .dout(n3095));
  jand g02866(.dina(n3095), .dinb(n3093), .dout(n3096));
  jnot g02867(.din(n3096), .dout(n3097));
  jand g02868(.dina(asqrt[41] ), .dinb(n2863), .dout(n3098));
  jand g02869(.dina(n3098), .dinb(n2850), .dout(n3099));
  jor  g02870(.dina(n3099), .dinb(n2895), .dout(n3100));
  jor  g02871(.dina(n3100), .dinb(n3097), .dout(n3101));
  jor  g02872(.dina(n3101), .dinb(n3089), .dout(n3102));
  jand g02873(.dina(n3102), .dinb(n194), .dout(n3103));
  jand g02874(.dina(n3097), .dinb(n3089), .dout(n3104));
  jor  g02875(.dina(n3098), .dinb(n2850), .dout(n3105));
  jand g02876(.dina(n2863), .dinb(n2850), .dout(n3106));
  jor  g02877(.dina(n3106), .dinb(n194), .dout(n3107));
  jnot g02878(.din(n3107), .dout(n3108));
  jand g02879(.dina(n3108), .dinb(n3105), .dout(n3109));
  jor  g02880(.dina(n3109), .dinb(n3104), .dout(n3112));
  jor  g02881(.dina(n3112), .dinb(n3103), .dout(asqrt[40] ));
  jand g02882(.dina(asqrt[40] ), .dinb(a[80] ), .dout(n3114));
  jnot g02883(.din(a[78] ), .dout(n3115));
  jnot g02884(.din(a[79] ), .dout(n3116));
  jand g02885(.dina(n2878), .dinb(n3116), .dout(n3117));
  jand g02886(.dina(n3117), .dinb(n3115), .dout(n3118));
  jor  g02887(.dina(n3118), .dinb(n3114), .dout(n3119));
  jand g02888(.dina(n3119), .dinb(asqrt[41] ), .dout(n3120));
  jand g02889(.dina(asqrt[40] ), .dinb(n2878), .dout(n3121));
  jxor g02890(.dina(n3121), .dinb(n2879), .dout(n3122));
  jor  g02891(.dina(n3119), .dinb(asqrt[41] ), .dout(n3123));
  jand g02892(.dina(n3123), .dinb(n3122), .dout(n3124));
  jor  g02893(.dina(n3124), .dinb(n3120), .dout(n3125));
  jand g02894(.dina(n3125), .dinb(asqrt[42] ), .dout(n3126));
  jor  g02895(.dina(n3120), .dinb(asqrt[42] ), .dout(n3127));
  jor  g02896(.dina(n3127), .dinb(n3124), .dout(n3128));
  jand g02897(.dina(n3121), .dinb(n2879), .dout(n3129));
  jnot g02898(.din(n3103), .dout(n3130));
  jnot g02899(.din(n3104), .dout(n3131));
  jnot g02900(.din(n3109), .dout(n3132));
  jand g02901(.dina(n3132), .dinb(asqrt[41] ), .dout(n3133));
  jand g02902(.dina(n3133), .dinb(n3131), .dout(n3134));
  jand g02903(.dina(n3134), .dinb(n3130), .dout(n3135));
  jor  g02904(.dina(n3135), .dinb(n3129), .dout(n3136));
  jxor g02905(.dina(n3136), .dinb(n2640), .dout(n3137));
  jand g02906(.dina(n3137), .dinb(n3128), .dout(n3138));
  jor  g02907(.dina(n3138), .dinb(n3126), .dout(n3139));
  jand g02908(.dina(n3139), .dinb(asqrt[43] ), .dout(n3140));
  jor  g02909(.dina(n3139), .dinb(asqrt[43] ), .dout(n3141));
  jxor g02910(.dina(n2883), .dinb(n2870), .dout(n3142));
  jand g02911(.dina(n3142), .dinb(asqrt[40] ), .dout(n3143));
  jxor g02912(.dina(n3143), .dinb(n2886), .dout(n3144));
  jnot g02913(.din(n3144), .dout(n3145));
  jand g02914(.dina(n3145), .dinb(n3141), .dout(n3146));
  jor  g02915(.dina(n3146), .dinb(n3140), .dout(n3147));
  jand g02916(.dina(n3147), .dinb(asqrt[44] ), .dout(n3148));
  jnot g02917(.din(n2892), .dout(n3149));
  jand g02918(.dina(n3149), .dinb(n2890), .dout(n3150));
  jand g02919(.dina(n3150), .dinb(asqrt[40] ), .dout(n3151));
  jxor g02920(.dina(n3151), .dinb(n2900), .dout(n3152));
  jnot g02921(.din(n3152), .dout(n3153));
  jor  g02922(.dina(n3140), .dinb(asqrt[44] ), .dout(n3154));
  jor  g02923(.dina(n3154), .dinb(n3146), .dout(n3155));
  jand g02924(.dina(n3155), .dinb(n3153), .dout(n3156));
  jor  g02925(.dina(n3156), .dinb(n3148), .dout(n3157));
  jand g02926(.dina(n3157), .dinb(asqrt[45] ), .dout(n3158));
  jor  g02927(.dina(n3157), .dinb(asqrt[45] ), .dout(n3159));
  jnot g02928(.din(n2907), .dout(n3160));
  jxor g02929(.dina(n2902), .dinb(n2420), .dout(n3161));
  jand g02930(.dina(n3161), .dinb(asqrt[40] ), .dout(n3162));
  jxor g02931(.dina(n3162), .dinb(n3160), .dout(n3163));
  jand g02932(.dina(n3163), .dinb(n3159), .dout(n3164));
  jor  g02933(.dina(n3164), .dinb(n3158), .dout(n3165));
  jand g02934(.dina(n3165), .dinb(asqrt[46] ), .dout(n3166));
  jor  g02935(.dina(n3158), .dinb(asqrt[46] ), .dout(n3167));
  jor  g02936(.dina(n3167), .dinb(n3164), .dout(n3168));
  jnot g02937(.din(n2914), .dout(n3169));
  jnot g02938(.din(n2916), .dout(n3170));
  jand g02939(.dina(asqrt[40] ), .dinb(n2910), .dout(n3171));
  jand g02940(.dina(n3171), .dinb(n3170), .dout(n3172));
  jor  g02941(.dina(n3172), .dinb(n3169), .dout(n3173));
  jnot g02942(.din(n2917), .dout(n3174));
  jand g02943(.dina(n3171), .dinb(n3174), .dout(n3175));
  jnot g02944(.din(n3175), .dout(n3176));
  jand g02945(.dina(n3176), .dinb(n3173), .dout(n3177));
  jand g02946(.dina(n3177), .dinb(n3168), .dout(n3178));
  jor  g02947(.dina(n3178), .dinb(n3166), .dout(n3179));
  jand g02948(.dina(n3179), .dinb(asqrt[47] ), .dout(n3180));
  jor  g02949(.dina(n3179), .dinb(asqrt[47] ), .dout(n3181));
  jxor g02950(.dina(n2918), .dinb(n2005), .dout(n3182));
  jand g02951(.dina(n3182), .dinb(asqrt[40] ), .dout(n3183));
  jxor g02952(.dina(n3183), .dinb(n2923), .dout(n3184));
  jand g02953(.dina(n3184), .dinb(n3181), .dout(n3185));
  jor  g02954(.dina(n3185), .dinb(n3180), .dout(n3186));
  jand g02955(.dina(n3186), .dinb(asqrt[48] ), .dout(n3187));
  jnot g02956(.din(n2929), .dout(n3188));
  jand g02957(.dina(n3188), .dinb(n2927), .dout(n3189));
  jand g02958(.dina(n3189), .dinb(asqrt[40] ), .dout(n3190));
  jxor g02959(.dina(n3190), .dinb(n2937), .dout(n3191));
  jnot g02960(.din(n3191), .dout(n3192));
  jor  g02961(.dina(n3180), .dinb(asqrt[48] ), .dout(n3193));
  jor  g02962(.dina(n3193), .dinb(n3185), .dout(n3194));
  jand g02963(.dina(n3194), .dinb(n3192), .dout(n3195));
  jor  g02964(.dina(n3195), .dinb(n3187), .dout(n3196));
  jand g02965(.dina(n3196), .dinb(asqrt[49] ), .dout(n3197));
  jor  g02966(.dina(n3196), .dinb(asqrt[49] ), .dout(n3198));
  jxor g02967(.dina(n2939), .dinb(n1641), .dout(n3199));
  jand g02968(.dina(n3199), .dinb(asqrt[40] ), .dout(n3200));
  jxor g02969(.dina(n3200), .dinb(n2945), .dout(n3201));
  jand g02970(.dina(n3201), .dinb(n3198), .dout(n3202));
  jor  g02971(.dina(n3202), .dinb(n3197), .dout(n3203));
  jand g02972(.dina(n3203), .dinb(asqrt[50] ), .dout(n3204));
  jor  g02973(.dina(n3197), .dinb(asqrt[50] ), .dout(n3205));
  jor  g02974(.dina(n3205), .dinb(n3202), .dout(n3206));
  jnot g02975(.din(n2953), .dout(n3207));
  jnot g02976(.din(n2955), .dout(n3208));
  jand g02977(.dina(asqrt[40] ), .dinb(n2949), .dout(n3209));
  jand g02978(.dina(n3209), .dinb(n3208), .dout(n3210));
  jor  g02979(.dina(n3210), .dinb(n3207), .dout(n3211));
  jnot g02980(.din(n2956), .dout(n3212));
  jand g02981(.dina(n3209), .dinb(n3212), .dout(n3213));
  jnot g02982(.din(n3213), .dout(n3214));
  jand g02983(.dina(n3214), .dinb(n3211), .dout(n3215));
  jand g02984(.dina(n3215), .dinb(n3206), .dout(n3216));
  jor  g02985(.dina(n3216), .dinb(n3204), .dout(n3217));
  jand g02986(.dina(n3217), .dinb(asqrt[51] ), .dout(n3218));
  jxor g02987(.dina(n2957), .dinb(n1312), .dout(n3219));
  jand g02988(.dina(n3219), .dinb(asqrt[40] ), .dout(n3220));
  jxor g02989(.dina(n3220), .dinb(n2964), .dout(n3221));
  jnot g02990(.din(n3221), .dout(n3222));
  jor  g02991(.dina(n3217), .dinb(asqrt[51] ), .dout(n3223));
  jand g02992(.dina(n3223), .dinb(n3222), .dout(n3224));
  jor  g02993(.dina(n3224), .dinb(n3218), .dout(n3225));
  jand g02994(.dina(n3225), .dinb(asqrt[52] ), .dout(n3226));
  jnot g02995(.din(n2969), .dout(n3227));
  jand g02996(.dina(n3227), .dinb(n2967), .dout(n3228));
  jand g02997(.dina(n3228), .dinb(asqrt[40] ), .dout(n3229));
  jxor g02998(.dina(n3229), .dinb(n2977), .dout(n3230));
  jnot g02999(.din(n3230), .dout(n3231));
  jor  g03000(.dina(n3218), .dinb(asqrt[52] ), .dout(n3232));
  jor  g03001(.dina(n3232), .dinb(n3224), .dout(n3233));
  jand g03002(.dina(n3233), .dinb(n3231), .dout(n3234));
  jor  g03003(.dina(n3234), .dinb(n3226), .dout(n3235));
  jand g03004(.dina(n3235), .dinb(asqrt[53] ), .dout(n3236));
  jor  g03005(.dina(n3235), .dinb(asqrt[53] ), .dout(n3237));
  jnot g03006(.din(n2983), .dout(n3238));
  jnot g03007(.din(n2984), .dout(n3239));
  jand g03008(.dina(asqrt[40] ), .dinb(n2980), .dout(n3240));
  jand g03009(.dina(n3240), .dinb(n3239), .dout(n3241));
  jor  g03010(.dina(n3241), .dinb(n3238), .dout(n3242));
  jnot g03011(.din(n2985), .dout(n3243));
  jand g03012(.dina(n3240), .dinb(n3243), .dout(n3244));
  jnot g03013(.din(n3244), .dout(n3245));
  jand g03014(.dina(n3245), .dinb(n3242), .dout(n3246));
  jand g03015(.dina(n3246), .dinb(n3237), .dout(n3247));
  jor  g03016(.dina(n3247), .dinb(n3236), .dout(n3248));
  jand g03017(.dina(n3248), .dinb(asqrt[54] ), .dout(n3249));
  jor  g03018(.dina(n3236), .dinb(asqrt[54] ), .dout(n3250));
  jor  g03019(.dina(n3250), .dinb(n3247), .dout(n3251));
  jnot g03020(.din(n2991), .dout(n3252));
  jnot g03021(.din(n2993), .dout(n3253));
  jand g03022(.dina(asqrt[40] ), .dinb(n2987), .dout(n3254));
  jand g03023(.dina(n3254), .dinb(n3253), .dout(n3255));
  jor  g03024(.dina(n3255), .dinb(n3252), .dout(n3256));
  jnot g03025(.din(n2994), .dout(n3257));
  jand g03026(.dina(n3254), .dinb(n3257), .dout(n3258));
  jnot g03027(.din(n3258), .dout(n3259));
  jand g03028(.dina(n3259), .dinb(n3256), .dout(n3260));
  jand g03029(.dina(n3260), .dinb(n3251), .dout(n3261));
  jor  g03030(.dina(n3261), .dinb(n3249), .dout(n3262));
  jand g03031(.dina(n3262), .dinb(asqrt[55] ), .dout(n3263));
  jxor g03032(.dina(n2995), .dinb(n791), .dout(n3264));
  jand g03033(.dina(n3264), .dinb(asqrt[40] ), .dout(n3265));
  jxor g03034(.dina(n3265), .dinb(n3005), .dout(n3266));
  jnot g03035(.din(n3266), .dout(n3267));
  jor  g03036(.dina(n3262), .dinb(asqrt[55] ), .dout(n3268));
  jand g03037(.dina(n3268), .dinb(n3267), .dout(n3269));
  jor  g03038(.dina(n3269), .dinb(n3263), .dout(n3270));
  jand g03039(.dina(n3270), .dinb(asqrt[56] ), .dout(n3271));
  jnot g03040(.din(n3010), .dout(n3272));
  jand g03041(.dina(n3272), .dinb(n3008), .dout(n3273));
  jand g03042(.dina(n3273), .dinb(asqrt[40] ), .dout(n3274));
  jxor g03043(.dina(n3274), .dinb(n3018), .dout(n3275));
  jnot g03044(.din(n3275), .dout(n3276));
  jor  g03045(.dina(n3263), .dinb(asqrt[56] ), .dout(n3277));
  jor  g03046(.dina(n3277), .dinb(n3269), .dout(n3278));
  jand g03047(.dina(n3278), .dinb(n3276), .dout(n3279));
  jor  g03048(.dina(n3279), .dinb(n3271), .dout(n3280));
  jand g03049(.dina(n3280), .dinb(asqrt[57] ), .dout(n3281));
  jor  g03050(.dina(n3280), .dinb(asqrt[57] ), .dout(n3282));
  jnot g03051(.din(n3024), .dout(n3283));
  jnot g03052(.din(n3025), .dout(n3284));
  jand g03053(.dina(asqrt[40] ), .dinb(n3021), .dout(n3285));
  jand g03054(.dina(n3285), .dinb(n3284), .dout(n3286));
  jor  g03055(.dina(n3286), .dinb(n3283), .dout(n3287));
  jnot g03056(.din(n3026), .dout(n3288));
  jand g03057(.dina(n3285), .dinb(n3288), .dout(n3289));
  jnot g03058(.din(n3289), .dout(n3290));
  jand g03059(.dina(n3290), .dinb(n3287), .dout(n3291));
  jand g03060(.dina(n3291), .dinb(n3282), .dout(n3292));
  jor  g03061(.dina(n3292), .dinb(n3281), .dout(n3293));
  jand g03062(.dina(n3293), .dinb(asqrt[58] ), .dout(n3294));
  jor  g03063(.dina(n3281), .dinb(asqrt[58] ), .dout(n3295));
  jor  g03064(.dina(n3295), .dinb(n3292), .dout(n3296));
  jnot g03065(.din(n3032), .dout(n3297));
  jnot g03066(.din(n3034), .dout(n3298));
  jand g03067(.dina(asqrt[40] ), .dinb(n3028), .dout(n3299));
  jand g03068(.dina(n3299), .dinb(n3298), .dout(n3300));
  jor  g03069(.dina(n3300), .dinb(n3297), .dout(n3301));
  jnot g03070(.din(n3035), .dout(n3302));
  jand g03071(.dina(n3299), .dinb(n3302), .dout(n3303));
  jnot g03072(.din(n3303), .dout(n3304));
  jand g03073(.dina(n3304), .dinb(n3301), .dout(n3305));
  jand g03074(.dina(n3305), .dinb(n3296), .dout(n3306));
  jor  g03075(.dina(n3306), .dinb(n3294), .dout(n3307));
  jand g03076(.dina(n3307), .dinb(asqrt[59] ), .dout(n3308));
  jxor g03077(.dina(n3036), .dinb(n425), .dout(n3309));
  jand g03078(.dina(n3309), .dinb(asqrt[40] ), .dout(n3310));
  jxor g03079(.dina(n3310), .dinb(n3046), .dout(n3311));
  jnot g03080(.din(n3311), .dout(n3312));
  jor  g03081(.dina(n3307), .dinb(asqrt[59] ), .dout(n3313));
  jand g03082(.dina(n3313), .dinb(n3312), .dout(n3314));
  jor  g03083(.dina(n3314), .dinb(n3308), .dout(n3315));
  jand g03084(.dina(n3315), .dinb(asqrt[60] ), .dout(n3316));
  jnot g03085(.din(n3051), .dout(n3317));
  jand g03086(.dina(n3317), .dinb(n3049), .dout(n3318));
  jand g03087(.dina(n3318), .dinb(asqrt[40] ), .dout(n3319));
  jxor g03088(.dina(n3319), .dinb(n3059), .dout(n3320));
  jnot g03089(.din(n3320), .dout(n3321));
  jor  g03090(.dina(n3308), .dinb(asqrt[60] ), .dout(n3322));
  jor  g03091(.dina(n3322), .dinb(n3314), .dout(n3323));
  jand g03092(.dina(n3323), .dinb(n3321), .dout(n3324));
  jor  g03093(.dina(n3324), .dinb(n3316), .dout(n3325));
  jand g03094(.dina(n3325), .dinb(asqrt[61] ), .dout(n3326));
  jor  g03095(.dina(n3325), .dinb(asqrt[61] ), .dout(n3327));
  jnot g03096(.din(n3065), .dout(n3328));
  jnot g03097(.din(n3066), .dout(n3329));
  jand g03098(.dina(asqrt[40] ), .dinb(n3062), .dout(n3330));
  jand g03099(.dina(n3330), .dinb(n3329), .dout(n3331));
  jor  g03100(.dina(n3331), .dinb(n3328), .dout(n3332));
  jnot g03101(.din(n3067), .dout(n3333));
  jand g03102(.dina(n3330), .dinb(n3333), .dout(n3334));
  jnot g03103(.din(n3334), .dout(n3335));
  jand g03104(.dina(n3335), .dinb(n3332), .dout(n3336));
  jand g03105(.dina(n3336), .dinb(n3327), .dout(n3337));
  jor  g03106(.dina(n3337), .dinb(n3326), .dout(n3338));
  jand g03107(.dina(n3338), .dinb(asqrt[62] ), .dout(n3339));
  jor  g03108(.dina(n3326), .dinb(asqrt[62] ), .dout(n3340));
  jor  g03109(.dina(n3340), .dinb(n3337), .dout(n3341));
  jnot g03110(.din(n3073), .dout(n3342));
  jnot g03111(.din(n3075), .dout(n3343));
  jand g03112(.dina(asqrt[40] ), .dinb(n3069), .dout(n3344));
  jand g03113(.dina(n3344), .dinb(n3343), .dout(n3345));
  jor  g03114(.dina(n3345), .dinb(n3342), .dout(n3346));
  jnot g03115(.din(n3076), .dout(n3347));
  jand g03116(.dina(n3344), .dinb(n3347), .dout(n3348));
  jnot g03117(.din(n3348), .dout(n3349));
  jand g03118(.dina(n3349), .dinb(n3346), .dout(n3350));
  jand g03119(.dina(n3350), .dinb(n3341), .dout(n3351));
  jor  g03120(.dina(n3351), .dinb(n3339), .dout(n3352));
  jxor g03121(.dina(n3077), .dinb(n199), .dout(n3353));
  jand g03122(.dina(n3353), .dinb(asqrt[40] ), .dout(n3354));
  jxor g03123(.dina(n3354), .dinb(n3087), .dout(n3355));
  jnot g03124(.din(n3089), .dout(n3356));
  jand g03125(.dina(asqrt[40] ), .dinb(n3096), .dout(n3357));
  jand g03126(.dina(n3357), .dinb(n3356), .dout(n3358));
  jor  g03127(.dina(n3358), .dinb(n3104), .dout(n3359));
  jor  g03128(.dina(n3359), .dinb(n3355), .dout(n3360));
  jnot g03129(.din(n3360), .dout(n3361));
  jand g03130(.dina(n3361), .dinb(n3352), .dout(n3362));
  jor  g03131(.dina(n3362), .dinb(asqrt[63] ), .dout(n3363));
  jnot g03132(.din(n3355), .dout(n3364));
  jor  g03133(.dina(n3364), .dinb(n3352), .dout(n3365));
  jor  g03134(.dina(n3357), .dinb(n3356), .dout(n3366));
  jand g03135(.dina(n3096), .dinb(n3356), .dout(n3367));
  jor  g03136(.dina(n3367), .dinb(n194), .dout(n3368));
  jnot g03137(.din(n3368), .dout(n3369));
  jand g03138(.dina(n3369), .dinb(n3366), .dout(n3370));
  jnot g03139(.din(asqrt[40] ), .dout(n3371));
  jnot g03140(.din(n3370), .dout(n3374));
  jand g03141(.dina(n3374), .dinb(n3365), .dout(n3375));
  jand g03142(.dina(n3375), .dinb(n3363), .dout(n3376));
  jnot g03143(.din(n3376), .dout(asqrt[39] ));
  jor  g03144(.dina(n3376), .dinb(n3115), .dout(n3378));
  jnot g03145(.din(a[76] ), .dout(n3379));
  jnot g03146(.din(a[77] ), .dout(n3380));
  jand g03147(.dina(n3115), .dinb(n3380), .dout(n3381));
  jand g03148(.dina(n3381), .dinb(n3379), .dout(n3382));
  jnot g03149(.din(n3382), .dout(n3383));
  jand g03150(.dina(n3383), .dinb(n3378), .dout(n3384));
  jor  g03151(.dina(n3384), .dinb(n3371), .dout(n3385));
  jor  g03152(.dina(n3376), .dinb(a[78] ), .dout(n3386));
  jxor g03153(.dina(n3386), .dinb(n3116), .dout(n3387));
  jand g03154(.dina(n3384), .dinb(n3371), .dout(n3388));
  jor  g03155(.dina(n3388), .dinb(n3387), .dout(n3389));
  jand g03156(.dina(n3389), .dinb(n3385), .dout(n3390));
  jor  g03157(.dina(n3390), .dinb(n2875), .dout(n3391));
  jand g03158(.dina(n3385), .dinb(n2875), .dout(n3392));
  jand g03159(.dina(n3392), .dinb(n3389), .dout(n3393));
  jor  g03160(.dina(n3386), .dinb(a[79] ), .dout(n3394));
  jnot g03161(.din(n3363), .dout(n3395));
  jnot g03162(.din(n3365), .dout(n3396));
  jor  g03163(.dina(n3370), .dinb(n3371), .dout(n3397));
  jor  g03164(.dina(n3397), .dinb(n3396), .dout(n3398));
  jor  g03165(.dina(n3398), .dinb(n3395), .dout(n3399));
  jand g03166(.dina(n3399), .dinb(n3394), .dout(n3400));
  jxor g03167(.dina(n3400), .dinb(n2878), .dout(n3401));
  jor  g03168(.dina(n3401), .dinb(n3393), .dout(n3402));
  jand g03169(.dina(n3402), .dinb(n3391), .dout(n3403));
  jor  g03170(.dina(n3403), .dinb(n2870), .dout(n3404));
  jand g03171(.dina(n3403), .dinb(n2870), .dout(n3405));
  jxor g03172(.dina(n3119), .dinb(n2875), .dout(n3406));
  jor  g03173(.dina(n3406), .dinb(n3376), .dout(n3407));
  jxor g03174(.dina(n3407), .dinb(n3122), .dout(n3408));
  jor  g03175(.dina(n3408), .dinb(n3405), .dout(n3409));
  jand g03176(.dina(n3409), .dinb(n3404), .dout(n3410));
  jor  g03177(.dina(n3410), .dinb(n2425), .dout(n3411));
  jnot g03178(.din(n3128), .dout(n3412));
  jor  g03179(.dina(n3412), .dinb(n3126), .dout(n3413));
  jor  g03180(.dina(n3413), .dinb(n3376), .dout(n3414));
  jxor g03181(.dina(n3414), .dinb(n3137), .dout(n3415));
  jand g03182(.dina(n3404), .dinb(n2425), .dout(n3416));
  jand g03183(.dina(n3416), .dinb(n3409), .dout(n3417));
  jor  g03184(.dina(n3417), .dinb(n3415), .dout(n3418));
  jand g03185(.dina(n3418), .dinb(n3411), .dout(n3419));
  jor  g03186(.dina(n3419), .dinb(n2420), .dout(n3420));
  jand g03187(.dina(n3419), .dinb(n2420), .dout(n3421));
  jxor g03188(.dina(n3139), .dinb(n2425), .dout(n3422));
  jor  g03189(.dina(n3422), .dinb(n3376), .dout(n3423));
  jxor g03190(.dina(n3423), .dinb(n3144), .dout(n3424));
  jnot g03191(.din(n3424), .dout(n3425));
  jor  g03192(.dina(n3425), .dinb(n3421), .dout(n3426));
  jand g03193(.dina(n3426), .dinb(n3420), .dout(n3427));
  jor  g03194(.dina(n3427), .dinb(n2010), .dout(n3428));
  jand g03195(.dina(n3420), .dinb(n2010), .dout(n3429));
  jand g03196(.dina(n3429), .dinb(n3426), .dout(n3430));
  jnot g03197(.din(n3148), .dout(n3431));
  jand g03198(.dina(asqrt[39] ), .dinb(n3431), .dout(n3432));
  jand g03199(.dina(n3432), .dinb(n3155), .dout(n3433));
  jor  g03200(.dina(n3433), .dinb(n3153), .dout(n3434));
  jand g03201(.dina(n3432), .dinb(n3156), .dout(n3435));
  jnot g03202(.din(n3435), .dout(n3436));
  jand g03203(.dina(n3436), .dinb(n3434), .dout(n3437));
  jnot g03204(.din(n3437), .dout(n3438));
  jor  g03205(.dina(n3438), .dinb(n3430), .dout(n3439));
  jand g03206(.dina(n3439), .dinb(n3428), .dout(n3440));
  jor  g03207(.dina(n3440), .dinb(n2005), .dout(n3441));
  jand g03208(.dina(n3440), .dinb(n2005), .dout(n3442));
  jnot g03209(.din(n3163), .dout(n3443));
  jxor g03210(.dina(n3157), .dinb(n2010), .dout(n3444));
  jor  g03211(.dina(n3444), .dinb(n3376), .dout(n3445));
  jxor g03212(.dina(n3445), .dinb(n3443), .dout(n3446));
  jnot g03213(.din(n3446), .dout(n3447));
  jor  g03214(.dina(n3447), .dinb(n3442), .dout(n3448));
  jand g03215(.dina(n3448), .dinb(n3441), .dout(n3449));
  jor  g03216(.dina(n3449), .dinb(n1646), .dout(n3450));
  jnot g03217(.din(n3168), .dout(n3451));
  jor  g03218(.dina(n3451), .dinb(n3166), .dout(n3452));
  jor  g03219(.dina(n3452), .dinb(n3376), .dout(n3453));
  jxor g03220(.dina(n3453), .dinb(n3177), .dout(n3454));
  jand g03221(.dina(n3441), .dinb(n1646), .dout(n3455));
  jand g03222(.dina(n3455), .dinb(n3448), .dout(n3456));
  jor  g03223(.dina(n3456), .dinb(n3454), .dout(n3457));
  jand g03224(.dina(n3457), .dinb(n3450), .dout(n3458));
  jor  g03225(.dina(n3458), .dinb(n1641), .dout(n3459));
  jand g03226(.dina(n3458), .dinb(n1641), .dout(n3460));
  jnot g03227(.din(n3184), .dout(n3461));
  jxor g03228(.dina(n3179), .dinb(n1646), .dout(n3462));
  jor  g03229(.dina(n3462), .dinb(n3376), .dout(n3463));
  jxor g03230(.dina(n3463), .dinb(n3461), .dout(n3464));
  jnot g03231(.din(n3464), .dout(n3465));
  jor  g03232(.dina(n3465), .dinb(n3460), .dout(n3466));
  jand g03233(.dina(n3466), .dinb(n3459), .dout(n3467));
  jor  g03234(.dina(n3467), .dinb(n1317), .dout(n3468));
  jand g03235(.dina(n3459), .dinb(n1317), .dout(n3469));
  jand g03236(.dina(n3469), .dinb(n3466), .dout(n3470));
  jnot g03237(.din(n3187), .dout(n3471));
  jand g03238(.dina(asqrt[39] ), .dinb(n3471), .dout(n3472));
  jand g03239(.dina(n3472), .dinb(n3194), .dout(n3473));
  jor  g03240(.dina(n3473), .dinb(n3192), .dout(n3474));
  jand g03241(.dina(n3472), .dinb(n3195), .dout(n3475));
  jnot g03242(.din(n3475), .dout(n3476));
  jand g03243(.dina(n3476), .dinb(n3474), .dout(n3477));
  jnot g03244(.din(n3477), .dout(n3478));
  jor  g03245(.dina(n3478), .dinb(n3470), .dout(n3479));
  jand g03246(.dina(n3479), .dinb(n3468), .dout(n3480));
  jor  g03247(.dina(n3480), .dinb(n1312), .dout(n3481));
  jxor g03248(.dina(n3196), .dinb(n1317), .dout(n3482));
  jor  g03249(.dina(n3482), .dinb(n3376), .dout(n3483));
  jxor g03250(.dina(n3483), .dinb(n3201), .dout(n3484));
  jand g03251(.dina(n3480), .dinb(n1312), .dout(n3485));
  jor  g03252(.dina(n3485), .dinb(n3484), .dout(n3486));
  jand g03253(.dina(n3486), .dinb(n3481), .dout(n3487));
  jor  g03254(.dina(n3487), .dinb(n1039), .dout(n3488));
  jnot g03255(.din(n3206), .dout(n3489));
  jor  g03256(.dina(n3489), .dinb(n3204), .dout(n3490));
  jor  g03257(.dina(n3490), .dinb(n3376), .dout(n3491));
  jxor g03258(.dina(n3491), .dinb(n3215), .dout(n3492));
  jand g03259(.dina(n3481), .dinb(n1039), .dout(n3493));
  jand g03260(.dina(n3493), .dinb(n3486), .dout(n3494));
  jor  g03261(.dina(n3494), .dinb(n3492), .dout(n3495));
  jand g03262(.dina(n3495), .dinb(n3488), .dout(n3496));
  jor  g03263(.dina(n3496), .dinb(n1034), .dout(n3497));
  jand g03264(.dina(n3496), .dinb(n1034), .dout(n3498));
  jnot g03265(.din(n3218), .dout(n3499));
  jand g03266(.dina(asqrt[39] ), .dinb(n3499), .dout(n3500));
  jand g03267(.dina(n3500), .dinb(n3223), .dout(n3501));
  jor  g03268(.dina(n3501), .dinb(n3222), .dout(n3502));
  jand g03269(.dina(n3500), .dinb(n3224), .dout(n3503));
  jnot g03270(.din(n3503), .dout(n3504));
  jand g03271(.dina(n3504), .dinb(n3502), .dout(n3505));
  jnot g03272(.din(n3505), .dout(n3506));
  jor  g03273(.dina(n3506), .dinb(n3498), .dout(n3507));
  jand g03274(.dina(n3507), .dinb(n3497), .dout(n3508));
  jor  g03275(.dina(n3508), .dinb(n796), .dout(n3509));
  jand g03276(.dina(n3497), .dinb(n796), .dout(n3510));
  jand g03277(.dina(n3510), .dinb(n3507), .dout(n3511));
  jnot g03278(.din(n3226), .dout(n3512));
  jand g03279(.dina(asqrt[39] ), .dinb(n3512), .dout(n3513));
  jand g03280(.dina(n3513), .dinb(n3233), .dout(n3514));
  jor  g03281(.dina(n3514), .dinb(n3231), .dout(n3515));
  jand g03282(.dina(n3513), .dinb(n3234), .dout(n3516));
  jnot g03283(.din(n3516), .dout(n3517));
  jand g03284(.dina(n3517), .dinb(n3515), .dout(n3518));
  jnot g03285(.din(n3518), .dout(n3519));
  jor  g03286(.dina(n3519), .dinb(n3511), .dout(n3520));
  jand g03287(.dina(n3520), .dinb(n3509), .dout(n3521));
  jor  g03288(.dina(n3521), .dinb(n791), .dout(n3522));
  jxor g03289(.dina(n3235), .dinb(n796), .dout(n3523));
  jor  g03290(.dina(n3523), .dinb(n3376), .dout(n3524));
  jxor g03291(.dina(n3524), .dinb(n3246), .dout(n3525));
  jand g03292(.dina(n3521), .dinb(n791), .dout(n3526));
  jor  g03293(.dina(n3526), .dinb(n3525), .dout(n3527));
  jand g03294(.dina(n3527), .dinb(n3522), .dout(n3528));
  jor  g03295(.dina(n3528), .dinb(n595), .dout(n3529));
  jnot g03296(.din(n3251), .dout(n3530));
  jor  g03297(.dina(n3530), .dinb(n3249), .dout(n3531));
  jor  g03298(.dina(n3531), .dinb(n3376), .dout(n3532));
  jxor g03299(.dina(n3532), .dinb(n3260), .dout(n3533));
  jand g03300(.dina(n3522), .dinb(n595), .dout(n3534));
  jand g03301(.dina(n3534), .dinb(n3527), .dout(n3535));
  jor  g03302(.dina(n3535), .dinb(n3533), .dout(n3536));
  jand g03303(.dina(n3536), .dinb(n3529), .dout(n3537));
  jor  g03304(.dina(n3537), .dinb(n590), .dout(n3538));
  jand g03305(.dina(n3537), .dinb(n590), .dout(n3539));
  jnot g03306(.din(n3263), .dout(n3540));
  jand g03307(.dina(asqrt[39] ), .dinb(n3540), .dout(n3541));
  jand g03308(.dina(n3541), .dinb(n3268), .dout(n3542));
  jor  g03309(.dina(n3542), .dinb(n3267), .dout(n3543));
  jand g03310(.dina(n3541), .dinb(n3269), .dout(n3544));
  jnot g03311(.din(n3544), .dout(n3545));
  jand g03312(.dina(n3545), .dinb(n3543), .dout(n3546));
  jnot g03313(.din(n3546), .dout(n3547));
  jor  g03314(.dina(n3547), .dinb(n3539), .dout(n3548));
  jand g03315(.dina(n3548), .dinb(n3538), .dout(n3549));
  jor  g03316(.dina(n3549), .dinb(n430), .dout(n3550));
  jand g03317(.dina(n3538), .dinb(n430), .dout(n3551));
  jand g03318(.dina(n3551), .dinb(n3548), .dout(n3552));
  jnot g03319(.din(n3271), .dout(n3553));
  jand g03320(.dina(asqrt[39] ), .dinb(n3553), .dout(n3554));
  jand g03321(.dina(n3554), .dinb(n3278), .dout(n3555));
  jor  g03322(.dina(n3555), .dinb(n3276), .dout(n3556));
  jand g03323(.dina(n3554), .dinb(n3279), .dout(n3557));
  jnot g03324(.din(n3557), .dout(n3558));
  jand g03325(.dina(n3558), .dinb(n3556), .dout(n3559));
  jnot g03326(.din(n3559), .dout(n3560));
  jor  g03327(.dina(n3560), .dinb(n3552), .dout(n3561));
  jand g03328(.dina(n3561), .dinb(n3550), .dout(n3562));
  jor  g03329(.dina(n3562), .dinb(n425), .dout(n3563));
  jxor g03330(.dina(n3280), .dinb(n430), .dout(n3564));
  jor  g03331(.dina(n3564), .dinb(n3376), .dout(n3565));
  jxor g03332(.dina(n3565), .dinb(n3291), .dout(n3566));
  jand g03333(.dina(n3562), .dinb(n425), .dout(n3567));
  jor  g03334(.dina(n3567), .dinb(n3566), .dout(n3568));
  jand g03335(.dina(n3568), .dinb(n3563), .dout(n3569));
  jor  g03336(.dina(n3569), .dinb(n305), .dout(n3570));
  jnot g03337(.din(n3296), .dout(n3571));
  jor  g03338(.dina(n3571), .dinb(n3294), .dout(n3572));
  jor  g03339(.dina(n3572), .dinb(n3376), .dout(n3573));
  jxor g03340(.dina(n3573), .dinb(n3305), .dout(n3574));
  jand g03341(.dina(n3563), .dinb(n305), .dout(n3575));
  jand g03342(.dina(n3575), .dinb(n3568), .dout(n3576));
  jor  g03343(.dina(n3576), .dinb(n3574), .dout(n3577));
  jand g03344(.dina(n3577), .dinb(n3570), .dout(n3578));
  jor  g03345(.dina(n3578), .dinb(n290), .dout(n3579));
  jand g03346(.dina(n3578), .dinb(n290), .dout(n3580));
  jnot g03347(.din(n3308), .dout(n3581));
  jand g03348(.dina(asqrt[39] ), .dinb(n3581), .dout(n3582));
  jand g03349(.dina(n3582), .dinb(n3313), .dout(n3583));
  jor  g03350(.dina(n3583), .dinb(n3312), .dout(n3584));
  jand g03351(.dina(n3582), .dinb(n3314), .dout(n3585));
  jnot g03352(.din(n3585), .dout(n3586));
  jand g03353(.dina(n3586), .dinb(n3584), .dout(n3587));
  jnot g03354(.din(n3587), .dout(n3588));
  jor  g03355(.dina(n3588), .dinb(n3580), .dout(n3589));
  jand g03356(.dina(n3589), .dinb(n3579), .dout(n3590));
  jor  g03357(.dina(n3590), .dinb(n223), .dout(n3591));
  jand g03358(.dina(n3579), .dinb(n223), .dout(n3592));
  jand g03359(.dina(n3592), .dinb(n3589), .dout(n3593));
  jnot g03360(.din(n3316), .dout(n3594));
  jand g03361(.dina(asqrt[39] ), .dinb(n3594), .dout(n3595));
  jand g03362(.dina(n3595), .dinb(n3323), .dout(n3596));
  jor  g03363(.dina(n3596), .dinb(n3321), .dout(n3597));
  jand g03364(.dina(n3595), .dinb(n3324), .dout(n3598));
  jnot g03365(.din(n3598), .dout(n3599));
  jand g03366(.dina(n3599), .dinb(n3597), .dout(n3600));
  jnot g03367(.din(n3600), .dout(n3601));
  jor  g03368(.dina(n3601), .dinb(n3593), .dout(n3602));
  jand g03369(.dina(n3602), .dinb(n3591), .dout(n3603));
  jor  g03370(.dina(n3603), .dinb(n199), .dout(n3604));
  jand g03371(.dina(n3603), .dinb(n199), .dout(n3605));
  jxor g03372(.dina(n3325), .dinb(n223), .dout(n3606));
  jor  g03373(.dina(n3606), .dinb(n3376), .dout(n3607));
  jxor g03374(.dina(n3607), .dinb(n3336), .dout(n3608));
  jor  g03375(.dina(n3608), .dinb(n3605), .dout(n3609));
  jand g03376(.dina(n3609), .dinb(n3604), .dout(n3610));
  jnot g03377(.din(n3341), .dout(n3611));
  jor  g03378(.dina(n3611), .dinb(n3339), .dout(n3612));
  jor  g03379(.dina(n3612), .dinb(n3376), .dout(n3613));
  jxor g03380(.dina(n3613), .dinb(n3350), .dout(n3614));
  jand g03381(.dina(asqrt[39] ), .dinb(n3364), .dout(n3615));
  jand g03382(.dina(n3615), .dinb(n3352), .dout(n3616));
  jor  g03383(.dina(n3616), .dinb(n3396), .dout(n3617));
  jor  g03384(.dina(n3617), .dinb(n3614), .dout(n3618));
  jor  g03385(.dina(n3618), .dinb(n3610), .dout(n3619));
  jand g03386(.dina(n3619), .dinb(n194), .dout(n3620));
  jand g03387(.dina(n3614), .dinb(n3610), .dout(n3621));
  jor  g03388(.dina(n3615), .dinb(n3352), .dout(n3622));
  jand g03389(.dina(n3364), .dinb(n3352), .dout(n3623));
  jor  g03390(.dina(n3623), .dinb(n194), .dout(n3624));
  jnot g03391(.din(n3624), .dout(n3625));
  jand g03392(.dina(n3625), .dinb(n3622), .dout(n3626));
  jor  g03393(.dina(n3626), .dinb(n3621), .dout(n3629));
  jor  g03394(.dina(n3629), .dinb(n3620), .dout(asqrt[38] ));
  jand g03395(.dina(asqrt[38] ), .dinb(a[76] ), .dout(n3631));
  jnot g03396(.din(a[74] ), .dout(n3632));
  jnot g03397(.din(a[75] ), .dout(n3633));
  jand g03398(.dina(n3379), .dinb(n3633), .dout(n3634));
  jand g03399(.dina(n3634), .dinb(n3632), .dout(n3635));
  jor  g03400(.dina(n3635), .dinb(n3631), .dout(n3636));
  jand g03401(.dina(n3636), .dinb(asqrt[39] ), .dout(n3637));
  jand g03402(.dina(asqrt[38] ), .dinb(n3379), .dout(n3638));
  jxor g03403(.dina(n3638), .dinb(n3380), .dout(n3639));
  jor  g03404(.dina(n3636), .dinb(asqrt[39] ), .dout(n3640));
  jand g03405(.dina(n3640), .dinb(n3639), .dout(n3641));
  jor  g03406(.dina(n3641), .dinb(n3637), .dout(n3642));
  jand g03407(.dina(n3642), .dinb(asqrt[40] ), .dout(n3643));
  jor  g03408(.dina(n3637), .dinb(asqrt[40] ), .dout(n3644));
  jor  g03409(.dina(n3644), .dinb(n3641), .dout(n3645));
  jand g03410(.dina(n3638), .dinb(n3380), .dout(n3646));
  jnot g03411(.din(n3620), .dout(n3647));
  jnot g03412(.din(n3621), .dout(n3648));
  jnot g03413(.din(n3626), .dout(n3649));
  jand g03414(.dina(n3649), .dinb(asqrt[39] ), .dout(n3650));
  jand g03415(.dina(n3650), .dinb(n3648), .dout(n3651));
  jand g03416(.dina(n3651), .dinb(n3647), .dout(n3652));
  jor  g03417(.dina(n3652), .dinb(n3646), .dout(n3653));
  jxor g03418(.dina(n3653), .dinb(n3115), .dout(n3654));
  jand g03419(.dina(n3654), .dinb(n3645), .dout(n3655));
  jor  g03420(.dina(n3655), .dinb(n3643), .dout(n3656));
  jand g03421(.dina(n3656), .dinb(asqrt[41] ), .dout(n3657));
  jor  g03422(.dina(n3656), .dinb(asqrt[41] ), .dout(n3658));
  jxor g03423(.dina(n3384), .dinb(n3371), .dout(n3659));
  jand g03424(.dina(n3659), .dinb(asqrt[38] ), .dout(n3660));
  jxor g03425(.dina(n3660), .dinb(n3387), .dout(n3661));
  jnot g03426(.din(n3661), .dout(n3662));
  jand g03427(.dina(n3662), .dinb(n3658), .dout(n3663));
  jor  g03428(.dina(n3663), .dinb(n3657), .dout(n3664));
  jand g03429(.dina(n3664), .dinb(asqrt[42] ), .dout(n3665));
  jnot g03430(.din(n3393), .dout(n3666));
  jand g03431(.dina(n3666), .dinb(n3391), .dout(n3667));
  jand g03432(.dina(n3667), .dinb(asqrt[38] ), .dout(n3668));
  jxor g03433(.dina(n3668), .dinb(n3401), .dout(n3669));
  jnot g03434(.din(n3669), .dout(n3670));
  jor  g03435(.dina(n3657), .dinb(asqrt[42] ), .dout(n3671));
  jor  g03436(.dina(n3671), .dinb(n3663), .dout(n3672));
  jand g03437(.dina(n3672), .dinb(n3670), .dout(n3673));
  jor  g03438(.dina(n3673), .dinb(n3665), .dout(n3674));
  jand g03439(.dina(n3674), .dinb(asqrt[43] ), .dout(n3675));
  jor  g03440(.dina(n3674), .dinb(asqrt[43] ), .dout(n3676));
  jnot g03441(.din(n3408), .dout(n3677));
  jxor g03442(.dina(n3403), .dinb(n2870), .dout(n3678));
  jand g03443(.dina(n3678), .dinb(asqrt[38] ), .dout(n3679));
  jxor g03444(.dina(n3679), .dinb(n3677), .dout(n3680));
  jand g03445(.dina(n3680), .dinb(n3676), .dout(n3681));
  jor  g03446(.dina(n3681), .dinb(n3675), .dout(n3682));
  jand g03447(.dina(n3682), .dinb(asqrt[44] ), .dout(n3683));
  jor  g03448(.dina(n3675), .dinb(asqrt[44] ), .dout(n3684));
  jor  g03449(.dina(n3684), .dinb(n3681), .dout(n3685));
  jnot g03450(.din(n3415), .dout(n3686));
  jnot g03451(.din(n3417), .dout(n3687));
  jand g03452(.dina(asqrt[38] ), .dinb(n3411), .dout(n3688));
  jand g03453(.dina(n3688), .dinb(n3687), .dout(n3689));
  jor  g03454(.dina(n3689), .dinb(n3686), .dout(n3690));
  jnot g03455(.din(n3418), .dout(n3691));
  jand g03456(.dina(n3688), .dinb(n3691), .dout(n3692));
  jnot g03457(.din(n3692), .dout(n3693));
  jand g03458(.dina(n3693), .dinb(n3690), .dout(n3694));
  jand g03459(.dina(n3694), .dinb(n3685), .dout(n3695));
  jor  g03460(.dina(n3695), .dinb(n3683), .dout(n3696));
  jand g03461(.dina(n3696), .dinb(asqrt[45] ), .dout(n3697));
  jor  g03462(.dina(n3696), .dinb(asqrt[45] ), .dout(n3698));
  jxor g03463(.dina(n3419), .dinb(n2420), .dout(n3699));
  jand g03464(.dina(n3699), .dinb(asqrt[38] ), .dout(n3700));
  jxor g03465(.dina(n3700), .dinb(n3424), .dout(n3701));
  jand g03466(.dina(n3701), .dinb(n3698), .dout(n3702));
  jor  g03467(.dina(n3702), .dinb(n3697), .dout(n3703));
  jand g03468(.dina(n3703), .dinb(asqrt[46] ), .dout(n3704));
  jnot g03469(.din(n3430), .dout(n3705));
  jand g03470(.dina(n3705), .dinb(n3428), .dout(n3706));
  jand g03471(.dina(n3706), .dinb(asqrt[38] ), .dout(n3707));
  jxor g03472(.dina(n3707), .dinb(n3438), .dout(n3708));
  jnot g03473(.din(n3708), .dout(n3709));
  jor  g03474(.dina(n3697), .dinb(asqrt[46] ), .dout(n3710));
  jor  g03475(.dina(n3710), .dinb(n3702), .dout(n3711));
  jand g03476(.dina(n3711), .dinb(n3709), .dout(n3712));
  jor  g03477(.dina(n3712), .dinb(n3704), .dout(n3713));
  jand g03478(.dina(n3713), .dinb(asqrt[47] ), .dout(n3714));
  jor  g03479(.dina(n3713), .dinb(asqrt[47] ), .dout(n3715));
  jxor g03480(.dina(n3440), .dinb(n2005), .dout(n3716));
  jand g03481(.dina(n3716), .dinb(asqrt[38] ), .dout(n3717));
  jxor g03482(.dina(n3717), .dinb(n3446), .dout(n3718));
  jand g03483(.dina(n3718), .dinb(n3715), .dout(n3719));
  jor  g03484(.dina(n3719), .dinb(n3714), .dout(n3720));
  jand g03485(.dina(n3720), .dinb(asqrt[48] ), .dout(n3721));
  jor  g03486(.dina(n3714), .dinb(asqrt[48] ), .dout(n3722));
  jor  g03487(.dina(n3722), .dinb(n3719), .dout(n3723));
  jnot g03488(.din(n3454), .dout(n3724));
  jnot g03489(.din(n3456), .dout(n3725));
  jand g03490(.dina(asqrt[38] ), .dinb(n3450), .dout(n3726));
  jand g03491(.dina(n3726), .dinb(n3725), .dout(n3727));
  jor  g03492(.dina(n3727), .dinb(n3724), .dout(n3728));
  jnot g03493(.din(n3457), .dout(n3729));
  jand g03494(.dina(n3726), .dinb(n3729), .dout(n3730));
  jnot g03495(.din(n3730), .dout(n3731));
  jand g03496(.dina(n3731), .dinb(n3728), .dout(n3732));
  jand g03497(.dina(n3732), .dinb(n3723), .dout(n3733));
  jor  g03498(.dina(n3733), .dinb(n3721), .dout(n3734));
  jand g03499(.dina(n3734), .dinb(asqrt[49] ), .dout(n3735));
  jxor g03500(.dina(n3458), .dinb(n1641), .dout(n3736));
  jand g03501(.dina(n3736), .dinb(asqrt[38] ), .dout(n3737));
  jxor g03502(.dina(n3737), .dinb(n3465), .dout(n3738));
  jnot g03503(.din(n3738), .dout(n3739));
  jor  g03504(.dina(n3734), .dinb(asqrt[49] ), .dout(n3740));
  jand g03505(.dina(n3740), .dinb(n3739), .dout(n3741));
  jor  g03506(.dina(n3741), .dinb(n3735), .dout(n3742));
  jand g03507(.dina(n3742), .dinb(asqrt[50] ), .dout(n3743));
  jnot g03508(.din(n3470), .dout(n3744));
  jand g03509(.dina(n3744), .dinb(n3468), .dout(n3745));
  jand g03510(.dina(n3745), .dinb(asqrt[38] ), .dout(n3746));
  jxor g03511(.dina(n3746), .dinb(n3478), .dout(n3747));
  jnot g03512(.din(n3747), .dout(n3748));
  jor  g03513(.dina(n3735), .dinb(asqrt[50] ), .dout(n3749));
  jor  g03514(.dina(n3749), .dinb(n3741), .dout(n3750));
  jand g03515(.dina(n3750), .dinb(n3748), .dout(n3751));
  jor  g03516(.dina(n3751), .dinb(n3743), .dout(n3752));
  jand g03517(.dina(n3752), .dinb(asqrt[51] ), .dout(n3753));
  jor  g03518(.dina(n3752), .dinb(asqrt[51] ), .dout(n3754));
  jnot g03519(.din(n3484), .dout(n3755));
  jnot g03520(.din(n3485), .dout(n3756));
  jand g03521(.dina(asqrt[38] ), .dinb(n3481), .dout(n3757));
  jand g03522(.dina(n3757), .dinb(n3756), .dout(n3758));
  jor  g03523(.dina(n3758), .dinb(n3755), .dout(n3759));
  jnot g03524(.din(n3486), .dout(n3760));
  jand g03525(.dina(n3757), .dinb(n3760), .dout(n3761));
  jnot g03526(.din(n3761), .dout(n3762));
  jand g03527(.dina(n3762), .dinb(n3759), .dout(n3763));
  jand g03528(.dina(n3763), .dinb(n3754), .dout(n3764));
  jor  g03529(.dina(n3764), .dinb(n3753), .dout(n3765));
  jand g03530(.dina(n3765), .dinb(asqrt[52] ), .dout(n3766));
  jor  g03531(.dina(n3753), .dinb(asqrt[52] ), .dout(n3767));
  jor  g03532(.dina(n3767), .dinb(n3764), .dout(n3768));
  jnot g03533(.din(n3492), .dout(n3769));
  jnot g03534(.din(n3494), .dout(n3770));
  jand g03535(.dina(asqrt[38] ), .dinb(n3488), .dout(n3771));
  jand g03536(.dina(n3771), .dinb(n3770), .dout(n3772));
  jor  g03537(.dina(n3772), .dinb(n3769), .dout(n3773));
  jnot g03538(.din(n3495), .dout(n3774));
  jand g03539(.dina(n3771), .dinb(n3774), .dout(n3775));
  jnot g03540(.din(n3775), .dout(n3776));
  jand g03541(.dina(n3776), .dinb(n3773), .dout(n3777));
  jand g03542(.dina(n3777), .dinb(n3768), .dout(n3778));
  jor  g03543(.dina(n3778), .dinb(n3766), .dout(n3779));
  jand g03544(.dina(n3779), .dinb(asqrt[53] ), .dout(n3780));
  jxor g03545(.dina(n3496), .dinb(n1034), .dout(n3781));
  jand g03546(.dina(n3781), .dinb(asqrt[38] ), .dout(n3782));
  jxor g03547(.dina(n3782), .dinb(n3506), .dout(n3783));
  jnot g03548(.din(n3783), .dout(n3784));
  jor  g03549(.dina(n3779), .dinb(asqrt[53] ), .dout(n3785));
  jand g03550(.dina(n3785), .dinb(n3784), .dout(n3786));
  jor  g03551(.dina(n3786), .dinb(n3780), .dout(n3787));
  jand g03552(.dina(n3787), .dinb(asqrt[54] ), .dout(n3788));
  jnot g03553(.din(n3511), .dout(n3789));
  jand g03554(.dina(n3789), .dinb(n3509), .dout(n3790));
  jand g03555(.dina(n3790), .dinb(asqrt[38] ), .dout(n3791));
  jxor g03556(.dina(n3791), .dinb(n3519), .dout(n3792));
  jnot g03557(.din(n3792), .dout(n3793));
  jor  g03558(.dina(n3780), .dinb(asqrt[54] ), .dout(n3794));
  jor  g03559(.dina(n3794), .dinb(n3786), .dout(n3795));
  jand g03560(.dina(n3795), .dinb(n3793), .dout(n3796));
  jor  g03561(.dina(n3796), .dinb(n3788), .dout(n3797));
  jand g03562(.dina(n3797), .dinb(asqrt[55] ), .dout(n3798));
  jor  g03563(.dina(n3797), .dinb(asqrt[55] ), .dout(n3799));
  jnot g03564(.din(n3525), .dout(n3800));
  jnot g03565(.din(n3526), .dout(n3801));
  jand g03566(.dina(asqrt[38] ), .dinb(n3522), .dout(n3802));
  jand g03567(.dina(n3802), .dinb(n3801), .dout(n3803));
  jor  g03568(.dina(n3803), .dinb(n3800), .dout(n3804));
  jnot g03569(.din(n3527), .dout(n3805));
  jand g03570(.dina(n3802), .dinb(n3805), .dout(n3806));
  jnot g03571(.din(n3806), .dout(n3807));
  jand g03572(.dina(n3807), .dinb(n3804), .dout(n3808));
  jand g03573(.dina(n3808), .dinb(n3799), .dout(n3809));
  jor  g03574(.dina(n3809), .dinb(n3798), .dout(n3810));
  jand g03575(.dina(n3810), .dinb(asqrt[56] ), .dout(n3811));
  jor  g03576(.dina(n3798), .dinb(asqrt[56] ), .dout(n3812));
  jor  g03577(.dina(n3812), .dinb(n3809), .dout(n3813));
  jnot g03578(.din(n3533), .dout(n3814));
  jnot g03579(.din(n3535), .dout(n3815));
  jand g03580(.dina(asqrt[38] ), .dinb(n3529), .dout(n3816));
  jand g03581(.dina(n3816), .dinb(n3815), .dout(n3817));
  jor  g03582(.dina(n3817), .dinb(n3814), .dout(n3818));
  jnot g03583(.din(n3536), .dout(n3819));
  jand g03584(.dina(n3816), .dinb(n3819), .dout(n3820));
  jnot g03585(.din(n3820), .dout(n3821));
  jand g03586(.dina(n3821), .dinb(n3818), .dout(n3822));
  jand g03587(.dina(n3822), .dinb(n3813), .dout(n3823));
  jor  g03588(.dina(n3823), .dinb(n3811), .dout(n3824));
  jand g03589(.dina(n3824), .dinb(asqrt[57] ), .dout(n3825));
  jxor g03590(.dina(n3537), .dinb(n590), .dout(n3826));
  jand g03591(.dina(n3826), .dinb(asqrt[38] ), .dout(n3827));
  jxor g03592(.dina(n3827), .dinb(n3547), .dout(n3828));
  jnot g03593(.din(n3828), .dout(n3829));
  jor  g03594(.dina(n3824), .dinb(asqrt[57] ), .dout(n3830));
  jand g03595(.dina(n3830), .dinb(n3829), .dout(n3831));
  jor  g03596(.dina(n3831), .dinb(n3825), .dout(n3832));
  jand g03597(.dina(n3832), .dinb(asqrt[58] ), .dout(n3833));
  jnot g03598(.din(n3552), .dout(n3834));
  jand g03599(.dina(n3834), .dinb(n3550), .dout(n3835));
  jand g03600(.dina(n3835), .dinb(asqrt[38] ), .dout(n3836));
  jxor g03601(.dina(n3836), .dinb(n3560), .dout(n3837));
  jnot g03602(.din(n3837), .dout(n3838));
  jor  g03603(.dina(n3825), .dinb(asqrt[58] ), .dout(n3839));
  jor  g03604(.dina(n3839), .dinb(n3831), .dout(n3840));
  jand g03605(.dina(n3840), .dinb(n3838), .dout(n3841));
  jor  g03606(.dina(n3841), .dinb(n3833), .dout(n3842));
  jand g03607(.dina(n3842), .dinb(asqrt[59] ), .dout(n3843));
  jor  g03608(.dina(n3842), .dinb(asqrt[59] ), .dout(n3844));
  jnot g03609(.din(n3566), .dout(n3845));
  jnot g03610(.din(n3567), .dout(n3846));
  jand g03611(.dina(asqrt[38] ), .dinb(n3563), .dout(n3847));
  jand g03612(.dina(n3847), .dinb(n3846), .dout(n3848));
  jor  g03613(.dina(n3848), .dinb(n3845), .dout(n3849));
  jnot g03614(.din(n3568), .dout(n3850));
  jand g03615(.dina(n3847), .dinb(n3850), .dout(n3851));
  jnot g03616(.din(n3851), .dout(n3852));
  jand g03617(.dina(n3852), .dinb(n3849), .dout(n3853));
  jand g03618(.dina(n3853), .dinb(n3844), .dout(n3854));
  jor  g03619(.dina(n3854), .dinb(n3843), .dout(n3855));
  jand g03620(.dina(n3855), .dinb(asqrt[60] ), .dout(n3856));
  jor  g03621(.dina(n3843), .dinb(asqrt[60] ), .dout(n3857));
  jor  g03622(.dina(n3857), .dinb(n3854), .dout(n3858));
  jnot g03623(.din(n3574), .dout(n3859));
  jnot g03624(.din(n3576), .dout(n3860));
  jand g03625(.dina(asqrt[38] ), .dinb(n3570), .dout(n3861));
  jand g03626(.dina(n3861), .dinb(n3860), .dout(n3862));
  jor  g03627(.dina(n3862), .dinb(n3859), .dout(n3863));
  jnot g03628(.din(n3577), .dout(n3864));
  jand g03629(.dina(n3861), .dinb(n3864), .dout(n3865));
  jnot g03630(.din(n3865), .dout(n3866));
  jand g03631(.dina(n3866), .dinb(n3863), .dout(n3867));
  jand g03632(.dina(n3867), .dinb(n3858), .dout(n3868));
  jor  g03633(.dina(n3868), .dinb(n3856), .dout(n3869));
  jand g03634(.dina(n3869), .dinb(asqrt[61] ), .dout(n3870));
  jxor g03635(.dina(n3578), .dinb(n290), .dout(n3871));
  jand g03636(.dina(n3871), .dinb(asqrt[38] ), .dout(n3872));
  jxor g03637(.dina(n3872), .dinb(n3588), .dout(n3873));
  jnot g03638(.din(n3873), .dout(n3874));
  jor  g03639(.dina(n3869), .dinb(asqrt[61] ), .dout(n3875));
  jand g03640(.dina(n3875), .dinb(n3874), .dout(n3876));
  jor  g03641(.dina(n3876), .dinb(n3870), .dout(n3877));
  jand g03642(.dina(n3877), .dinb(asqrt[62] ), .dout(n3878));
  jnot g03643(.din(n3593), .dout(n3879));
  jand g03644(.dina(n3879), .dinb(n3591), .dout(n3880));
  jand g03645(.dina(n3880), .dinb(asqrt[38] ), .dout(n3881));
  jxor g03646(.dina(n3881), .dinb(n3601), .dout(n3882));
  jnot g03647(.din(n3882), .dout(n3883));
  jor  g03648(.dina(n3870), .dinb(asqrt[62] ), .dout(n3884));
  jor  g03649(.dina(n3884), .dinb(n3876), .dout(n3885));
  jand g03650(.dina(n3885), .dinb(n3883), .dout(n3886));
  jor  g03651(.dina(n3886), .dinb(n3878), .dout(n3887));
  jxor g03652(.dina(n3603), .dinb(n199), .dout(n3888));
  jand g03653(.dina(n3888), .dinb(asqrt[38] ), .dout(n3889));
  jxor g03654(.dina(n3889), .dinb(n3608), .dout(n3890));
  jnot g03655(.din(n3610), .dout(n3891));
  jnot g03656(.din(n3614), .dout(n3892));
  jand g03657(.dina(asqrt[38] ), .dinb(n3892), .dout(n3893));
  jand g03658(.dina(n3893), .dinb(n3891), .dout(n3894));
  jor  g03659(.dina(n3894), .dinb(n3621), .dout(n3895));
  jor  g03660(.dina(n3895), .dinb(n3890), .dout(n3896));
  jnot g03661(.din(n3896), .dout(n3897));
  jand g03662(.dina(n3897), .dinb(n3887), .dout(n3898));
  jor  g03663(.dina(n3898), .dinb(asqrt[63] ), .dout(n3899));
  jnot g03664(.din(n3890), .dout(n3900));
  jor  g03665(.dina(n3900), .dinb(n3887), .dout(n3901));
  jor  g03666(.dina(n3893), .dinb(n3891), .dout(n3902));
  jand g03667(.dina(n3892), .dinb(n3891), .dout(n3903));
  jor  g03668(.dina(n3903), .dinb(n194), .dout(n3904));
  jnot g03669(.din(n3904), .dout(n3905));
  jand g03670(.dina(n3905), .dinb(n3902), .dout(n3906));
  jnot g03671(.din(asqrt[38] ), .dout(n3907));
  jnot g03672(.din(n3906), .dout(n3910));
  jand g03673(.dina(n3910), .dinb(n3901), .dout(n3911));
  jand g03674(.dina(n3911), .dinb(n3899), .dout(n3912));
  jnot g03675(.din(n3912), .dout(asqrt[37] ));
  jor  g03676(.dina(n3912), .dinb(n3632), .dout(n3914));
  jnot g03677(.din(a[72] ), .dout(n3915));
  jnot g03678(.din(a[73] ), .dout(n3916));
  jand g03679(.dina(n3632), .dinb(n3916), .dout(n3917));
  jand g03680(.dina(n3917), .dinb(n3915), .dout(n3918));
  jnot g03681(.din(n3918), .dout(n3919));
  jand g03682(.dina(n3919), .dinb(n3914), .dout(n3920));
  jor  g03683(.dina(n3920), .dinb(n3907), .dout(n3921));
  jor  g03684(.dina(n3912), .dinb(a[74] ), .dout(n3922));
  jxor g03685(.dina(n3922), .dinb(n3633), .dout(n3923));
  jand g03686(.dina(n3920), .dinb(n3907), .dout(n3924));
  jor  g03687(.dina(n3924), .dinb(n3923), .dout(n3925));
  jand g03688(.dina(n3925), .dinb(n3921), .dout(n3926));
  jor  g03689(.dina(n3926), .dinb(n3376), .dout(n3927));
  jand g03690(.dina(n3921), .dinb(n3376), .dout(n3928));
  jand g03691(.dina(n3928), .dinb(n3925), .dout(n3929));
  jor  g03692(.dina(n3922), .dinb(a[75] ), .dout(n3930));
  jnot g03693(.din(n3899), .dout(n3931));
  jnot g03694(.din(n3901), .dout(n3932));
  jor  g03695(.dina(n3906), .dinb(n3907), .dout(n3933));
  jor  g03696(.dina(n3933), .dinb(n3932), .dout(n3934));
  jor  g03697(.dina(n3934), .dinb(n3931), .dout(n3935));
  jand g03698(.dina(n3935), .dinb(n3930), .dout(n3936));
  jxor g03699(.dina(n3936), .dinb(n3379), .dout(n3937));
  jor  g03700(.dina(n3937), .dinb(n3929), .dout(n3938));
  jand g03701(.dina(n3938), .dinb(n3927), .dout(n3939));
  jor  g03702(.dina(n3939), .dinb(n3371), .dout(n3940));
  jand g03703(.dina(n3939), .dinb(n3371), .dout(n3941));
  jxor g03704(.dina(n3636), .dinb(n3376), .dout(n3942));
  jor  g03705(.dina(n3942), .dinb(n3912), .dout(n3943));
  jxor g03706(.dina(n3943), .dinb(n3639), .dout(n3944));
  jor  g03707(.dina(n3944), .dinb(n3941), .dout(n3945));
  jand g03708(.dina(n3945), .dinb(n3940), .dout(n3946));
  jor  g03709(.dina(n3946), .dinb(n2875), .dout(n3947));
  jnot g03710(.din(n3645), .dout(n3948));
  jor  g03711(.dina(n3948), .dinb(n3643), .dout(n3949));
  jor  g03712(.dina(n3949), .dinb(n3912), .dout(n3950));
  jxor g03713(.dina(n3950), .dinb(n3654), .dout(n3951));
  jand g03714(.dina(n3940), .dinb(n2875), .dout(n3952));
  jand g03715(.dina(n3952), .dinb(n3945), .dout(n3953));
  jor  g03716(.dina(n3953), .dinb(n3951), .dout(n3954));
  jand g03717(.dina(n3954), .dinb(n3947), .dout(n3955));
  jor  g03718(.dina(n3955), .dinb(n2870), .dout(n3956));
  jand g03719(.dina(n3955), .dinb(n2870), .dout(n3957));
  jxor g03720(.dina(n3656), .dinb(n2875), .dout(n3958));
  jor  g03721(.dina(n3958), .dinb(n3912), .dout(n3959));
  jxor g03722(.dina(n3959), .dinb(n3661), .dout(n3960));
  jnot g03723(.din(n3960), .dout(n3961));
  jor  g03724(.dina(n3961), .dinb(n3957), .dout(n3962));
  jand g03725(.dina(n3962), .dinb(n3956), .dout(n3963));
  jor  g03726(.dina(n3963), .dinb(n2425), .dout(n3964));
  jand g03727(.dina(n3956), .dinb(n2425), .dout(n3965));
  jand g03728(.dina(n3965), .dinb(n3962), .dout(n3966));
  jnot g03729(.din(n3665), .dout(n3967));
  jand g03730(.dina(asqrt[37] ), .dinb(n3967), .dout(n3968));
  jand g03731(.dina(n3968), .dinb(n3672), .dout(n3969));
  jor  g03732(.dina(n3969), .dinb(n3670), .dout(n3970));
  jand g03733(.dina(n3968), .dinb(n3673), .dout(n3971));
  jnot g03734(.din(n3971), .dout(n3972));
  jand g03735(.dina(n3972), .dinb(n3970), .dout(n3973));
  jnot g03736(.din(n3973), .dout(n3974));
  jor  g03737(.dina(n3974), .dinb(n3966), .dout(n3975));
  jand g03738(.dina(n3975), .dinb(n3964), .dout(n3976));
  jor  g03739(.dina(n3976), .dinb(n2420), .dout(n3977));
  jand g03740(.dina(n3976), .dinb(n2420), .dout(n3978));
  jnot g03741(.din(n3680), .dout(n3979));
  jxor g03742(.dina(n3674), .dinb(n2425), .dout(n3980));
  jor  g03743(.dina(n3980), .dinb(n3912), .dout(n3981));
  jxor g03744(.dina(n3981), .dinb(n3979), .dout(n3982));
  jnot g03745(.din(n3982), .dout(n3983));
  jor  g03746(.dina(n3983), .dinb(n3978), .dout(n3984));
  jand g03747(.dina(n3984), .dinb(n3977), .dout(n3985));
  jor  g03748(.dina(n3985), .dinb(n2010), .dout(n3986));
  jnot g03749(.din(n3685), .dout(n3987));
  jor  g03750(.dina(n3987), .dinb(n3683), .dout(n3988));
  jor  g03751(.dina(n3988), .dinb(n3912), .dout(n3989));
  jxor g03752(.dina(n3989), .dinb(n3694), .dout(n3990));
  jand g03753(.dina(n3977), .dinb(n2010), .dout(n3991));
  jand g03754(.dina(n3991), .dinb(n3984), .dout(n3992));
  jor  g03755(.dina(n3992), .dinb(n3990), .dout(n3993));
  jand g03756(.dina(n3993), .dinb(n3986), .dout(n3994));
  jor  g03757(.dina(n3994), .dinb(n2005), .dout(n3995));
  jand g03758(.dina(n3994), .dinb(n2005), .dout(n3996));
  jnot g03759(.din(n3701), .dout(n3997));
  jxor g03760(.dina(n3696), .dinb(n2010), .dout(n3998));
  jor  g03761(.dina(n3998), .dinb(n3912), .dout(n3999));
  jxor g03762(.dina(n3999), .dinb(n3997), .dout(n4000));
  jnot g03763(.din(n4000), .dout(n4001));
  jor  g03764(.dina(n4001), .dinb(n3996), .dout(n4002));
  jand g03765(.dina(n4002), .dinb(n3995), .dout(n4003));
  jor  g03766(.dina(n4003), .dinb(n1646), .dout(n4004));
  jand g03767(.dina(n3995), .dinb(n1646), .dout(n4005));
  jand g03768(.dina(n4005), .dinb(n4002), .dout(n4006));
  jnot g03769(.din(n3704), .dout(n4007));
  jand g03770(.dina(asqrt[37] ), .dinb(n4007), .dout(n4008));
  jand g03771(.dina(n4008), .dinb(n3711), .dout(n4009));
  jor  g03772(.dina(n4009), .dinb(n3709), .dout(n4010));
  jand g03773(.dina(n4008), .dinb(n3712), .dout(n4011));
  jnot g03774(.din(n4011), .dout(n4012));
  jand g03775(.dina(n4012), .dinb(n4010), .dout(n4013));
  jnot g03776(.din(n4013), .dout(n4014));
  jor  g03777(.dina(n4014), .dinb(n4006), .dout(n4015));
  jand g03778(.dina(n4015), .dinb(n4004), .dout(n4016));
  jor  g03779(.dina(n4016), .dinb(n1641), .dout(n4017));
  jxor g03780(.dina(n3713), .dinb(n1646), .dout(n4018));
  jor  g03781(.dina(n4018), .dinb(n3912), .dout(n4019));
  jxor g03782(.dina(n4019), .dinb(n3718), .dout(n4020));
  jand g03783(.dina(n4016), .dinb(n1641), .dout(n4021));
  jor  g03784(.dina(n4021), .dinb(n4020), .dout(n4022));
  jand g03785(.dina(n4022), .dinb(n4017), .dout(n4023));
  jor  g03786(.dina(n4023), .dinb(n1317), .dout(n4024));
  jnot g03787(.din(n3723), .dout(n4025));
  jor  g03788(.dina(n4025), .dinb(n3721), .dout(n4026));
  jor  g03789(.dina(n4026), .dinb(n3912), .dout(n4027));
  jxor g03790(.dina(n4027), .dinb(n3732), .dout(n4028));
  jand g03791(.dina(n4017), .dinb(n1317), .dout(n4029));
  jand g03792(.dina(n4029), .dinb(n4022), .dout(n4030));
  jor  g03793(.dina(n4030), .dinb(n4028), .dout(n4031));
  jand g03794(.dina(n4031), .dinb(n4024), .dout(n4032));
  jor  g03795(.dina(n4032), .dinb(n1312), .dout(n4033));
  jand g03796(.dina(n4032), .dinb(n1312), .dout(n4034));
  jnot g03797(.din(n3735), .dout(n4035));
  jand g03798(.dina(asqrt[37] ), .dinb(n4035), .dout(n4036));
  jand g03799(.dina(n4036), .dinb(n3740), .dout(n4037));
  jor  g03800(.dina(n4037), .dinb(n3739), .dout(n4038));
  jand g03801(.dina(n4036), .dinb(n3741), .dout(n4039));
  jnot g03802(.din(n4039), .dout(n4040));
  jand g03803(.dina(n4040), .dinb(n4038), .dout(n4041));
  jnot g03804(.din(n4041), .dout(n4042));
  jor  g03805(.dina(n4042), .dinb(n4034), .dout(n4043));
  jand g03806(.dina(n4043), .dinb(n4033), .dout(n4044));
  jor  g03807(.dina(n4044), .dinb(n1039), .dout(n4045));
  jand g03808(.dina(n4033), .dinb(n1039), .dout(n4046));
  jand g03809(.dina(n4046), .dinb(n4043), .dout(n4047));
  jnot g03810(.din(n3743), .dout(n4048));
  jand g03811(.dina(asqrt[37] ), .dinb(n4048), .dout(n4049));
  jand g03812(.dina(n4049), .dinb(n3750), .dout(n4050));
  jor  g03813(.dina(n4050), .dinb(n3748), .dout(n4051));
  jand g03814(.dina(n4049), .dinb(n3751), .dout(n4052));
  jnot g03815(.din(n4052), .dout(n4053));
  jand g03816(.dina(n4053), .dinb(n4051), .dout(n4054));
  jnot g03817(.din(n4054), .dout(n4055));
  jor  g03818(.dina(n4055), .dinb(n4047), .dout(n4056));
  jand g03819(.dina(n4056), .dinb(n4045), .dout(n4057));
  jor  g03820(.dina(n4057), .dinb(n1034), .dout(n4058));
  jxor g03821(.dina(n3752), .dinb(n1039), .dout(n4059));
  jor  g03822(.dina(n4059), .dinb(n3912), .dout(n4060));
  jxor g03823(.dina(n4060), .dinb(n3763), .dout(n4061));
  jand g03824(.dina(n4057), .dinb(n1034), .dout(n4062));
  jor  g03825(.dina(n4062), .dinb(n4061), .dout(n4063));
  jand g03826(.dina(n4063), .dinb(n4058), .dout(n4064));
  jor  g03827(.dina(n4064), .dinb(n796), .dout(n4065));
  jnot g03828(.din(n3768), .dout(n4066));
  jor  g03829(.dina(n4066), .dinb(n3766), .dout(n4067));
  jor  g03830(.dina(n4067), .dinb(n3912), .dout(n4068));
  jxor g03831(.dina(n4068), .dinb(n3777), .dout(n4069));
  jand g03832(.dina(n4058), .dinb(n796), .dout(n4070));
  jand g03833(.dina(n4070), .dinb(n4063), .dout(n4071));
  jor  g03834(.dina(n4071), .dinb(n4069), .dout(n4072));
  jand g03835(.dina(n4072), .dinb(n4065), .dout(n4073));
  jor  g03836(.dina(n4073), .dinb(n791), .dout(n4074));
  jand g03837(.dina(n4073), .dinb(n791), .dout(n4075));
  jnot g03838(.din(n3780), .dout(n4076));
  jand g03839(.dina(asqrt[37] ), .dinb(n4076), .dout(n4077));
  jand g03840(.dina(n4077), .dinb(n3785), .dout(n4078));
  jor  g03841(.dina(n4078), .dinb(n3784), .dout(n4079));
  jand g03842(.dina(n4077), .dinb(n3786), .dout(n4080));
  jnot g03843(.din(n4080), .dout(n4081));
  jand g03844(.dina(n4081), .dinb(n4079), .dout(n4082));
  jnot g03845(.din(n4082), .dout(n4083));
  jor  g03846(.dina(n4083), .dinb(n4075), .dout(n4084));
  jand g03847(.dina(n4084), .dinb(n4074), .dout(n4085));
  jor  g03848(.dina(n4085), .dinb(n595), .dout(n4086));
  jand g03849(.dina(n4074), .dinb(n595), .dout(n4087));
  jand g03850(.dina(n4087), .dinb(n4084), .dout(n4088));
  jnot g03851(.din(n3788), .dout(n4089));
  jand g03852(.dina(asqrt[37] ), .dinb(n4089), .dout(n4090));
  jand g03853(.dina(n4090), .dinb(n3795), .dout(n4091));
  jor  g03854(.dina(n4091), .dinb(n3793), .dout(n4092));
  jand g03855(.dina(n4090), .dinb(n3796), .dout(n4093));
  jnot g03856(.din(n4093), .dout(n4094));
  jand g03857(.dina(n4094), .dinb(n4092), .dout(n4095));
  jnot g03858(.din(n4095), .dout(n4096));
  jor  g03859(.dina(n4096), .dinb(n4088), .dout(n4097));
  jand g03860(.dina(n4097), .dinb(n4086), .dout(n4098));
  jor  g03861(.dina(n4098), .dinb(n590), .dout(n4099));
  jxor g03862(.dina(n3797), .dinb(n595), .dout(n4100));
  jor  g03863(.dina(n4100), .dinb(n3912), .dout(n4101));
  jxor g03864(.dina(n4101), .dinb(n3808), .dout(n4102));
  jand g03865(.dina(n4098), .dinb(n590), .dout(n4103));
  jor  g03866(.dina(n4103), .dinb(n4102), .dout(n4104));
  jand g03867(.dina(n4104), .dinb(n4099), .dout(n4105));
  jor  g03868(.dina(n4105), .dinb(n430), .dout(n4106));
  jnot g03869(.din(n3813), .dout(n4107));
  jor  g03870(.dina(n4107), .dinb(n3811), .dout(n4108));
  jor  g03871(.dina(n4108), .dinb(n3912), .dout(n4109));
  jxor g03872(.dina(n4109), .dinb(n3822), .dout(n4110));
  jand g03873(.dina(n4099), .dinb(n430), .dout(n4111));
  jand g03874(.dina(n4111), .dinb(n4104), .dout(n4112));
  jor  g03875(.dina(n4112), .dinb(n4110), .dout(n4113));
  jand g03876(.dina(n4113), .dinb(n4106), .dout(n4114));
  jor  g03877(.dina(n4114), .dinb(n425), .dout(n4115));
  jand g03878(.dina(n4114), .dinb(n425), .dout(n4116));
  jnot g03879(.din(n3825), .dout(n4117));
  jand g03880(.dina(asqrt[37] ), .dinb(n4117), .dout(n4118));
  jand g03881(.dina(n4118), .dinb(n3830), .dout(n4119));
  jor  g03882(.dina(n4119), .dinb(n3829), .dout(n4120));
  jand g03883(.dina(n4118), .dinb(n3831), .dout(n4121));
  jnot g03884(.din(n4121), .dout(n4122));
  jand g03885(.dina(n4122), .dinb(n4120), .dout(n4123));
  jnot g03886(.din(n4123), .dout(n4124));
  jor  g03887(.dina(n4124), .dinb(n4116), .dout(n4125));
  jand g03888(.dina(n4125), .dinb(n4115), .dout(n4126));
  jor  g03889(.dina(n4126), .dinb(n305), .dout(n4127));
  jand g03890(.dina(n4115), .dinb(n305), .dout(n4128));
  jand g03891(.dina(n4128), .dinb(n4125), .dout(n4129));
  jnot g03892(.din(n3833), .dout(n4130));
  jand g03893(.dina(asqrt[37] ), .dinb(n4130), .dout(n4131));
  jand g03894(.dina(n4131), .dinb(n3840), .dout(n4132));
  jor  g03895(.dina(n4132), .dinb(n3838), .dout(n4133));
  jand g03896(.dina(n4131), .dinb(n3841), .dout(n4134));
  jnot g03897(.din(n4134), .dout(n4135));
  jand g03898(.dina(n4135), .dinb(n4133), .dout(n4136));
  jnot g03899(.din(n4136), .dout(n4137));
  jor  g03900(.dina(n4137), .dinb(n4129), .dout(n4138));
  jand g03901(.dina(n4138), .dinb(n4127), .dout(n4139));
  jor  g03902(.dina(n4139), .dinb(n290), .dout(n4140));
  jxor g03903(.dina(n3842), .dinb(n305), .dout(n4141));
  jor  g03904(.dina(n4141), .dinb(n3912), .dout(n4142));
  jxor g03905(.dina(n4142), .dinb(n3853), .dout(n4143));
  jand g03906(.dina(n4139), .dinb(n290), .dout(n4144));
  jor  g03907(.dina(n4144), .dinb(n4143), .dout(n4145));
  jand g03908(.dina(n4145), .dinb(n4140), .dout(n4146));
  jor  g03909(.dina(n4146), .dinb(n223), .dout(n4147));
  jnot g03910(.din(n3858), .dout(n4148));
  jor  g03911(.dina(n4148), .dinb(n3856), .dout(n4149));
  jor  g03912(.dina(n4149), .dinb(n3912), .dout(n4150));
  jxor g03913(.dina(n4150), .dinb(n3867), .dout(n4151));
  jand g03914(.dina(n4140), .dinb(n223), .dout(n4152));
  jand g03915(.dina(n4152), .dinb(n4145), .dout(n4153));
  jor  g03916(.dina(n4153), .dinb(n4151), .dout(n4154));
  jand g03917(.dina(n4154), .dinb(n4147), .dout(n4155));
  jor  g03918(.dina(n4155), .dinb(n199), .dout(n4156));
  jand g03919(.dina(n4155), .dinb(n199), .dout(n4157));
  jnot g03920(.din(n3870), .dout(n4158));
  jand g03921(.dina(asqrt[37] ), .dinb(n4158), .dout(n4159));
  jand g03922(.dina(n4159), .dinb(n3875), .dout(n4160));
  jor  g03923(.dina(n4160), .dinb(n3874), .dout(n4161));
  jand g03924(.dina(n4159), .dinb(n3876), .dout(n4162));
  jnot g03925(.din(n4162), .dout(n4163));
  jand g03926(.dina(n4163), .dinb(n4161), .dout(n4164));
  jnot g03927(.din(n4164), .dout(n4165));
  jor  g03928(.dina(n4165), .dinb(n4157), .dout(n4166));
  jand g03929(.dina(n4166), .dinb(n4156), .dout(n4167));
  jnot g03930(.din(n3878), .dout(n4168));
  jand g03931(.dina(asqrt[37] ), .dinb(n4168), .dout(n4169));
  jand g03932(.dina(n4169), .dinb(n3885), .dout(n4170));
  jor  g03933(.dina(n4170), .dinb(n3883), .dout(n4171));
  jand g03934(.dina(n4169), .dinb(n3886), .dout(n4172));
  jnot g03935(.din(n4172), .dout(n4173));
  jand g03936(.dina(n4173), .dinb(n4171), .dout(n4174));
  jnot g03937(.din(n4174), .dout(n4175));
  jand g03938(.dina(asqrt[37] ), .dinb(n3900), .dout(n4176));
  jand g03939(.dina(n4176), .dinb(n3887), .dout(n4177));
  jor  g03940(.dina(n4177), .dinb(n3932), .dout(n4178));
  jor  g03941(.dina(n4178), .dinb(n4175), .dout(n4179));
  jor  g03942(.dina(n4179), .dinb(n4167), .dout(n4180));
  jand g03943(.dina(n4180), .dinb(n194), .dout(n4181));
  jand g03944(.dina(n4175), .dinb(n4167), .dout(n4182));
  jor  g03945(.dina(n4176), .dinb(n3887), .dout(n4183));
  jand g03946(.dina(n3900), .dinb(n3887), .dout(n4184));
  jor  g03947(.dina(n4184), .dinb(n194), .dout(n4185));
  jnot g03948(.din(n4185), .dout(n4186));
  jand g03949(.dina(n4186), .dinb(n4183), .dout(n4187));
  jor  g03950(.dina(n4187), .dinb(n4182), .dout(n4190));
  jor  g03951(.dina(n4190), .dinb(n4181), .dout(asqrt[36] ));
  jand g03952(.dina(asqrt[36] ), .dinb(a[72] ), .dout(n4192));
  jnot g03953(.din(a[70] ), .dout(n4193));
  jnot g03954(.din(a[71] ), .dout(n4194));
  jand g03955(.dina(n3915), .dinb(n4194), .dout(n4195));
  jand g03956(.dina(n4195), .dinb(n4193), .dout(n4196));
  jor  g03957(.dina(n4196), .dinb(n4192), .dout(n4197));
  jand g03958(.dina(n4197), .dinb(asqrt[37] ), .dout(n4198));
  jand g03959(.dina(asqrt[36] ), .dinb(n3915), .dout(n4199));
  jxor g03960(.dina(n4199), .dinb(n3916), .dout(n4200));
  jor  g03961(.dina(n4197), .dinb(asqrt[37] ), .dout(n4201));
  jand g03962(.dina(n4201), .dinb(n4200), .dout(n4202));
  jor  g03963(.dina(n4202), .dinb(n4198), .dout(n4203));
  jand g03964(.dina(n4203), .dinb(asqrt[38] ), .dout(n4204));
  jor  g03965(.dina(n4198), .dinb(asqrt[38] ), .dout(n4205));
  jor  g03966(.dina(n4205), .dinb(n4202), .dout(n4206));
  jand g03967(.dina(n4199), .dinb(n3916), .dout(n4207));
  jnot g03968(.din(n4181), .dout(n4208));
  jnot g03969(.din(n4182), .dout(n4209));
  jnot g03970(.din(n4187), .dout(n4210));
  jand g03971(.dina(n4210), .dinb(asqrt[37] ), .dout(n4211));
  jand g03972(.dina(n4211), .dinb(n4209), .dout(n4212));
  jand g03973(.dina(n4212), .dinb(n4208), .dout(n4213));
  jor  g03974(.dina(n4213), .dinb(n4207), .dout(n4214));
  jxor g03975(.dina(n4214), .dinb(n3632), .dout(n4215));
  jand g03976(.dina(n4215), .dinb(n4206), .dout(n4216));
  jor  g03977(.dina(n4216), .dinb(n4204), .dout(n4217));
  jand g03978(.dina(n4217), .dinb(asqrt[39] ), .dout(n4218));
  jor  g03979(.dina(n4217), .dinb(asqrt[39] ), .dout(n4219));
  jxor g03980(.dina(n3920), .dinb(n3907), .dout(n4220));
  jand g03981(.dina(n4220), .dinb(asqrt[36] ), .dout(n4221));
  jxor g03982(.dina(n4221), .dinb(n3923), .dout(n4222));
  jnot g03983(.din(n4222), .dout(n4223));
  jand g03984(.dina(n4223), .dinb(n4219), .dout(n4224));
  jor  g03985(.dina(n4224), .dinb(n4218), .dout(n4225));
  jand g03986(.dina(n4225), .dinb(asqrt[40] ), .dout(n4226));
  jnot g03987(.din(n3929), .dout(n4227));
  jand g03988(.dina(n4227), .dinb(n3927), .dout(n4228));
  jand g03989(.dina(n4228), .dinb(asqrt[36] ), .dout(n4229));
  jxor g03990(.dina(n4229), .dinb(n3937), .dout(n4230));
  jnot g03991(.din(n4230), .dout(n4231));
  jor  g03992(.dina(n4218), .dinb(asqrt[40] ), .dout(n4232));
  jor  g03993(.dina(n4232), .dinb(n4224), .dout(n4233));
  jand g03994(.dina(n4233), .dinb(n4231), .dout(n4234));
  jor  g03995(.dina(n4234), .dinb(n4226), .dout(n4235));
  jand g03996(.dina(n4235), .dinb(asqrt[41] ), .dout(n4236));
  jor  g03997(.dina(n4235), .dinb(asqrt[41] ), .dout(n4237));
  jnot g03998(.din(n3944), .dout(n4238));
  jxor g03999(.dina(n3939), .dinb(n3371), .dout(n4239));
  jand g04000(.dina(n4239), .dinb(asqrt[36] ), .dout(n4240));
  jxor g04001(.dina(n4240), .dinb(n4238), .dout(n4241));
  jand g04002(.dina(n4241), .dinb(n4237), .dout(n4242));
  jor  g04003(.dina(n4242), .dinb(n4236), .dout(n4243));
  jand g04004(.dina(n4243), .dinb(asqrt[42] ), .dout(n4244));
  jor  g04005(.dina(n4236), .dinb(asqrt[42] ), .dout(n4245));
  jor  g04006(.dina(n4245), .dinb(n4242), .dout(n4246));
  jnot g04007(.din(n3951), .dout(n4247));
  jnot g04008(.din(n3953), .dout(n4248));
  jand g04009(.dina(asqrt[36] ), .dinb(n3947), .dout(n4249));
  jand g04010(.dina(n4249), .dinb(n4248), .dout(n4250));
  jor  g04011(.dina(n4250), .dinb(n4247), .dout(n4251));
  jnot g04012(.din(n3954), .dout(n4252));
  jand g04013(.dina(n4249), .dinb(n4252), .dout(n4253));
  jnot g04014(.din(n4253), .dout(n4254));
  jand g04015(.dina(n4254), .dinb(n4251), .dout(n4255));
  jand g04016(.dina(n4255), .dinb(n4246), .dout(n4256));
  jor  g04017(.dina(n4256), .dinb(n4244), .dout(n4257));
  jand g04018(.dina(n4257), .dinb(asqrt[43] ), .dout(n4258));
  jor  g04019(.dina(n4257), .dinb(asqrt[43] ), .dout(n4259));
  jxor g04020(.dina(n3955), .dinb(n2870), .dout(n4260));
  jand g04021(.dina(n4260), .dinb(asqrt[36] ), .dout(n4261));
  jxor g04022(.dina(n4261), .dinb(n3960), .dout(n4262));
  jand g04023(.dina(n4262), .dinb(n4259), .dout(n4263));
  jor  g04024(.dina(n4263), .dinb(n4258), .dout(n4264));
  jand g04025(.dina(n4264), .dinb(asqrt[44] ), .dout(n4265));
  jnot g04026(.din(n3966), .dout(n4266));
  jand g04027(.dina(n4266), .dinb(n3964), .dout(n4267));
  jand g04028(.dina(n4267), .dinb(asqrt[36] ), .dout(n4268));
  jxor g04029(.dina(n4268), .dinb(n3974), .dout(n4269));
  jnot g04030(.din(n4269), .dout(n4270));
  jor  g04031(.dina(n4258), .dinb(asqrt[44] ), .dout(n4271));
  jor  g04032(.dina(n4271), .dinb(n4263), .dout(n4272));
  jand g04033(.dina(n4272), .dinb(n4270), .dout(n4273));
  jor  g04034(.dina(n4273), .dinb(n4265), .dout(n4274));
  jand g04035(.dina(n4274), .dinb(asqrt[45] ), .dout(n4275));
  jor  g04036(.dina(n4274), .dinb(asqrt[45] ), .dout(n4276));
  jxor g04037(.dina(n3976), .dinb(n2420), .dout(n4277));
  jand g04038(.dina(n4277), .dinb(asqrt[36] ), .dout(n4278));
  jxor g04039(.dina(n4278), .dinb(n3982), .dout(n4279));
  jand g04040(.dina(n4279), .dinb(n4276), .dout(n4280));
  jor  g04041(.dina(n4280), .dinb(n4275), .dout(n4281));
  jand g04042(.dina(n4281), .dinb(asqrt[46] ), .dout(n4282));
  jor  g04043(.dina(n4275), .dinb(asqrt[46] ), .dout(n4283));
  jor  g04044(.dina(n4283), .dinb(n4280), .dout(n4284));
  jnot g04045(.din(n3990), .dout(n4285));
  jnot g04046(.din(n3992), .dout(n4286));
  jand g04047(.dina(asqrt[36] ), .dinb(n3986), .dout(n4287));
  jand g04048(.dina(n4287), .dinb(n4286), .dout(n4288));
  jor  g04049(.dina(n4288), .dinb(n4285), .dout(n4289));
  jnot g04050(.din(n3993), .dout(n4290));
  jand g04051(.dina(n4287), .dinb(n4290), .dout(n4291));
  jnot g04052(.din(n4291), .dout(n4292));
  jand g04053(.dina(n4292), .dinb(n4289), .dout(n4293));
  jand g04054(.dina(n4293), .dinb(n4284), .dout(n4294));
  jor  g04055(.dina(n4294), .dinb(n4282), .dout(n4295));
  jand g04056(.dina(n4295), .dinb(asqrt[47] ), .dout(n4296));
  jxor g04057(.dina(n3994), .dinb(n2005), .dout(n4297));
  jand g04058(.dina(n4297), .dinb(asqrt[36] ), .dout(n4298));
  jxor g04059(.dina(n4298), .dinb(n4001), .dout(n4299));
  jnot g04060(.din(n4299), .dout(n4300));
  jor  g04061(.dina(n4295), .dinb(asqrt[47] ), .dout(n4301));
  jand g04062(.dina(n4301), .dinb(n4300), .dout(n4302));
  jor  g04063(.dina(n4302), .dinb(n4296), .dout(n4303));
  jand g04064(.dina(n4303), .dinb(asqrt[48] ), .dout(n4304));
  jnot g04065(.din(n4006), .dout(n4305));
  jand g04066(.dina(n4305), .dinb(n4004), .dout(n4306));
  jand g04067(.dina(n4306), .dinb(asqrt[36] ), .dout(n4307));
  jxor g04068(.dina(n4307), .dinb(n4014), .dout(n4308));
  jnot g04069(.din(n4308), .dout(n4309));
  jor  g04070(.dina(n4296), .dinb(asqrt[48] ), .dout(n4310));
  jor  g04071(.dina(n4310), .dinb(n4302), .dout(n4311));
  jand g04072(.dina(n4311), .dinb(n4309), .dout(n4312));
  jor  g04073(.dina(n4312), .dinb(n4304), .dout(n4313));
  jand g04074(.dina(n4313), .dinb(asqrt[49] ), .dout(n4314));
  jor  g04075(.dina(n4313), .dinb(asqrt[49] ), .dout(n4315));
  jnot g04076(.din(n4020), .dout(n4316));
  jnot g04077(.din(n4021), .dout(n4317));
  jand g04078(.dina(asqrt[36] ), .dinb(n4017), .dout(n4318));
  jand g04079(.dina(n4318), .dinb(n4317), .dout(n4319));
  jor  g04080(.dina(n4319), .dinb(n4316), .dout(n4320));
  jnot g04081(.din(n4022), .dout(n4321));
  jand g04082(.dina(n4318), .dinb(n4321), .dout(n4322));
  jnot g04083(.din(n4322), .dout(n4323));
  jand g04084(.dina(n4323), .dinb(n4320), .dout(n4324));
  jand g04085(.dina(n4324), .dinb(n4315), .dout(n4325));
  jor  g04086(.dina(n4325), .dinb(n4314), .dout(n4326));
  jand g04087(.dina(n4326), .dinb(asqrt[50] ), .dout(n4327));
  jor  g04088(.dina(n4314), .dinb(asqrt[50] ), .dout(n4328));
  jor  g04089(.dina(n4328), .dinb(n4325), .dout(n4329));
  jnot g04090(.din(n4028), .dout(n4330));
  jnot g04091(.din(n4030), .dout(n4331));
  jand g04092(.dina(asqrt[36] ), .dinb(n4024), .dout(n4332));
  jand g04093(.dina(n4332), .dinb(n4331), .dout(n4333));
  jor  g04094(.dina(n4333), .dinb(n4330), .dout(n4334));
  jnot g04095(.din(n4031), .dout(n4335));
  jand g04096(.dina(n4332), .dinb(n4335), .dout(n4336));
  jnot g04097(.din(n4336), .dout(n4337));
  jand g04098(.dina(n4337), .dinb(n4334), .dout(n4338));
  jand g04099(.dina(n4338), .dinb(n4329), .dout(n4339));
  jor  g04100(.dina(n4339), .dinb(n4327), .dout(n4340));
  jand g04101(.dina(n4340), .dinb(asqrt[51] ), .dout(n4341));
  jxor g04102(.dina(n4032), .dinb(n1312), .dout(n4342));
  jand g04103(.dina(n4342), .dinb(asqrt[36] ), .dout(n4343));
  jxor g04104(.dina(n4343), .dinb(n4042), .dout(n4344));
  jnot g04105(.din(n4344), .dout(n4345));
  jor  g04106(.dina(n4340), .dinb(asqrt[51] ), .dout(n4346));
  jand g04107(.dina(n4346), .dinb(n4345), .dout(n4347));
  jor  g04108(.dina(n4347), .dinb(n4341), .dout(n4348));
  jand g04109(.dina(n4348), .dinb(asqrt[52] ), .dout(n4349));
  jnot g04110(.din(n4047), .dout(n4350));
  jand g04111(.dina(n4350), .dinb(n4045), .dout(n4351));
  jand g04112(.dina(n4351), .dinb(asqrt[36] ), .dout(n4352));
  jxor g04113(.dina(n4352), .dinb(n4055), .dout(n4353));
  jnot g04114(.din(n4353), .dout(n4354));
  jor  g04115(.dina(n4341), .dinb(asqrt[52] ), .dout(n4355));
  jor  g04116(.dina(n4355), .dinb(n4347), .dout(n4356));
  jand g04117(.dina(n4356), .dinb(n4354), .dout(n4357));
  jor  g04118(.dina(n4357), .dinb(n4349), .dout(n4358));
  jand g04119(.dina(n4358), .dinb(asqrt[53] ), .dout(n4359));
  jor  g04120(.dina(n4358), .dinb(asqrt[53] ), .dout(n4360));
  jnot g04121(.din(n4061), .dout(n4361));
  jnot g04122(.din(n4062), .dout(n4362));
  jand g04123(.dina(asqrt[36] ), .dinb(n4058), .dout(n4363));
  jand g04124(.dina(n4363), .dinb(n4362), .dout(n4364));
  jor  g04125(.dina(n4364), .dinb(n4361), .dout(n4365));
  jnot g04126(.din(n4063), .dout(n4366));
  jand g04127(.dina(n4363), .dinb(n4366), .dout(n4367));
  jnot g04128(.din(n4367), .dout(n4368));
  jand g04129(.dina(n4368), .dinb(n4365), .dout(n4369));
  jand g04130(.dina(n4369), .dinb(n4360), .dout(n4370));
  jor  g04131(.dina(n4370), .dinb(n4359), .dout(n4371));
  jand g04132(.dina(n4371), .dinb(asqrt[54] ), .dout(n4372));
  jor  g04133(.dina(n4359), .dinb(asqrt[54] ), .dout(n4373));
  jor  g04134(.dina(n4373), .dinb(n4370), .dout(n4374));
  jnot g04135(.din(n4069), .dout(n4375));
  jnot g04136(.din(n4071), .dout(n4376));
  jand g04137(.dina(asqrt[36] ), .dinb(n4065), .dout(n4377));
  jand g04138(.dina(n4377), .dinb(n4376), .dout(n4378));
  jor  g04139(.dina(n4378), .dinb(n4375), .dout(n4379));
  jnot g04140(.din(n4072), .dout(n4380));
  jand g04141(.dina(n4377), .dinb(n4380), .dout(n4381));
  jnot g04142(.din(n4381), .dout(n4382));
  jand g04143(.dina(n4382), .dinb(n4379), .dout(n4383));
  jand g04144(.dina(n4383), .dinb(n4374), .dout(n4384));
  jor  g04145(.dina(n4384), .dinb(n4372), .dout(n4385));
  jand g04146(.dina(n4385), .dinb(asqrt[55] ), .dout(n4386));
  jxor g04147(.dina(n4073), .dinb(n791), .dout(n4387));
  jand g04148(.dina(n4387), .dinb(asqrt[36] ), .dout(n4388));
  jxor g04149(.dina(n4388), .dinb(n4083), .dout(n4389));
  jnot g04150(.din(n4389), .dout(n4390));
  jor  g04151(.dina(n4385), .dinb(asqrt[55] ), .dout(n4391));
  jand g04152(.dina(n4391), .dinb(n4390), .dout(n4392));
  jor  g04153(.dina(n4392), .dinb(n4386), .dout(n4393));
  jand g04154(.dina(n4393), .dinb(asqrt[56] ), .dout(n4394));
  jnot g04155(.din(n4088), .dout(n4395));
  jand g04156(.dina(n4395), .dinb(n4086), .dout(n4396));
  jand g04157(.dina(n4396), .dinb(asqrt[36] ), .dout(n4397));
  jxor g04158(.dina(n4397), .dinb(n4096), .dout(n4398));
  jnot g04159(.din(n4398), .dout(n4399));
  jor  g04160(.dina(n4386), .dinb(asqrt[56] ), .dout(n4400));
  jor  g04161(.dina(n4400), .dinb(n4392), .dout(n4401));
  jand g04162(.dina(n4401), .dinb(n4399), .dout(n4402));
  jor  g04163(.dina(n4402), .dinb(n4394), .dout(n4403));
  jand g04164(.dina(n4403), .dinb(asqrt[57] ), .dout(n4404));
  jor  g04165(.dina(n4403), .dinb(asqrt[57] ), .dout(n4405));
  jnot g04166(.din(n4102), .dout(n4406));
  jnot g04167(.din(n4103), .dout(n4407));
  jand g04168(.dina(asqrt[36] ), .dinb(n4099), .dout(n4408));
  jand g04169(.dina(n4408), .dinb(n4407), .dout(n4409));
  jor  g04170(.dina(n4409), .dinb(n4406), .dout(n4410));
  jnot g04171(.din(n4104), .dout(n4411));
  jand g04172(.dina(n4408), .dinb(n4411), .dout(n4412));
  jnot g04173(.din(n4412), .dout(n4413));
  jand g04174(.dina(n4413), .dinb(n4410), .dout(n4414));
  jand g04175(.dina(n4414), .dinb(n4405), .dout(n4415));
  jor  g04176(.dina(n4415), .dinb(n4404), .dout(n4416));
  jand g04177(.dina(n4416), .dinb(asqrt[58] ), .dout(n4417));
  jor  g04178(.dina(n4404), .dinb(asqrt[58] ), .dout(n4418));
  jor  g04179(.dina(n4418), .dinb(n4415), .dout(n4419));
  jnot g04180(.din(n4110), .dout(n4420));
  jnot g04181(.din(n4112), .dout(n4421));
  jand g04182(.dina(asqrt[36] ), .dinb(n4106), .dout(n4422));
  jand g04183(.dina(n4422), .dinb(n4421), .dout(n4423));
  jor  g04184(.dina(n4423), .dinb(n4420), .dout(n4424));
  jnot g04185(.din(n4113), .dout(n4425));
  jand g04186(.dina(n4422), .dinb(n4425), .dout(n4426));
  jnot g04187(.din(n4426), .dout(n4427));
  jand g04188(.dina(n4427), .dinb(n4424), .dout(n4428));
  jand g04189(.dina(n4428), .dinb(n4419), .dout(n4429));
  jor  g04190(.dina(n4429), .dinb(n4417), .dout(n4430));
  jand g04191(.dina(n4430), .dinb(asqrt[59] ), .dout(n4431));
  jxor g04192(.dina(n4114), .dinb(n425), .dout(n4432));
  jand g04193(.dina(n4432), .dinb(asqrt[36] ), .dout(n4433));
  jxor g04194(.dina(n4433), .dinb(n4124), .dout(n4434));
  jnot g04195(.din(n4434), .dout(n4435));
  jor  g04196(.dina(n4430), .dinb(asqrt[59] ), .dout(n4436));
  jand g04197(.dina(n4436), .dinb(n4435), .dout(n4437));
  jor  g04198(.dina(n4437), .dinb(n4431), .dout(n4438));
  jand g04199(.dina(n4438), .dinb(asqrt[60] ), .dout(n4439));
  jnot g04200(.din(n4129), .dout(n4440));
  jand g04201(.dina(n4440), .dinb(n4127), .dout(n4441));
  jand g04202(.dina(n4441), .dinb(asqrt[36] ), .dout(n4442));
  jxor g04203(.dina(n4442), .dinb(n4137), .dout(n4443));
  jnot g04204(.din(n4443), .dout(n4444));
  jor  g04205(.dina(n4431), .dinb(asqrt[60] ), .dout(n4445));
  jor  g04206(.dina(n4445), .dinb(n4437), .dout(n4446));
  jand g04207(.dina(n4446), .dinb(n4444), .dout(n4447));
  jor  g04208(.dina(n4447), .dinb(n4439), .dout(n4448));
  jand g04209(.dina(n4448), .dinb(asqrt[61] ), .dout(n4449));
  jor  g04210(.dina(n4448), .dinb(asqrt[61] ), .dout(n4450));
  jnot g04211(.din(n4143), .dout(n4451));
  jnot g04212(.din(n4144), .dout(n4452));
  jand g04213(.dina(asqrt[36] ), .dinb(n4140), .dout(n4453));
  jand g04214(.dina(n4453), .dinb(n4452), .dout(n4454));
  jor  g04215(.dina(n4454), .dinb(n4451), .dout(n4455));
  jnot g04216(.din(n4145), .dout(n4456));
  jand g04217(.dina(n4453), .dinb(n4456), .dout(n4457));
  jnot g04218(.din(n4457), .dout(n4458));
  jand g04219(.dina(n4458), .dinb(n4455), .dout(n4459));
  jand g04220(.dina(n4459), .dinb(n4450), .dout(n4460));
  jor  g04221(.dina(n4460), .dinb(n4449), .dout(n4461));
  jand g04222(.dina(n4461), .dinb(asqrt[62] ), .dout(n4462));
  jor  g04223(.dina(n4449), .dinb(asqrt[62] ), .dout(n4463));
  jor  g04224(.dina(n4463), .dinb(n4460), .dout(n4464));
  jnot g04225(.din(n4151), .dout(n4465));
  jnot g04226(.din(n4153), .dout(n4466));
  jand g04227(.dina(asqrt[36] ), .dinb(n4147), .dout(n4467));
  jand g04228(.dina(n4467), .dinb(n4466), .dout(n4468));
  jor  g04229(.dina(n4468), .dinb(n4465), .dout(n4469));
  jnot g04230(.din(n4154), .dout(n4470));
  jand g04231(.dina(n4467), .dinb(n4470), .dout(n4471));
  jnot g04232(.din(n4471), .dout(n4472));
  jand g04233(.dina(n4472), .dinb(n4469), .dout(n4473));
  jand g04234(.dina(n4473), .dinb(n4464), .dout(n4474));
  jor  g04235(.dina(n4474), .dinb(n4462), .dout(n4475));
  jxor g04236(.dina(n4155), .dinb(n199), .dout(n4476));
  jand g04237(.dina(n4476), .dinb(asqrt[36] ), .dout(n4477));
  jxor g04238(.dina(n4477), .dinb(n4165), .dout(n4478));
  jnot g04239(.din(n4167), .dout(n4479));
  jand g04240(.dina(asqrt[36] ), .dinb(n4174), .dout(n4480));
  jand g04241(.dina(n4480), .dinb(n4479), .dout(n4481));
  jor  g04242(.dina(n4481), .dinb(n4182), .dout(n4482));
  jor  g04243(.dina(n4482), .dinb(n4478), .dout(n4483));
  jnot g04244(.din(n4483), .dout(n4484));
  jand g04245(.dina(n4484), .dinb(n4475), .dout(n4485));
  jor  g04246(.dina(n4485), .dinb(asqrt[63] ), .dout(n4486));
  jnot g04247(.din(n4478), .dout(n4487));
  jor  g04248(.dina(n4487), .dinb(n4475), .dout(n4488));
  jor  g04249(.dina(n4480), .dinb(n4479), .dout(n4489));
  jand g04250(.dina(n4174), .dinb(n4479), .dout(n4490));
  jor  g04251(.dina(n4490), .dinb(n194), .dout(n4491));
  jnot g04252(.din(n4491), .dout(n4492));
  jand g04253(.dina(n4492), .dinb(n4489), .dout(n4493));
  jnot g04254(.din(asqrt[36] ), .dout(n4494));
  jnot g04255(.din(n4493), .dout(n4497));
  jand g04256(.dina(n4497), .dinb(n4488), .dout(n4498));
  jand g04257(.dina(n4498), .dinb(n4486), .dout(n4499));
  jnot g04258(.din(n4499), .dout(asqrt[35] ));
  jor  g04259(.dina(n4499), .dinb(n4193), .dout(n4501));
  jnot g04260(.din(a[68] ), .dout(n4502));
  jnot g04261(.din(a[69] ), .dout(n4503));
  jand g04262(.dina(n4193), .dinb(n4503), .dout(n4504));
  jand g04263(.dina(n4504), .dinb(n4502), .dout(n4505));
  jnot g04264(.din(n4505), .dout(n4506));
  jand g04265(.dina(n4506), .dinb(n4501), .dout(n4507));
  jor  g04266(.dina(n4507), .dinb(n4494), .dout(n4508));
  jor  g04267(.dina(n4499), .dinb(a[70] ), .dout(n4509));
  jxor g04268(.dina(n4509), .dinb(n4194), .dout(n4510));
  jand g04269(.dina(n4507), .dinb(n4494), .dout(n4511));
  jor  g04270(.dina(n4511), .dinb(n4510), .dout(n4512));
  jand g04271(.dina(n4512), .dinb(n4508), .dout(n4513));
  jor  g04272(.dina(n4513), .dinb(n3912), .dout(n4514));
  jand g04273(.dina(n4508), .dinb(n3912), .dout(n4515));
  jand g04274(.dina(n4515), .dinb(n4512), .dout(n4516));
  jor  g04275(.dina(n4509), .dinb(a[71] ), .dout(n4517));
  jnot g04276(.din(n4486), .dout(n4518));
  jnot g04277(.din(n4488), .dout(n4519));
  jor  g04278(.dina(n4493), .dinb(n4494), .dout(n4520));
  jor  g04279(.dina(n4520), .dinb(n4519), .dout(n4521));
  jor  g04280(.dina(n4521), .dinb(n4518), .dout(n4522));
  jand g04281(.dina(n4522), .dinb(n4517), .dout(n4523));
  jxor g04282(.dina(n4523), .dinb(n3915), .dout(n4524));
  jor  g04283(.dina(n4524), .dinb(n4516), .dout(n4525));
  jand g04284(.dina(n4525), .dinb(n4514), .dout(n4526));
  jor  g04285(.dina(n4526), .dinb(n3907), .dout(n4527));
  jand g04286(.dina(n4526), .dinb(n3907), .dout(n4528));
  jxor g04287(.dina(n4197), .dinb(n3912), .dout(n4529));
  jor  g04288(.dina(n4529), .dinb(n4499), .dout(n4530));
  jxor g04289(.dina(n4530), .dinb(n4200), .dout(n4531));
  jor  g04290(.dina(n4531), .dinb(n4528), .dout(n4532));
  jand g04291(.dina(n4532), .dinb(n4527), .dout(n4533));
  jor  g04292(.dina(n4533), .dinb(n3376), .dout(n4534));
  jnot g04293(.din(n4206), .dout(n4535));
  jor  g04294(.dina(n4535), .dinb(n4204), .dout(n4536));
  jor  g04295(.dina(n4536), .dinb(n4499), .dout(n4537));
  jxor g04296(.dina(n4537), .dinb(n4215), .dout(n4538));
  jand g04297(.dina(n4527), .dinb(n3376), .dout(n4539));
  jand g04298(.dina(n4539), .dinb(n4532), .dout(n4540));
  jor  g04299(.dina(n4540), .dinb(n4538), .dout(n4541));
  jand g04300(.dina(n4541), .dinb(n4534), .dout(n4542));
  jor  g04301(.dina(n4542), .dinb(n3371), .dout(n4543));
  jand g04302(.dina(n4542), .dinb(n3371), .dout(n4544));
  jxor g04303(.dina(n4217), .dinb(n3376), .dout(n4545));
  jor  g04304(.dina(n4545), .dinb(n4499), .dout(n4546));
  jxor g04305(.dina(n4546), .dinb(n4222), .dout(n4547));
  jnot g04306(.din(n4547), .dout(n4548));
  jor  g04307(.dina(n4548), .dinb(n4544), .dout(n4549));
  jand g04308(.dina(n4549), .dinb(n4543), .dout(n4550));
  jor  g04309(.dina(n4550), .dinb(n2875), .dout(n4551));
  jand g04310(.dina(n4543), .dinb(n2875), .dout(n4552));
  jand g04311(.dina(n4552), .dinb(n4549), .dout(n4553));
  jnot g04312(.din(n4226), .dout(n4554));
  jand g04313(.dina(asqrt[35] ), .dinb(n4554), .dout(n4555));
  jand g04314(.dina(n4555), .dinb(n4233), .dout(n4556));
  jor  g04315(.dina(n4556), .dinb(n4231), .dout(n4557));
  jand g04316(.dina(n4555), .dinb(n4234), .dout(n4558));
  jnot g04317(.din(n4558), .dout(n4559));
  jand g04318(.dina(n4559), .dinb(n4557), .dout(n4560));
  jnot g04319(.din(n4560), .dout(n4561));
  jor  g04320(.dina(n4561), .dinb(n4553), .dout(n4562));
  jand g04321(.dina(n4562), .dinb(n4551), .dout(n4563));
  jor  g04322(.dina(n4563), .dinb(n2870), .dout(n4564));
  jand g04323(.dina(n4563), .dinb(n2870), .dout(n4565));
  jnot g04324(.din(n4241), .dout(n4566));
  jxor g04325(.dina(n4235), .dinb(n2875), .dout(n4567));
  jor  g04326(.dina(n4567), .dinb(n4499), .dout(n4568));
  jxor g04327(.dina(n4568), .dinb(n4566), .dout(n4569));
  jnot g04328(.din(n4569), .dout(n4570));
  jor  g04329(.dina(n4570), .dinb(n4565), .dout(n4571));
  jand g04330(.dina(n4571), .dinb(n4564), .dout(n4572));
  jor  g04331(.dina(n4572), .dinb(n2425), .dout(n4573));
  jnot g04332(.din(n4246), .dout(n4574));
  jor  g04333(.dina(n4574), .dinb(n4244), .dout(n4575));
  jor  g04334(.dina(n4575), .dinb(n4499), .dout(n4576));
  jxor g04335(.dina(n4576), .dinb(n4255), .dout(n4577));
  jand g04336(.dina(n4564), .dinb(n2425), .dout(n4578));
  jand g04337(.dina(n4578), .dinb(n4571), .dout(n4579));
  jor  g04338(.dina(n4579), .dinb(n4577), .dout(n4580));
  jand g04339(.dina(n4580), .dinb(n4573), .dout(n4581));
  jor  g04340(.dina(n4581), .dinb(n2420), .dout(n4582));
  jand g04341(.dina(n4581), .dinb(n2420), .dout(n4583));
  jnot g04342(.din(n4262), .dout(n4584));
  jxor g04343(.dina(n4257), .dinb(n2425), .dout(n4585));
  jor  g04344(.dina(n4585), .dinb(n4499), .dout(n4586));
  jxor g04345(.dina(n4586), .dinb(n4584), .dout(n4587));
  jnot g04346(.din(n4587), .dout(n4588));
  jor  g04347(.dina(n4588), .dinb(n4583), .dout(n4589));
  jand g04348(.dina(n4589), .dinb(n4582), .dout(n4590));
  jor  g04349(.dina(n4590), .dinb(n2010), .dout(n4591));
  jand g04350(.dina(n4582), .dinb(n2010), .dout(n4592));
  jand g04351(.dina(n4592), .dinb(n4589), .dout(n4593));
  jnot g04352(.din(n4265), .dout(n4594));
  jand g04353(.dina(asqrt[35] ), .dinb(n4594), .dout(n4595));
  jand g04354(.dina(n4595), .dinb(n4272), .dout(n4596));
  jor  g04355(.dina(n4596), .dinb(n4270), .dout(n4597));
  jand g04356(.dina(n4595), .dinb(n4273), .dout(n4598));
  jnot g04357(.din(n4598), .dout(n4599));
  jand g04358(.dina(n4599), .dinb(n4597), .dout(n4600));
  jnot g04359(.din(n4600), .dout(n4601));
  jor  g04360(.dina(n4601), .dinb(n4593), .dout(n4602));
  jand g04361(.dina(n4602), .dinb(n4591), .dout(n4603));
  jor  g04362(.dina(n4603), .dinb(n2005), .dout(n4604));
  jxor g04363(.dina(n4274), .dinb(n2010), .dout(n4605));
  jor  g04364(.dina(n4605), .dinb(n4499), .dout(n4606));
  jxor g04365(.dina(n4606), .dinb(n4279), .dout(n4607));
  jand g04366(.dina(n4603), .dinb(n2005), .dout(n4608));
  jor  g04367(.dina(n4608), .dinb(n4607), .dout(n4609));
  jand g04368(.dina(n4609), .dinb(n4604), .dout(n4610));
  jor  g04369(.dina(n4610), .dinb(n1646), .dout(n4611));
  jnot g04370(.din(n4284), .dout(n4612));
  jor  g04371(.dina(n4612), .dinb(n4282), .dout(n4613));
  jor  g04372(.dina(n4613), .dinb(n4499), .dout(n4614));
  jxor g04373(.dina(n4614), .dinb(n4293), .dout(n4615));
  jand g04374(.dina(n4604), .dinb(n1646), .dout(n4616));
  jand g04375(.dina(n4616), .dinb(n4609), .dout(n4617));
  jor  g04376(.dina(n4617), .dinb(n4615), .dout(n4618));
  jand g04377(.dina(n4618), .dinb(n4611), .dout(n4619));
  jor  g04378(.dina(n4619), .dinb(n1641), .dout(n4620));
  jand g04379(.dina(n4619), .dinb(n1641), .dout(n4621));
  jnot g04380(.din(n4296), .dout(n4622));
  jand g04381(.dina(asqrt[35] ), .dinb(n4622), .dout(n4623));
  jand g04382(.dina(n4623), .dinb(n4301), .dout(n4624));
  jor  g04383(.dina(n4624), .dinb(n4300), .dout(n4625));
  jand g04384(.dina(n4623), .dinb(n4302), .dout(n4626));
  jnot g04385(.din(n4626), .dout(n4627));
  jand g04386(.dina(n4627), .dinb(n4625), .dout(n4628));
  jnot g04387(.din(n4628), .dout(n4629));
  jor  g04388(.dina(n4629), .dinb(n4621), .dout(n4630));
  jand g04389(.dina(n4630), .dinb(n4620), .dout(n4631));
  jor  g04390(.dina(n4631), .dinb(n1317), .dout(n4632));
  jand g04391(.dina(n4620), .dinb(n1317), .dout(n4633));
  jand g04392(.dina(n4633), .dinb(n4630), .dout(n4634));
  jnot g04393(.din(n4304), .dout(n4635));
  jand g04394(.dina(asqrt[35] ), .dinb(n4635), .dout(n4636));
  jand g04395(.dina(n4636), .dinb(n4311), .dout(n4637));
  jor  g04396(.dina(n4637), .dinb(n4309), .dout(n4638));
  jand g04397(.dina(n4636), .dinb(n4312), .dout(n4639));
  jnot g04398(.din(n4639), .dout(n4640));
  jand g04399(.dina(n4640), .dinb(n4638), .dout(n4641));
  jnot g04400(.din(n4641), .dout(n4642));
  jor  g04401(.dina(n4642), .dinb(n4634), .dout(n4643));
  jand g04402(.dina(n4643), .dinb(n4632), .dout(n4644));
  jor  g04403(.dina(n4644), .dinb(n1312), .dout(n4645));
  jxor g04404(.dina(n4313), .dinb(n1317), .dout(n4646));
  jor  g04405(.dina(n4646), .dinb(n4499), .dout(n4647));
  jxor g04406(.dina(n4647), .dinb(n4324), .dout(n4648));
  jand g04407(.dina(n4644), .dinb(n1312), .dout(n4649));
  jor  g04408(.dina(n4649), .dinb(n4648), .dout(n4650));
  jand g04409(.dina(n4650), .dinb(n4645), .dout(n4651));
  jor  g04410(.dina(n4651), .dinb(n1039), .dout(n4652));
  jnot g04411(.din(n4329), .dout(n4653));
  jor  g04412(.dina(n4653), .dinb(n4327), .dout(n4654));
  jor  g04413(.dina(n4654), .dinb(n4499), .dout(n4655));
  jxor g04414(.dina(n4655), .dinb(n4338), .dout(n4656));
  jand g04415(.dina(n4645), .dinb(n1039), .dout(n4657));
  jand g04416(.dina(n4657), .dinb(n4650), .dout(n4658));
  jor  g04417(.dina(n4658), .dinb(n4656), .dout(n4659));
  jand g04418(.dina(n4659), .dinb(n4652), .dout(n4660));
  jor  g04419(.dina(n4660), .dinb(n1034), .dout(n4661));
  jand g04420(.dina(n4660), .dinb(n1034), .dout(n4662));
  jnot g04421(.din(n4341), .dout(n4663));
  jand g04422(.dina(asqrt[35] ), .dinb(n4663), .dout(n4664));
  jand g04423(.dina(n4664), .dinb(n4346), .dout(n4665));
  jor  g04424(.dina(n4665), .dinb(n4345), .dout(n4666));
  jand g04425(.dina(n4664), .dinb(n4347), .dout(n4667));
  jnot g04426(.din(n4667), .dout(n4668));
  jand g04427(.dina(n4668), .dinb(n4666), .dout(n4669));
  jnot g04428(.din(n4669), .dout(n4670));
  jor  g04429(.dina(n4670), .dinb(n4662), .dout(n4671));
  jand g04430(.dina(n4671), .dinb(n4661), .dout(n4672));
  jor  g04431(.dina(n4672), .dinb(n796), .dout(n4673));
  jand g04432(.dina(n4661), .dinb(n796), .dout(n4674));
  jand g04433(.dina(n4674), .dinb(n4671), .dout(n4675));
  jnot g04434(.din(n4349), .dout(n4676));
  jand g04435(.dina(asqrt[35] ), .dinb(n4676), .dout(n4677));
  jand g04436(.dina(n4677), .dinb(n4356), .dout(n4678));
  jor  g04437(.dina(n4678), .dinb(n4354), .dout(n4679));
  jand g04438(.dina(n4677), .dinb(n4357), .dout(n4680));
  jnot g04439(.din(n4680), .dout(n4681));
  jand g04440(.dina(n4681), .dinb(n4679), .dout(n4682));
  jnot g04441(.din(n4682), .dout(n4683));
  jor  g04442(.dina(n4683), .dinb(n4675), .dout(n4684));
  jand g04443(.dina(n4684), .dinb(n4673), .dout(n4685));
  jor  g04444(.dina(n4685), .dinb(n791), .dout(n4686));
  jxor g04445(.dina(n4358), .dinb(n796), .dout(n4687));
  jor  g04446(.dina(n4687), .dinb(n4499), .dout(n4688));
  jxor g04447(.dina(n4688), .dinb(n4369), .dout(n4689));
  jand g04448(.dina(n4685), .dinb(n791), .dout(n4690));
  jor  g04449(.dina(n4690), .dinb(n4689), .dout(n4691));
  jand g04450(.dina(n4691), .dinb(n4686), .dout(n4692));
  jor  g04451(.dina(n4692), .dinb(n595), .dout(n4693));
  jnot g04452(.din(n4374), .dout(n4694));
  jor  g04453(.dina(n4694), .dinb(n4372), .dout(n4695));
  jor  g04454(.dina(n4695), .dinb(n4499), .dout(n4696));
  jxor g04455(.dina(n4696), .dinb(n4383), .dout(n4697));
  jand g04456(.dina(n4686), .dinb(n595), .dout(n4698));
  jand g04457(.dina(n4698), .dinb(n4691), .dout(n4699));
  jor  g04458(.dina(n4699), .dinb(n4697), .dout(n4700));
  jand g04459(.dina(n4700), .dinb(n4693), .dout(n4701));
  jor  g04460(.dina(n4701), .dinb(n590), .dout(n4702));
  jand g04461(.dina(n4701), .dinb(n590), .dout(n4703));
  jnot g04462(.din(n4386), .dout(n4704));
  jand g04463(.dina(asqrt[35] ), .dinb(n4704), .dout(n4705));
  jand g04464(.dina(n4705), .dinb(n4391), .dout(n4706));
  jor  g04465(.dina(n4706), .dinb(n4390), .dout(n4707));
  jand g04466(.dina(n4705), .dinb(n4392), .dout(n4708));
  jnot g04467(.din(n4708), .dout(n4709));
  jand g04468(.dina(n4709), .dinb(n4707), .dout(n4710));
  jnot g04469(.din(n4710), .dout(n4711));
  jor  g04470(.dina(n4711), .dinb(n4703), .dout(n4712));
  jand g04471(.dina(n4712), .dinb(n4702), .dout(n4713));
  jor  g04472(.dina(n4713), .dinb(n430), .dout(n4714));
  jand g04473(.dina(n4702), .dinb(n430), .dout(n4715));
  jand g04474(.dina(n4715), .dinb(n4712), .dout(n4716));
  jnot g04475(.din(n4394), .dout(n4717));
  jand g04476(.dina(asqrt[35] ), .dinb(n4717), .dout(n4718));
  jand g04477(.dina(n4718), .dinb(n4401), .dout(n4719));
  jor  g04478(.dina(n4719), .dinb(n4399), .dout(n4720));
  jand g04479(.dina(n4718), .dinb(n4402), .dout(n4721));
  jnot g04480(.din(n4721), .dout(n4722));
  jand g04481(.dina(n4722), .dinb(n4720), .dout(n4723));
  jnot g04482(.din(n4723), .dout(n4724));
  jor  g04483(.dina(n4724), .dinb(n4716), .dout(n4725));
  jand g04484(.dina(n4725), .dinb(n4714), .dout(n4726));
  jor  g04485(.dina(n4726), .dinb(n425), .dout(n4727));
  jxor g04486(.dina(n4403), .dinb(n430), .dout(n4728));
  jor  g04487(.dina(n4728), .dinb(n4499), .dout(n4729));
  jxor g04488(.dina(n4729), .dinb(n4414), .dout(n4730));
  jand g04489(.dina(n4726), .dinb(n425), .dout(n4731));
  jor  g04490(.dina(n4731), .dinb(n4730), .dout(n4732));
  jand g04491(.dina(n4732), .dinb(n4727), .dout(n4733));
  jor  g04492(.dina(n4733), .dinb(n305), .dout(n4734));
  jnot g04493(.din(n4419), .dout(n4735));
  jor  g04494(.dina(n4735), .dinb(n4417), .dout(n4736));
  jor  g04495(.dina(n4736), .dinb(n4499), .dout(n4737));
  jxor g04496(.dina(n4737), .dinb(n4428), .dout(n4738));
  jand g04497(.dina(n4727), .dinb(n305), .dout(n4739));
  jand g04498(.dina(n4739), .dinb(n4732), .dout(n4740));
  jor  g04499(.dina(n4740), .dinb(n4738), .dout(n4741));
  jand g04500(.dina(n4741), .dinb(n4734), .dout(n4742));
  jor  g04501(.dina(n4742), .dinb(n290), .dout(n4743));
  jand g04502(.dina(n4742), .dinb(n290), .dout(n4744));
  jnot g04503(.din(n4431), .dout(n4745));
  jand g04504(.dina(asqrt[35] ), .dinb(n4745), .dout(n4746));
  jand g04505(.dina(n4746), .dinb(n4436), .dout(n4747));
  jor  g04506(.dina(n4747), .dinb(n4435), .dout(n4748));
  jand g04507(.dina(n4746), .dinb(n4437), .dout(n4749));
  jnot g04508(.din(n4749), .dout(n4750));
  jand g04509(.dina(n4750), .dinb(n4748), .dout(n4751));
  jnot g04510(.din(n4751), .dout(n4752));
  jor  g04511(.dina(n4752), .dinb(n4744), .dout(n4753));
  jand g04512(.dina(n4753), .dinb(n4743), .dout(n4754));
  jor  g04513(.dina(n4754), .dinb(n223), .dout(n4755));
  jand g04514(.dina(n4743), .dinb(n223), .dout(n4756));
  jand g04515(.dina(n4756), .dinb(n4753), .dout(n4757));
  jnot g04516(.din(n4439), .dout(n4758));
  jand g04517(.dina(asqrt[35] ), .dinb(n4758), .dout(n4759));
  jand g04518(.dina(n4759), .dinb(n4446), .dout(n4760));
  jor  g04519(.dina(n4760), .dinb(n4444), .dout(n4761));
  jand g04520(.dina(n4759), .dinb(n4447), .dout(n4762));
  jnot g04521(.din(n4762), .dout(n4763));
  jand g04522(.dina(n4763), .dinb(n4761), .dout(n4764));
  jnot g04523(.din(n4764), .dout(n4765));
  jor  g04524(.dina(n4765), .dinb(n4757), .dout(n4766));
  jand g04525(.dina(n4766), .dinb(n4755), .dout(n4767));
  jor  g04526(.dina(n4767), .dinb(n199), .dout(n4768));
  jand g04527(.dina(n4767), .dinb(n199), .dout(n4769));
  jxor g04528(.dina(n4448), .dinb(n223), .dout(n4770));
  jor  g04529(.dina(n4770), .dinb(n4499), .dout(n4771));
  jxor g04530(.dina(n4771), .dinb(n4459), .dout(n4772));
  jor  g04531(.dina(n4772), .dinb(n4769), .dout(n4773));
  jand g04532(.dina(n4773), .dinb(n4768), .dout(n4774));
  jnot g04533(.din(n4464), .dout(n4775));
  jor  g04534(.dina(n4775), .dinb(n4462), .dout(n4776));
  jor  g04535(.dina(n4776), .dinb(n4499), .dout(n4777));
  jxor g04536(.dina(n4777), .dinb(n4473), .dout(n4778));
  jand g04537(.dina(asqrt[35] ), .dinb(n4487), .dout(n4779));
  jand g04538(.dina(n4779), .dinb(n4475), .dout(n4780));
  jor  g04539(.dina(n4780), .dinb(n4519), .dout(n4781));
  jor  g04540(.dina(n4781), .dinb(n4778), .dout(n4782));
  jor  g04541(.dina(n4782), .dinb(n4774), .dout(n4783));
  jand g04542(.dina(n4783), .dinb(n194), .dout(n4784));
  jand g04543(.dina(n4778), .dinb(n4774), .dout(n4785));
  jor  g04544(.dina(n4779), .dinb(n4475), .dout(n4786));
  jand g04545(.dina(n4487), .dinb(n4475), .dout(n4787));
  jor  g04546(.dina(n4787), .dinb(n194), .dout(n4788));
  jnot g04547(.din(n4788), .dout(n4789));
  jand g04548(.dina(n4789), .dinb(n4786), .dout(n4790));
  jor  g04549(.dina(n4790), .dinb(n4785), .dout(n4793));
  jor  g04550(.dina(n4793), .dinb(n4784), .dout(asqrt[34] ));
  jand g04551(.dina(asqrt[34] ), .dinb(a[68] ), .dout(n4795));
  jnot g04552(.din(a[66] ), .dout(n4796));
  jnot g04553(.din(a[67] ), .dout(n4797));
  jand g04554(.dina(n4502), .dinb(n4797), .dout(n4798));
  jand g04555(.dina(n4798), .dinb(n4796), .dout(n4799));
  jor  g04556(.dina(n4799), .dinb(n4795), .dout(n4800));
  jand g04557(.dina(n4800), .dinb(asqrt[35] ), .dout(n4801));
  jand g04558(.dina(asqrt[34] ), .dinb(n4502), .dout(n4802));
  jxor g04559(.dina(n4802), .dinb(n4503), .dout(n4803));
  jor  g04560(.dina(n4800), .dinb(asqrt[35] ), .dout(n4804));
  jand g04561(.dina(n4804), .dinb(n4803), .dout(n4805));
  jor  g04562(.dina(n4805), .dinb(n4801), .dout(n4806));
  jand g04563(.dina(n4806), .dinb(asqrt[36] ), .dout(n4807));
  jor  g04564(.dina(n4801), .dinb(asqrt[36] ), .dout(n4808));
  jor  g04565(.dina(n4808), .dinb(n4805), .dout(n4809));
  jand g04566(.dina(n4802), .dinb(n4503), .dout(n4810));
  jnot g04567(.din(n4784), .dout(n4811));
  jnot g04568(.din(n4785), .dout(n4812));
  jnot g04569(.din(n4790), .dout(n4813));
  jand g04570(.dina(n4813), .dinb(asqrt[35] ), .dout(n4814));
  jand g04571(.dina(n4814), .dinb(n4812), .dout(n4815));
  jand g04572(.dina(n4815), .dinb(n4811), .dout(n4816));
  jor  g04573(.dina(n4816), .dinb(n4810), .dout(n4817));
  jxor g04574(.dina(n4817), .dinb(n4193), .dout(n4818));
  jand g04575(.dina(n4818), .dinb(n4809), .dout(n4819));
  jor  g04576(.dina(n4819), .dinb(n4807), .dout(n4820));
  jand g04577(.dina(n4820), .dinb(asqrt[37] ), .dout(n4821));
  jor  g04578(.dina(n4820), .dinb(asqrt[37] ), .dout(n4822));
  jxor g04579(.dina(n4507), .dinb(n4494), .dout(n4823));
  jand g04580(.dina(n4823), .dinb(asqrt[34] ), .dout(n4824));
  jxor g04581(.dina(n4824), .dinb(n4510), .dout(n4825));
  jnot g04582(.din(n4825), .dout(n4826));
  jand g04583(.dina(n4826), .dinb(n4822), .dout(n4827));
  jor  g04584(.dina(n4827), .dinb(n4821), .dout(n4828));
  jand g04585(.dina(n4828), .dinb(asqrt[38] ), .dout(n4829));
  jnot g04586(.din(n4516), .dout(n4830));
  jand g04587(.dina(n4830), .dinb(n4514), .dout(n4831));
  jand g04588(.dina(n4831), .dinb(asqrt[34] ), .dout(n4832));
  jxor g04589(.dina(n4832), .dinb(n4524), .dout(n4833));
  jnot g04590(.din(n4833), .dout(n4834));
  jor  g04591(.dina(n4821), .dinb(asqrt[38] ), .dout(n4835));
  jor  g04592(.dina(n4835), .dinb(n4827), .dout(n4836));
  jand g04593(.dina(n4836), .dinb(n4834), .dout(n4837));
  jor  g04594(.dina(n4837), .dinb(n4829), .dout(n4838));
  jand g04595(.dina(n4838), .dinb(asqrt[39] ), .dout(n4839));
  jor  g04596(.dina(n4838), .dinb(asqrt[39] ), .dout(n4840));
  jnot g04597(.din(n4531), .dout(n4841));
  jxor g04598(.dina(n4526), .dinb(n3907), .dout(n4842));
  jand g04599(.dina(n4842), .dinb(asqrt[34] ), .dout(n4843));
  jxor g04600(.dina(n4843), .dinb(n4841), .dout(n4844));
  jand g04601(.dina(n4844), .dinb(n4840), .dout(n4845));
  jor  g04602(.dina(n4845), .dinb(n4839), .dout(n4846));
  jand g04603(.dina(n4846), .dinb(asqrt[40] ), .dout(n4847));
  jor  g04604(.dina(n4839), .dinb(asqrt[40] ), .dout(n4848));
  jor  g04605(.dina(n4848), .dinb(n4845), .dout(n4849));
  jnot g04606(.din(n4538), .dout(n4850));
  jnot g04607(.din(n4540), .dout(n4851));
  jand g04608(.dina(asqrt[34] ), .dinb(n4534), .dout(n4852));
  jand g04609(.dina(n4852), .dinb(n4851), .dout(n4853));
  jor  g04610(.dina(n4853), .dinb(n4850), .dout(n4854));
  jnot g04611(.din(n4541), .dout(n4855));
  jand g04612(.dina(n4852), .dinb(n4855), .dout(n4856));
  jnot g04613(.din(n4856), .dout(n4857));
  jand g04614(.dina(n4857), .dinb(n4854), .dout(n4858));
  jand g04615(.dina(n4858), .dinb(n4849), .dout(n4859));
  jor  g04616(.dina(n4859), .dinb(n4847), .dout(n4860));
  jand g04617(.dina(n4860), .dinb(asqrt[41] ), .dout(n4861));
  jor  g04618(.dina(n4860), .dinb(asqrt[41] ), .dout(n4862));
  jxor g04619(.dina(n4542), .dinb(n3371), .dout(n4863));
  jand g04620(.dina(n4863), .dinb(asqrt[34] ), .dout(n4864));
  jxor g04621(.dina(n4864), .dinb(n4547), .dout(n4865));
  jand g04622(.dina(n4865), .dinb(n4862), .dout(n4866));
  jor  g04623(.dina(n4866), .dinb(n4861), .dout(n4867));
  jand g04624(.dina(n4867), .dinb(asqrt[42] ), .dout(n4868));
  jnot g04625(.din(n4553), .dout(n4869));
  jand g04626(.dina(n4869), .dinb(n4551), .dout(n4870));
  jand g04627(.dina(n4870), .dinb(asqrt[34] ), .dout(n4871));
  jxor g04628(.dina(n4871), .dinb(n4561), .dout(n4872));
  jnot g04629(.din(n4872), .dout(n4873));
  jor  g04630(.dina(n4861), .dinb(asqrt[42] ), .dout(n4874));
  jor  g04631(.dina(n4874), .dinb(n4866), .dout(n4875));
  jand g04632(.dina(n4875), .dinb(n4873), .dout(n4876));
  jor  g04633(.dina(n4876), .dinb(n4868), .dout(n4877));
  jand g04634(.dina(n4877), .dinb(asqrt[43] ), .dout(n4878));
  jor  g04635(.dina(n4877), .dinb(asqrt[43] ), .dout(n4879));
  jxor g04636(.dina(n4563), .dinb(n2870), .dout(n4880));
  jand g04637(.dina(n4880), .dinb(asqrt[34] ), .dout(n4881));
  jxor g04638(.dina(n4881), .dinb(n4569), .dout(n4882));
  jand g04639(.dina(n4882), .dinb(n4879), .dout(n4883));
  jor  g04640(.dina(n4883), .dinb(n4878), .dout(n4884));
  jand g04641(.dina(n4884), .dinb(asqrt[44] ), .dout(n4885));
  jor  g04642(.dina(n4878), .dinb(asqrt[44] ), .dout(n4886));
  jor  g04643(.dina(n4886), .dinb(n4883), .dout(n4887));
  jnot g04644(.din(n4577), .dout(n4888));
  jnot g04645(.din(n4579), .dout(n4889));
  jand g04646(.dina(asqrt[34] ), .dinb(n4573), .dout(n4890));
  jand g04647(.dina(n4890), .dinb(n4889), .dout(n4891));
  jor  g04648(.dina(n4891), .dinb(n4888), .dout(n4892));
  jnot g04649(.din(n4580), .dout(n4893));
  jand g04650(.dina(n4890), .dinb(n4893), .dout(n4894));
  jnot g04651(.din(n4894), .dout(n4895));
  jand g04652(.dina(n4895), .dinb(n4892), .dout(n4896));
  jand g04653(.dina(n4896), .dinb(n4887), .dout(n4897));
  jor  g04654(.dina(n4897), .dinb(n4885), .dout(n4898));
  jand g04655(.dina(n4898), .dinb(asqrt[45] ), .dout(n4899));
  jxor g04656(.dina(n4581), .dinb(n2420), .dout(n4900));
  jand g04657(.dina(n4900), .dinb(asqrt[34] ), .dout(n4901));
  jxor g04658(.dina(n4901), .dinb(n4588), .dout(n4902));
  jnot g04659(.din(n4902), .dout(n4903));
  jor  g04660(.dina(n4898), .dinb(asqrt[45] ), .dout(n4904));
  jand g04661(.dina(n4904), .dinb(n4903), .dout(n4905));
  jor  g04662(.dina(n4905), .dinb(n4899), .dout(n4906));
  jand g04663(.dina(n4906), .dinb(asqrt[46] ), .dout(n4907));
  jnot g04664(.din(n4593), .dout(n4908));
  jand g04665(.dina(n4908), .dinb(n4591), .dout(n4909));
  jand g04666(.dina(n4909), .dinb(asqrt[34] ), .dout(n4910));
  jxor g04667(.dina(n4910), .dinb(n4601), .dout(n4911));
  jnot g04668(.din(n4911), .dout(n4912));
  jor  g04669(.dina(n4899), .dinb(asqrt[46] ), .dout(n4913));
  jor  g04670(.dina(n4913), .dinb(n4905), .dout(n4914));
  jand g04671(.dina(n4914), .dinb(n4912), .dout(n4915));
  jor  g04672(.dina(n4915), .dinb(n4907), .dout(n4916));
  jand g04673(.dina(n4916), .dinb(asqrt[47] ), .dout(n4917));
  jor  g04674(.dina(n4916), .dinb(asqrt[47] ), .dout(n4918));
  jnot g04675(.din(n4607), .dout(n4919));
  jnot g04676(.din(n4608), .dout(n4920));
  jand g04677(.dina(asqrt[34] ), .dinb(n4604), .dout(n4921));
  jand g04678(.dina(n4921), .dinb(n4920), .dout(n4922));
  jor  g04679(.dina(n4922), .dinb(n4919), .dout(n4923));
  jnot g04680(.din(n4609), .dout(n4924));
  jand g04681(.dina(n4921), .dinb(n4924), .dout(n4925));
  jnot g04682(.din(n4925), .dout(n4926));
  jand g04683(.dina(n4926), .dinb(n4923), .dout(n4927));
  jand g04684(.dina(n4927), .dinb(n4918), .dout(n4928));
  jor  g04685(.dina(n4928), .dinb(n4917), .dout(n4929));
  jand g04686(.dina(n4929), .dinb(asqrt[48] ), .dout(n4930));
  jor  g04687(.dina(n4917), .dinb(asqrt[48] ), .dout(n4931));
  jor  g04688(.dina(n4931), .dinb(n4928), .dout(n4932));
  jnot g04689(.din(n4615), .dout(n4933));
  jnot g04690(.din(n4617), .dout(n4934));
  jand g04691(.dina(asqrt[34] ), .dinb(n4611), .dout(n4935));
  jand g04692(.dina(n4935), .dinb(n4934), .dout(n4936));
  jor  g04693(.dina(n4936), .dinb(n4933), .dout(n4937));
  jnot g04694(.din(n4618), .dout(n4938));
  jand g04695(.dina(n4935), .dinb(n4938), .dout(n4939));
  jnot g04696(.din(n4939), .dout(n4940));
  jand g04697(.dina(n4940), .dinb(n4937), .dout(n4941));
  jand g04698(.dina(n4941), .dinb(n4932), .dout(n4942));
  jor  g04699(.dina(n4942), .dinb(n4930), .dout(n4943));
  jand g04700(.dina(n4943), .dinb(asqrt[49] ), .dout(n4944));
  jxor g04701(.dina(n4619), .dinb(n1641), .dout(n4945));
  jand g04702(.dina(n4945), .dinb(asqrt[34] ), .dout(n4946));
  jxor g04703(.dina(n4946), .dinb(n4629), .dout(n4947));
  jnot g04704(.din(n4947), .dout(n4948));
  jor  g04705(.dina(n4943), .dinb(asqrt[49] ), .dout(n4949));
  jand g04706(.dina(n4949), .dinb(n4948), .dout(n4950));
  jor  g04707(.dina(n4950), .dinb(n4944), .dout(n4951));
  jand g04708(.dina(n4951), .dinb(asqrt[50] ), .dout(n4952));
  jnot g04709(.din(n4634), .dout(n4953));
  jand g04710(.dina(n4953), .dinb(n4632), .dout(n4954));
  jand g04711(.dina(n4954), .dinb(asqrt[34] ), .dout(n4955));
  jxor g04712(.dina(n4955), .dinb(n4642), .dout(n4956));
  jnot g04713(.din(n4956), .dout(n4957));
  jor  g04714(.dina(n4944), .dinb(asqrt[50] ), .dout(n4958));
  jor  g04715(.dina(n4958), .dinb(n4950), .dout(n4959));
  jand g04716(.dina(n4959), .dinb(n4957), .dout(n4960));
  jor  g04717(.dina(n4960), .dinb(n4952), .dout(n4961));
  jand g04718(.dina(n4961), .dinb(asqrt[51] ), .dout(n4962));
  jor  g04719(.dina(n4961), .dinb(asqrt[51] ), .dout(n4963));
  jnot g04720(.din(n4648), .dout(n4964));
  jnot g04721(.din(n4649), .dout(n4965));
  jand g04722(.dina(asqrt[34] ), .dinb(n4645), .dout(n4966));
  jand g04723(.dina(n4966), .dinb(n4965), .dout(n4967));
  jor  g04724(.dina(n4967), .dinb(n4964), .dout(n4968));
  jnot g04725(.din(n4650), .dout(n4969));
  jand g04726(.dina(n4966), .dinb(n4969), .dout(n4970));
  jnot g04727(.din(n4970), .dout(n4971));
  jand g04728(.dina(n4971), .dinb(n4968), .dout(n4972));
  jand g04729(.dina(n4972), .dinb(n4963), .dout(n4973));
  jor  g04730(.dina(n4973), .dinb(n4962), .dout(n4974));
  jand g04731(.dina(n4974), .dinb(asqrt[52] ), .dout(n4975));
  jor  g04732(.dina(n4962), .dinb(asqrt[52] ), .dout(n4976));
  jor  g04733(.dina(n4976), .dinb(n4973), .dout(n4977));
  jnot g04734(.din(n4656), .dout(n4978));
  jnot g04735(.din(n4658), .dout(n4979));
  jand g04736(.dina(asqrt[34] ), .dinb(n4652), .dout(n4980));
  jand g04737(.dina(n4980), .dinb(n4979), .dout(n4981));
  jor  g04738(.dina(n4981), .dinb(n4978), .dout(n4982));
  jnot g04739(.din(n4659), .dout(n4983));
  jand g04740(.dina(n4980), .dinb(n4983), .dout(n4984));
  jnot g04741(.din(n4984), .dout(n4985));
  jand g04742(.dina(n4985), .dinb(n4982), .dout(n4986));
  jand g04743(.dina(n4986), .dinb(n4977), .dout(n4987));
  jor  g04744(.dina(n4987), .dinb(n4975), .dout(n4988));
  jand g04745(.dina(n4988), .dinb(asqrt[53] ), .dout(n4989));
  jxor g04746(.dina(n4660), .dinb(n1034), .dout(n4990));
  jand g04747(.dina(n4990), .dinb(asqrt[34] ), .dout(n4991));
  jxor g04748(.dina(n4991), .dinb(n4670), .dout(n4992));
  jnot g04749(.din(n4992), .dout(n4993));
  jor  g04750(.dina(n4988), .dinb(asqrt[53] ), .dout(n4994));
  jand g04751(.dina(n4994), .dinb(n4993), .dout(n4995));
  jor  g04752(.dina(n4995), .dinb(n4989), .dout(n4996));
  jand g04753(.dina(n4996), .dinb(asqrt[54] ), .dout(n4997));
  jnot g04754(.din(n4675), .dout(n4998));
  jand g04755(.dina(n4998), .dinb(n4673), .dout(n4999));
  jand g04756(.dina(n4999), .dinb(asqrt[34] ), .dout(n5000));
  jxor g04757(.dina(n5000), .dinb(n4683), .dout(n5001));
  jnot g04758(.din(n5001), .dout(n5002));
  jor  g04759(.dina(n4989), .dinb(asqrt[54] ), .dout(n5003));
  jor  g04760(.dina(n5003), .dinb(n4995), .dout(n5004));
  jand g04761(.dina(n5004), .dinb(n5002), .dout(n5005));
  jor  g04762(.dina(n5005), .dinb(n4997), .dout(n5006));
  jand g04763(.dina(n5006), .dinb(asqrt[55] ), .dout(n5007));
  jor  g04764(.dina(n5006), .dinb(asqrt[55] ), .dout(n5008));
  jnot g04765(.din(n4689), .dout(n5009));
  jnot g04766(.din(n4690), .dout(n5010));
  jand g04767(.dina(asqrt[34] ), .dinb(n4686), .dout(n5011));
  jand g04768(.dina(n5011), .dinb(n5010), .dout(n5012));
  jor  g04769(.dina(n5012), .dinb(n5009), .dout(n5013));
  jnot g04770(.din(n4691), .dout(n5014));
  jand g04771(.dina(n5011), .dinb(n5014), .dout(n5015));
  jnot g04772(.din(n5015), .dout(n5016));
  jand g04773(.dina(n5016), .dinb(n5013), .dout(n5017));
  jand g04774(.dina(n5017), .dinb(n5008), .dout(n5018));
  jor  g04775(.dina(n5018), .dinb(n5007), .dout(n5019));
  jand g04776(.dina(n5019), .dinb(asqrt[56] ), .dout(n5020));
  jor  g04777(.dina(n5007), .dinb(asqrt[56] ), .dout(n5021));
  jor  g04778(.dina(n5021), .dinb(n5018), .dout(n5022));
  jnot g04779(.din(n4697), .dout(n5023));
  jnot g04780(.din(n4699), .dout(n5024));
  jand g04781(.dina(asqrt[34] ), .dinb(n4693), .dout(n5025));
  jand g04782(.dina(n5025), .dinb(n5024), .dout(n5026));
  jor  g04783(.dina(n5026), .dinb(n5023), .dout(n5027));
  jnot g04784(.din(n4700), .dout(n5028));
  jand g04785(.dina(n5025), .dinb(n5028), .dout(n5029));
  jnot g04786(.din(n5029), .dout(n5030));
  jand g04787(.dina(n5030), .dinb(n5027), .dout(n5031));
  jand g04788(.dina(n5031), .dinb(n5022), .dout(n5032));
  jor  g04789(.dina(n5032), .dinb(n5020), .dout(n5033));
  jand g04790(.dina(n5033), .dinb(asqrt[57] ), .dout(n5034));
  jxor g04791(.dina(n4701), .dinb(n590), .dout(n5035));
  jand g04792(.dina(n5035), .dinb(asqrt[34] ), .dout(n5036));
  jxor g04793(.dina(n5036), .dinb(n4711), .dout(n5037));
  jnot g04794(.din(n5037), .dout(n5038));
  jor  g04795(.dina(n5033), .dinb(asqrt[57] ), .dout(n5039));
  jand g04796(.dina(n5039), .dinb(n5038), .dout(n5040));
  jor  g04797(.dina(n5040), .dinb(n5034), .dout(n5041));
  jand g04798(.dina(n5041), .dinb(asqrt[58] ), .dout(n5042));
  jnot g04799(.din(n4716), .dout(n5043));
  jand g04800(.dina(n5043), .dinb(n4714), .dout(n5044));
  jand g04801(.dina(n5044), .dinb(asqrt[34] ), .dout(n5045));
  jxor g04802(.dina(n5045), .dinb(n4724), .dout(n5046));
  jnot g04803(.din(n5046), .dout(n5047));
  jor  g04804(.dina(n5034), .dinb(asqrt[58] ), .dout(n5048));
  jor  g04805(.dina(n5048), .dinb(n5040), .dout(n5049));
  jand g04806(.dina(n5049), .dinb(n5047), .dout(n5050));
  jor  g04807(.dina(n5050), .dinb(n5042), .dout(n5051));
  jand g04808(.dina(n5051), .dinb(asqrt[59] ), .dout(n5052));
  jor  g04809(.dina(n5051), .dinb(asqrt[59] ), .dout(n5053));
  jnot g04810(.din(n4730), .dout(n5054));
  jnot g04811(.din(n4731), .dout(n5055));
  jand g04812(.dina(asqrt[34] ), .dinb(n4727), .dout(n5056));
  jand g04813(.dina(n5056), .dinb(n5055), .dout(n5057));
  jor  g04814(.dina(n5057), .dinb(n5054), .dout(n5058));
  jnot g04815(.din(n4732), .dout(n5059));
  jand g04816(.dina(n5056), .dinb(n5059), .dout(n5060));
  jnot g04817(.din(n5060), .dout(n5061));
  jand g04818(.dina(n5061), .dinb(n5058), .dout(n5062));
  jand g04819(.dina(n5062), .dinb(n5053), .dout(n5063));
  jor  g04820(.dina(n5063), .dinb(n5052), .dout(n5064));
  jand g04821(.dina(n5064), .dinb(asqrt[60] ), .dout(n5065));
  jor  g04822(.dina(n5052), .dinb(asqrt[60] ), .dout(n5066));
  jor  g04823(.dina(n5066), .dinb(n5063), .dout(n5067));
  jnot g04824(.din(n4738), .dout(n5068));
  jnot g04825(.din(n4740), .dout(n5069));
  jand g04826(.dina(asqrt[34] ), .dinb(n4734), .dout(n5070));
  jand g04827(.dina(n5070), .dinb(n5069), .dout(n5071));
  jor  g04828(.dina(n5071), .dinb(n5068), .dout(n5072));
  jnot g04829(.din(n4741), .dout(n5073));
  jand g04830(.dina(n5070), .dinb(n5073), .dout(n5074));
  jnot g04831(.din(n5074), .dout(n5075));
  jand g04832(.dina(n5075), .dinb(n5072), .dout(n5076));
  jand g04833(.dina(n5076), .dinb(n5067), .dout(n5077));
  jor  g04834(.dina(n5077), .dinb(n5065), .dout(n5078));
  jand g04835(.dina(n5078), .dinb(asqrt[61] ), .dout(n5079));
  jxor g04836(.dina(n4742), .dinb(n290), .dout(n5080));
  jand g04837(.dina(n5080), .dinb(asqrt[34] ), .dout(n5081));
  jxor g04838(.dina(n5081), .dinb(n4752), .dout(n5082));
  jnot g04839(.din(n5082), .dout(n5083));
  jor  g04840(.dina(n5078), .dinb(asqrt[61] ), .dout(n5084));
  jand g04841(.dina(n5084), .dinb(n5083), .dout(n5085));
  jor  g04842(.dina(n5085), .dinb(n5079), .dout(n5086));
  jand g04843(.dina(n5086), .dinb(asqrt[62] ), .dout(n5087));
  jnot g04844(.din(n4757), .dout(n5088));
  jand g04845(.dina(n5088), .dinb(n4755), .dout(n5089));
  jand g04846(.dina(n5089), .dinb(asqrt[34] ), .dout(n5090));
  jxor g04847(.dina(n5090), .dinb(n4765), .dout(n5091));
  jnot g04848(.din(n5091), .dout(n5092));
  jor  g04849(.dina(n5079), .dinb(asqrt[62] ), .dout(n5093));
  jor  g04850(.dina(n5093), .dinb(n5085), .dout(n5094));
  jand g04851(.dina(n5094), .dinb(n5092), .dout(n5095));
  jor  g04852(.dina(n5095), .dinb(n5087), .dout(n5096));
  jxor g04853(.dina(n4767), .dinb(n199), .dout(n5097));
  jand g04854(.dina(n5097), .dinb(asqrt[34] ), .dout(n5098));
  jxor g04855(.dina(n5098), .dinb(n4772), .dout(n5099));
  jnot g04856(.din(n4774), .dout(n5100));
  jnot g04857(.din(n4778), .dout(n5101));
  jand g04858(.dina(asqrt[34] ), .dinb(n5101), .dout(n5102));
  jand g04859(.dina(n5102), .dinb(n5100), .dout(n5103));
  jor  g04860(.dina(n5103), .dinb(n4785), .dout(n5104));
  jor  g04861(.dina(n5104), .dinb(n5099), .dout(n5105));
  jnot g04862(.din(n5105), .dout(n5106));
  jand g04863(.dina(n5106), .dinb(n5096), .dout(n5107));
  jor  g04864(.dina(n5107), .dinb(asqrt[63] ), .dout(n5108));
  jnot g04865(.din(n5099), .dout(n5109));
  jor  g04866(.dina(n5109), .dinb(n5096), .dout(n5110));
  jor  g04867(.dina(n5102), .dinb(n5100), .dout(n5111));
  jand g04868(.dina(n5101), .dinb(n5100), .dout(n5112));
  jor  g04869(.dina(n5112), .dinb(n194), .dout(n5113));
  jnot g04870(.din(n5113), .dout(n5114));
  jand g04871(.dina(n5114), .dinb(n5111), .dout(n5115));
  jnot g04872(.din(asqrt[34] ), .dout(n5116));
  jnot g04873(.din(n5115), .dout(n5119));
  jand g04874(.dina(n5119), .dinb(n5110), .dout(n5120));
  jand g04875(.dina(n5120), .dinb(n5108), .dout(n5121));
  jnot g04876(.din(n5121), .dout(asqrt[33] ));
  jor  g04877(.dina(n5121), .dinb(n4796), .dout(n5123));
  jnot g04878(.din(a[64] ), .dout(n5124));
  jnot g04879(.din(a[65] ), .dout(n5125));
  jand g04880(.dina(n4796), .dinb(n5125), .dout(n5126));
  jand g04881(.dina(n5126), .dinb(n5124), .dout(n5127));
  jnot g04882(.din(n5127), .dout(n5128));
  jand g04883(.dina(n5128), .dinb(n5123), .dout(n5129));
  jor  g04884(.dina(n5129), .dinb(n5116), .dout(n5130));
  jor  g04885(.dina(n5121), .dinb(a[66] ), .dout(n5131));
  jxor g04886(.dina(n5131), .dinb(n4797), .dout(n5132));
  jand g04887(.dina(n5129), .dinb(n5116), .dout(n5133));
  jor  g04888(.dina(n5133), .dinb(n5132), .dout(n5134));
  jand g04889(.dina(n5134), .dinb(n5130), .dout(n5135));
  jor  g04890(.dina(n5135), .dinb(n4499), .dout(n5136));
  jand g04891(.dina(n5130), .dinb(n4499), .dout(n5137));
  jand g04892(.dina(n5137), .dinb(n5134), .dout(n5138));
  jor  g04893(.dina(n5131), .dinb(a[67] ), .dout(n5139));
  jnot g04894(.din(n5108), .dout(n5140));
  jnot g04895(.din(n5110), .dout(n5141));
  jor  g04896(.dina(n5115), .dinb(n5116), .dout(n5142));
  jor  g04897(.dina(n5142), .dinb(n5141), .dout(n5143));
  jor  g04898(.dina(n5143), .dinb(n5140), .dout(n5144));
  jand g04899(.dina(n5144), .dinb(n5139), .dout(n5145));
  jxor g04900(.dina(n5145), .dinb(n4502), .dout(n5146));
  jor  g04901(.dina(n5146), .dinb(n5138), .dout(n5147));
  jand g04902(.dina(n5147), .dinb(n5136), .dout(n5148));
  jor  g04903(.dina(n5148), .dinb(n4494), .dout(n5149));
  jand g04904(.dina(n5148), .dinb(n4494), .dout(n5150));
  jxor g04905(.dina(n4800), .dinb(n4499), .dout(n5151));
  jor  g04906(.dina(n5151), .dinb(n5121), .dout(n5152));
  jxor g04907(.dina(n5152), .dinb(n4803), .dout(n5153));
  jor  g04908(.dina(n5153), .dinb(n5150), .dout(n5154));
  jand g04909(.dina(n5154), .dinb(n5149), .dout(n5155));
  jor  g04910(.dina(n5155), .dinb(n3912), .dout(n5156));
  jnot g04911(.din(n4809), .dout(n5157));
  jor  g04912(.dina(n5157), .dinb(n4807), .dout(n5158));
  jor  g04913(.dina(n5158), .dinb(n5121), .dout(n5159));
  jxor g04914(.dina(n5159), .dinb(n4818), .dout(n5160));
  jand g04915(.dina(n5149), .dinb(n3912), .dout(n5161));
  jand g04916(.dina(n5161), .dinb(n5154), .dout(n5162));
  jor  g04917(.dina(n5162), .dinb(n5160), .dout(n5163));
  jand g04918(.dina(n5163), .dinb(n5156), .dout(n5164));
  jor  g04919(.dina(n5164), .dinb(n3907), .dout(n5165));
  jand g04920(.dina(n5164), .dinb(n3907), .dout(n5166));
  jxor g04921(.dina(n4820), .dinb(n3912), .dout(n5167));
  jor  g04922(.dina(n5167), .dinb(n5121), .dout(n5168));
  jxor g04923(.dina(n5168), .dinb(n4825), .dout(n5169));
  jnot g04924(.din(n5169), .dout(n5170));
  jor  g04925(.dina(n5170), .dinb(n5166), .dout(n5171));
  jand g04926(.dina(n5171), .dinb(n5165), .dout(n5172));
  jor  g04927(.dina(n5172), .dinb(n3376), .dout(n5173));
  jand g04928(.dina(n5165), .dinb(n3376), .dout(n5174));
  jand g04929(.dina(n5174), .dinb(n5171), .dout(n5175));
  jnot g04930(.din(n4829), .dout(n5176));
  jand g04931(.dina(asqrt[33] ), .dinb(n5176), .dout(n5177));
  jand g04932(.dina(n5177), .dinb(n4836), .dout(n5178));
  jor  g04933(.dina(n5178), .dinb(n4834), .dout(n5179));
  jand g04934(.dina(n5177), .dinb(n4837), .dout(n5180));
  jnot g04935(.din(n5180), .dout(n5181));
  jand g04936(.dina(n5181), .dinb(n5179), .dout(n5182));
  jnot g04937(.din(n5182), .dout(n5183));
  jor  g04938(.dina(n5183), .dinb(n5175), .dout(n5184));
  jand g04939(.dina(n5184), .dinb(n5173), .dout(n5185));
  jor  g04940(.dina(n5185), .dinb(n3371), .dout(n5186));
  jand g04941(.dina(n5185), .dinb(n3371), .dout(n5187));
  jnot g04942(.din(n4844), .dout(n5188));
  jxor g04943(.dina(n4838), .dinb(n3376), .dout(n5189));
  jor  g04944(.dina(n5189), .dinb(n5121), .dout(n5190));
  jxor g04945(.dina(n5190), .dinb(n5188), .dout(n5191));
  jnot g04946(.din(n5191), .dout(n5192));
  jor  g04947(.dina(n5192), .dinb(n5187), .dout(n5193));
  jand g04948(.dina(n5193), .dinb(n5186), .dout(n5194));
  jor  g04949(.dina(n5194), .dinb(n2875), .dout(n5195));
  jnot g04950(.din(n4849), .dout(n5196));
  jor  g04951(.dina(n5196), .dinb(n4847), .dout(n5197));
  jor  g04952(.dina(n5197), .dinb(n5121), .dout(n5198));
  jxor g04953(.dina(n5198), .dinb(n4858), .dout(n5199));
  jand g04954(.dina(n5186), .dinb(n2875), .dout(n5200));
  jand g04955(.dina(n5200), .dinb(n5193), .dout(n5201));
  jor  g04956(.dina(n5201), .dinb(n5199), .dout(n5202));
  jand g04957(.dina(n5202), .dinb(n5195), .dout(n5203));
  jor  g04958(.dina(n5203), .dinb(n2870), .dout(n5204));
  jand g04959(.dina(n5203), .dinb(n2870), .dout(n5205));
  jnot g04960(.din(n4865), .dout(n5206));
  jxor g04961(.dina(n4860), .dinb(n2875), .dout(n5207));
  jor  g04962(.dina(n5207), .dinb(n5121), .dout(n5208));
  jxor g04963(.dina(n5208), .dinb(n5206), .dout(n5209));
  jnot g04964(.din(n5209), .dout(n5210));
  jor  g04965(.dina(n5210), .dinb(n5205), .dout(n5211));
  jand g04966(.dina(n5211), .dinb(n5204), .dout(n5212));
  jor  g04967(.dina(n5212), .dinb(n2425), .dout(n5213));
  jand g04968(.dina(n5204), .dinb(n2425), .dout(n5214));
  jand g04969(.dina(n5214), .dinb(n5211), .dout(n5215));
  jnot g04970(.din(n4868), .dout(n5216));
  jand g04971(.dina(asqrt[33] ), .dinb(n5216), .dout(n5217));
  jand g04972(.dina(n5217), .dinb(n4875), .dout(n5218));
  jor  g04973(.dina(n5218), .dinb(n4873), .dout(n5219));
  jand g04974(.dina(n5217), .dinb(n4876), .dout(n5220));
  jnot g04975(.din(n5220), .dout(n5221));
  jand g04976(.dina(n5221), .dinb(n5219), .dout(n5222));
  jnot g04977(.din(n5222), .dout(n5223));
  jor  g04978(.dina(n5223), .dinb(n5215), .dout(n5224));
  jand g04979(.dina(n5224), .dinb(n5213), .dout(n5225));
  jor  g04980(.dina(n5225), .dinb(n2420), .dout(n5226));
  jxor g04981(.dina(n4877), .dinb(n2425), .dout(n5227));
  jor  g04982(.dina(n5227), .dinb(n5121), .dout(n5228));
  jxor g04983(.dina(n5228), .dinb(n4882), .dout(n5229));
  jand g04984(.dina(n5225), .dinb(n2420), .dout(n5230));
  jor  g04985(.dina(n5230), .dinb(n5229), .dout(n5231));
  jand g04986(.dina(n5231), .dinb(n5226), .dout(n5232));
  jor  g04987(.dina(n5232), .dinb(n2010), .dout(n5233));
  jnot g04988(.din(n4887), .dout(n5234));
  jor  g04989(.dina(n5234), .dinb(n4885), .dout(n5235));
  jor  g04990(.dina(n5235), .dinb(n5121), .dout(n5236));
  jxor g04991(.dina(n5236), .dinb(n4896), .dout(n5237));
  jand g04992(.dina(n5226), .dinb(n2010), .dout(n5238));
  jand g04993(.dina(n5238), .dinb(n5231), .dout(n5239));
  jor  g04994(.dina(n5239), .dinb(n5237), .dout(n5240));
  jand g04995(.dina(n5240), .dinb(n5233), .dout(n5241));
  jor  g04996(.dina(n5241), .dinb(n2005), .dout(n5242));
  jand g04997(.dina(n5241), .dinb(n2005), .dout(n5243));
  jnot g04998(.din(n4899), .dout(n5244));
  jand g04999(.dina(asqrt[33] ), .dinb(n5244), .dout(n5245));
  jand g05000(.dina(n5245), .dinb(n4904), .dout(n5246));
  jor  g05001(.dina(n5246), .dinb(n4903), .dout(n5247));
  jand g05002(.dina(n5245), .dinb(n4905), .dout(n5248));
  jnot g05003(.din(n5248), .dout(n5249));
  jand g05004(.dina(n5249), .dinb(n5247), .dout(n5250));
  jnot g05005(.din(n5250), .dout(n5251));
  jor  g05006(.dina(n5251), .dinb(n5243), .dout(n5252));
  jand g05007(.dina(n5252), .dinb(n5242), .dout(n5253));
  jor  g05008(.dina(n5253), .dinb(n1646), .dout(n5254));
  jand g05009(.dina(n5242), .dinb(n1646), .dout(n5255));
  jand g05010(.dina(n5255), .dinb(n5252), .dout(n5256));
  jnot g05011(.din(n4907), .dout(n5257));
  jand g05012(.dina(asqrt[33] ), .dinb(n5257), .dout(n5258));
  jand g05013(.dina(n5258), .dinb(n4914), .dout(n5259));
  jor  g05014(.dina(n5259), .dinb(n4912), .dout(n5260));
  jand g05015(.dina(n5258), .dinb(n4915), .dout(n5261));
  jnot g05016(.din(n5261), .dout(n5262));
  jand g05017(.dina(n5262), .dinb(n5260), .dout(n5263));
  jnot g05018(.din(n5263), .dout(n5264));
  jor  g05019(.dina(n5264), .dinb(n5256), .dout(n5265));
  jand g05020(.dina(n5265), .dinb(n5254), .dout(n5266));
  jor  g05021(.dina(n5266), .dinb(n1641), .dout(n5267));
  jxor g05022(.dina(n4916), .dinb(n1646), .dout(n5268));
  jor  g05023(.dina(n5268), .dinb(n5121), .dout(n5269));
  jxor g05024(.dina(n5269), .dinb(n4927), .dout(n5270));
  jand g05025(.dina(n5266), .dinb(n1641), .dout(n5271));
  jor  g05026(.dina(n5271), .dinb(n5270), .dout(n5272));
  jand g05027(.dina(n5272), .dinb(n5267), .dout(n5273));
  jor  g05028(.dina(n5273), .dinb(n1317), .dout(n5274));
  jnot g05029(.din(n4932), .dout(n5275));
  jor  g05030(.dina(n5275), .dinb(n4930), .dout(n5276));
  jor  g05031(.dina(n5276), .dinb(n5121), .dout(n5277));
  jxor g05032(.dina(n5277), .dinb(n4941), .dout(n5278));
  jand g05033(.dina(n5267), .dinb(n1317), .dout(n5279));
  jand g05034(.dina(n5279), .dinb(n5272), .dout(n5280));
  jor  g05035(.dina(n5280), .dinb(n5278), .dout(n5281));
  jand g05036(.dina(n5281), .dinb(n5274), .dout(n5282));
  jor  g05037(.dina(n5282), .dinb(n1312), .dout(n5283));
  jand g05038(.dina(n5282), .dinb(n1312), .dout(n5284));
  jnot g05039(.din(n4944), .dout(n5285));
  jand g05040(.dina(asqrt[33] ), .dinb(n5285), .dout(n5286));
  jand g05041(.dina(n5286), .dinb(n4949), .dout(n5287));
  jor  g05042(.dina(n5287), .dinb(n4948), .dout(n5288));
  jand g05043(.dina(n5286), .dinb(n4950), .dout(n5289));
  jnot g05044(.din(n5289), .dout(n5290));
  jand g05045(.dina(n5290), .dinb(n5288), .dout(n5291));
  jnot g05046(.din(n5291), .dout(n5292));
  jor  g05047(.dina(n5292), .dinb(n5284), .dout(n5293));
  jand g05048(.dina(n5293), .dinb(n5283), .dout(n5294));
  jor  g05049(.dina(n5294), .dinb(n1039), .dout(n5295));
  jand g05050(.dina(n5283), .dinb(n1039), .dout(n5296));
  jand g05051(.dina(n5296), .dinb(n5293), .dout(n5297));
  jnot g05052(.din(n4952), .dout(n5298));
  jand g05053(.dina(asqrt[33] ), .dinb(n5298), .dout(n5299));
  jand g05054(.dina(n5299), .dinb(n4959), .dout(n5300));
  jor  g05055(.dina(n5300), .dinb(n4957), .dout(n5301));
  jand g05056(.dina(n5299), .dinb(n4960), .dout(n5302));
  jnot g05057(.din(n5302), .dout(n5303));
  jand g05058(.dina(n5303), .dinb(n5301), .dout(n5304));
  jnot g05059(.din(n5304), .dout(n5305));
  jor  g05060(.dina(n5305), .dinb(n5297), .dout(n5306));
  jand g05061(.dina(n5306), .dinb(n5295), .dout(n5307));
  jor  g05062(.dina(n5307), .dinb(n1034), .dout(n5308));
  jxor g05063(.dina(n4961), .dinb(n1039), .dout(n5309));
  jor  g05064(.dina(n5309), .dinb(n5121), .dout(n5310));
  jxor g05065(.dina(n5310), .dinb(n4972), .dout(n5311));
  jand g05066(.dina(n5307), .dinb(n1034), .dout(n5312));
  jor  g05067(.dina(n5312), .dinb(n5311), .dout(n5313));
  jand g05068(.dina(n5313), .dinb(n5308), .dout(n5314));
  jor  g05069(.dina(n5314), .dinb(n796), .dout(n5315));
  jnot g05070(.din(n4977), .dout(n5316));
  jor  g05071(.dina(n5316), .dinb(n4975), .dout(n5317));
  jor  g05072(.dina(n5317), .dinb(n5121), .dout(n5318));
  jxor g05073(.dina(n5318), .dinb(n4986), .dout(n5319));
  jand g05074(.dina(n5308), .dinb(n796), .dout(n5320));
  jand g05075(.dina(n5320), .dinb(n5313), .dout(n5321));
  jor  g05076(.dina(n5321), .dinb(n5319), .dout(n5322));
  jand g05077(.dina(n5322), .dinb(n5315), .dout(n5323));
  jor  g05078(.dina(n5323), .dinb(n791), .dout(n5324));
  jand g05079(.dina(n5323), .dinb(n791), .dout(n5325));
  jnot g05080(.din(n4989), .dout(n5326));
  jand g05081(.dina(asqrt[33] ), .dinb(n5326), .dout(n5327));
  jand g05082(.dina(n5327), .dinb(n4994), .dout(n5328));
  jor  g05083(.dina(n5328), .dinb(n4993), .dout(n5329));
  jand g05084(.dina(n5327), .dinb(n4995), .dout(n5330));
  jnot g05085(.din(n5330), .dout(n5331));
  jand g05086(.dina(n5331), .dinb(n5329), .dout(n5332));
  jnot g05087(.din(n5332), .dout(n5333));
  jor  g05088(.dina(n5333), .dinb(n5325), .dout(n5334));
  jand g05089(.dina(n5334), .dinb(n5324), .dout(n5335));
  jor  g05090(.dina(n5335), .dinb(n595), .dout(n5336));
  jand g05091(.dina(n5324), .dinb(n595), .dout(n5337));
  jand g05092(.dina(n5337), .dinb(n5334), .dout(n5338));
  jnot g05093(.din(n4997), .dout(n5339));
  jand g05094(.dina(asqrt[33] ), .dinb(n5339), .dout(n5340));
  jand g05095(.dina(n5340), .dinb(n5004), .dout(n5341));
  jor  g05096(.dina(n5341), .dinb(n5002), .dout(n5342));
  jand g05097(.dina(n5340), .dinb(n5005), .dout(n5343));
  jnot g05098(.din(n5343), .dout(n5344));
  jand g05099(.dina(n5344), .dinb(n5342), .dout(n5345));
  jnot g05100(.din(n5345), .dout(n5346));
  jor  g05101(.dina(n5346), .dinb(n5338), .dout(n5347));
  jand g05102(.dina(n5347), .dinb(n5336), .dout(n5348));
  jor  g05103(.dina(n5348), .dinb(n590), .dout(n5349));
  jxor g05104(.dina(n5006), .dinb(n595), .dout(n5350));
  jor  g05105(.dina(n5350), .dinb(n5121), .dout(n5351));
  jxor g05106(.dina(n5351), .dinb(n5017), .dout(n5352));
  jand g05107(.dina(n5348), .dinb(n590), .dout(n5353));
  jor  g05108(.dina(n5353), .dinb(n5352), .dout(n5354));
  jand g05109(.dina(n5354), .dinb(n5349), .dout(n5355));
  jor  g05110(.dina(n5355), .dinb(n430), .dout(n5356));
  jnot g05111(.din(n5022), .dout(n5357));
  jor  g05112(.dina(n5357), .dinb(n5020), .dout(n5358));
  jor  g05113(.dina(n5358), .dinb(n5121), .dout(n5359));
  jxor g05114(.dina(n5359), .dinb(n5031), .dout(n5360));
  jand g05115(.dina(n5349), .dinb(n430), .dout(n5361));
  jand g05116(.dina(n5361), .dinb(n5354), .dout(n5362));
  jor  g05117(.dina(n5362), .dinb(n5360), .dout(n5363));
  jand g05118(.dina(n5363), .dinb(n5356), .dout(n5364));
  jor  g05119(.dina(n5364), .dinb(n425), .dout(n5365));
  jand g05120(.dina(n5364), .dinb(n425), .dout(n5366));
  jnot g05121(.din(n5034), .dout(n5367));
  jand g05122(.dina(asqrt[33] ), .dinb(n5367), .dout(n5368));
  jand g05123(.dina(n5368), .dinb(n5039), .dout(n5369));
  jor  g05124(.dina(n5369), .dinb(n5038), .dout(n5370));
  jand g05125(.dina(n5368), .dinb(n5040), .dout(n5371));
  jnot g05126(.din(n5371), .dout(n5372));
  jand g05127(.dina(n5372), .dinb(n5370), .dout(n5373));
  jnot g05128(.din(n5373), .dout(n5374));
  jor  g05129(.dina(n5374), .dinb(n5366), .dout(n5375));
  jand g05130(.dina(n5375), .dinb(n5365), .dout(n5376));
  jor  g05131(.dina(n5376), .dinb(n305), .dout(n5377));
  jand g05132(.dina(n5365), .dinb(n305), .dout(n5378));
  jand g05133(.dina(n5378), .dinb(n5375), .dout(n5379));
  jnot g05134(.din(n5042), .dout(n5380));
  jand g05135(.dina(asqrt[33] ), .dinb(n5380), .dout(n5381));
  jand g05136(.dina(n5381), .dinb(n5049), .dout(n5382));
  jor  g05137(.dina(n5382), .dinb(n5047), .dout(n5383));
  jand g05138(.dina(n5381), .dinb(n5050), .dout(n5384));
  jnot g05139(.din(n5384), .dout(n5385));
  jand g05140(.dina(n5385), .dinb(n5383), .dout(n5386));
  jnot g05141(.din(n5386), .dout(n5387));
  jor  g05142(.dina(n5387), .dinb(n5379), .dout(n5388));
  jand g05143(.dina(n5388), .dinb(n5377), .dout(n5389));
  jor  g05144(.dina(n5389), .dinb(n290), .dout(n5390));
  jxor g05145(.dina(n5051), .dinb(n305), .dout(n5391));
  jor  g05146(.dina(n5391), .dinb(n5121), .dout(n5392));
  jxor g05147(.dina(n5392), .dinb(n5062), .dout(n5393));
  jand g05148(.dina(n5389), .dinb(n290), .dout(n5394));
  jor  g05149(.dina(n5394), .dinb(n5393), .dout(n5395));
  jand g05150(.dina(n5395), .dinb(n5390), .dout(n5396));
  jor  g05151(.dina(n5396), .dinb(n223), .dout(n5397));
  jnot g05152(.din(n5067), .dout(n5398));
  jor  g05153(.dina(n5398), .dinb(n5065), .dout(n5399));
  jor  g05154(.dina(n5399), .dinb(n5121), .dout(n5400));
  jxor g05155(.dina(n5400), .dinb(n5076), .dout(n5401));
  jand g05156(.dina(n5390), .dinb(n223), .dout(n5402));
  jand g05157(.dina(n5402), .dinb(n5395), .dout(n5403));
  jor  g05158(.dina(n5403), .dinb(n5401), .dout(n5404));
  jand g05159(.dina(n5404), .dinb(n5397), .dout(n5405));
  jor  g05160(.dina(n5405), .dinb(n199), .dout(n5406));
  jand g05161(.dina(n5405), .dinb(n199), .dout(n5407));
  jnot g05162(.din(n5079), .dout(n5408));
  jand g05163(.dina(asqrt[33] ), .dinb(n5408), .dout(n5409));
  jand g05164(.dina(n5409), .dinb(n5084), .dout(n5410));
  jor  g05165(.dina(n5410), .dinb(n5083), .dout(n5411));
  jand g05166(.dina(n5409), .dinb(n5085), .dout(n5412));
  jnot g05167(.din(n5412), .dout(n5413));
  jand g05168(.dina(n5413), .dinb(n5411), .dout(n5414));
  jnot g05169(.din(n5414), .dout(n5415));
  jor  g05170(.dina(n5415), .dinb(n5407), .dout(n5416));
  jand g05171(.dina(n5416), .dinb(n5406), .dout(n5417));
  jnot g05172(.din(n5087), .dout(n5418));
  jand g05173(.dina(asqrt[33] ), .dinb(n5418), .dout(n5419));
  jand g05174(.dina(n5419), .dinb(n5094), .dout(n5420));
  jor  g05175(.dina(n5420), .dinb(n5092), .dout(n5421));
  jand g05176(.dina(n5419), .dinb(n5095), .dout(n5422));
  jnot g05177(.din(n5422), .dout(n5423));
  jand g05178(.dina(n5423), .dinb(n5421), .dout(n5424));
  jnot g05179(.din(n5424), .dout(n5425));
  jand g05180(.dina(asqrt[33] ), .dinb(n5109), .dout(n5426));
  jand g05181(.dina(n5426), .dinb(n5096), .dout(n5427));
  jor  g05182(.dina(n5427), .dinb(n5141), .dout(n5428));
  jor  g05183(.dina(n5428), .dinb(n5425), .dout(n5429));
  jor  g05184(.dina(n5429), .dinb(n5417), .dout(n5430));
  jand g05185(.dina(n5430), .dinb(n194), .dout(n5431));
  jand g05186(.dina(n5425), .dinb(n5417), .dout(n5432));
  jor  g05187(.dina(n5426), .dinb(n5096), .dout(n5433));
  jand g05188(.dina(n5109), .dinb(n5096), .dout(n5434));
  jor  g05189(.dina(n5434), .dinb(n194), .dout(n5435));
  jnot g05190(.din(n5435), .dout(n5436));
  jand g05191(.dina(n5436), .dinb(n5433), .dout(n5437));
  jor  g05192(.dina(n5437), .dinb(n5432), .dout(n5440));
  jor  g05193(.dina(n5440), .dinb(n5431), .dout(asqrt[32] ));
  jand g05194(.dina(asqrt[32] ), .dinb(a[64] ), .dout(n5442));
  jnot g05195(.din(a[62] ), .dout(n5443));
  jand g05196(.dina(n5124), .dinb(n200), .dout(n5444));
  jand g05197(.dina(n5444), .dinb(n5443), .dout(n5445));
  jor  g05198(.dina(n5445), .dinb(n5442), .dout(n5446));
  jand g05199(.dina(n5446), .dinb(asqrt[33] ), .dout(n5447));
  jand g05200(.dina(asqrt[32] ), .dinb(n5124), .dout(n5448));
  jxor g05201(.dina(n5448), .dinb(n5125), .dout(n5449));
  jor  g05202(.dina(n5446), .dinb(asqrt[33] ), .dout(n5450));
  jand g05203(.dina(n5450), .dinb(n5449), .dout(n5451));
  jor  g05204(.dina(n5451), .dinb(n5447), .dout(n5452));
  jand g05205(.dina(n5452), .dinb(asqrt[34] ), .dout(n5453));
  jor  g05206(.dina(n5447), .dinb(asqrt[34] ), .dout(n5454));
  jor  g05207(.dina(n5454), .dinb(n5451), .dout(n5455));
  jand g05208(.dina(n5448), .dinb(n5125), .dout(n5456));
  jnot g05209(.din(n5431), .dout(n5457));
  jnot g05210(.din(n5432), .dout(n5458));
  jnot g05211(.din(n5437), .dout(n5459));
  jand g05212(.dina(n5459), .dinb(asqrt[33] ), .dout(n5460));
  jand g05213(.dina(n5460), .dinb(n5458), .dout(n5461));
  jand g05214(.dina(n5461), .dinb(n5457), .dout(n5462));
  jor  g05215(.dina(n5462), .dinb(n5456), .dout(n5463));
  jxor g05216(.dina(n5463), .dinb(n4796), .dout(n5464));
  jand g05217(.dina(n5464), .dinb(n5455), .dout(n5465));
  jor  g05218(.dina(n5465), .dinb(n5453), .dout(n5466));
  jand g05219(.dina(n5466), .dinb(asqrt[35] ), .dout(n5467));
  jor  g05220(.dina(n5466), .dinb(asqrt[35] ), .dout(n5468));
  jxor g05221(.dina(n5129), .dinb(n5116), .dout(n5469));
  jand g05222(.dina(n5469), .dinb(asqrt[32] ), .dout(n5470));
  jxor g05223(.dina(n5470), .dinb(n5132), .dout(n5471));
  jnot g05224(.din(n5471), .dout(n5472));
  jand g05225(.dina(n5472), .dinb(n5468), .dout(n5473));
  jor  g05226(.dina(n5473), .dinb(n5467), .dout(n5474));
  jand g05227(.dina(n5474), .dinb(asqrt[36] ), .dout(n5475));
  jnot g05228(.din(n5138), .dout(n5476));
  jand g05229(.dina(n5476), .dinb(n5136), .dout(n5477));
  jand g05230(.dina(n5477), .dinb(asqrt[32] ), .dout(n5478));
  jxor g05231(.dina(n5478), .dinb(n5146), .dout(n5479));
  jnot g05232(.din(n5479), .dout(n5480));
  jor  g05233(.dina(n5467), .dinb(asqrt[36] ), .dout(n5481));
  jor  g05234(.dina(n5481), .dinb(n5473), .dout(n5482));
  jand g05235(.dina(n5482), .dinb(n5480), .dout(n5483));
  jor  g05236(.dina(n5483), .dinb(n5475), .dout(n5484));
  jand g05237(.dina(n5484), .dinb(asqrt[37] ), .dout(n5485));
  jor  g05238(.dina(n5484), .dinb(asqrt[37] ), .dout(n5486));
  jnot g05239(.din(n5153), .dout(n5487));
  jxor g05240(.dina(n5148), .dinb(n4494), .dout(n5488));
  jand g05241(.dina(n5488), .dinb(asqrt[32] ), .dout(n5489));
  jxor g05242(.dina(n5489), .dinb(n5487), .dout(n5490));
  jand g05243(.dina(n5490), .dinb(n5486), .dout(n5491));
  jor  g05244(.dina(n5491), .dinb(n5485), .dout(n5492));
  jand g05245(.dina(n5492), .dinb(asqrt[38] ), .dout(n5493));
  jor  g05246(.dina(n5485), .dinb(asqrt[38] ), .dout(n5494));
  jor  g05247(.dina(n5494), .dinb(n5491), .dout(n5495));
  jnot g05248(.din(n5160), .dout(n5496));
  jnot g05249(.din(n5162), .dout(n5497));
  jand g05250(.dina(asqrt[32] ), .dinb(n5156), .dout(n5498));
  jand g05251(.dina(n5498), .dinb(n5497), .dout(n5499));
  jor  g05252(.dina(n5499), .dinb(n5496), .dout(n5500));
  jnot g05253(.din(n5163), .dout(n5501));
  jand g05254(.dina(n5498), .dinb(n5501), .dout(n5502));
  jnot g05255(.din(n5502), .dout(n5503));
  jand g05256(.dina(n5503), .dinb(n5500), .dout(n5504));
  jand g05257(.dina(n5504), .dinb(n5495), .dout(n5505));
  jor  g05258(.dina(n5505), .dinb(n5493), .dout(n5506));
  jand g05259(.dina(n5506), .dinb(asqrt[39] ), .dout(n5507));
  jor  g05260(.dina(n5506), .dinb(asqrt[39] ), .dout(n5508));
  jxor g05261(.dina(n5164), .dinb(n3907), .dout(n5509));
  jand g05262(.dina(n5509), .dinb(asqrt[32] ), .dout(n5510));
  jxor g05263(.dina(n5510), .dinb(n5169), .dout(n5511));
  jand g05264(.dina(n5511), .dinb(n5508), .dout(n5512));
  jor  g05265(.dina(n5512), .dinb(n5507), .dout(n5513));
  jand g05266(.dina(n5513), .dinb(asqrt[40] ), .dout(n5514));
  jnot g05267(.din(n5175), .dout(n5515));
  jand g05268(.dina(n5515), .dinb(n5173), .dout(n5516));
  jand g05269(.dina(n5516), .dinb(asqrt[32] ), .dout(n5517));
  jxor g05270(.dina(n5517), .dinb(n5183), .dout(n5518));
  jnot g05271(.din(n5518), .dout(n5519));
  jor  g05272(.dina(n5507), .dinb(asqrt[40] ), .dout(n5520));
  jor  g05273(.dina(n5520), .dinb(n5512), .dout(n5521));
  jand g05274(.dina(n5521), .dinb(n5519), .dout(n5522));
  jor  g05275(.dina(n5522), .dinb(n5514), .dout(n5523));
  jand g05276(.dina(n5523), .dinb(asqrt[41] ), .dout(n5524));
  jor  g05277(.dina(n5523), .dinb(asqrt[41] ), .dout(n5525));
  jxor g05278(.dina(n5185), .dinb(n3371), .dout(n5526));
  jand g05279(.dina(n5526), .dinb(asqrt[32] ), .dout(n5527));
  jxor g05280(.dina(n5527), .dinb(n5191), .dout(n5528));
  jand g05281(.dina(n5528), .dinb(n5525), .dout(n5529));
  jor  g05282(.dina(n5529), .dinb(n5524), .dout(n5530));
  jand g05283(.dina(n5530), .dinb(asqrt[42] ), .dout(n5531));
  jor  g05284(.dina(n5524), .dinb(asqrt[42] ), .dout(n5532));
  jor  g05285(.dina(n5532), .dinb(n5529), .dout(n5533));
  jnot g05286(.din(n5199), .dout(n5534));
  jnot g05287(.din(n5201), .dout(n5535));
  jand g05288(.dina(asqrt[32] ), .dinb(n5195), .dout(n5536));
  jand g05289(.dina(n5536), .dinb(n5535), .dout(n5537));
  jor  g05290(.dina(n5537), .dinb(n5534), .dout(n5538));
  jnot g05291(.din(n5202), .dout(n5539));
  jand g05292(.dina(n5536), .dinb(n5539), .dout(n5540));
  jnot g05293(.din(n5540), .dout(n5541));
  jand g05294(.dina(n5541), .dinb(n5538), .dout(n5542));
  jand g05295(.dina(n5542), .dinb(n5533), .dout(n5543));
  jor  g05296(.dina(n5543), .dinb(n5531), .dout(n5544));
  jand g05297(.dina(n5544), .dinb(asqrt[43] ), .dout(n5545));
  jxor g05298(.dina(n5203), .dinb(n2870), .dout(n5546));
  jand g05299(.dina(n5546), .dinb(asqrt[32] ), .dout(n5547));
  jxor g05300(.dina(n5547), .dinb(n5210), .dout(n5548));
  jnot g05301(.din(n5548), .dout(n5549));
  jor  g05302(.dina(n5544), .dinb(asqrt[43] ), .dout(n5550));
  jand g05303(.dina(n5550), .dinb(n5549), .dout(n5551));
  jor  g05304(.dina(n5551), .dinb(n5545), .dout(n5552));
  jand g05305(.dina(n5552), .dinb(asqrt[44] ), .dout(n5553));
  jnot g05306(.din(n5215), .dout(n5554));
  jand g05307(.dina(n5554), .dinb(n5213), .dout(n5555));
  jand g05308(.dina(n5555), .dinb(asqrt[32] ), .dout(n5556));
  jxor g05309(.dina(n5556), .dinb(n5223), .dout(n5557));
  jnot g05310(.din(n5557), .dout(n5558));
  jor  g05311(.dina(n5545), .dinb(asqrt[44] ), .dout(n5559));
  jor  g05312(.dina(n5559), .dinb(n5551), .dout(n5560));
  jand g05313(.dina(n5560), .dinb(n5558), .dout(n5561));
  jor  g05314(.dina(n5561), .dinb(n5553), .dout(n5562));
  jand g05315(.dina(n5562), .dinb(asqrt[45] ), .dout(n5563));
  jor  g05316(.dina(n5562), .dinb(asqrt[45] ), .dout(n5564));
  jnot g05317(.din(n5229), .dout(n5565));
  jnot g05318(.din(n5230), .dout(n5566));
  jand g05319(.dina(asqrt[32] ), .dinb(n5226), .dout(n5567));
  jand g05320(.dina(n5567), .dinb(n5566), .dout(n5568));
  jor  g05321(.dina(n5568), .dinb(n5565), .dout(n5569));
  jnot g05322(.din(n5231), .dout(n5570));
  jand g05323(.dina(n5567), .dinb(n5570), .dout(n5571));
  jnot g05324(.din(n5571), .dout(n5572));
  jand g05325(.dina(n5572), .dinb(n5569), .dout(n5573));
  jand g05326(.dina(n5573), .dinb(n5564), .dout(n5574));
  jor  g05327(.dina(n5574), .dinb(n5563), .dout(n5575));
  jand g05328(.dina(n5575), .dinb(asqrt[46] ), .dout(n5576));
  jor  g05329(.dina(n5563), .dinb(asqrt[46] ), .dout(n5577));
  jor  g05330(.dina(n5577), .dinb(n5574), .dout(n5578));
  jnot g05331(.din(n5237), .dout(n5579));
  jnot g05332(.din(n5239), .dout(n5580));
  jand g05333(.dina(asqrt[32] ), .dinb(n5233), .dout(n5581));
  jand g05334(.dina(n5581), .dinb(n5580), .dout(n5582));
  jor  g05335(.dina(n5582), .dinb(n5579), .dout(n5583));
  jnot g05336(.din(n5240), .dout(n5584));
  jand g05337(.dina(n5581), .dinb(n5584), .dout(n5585));
  jnot g05338(.din(n5585), .dout(n5586));
  jand g05339(.dina(n5586), .dinb(n5583), .dout(n5587));
  jand g05340(.dina(n5587), .dinb(n5578), .dout(n5588));
  jor  g05341(.dina(n5588), .dinb(n5576), .dout(n5589));
  jand g05342(.dina(n5589), .dinb(asqrt[47] ), .dout(n5590));
  jxor g05343(.dina(n5241), .dinb(n2005), .dout(n5591));
  jand g05344(.dina(n5591), .dinb(asqrt[32] ), .dout(n5592));
  jxor g05345(.dina(n5592), .dinb(n5251), .dout(n5593));
  jnot g05346(.din(n5593), .dout(n5594));
  jor  g05347(.dina(n5589), .dinb(asqrt[47] ), .dout(n5595));
  jand g05348(.dina(n5595), .dinb(n5594), .dout(n5596));
  jor  g05349(.dina(n5596), .dinb(n5590), .dout(n5597));
  jand g05350(.dina(n5597), .dinb(asqrt[48] ), .dout(n5598));
  jnot g05351(.din(n5256), .dout(n5599));
  jand g05352(.dina(n5599), .dinb(n5254), .dout(n5600));
  jand g05353(.dina(n5600), .dinb(asqrt[32] ), .dout(n5601));
  jxor g05354(.dina(n5601), .dinb(n5264), .dout(n5602));
  jnot g05355(.din(n5602), .dout(n5603));
  jor  g05356(.dina(n5590), .dinb(asqrt[48] ), .dout(n5604));
  jor  g05357(.dina(n5604), .dinb(n5596), .dout(n5605));
  jand g05358(.dina(n5605), .dinb(n5603), .dout(n5606));
  jor  g05359(.dina(n5606), .dinb(n5598), .dout(n5607));
  jand g05360(.dina(n5607), .dinb(asqrt[49] ), .dout(n5608));
  jor  g05361(.dina(n5607), .dinb(asqrt[49] ), .dout(n5609));
  jnot g05362(.din(n5270), .dout(n5610));
  jnot g05363(.din(n5271), .dout(n5611));
  jand g05364(.dina(asqrt[32] ), .dinb(n5267), .dout(n5612));
  jand g05365(.dina(n5612), .dinb(n5611), .dout(n5613));
  jor  g05366(.dina(n5613), .dinb(n5610), .dout(n5614));
  jnot g05367(.din(n5272), .dout(n5615));
  jand g05368(.dina(n5612), .dinb(n5615), .dout(n5616));
  jnot g05369(.din(n5616), .dout(n5617));
  jand g05370(.dina(n5617), .dinb(n5614), .dout(n5618));
  jand g05371(.dina(n5618), .dinb(n5609), .dout(n5619));
  jor  g05372(.dina(n5619), .dinb(n5608), .dout(n5620));
  jand g05373(.dina(n5620), .dinb(asqrt[50] ), .dout(n5621));
  jor  g05374(.dina(n5608), .dinb(asqrt[50] ), .dout(n5622));
  jor  g05375(.dina(n5622), .dinb(n5619), .dout(n5623));
  jnot g05376(.din(n5278), .dout(n5624));
  jnot g05377(.din(n5280), .dout(n5625));
  jand g05378(.dina(asqrt[32] ), .dinb(n5274), .dout(n5626));
  jand g05379(.dina(n5626), .dinb(n5625), .dout(n5627));
  jor  g05380(.dina(n5627), .dinb(n5624), .dout(n5628));
  jnot g05381(.din(n5281), .dout(n5629));
  jand g05382(.dina(n5626), .dinb(n5629), .dout(n5630));
  jnot g05383(.din(n5630), .dout(n5631));
  jand g05384(.dina(n5631), .dinb(n5628), .dout(n5632));
  jand g05385(.dina(n5632), .dinb(n5623), .dout(n5633));
  jor  g05386(.dina(n5633), .dinb(n5621), .dout(n5634));
  jand g05387(.dina(n5634), .dinb(asqrt[51] ), .dout(n5635));
  jxor g05388(.dina(n5282), .dinb(n1312), .dout(n5636));
  jand g05389(.dina(n5636), .dinb(asqrt[32] ), .dout(n5637));
  jxor g05390(.dina(n5637), .dinb(n5292), .dout(n5638));
  jnot g05391(.din(n5638), .dout(n5639));
  jor  g05392(.dina(n5634), .dinb(asqrt[51] ), .dout(n5640));
  jand g05393(.dina(n5640), .dinb(n5639), .dout(n5641));
  jor  g05394(.dina(n5641), .dinb(n5635), .dout(n5642));
  jand g05395(.dina(n5642), .dinb(asqrt[52] ), .dout(n5643));
  jnot g05396(.din(n5297), .dout(n5644));
  jand g05397(.dina(n5644), .dinb(n5295), .dout(n5645));
  jand g05398(.dina(n5645), .dinb(asqrt[32] ), .dout(n5646));
  jxor g05399(.dina(n5646), .dinb(n5305), .dout(n5647));
  jnot g05400(.din(n5647), .dout(n5648));
  jor  g05401(.dina(n5635), .dinb(asqrt[52] ), .dout(n5649));
  jor  g05402(.dina(n5649), .dinb(n5641), .dout(n5650));
  jand g05403(.dina(n5650), .dinb(n5648), .dout(n5651));
  jor  g05404(.dina(n5651), .dinb(n5643), .dout(n5652));
  jand g05405(.dina(n5652), .dinb(asqrt[53] ), .dout(n5653));
  jor  g05406(.dina(n5652), .dinb(asqrt[53] ), .dout(n5654));
  jnot g05407(.din(n5311), .dout(n5655));
  jnot g05408(.din(n5312), .dout(n5656));
  jand g05409(.dina(asqrt[32] ), .dinb(n5308), .dout(n5657));
  jand g05410(.dina(n5657), .dinb(n5656), .dout(n5658));
  jor  g05411(.dina(n5658), .dinb(n5655), .dout(n5659));
  jnot g05412(.din(n5313), .dout(n5660));
  jand g05413(.dina(n5657), .dinb(n5660), .dout(n5661));
  jnot g05414(.din(n5661), .dout(n5662));
  jand g05415(.dina(n5662), .dinb(n5659), .dout(n5663));
  jand g05416(.dina(n5663), .dinb(n5654), .dout(n5664));
  jor  g05417(.dina(n5664), .dinb(n5653), .dout(n5665));
  jand g05418(.dina(n5665), .dinb(asqrt[54] ), .dout(n5666));
  jor  g05419(.dina(n5653), .dinb(asqrt[54] ), .dout(n5667));
  jor  g05420(.dina(n5667), .dinb(n5664), .dout(n5668));
  jnot g05421(.din(n5319), .dout(n5669));
  jnot g05422(.din(n5321), .dout(n5670));
  jand g05423(.dina(asqrt[32] ), .dinb(n5315), .dout(n5671));
  jand g05424(.dina(n5671), .dinb(n5670), .dout(n5672));
  jor  g05425(.dina(n5672), .dinb(n5669), .dout(n5673));
  jnot g05426(.din(n5322), .dout(n5674));
  jand g05427(.dina(n5671), .dinb(n5674), .dout(n5675));
  jnot g05428(.din(n5675), .dout(n5676));
  jand g05429(.dina(n5676), .dinb(n5673), .dout(n5677));
  jand g05430(.dina(n5677), .dinb(n5668), .dout(n5678));
  jor  g05431(.dina(n5678), .dinb(n5666), .dout(n5679));
  jand g05432(.dina(n5679), .dinb(asqrt[55] ), .dout(n5680));
  jxor g05433(.dina(n5323), .dinb(n791), .dout(n5681));
  jand g05434(.dina(n5681), .dinb(asqrt[32] ), .dout(n5682));
  jxor g05435(.dina(n5682), .dinb(n5333), .dout(n5683));
  jnot g05436(.din(n5683), .dout(n5684));
  jor  g05437(.dina(n5679), .dinb(asqrt[55] ), .dout(n5685));
  jand g05438(.dina(n5685), .dinb(n5684), .dout(n5686));
  jor  g05439(.dina(n5686), .dinb(n5680), .dout(n5687));
  jand g05440(.dina(n5687), .dinb(asqrt[56] ), .dout(n5688));
  jnot g05441(.din(n5338), .dout(n5689));
  jand g05442(.dina(n5689), .dinb(n5336), .dout(n5690));
  jand g05443(.dina(n5690), .dinb(asqrt[32] ), .dout(n5691));
  jxor g05444(.dina(n5691), .dinb(n5346), .dout(n5692));
  jnot g05445(.din(n5692), .dout(n5693));
  jor  g05446(.dina(n5680), .dinb(asqrt[56] ), .dout(n5694));
  jor  g05447(.dina(n5694), .dinb(n5686), .dout(n5695));
  jand g05448(.dina(n5695), .dinb(n5693), .dout(n5696));
  jor  g05449(.dina(n5696), .dinb(n5688), .dout(n5697));
  jand g05450(.dina(n5697), .dinb(asqrt[57] ), .dout(n5698));
  jor  g05451(.dina(n5697), .dinb(asqrt[57] ), .dout(n5699));
  jnot g05452(.din(n5352), .dout(n5700));
  jnot g05453(.din(n5353), .dout(n5701));
  jand g05454(.dina(asqrt[32] ), .dinb(n5349), .dout(n5702));
  jand g05455(.dina(n5702), .dinb(n5701), .dout(n5703));
  jor  g05456(.dina(n5703), .dinb(n5700), .dout(n5704));
  jnot g05457(.din(n5354), .dout(n5705));
  jand g05458(.dina(n5702), .dinb(n5705), .dout(n5706));
  jnot g05459(.din(n5706), .dout(n5707));
  jand g05460(.dina(n5707), .dinb(n5704), .dout(n5708));
  jand g05461(.dina(n5708), .dinb(n5699), .dout(n5709));
  jor  g05462(.dina(n5709), .dinb(n5698), .dout(n5710));
  jand g05463(.dina(n5710), .dinb(asqrt[58] ), .dout(n5711));
  jor  g05464(.dina(n5698), .dinb(asqrt[58] ), .dout(n5712));
  jor  g05465(.dina(n5712), .dinb(n5709), .dout(n5713));
  jnot g05466(.din(n5360), .dout(n5714));
  jnot g05467(.din(n5362), .dout(n5715));
  jand g05468(.dina(asqrt[32] ), .dinb(n5356), .dout(n5716));
  jand g05469(.dina(n5716), .dinb(n5715), .dout(n5717));
  jor  g05470(.dina(n5717), .dinb(n5714), .dout(n5718));
  jnot g05471(.din(n5363), .dout(n5719));
  jand g05472(.dina(n5716), .dinb(n5719), .dout(n5720));
  jnot g05473(.din(n5720), .dout(n5721));
  jand g05474(.dina(n5721), .dinb(n5718), .dout(n5722));
  jand g05475(.dina(n5722), .dinb(n5713), .dout(n5723));
  jor  g05476(.dina(n5723), .dinb(n5711), .dout(n5724));
  jand g05477(.dina(n5724), .dinb(asqrt[59] ), .dout(n5725));
  jxor g05478(.dina(n5364), .dinb(n425), .dout(n5726));
  jand g05479(.dina(n5726), .dinb(asqrt[32] ), .dout(n5727));
  jxor g05480(.dina(n5727), .dinb(n5374), .dout(n5728));
  jnot g05481(.din(n5728), .dout(n5729));
  jor  g05482(.dina(n5724), .dinb(asqrt[59] ), .dout(n5730));
  jand g05483(.dina(n5730), .dinb(n5729), .dout(n5731));
  jor  g05484(.dina(n5731), .dinb(n5725), .dout(n5732));
  jand g05485(.dina(n5732), .dinb(asqrt[60] ), .dout(n5733));
  jnot g05486(.din(n5379), .dout(n5734));
  jand g05487(.dina(n5734), .dinb(n5377), .dout(n5735));
  jand g05488(.dina(n5735), .dinb(asqrt[32] ), .dout(n5736));
  jxor g05489(.dina(n5736), .dinb(n5387), .dout(n5737));
  jnot g05490(.din(n5737), .dout(n5738));
  jor  g05491(.dina(n5725), .dinb(asqrt[60] ), .dout(n5739));
  jor  g05492(.dina(n5739), .dinb(n5731), .dout(n5740));
  jand g05493(.dina(n5740), .dinb(n5738), .dout(n5741));
  jor  g05494(.dina(n5741), .dinb(n5733), .dout(n5742));
  jand g05495(.dina(n5742), .dinb(asqrt[61] ), .dout(n5743));
  jor  g05496(.dina(n5742), .dinb(asqrt[61] ), .dout(n5744));
  jnot g05497(.din(n5393), .dout(n5745));
  jnot g05498(.din(n5394), .dout(n5746));
  jand g05499(.dina(asqrt[32] ), .dinb(n5390), .dout(n5747));
  jand g05500(.dina(n5747), .dinb(n5746), .dout(n5748));
  jor  g05501(.dina(n5748), .dinb(n5745), .dout(n5749));
  jnot g05502(.din(n5395), .dout(n5750));
  jand g05503(.dina(n5747), .dinb(n5750), .dout(n5751));
  jnot g05504(.din(n5751), .dout(n5752));
  jand g05505(.dina(n5752), .dinb(n5749), .dout(n5753));
  jand g05506(.dina(n5753), .dinb(n5744), .dout(n5754));
  jor  g05507(.dina(n5754), .dinb(n5743), .dout(n5755));
  jand g05508(.dina(n5755), .dinb(asqrt[62] ), .dout(n5756));
  jor  g05509(.dina(n5743), .dinb(asqrt[62] ), .dout(n5757));
  jor  g05510(.dina(n5757), .dinb(n5754), .dout(n5758));
  jnot g05511(.din(n5401), .dout(n5759));
  jnot g05512(.din(n5403), .dout(n5760));
  jand g05513(.dina(asqrt[32] ), .dinb(n5397), .dout(n5761));
  jand g05514(.dina(n5761), .dinb(n5760), .dout(n5762));
  jor  g05515(.dina(n5762), .dinb(n5759), .dout(n5763));
  jnot g05516(.din(n5404), .dout(n5764));
  jand g05517(.dina(n5761), .dinb(n5764), .dout(n5765));
  jnot g05518(.din(n5765), .dout(n5766));
  jand g05519(.dina(n5766), .dinb(n5763), .dout(n5767));
  jand g05520(.dina(n5767), .dinb(n5758), .dout(n5768));
  jor  g05521(.dina(n5768), .dinb(n5756), .dout(n5769));
  jxor g05522(.dina(n5405), .dinb(n199), .dout(n5770));
  jand g05523(.dina(n5770), .dinb(asqrt[32] ), .dout(n5771));
  jxor g05524(.dina(n5771), .dinb(n5415), .dout(n5772));
  jnot g05525(.din(n5417), .dout(n5773));
  jand g05526(.dina(asqrt[32] ), .dinb(n5424), .dout(n5774));
  jand g05527(.dina(n5774), .dinb(n5773), .dout(n5775));
  jor  g05528(.dina(n5775), .dinb(n5432), .dout(n5776));
  jor  g05529(.dina(n5776), .dinb(n5772), .dout(n5777));
  jnot g05530(.din(n5777), .dout(n5778));
  jand g05531(.dina(n5778), .dinb(n5769), .dout(n5779));
  jor  g05532(.dina(n5779), .dinb(asqrt[63] ), .dout(n5780));
  jnot g05533(.din(n5772), .dout(n5781));
  jor  g05534(.dina(n5781), .dinb(n5769), .dout(n5782));
  jor  g05535(.dina(n5774), .dinb(n5773), .dout(n5783));
  jand g05536(.dina(n5424), .dinb(n5773), .dout(n5784));
  jor  g05537(.dina(n5784), .dinb(n194), .dout(n5785));
  jnot g05538(.din(n5785), .dout(n5786));
  jand g05539(.dina(n5786), .dinb(n5783), .dout(n5787));
  jnot g05540(.din(asqrt[32] ), .dout(n5788));
  jnot g05541(.din(n5787), .dout(n5791));
  jand g05542(.dina(n5791), .dinb(n5782), .dout(n5792));
  jand g05543(.dina(n5792), .dinb(n5780), .dout(n5793));
  jor  g05544(.dina(n5793), .dinb(a[62] ), .dout(n5794));
  jxor g05545(.dina(n5794), .dinb(n200), .dout(n5795));
  jor  g05546(.dina(n5793), .dinb(n5443), .dout(n5796));
  jnot g05547(.din(a[60] ), .dout(n5797));
  jnot g05548(.din(a[61] ), .dout(n5798));
  jand g05549(.dina(n5443), .dinb(n5798), .dout(n5799));
  jand g05550(.dina(n5799), .dinb(n5797), .dout(n5800));
  jnot g05551(.din(n5800), .dout(n5801));
  jand g05552(.dina(n5801), .dinb(n5796), .dout(n5802));
  jor  g05553(.dina(n5802), .dinb(n5788), .dout(n5803));
  jand g05554(.dina(n5802), .dinb(n5788), .dout(n5804));
  jor  g05555(.dina(n5804), .dinb(n5795), .dout(n5805));
  jand g05556(.dina(n5805), .dinb(n5803), .dout(n5806));
  jor  g05557(.dina(n5806), .dinb(n5121), .dout(n5807));
  jor  g05558(.dina(n5794), .dinb(a[63] ), .dout(n5808));
  jnot g05559(.din(n5780), .dout(n5809));
  jnot g05560(.din(n5782), .dout(n5810));
  jor  g05561(.dina(n5787), .dinb(n5788), .dout(n5811));
  jor  g05562(.dina(n5811), .dinb(n5810), .dout(n5812));
  jor  g05563(.dina(n5812), .dinb(n5809), .dout(n5813));
  jand g05564(.dina(n5813), .dinb(n5808), .dout(n5814));
  jxor g05565(.dina(n5814), .dinb(n5124), .dout(n5815));
  jand g05566(.dina(n5803), .dinb(n5121), .dout(n5816));
  jand g05567(.dina(n5816), .dinb(n5805), .dout(n5817));
  jor  g05568(.dina(n5817), .dinb(n5815), .dout(n5818));
  jand g05569(.dina(n5818), .dinb(n5807), .dout(n5819));
  jor  g05570(.dina(n5819), .dinb(n5116), .dout(n5820));
  jand g05571(.dina(n5819), .dinb(n5116), .dout(n5821));
  jxor g05572(.dina(n5446), .dinb(n5121), .dout(n5822));
  jor  g05573(.dina(n5822), .dinb(n5793), .dout(n5823));
  jxor g05574(.dina(n5823), .dinb(n5449), .dout(n5824));
  jor  g05575(.dina(n5824), .dinb(n5821), .dout(n5825));
  jand g05576(.dina(n5825), .dinb(n5820), .dout(n5826));
  jor  g05577(.dina(n5826), .dinb(n4499), .dout(n5827));
  jnot g05578(.din(n5455), .dout(n5828));
  jor  g05579(.dina(n5828), .dinb(n5453), .dout(n5829));
  jor  g05580(.dina(n5829), .dinb(n5793), .dout(n5830));
  jxor g05581(.dina(n5830), .dinb(n5464), .dout(n5831));
  jand g05582(.dina(n5820), .dinb(n4499), .dout(n5832));
  jand g05583(.dina(n5832), .dinb(n5825), .dout(n5833));
  jor  g05584(.dina(n5833), .dinb(n5831), .dout(n5834));
  jand g05585(.dina(n5834), .dinb(n5827), .dout(n5835));
  jor  g05586(.dina(n5835), .dinb(n4494), .dout(n5836));
  jand g05587(.dina(n5835), .dinb(n4494), .dout(n5837));
  jxor g05588(.dina(n5466), .dinb(n4499), .dout(n5838));
  jor  g05589(.dina(n5838), .dinb(n5793), .dout(n5839));
  jxor g05590(.dina(n5839), .dinb(n5471), .dout(n5840));
  jnot g05591(.din(n5840), .dout(n5841));
  jor  g05592(.dina(n5841), .dinb(n5837), .dout(n5842));
  jand g05593(.dina(n5842), .dinb(n5836), .dout(n5843));
  jor  g05594(.dina(n5843), .dinb(n3912), .dout(n5844));
  jand g05595(.dina(n5836), .dinb(n3912), .dout(n5845));
  jand g05596(.dina(n5845), .dinb(n5842), .dout(n5846));
  jnot g05597(.din(n5475), .dout(n5847));
  jnot g05598(.din(n5793), .dout(asqrt[31] ));
  jand g05599(.dina(asqrt[31] ), .dinb(n5847), .dout(n5849));
  jand g05600(.dina(n5849), .dinb(n5482), .dout(n5850));
  jor  g05601(.dina(n5850), .dinb(n5480), .dout(n5851));
  jand g05602(.dina(n5849), .dinb(n5483), .dout(n5852));
  jnot g05603(.din(n5852), .dout(n5853));
  jand g05604(.dina(n5853), .dinb(n5851), .dout(n5854));
  jnot g05605(.din(n5854), .dout(n5855));
  jor  g05606(.dina(n5855), .dinb(n5846), .dout(n5856));
  jand g05607(.dina(n5856), .dinb(n5844), .dout(n5857));
  jor  g05608(.dina(n5857), .dinb(n3907), .dout(n5858));
  jand g05609(.dina(n5857), .dinb(n3907), .dout(n5859));
  jnot g05610(.din(n5490), .dout(n5860));
  jxor g05611(.dina(n5484), .dinb(n3912), .dout(n5861));
  jor  g05612(.dina(n5861), .dinb(n5793), .dout(n5862));
  jxor g05613(.dina(n5862), .dinb(n5860), .dout(n5863));
  jnot g05614(.din(n5863), .dout(n5864));
  jor  g05615(.dina(n5864), .dinb(n5859), .dout(n5865));
  jand g05616(.dina(n5865), .dinb(n5858), .dout(n5866));
  jor  g05617(.dina(n5866), .dinb(n3376), .dout(n5867));
  jnot g05618(.din(n5495), .dout(n5868));
  jor  g05619(.dina(n5868), .dinb(n5493), .dout(n5869));
  jor  g05620(.dina(n5869), .dinb(n5793), .dout(n5870));
  jxor g05621(.dina(n5870), .dinb(n5504), .dout(n5871));
  jand g05622(.dina(n5858), .dinb(n3376), .dout(n5872));
  jand g05623(.dina(n5872), .dinb(n5865), .dout(n5873));
  jor  g05624(.dina(n5873), .dinb(n5871), .dout(n5874));
  jand g05625(.dina(n5874), .dinb(n5867), .dout(n5875));
  jor  g05626(.dina(n5875), .dinb(n3371), .dout(n5876));
  jand g05627(.dina(n5875), .dinb(n3371), .dout(n5877));
  jnot g05628(.din(n5511), .dout(n5878));
  jxor g05629(.dina(n5506), .dinb(n3376), .dout(n5879));
  jor  g05630(.dina(n5879), .dinb(n5793), .dout(n5880));
  jxor g05631(.dina(n5880), .dinb(n5878), .dout(n5881));
  jnot g05632(.din(n5881), .dout(n5882));
  jor  g05633(.dina(n5882), .dinb(n5877), .dout(n5883));
  jand g05634(.dina(n5883), .dinb(n5876), .dout(n5884));
  jor  g05635(.dina(n5884), .dinb(n2875), .dout(n5885));
  jand g05636(.dina(n5876), .dinb(n2875), .dout(n5886));
  jand g05637(.dina(n5886), .dinb(n5883), .dout(n5887));
  jnot g05638(.din(n5514), .dout(n5888));
  jand g05639(.dina(asqrt[31] ), .dinb(n5888), .dout(n5889));
  jand g05640(.dina(n5889), .dinb(n5521), .dout(n5890));
  jor  g05641(.dina(n5890), .dinb(n5519), .dout(n5891));
  jand g05642(.dina(n5889), .dinb(n5522), .dout(n5892));
  jnot g05643(.din(n5892), .dout(n5893));
  jand g05644(.dina(n5893), .dinb(n5891), .dout(n5894));
  jnot g05645(.din(n5894), .dout(n5895));
  jor  g05646(.dina(n5895), .dinb(n5887), .dout(n5896));
  jand g05647(.dina(n5896), .dinb(n5885), .dout(n5897));
  jor  g05648(.dina(n5897), .dinb(n2870), .dout(n5898));
  jxor g05649(.dina(n5523), .dinb(n2875), .dout(n5899));
  jor  g05650(.dina(n5899), .dinb(n5793), .dout(n5900));
  jxor g05651(.dina(n5900), .dinb(n5528), .dout(n5901));
  jand g05652(.dina(n5897), .dinb(n2870), .dout(n5902));
  jor  g05653(.dina(n5902), .dinb(n5901), .dout(n5903));
  jand g05654(.dina(n5903), .dinb(n5898), .dout(n5904));
  jor  g05655(.dina(n5904), .dinb(n2425), .dout(n5905));
  jnot g05656(.din(n5533), .dout(n5906));
  jor  g05657(.dina(n5906), .dinb(n5531), .dout(n5907));
  jor  g05658(.dina(n5907), .dinb(n5793), .dout(n5908));
  jxor g05659(.dina(n5908), .dinb(n5542), .dout(n5909));
  jand g05660(.dina(n5898), .dinb(n2425), .dout(n5910));
  jand g05661(.dina(n5910), .dinb(n5903), .dout(n5911));
  jor  g05662(.dina(n5911), .dinb(n5909), .dout(n5912));
  jand g05663(.dina(n5912), .dinb(n5905), .dout(n5913));
  jor  g05664(.dina(n5913), .dinb(n2420), .dout(n5914));
  jand g05665(.dina(n5913), .dinb(n2420), .dout(n5915));
  jnot g05666(.din(n5545), .dout(n5916));
  jand g05667(.dina(asqrt[31] ), .dinb(n5916), .dout(n5917));
  jand g05668(.dina(n5917), .dinb(n5550), .dout(n5918));
  jor  g05669(.dina(n5918), .dinb(n5549), .dout(n5919));
  jand g05670(.dina(n5917), .dinb(n5551), .dout(n5920));
  jnot g05671(.din(n5920), .dout(n5921));
  jand g05672(.dina(n5921), .dinb(n5919), .dout(n5922));
  jnot g05673(.din(n5922), .dout(n5923));
  jor  g05674(.dina(n5923), .dinb(n5915), .dout(n5924));
  jand g05675(.dina(n5924), .dinb(n5914), .dout(n5925));
  jor  g05676(.dina(n5925), .dinb(n2010), .dout(n5926));
  jand g05677(.dina(n5914), .dinb(n2010), .dout(n5927));
  jand g05678(.dina(n5927), .dinb(n5924), .dout(n5928));
  jnot g05679(.din(n5553), .dout(n5929));
  jand g05680(.dina(asqrt[31] ), .dinb(n5929), .dout(n5930));
  jand g05681(.dina(n5930), .dinb(n5560), .dout(n5931));
  jor  g05682(.dina(n5931), .dinb(n5558), .dout(n5932));
  jand g05683(.dina(n5930), .dinb(n5561), .dout(n5933));
  jnot g05684(.din(n5933), .dout(n5934));
  jand g05685(.dina(n5934), .dinb(n5932), .dout(n5935));
  jnot g05686(.din(n5935), .dout(n5936));
  jor  g05687(.dina(n5936), .dinb(n5928), .dout(n5937));
  jand g05688(.dina(n5937), .dinb(n5926), .dout(n5938));
  jor  g05689(.dina(n5938), .dinb(n2005), .dout(n5939));
  jxor g05690(.dina(n5562), .dinb(n2010), .dout(n5940));
  jor  g05691(.dina(n5940), .dinb(n5793), .dout(n5941));
  jxor g05692(.dina(n5941), .dinb(n5573), .dout(n5942));
  jand g05693(.dina(n5938), .dinb(n2005), .dout(n5943));
  jor  g05694(.dina(n5943), .dinb(n5942), .dout(n5944));
  jand g05695(.dina(n5944), .dinb(n5939), .dout(n5945));
  jor  g05696(.dina(n5945), .dinb(n1646), .dout(n5946));
  jnot g05697(.din(n5578), .dout(n5947));
  jor  g05698(.dina(n5947), .dinb(n5576), .dout(n5948));
  jor  g05699(.dina(n5948), .dinb(n5793), .dout(n5949));
  jxor g05700(.dina(n5949), .dinb(n5587), .dout(n5950));
  jand g05701(.dina(n5939), .dinb(n1646), .dout(n5951));
  jand g05702(.dina(n5951), .dinb(n5944), .dout(n5952));
  jor  g05703(.dina(n5952), .dinb(n5950), .dout(n5953));
  jand g05704(.dina(n5953), .dinb(n5946), .dout(n5954));
  jor  g05705(.dina(n5954), .dinb(n1641), .dout(n5955));
  jand g05706(.dina(n5954), .dinb(n1641), .dout(n5956));
  jnot g05707(.din(n5590), .dout(n5957));
  jand g05708(.dina(asqrt[31] ), .dinb(n5957), .dout(n5958));
  jand g05709(.dina(n5958), .dinb(n5595), .dout(n5959));
  jor  g05710(.dina(n5959), .dinb(n5594), .dout(n5960));
  jand g05711(.dina(n5958), .dinb(n5596), .dout(n5961));
  jnot g05712(.din(n5961), .dout(n5962));
  jand g05713(.dina(n5962), .dinb(n5960), .dout(n5963));
  jnot g05714(.din(n5963), .dout(n5964));
  jor  g05715(.dina(n5964), .dinb(n5956), .dout(n5965));
  jand g05716(.dina(n5965), .dinb(n5955), .dout(n5966));
  jor  g05717(.dina(n5966), .dinb(n1317), .dout(n5967));
  jand g05718(.dina(n5955), .dinb(n1317), .dout(n5968));
  jand g05719(.dina(n5968), .dinb(n5965), .dout(n5969));
  jnot g05720(.din(n5598), .dout(n5970));
  jand g05721(.dina(asqrt[31] ), .dinb(n5970), .dout(n5971));
  jand g05722(.dina(n5971), .dinb(n5605), .dout(n5972));
  jor  g05723(.dina(n5972), .dinb(n5603), .dout(n5973));
  jand g05724(.dina(n5971), .dinb(n5606), .dout(n5974));
  jnot g05725(.din(n5974), .dout(n5975));
  jand g05726(.dina(n5975), .dinb(n5973), .dout(n5976));
  jnot g05727(.din(n5976), .dout(n5977));
  jor  g05728(.dina(n5977), .dinb(n5969), .dout(n5978));
  jand g05729(.dina(n5978), .dinb(n5967), .dout(n5979));
  jor  g05730(.dina(n5979), .dinb(n1312), .dout(n5980));
  jxor g05731(.dina(n5607), .dinb(n1317), .dout(n5981));
  jor  g05732(.dina(n5981), .dinb(n5793), .dout(n5982));
  jxor g05733(.dina(n5982), .dinb(n5618), .dout(n5983));
  jand g05734(.dina(n5979), .dinb(n1312), .dout(n5984));
  jor  g05735(.dina(n5984), .dinb(n5983), .dout(n5985));
  jand g05736(.dina(n5985), .dinb(n5980), .dout(n5986));
  jor  g05737(.dina(n5986), .dinb(n1039), .dout(n5987));
  jnot g05738(.din(n5623), .dout(n5988));
  jor  g05739(.dina(n5988), .dinb(n5621), .dout(n5989));
  jor  g05740(.dina(n5989), .dinb(n5793), .dout(n5990));
  jxor g05741(.dina(n5990), .dinb(n5632), .dout(n5991));
  jand g05742(.dina(n5980), .dinb(n1039), .dout(n5992));
  jand g05743(.dina(n5992), .dinb(n5985), .dout(n5993));
  jor  g05744(.dina(n5993), .dinb(n5991), .dout(n5994));
  jand g05745(.dina(n5994), .dinb(n5987), .dout(n5995));
  jor  g05746(.dina(n5995), .dinb(n1034), .dout(n5996));
  jand g05747(.dina(n5995), .dinb(n1034), .dout(n5997));
  jnot g05748(.din(n5635), .dout(n5998));
  jand g05749(.dina(asqrt[31] ), .dinb(n5998), .dout(n5999));
  jand g05750(.dina(n5999), .dinb(n5640), .dout(n6000));
  jor  g05751(.dina(n6000), .dinb(n5639), .dout(n6001));
  jand g05752(.dina(n5999), .dinb(n5641), .dout(n6002));
  jnot g05753(.din(n6002), .dout(n6003));
  jand g05754(.dina(n6003), .dinb(n6001), .dout(n6004));
  jnot g05755(.din(n6004), .dout(n6005));
  jor  g05756(.dina(n6005), .dinb(n5997), .dout(n6006));
  jand g05757(.dina(n6006), .dinb(n5996), .dout(n6007));
  jor  g05758(.dina(n6007), .dinb(n796), .dout(n6008));
  jand g05759(.dina(n5996), .dinb(n796), .dout(n6009));
  jand g05760(.dina(n6009), .dinb(n6006), .dout(n6010));
  jnot g05761(.din(n5643), .dout(n6011));
  jand g05762(.dina(asqrt[31] ), .dinb(n6011), .dout(n6012));
  jand g05763(.dina(n6012), .dinb(n5650), .dout(n6013));
  jor  g05764(.dina(n6013), .dinb(n5648), .dout(n6014));
  jand g05765(.dina(n6012), .dinb(n5651), .dout(n6015));
  jnot g05766(.din(n6015), .dout(n6016));
  jand g05767(.dina(n6016), .dinb(n6014), .dout(n6017));
  jnot g05768(.din(n6017), .dout(n6018));
  jor  g05769(.dina(n6018), .dinb(n6010), .dout(n6019));
  jand g05770(.dina(n6019), .dinb(n6008), .dout(n6020));
  jor  g05771(.dina(n6020), .dinb(n791), .dout(n6021));
  jxor g05772(.dina(n5652), .dinb(n796), .dout(n6022));
  jor  g05773(.dina(n6022), .dinb(n5793), .dout(n6023));
  jxor g05774(.dina(n6023), .dinb(n5663), .dout(n6024));
  jand g05775(.dina(n6020), .dinb(n791), .dout(n6025));
  jor  g05776(.dina(n6025), .dinb(n6024), .dout(n6026));
  jand g05777(.dina(n6026), .dinb(n6021), .dout(n6027));
  jor  g05778(.dina(n6027), .dinb(n595), .dout(n6028));
  jnot g05779(.din(n5668), .dout(n6029));
  jor  g05780(.dina(n6029), .dinb(n5666), .dout(n6030));
  jor  g05781(.dina(n6030), .dinb(n5793), .dout(n6031));
  jxor g05782(.dina(n6031), .dinb(n5677), .dout(n6032));
  jand g05783(.dina(n6021), .dinb(n595), .dout(n6033));
  jand g05784(.dina(n6033), .dinb(n6026), .dout(n6034));
  jor  g05785(.dina(n6034), .dinb(n6032), .dout(n6035));
  jand g05786(.dina(n6035), .dinb(n6028), .dout(n6036));
  jor  g05787(.dina(n6036), .dinb(n590), .dout(n6037));
  jand g05788(.dina(n6036), .dinb(n590), .dout(n6038));
  jnot g05789(.din(n5680), .dout(n6039));
  jand g05790(.dina(asqrt[31] ), .dinb(n6039), .dout(n6040));
  jand g05791(.dina(n6040), .dinb(n5685), .dout(n6041));
  jor  g05792(.dina(n6041), .dinb(n5684), .dout(n6042));
  jand g05793(.dina(n6040), .dinb(n5686), .dout(n6043));
  jnot g05794(.din(n6043), .dout(n6044));
  jand g05795(.dina(n6044), .dinb(n6042), .dout(n6045));
  jnot g05796(.din(n6045), .dout(n6046));
  jor  g05797(.dina(n6046), .dinb(n6038), .dout(n6047));
  jand g05798(.dina(n6047), .dinb(n6037), .dout(n6048));
  jor  g05799(.dina(n6048), .dinb(n430), .dout(n6049));
  jand g05800(.dina(n6037), .dinb(n430), .dout(n6050));
  jand g05801(.dina(n6050), .dinb(n6047), .dout(n6051));
  jnot g05802(.din(n5688), .dout(n6052));
  jand g05803(.dina(asqrt[31] ), .dinb(n6052), .dout(n6053));
  jand g05804(.dina(n6053), .dinb(n5695), .dout(n6054));
  jor  g05805(.dina(n6054), .dinb(n5693), .dout(n6055));
  jand g05806(.dina(n6053), .dinb(n5696), .dout(n6056));
  jnot g05807(.din(n6056), .dout(n6057));
  jand g05808(.dina(n6057), .dinb(n6055), .dout(n6058));
  jnot g05809(.din(n6058), .dout(n6059));
  jor  g05810(.dina(n6059), .dinb(n6051), .dout(n6060));
  jand g05811(.dina(n6060), .dinb(n6049), .dout(n6061));
  jor  g05812(.dina(n6061), .dinb(n425), .dout(n6062));
  jxor g05813(.dina(n5697), .dinb(n430), .dout(n6063));
  jor  g05814(.dina(n6063), .dinb(n5793), .dout(n6064));
  jxor g05815(.dina(n6064), .dinb(n5708), .dout(n6065));
  jand g05816(.dina(n6061), .dinb(n425), .dout(n6066));
  jor  g05817(.dina(n6066), .dinb(n6065), .dout(n6067));
  jand g05818(.dina(n6067), .dinb(n6062), .dout(n6068));
  jor  g05819(.dina(n6068), .dinb(n305), .dout(n6069));
  jnot g05820(.din(n5713), .dout(n6070));
  jor  g05821(.dina(n6070), .dinb(n5711), .dout(n6071));
  jor  g05822(.dina(n6071), .dinb(n5793), .dout(n6072));
  jxor g05823(.dina(n6072), .dinb(n5722), .dout(n6073));
  jand g05824(.dina(n6062), .dinb(n305), .dout(n6074));
  jand g05825(.dina(n6074), .dinb(n6067), .dout(n6075));
  jor  g05826(.dina(n6075), .dinb(n6073), .dout(n6076));
  jand g05827(.dina(n6076), .dinb(n6069), .dout(n6077));
  jor  g05828(.dina(n6077), .dinb(n290), .dout(n6078));
  jand g05829(.dina(n6077), .dinb(n290), .dout(n6079));
  jnot g05830(.din(n5725), .dout(n6080));
  jand g05831(.dina(asqrt[31] ), .dinb(n6080), .dout(n6081));
  jand g05832(.dina(n6081), .dinb(n5730), .dout(n6082));
  jor  g05833(.dina(n6082), .dinb(n5729), .dout(n6083));
  jand g05834(.dina(n6081), .dinb(n5731), .dout(n6084));
  jnot g05835(.din(n6084), .dout(n6085));
  jand g05836(.dina(n6085), .dinb(n6083), .dout(n6086));
  jnot g05837(.din(n6086), .dout(n6087));
  jor  g05838(.dina(n6087), .dinb(n6079), .dout(n6088));
  jand g05839(.dina(n6088), .dinb(n6078), .dout(n6089));
  jor  g05840(.dina(n6089), .dinb(n223), .dout(n6090));
  jand g05841(.dina(n6078), .dinb(n223), .dout(n6091));
  jand g05842(.dina(n6091), .dinb(n6088), .dout(n6092));
  jnot g05843(.din(n5733), .dout(n6093));
  jand g05844(.dina(asqrt[31] ), .dinb(n6093), .dout(n6094));
  jand g05845(.dina(n6094), .dinb(n5740), .dout(n6095));
  jor  g05846(.dina(n6095), .dinb(n5738), .dout(n6096));
  jand g05847(.dina(n6094), .dinb(n5741), .dout(n6097));
  jnot g05848(.din(n6097), .dout(n6098));
  jand g05849(.dina(n6098), .dinb(n6096), .dout(n6099));
  jnot g05850(.din(n6099), .dout(n6100));
  jor  g05851(.dina(n6100), .dinb(n6092), .dout(n6101));
  jand g05852(.dina(n6101), .dinb(n6090), .dout(n6102));
  jor  g05853(.dina(n6102), .dinb(n199), .dout(n6103));
  jand g05854(.dina(n6102), .dinb(n199), .dout(n6104));
  jxor g05855(.dina(n5742), .dinb(n223), .dout(n6105));
  jor  g05856(.dina(n6105), .dinb(n5793), .dout(n6106));
  jxor g05857(.dina(n6106), .dinb(n5753), .dout(n6107));
  jor  g05858(.dina(n6107), .dinb(n6104), .dout(n6108));
  jand g05859(.dina(n6108), .dinb(n6103), .dout(n6109));
  jnot g05860(.din(n5758), .dout(n6110));
  jor  g05861(.dina(n6110), .dinb(n5756), .dout(n6111));
  jor  g05862(.dina(n6111), .dinb(n5793), .dout(n6112));
  jxor g05863(.dina(n6112), .dinb(n5767), .dout(n6113));
  jand g05864(.dina(asqrt[31] ), .dinb(n5781), .dout(n6114));
  jand g05865(.dina(n6114), .dinb(n5769), .dout(n6115));
  jor  g05866(.dina(n6115), .dinb(n5810), .dout(n6116));
  jor  g05867(.dina(n6116), .dinb(n6113), .dout(n6117));
  jor  g05868(.dina(n6117), .dinb(n6109), .dout(n6118));
  jand g05869(.dina(n6118), .dinb(n194), .dout(n6119));
  jand g05870(.dina(n6113), .dinb(n6109), .dout(n6120));
  jor  g05871(.dina(n6114), .dinb(n5769), .dout(n6121));
  jand g05872(.dina(n5781), .dinb(n5769), .dout(n6122));
  jor  g05873(.dina(n6122), .dinb(n194), .dout(n6123));
  jnot g05874(.din(n6123), .dout(n6124));
  jand g05875(.dina(n6124), .dinb(n6121), .dout(n6125));
  jor  g05876(.dina(n6125), .dinb(n6120), .dout(n6128));
  jor  g05877(.dina(n6128), .dinb(n6119), .dout(asqrt[30] ));
  jxor g05878(.dina(n5802), .dinb(n5788), .dout(n6130));
  jand g05879(.dina(n6130), .dinb(asqrt[30] ), .dout(n6131));
  jxor g05880(.dina(n6131), .dinb(n5795), .dout(n6132));
  jand g05881(.dina(asqrt[30] ), .dinb(a[60] ), .dout(n6133));
  jnot g05882(.din(a[58] ), .dout(n6134));
  jnot g05883(.din(a[59] ), .dout(n6135));
  jand g05884(.dina(n5797), .dinb(n6135), .dout(n6136));
  jand g05885(.dina(n6136), .dinb(n6134), .dout(n6137));
  jor  g05886(.dina(n6137), .dinb(n6133), .dout(n6138));
  jand g05887(.dina(n6138), .dinb(asqrt[31] ), .dout(n6139));
  jand g05888(.dina(asqrt[30] ), .dinb(n5797), .dout(n6140));
  jxor g05889(.dina(n6140), .dinb(n5798), .dout(n6141));
  jor  g05890(.dina(n6138), .dinb(asqrt[31] ), .dout(n6142));
  jand g05891(.dina(n6142), .dinb(n6141), .dout(n6143));
  jor  g05892(.dina(n6143), .dinb(n6139), .dout(n6144));
  jand g05893(.dina(n6144), .dinb(asqrt[32] ), .dout(n6145));
  jand g05894(.dina(n6140), .dinb(n5798), .dout(n6146));
  jnot g05895(.din(n6119), .dout(n6147));
  jnot g05896(.din(n6120), .dout(n6148));
  jnot g05897(.din(n6125), .dout(n6149));
  jand g05898(.dina(n6149), .dinb(asqrt[31] ), .dout(n6150));
  jand g05899(.dina(n6150), .dinb(n6148), .dout(n6151));
  jand g05900(.dina(n6151), .dinb(n6147), .dout(n6152));
  jor  g05901(.dina(n6152), .dinb(n6146), .dout(n6153));
  jxor g05902(.dina(n6153), .dinb(n5443), .dout(n6154));
  jor  g05903(.dina(n6139), .dinb(asqrt[32] ), .dout(n6155));
  jor  g05904(.dina(n6155), .dinb(n6143), .dout(n6156));
  jand g05905(.dina(n6156), .dinb(n6154), .dout(n6157));
  jor  g05906(.dina(n6157), .dinb(n6145), .dout(n6158));
  jand g05907(.dina(n6158), .dinb(asqrt[33] ), .dout(n6159));
  jnot g05908(.din(n6132), .dout(n6160));
  jor  g05909(.dina(n6158), .dinb(asqrt[33] ), .dout(n6161));
  jand g05910(.dina(n6161), .dinb(n6160), .dout(n6162));
  jor  g05911(.dina(n6162), .dinb(n6159), .dout(n6163));
  jand g05912(.dina(n6163), .dinb(asqrt[34] ), .dout(n6164));
  jor  g05913(.dina(n6159), .dinb(asqrt[34] ), .dout(n6165));
  jor  g05914(.dina(n6165), .dinb(n6162), .dout(n6166));
  jnot g05915(.din(n5815), .dout(n6167));
  jnot g05916(.din(n5817), .dout(n6168));
  jand g05917(.dina(asqrt[30] ), .dinb(n5807), .dout(n6169));
  jand g05918(.dina(n6169), .dinb(n6168), .dout(n6170));
  jor  g05919(.dina(n6170), .dinb(n6167), .dout(n6171));
  jnot g05920(.din(n5818), .dout(n6172));
  jand g05921(.dina(n6169), .dinb(n6172), .dout(n6173));
  jnot g05922(.din(n6173), .dout(n6174));
  jand g05923(.dina(n6174), .dinb(n6171), .dout(n6175));
  jand g05924(.dina(n6175), .dinb(n6166), .dout(n6176));
  jor  g05925(.dina(n6176), .dinb(n6164), .dout(n6177));
  jand g05926(.dina(n6177), .dinb(asqrt[35] ), .dout(n6178));
  jor  g05927(.dina(n6177), .dinb(asqrt[35] ), .dout(n6179));
  jnot g05928(.din(n5824), .dout(n6180));
  jxor g05929(.dina(n5819), .dinb(n5116), .dout(n6181));
  jand g05930(.dina(n6181), .dinb(asqrt[30] ), .dout(n6182));
  jxor g05931(.dina(n6182), .dinb(n6180), .dout(n6183));
  jand g05932(.dina(n6183), .dinb(n6179), .dout(n6184));
  jor  g05933(.dina(n6184), .dinb(n6178), .dout(n6185));
  jand g05934(.dina(n6185), .dinb(asqrt[36] ), .dout(n6186));
  jor  g05935(.dina(n6178), .dinb(asqrt[36] ), .dout(n6187));
  jor  g05936(.dina(n6187), .dinb(n6184), .dout(n6188));
  jnot g05937(.din(n5831), .dout(n6189));
  jnot g05938(.din(n5833), .dout(n6190));
  jand g05939(.dina(asqrt[30] ), .dinb(n5827), .dout(n6191));
  jand g05940(.dina(n6191), .dinb(n6190), .dout(n6192));
  jor  g05941(.dina(n6192), .dinb(n6189), .dout(n6193));
  jnot g05942(.din(n5834), .dout(n6194));
  jand g05943(.dina(n6191), .dinb(n6194), .dout(n6195));
  jnot g05944(.din(n6195), .dout(n6196));
  jand g05945(.dina(n6196), .dinb(n6193), .dout(n6197));
  jand g05946(.dina(n6197), .dinb(n6188), .dout(n6198));
  jor  g05947(.dina(n6198), .dinb(n6186), .dout(n6199));
  jand g05948(.dina(n6199), .dinb(asqrt[37] ), .dout(n6200));
  jor  g05949(.dina(n6199), .dinb(asqrt[37] ), .dout(n6201));
  jxor g05950(.dina(n5835), .dinb(n4494), .dout(n6202));
  jand g05951(.dina(n6202), .dinb(asqrt[30] ), .dout(n6203));
  jxor g05952(.dina(n6203), .dinb(n5840), .dout(n6204));
  jand g05953(.dina(n6204), .dinb(n6201), .dout(n6205));
  jor  g05954(.dina(n6205), .dinb(n6200), .dout(n6206));
  jand g05955(.dina(n6206), .dinb(asqrt[38] ), .dout(n6207));
  jnot g05956(.din(n5846), .dout(n6208));
  jand g05957(.dina(n6208), .dinb(n5844), .dout(n6209));
  jand g05958(.dina(n6209), .dinb(asqrt[30] ), .dout(n6210));
  jxor g05959(.dina(n6210), .dinb(n5855), .dout(n6211));
  jnot g05960(.din(n6211), .dout(n6212));
  jor  g05961(.dina(n6200), .dinb(asqrt[38] ), .dout(n6213));
  jor  g05962(.dina(n6213), .dinb(n6205), .dout(n6214));
  jand g05963(.dina(n6214), .dinb(n6212), .dout(n6215));
  jor  g05964(.dina(n6215), .dinb(n6207), .dout(n6216));
  jand g05965(.dina(n6216), .dinb(asqrt[39] ), .dout(n6217));
  jor  g05966(.dina(n6216), .dinb(asqrt[39] ), .dout(n6218));
  jxor g05967(.dina(n5857), .dinb(n3907), .dout(n6219));
  jand g05968(.dina(n6219), .dinb(asqrt[30] ), .dout(n6220));
  jxor g05969(.dina(n6220), .dinb(n5863), .dout(n6221));
  jand g05970(.dina(n6221), .dinb(n6218), .dout(n6222));
  jor  g05971(.dina(n6222), .dinb(n6217), .dout(n6223));
  jand g05972(.dina(n6223), .dinb(asqrt[40] ), .dout(n6224));
  jor  g05973(.dina(n6217), .dinb(asqrt[40] ), .dout(n6225));
  jor  g05974(.dina(n6225), .dinb(n6222), .dout(n6226));
  jnot g05975(.din(n5871), .dout(n6227));
  jnot g05976(.din(n5873), .dout(n6228));
  jand g05977(.dina(asqrt[30] ), .dinb(n5867), .dout(n6229));
  jand g05978(.dina(n6229), .dinb(n6228), .dout(n6230));
  jor  g05979(.dina(n6230), .dinb(n6227), .dout(n6231));
  jnot g05980(.din(n5874), .dout(n6232));
  jand g05981(.dina(n6229), .dinb(n6232), .dout(n6233));
  jnot g05982(.din(n6233), .dout(n6234));
  jand g05983(.dina(n6234), .dinb(n6231), .dout(n6235));
  jand g05984(.dina(n6235), .dinb(n6226), .dout(n6236));
  jor  g05985(.dina(n6236), .dinb(n6224), .dout(n6237));
  jand g05986(.dina(n6237), .dinb(asqrt[41] ), .dout(n6238));
  jxor g05987(.dina(n5875), .dinb(n3371), .dout(n6239));
  jand g05988(.dina(n6239), .dinb(asqrt[30] ), .dout(n6240));
  jxor g05989(.dina(n6240), .dinb(n5882), .dout(n6241));
  jnot g05990(.din(n6241), .dout(n6242));
  jor  g05991(.dina(n6237), .dinb(asqrt[41] ), .dout(n6243));
  jand g05992(.dina(n6243), .dinb(n6242), .dout(n6244));
  jor  g05993(.dina(n6244), .dinb(n6238), .dout(n6245));
  jand g05994(.dina(n6245), .dinb(asqrt[42] ), .dout(n6246));
  jnot g05995(.din(n5887), .dout(n6247));
  jand g05996(.dina(n6247), .dinb(n5885), .dout(n6248));
  jand g05997(.dina(n6248), .dinb(asqrt[30] ), .dout(n6249));
  jxor g05998(.dina(n6249), .dinb(n5895), .dout(n6250));
  jnot g05999(.din(n6250), .dout(n6251));
  jor  g06000(.dina(n6238), .dinb(asqrt[42] ), .dout(n6252));
  jor  g06001(.dina(n6252), .dinb(n6244), .dout(n6253));
  jand g06002(.dina(n6253), .dinb(n6251), .dout(n6254));
  jor  g06003(.dina(n6254), .dinb(n6246), .dout(n6255));
  jand g06004(.dina(n6255), .dinb(asqrt[43] ), .dout(n6256));
  jor  g06005(.dina(n6255), .dinb(asqrt[43] ), .dout(n6257));
  jnot g06006(.din(n5901), .dout(n6258));
  jnot g06007(.din(n5902), .dout(n6259));
  jand g06008(.dina(asqrt[30] ), .dinb(n5898), .dout(n6260));
  jand g06009(.dina(n6260), .dinb(n6259), .dout(n6261));
  jor  g06010(.dina(n6261), .dinb(n6258), .dout(n6262));
  jnot g06011(.din(n5903), .dout(n6263));
  jand g06012(.dina(n6260), .dinb(n6263), .dout(n6264));
  jnot g06013(.din(n6264), .dout(n6265));
  jand g06014(.dina(n6265), .dinb(n6262), .dout(n6266));
  jand g06015(.dina(n6266), .dinb(n6257), .dout(n6267));
  jor  g06016(.dina(n6267), .dinb(n6256), .dout(n6268));
  jand g06017(.dina(n6268), .dinb(asqrt[44] ), .dout(n6269));
  jor  g06018(.dina(n6256), .dinb(asqrt[44] ), .dout(n6270));
  jor  g06019(.dina(n6270), .dinb(n6267), .dout(n6271));
  jnot g06020(.din(n5909), .dout(n6272));
  jnot g06021(.din(n5911), .dout(n6273));
  jand g06022(.dina(asqrt[30] ), .dinb(n5905), .dout(n6274));
  jand g06023(.dina(n6274), .dinb(n6273), .dout(n6275));
  jor  g06024(.dina(n6275), .dinb(n6272), .dout(n6276));
  jnot g06025(.din(n5912), .dout(n6277));
  jand g06026(.dina(n6274), .dinb(n6277), .dout(n6278));
  jnot g06027(.din(n6278), .dout(n6279));
  jand g06028(.dina(n6279), .dinb(n6276), .dout(n6280));
  jand g06029(.dina(n6280), .dinb(n6271), .dout(n6281));
  jor  g06030(.dina(n6281), .dinb(n6269), .dout(n6282));
  jand g06031(.dina(n6282), .dinb(asqrt[45] ), .dout(n6283));
  jxor g06032(.dina(n5913), .dinb(n2420), .dout(n6284));
  jand g06033(.dina(n6284), .dinb(asqrt[30] ), .dout(n6285));
  jxor g06034(.dina(n6285), .dinb(n5923), .dout(n6286));
  jnot g06035(.din(n6286), .dout(n6287));
  jor  g06036(.dina(n6282), .dinb(asqrt[45] ), .dout(n6288));
  jand g06037(.dina(n6288), .dinb(n6287), .dout(n6289));
  jor  g06038(.dina(n6289), .dinb(n6283), .dout(n6290));
  jand g06039(.dina(n6290), .dinb(asqrt[46] ), .dout(n6291));
  jnot g06040(.din(n5928), .dout(n6292));
  jand g06041(.dina(n6292), .dinb(n5926), .dout(n6293));
  jand g06042(.dina(n6293), .dinb(asqrt[30] ), .dout(n6294));
  jxor g06043(.dina(n6294), .dinb(n5936), .dout(n6295));
  jnot g06044(.din(n6295), .dout(n6296));
  jor  g06045(.dina(n6283), .dinb(asqrt[46] ), .dout(n6297));
  jor  g06046(.dina(n6297), .dinb(n6289), .dout(n6298));
  jand g06047(.dina(n6298), .dinb(n6296), .dout(n6299));
  jor  g06048(.dina(n6299), .dinb(n6291), .dout(n6300));
  jand g06049(.dina(n6300), .dinb(asqrt[47] ), .dout(n6301));
  jor  g06050(.dina(n6300), .dinb(asqrt[47] ), .dout(n6302));
  jnot g06051(.din(n5942), .dout(n6303));
  jnot g06052(.din(n5943), .dout(n6304));
  jand g06053(.dina(asqrt[30] ), .dinb(n5939), .dout(n6305));
  jand g06054(.dina(n6305), .dinb(n6304), .dout(n6306));
  jor  g06055(.dina(n6306), .dinb(n6303), .dout(n6307));
  jnot g06056(.din(n5944), .dout(n6308));
  jand g06057(.dina(n6305), .dinb(n6308), .dout(n6309));
  jnot g06058(.din(n6309), .dout(n6310));
  jand g06059(.dina(n6310), .dinb(n6307), .dout(n6311));
  jand g06060(.dina(n6311), .dinb(n6302), .dout(n6312));
  jor  g06061(.dina(n6312), .dinb(n6301), .dout(n6313));
  jand g06062(.dina(n6313), .dinb(asqrt[48] ), .dout(n6314));
  jor  g06063(.dina(n6301), .dinb(asqrt[48] ), .dout(n6315));
  jor  g06064(.dina(n6315), .dinb(n6312), .dout(n6316));
  jnot g06065(.din(n5950), .dout(n6317));
  jnot g06066(.din(n5952), .dout(n6318));
  jand g06067(.dina(asqrt[30] ), .dinb(n5946), .dout(n6319));
  jand g06068(.dina(n6319), .dinb(n6318), .dout(n6320));
  jor  g06069(.dina(n6320), .dinb(n6317), .dout(n6321));
  jnot g06070(.din(n5953), .dout(n6322));
  jand g06071(.dina(n6319), .dinb(n6322), .dout(n6323));
  jnot g06072(.din(n6323), .dout(n6324));
  jand g06073(.dina(n6324), .dinb(n6321), .dout(n6325));
  jand g06074(.dina(n6325), .dinb(n6316), .dout(n6326));
  jor  g06075(.dina(n6326), .dinb(n6314), .dout(n6327));
  jand g06076(.dina(n6327), .dinb(asqrt[49] ), .dout(n6328));
  jxor g06077(.dina(n5954), .dinb(n1641), .dout(n6329));
  jand g06078(.dina(n6329), .dinb(asqrt[30] ), .dout(n6330));
  jxor g06079(.dina(n6330), .dinb(n5964), .dout(n6331));
  jnot g06080(.din(n6331), .dout(n6332));
  jor  g06081(.dina(n6327), .dinb(asqrt[49] ), .dout(n6333));
  jand g06082(.dina(n6333), .dinb(n6332), .dout(n6334));
  jor  g06083(.dina(n6334), .dinb(n6328), .dout(n6335));
  jand g06084(.dina(n6335), .dinb(asqrt[50] ), .dout(n6336));
  jnot g06085(.din(n5969), .dout(n6337));
  jand g06086(.dina(n6337), .dinb(n5967), .dout(n6338));
  jand g06087(.dina(n6338), .dinb(asqrt[30] ), .dout(n6339));
  jxor g06088(.dina(n6339), .dinb(n5977), .dout(n6340));
  jnot g06089(.din(n6340), .dout(n6341));
  jor  g06090(.dina(n6328), .dinb(asqrt[50] ), .dout(n6342));
  jor  g06091(.dina(n6342), .dinb(n6334), .dout(n6343));
  jand g06092(.dina(n6343), .dinb(n6341), .dout(n6344));
  jor  g06093(.dina(n6344), .dinb(n6336), .dout(n6345));
  jand g06094(.dina(n6345), .dinb(asqrt[51] ), .dout(n6346));
  jor  g06095(.dina(n6345), .dinb(asqrt[51] ), .dout(n6347));
  jnot g06096(.din(n5983), .dout(n6348));
  jnot g06097(.din(n5984), .dout(n6349));
  jand g06098(.dina(asqrt[30] ), .dinb(n5980), .dout(n6350));
  jand g06099(.dina(n6350), .dinb(n6349), .dout(n6351));
  jor  g06100(.dina(n6351), .dinb(n6348), .dout(n6352));
  jnot g06101(.din(n5985), .dout(n6353));
  jand g06102(.dina(n6350), .dinb(n6353), .dout(n6354));
  jnot g06103(.din(n6354), .dout(n6355));
  jand g06104(.dina(n6355), .dinb(n6352), .dout(n6356));
  jand g06105(.dina(n6356), .dinb(n6347), .dout(n6357));
  jor  g06106(.dina(n6357), .dinb(n6346), .dout(n6358));
  jand g06107(.dina(n6358), .dinb(asqrt[52] ), .dout(n6359));
  jor  g06108(.dina(n6346), .dinb(asqrt[52] ), .dout(n6360));
  jor  g06109(.dina(n6360), .dinb(n6357), .dout(n6361));
  jnot g06110(.din(n5991), .dout(n6362));
  jnot g06111(.din(n5993), .dout(n6363));
  jand g06112(.dina(asqrt[30] ), .dinb(n5987), .dout(n6364));
  jand g06113(.dina(n6364), .dinb(n6363), .dout(n6365));
  jor  g06114(.dina(n6365), .dinb(n6362), .dout(n6366));
  jnot g06115(.din(n5994), .dout(n6367));
  jand g06116(.dina(n6364), .dinb(n6367), .dout(n6368));
  jnot g06117(.din(n6368), .dout(n6369));
  jand g06118(.dina(n6369), .dinb(n6366), .dout(n6370));
  jand g06119(.dina(n6370), .dinb(n6361), .dout(n6371));
  jor  g06120(.dina(n6371), .dinb(n6359), .dout(n6372));
  jand g06121(.dina(n6372), .dinb(asqrt[53] ), .dout(n6373));
  jxor g06122(.dina(n5995), .dinb(n1034), .dout(n6374));
  jand g06123(.dina(n6374), .dinb(asqrt[30] ), .dout(n6375));
  jxor g06124(.dina(n6375), .dinb(n6005), .dout(n6376));
  jnot g06125(.din(n6376), .dout(n6377));
  jor  g06126(.dina(n6372), .dinb(asqrt[53] ), .dout(n6378));
  jand g06127(.dina(n6378), .dinb(n6377), .dout(n6379));
  jor  g06128(.dina(n6379), .dinb(n6373), .dout(n6380));
  jand g06129(.dina(n6380), .dinb(asqrt[54] ), .dout(n6381));
  jnot g06130(.din(n6010), .dout(n6382));
  jand g06131(.dina(n6382), .dinb(n6008), .dout(n6383));
  jand g06132(.dina(n6383), .dinb(asqrt[30] ), .dout(n6384));
  jxor g06133(.dina(n6384), .dinb(n6018), .dout(n6385));
  jnot g06134(.din(n6385), .dout(n6386));
  jor  g06135(.dina(n6373), .dinb(asqrt[54] ), .dout(n6387));
  jor  g06136(.dina(n6387), .dinb(n6379), .dout(n6388));
  jand g06137(.dina(n6388), .dinb(n6386), .dout(n6389));
  jor  g06138(.dina(n6389), .dinb(n6381), .dout(n6390));
  jand g06139(.dina(n6390), .dinb(asqrt[55] ), .dout(n6391));
  jor  g06140(.dina(n6390), .dinb(asqrt[55] ), .dout(n6392));
  jnot g06141(.din(n6024), .dout(n6393));
  jnot g06142(.din(n6025), .dout(n6394));
  jand g06143(.dina(asqrt[30] ), .dinb(n6021), .dout(n6395));
  jand g06144(.dina(n6395), .dinb(n6394), .dout(n6396));
  jor  g06145(.dina(n6396), .dinb(n6393), .dout(n6397));
  jnot g06146(.din(n6026), .dout(n6398));
  jand g06147(.dina(n6395), .dinb(n6398), .dout(n6399));
  jnot g06148(.din(n6399), .dout(n6400));
  jand g06149(.dina(n6400), .dinb(n6397), .dout(n6401));
  jand g06150(.dina(n6401), .dinb(n6392), .dout(n6402));
  jor  g06151(.dina(n6402), .dinb(n6391), .dout(n6403));
  jand g06152(.dina(n6403), .dinb(asqrt[56] ), .dout(n6404));
  jor  g06153(.dina(n6391), .dinb(asqrt[56] ), .dout(n6405));
  jor  g06154(.dina(n6405), .dinb(n6402), .dout(n6406));
  jnot g06155(.din(n6032), .dout(n6407));
  jnot g06156(.din(n6034), .dout(n6408));
  jand g06157(.dina(asqrt[30] ), .dinb(n6028), .dout(n6409));
  jand g06158(.dina(n6409), .dinb(n6408), .dout(n6410));
  jor  g06159(.dina(n6410), .dinb(n6407), .dout(n6411));
  jnot g06160(.din(n6035), .dout(n6412));
  jand g06161(.dina(n6409), .dinb(n6412), .dout(n6413));
  jnot g06162(.din(n6413), .dout(n6414));
  jand g06163(.dina(n6414), .dinb(n6411), .dout(n6415));
  jand g06164(.dina(n6415), .dinb(n6406), .dout(n6416));
  jor  g06165(.dina(n6416), .dinb(n6404), .dout(n6417));
  jand g06166(.dina(n6417), .dinb(asqrt[57] ), .dout(n6418));
  jxor g06167(.dina(n6036), .dinb(n590), .dout(n6419));
  jand g06168(.dina(n6419), .dinb(asqrt[30] ), .dout(n6420));
  jxor g06169(.dina(n6420), .dinb(n6046), .dout(n6421));
  jnot g06170(.din(n6421), .dout(n6422));
  jor  g06171(.dina(n6417), .dinb(asqrt[57] ), .dout(n6423));
  jand g06172(.dina(n6423), .dinb(n6422), .dout(n6424));
  jor  g06173(.dina(n6424), .dinb(n6418), .dout(n6425));
  jand g06174(.dina(n6425), .dinb(asqrt[58] ), .dout(n6426));
  jnot g06175(.din(n6051), .dout(n6427));
  jand g06176(.dina(n6427), .dinb(n6049), .dout(n6428));
  jand g06177(.dina(n6428), .dinb(asqrt[30] ), .dout(n6429));
  jxor g06178(.dina(n6429), .dinb(n6059), .dout(n6430));
  jnot g06179(.din(n6430), .dout(n6431));
  jor  g06180(.dina(n6418), .dinb(asqrt[58] ), .dout(n6432));
  jor  g06181(.dina(n6432), .dinb(n6424), .dout(n6433));
  jand g06182(.dina(n6433), .dinb(n6431), .dout(n6434));
  jor  g06183(.dina(n6434), .dinb(n6426), .dout(n6435));
  jand g06184(.dina(n6435), .dinb(asqrt[59] ), .dout(n6436));
  jor  g06185(.dina(n6435), .dinb(asqrt[59] ), .dout(n6437));
  jnot g06186(.din(n6065), .dout(n6438));
  jnot g06187(.din(n6066), .dout(n6439));
  jand g06188(.dina(asqrt[30] ), .dinb(n6062), .dout(n6440));
  jand g06189(.dina(n6440), .dinb(n6439), .dout(n6441));
  jor  g06190(.dina(n6441), .dinb(n6438), .dout(n6442));
  jnot g06191(.din(n6067), .dout(n6443));
  jand g06192(.dina(n6440), .dinb(n6443), .dout(n6444));
  jnot g06193(.din(n6444), .dout(n6445));
  jand g06194(.dina(n6445), .dinb(n6442), .dout(n6446));
  jand g06195(.dina(n6446), .dinb(n6437), .dout(n6447));
  jor  g06196(.dina(n6447), .dinb(n6436), .dout(n6448));
  jand g06197(.dina(n6448), .dinb(asqrt[60] ), .dout(n6449));
  jor  g06198(.dina(n6436), .dinb(asqrt[60] ), .dout(n6450));
  jor  g06199(.dina(n6450), .dinb(n6447), .dout(n6451));
  jnot g06200(.din(n6073), .dout(n6452));
  jnot g06201(.din(n6075), .dout(n6453));
  jand g06202(.dina(asqrt[30] ), .dinb(n6069), .dout(n6454));
  jand g06203(.dina(n6454), .dinb(n6453), .dout(n6455));
  jor  g06204(.dina(n6455), .dinb(n6452), .dout(n6456));
  jnot g06205(.din(n6076), .dout(n6457));
  jand g06206(.dina(n6454), .dinb(n6457), .dout(n6458));
  jnot g06207(.din(n6458), .dout(n6459));
  jand g06208(.dina(n6459), .dinb(n6456), .dout(n6460));
  jand g06209(.dina(n6460), .dinb(n6451), .dout(n6461));
  jor  g06210(.dina(n6461), .dinb(n6449), .dout(n6462));
  jand g06211(.dina(n6462), .dinb(asqrt[61] ), .dout(n6463));
  jxor g06212(.dina(n6077), .dinb(n290), .dout(n6464));
  jand g06213(.dina(n6464), .dinb(asqrt[30] ), .dout(n6465));
  jxor g06214(.dina(n6465), .dinb(n6087), .dout(n6466));
  jnot g06215(.din(n6466), .dout(n6467));
  jor  g06216(.dina(n6462), .dinb(asqrt[61] ), .dout(n6468));
  jand g06217(.dina(n6468), .dinb(n6467), .dout(n6469));
  jor  g06218(.dina(n6469), .dinb(n6463), .dout(n6470));
  jand g06219(.dina(n6470), .dinb(asqrt[62] ), .dout(n6471));
  jnot g06220(.din(n6092), .dout(n6472));
  jand g06221(.dina(n6472), .dinb(n6090), .dout(n6473));
  jand g06222(.dina(n6473), .dinb(asqrt[30] ), .dout(n6474));
  jxor g06223(.dina(n6474), .dinb(n6100), .dout(n6475));
  jnot g06224(.din(n6475), .dout(n6476));
  jor  g06225(.dina(n6463), .dinb(asqrt[62] ), .dout(n6477));
  jor  g06226(.dina(n6477), .dinb(n6469), .dout(n6478));
  jand g06227(.dina(n6478), .dinb(n6476), .dout(n6479));
  jor  g06228(.dina(n6479), .dinb(n6471), .dout(n6480));
  jxor g06229(.dina(n6102), .dinb(n199), .dout(n6481));
  jand g06230(.dina(n6481), .dinb(asqrt[30] ), .dout(n6482));
  jxor g06231(.dina(n6482), .dinb(n6107), .dout(n6483));
  jnot g06232(.din(n6109), .dout(n6484));
  jnot g06233(.din(n6113), .dout(n6485));
  jand g06234(.dina(asqrt[30] ), .dinb(n6485), .dout(n6486));
  jand g06235(.dina(n6486), .dinb(n6484), .dout(n6487));
  jor  g06236(.dina(n6487), .dinb(n6120), .dout(n6488));
  jor  g06237(.dina(n6488), .dinb(n6483), .dout(n6489));
  jnot g06238(.din(n6489), .dout(n6490));
  jand g06239(.dina(n6490), .dinb(n6480), .dout(n6491));
  jor  g06240(.dina(n6491), .dinb(asqrt[63] ), .dout(n6492));
  jnot g06241(.din(n6483), .dout(n6493));
  jor  g06242(.dina(n6493), .dinb(n6480), .dout(n6494));
  jor  g06243(.dina(n6486), .dinb(n6484), .dout(n6495));
  jand g06244(.dina(n6485), .dinb(n6484), .dout(n6496));
  jor  g06245(.dina(n6496), .dinb(n194), .dout(n6497));
  jnot g06246(.din(n6497), .dout(n6498));
  jand g06247(.dina(n6498), .dinb(n6495), .dout(n6499));
  jnot g06248(.din(asqrt[30] ), .dout(n6500));
  jnot g06249(.din(n6499), .dout(n6503));
  jand g06250(.dina(n6503), .dinb(n6494), .dout(n6504));
  jand g06251(.dina(n6504), .dinb(n6492), .dout(n6505));
  jxor g06252(.dina(n6158), .dinb(n5121), .dout(n6506));
  jor  g06253(.dina(n6506), .dinb(n6505), .dout(n6507));
  jxor g06254(.dina(n6507), .dinb(n6132), .dout(n6508));
  jor  g06255(.dina(n6505), .dinb(n6134), .dout(n6509));
  jnot g06256(.din(a[56] ), .dout(n6510));
  jnot g06257(.din(a[57] ), .dout(n6511));
  jand g06258(.dina(n6134), .dinb(n6511), .dout(n6512));
  jand g06259(.dina(n6512), .dinb(n6510), .dout(n6513));
  jnot g06260(.din(n6513), .dout(n6514));
  jand g06261(.dina(n6514), .dinb(n6509), .dout(n6515));
  jor  g06262(.dina(n6515), .dinb(n6500), .dout(n6516));
  jor  g06263(.dina(n6505), .dinb(a[58] ), .dout(n6517));
  jxor g06264(.dina(n6517), .dinb(n6135), .dout(n6518));
  jand g06265(.dina(n6515), .dinb(n6500), .dout(n6519));
  jor  g06266(.dina(n6519), .dinb(n6518), .dout(n6520));
  jand g06267(.dina(n6520), .dinb(n6516), .dout(n6521));
  jor  g06268(.dina(n6521), .dinb(n5793), .dout(n6522));
  jand g06269(.dina(n6516), .dinb(n5793), .dout(n6523));
  jand g06270(.dina(n6523), .dinb(n6520), .dout(n6524));
  jor  g06271(.dina(n6517), .dinb(a[59] ), .dout(n6525));
  jnot g06272(.din(n6492), .dout(n6526));
  jnot g06273(.din(n6494), .dout(n6527));
  jor  g06274(.dina(n6499), .dinb(n6500), .dout(n6528));
  jor  g06275(.dina(n6528), .dinb(n6527), .dout(n6529));
  jor  g06276(.dina(n6529), .dinb(n6526), .dout(n6530));
  jand g06277(.dina(n6530), .dinb(n6525), .dout(n6531));
  jxor g06278(.dina(n6531), .dinb(n5797), .dout(n6532));
  jor  g06279(.dina(n6532), .dinb(n6524), .dout(n6533));
  jand g06280(.dina(n6533), .dinb(n6522), .dout(n6534));
  jor  g06281(.dina(n6534), .dinb(n5788), .dout(n6535));
  jand g06282(.dina(n6534), .dinb(n5788), .dout(n6536));
  jxor g06283(.dina(n6138), .dinb(n5793), .dout(n6537));
  jor  g06284(.dina(n6537), .dinb(n6505), .dout(n6538));
  jxor g06285(.dina(n6538), .dinb(n6141), .dout(n6539));
  jor  g06286(.dina(n6539), .dinb(n6536), .dout(n6540));
  jand g06287(.dina(n6540), .dinb(n6535), .dout(n6541));
  jor  g06288(.dina(n6541), .dinb(n5121), .dout(n6542));
  jand g06289(.dina(n6535), .dinb(n5121), .dout(n6543));
  jand g06290(.dina(n6543), .dinb(n6540), .dout(n6544));
  jnot g06291(.din(n6145), .dout(n6545));
  jnot g06292(.din(n6505), .dout(asqrt[29] ));
  jand g06293(.dina(asqrt[29] ), .dinb(n6545), .dout(n6547));
  jand g06294(.dina(n6547), .dinb(n6156), .dout(n6548));
  jor  g06295(.dina(n6548), .dinb(n6154), .dout(n6549));
  jand g06296(.dina(n6547), .dinb(n6157), .dout(n6550));
  jnot g06297(.din(n6550), .dout(n6551));
  jand g06298(.dina(n6551), .dinb(n6549), .dout(n6552));
  jnot g06299(.din(n6552), .dout(n6553));
  jor  g06300(.dina(n6553), .dinb(n6544), .dout(n6554));
  jand g06301(.dina(n6554), .dinb(n6542), .dout(n6555));
  jor  g06302(.dina(n6555), .dinb(n5116), .dout(n6556));
  jnot g06303(.din(n6508), .dout(n6557));
  jand g06304(.dina(n6555), .dinb(n5116), .dout(n6558));
  jor  g06305(.dina(n6558), .dinb(n6557), .dout(n6559));
  jand g06306(.dina(n6559), .dinb(n6556), .dout(n6560));
  jor  g06307(.dina(n6560), .dinb(n4499), .dout(n6561));
  jnot g06308(.din(n6166), .dout(n6562));
  jor  g06309(.dina(n6562), .dinb(n6164), .dout(n6563));
  jor  g06310(.dina(n6563), .dinb(n6505), .dout(n6564));
  jxor g06311(.dina(n6564), .dinb(n6175), .dout(n6565));
  jand g06312(.dina(n6556), .dinb(n4499), .dout(n6566));
  jand g06313(.dina(n6566), .dinb(n6559), .dout(n6567));
  jor  g06314(.dina(n6567), .dinb(n6565), .dout(n6568));
  jand g06315(.dina(n6568), .dinb(n6561), .dout(n6569));
  jor  g06316(.dina(n6569), .dinb(n4494), .dout(n6570));
  jand g06317(.dina(n6569), .dinb(n4494), .dout(n6571));
  jnot g06318(.din(n6183), .dout(n6572));
  jxor g06319(.dina(n6177), .dinb(n4499), .dout(n6573));
  jor  g06320(.dina(n6573), .dinb(n6505), .dout(n6574));
  jxor g06321(.dina(n6574), .dinb(n6572), .dout(n6575));
  jnot g06322(.din(n6575), .dout(n6576));
  jor  g06323(.dina(n6576), .dinb(n6571), .dout(n6577));
  jand g06324(.dina(n6577), .dinb(n6570), .dout(n6578));
  jor  g06325(.dina(n6578), .dinb(n3912), .dout(n6579));
  jnot g06326(.din(n6188), .dout(n6580));
  jor  g06327(.dina(n6580), .dinb(n6186), .dout(n6581));
  jor  g06328(.dina(n6581), .dinb(n6505), .dout(n6582));
  jxor g06329(.dina(n6582), .dinb(n6197), .dout(n6583));
  jand g06330(.dina(n6570), .dinb(n3912), .dout(n6584));
  jand g06331(.dina(n6584), .dinb(n6577), .dout(n6585));
  jor  g06332(.dina(n6585), .dinb(n6583), .dout(n6586));
  jand g06333(.dina(n6586), .dinb(n6579), .dout(n6587));
  jor  g06334(.dina(n6587), .dinb(n3907), .dout(n6588));
  jand g06335(.dina(n6587), .dinb(n3907), .dout(n6589));
  jnot g06336(.din(n6204), .dout(n6590));
  jxor g06337(.dina(n6199), .dinb(n3912), .dout(n6591));
  jor  g06338(.dina(n6591), .dinb(n6505), .dout(n6592));
  jxor g06339(.dina(n6592), .dinb(n6590), .dout(n6593));
  jnot g06340(.din(n6593), .dout(n6594));
  jor  g06341(.dina(n6594), .dinb(n6589), .dout(n6595));
  jand g06342(.dina(n6595), .dinb(n6588), .dout(n6596));
  jor  g06343(.dina(n6596), .dinb(n3376), .dout(n6597));
  jand g06344(.dina(n6588), .dinb(n3376), .dout(n6598));
  jand g06345(.dina(n6598), .dinb(n6595), .dout(n6599));
  jnot g06346(.din(n6207), .dout(n6600));
  jand g06347(.dina(asqrt[29] ), .dinb(n6600), .dout(n6601));
  jand g06348(.dina(n6601), .dinb(n6214), .dout(n6602));
  jor  g06349(.dina(n6602), .dinb(n6212), .dout(n6603));
  jand g06350(.dina(n6601), .dinb(n6215), .dout(n6604));
  jnot g06351(.din(n6604), .dout(n6605));
  jand g06352(.dina(n6605), .dinb(n6603), .dout(n6606));
  jnot g06353(.din(n6606), .dout(n6607));
  jor  g06354(.dina(n6607), .dinb(n6599), .dout(n6608));
  jand g06355(.dina(n6608), .dinb(n6597), .dout(n6609));
  jor  g06356(.dina(n6609), .dinb(n3371), .dout(n6610));
  jxor g06357(.dina(n6216), .dinb(n3376), .dout(n6611));
  jor  g06358(.dina(n6611), .dinb(n6505), .dout(n6612));
  jxor g06359(.dina(n6612), .dinb(n6221), .dout(n6613));
  jand g06360(.dina(n6609), .dinb(n3371), .dout(n6614));
  jor  g06361(.dina(n6614), .dinb(n6613), .dout(n6615));
  jand g06362(.dina(n6615), .dinb(n6610), .dout(n6616));
  jor  g06363(.dina(n6616), .dinb(n2875), .dout(n6617));
  jnot g06364(.din(n6226), .dout(n6618));
  jor  g06365(.dina(n6618), .dinb(n6224), .dout(n6619));
  jor  g06366(.dina(n6619), .dinb(n6505), .dout(n6620));
  jxor g06367(.dina(n6620), .dinb(n6235), .dout(n6621));
  jand g06368(.dina(n6610), .dinb(n2875), .dout(n6622));
  jand g06369(.dina(n6622), .dinb(n6615), .dout(n6623));
  jor  g06370(.dina(n6623), .dinb(n6621), .dout(n6624));
  jand g06371(.dina(n6624), .dinb(n6617), .dout(n6625));
  jor  g06372(.dina(n6625), .dinb(n2870), .dout(n6626));
  jand g06373(.dina(n6625), .dinb(n2870), .dout(n6627));
  jnot g06374(.din(n6238), .dout(n6628));
  jand g06375(.dina(asqrt[29] ), .dinb(n6628), .dout(n6629));
  jand g06376(.dina(n6629), .dinb(n6243), .dout(n6630));
  jor  g06377(.dina(n6630), .dinb(n6242), .dout(n6631));
  jand g06378(.dina(n6629), .dinb(n6244), .dout(n6632));
  jnot g06379(.din(n6632), .dout(n6633));
  jand g06380(.dina(n6633), .dinb(n6631), .dout(n6634));
  jnot g06381(.din(n6634), .dout(n6635));
  jor  g06382(.dina(n6635), .dinb(n6627), .dout(n6636));
  jand g06383(.dina(n6636), .dinb(n6626), .dout(n6637));
  jor  g06384(.dina(n6637), .dinb(n2425), .dout(n6638));
  jand g06385(.dina(n6626), .dinb(n2425), .dout(n6639));
  jand g06386(.dina(n6639), .dinb(n6636), .dout(n6640));
  jnot g06387(.din(n6246), .dout(n6641));
  jand g06388(.dina(asqrt[29] ), .dinb(n6641), .dout(n6642));
  jand g06389(.dina(n6642), .dinb(n6253), .dout(n6643));
  jor  g06390(.dina(n6643), .dinb(n6251), .dout(n6644));
  jand g06391(.dina(n6642), .dinb(n6254), .dout(n6645));
  jnot g06392(.din(n6645), .dout(n6646));
  jand g06393(.dina(n6646), .dinb(n6644), .dout(n6647));
  jnot g06394(.din(n6647), .dout(n6648));
  jor  g06395(.dina(n6648), .dinb(n6640), .dout(n6649));
  jand g06396(.dina(n6649), .dinb(n6638), .dout(n6650));
  jor  g06397(.dina(n6650), .dinb(n2420), .dout(n6651));
  jxor g06398(.dina(n6255), .dinb(n2425), .dout(n6652));
  jor  g06399(.dina(n6652), .dinb(n6505), .dout(n6653));
  jxor g06400(.dina(n6653), .dinb(n6266), .dout(n6654));
  jand g06401(.dina(n6650), .dinb(n2420), .dout(n6655));
  jor  g06402(.dina(n6655), .dinb(n6654), .dout(n6656));
  jand g06403(.dina(n6656), .dinb(n6651), .dout(n6657));
  jor  g06404(.dina(n6657), .dinb(n2010), .dout(n6658));
  jnot g06405(.din(n6271), .dout(n6659));
  jor  g06406(.dina(n6659), .dinb(n6269), .dout(n6660));
  jor  g06407(.dina(n6660), .dinb(n6505), .dout(n6661));
  jxor g06408(.dina(n6661), .dinb(n6280), .dout(n6662));
  jand g06409(.dina(n6651), .dinb(n2010), .dout(n6663));
  jand g06410(.dina(n6663), .dinb(n6656), .dout(n6664));
  jor  g06411(.dina(n6664), .dinb(n6662), .dout(n6665));
  jand g06412(.dina(n6665), .dinb(n6658), .dout(n6666));
  jor  g06413(.dina(n6666), .dinb(n2005), .dout(n6667));
  jand g06414(.dina(n6666), .dinb(n2005), .dout(n6668));
  jnot g06415(.din(n6283), .dout(n6669));
  jand g06416(.dina(asqrt[29] ), .dinb(n6669), .dout(n6670));
  jand g06417(.dina(n6670), .dinb(n6288), .dout(n6671));
  jor  g06418(.dina(n6671), .dinb(n6287), .dout(n6672));
  jand g06419(.dina(n6670), .dinb(n6289), .dout(n6673));
  jnot g06420(.din(n6673), .dout(n6674));
  jand g06421(.dina(n6674), .dinb(n6672), .dout(n6675));
  jnot g06422(.din(n6675), .dout(n6676));
  jor  g06423(.dina(n6676), .dinb(n6668), .dout(n6677));
  jand g06424(.dina(n6677), .dinb(n6667), .dout(n6678));
  jor  g06425(.dina(n6678), .dinb(n1646), .dout(n6679));
  jand g06426(.dina(n6667), .dinb(n1646), .dout(n6680));
  jand g06427(.dina(n6680), .dinb(n6677), .dout(n6681));
  jnot g06428(.din(n6291), .dout(n6682));
  jand g06429(.dina(asqrt[29] ), .dinb(n6682), .dout(n6683));
  jand g06430(.dina(n6683), .dinb(n6298), .dout(n6684));
  jor  g06431(.dina(n6684), .dinb(n6296), .dout(n6685));
  jand g06432(.dina(n6683), .dinb(n6299), .dout(n6686));
  jnot g06433(.din(n6686), .dout(n6687));
  jand g06434(.dina(n6687), .dinb(n6685), .dout(n6688));
  jnot g06435(.din(n6688), .dout(n6689));
  jor  g06436(.dina(n6689), .dinb(n6681), .dout(n6690));
  jand g06437(.dina(n6690), .dinb(n6679), .dout(n6691));
  jor  g06438(.dina(n6691), .dinb(n1641), .dout(n6692));
  jxor g06439(.dina(n6300), .dinb(n1646), .dout(n6693));
  jor  g06440(.dina(n6693), .dinb(n6505), .dout(n6694));
  jxor g06441(.dina(n6694), .dinb(n6311), .dout(n6695));
  jand g06442(.dina(n6691), .dinb(n1641), .dout(n6696));
  jor  g06443(.dina(n6696), .dinb(n6695), .dout(n6697));
  jand g06444(.dina(n6697), .dinb(n6692), .dout(n6698));
  jor  g06445(.dina(n6698), .dinb(n1317), .dout(n6699));
  jnot g06446(.din(n6316), .dout(n6700));
  jor  g06447(.dina(n6700), .dinb(n6314), .dout(n6701));
  jor  g06448(.dina(n6701), .dinb(n6505), .dout(n6702));
  jxor g06449(.dina(n6702), .dinb(n6325), .dout(n6703));
  jand g06450(.dina(n6692), .dinb(n1317), .dout(n6704));
  jand g06451(.dina(n6704), .dinb(n6697), .dout(n6705));
  jor  g06452(.dina(n6705), .dinb(n6703), .dout(n6706));
  jand g06453(.dina(n6706), .dinb(n6699), .dout(n6707));
  jor  g06454(.dina(n6707), .dinb(n1312), .dout(n6708));
  jand g06455(.dina(n6707), .dinb(n1312), .dout(n6709));
  jnot g06456(.din(n6328), .dout(n6710));
  jand g06457(.dina(asqrt[29] ), .dinb(n6710), .dout(n6711));
  jand g06458(.dina(n6711), .dinb(n6333), .dout(n6712));
  jor  g06459(.dina(n6712), .dinb(n6332), .dout(n6713));
  jand g06460(.dina(n6711), .dinb(n6334), .dout(n6714));
  jnot g06461(.din(n6714), .dout(n6715));
  jand g06462(.dina(n6715), .dinb(n6713), .dout(n6716));
  jnot g06463(.din(n6716), .dout(n6717));
  jor  g06464(.dina(n6717), .dinb(n6709), .dout(n6718));
  jand g06465(.dina(n6718), .dinb(n6708), .dout(n6719));
  jor  g06466(.dina(n6719), .dinb(n1039), .dout(n6720));
  jand g06467(.dina(n6708), .dinb(n1039), .dout(n6721));
  jand g06468(.dina(n6721), .dinb(n6718), .dout(n6722));
  jnot g06469(.din(n6336), .dout(n6723));
  jand g06470(.dina(asqrt[29] ), .dinb(n6723), .dout(n6724));
  jand g06471(.dina(n6724), .dinb(n6343), .dout(n6725));
  jor  g06472(.dina(n6725), .dinb(n6341), .dout(n6726));
  jand g06473(.dina(n6724), .dinb(n6344), .dout(n6727));
  jnot g06474(.din(n6727), .dout(n6728));
  jand g06475(.dina(n6728), .dinb(n6726), .dout(n6729));
  jnot g06476(.din(n6729), .dout(n6730));
  jor  g06477(.dina(n6730), .dinb(n6722), .dout(n6731));
  jand g06478(.dina(n6731), .dinb(n6720), .dout(n6732));
  jor  g06479(.dina(n6732), .dinb(n1034), .dout(n6733));
  jxor g06480(.dina(n6345), .dinb(n1039), .dout(n6734));
  jor  g06481(.dina(n6734), .dinb(n6505), .dout(n6735));
  jxor g06482(.dina(n6735), .dinb(n6356), .dout(n6736));
  jand g06483(.dina(n6732), .dinb(n1034), .dout(n6737));
  jor  g06484(.dina(n6737), .dinb(n6736), .dout(n6738));
  jand g06485(.dina(n6738), .dinb(n6733), .dout(n6739));
  jor  g06486(.dina(n6739), .dinb(n796), .dout(n6740));
  jnot g06487(.din(n6361), .dout(n6741));
  jor  g06488(.dina(n6741), .dinb(n6359), .dout(n6742));
  jor  g06489(.dina(n6742), .dinb(n6505), .dout(n6743));
  jxor g06490(.dina(n6743), .dinb(n6370), .dout(n6744));
  jand g06491(.dina(n6733), .dinb(n796), .dout(n6745));
  jand g06492(.dina(n6745), .dinb(n6738), .dout(n6746));
  jor  g06493(.dina(n6746), .dinb(n6744), .dout(n6747));
  jand g06494(.dina(n6747), .dinb(n6740), .dout(n6748));
  jor  g06495(.dina(n6748), .dinb(n791), .dout(n6749));
  jand g06496(.dina(n6748), .dinb(n791), .dout(n6750));
  jnot g06497(.din(n6373), .dout(n6751));
  jand g06498(.dina(asqrt[29] ), .dinb(n6751), .dout(n6752));
  jand g06499(.dina(n6752), .dinb(n6378), .dout(n6753));
  jor  g06500(.dina(n6753), .dinb(n6377), .dout(n6754));
  jand g06501(.dina(n6752), .dinb(n6379), .dout(n6755));
  jnot g06502(.din(n6755), .dout(n6756));
  jand g06503(.dina(n6756), .dinb(n6754), .dout(n6757));
  jnot g06504(.din(n6757), .dout(n6758));
  jor  g06505(.dina(n6758), .dinb(n6750), .dout(n6759));
  jand g06506(.dina(n6759), .dinb(n6749), .dout(n6760));
  jor  g06507(.dina(n6760), .dinb(n595), .dout(n6761));
  jand g06508(.dina(n6749), .dinb(n595), .dout(n6762));
  jand g06509(.dina(n6762), .dinb(n6759), .dout(n6763));
  jnot g06510(.din(n6381), .dout(n6764));
  jand g06511(.dina(asqrt[29] ), .dinb(n6764), .dout(n6765));
  jand g06512(.dina(n6765), .dinb(n6388), .dout(n6766));
  jor  g06513(.dina(n6766), .dinb(n6386), .dout(n6767));
  jand g06514(.dina(n6765), .dinb(n6389), .dout(n6768));
  jnot g06515(.din(n6768), .dout(n6769));
  jand g06516(.dina(n6769), .dinb(n6767), .dout(n6770));
  jnot g06517(.din(n6770), .dout(n6771));
  jor  g06518(.dina(n6771), .dinb(n6763), .dout(n6772));
  jand g06519(.dina(n6772), .dinb(n6761), .dout(n6773));
  jor  g06520(.dina(n6773), .dinb(n590), .dout(n6774));
  jxor g06521(.dina(n6390), .dinb(n595), .dout(n6775));
  jor  g06522(.dina(n6775), .dinb(n6505), .dout(n6776));
  jxor g06523(.dina(n6776), .dinb(n6401), .dout(n6777));
  jand g06524(.dina(n6773), .dinb(n590), .dout(n6778));
  jor  g06525(.dina(n6778), .dinb(n6777), .dout(n6779));
  jand g06526(.dina(n6779), .dinb(n6774), .dout(n6780));
  jor  g06527(.dina(n6780), .dinb(n430), .dout(n6781));
  jnot g06528(.din(n6406), .dout(n6782));
  jor  g06529(.dina(n6782), .dinb(n6404), .dout(n6783));
  jor  g06530(.dina(n6783), .dinb(n6505), .dout(n6784));
  jxor g06531(.dina(n6784), .dinb(n6415), .dout(n6785));
  jand g06532(.dina(n6774), .dinb(n430), .dout(n6786));
  jand g06533(.dina(n6786), .dinb(n6779), .dout(n6787));
  jor  g06534(.dina(n6787), .dinb(n6785), .dout(n6788));
  jand g06535(.dina(n6788), .dinb(n6781), .dout(n6789));
  jor  g06536(.dina(n6789), .dinb(n425), .dout(n6790));
  jand g06537(.dina(n6789), .dinb(n425), .dout(n6791));
  jnot g06538(.din(n6418), .dout(n6792));
  jand g06539(.dina(asqrt[29] ), .dinb(n6792), .dout(n6793));
  jand g06540(.dina(n6793), .dinb(n6423), .dout(n6794));
  jor  g06541(.dina(n6794), .dinb(n6422), .dout(n6795));
  jand g06542(.dina(n6793), .dinb(n6424), .dout(n6796));
  jnot g06543(.din(n6796), .dout(n6797));
  jand g06544(.dina(n6797), .dinb(n6795), .dout(n6798));
  jnot g06545(.din(n6798), .dout(n6799));
  jor  g06546(.dina(n6799), .dinb(n6791), .dout(n6800));
  jand g06547(.dina(n6800), .dinb(n6790), .dout(n6801));
  jor  g06548(.dina(n6801), .dinb(n305), .dout(n6802));
  jand g06549(.dina(n6790), .dinb(n305), .dout(n6803));
  jand g06550(.dina(n6803), .dinb(n6800), .dout(n6804));
  jnot g06551(.din(n6426), .dout(n6805));
  jand g06552(.dina(asqrt[29] ), .dinb(n6805), .dout(n6806));
  jand g06553(.dina(n6806), .dinb(n6433), .dout(n6807));
  jor  g06554(.dina(n6807), .dinb(n6431), .dout(n6808));
  jand g06555(.dina(n6806), .dinb(n6434), .dout(n6809));
  jnot g06556(.din(n6809), .dout(n6810));
  jand g06557(.dina(n6810), .dinb(n6808), .dout(n6811));
  jnot g06558(.din(n6811), .dout(n6812));
  jor  g06559(.dina(n6812), .dinb(n6804), .dout(n6813));
  jand g06560(.dina(n6813), .dinb(n6802), .dout(n6814));
  jor  g06561(.dina(n6814), .dinb(n290), .dout(n6815));
  jxor g06562(.dina(n6435), .dinb(n305), .dout(n6816));
  jor  g06563(.dina(n6816), .dinb(n6505), .dout(n6817));
  jxor g06564(.dina(n6817), .dinb(n6446), .dout(n6818));
  jand g06565(.dina(n6814), .dinb(n290), .dout(n6819));
  jor  g06566(.dina(n6819), .dinb(n6818), .dout(n6820));
  jand g06567(.dina(n6820), .dinb(n6815), .dout(n6821));
  jor  g06568(.dina(n6821), .dinb(n223), .dout(n6822));
  jnot g06569(.din(n6451), .dout(n6823));
  jor  g06570(.dina(n6823), .dinb(n6449), .dout(n6824));
  jor  g06571(.dina(n6824), .dinb(n6505), .dout(n6825));
  jxor g06572(.dina(n6825), .dinb(n6460), .dout(n6826));
  jand g06573(.dina(n6815), .dinb(n223), .dout(n6827));
  jand g06574(.dina(n6827), .dinb(n6820), .dout(n6828));
  jor  g06575(.dina(n6828), .dinb(n6826), .dout(n6829));
  jand g06576(.dina(n6829), .dinb(n6822), .dout(n6830));
  jor  g06577(.dina(n6830), .dinb(n199), .dout(n6831));
  jand g06578(.dina(n6830), .dinb(n199), .dout(n6832));
  jnot g06579(.din(n6463), .dout(n6833));
  jand g06580(.dina(asqrt[29] ), .dinb(n6833), .dout(n6834));
  jand g06581(.dina(n6834), .dinb(n6468), .dout(n6835));
  jor  g06582(.dina(n6835), .dinb(n6467), .dout(n6836));
  jand g06583(.dina(n6834), .dinb(n6469), .dout(n6837));
  jnot g06584(.din(n6837), .dout(n6838));
  jand g06585(.dina(n6838), .dinb(n6836), .dout(n6839));
  jnot g06586(.din(n6839), .dout(n6840));
  jor  g06587(.dina(n6840), .dinb(n6832), .dout(n6841));
  jand g06588(.dina(n6841), .dinb(n6831), .dout(n6842));
  jnot g06589(.din(n6471), .dout(n6843));
  jand g06590(.dina(asqrt[29] ), .dinb(n6843), .dout(n6844));
  jand g06591(.dina(n6844), .dinb(n6478), .dout(n6845));
  jor  g06592(.dina(n6845), .dinb(n6476), .dout(n6846));
  jand g06593(.dina(n6844), .dinb(n6479), .dout(n6847));
  jnot g06594(.din(n6847), .dout(n6848));
  jand g06595(.dina(n6848), .dinb(n6846), .dout(n6849));
  jnot g06596(.din(n6849), .dout(n6850));
  jand g06597(.dina(asqrt[29] ), .dinb(n6493), .dout(n6851));
  jand g06598(.dina(n6851), .dinb(n6480), .dout(n6852));
  jor  g06599(.dina(n6852), .dinb(n6527), .dout(n6853));
  jor  g06600(.dina(n6853), .dinb(n6850), .dout(n6854));
  jor  g06601(.dina(n6854), .dinb(n6842), .dout(n6855));
  jand g06602(.dina(n6855), .dinb(n194), .dout(n6856));
  jand g06603(.dina(n6850), .dinb(n6842), .dout(n6857));
  jor  g06604(.dina(n6851), .dinb(n6480), .dout(n6858));
  jand g06605(.dina(n6493), .dinb(n6480), .dout(n6859));
  jor  g06606(.dina(n6859), .dinb(n194), .dout(n6860));
  jnot g06607(.din(n6860), .dout(n6861));
  jand g06608(.dina(n6861), .dinb(n6858), .dout(n6862));
  jor  g06609(.dina(n6862), .dinb(n6857), .dout(n6865));
  jor  g06610(.dina(n6865), .dinb(n6856), .dout(asqrt[28] ));
  jxor g06611(.dina(n6555), .dinb(n5116), .dout(n6867));
  jand g06612(.dina(n6867), .dinb(asqrt[28] ), .dout(n6868));
  jxor g06613(.dina(n6868), .dinb(n6508), .dout(n6869));
  jnot g06614(.din(n6869), .dout(n6870));
  jand g06615(.dina(asqrt[28] ), .dinb(a[56] ), .dout(n6871));
  jnot g06616(.din(a[54] ), .dout(n6872));
  jnot g06617(.din(a[55] ), .dout(n6873));
  jand g06618(.dina(n6510), .dinb(n6873), .dout(n6874));
  jand g06619(.dina(n6874), .dinb(n6872), .dout(n6875));
  jor  g06620(.dina(n6875), .dinb(n6871), .dout(n6876));
  jand g06621(.dina(n6876), .dinb(asqrt[29] ), .dout(n6877));
  jand g06622(.dina(asqrt[28] ), .dinb(n6510), .dout(n6878));
  jxor g06623(.dina(n6878), .dinb(n6511), .dout(n6879));
  jor  g06624(.dina(n6876), .dinb(asqrt[29] ), .dout(n6880));
  jand g06625(.dina(n6880), .dinb(n6879), .dout(n6881));
  jor  g06626(.dina(n6881), .dinb(n6877), .dout(n6882));
  jand g06627(.dina(n6882), .dinb(asqrt[30] ), .dout(n6883));
  jor  g06628(.dina(n6877), .dinb(asqrt[30] ), .dout(n6884));
  jor  g06629(.dina(n6884), .dinb(n6881), .dout(n6885));
  jand g06630(.dina(n6878), .dinb(n6511), .dout(n6886));
  jnot g06631(.din(n6856), .dout(n6887));
  jnot g06632(.din(n6857), .dout(n6888));
  jnot g06633(.din(n6862), .dout(n6889));
  jand g06634(.dina(n6889), .dinb(asqrt[29] ), .dout(n6890));
  jand g06635(.dina(n6890), .dinb(n6888), .dout(n6891));
  jand g06636(.dina(n6891), .dinb(n6887), .dout(n6892));
  jor  g06637(.dina(n6892), .dinb(n6886), .dout(n6893));
  jxor g06638(.dina(n6893), .dinb(n6134), .dout(n6894));
  jand g06639(.dina(n6894), .dinb(n6885), .dout(n6895));
  jor  g06640(.dina(n6895), .dinb(n6883), .dout(n6896));
  jand g06641(.dina(n6896), .dinb(asqrt[31] ), .dout(n6897));
  jor  g06642(.dina(n6896), .dinb(asqrt[31] ), .dout(n6898));
  jxor g06643(.dina(n6515), .dinb(n6500), .dout(n6899));
  jand g06644(.dina(n6899), .dinb(asqrt[28] ), .dout(n6900));
  jxor g06645(.dina(n6900), .dinb(n6518), .dout(n6901));
  jnot g06646(.din(n6901), .dout(n6902));
  jand g06647(.dina(n6902), .dinb(n6898), .dout(n6903));
  jor  g06648(.dina(n6903), .dinb(n6897), .dout(n6904));
  jand g06649(.dina(n6904), .dinb(asqrt[32] ), .dout(n6905));
  jnot g06650(.din(n6524), .dout(n6906));
  jand g06651(.dina(n6906), .dinb(n6522), .dout(n6907));
  jand g06652(.dina(n6907), .dinb(asqrt[28] ), .dout(n6908));
  jxor g06653(.dina(n6908), .dinb(n6532), .dout(n6909));
  jnot g06654(.din(n6909), .dout(n6910));
  jor  g06655(.dina(n6897), .dinb(asqrt[32] ), .dout(n6911));
  jor  g06656(.dina(n6911), .dinb(n6903), .dout(n6912));
  jand g06657(.dina(n6912), .dinb(n6910), .dout(n6913));
  jor  g06658(.dina(n6913), .dinb(n6905), .dout(n6914));
  jand g06659(.dina(n6914), .dinb(asqrt[33] ), .dout(n6915));
  jor  g06660(.dina(n6914), .dinb(asqrt[33] ), .dout(n6916));
  jnot g06661(.din(n6539), .dout(n6917));
  jxor g06662(.dina(n6534), .dinb(n5788), .dout(n6918));
  jand g06663(.dina(n6918), .dinb(asqrt[28] ), .dout(n6919));
  jxor g06664(.dina(n6919), .dinb(n6917), .dout(n6920));
  jand g06665(.dina(n6920), .dinb(n6916), .dout(n6921));
  jor  g06666(.dina(n6921), .dinb(n6915), .dout(n6922));
  jand g06667(.dina(n6922), .dinb(asqrt[34] ), .dout(n6923));
  jnot g06668(.din(n6544), .dout(n6924));
  jand g06669(.dina(n6924), .dinb(n6542), .dout(n6925));
  jand g06670(.dina(n6925), .dinb(asqrt[28] ), .dout(n6926));
  jxor g06671(.dina(n6926), .dinb(n6553), .dout(n6927));
  jnot g06672(.din(n6927), .dout(n6928));
  jor  g06673(.dina(n6915), .dinb(asqrt[34] ), .dout(n6929));
  jor  g06674(.dina(n6929), .dinb(n6921), .dout(n6930));
  jand g06675(.dina(n6930), .dinb(n6928), .dout(n6931));
  jor  g06676(.dina(n6931), .dinb(n6923), .dout(n6932));
  jand g06677(.dina(n6932), .dinb(asqrt[35] ), .dout(n6933));
  jor  g06678(.dina(n6932), .dinb(asqrt[35] ), .dout(n6934));
  jand g06679(.dina(n6934), .dinb(n6869), .dout(n6935));
  jor  g06680(.dina(n6935), .dinb(n6933), .dout(n6936));
  jand g06681(.dina(n6936), .dinb(asqrt[36] ), .dout(n6937));
  jor  g06682(.dina(n6933), .dinb(asqrt[36] ), .dout(n6938));
  jor  g06683(.dina(n6938), .dinb(n6935), .dout(n6939));
  jnot g06684(.din(n6565), .dout(n6940));
  jnot g06685(.din(n6567), .dout(n6941));
  jand g06686(.dina(asqrt[28] ), .dinb(n6561), .dout(n6942));
  jand g06687(.dina(n6942), .dinb(n6941), .dout(n6943));
  jor  g06688(.dina(n6943), .dinb(n6940), .dout(n6944));
  jnot g06689(.din(n6568), .dout(n6945));
  jand g06690(.dina(n6942), .dinb(n6945), .dout(n6946));
  jnot g06691(.din(n6946), .dout(n6947));
  jand g06692(.dina(n6947), .dinb(n6944), .dout(n6948));
  jand g06693(.dina(n6948), .dinb(n6939), .dout(n6949));
  jor  g06694(.dina(n6949), .dinb(n6937), .dout(n6950));
  jand g06695(.dina(n6950), .dinb(asqrt[37] ), .dout(n6951));
  jor  g06696(.dina(n6950), .dinb(asqrt[37] ), .dout(n6952));
  jxor g06697(.dina(n6569), .dinb(n4494), .dout(n6953));
  jand g06698(.dina(n6953), .dinb(asqrt[28] ), .dout(n6954));
  jxor g06699(.dina(n6954), .dinb(n6575), .dout(n6955));
  jand g06700(.dina(n6955), .dinb(n6952), .dout(n6956));
  jor  g06701(.dina(n6956), .dinb(n6951), .dout(n6957));
  jand g06702(.dina(n6957), .dinb(asqrt[38] ), .dout(n6958));
  jor  g06703(.dina(n6951), .dinb(asqrt[38] ), .dout(n6959));
  jor  g06704(.dina(n6959), .dinb(n6956), .dout(n6960));
  jnot g06705(.din(n6583), .dout(n6961));
  jnot g06706(.din(n6585), .dout(n6962));
  jand g06707(.dina(asqrt[28] ), .dinb(n6579), .dout(n6963));
  jand g06708(.dina(n6963), .dinb(n6962), .dout(n6964));
  jor  g06709(.dina(n6964), .dinb(n6961), .dout(n6965));
  jnot g06710(.din(n6586), .dout(n6966));
  jand g06711(.dina(n6963), .dinb(n6966), .dout(n6967));
  jnot g06712(.din(n6967), .dout(n6968));
  jand g06713(.dina(n6968), .dinb(n6965), .dout(n6969));
  jand g06714(.dina(n6969), .dinb(n6960), .dout(n6970));
  jor  g06715(.dina(n6970), .dinb(n6958), .dout(n6971));
  jand g06716(.dina(n6971), .dinb(asqrt[39] ), .dout(n6972));
  jxor g06717(.dina(n6587), .dinb(n3907), .dout(n6973));
  jand g06718(.dina(n6973), .dinb(asqrt[28] ), .dout(n6974));
  jxor g06719(.dina(n6974), .dinb(n6594), .dout(n6975));
  jnot g06720(.din(n6975), .dout(n6976));
  jor  g06721(.dina(n6971), .dinb(asqrt[39] ), .dout(n6977));
  jand g06722(.dina(n6977), .dinb(n6976), .dout(n6978));
  jor  g06723(.dina(n6978), .dinb(n6972), .dout(n6979));
  jand g06724(.dina(n6979), .dinb(asqrt[40] ), .dout(n6980));
  jnot g06725(.din(n6599), .dout(n6981));
  jand g06726(.dina(n6981), .dinb(n6597), .dout(n6982));
  jand g06727(.dina(n6982), .dinb(asqrt[28] ), .dout(n6983));
  jxor g06728(.dina(n6983), .dinb(n6607), .dout(n6984));
  jnot g06729(.din(n6984), .dout(n6985));
  jor  g06730(.dina(n6972), .dinb(asqrt[40] ), .dout(n6986));
  jor  g06731(.dina(n6986), .dinb(n6978), .dout(n6987));
  jand g06732(.dina(n6987), .dinb(n6985), .dout(n6988));
  jor  g06733(.dina(n6988), .dinb(n6980), .dout(n6989));
  jand g06734(.dina(n6989), .dinb(asqrt[41] ), .dout(n6990));
  jor  g06735(.dina(n6989), .dinb(asqrt[41] ), .dout(n6991));
  jnot g06736(.din(n6613), .dout(n6992));
  jnot g06737(.din(n6614), .dout(n6993));
  jand g06738(.dina(asqrt[28] ), .dinb(n6610), .dout(n6994));
  jand g06739(.dina(n6994), .dinb(n6993), .dout(n6995));
  jor  g06740(.dina(n6995), .dinb(n6992), .dout(n6996));
  jnot g06741(.din(n6615), .dout(n6997));
  jand g06742(.dina(n6994), .dinb(n6997), .dout(n6998));
  jnot g06743(.din(n6998), .dout(n6999));
  jand g06744(.dina(n6999), .dinb(n6996), .dout(n7000));
  jand g06745(.dina(n7000), .dinb(n6991), .dout(n7001));
  jor  g06746(.dina(n7001), .dinb(n6990), .dout(n7002));
  jand g06747(.dina(n7002), .dinb(asqrt[42] ), .dout(n7003));
  jor  g06748(.dina(n6990), .dinb(asqrt[42] ), .dout(n7004));
  jor  g06749(.dina(n7004), .dinb(n7001), .dout(n7005));
  jnot g06750(.din(n6621), .dout(n7006));
  jnot g06751(.din(n6623), .dout(n7007));
  jand g06752(.dina(asqrt[28] ), .dinb(n6617), .dout(n7008));
  jand g06753(.dina(n7008), .dinb(n7007), .dout(n7009));
  jor  g06754(.dina(n7009), .dinb(n7006), .dout(n7010));
  jnot g06755(.din(n6624), .dout(n7011));
  jand g06756(.dina(n7008), .dinb(n7011), .dout(n7012));
  jnot g06757(.din(n7012), .dout(n7013));
  jand g06758(.dina(n7013), .dinb(n7010), .dout(n7014));
  jand g06759(.dina(n7014), .dinb(n7005), .dout(n7015));
  jor  g06760(.dina(n7015), .dinb(n7003), .dout(n7016));
  jand g06761(.dina(n7016), .dinb(asqrt[43] ), .dout(n7017));
  jxor g06762(.dina(n6625), .dinb(n2870), .dout(n7018));
  jand g06763(.dina(n7018), .dinb(asqrt[28] ), .dout(n7019));
  jxor g06764(.dina(n7019), .dinb(n6635), .dout(n7020));
  jnot g06765(.din(n7020), .dout(n7021));
  jor  g06766(.dina(n7016), .dinb(asqrt[43] ), .dout(n7022));
  jand g06767(.dina(n7022), .dinb(n7021), .dout(n7023));
  jor  g06768(.dina(n7023), .dinb(n7017), .dout(n7024));
  jand g06769(.dina(n7024), .dinb(asqrt[44] ), .dout(n7025));
  jnot g06770(.din(n6640), .dout(n7026));
  jand g06771(.dina(n7026), .dinb(n6638), .dout(n7027));
  jand g06772(.dina(n7027), .dinb(asqrt[28] ), .dout(n7028));
  jxor g06773(.dina(n7028), .dinb(n6648), .dout(n7029));
  jnot g06774(.din(n7029), .dout(n7030));
  jor  g06775(.dina(n7017), .dinb(asqrt[44] ), .dout(n7031));
  jor  g06776(.dina(n7031), .dinb(n7023), .dout(n7032));
  jand g06777(.dina(n7032), .dinb(n7030), .dout(n7033));
  jor  g06778(.dina(n7033), .dinb(n7025), .dout(n7034));
  jand g06779(.dina(n7034), .dinb(asqrt[45] ), .dout(n7035));
  jor  g06780(.dina(n7034), .dinb(asqrt[45] ), .dout(n7036));
  jnot g06781(.din(n6654), .dout(n7037));
  jnot g06782(.din(n6655), .dout(n7038));
  jand g06783(.dina(asqrt[28] ), .dinb(n6651), .dout(n7039));
  jand g06784(.dina(n7039), .dinb(n7038), .dout(n7040));
  jor  g06785(.dina(n7040), .dinb(n7037), .dout(n7041));
  jnot g06786(.din(n6656), .dout(n7042));
  jand g06787(.dina(n7039), .dinb(n7042), .dout(n7043));
  jnot g06788(.din(n7043), .dout(n7044));
  jand g06789(.dina(n7044), .dinb(n7041), .dout(n7045));
  jand g06790(.dina(n7045), .dinb(n7036), .dout(n7046));
  jor  g06791(.dina(n7046), .dinb(n7035), .dout(n7047));
  jand g06792(.dina(n7047), .dinb(asqrt[46] ), .dout(n7048));
  jor  g06793(.dina(n7035), .dinb(asqrt[46] ), .dout(n7049));
  jor  g06794(.dina(n7049), .dinb(n7046), .dout(n7050));
  jnot g06795(.din(n6662), .dout(n7051));
  jnot g06796(.din(n6664), .dout(n7052));
  jand g06797(.dina(asqrt[28] ), .dinb(n6658), .dout(n7053));
  jand g06798(.dina(n7053), .dinb(n7052), .dout(n7054));
  jor  g06799(.dina(n7054), .dinb(n7051), .dout(n7055));
  jnot g06800(.din(n6665), .dout(n7056));
  jand g06801(.dina(n7053), .dinb(n7056), .dout(n7057));
  jnot g06802(.din(n7057), .dout(n7058));
  jand g06803(.dina(n7058), .dinb(n7055), .dout(n7059));
  jand g06804(.dina(n7059), .dinb(n7050), .dout(n7060));
  jor  g06805(.dina(n7060), .dinb(n7048), .dout(n7061));
  jand g06806(.dina(n7061), .dinb(asqrt[47] ), .dout(n7062));
  jxor g06807(.dina(n6666), .dinb(n2005), .dout(n7063));
  jand g06808(.dina(n7063), .dinb(asqrt[28] ), .dout(n7064));
  jxor g06809(.dina(n7064), .dinb(n6676), .dout(n7065));
  jnot g06810(.din(n7065), .dout(n7066));
  jor  g06811(.dina(n7061), .dinb(asqrt[47] ), .dout(n7067));
  jand g06812(.dina(n7067), .dinb(n7066), .dout(n7068));
  jor  g06813(.dina(n7068), .dinb(n7062), .dout(n7069));
  jand g06814(.dina(n7069), .dinb(asqrt[48] ), .dout(n7070));
  jnot g06815(.din(n6681), .dout(n7071));
  jand g06816(.dina(n7071), .dinb(n6679), .dout(n7072));
  jand g06817(.dina(n7072), .dinb(asqrt[28] ), .dout(n7073));
  jxor g06818(.dina(n7073), .dinb(n6689), .dout(n7074));
  jnot g06819(.din(n7074), .dout(n7075));
  jor  g06820(.dina(n7062), .dinb(asqrt[48] ), .dout(n7076));
  jor  g06821(.dina(n7076), .dinb(n7068), .dout(n7077));
  jand g06822(.dina(n7077), .dinb(n7075), .dout(n7078));
  jor  g06823(.dina(n7078), .dinb(n7070), .dout(n7079));
  jand g06824(.dina(n7079), .dinb(asqrt[49] ), .dout(n7080));
  jor  g06825(.dina(n7079), .dinb(asqrt[49] ), .dout(n7081));
  jnot g06826(.din(n6695), .dout(n7082));
  jnot g06827(.din(n6696), .dout(n7083));
  jand g06828(.dina(asqrt[28] ), .dinb(n6692), .dout(n7084));
  jand g06829(.dina(n7084), .dinb(n7083), .dout(n7085));
  jor  g06830(.dina(n7085), .dinb(n7082), .dout(n7086));
  jnot g06831(.din(n6697), .dout(n7087));
  jand g06832(.dina(n7084), .dinb(n7087), .dout(n7088));
  jnot g06833(.din(n7088), .dout(n7089));
  jand g06834(.dina(n7089), .dinb(n7086), .dout(n7090));
  jand g06835(.dina(n7090), .dinb(n7081), .dout(n7091));
  jor  g06836(.dina(n7091), .dinb(n7080), .dout(n7092));
  jand g06837(.dina(n7092), .dinb(asqrt[50] ), .dout(n7093));
  jor  g06838(.dina(n7080), .dinb(asqrt[50] ), .dout(n7094));
  jor  g06839(.dina(n7094), .dinb(n7091), .dout(n7095));
  jnot g06840(.din(n6703), .dout(n7096));
  jnot g06841(.din(n6705), .dout(n7097));
  jand g06842(.dina(asqrt[28] ), .dinb(n6699), .dout(n7098));
  jand g06843(.dina(n7098), .dinb(n7097), .dout(n7099));
  jor  g06844(.dina(n7099), .dinb(n7096), .dout(n7100));
  jnot g06845(.din(n6706), .dout(n7101));
  jand g06846(.dina(n7098), .dinb(n7101), .dout(n7102));
  jnot g06847(.din(n7102), .dout(n7103));
  jand g06848(.dina(n7103), .dinb(n7100), .dout(n7104));
  jand g06849(.dina(n7104), .dinb(n7095), .dout(n7105));
  jor  g06850(.dina(n7105), .dinb(n7093), .dout(n7106));
  jand g06851(.dina(n7106), .dinb(asqrt[51] ), .dout(n7107));
  jxor g06852(.dina(n6707), .dinb(n1312), .dout(n7108));
  jand g06853(.dina(n7108), .dinb(asqrt[28] ), .dout(n7109));
  jxor g06854(.dina(n7109), .dinb(n6717), .dout(n7110));
  jnot g06855(.din(n7110), .dout(n7111));
  jor  g06856(.dina(n7106), .dinb(asqrt[51] ), .dout(n7112));
  jand g06857(.dina(n7112), .dinb(n7111), .dout(n7113));
  jor  g06858(.dina(n7113), .dinb(n7107), .dout(n7114));
  jand g06859(.dina(n7114), .dinb(asqrt[52] ), .dout(n7115));
  jnot g06860(.din(n6722), .dout(n7116));
  jand g06861(.dina(n7116), .dinb(n6720), .dout(n7117));
  jand g06862(.dina(n7117), .dinb(asqrt[28] ), .dout(n7118));
  jxor g06863(.dina(n7118), .dinb(n6730), .dout(n7119));
  jnot g06864(.din(n7119), .dout(n7120));
  jor  g06865(.dina(n7107), .dinb(asqrt[52] ), .dout(n7121));
  jor  g06866(.dina(n7121), .dinb(n7113), .dout(n7122));
  jand g06867(.dina(n7122), .dinb(n7120), .dout(n7123));
  jor  g06868(.dina(n7123), .dinb(n7115), .dout(n7124));
  jand g06869(.dina(n7124), .dinb(asqrt[53] ), .dout(n7125));
  jor  g06870(.dina(n7124), .dinb(asqrt[53] ), .dout(n7126));
  jnot g06871(.din(n6736), .dout(n7127));
  jnot g06872(.din(n6737), .dout(n7128));
  jand g06873(.dina(asqrt[28] ), .dinb(n6733), .dout(n7129));
  jand g06874(.dina(n7129), .dinb(n7128), .dout(n7130));
  jor  g06875(.dina(n7130), .dinb(n7127), .dout(n7131));
  jnot g06876(.din(n6738), .dout(n7132));
  jand g06877(.dina(n7129), .dinb(n7132), .dout(n7133));
  jnot g06878(.din(n7133), .dout(n7134));
  jand g06879(.dina(n7134), .dinb(n7131), .dout(n7135));
  jand g06880(.dina(n7135), .dinb(n7126), .dout(n7136));
  jor  g06881(.dina(n7136), .dinb(n7125), .dout(n7137));
  jand g06882(.dina(n7137), .dinb(asqrt[54] ), .dout(n7138));
  jor  g06883(.dina(n7125), .dinb(asqrt[54] ), .dout(n7139));
  jor  g06884(.dina(n7139), .dinb(n7136), .dout(n7140));
  jnot g06885(.din(n6744), .dout(n7141));
  jnot g06886(.din(n6746), .dout(n7142));
  jand g06887(.dina(asqrt[28] ), .dinb(n6740), .dout(n7143));
  jand g06888(.dina(n7143), .dinb(n7142), .dout(n7144));
  jor  g06889(.dina(n7144), .dinb(n7141), .dout(n7145));
  jnot g06890(.din(n6747), .dout(n7146));
  jand g06891(.dina(n7143), .dinb(n7146), .dout(n7147));
  jnot g06892(.din(n7147), .dout(n7148));
  jand g06893(.dina(n7148), .dinb(n7145), .dout(n7149));
  jand g06894(.dina(n7149), .dinb(n7140), .dout(n7150));
  jor  g06895(.dina(n7150), .dinb(n7138), .dout(n7151));
  jand g06896(.dina(n7151), .dinb(asqrt[55] ), .dout(n7152));
  jxor g06897(.dina(n6748), .dinb(n791), .dout(n7153));
  jand g06898(.dina(n7153), .dinb(asqrt[28] ), .dout(n7154));
  jxor g06899(.dina(n7154), .dinb(n6758), .dout(n7155));
  jnot g06900(.din(n7155), .dout(n7156));
  jor  g06901(.dina(n7151), .dinb(asqrt[55] ), .dout(n7157));
  jand g06902(.dina(n7157), .dinb(n7156), .dout(n7158));
  jor  g06903(.dina(n7158), .dinb(n7152), .dout(n7159));
  jand g06904(.dina(n7159), .dinb(asqrt[56] ), .dout(n7160));
  jnot g06905(.din(n6763), .dout(n7161));
  jand g06906(.dina(n7161), .dinb(n6761), .dout(n7162));
  jand g06907(.dina(n7162), .dinb(asqrt[28] ), .dout(n7163));
  jxor g06908(.dina(n7163), .dinb(n6771), .dout(n7164));
  jnot g06909(.din(n7164), .dout(n7165));
  jor  g06910(.dina(n7152), .dinb(asqrt[56] ), .dout(n7166));
  jor  g06911(.dina(n7166), .dinb(n7158), .dout(n7167));
  jand g06912(.dina(n7167), .dinb(n7165), .dout(n7168));
  jor  g06913(.dina(n7168), .dinb(n7160), .dout(n7169));
  jand g06914(.dina(n7169), .dinb(asqrt[57] ), .dout(n7170));
  jor  g06915(.dina(n7169), .dinb(asqrt[57] ), .dout(n7171));
  jnot g06916(.din(n6777), .dout(n7172));
  jnot g06917(.din(n6778), .dout(n7173));
  jand g06918(.dina(asqrt[28] ), .dinb(n6774), .dout(n7174));
  jand g06919(.dina(n7174), .dinb(n7173), .dout(n7175));
  jor  g06920(.dina(n7175), .dinb(n7172), .dout(n7176));
  jnot g06921(.din(n6779), .dout(n7177));
  jand g06922(.dina(n7174), .dinb(n7177), .dout(n7178));
  jnot g06923(.din(n7178), .dout(n7179));
  jand g06924(.dina(n7179), .dinb(n7176), .dout(n7180));
  jand g06925(.dina(n7180), .dinb(n7171), .dout(n7181));
  jor  g06926(.dina(n7181), .dinb(n7170), .dout(n7182));
  jand g06927(.dina(n7182), .dinb(asqrt[58] ), .dout(n7183));
  jor  g06928(.dina(n7170), .dinb(asqrt[58] ), .dout(n7184));
  jor  g06929(.dina(n7184), .dinb(n7181), .dout(n7185));
  jnot g06930(.din(n6785), .dout(n7186));
  jnot g06931(.din(n6787), .dout(n7187));
  jand g06932(.dina(asqrt[28] ), .dinb(n6781), .dout(n7188));
  jand g06933(.dina(n7188), .dinb(n7187), .dout(n7189));
  jor  g06934(.dina(n7189), .dinb(n7186), .dout(n7190));
  jnot g06935(.din(n6788), .dout(n7191));
  jand g06936(.dina(n7188), .dinb(n7191), .dout(n7192));
  jnot g06937(.din(n7192), .dout(n7193));
  jand g06938(.dina(n7193), .dinb(n7190), .dout(n7194));
  jand g06939(.dina(n7194), .dinb(n7185), .dout(n7195));
  jor  g06940(.dina(n7195), .dinb(n7183), .dout(n7196));
  jand g06941(.dina(n7196), .dinb(asqrt[59] ), .dout(n7197));
  jxor g06942(.dina(n6789), .dinb(n425), .dout(n7198));
  jand g06943(.dina(n7198), .dinb(asqrt[28] ), .dout(n7199));
  jxor g06944(.dina(n7199), .dinb(n6799), .dout(n7200));
  jnot g06945(.din(n7200), .dout(n7201));
  jor  g06946(.dina(n7196), .dinb(asqrt[59] ), .dout(n7202));
  jand g06947(.dina(n7202), .dinb(n7201), .dout(n7203));
  jor  g06948(.dina(n7203), .dinb(n7197), .dout(n7204));
  jand g06949(.dina(n7204), .dinb(asqrt[60] ), .dout(n7205));
  jnot g06950(.din(n6804), .dout(n7206));
  jand g06951(.dina(n7206), .dinb(n6802), .dout(n7207));
  jand g06952(.dina(n7207), .dinb(asqrt[28] ), .dout(n7208));
  jxor g06953(.dina(n7208), .dinb(n6812), .dout(n7209));
  jnot g06954(.din(n7209), .dout(n7210));
  jor  g06955(.dina(n7197), .dinb(asqrt[60] ), .dout(n7211));
  jor  g06956(.dina(n7211), .dinb(n7203), .dout(n7212));
  jand g06957(.dina(n7212), .dinb(n7210), .dout(n7213));
  jor  g06958(.dina(n7213), .dinb(n7205), .dout(n7214));
  jand g06959(.dina(n7214), .dinb(asqrt[61] ), .dout(n7215));
  jor  g06960(.dina(n7214), .dinb(asqrt[61] ), .dout(n7216));
  jnot g06961(.din(n6818), .dout(n7217));
  jnot g06962(.din(n6819), .dout(n7218));
  jand g06963(.dina(asqrt[28] ), .dinb(n6815), .dout(n7219));
  jand g06964(.dina(n7219), .dinb(n7218), .dout(n7220));
  jor  g06965(.dina(n7220), .dinb(n7217), .dout(n7221));
  jnot g06966(.din(n6820), .dout(n7222));
  jand g06967(.dina(n7219), .dinb(n7222), .dout(n7223));
  jnot g06968(.din(n7223), .dout(n7224));
  jand g06969(.dina(n7224), .dinb(n7221), .dout(n7225));
  jand g06970(.dina(n7225), .dinb(n7216), .dout(n7226));
  jor  g06971(.dina(n7226), .dinb(n7215), .dout(n7227));
  jand g06972(.dina(n7227), .dinb(asqrt[62] ), .dout(n7228));
  jor  g06973(.dina(n7215), .dinb(asqrt[62] ), .dout(n7229));
  jor  g06974(.dina(n7229), .dinb(n7226), .dout(n7230));
  jnot g06975(.din(n6826), .dout(n7231));
  jnot g06976(.din(n6828), .dout(n7232));
  jand g06977(.dina(asqrt[28] ), .dinb(n6822), .dout(n7233));
  jand g06978(.dina(n7233), .dinb(n7232), .dout(n7234));
  jor  g06979(.dina(n7234), .dinb(n7231), .dout(n7235));
  jnot g06980(.din(n6829), .dout(n7236));
  jand g06981(.dina(n7233), .dinb(n7236), .dout(n7237));
  jnot g06982(.din(n7237), .dout(n7238));
  jand g06983(.dina(n7238), .dinb(n7235), .dout(n7239));
  jand g06984(.dina(n7239), .dinb(n7230), .dout(n7240));
  jor  g06985(.dina(n7240), .dinb(n7228), .dout(n7241));
  jxor g06986(.dina(n6830), .dinb(n199), .dout(n7242));
  jand g06987(.dina(n7242), .dinb(asqrt[28] ), .dout(n7243));
  jxor g06988(.dina(n7243), .dinb(n6840), .dout(n7244));
  jnot g06989(.din(n6842), .dout(n7245));
  jand g06990(.dina(asqrt[28] ), .dinb(n6849), .dout(n7246));
  jand g06991(.dina(n7246), .dinb(n7245), .dout(n7247));
  jor  g06992(.dina(n7247), .dinb(n6857), .dout(n7248));
  jor  g06993(.dina(n7248), .dinb(n7244), .dout(n7249));
  jnot g06994(.din(n7249), .dout(n7250));
  jand g06995(.dina(n7250), .dinb(n7241), .dout(n7251));
  jor  g06996(.dina(n7251), .dinb(asqrt[63] ), .dout(n7252));
  jnot g06997(.din(n7244), .dout(n7253));
  jor  g06998(.dina(n7253), .dinb(n7241), .dout(n7254));
  jor  g06999(.dina(n7246), .dinb(n7245), .dout(n7255));
  jand g07000(.dina(n6849), .dinb(n7245), .dout(n7256));
  jor  g07001(.dina(n7256), .dinb(n194), .dout(n7257));
  jnot g07002(.din(n7257), .dout(n7258));
  jand g07003(.dina(n7258), .dinb(n7255), .dout(n7259));
  jnot g07004(.din(asqrt[28] ), .dout(n7260));
  jnot g07005(.din(n7259), .dout(n7263));
  jand g07006(.dina(n7263), .dinb(n7254), .dout(n7264));
  jand g07007(.dina(n7264), .dinb(n7252), .dout(n7265));
  jxor g07008(.dina(n6932), .dinb(n4499), .dout(n7266));
  jor  g07009(.dina(n7266), .dinb(n7265), .dout(n7267));
  jxor g07010(.dina(n7267), .dinb(n6870), .dout(n7268));
  jnot g07011(.din(n7268), .dout(n7269));
  jor  g07012(.dina(n7265), .dinb(n6872), .dout(n7270));
  jnot g07013(.din(a[52] ), .dout(n7271));
  jnot g07014(.din(a[53] ), .dout(n7272));
  jand g07015(.dina(n6872), .dinb(n7272), .dout(n7273));
  jand g07016(.dina(n7273), .dinb(n7271), .dout(n7274));
  jnot g07017(.din(n7274), .dout(n7275));
  jand g07018(.dina(n7275), .dinb(n7270), .dout(n7276));
  jor  g07019(.dina(n7276), .dinb(n7260), .dout(n7277));
  jor  g07020(.dina(n7265), .dinb(a[54] ), .dout(n7278));
  jxor g07021(.dina(n7278), .dinb(n6873), .dout(n7279));
  jand g07022(.dina(n7276), .dinb(n7260), .dout(n7280));
  jor  g07023(.dina(n7280), .dinb(n7279), .dout(n7281));
  jand g07024(.dina(n7281), .dinb(n7277), .dout(n7282));
  jor  g07025(.dina(n7282), .dinb(n6505), .dout(n7283));
  jand g07026(.dina(n7277), .dinb(n6505), .dout(n7284));
  jand g07027(.dina(n7284), .dinb(n7281), .dout(n7285));
  jor  g07028(.dina(n7278), .dinb(a[55] ), .dout(n7286));
  jnot g07029(.din(n7252), .dout(n7287));
  jnot g07030(.din(n7254), .dout(n7288));
  jor  g07031(.dina(n7259), .dinb(n7260), .dout(n7289));
  jor  g07032(.dina(n7289), .dinb(n7288), .dout(n7290));
  jor  g07033(.dina(n7290), .dinb(n7287), .dout(n7291));
  jand g07034(.dina(n7291), .dinb(n7286), .dout(n7292));
  jxor g07035(.dina(n7292), .dinb(n6510), .dout(n7293));
  jor  g07036(.dina(n7293), .dinb(n7285), .dout(n7294));
  jand g07037(.dina(n7294), .dinb(n7283), .dout(n7295));
  jor  g07038(.dina(n7295), .dinb(n6500), .dout(n7296));
  jand g07039(.dina(n7295), .dinb(n6500), .dout(n7297));
  jxor g07040(.dina(n6876), .dinb(n6505), .dout(n7298));
  jor  g07041(.dina(n7298), .dinb(n7265), .dout(n7299));
  jxor g07042(.dina(n7299), .dinb(n6879), .dout(n7300));
  jor  g07043(.dina(n7300), .dinb(n7297), .dout(n7301));
  jand g07044(.dina(n7301), .dinb(n7296), .dout(n7302));
  jor  g07045(.dina(n7302), .dinb(n5793), .dout(n7303));
  jnot g07046(.din(n6885), .dout(n7304));
  jor  g07047(.dina(n7304), .dinb(n6883), .dout(n7305));
  jor  g07048(.dina(n7305), .dinb(n7265), .dout(n7306));
  jxor g07049(.dina(n7306), .dinb(n6894), .dout(n7307));
  jand g07050(.dina(n7296), .dinb(n5793), .dout(n7308));
  jand g07051(.dina(n7308), .dinb(n7301), .dout(n7309));
  jor  g07052(.dina(n7309), .dinb(n7307), .dout(n7310));
  jand g07053(.dina(n7310), .dinb(n7303), .dout(n7311));
  jor  g07054(.dina(n7311), .dinb(n5788), .dout(n7312));
  jand g07055(.dina(n7311), .dinb(n5788), .dout(n7313));
  jxor g07056(.dina(n6896), .dinb(n5793), .dout(n7314));
  jor  g07057(.dina(n7314), .dinb(n7265), .dout(n7315));
  jxor g07058(.dina(n7315), .dinb(n6901), .dout(n7316));
  jnot g07059(.din(n7316), .dout(n7317));
  jor  g07060(.dina(n7317), .dinb(n7313), .dout(n7318));
  jand g07061(.dina(n7318), .dinb(n7312), .dout(n7319));
  jor  g07062(.dina(n7319), .dinb(n5121), .dout(n7320));
  jand g07063(.dina(n7312), .dinb(n5121), .dout(n7321));
  jand g07064(.dina(n7321), .dinb(n7318), .dout(n7322));
  jnot g07065(.din(n6905), .dout(n7323));
  jnot g07066(.din(n7265), .dout(asqrt[27] ));
  jand g07067(.dina(asqrt[27] ), .dinb(n7323), .dout(n7325));
  jand g07068(.dina(n7325), .dinb(n6912), .dout(n7326));
  jor  g07069(.dina(n7326), .dinb(n6910), .dout(n7327));
  jand g07070(.dina(n7325), .dinb(n6913), .dout(n7328));
  jnot g07071(.din(n7328), .dout(n7329));
  jand g07072(.dina(n7329), .dinb(n7327), .dout(n7330));
  jnot g07073(.din(n7330), .dout(n7331));
  jor  g07074(.dina(n7331), .dinb(n7322), .dout(n7332));
  jand g07075(.dina(n7332), .dinb(n7320), .dout(n7333));
  jor  g07076(.dina(n7333), .dinb(n5116), .dout(n7334));
  jand g07077(.dina(n7333), .dinb(n5116), .dout(n7335));
  jnot g07078(.din(n6920), .dout(n7336));
  jxor g07079(.dina(n6914), .dinb(n5121), .dout(n7337));
  jor  g07080(.dina(n7337), .dinb(n7265), .dout(n7338));
  jxor g07081(.dina(n7338), .dinb(n7336), .dout(n7339));
  jnot g07082(.din(n7339), .dout(n7340));
  jor  g07083(.dina(n7340), .dinb(n7335), .dout(n7341));
  jand g07084(.dina(n7341), .dinb(n7334), .dout(n7342));
  jor  g07085(.dina(n7342), .dinb(n4499), .dout(n7343));
  jand g07086(.dina(n7334), .dinb(n4499), .dout(n7344));
  jand g07087(.dina(n7344), .dinb(n7341), .dout(n7345));
  jnot g07088(.din(n6923), .dout(n7346));
  jand g07089(.dina(asqrt[27] ), .dinb(n7346), .dout(n7347));
  jand g07090(.dina(n7347), .dinb(n6930), .dout(n7348));
  jor  g07091(.dina(n7348), .dinb(n6928), .dout(n7349));
  jand g07092(.dina(n7347), .dinb(n6931), .dout(n7350));
  jnot g07093(.din(n7350), .dout(n7351));
  jand g07094(.dina(n7351), .dinb(n7349), .dout(n7352));
  jnot g07095(.din(n7352), .dout(n7353));
  jor  g07096(.dina(n7353), .dinb(n7345), .dout(n7354));
  jand g07097(.dina(n7354), .dinb(n7343), .dout(n7355));
  jor  g07098(.dina(n7355), .dinb(n4494), .dout(n7356));
  jand g07099(.dina(n7355), .dinb(n4494), .dout(n7357));
  jor  g07100(.dina(n7357), .dinb(n7269), .dout(n7358));
  jand g07101(.dina(n7358), .dinb(n7356), .dout(n7359));
  jor  g07102(.dina(n7359), .dinb(n3912), .dout(n7360));
  jnot g07103(.din(n6939), .dout(n7361));
  jor  g07104(.dina(n7361), .dinb(n6937), .dout(n7362));
  jor  g07105(.dina(n7362), .dinb(n7265), .dout(n7363));
  jxor g07106(.dina(n7363), .dinb(n6948), .dout(n7364));
  jand g07107(.dina(n7356), .dinb(n3912), .dout(n7365));
  jand g07108(.dina(n7365), .dinb(n7358), .dout(n7366));
  jor  g07109(.dina(n7366), .dinb(n7364), .dout(n7367));
  jand g07110(.dina(n7367), .dinb(n7360), .dout(n7368));
  jor  g07111(.dina(n7368), .dinb(n3907), .dout(n7369));
  jxor g07112(.dina(n6950), .dinb(n3912), .dout(n7370));
  jor  g07113(.dina(n7370), .dinb(n7265), .dout(n7371));
  jxor g07114(.dina(n7371), .dinb(n6955), .dout(n7372));
  jand g07115(.dina(n7368), .dinb(n3907), .dout(n7373));
  jor  g07116(.dina(n7373), .dinb(n7372), .dout(n7374));
  jand g07117(.dina(n7374), .dinb(n7369), .dout(n7375));
  jor  g07118(.dina(n7375), .dinb(n3376), .dout(n7376));
  jnot g07119(.din(n6960), .dout(n7377));
  jor  g07120(.dina(n7377), .dinb(n6958), .dout(n7378));
  jor  g07121(.dina(n7378), .dinb(n7265), .dout(n7379));
  jxor g07122(.dina(n7379), .dinb(n6969), .dout(n7380));
  jand g07123(.dina(n7369), .dinb(n3376), .dout(n7381));
  jand g07124(.dina(n7381), .dinb(n7374), .dout(n7382));
  jor  g07125(.dina(n7382), .dinb(n7380), .dout(n7383));
  jand g07126(.dina(n7383), .dinb(n7376), .dout(n7384));
  jor  g07127(.dina(n7384), .dinb(n3371), .dout(n7385));
  jand g07128(.dina(n7384), .dinb(n3371), .dout(n7386));
  jnot g07129(.din(n6972), .dout(n7387));
  jand g07130(.dina(asqrt[27] ), .dinb(n7387), .dout(n7388));
  jand g07131(.dina(n7388), .dinb(n6977), .dout(n7389));
  jor  g07132(.dina(n7389), .dinb(n6976), .dout(n7390));
  jand g07133(.dina(n7388), .dinb(n6978), .dout(n7391));
  jnot g07134(.din(n7391), .dout(n7392));
  jand g07135(.dina(n7392), .dinb(n7390), .dout(n7393));
  jnot g07136(.din(n7393), .dout(n7394));
  jor  g07137(.dina(n7394), .dinb(n7386), .dout(n7395));
  jand g07138(.dina(n7395), .dinb(n7385), .dout(n7396));
  jor  g07139(.dina(n7396), .dinb(n2875), .dout(n7397));
  jand g07140(.dina(n7385), .dinb(n2875), .dout(n7398));
  jand g07141(.dina(n7398), .dinb(n7395), .dout(n7399));
  jnot g07142(.din(n6980), .dout(n7400));
  jand g07143(.dina(asqrt[27] ), .dinb(n7400), .dout(n7401));
  jand g07144(.dina(n7401), .dinb(n6987), .dout(n7402));
  jor  g07145(.dina(n7402), .dinb(n6985), .dout(n7403));
  jand g07146(.dina(n7401), .dinb(n6988), .dout(n7404));
  jnot g07147(.din(n7404), .dout(n7405));
  jand g07148(.dina(n7405), .dinb(n7403), .dout(n7406));
  jnot g07149(.din(n7406), .dout(n7407));
  jor  g07150(.dina(n7407), .dinb(n7399), .dout(n7408));
  jand g07151(.dina(n7408), .dinb(n7397), .dout(n7409));
  jor  g07152(.dina(n7409), .dinb(n2870), .dout(n7410));
  jxor g07153(.dina(n6989), .dinb(n2875), .dout(n7411));
  jor  g07154(.dina(n7411), .dinb(n7265), .dout(n7412));
  jxor g07155(.dina(n7412), .dinb(n7000), .dout(n7413));
  jand g07156(.dina(n7409), .dinb(n2870), .dout(n7414));
  jor  g07157(.dina(n7414), .dinb(n7413), .dout(n7415));
  jand g07158(.dina(n7415), .dinb(n7410), .dout(n7416));
  jor  g07159(.dina(n7416), .dinb(n2425), .dout(n7417));
  jnot g07160(.din(n7005), .dout(n7418));
  jor  g07161(.dina(n7418), .dinb(n7003), .dout(n7419));
  jor  g07162(.dina(n7419), .dinb(n7265), .dout(n7420));
  jxor g07163(.dina(n7420), .dinb(n7014), .dout(n7421));
  jand g07164(.dina(n7410), .dinb(n2425), .dout(n7422));
  jand g07165(.dina(n7422), .dinb(n7415), .dout(n7423));
  jor  g07166(.dina(n7423), .dinb(n7421), .dout(n7424));
  jand g07167(.dina(n7424), .dinb(n7417), .dout(n7425));
  jor  g07168(.dina(n7425), .dinb(n2420), .dout(n7426));
  jand g07169(.dina(n7425), .dinb(n2420), .dout(n7427));
  jnot g07170(.din(n7017), .dout(n7428));
  jand g07171(.dina(asqrt[27] ), .dinb(n7428), .dout(n7429));
  jand g07172(.dina(n7429), .dinb(n7022), .dout(n7430));
  jor  g07173(.dina(n7430), .dinb(n7021), .dout(n7431));
  jand g07174(.dina(n7429), .dinb(n7023), .dout(n7432));
  jnot g07175(.din(n7432), .dout(n7433));
  jand g07176(.dina(n7433), .dinb(n7431), .dout(n7434));
  jnot g07177(.din(n7434), .dout(n7435));
  jor  g07178(.dina(n7435), .dinb(n7427), .dout(n7436));
  jand g07179(.dina(n7436), .dinb(n7426), .dout(n7437));
  jor  g07180(.dina(n7437), .dinb(n2010), .dout(n7438));
  jand g07181(.dina(n7426), .dinb(n2010), .dout(n7439));
  jand g07182(.dina(n7439), .dinb(n7436), .dout(n7440));
  jnot g07183(.din(n7025), .dout(n7441));
  jand g07184(.dina(asqrt[27] ), .dinb(n7441), .dout(n7442));
  jand g07185(.dina(n7442), .dinb(n7032), .dout(n7443));
  jor  g07186(.dina(n7443), .dinb(n7030), .dout(n7444));
  jand g07187(.dina(n7442), .dinb(n7033), .dout(n7445));
  jnot g07188(.din(n7445), .dout(n7446));
  jand g07189(.dina(n7446), .dinb(n7444), .dout(n7447));
  jnot g07190(.din(n7447), .dout(n7448));
  jor  g07191(.dina(n7448), .dinb(n7440), .dout(n7449));
  jand g07192(.dina(n7449), .dinb(n7438), .dout(n7450));
  jor  g07193(.dina(n7450), .dinb(n2005), .dout(n7451));
  jxor g07194(.dina(n7034), .dinb(n2010), .dout(n7452));
  jor  g07195(.dina(n7452), .dinb(n7265), .dout(n7453));
  jxor g07196(.dina(n7453), .dinb(n7045), .dout(n7454));
  jand g07197(.dina(n7450), .dinb(n2005), .dout(n7455));
  jor  g07198(.dina(n7455), .dinb(n7454), .dout(n7456));
  jand g07199(.dina(n7456), .dinb(n7451), .dout(n7457));
  jor  g07200(.dina(n7457), .dinb(n1646), .dout(n7458));
  jnot g07201(.din(n7050), .dout(n7459));
  jor  g07202(.dina(n7459), .dinb(n7048), .dout(n7460));
  jor  g07203(.dina(n7460), .dinb(n7265), .dout(n7461));
  jxor g07204(.dina(n7461), .dinb(n7059), .dout(n7462));
  jand g07205(.dina(n7451), .dinb(n1646), .dout(n7463));
  jand g07206(.dina(n7463), .dinb(n7456), .dout(n7464));
  jor  g07207(.dina(n7464), .dinb(n7462), .dout(n7465));
  jand g07208(.dina(n7465), .dinb(n7458), .dout(n7466));
  jor  g07209(.dina(n7466), .dinb(n1641), .dout(n7467));
  jand g07210(.dina(n7466), .dinb(n1641), .dout(n7468));
  jnot g07211(.din(n7062), .dout(n7469));
  jand g07212(.dina(asqrt[27] ), .dinb(n7469), .dout(n7470));
  jand g07213(.dina(n7470), .dinb(n7067), .dout(n7471));
  jor  g07214(.dina(n7471), .dinb(n7066), .dout(n7472));
  jand g07215(.dina(n7470), .dinb(n7068), .dout(n7473));
  jnot g07216(.din(n7473), .dout(n7474));
  jand g07217(.dina(n7474), .dinb(n7472), .dout(n7475));
  jnot g07218(.din(n7475), .dout(n7476));
  jor  g07219(.dina(n7476), .dinb(n7468), .dout(n7477));
  jand g07220(.dina(n7477), .dinb(n7467), .dout(n7478));
  jor  g07221(.dina(n7478), .dinb(n1317), .dout(n7479));
  jand g07222(.dina(n7467), .dinb(n1317), .dout(n7480));
  jand g07223(.dina(n7480), .dinb(n7477), .dout(n7481));
  jnot g07224(.din(n7070), .dout(n7482));
  jand g07225(.dina(asqrt[27] ), .dinb(n7482), .dout(n7483));
  jand g07226(.dina(n7483), .dinb(n7077), .dout(n7484));
  jor  g07227(.dina(n7484), .dinb(n7075), .dout(n7485));
  jand g07228(.dina(n7483), .dinb(n7078), .dout(n7486));
  jnot g07229(.din(n7486), .dout(n7487));
  jand g07230(.dina(n7487), .dinb(n7485), .dout(n7488));
  jnot g07231(.din(n7488), .dout(n7489));
  jor  g07232(.dina(n7489), .dinb(n7481), .dout(n7490));
  jand g07233(.dina(n7490), .dinb(n7479), .dout(n7491));
  jor  g07234(.dina(n7491), .dinb(n1312), .dout(n7492));
  jxor g07235(.dina(n7079), .dinb(n1317), .dout(n7493));
  jor  g07236(.dina(n7493), .dinb(n7265), .dout(n7494));
  jxor g07237(.dina(n7494), .dinb(n7090), .dout(n7495));
  jand g07238(.dina(n7491), .dinb(n1312), .dout(n7496));
  jor  g07239(.dina(n7496), .dinb(n7495), .dout(n7497));
  jand g07240(.dina(n7497), .dinb(n7492), .dout(n7498));
  jor  g07241(.dina(n7498), .dinb(n1039), .dout(n7499));
  jnot g07242(.din(n7095), .dout(n7500));
  jor  g07243(.dina(n7500), .dinb(n7093), .dout(n7501));
  jor  g07244(.dina(n7501), .dinb(n7265), .dout(n7502));
  jxor g07245(.dina(n7502), .dinb(n7104), .dout(n7503));
  jand g07246(.dina(n7492), .dinb(n1039), .dout(n7504));
  jand g07247(.dina(n7504), .dinb(n7497), .dout(n7505));
  jor  g07248(.dina(n7505), .dinb(n7503), .dout(n7506));
  jand g07249(.dina(n7506), .dinb(n7499), .dout(n7507));
  jor  g07250(.dina(n7507), .dinb(n1034), .dout(n7508));
  jand g07251(.dina(n7507), .dinb(n1034), .dout(n7509));
  jnot g07252(.din(n7107), .dout(n7510));
  jand g07253(.dina(asqrt[27] ), .dinb(n7510), .dout(n7511));
  jand g07254(.dina(n7511), .dinb(n7112), .dout(n7512));
  jor  g07255(.dina(n7512), .dinb(n7111), .dout(n7513));
  jand g07256(.dina(n7511), .dinb(n7113), .dout(n7514));
  jnot g07257(.din(n7514), .dout(n7515));
  jand g07258(.dina(n7515), .dinb(n7513), .dout(n7516));
  jnot g07259(.din(n7516), .dout(n7517));
  jor  g07260(.dina(n7517), .dinb(n7509), .dout(n7518));
  jand g07261(.dina(n7518), .dinb(n7508), .dout(n7519));
  jor  g07262(.dina(n7519), .dinb(n796), .dout(n7520));
  jand g07263(.dina(n7508), .dinb(n796), .dout(n7521));
  jand g07264(.dina(n7521), .dinb(n7518), .dout(n7522));
  jnot g07265(.din(n7115), .dout(n7523));
  jand g07266(.dina(asqrt[27] ), .dinb(n7523), .dout(n7524));
  jand g07267(.dina(n7524), .dinb(n7122), .dout(n7525));
  jor  g07268(.dina(n7525), .dinb(n7120), .dout(n7526));
  jand g07269(.dina(n7524), .dinb(n7123), .dout(n7527));
  jnot g07270(.din(n7527), .dout(n7528));
  jand g07271(.dina(n7528), .dinb(n7526), .dout(n7529));
  jnot g07272(.din(n7529), .dout(n7530));
  jor  g07273(.dina(n7530), .dinb(n7522), .dout(n7531));
  jand g07274(.dina(n7531), .dinb(n7520), .dout(n7532));
  jor  g07275(.dina(n7532), .dinb(n791), .dout(n7533));
  jxor g07276(.dina(n7124), .dinb(n796), .dout(n7534));
  jor  g07277(.dina(n7534), .dinb(n7265), .dout(n7535));
  jxor g07278(.dina(n7535), .dinb(n7135), .dout(n7536));
  jand g07279(.dina(n7532), .dinb(n791), .dout(n7537));
  jor  g07280(.dina(n7537), .dinb(n7536), .dout(n7538));
  jand g07281(.dina(n7538), .dinb(n7533), .dout(n7539));
  jor  g07282(.dina(n7539), .dinb(n595), .dout(n7540));
  jnot g07283(.din(n7140), .dout(n7541));
  jor  g07284(.dina(n7541), .dinb(n7138), .dout(n7542));
  jor  g07285(.dina(n7542), .dinb(n7265), .dout(n7543));
  jxor g07286(.dina(n7543), .dinb(n7149), .dout(n7544));
  jand g07287(.dina(n7533), .dinb(n595), .dout(n7545));
  jand g07288(.dina(n7545), .dinb(n7538), .dout(n7546));
  jor  g07289(.dina(n7546), .dinb(n7544), .dout(n7547));
  jand g07290(.dina(n7547), .dinb(n7540), .dout(n7548));
  jor  g07291(.dina(n7548), .dinb(n590), .dout(n7549));
  jand g07292(.dina(n7548), .dinb(n590), .dout(n7550));
  jnot g07293(.din(n7152), .dout(n7551));
  jand g07294(.dina(asqrt[27] ), .dinb(n7551), .dout(n7552));
  jand g07295(.dina(n7552), .dinb(n7157), .dout(n7553));
  jor  g07296(.dina(n7553), .dinb(n7156), .dout(n7554));
  jand g07297(.dina(n7552), .dinb(n7158), .dout(n7555));
  jnot g07298(.din(n7555), .dout(n7556));
  jand g07299(.dina(n7556), .dinb(n7554), .dout(n7557));
  jnot g07300(.din(n7557), .dout(n7558));
  jor  g07301(.dina(n7558), .dinb(n7550), .dout(n7559));
  jand g07302(.dina(n7559), .dinb(n7549), .dout(n7560));
  jor  g07303(.dina(n7560), .dinb(n430), .dout(n7561));
  jand g07304(.dina(n7549), .dinb(n430), .dout(n7562));
  jand g07305(.dina(n7562), .dinb(n7559), .dout(n7563));
  jnot g07306(.din(n7160), .dout(n7564));
  jand g07307(.dina(asqrt[27] ), .dinb(n7564), .dout(n7565));
  jand g07308(.dina(n7565), .dinb(n7167), .dout(n7566));
  jor  g07309(.dina(n7566), .dinb(n7165), .dout(n7567));
  jand g07310(.dina(n7565), .dinb(n7168), .dout(n7568));
  jnot g07311(.din(n7568), .dout(n7569));
  jand g07312(.dina(n7569), .dinb(n7567), .dout(n7570));
  jnot g07313(.din(n7570), .dout(n7571));
  jor  g07314(.dina(n7571), .dinb(n7563), .dout(n7572));
  jand g07315(.dina(n7572), .dinb(n7561), .dout(n7573));
  jor  g07316(.dina(n7573), .dinb(n425), .dout(n7574));
  jxor g07317(.dina(n7169), .dinb(n430), .dout(n7575));
  jor  g07318(.dina(n7575), .dinb(n7265), .dout(n7576));
  jxor g07319(.dina(n7576), .dinb(n7180), .dout(n7577));
  jand g07320(.dina(n7573), .dinb(n425), .dout(n7578));
  jor  g07321(.dina(n7578), .dinb(n7577), .dout(n7579));
  jand g07322(.dina(n7579), .dinb(n7574), .dout(n7580));
  jor  g07323(.dina(n7580), .dinb(n305), .dout(n7581));
  jnot g07324(.din(n7185), .dout(n7582));
  jor  g07325(.dina(n7582), .dinb(n7183), .dout(n7583));
  jor  g07326(.dina(n7583), .dinb(n7265), .dout(n7584));
  jxor g07327(.dina(n7584), .dinb(n7194), .dout(n7585));
  jand g07328(.dina(n7574), .dinb(n305), .dout(n7586));
  jand g07329(.dina(n7586), .dinb(n7579), .dout(n7587));
  jor  g07330(.dina(n7587), .dinb(n7585), .dout(n7588));
  jand g07331(.dina(n7588), .dinb(n7581), .dout(n7589));
  jor  g07332(.dina(n7589), .dinb(n290), .dout(n7590));
  jand g07333(.dina(n7589), .dinb(n290), .dout(n7591));
  jnot g07334(.din(n7197), .dout(n7592));
  jand g07335(.dina(asqrt[27] ), .dinb(n7592), .dout(n7593));
  jand g07336(.dina(n7593), .dinb(n7202), .dout(n7594));
  jor  g07337(.dina(n7594), .dinb(n7201), .dout(n7595));
  jand g07338(.dina(n7593), .dinb(n7203), .dout(n7596));
  jnot g07339(.din(n7596), .dout(n7597));
  jand g07340(.dina(n7597), .dinb(n7595), .dout(n7598));
  jnot g07341(.din(n7598), .dout(n7599));
  jor  g07342(.dina(n7599), .dinb(n7591), .dout(n7600));
  jand g07343(.dina(n7600), .dinb(n7590), .dout(n7601));
  jor  g07344(.dina(n7601), .dinb(n223), .dout(n7602));
  jand g07345(.dina(n7590), .dinb(n223), .dout(n7603));
  jand g07346(.dina(n7603), .dinb(n7600), .dout(n7604));
  jnot g07347(.din(n7205), .dout(n7605));
  jand g07348(.dina(asqrt[27] ), .dinb(n7605), .dout(n7606));
  jand g07349(.dina(n7606), .dinb(n7212), .dout(n7607));
  jor  g07350(.dina(n7607), .dinb(n7210), .dout(n7608));
  jand g07351(.dina(n7606), .dinb(n7213), .dout(n7609));
  jnot g07352(.din(n7609), .dout(n7610));
  jand g07353(.dina(n7610), .dinb(n7608), .dout(n7611));
  jnot g07354(.din(n7611), .dout(n7612));
  jor  g07355(.dina(n7612), .dinb(n7604), .dout(n7613));
  jand g07356(.dina(n7613), .dinb(n7602), .dout(n7614));
  jor  g07357(.dina(n7614), .dinb(n199), .dout(n7615));
  jand g07358(.dina(n7614), .dinb(n199), .dout(n7616));
  jxor g07359(.dina(n7214), .dinb(n223), .dout(n7617));
  jor  g07360(.dina(n7617), .dinb(n7265), .dout(n7618));
  jxor g07361(.dina(n7618), .dinb(n7225), .dout(n7619));
  jor  g07362(.dina(n7619), .dinb(n7616), .dout(n7620));
  jand g07363(.dina(n7620), .dinb(n7615), .dout(n7621));
  jnot g07364(.din(n7230), .dout(n7622));
  jor  g07365(.dina(n7622), .dinb(n7228), .dout(n7623));
  jor  g07366(.dina(n7623), .dinb(n7265), .dout(n7624));
  jxor g07367(.dina(n7624), .dinb(n7239), .dout(n7625));
  jand g07368(.dina(asqrt[27] ), .dinb(n7253), .dout(n7626));
  jand g07369(.dina(n7626), .dinb(n7241), .dout(n7627));
  jor  g07370(.dina(n7627), .dinb(n7288), .dout(n7628));
  jor  g07371(.dina(n7628), .dinb(n7625), .dout(n7629));
  jor  g07372(.dina(n7629), .dinb(n7621), .dout(n7630));
  jand g07373(.dina(n7630), .dinb(n194), .dout(n7631));
  jand g07374(.dina(n7625), .dinb(n7621), .dout(n7632));
  jor  g07375(.dina(n7626), .dinb(n7241), .dout(n7633));
  jand g07376(.dina(n7253), .dinb(n7241), .dout(n7634));
  jor  g07377(.dina(n7634), .dinb(n194), .dout(n7635));
  jnot g07378(.din(n7635), .dout(n7636));
  jand g07379(.dina(n7636), .dinb(n7633), .dout(n7637));
  jor  g07380(.dina(n7637), .dinb(n7632), .dout(n7640));
  jor  g07381(.dina(n7640), .dinb(n7631), .dout(asqrt[26] ));
  jxor g07382(.dina(n7355), .dinb(n4494), .dout(n7642));
  jand g07383(.dina(n7642), .dinb(asqrt[26] ), .dout(n7643));
  jxor g07384(.dina(n7643), .dinb(n7269), .dout(n7644));
  jnot g07385(.din(n7644), .dout(n7645));
  jand g07386(.dina(asqrt[26] ), .dinb(a[52] ), .dout(n7646));
  jnot g07387(.din(a[50] ), .dout(n7647));
  jnot g07388(.din(a[51] ), .dout(n7648));
  jand g07389(.dina(n7271), .dinb(n7648), .dout(n7649));
  jand g07390(.dina(n7649), .dinb(n7647), .dout(n7650));
  jor  g07391(.dina(n7650), .dinb(n7646), .dout(n7651));
  jand g07392(.dina(n7651), .dinb(asqrt[27] ), .dout(n7652));
  jand g07393(.dina(asqrt[26] ), .dinb(n7271), .dout(n7653));
  jxor g07394(.dina(n7653), .dinb(n7272), .dout(n7654));
  jor  g07395(.dina(n7651), .dinb(asqrt[27] ), .dout(n7655));
  jand g07396(.dina(n7655), .dinb(n7654), .dout(n7656));
  jor  g07397(.dina(n7656), .dinb(n7652), .dout(n7657));
  jand g07398(.dina(n7657), .dinb(asqrt[28] ), .dout(n7658));
  jor  g07399(.dina(n7652), .dinb(asqrt[28] ), .dout(n7659));
  jor  g07400(.dina(n7659), .dinb(n7656), .dout(n7660));
  jand g07401(.dina(n7653), .dinb(n7272), .dout(n7661));
  jnot g07402(.din(n7631), .dout(n7662));
  jnot g07403(.din(n7632), .dout(n7663));
  jnot g07404(.din(n7637), .dout(n7664));
  jand g07405(.dina(n7664), .dinb(asqrt[27] ), .dout(n7665));
  jand g07406(.dina(n7665), .dinb(n7663), .dout(n7666));
  jand g07407(.dina(n7666), .dinb(n7662), .dout(n7667));
  jor  g07408(.dina(n7667), .dinb(n7661), .dout(n7668));
  jxor g07409(.dina(n7668), .dinb(n6872), .dout(n7669));
  jand g07410(.dina(n7669), .dinb(n7660), .dout(n7670));
  jor  g07411(.dina(n7670), .dinb(n7658), .dout(n7671));
  jand g07412(.dina(n7671), .dinb(asqrt[29] ), .dout(n7672));
  jor  g07413(.dina(n7671), .dinb(asqrt[29] ), .dout(n7673));
  jxor g07414(.dina(n7276), .dinb(n7260), .dout(n7674));
  jand g07415(.dina(n7674), .dinb(asqrt[26] ), .dout(n7675));
  jxor g07416(.dina(n7675), .dinb(n7279), .dout(n7676));
  jnot g07417(.din(n7676), .dout(n7677));
  jand g07418(.dina(n7677), .dinb(n7673), .dout(n7678));
  jor  g07419(.dina(n7678), .dinb(n7672), .dout(n7679));
  jand g07420(.dina(n7679), .dinb(asqrt[30] ), .dout(n7680));
  jnot g07421(.din(n7285), .dout(n7681));
  jand g07422(.dina(n7681), .dinb(n7283), .dout(n7682));
  jand g07423(.dina(n7682), .dinb(asqrt[26] ), .dout(n7683));
  jxor g07424(.dina(n7683), .dinb(n7293), .dout(n7684));
  jnot g07425(.din(n7684), .dout(n7685));
  jor  g07426(.dina(n7672), .dinb(asqrt[30] ), .dout(n7686));
  jor  g07427(.dina(n7686), .dinb(n7678), .dout(n7687));
  jand g07428(.dina(n7687), .dinb(n7685), .dout(n7688));
  jor  g07429(.dina(n7688), .dinb(n7680), .dout(n7689));
  jand g07430(.dina(n7689), .dinb(asqrt[31] ), .dout(n7690));
  jor  g07431(.dina(n7689), .dinb(asqrt[31] ), .dout(n7691));
  jnot g07432(.din(n7300), .dout(n7692));
  jxor g07433(.dina(n7295), .dinb(n6500), .dout(n7693));
  jand g07434(.dina(n7693), .dinb(asqrt[26] ), .dout(n7694));
  jxor g07435(.dina(n7694), .dinb(n7692), .dout(n7695));
  jand g07436(.dina(n7695), .dinb(n7691), .dout(n7696));
  jor  g07437(.dina(n7696), .dinb(n7690), .dout(n7697));
  jand g07438(.dina(n7697), .dinb(asqrt[32] ), .dout(n7698));
  jor  g07439(.dina(n7690), .dinb(asqrt[32] ), .dout(n7699));
  jor  g07440(.dina(n7699), .dinb(n7696), .dout(n7700));
  jnot g07441(.din(n7307), .dout(n7701));
  jnot g07442(.din(n7309), .dout(n7702));
  jand g07443(.dina(asqrt[26] ), .dinb(n7303), .dout(n7703));
  jand g07444(.dina(n7703), .dinb(n7702), .dout(n7704));
  jor  g07445(.dina(n7704), .dinb(n7701), .dout(n7705));
  jnot g07446(.din(n7310), .dout(n7706));
  jand g07447(.dina(n7703), .dinb(n7706), .dout(n7707));
  jnot g07448(.din(n7707), .dout(n7708));
  jand g07449(.dina(n7708), .dinb(n7705), .dout(n7709));
  jand g07450(.dina(n7709), .dinb(n7700), .dout(n7710));
  jor  g07451(.dina(n7710), .dinb(n7698), .dout(n7711));
  jand g07452(.dina(n7711), .dinb(asqrt[33] ), .dout(n7712));
  jor  g07453(.dina(n7711), .dinb(asqrt[33] ), .dout(n7713));
  jxor g07454(.dina(n7311), .dinb(n5788), .dout(n7714));
  jand g07455(.dina(n7714), .dinb(asqrt[26] ), .dout(n7715));
  jxor g07456(.dina(n7715), .dinb(n7316), .dout(n7716));
  jand g07457(.dina(n7716), .dinb(n7713), .dout(n7717));
  jor  g07458(.dina(n7717), .dinb(n7712), .dout(n7718));
  jand g07459(.dina(n7718), .dinb(asqrt[34] ), .dout(n7719));
  jnot g07460(.din(n7322), .dout(n7720));
  jand g07461(.dina(n7720), .dinb(n7320), .dout(n7721));
  jand g07462(.dina(n7721), .dinb(asqrt[26] ), .dout(n7722));
  jxor g07463(.dina(n7722), .dinb(n7331), .dout(n7723));
  jnot g07464(.din(n7723), .dout(n7724));
  jor  g07465(.dina(n7712), .dinb(asqrt[34] ), .dout(n7725));
  jor  g07466(.dina(n7725), .dinb(n7717), .dout(n7726));
  jand g07467(.dina(n7726), .dinb(n7724), .dout(n7727));
  jor  g07468(.dina(n7727), .dinb(n7719), .dout(n7728));
  jand g07469(.dina(n7728), .dinb(asqrt[35] ), .dout(n7729));
  jor  g07470(.dina(n7728), .dinb(asqrt[35] ), .dout(n7730));
  jxor g07471(.dina(n7333), .dinb(n5116), .dout(n7731));
  jand g07472(.dina(n7731), .dinb(asqrt[26] ), .dout(n7732));
  jxor g07473(.dina(n7732), .dinb(n7339), .dout(n7733));
  jand g07474(.dina(n7733), .dinb(n7730), .dout(n7734));
  jor  g07475(.dina(n7734), .dinb(n7729), .dout(n7735));
  jand g07476(.dina(n7735), .dinb(asqrt[36] ), .dout(n7736));
  jnot g07477(.din(n7345), .dout(n7737));
  jand g07478(.dina(n7737), .dinb(n7343), .dout(n7738));
  jand g07479(.dina(n7738), .dinb(asqrt[26] ), .dout(n7739));
  jxor g07480(.dina(n7739), .dinb(n7353), .dout(n7740));
  jnot g07481(.din(n7740), .dout(n7741));
  jor  g07482(.dina(n7729), .dinb(asqrt[36] ), .dout(n7742));
  jor  g07483(.dina(n7742), .dinb(n7734), .dout(n7743));
  jand g07484(.dina(n7743), .dinb(n7741), .dout(n7744));
  jor  g07485(.dina(n7744), .dinb(n7736), .dout(n7745));
  jand g07486(.dina(n7745), .dinb(asqrt[37] ), .dout(n7746));
  jor  g07487(.dina(n7745), .dinb(asqrt[37] ), .dout(n7747));
  jand g07488(.dina(n7747), .dinb(n7645), .dout(n7748));
  jor  g07489(.dina(n7748), .dinb(n7746), .dout(n7749));
  jand g07490(.dina(n7749), .dinb(asqrt[38] ), .dout(n7750));
  jor  g07491(.dina(n7746), .dinb(asqrt[38] ), .dout(n7751));
  jor  g07492(.dina(n7751), .dinb(n7748), .dout(n7752));
  jnot g07493(.din(n7364), .dout(n7753));
  jnot g07494(.din(n7366), .dout(n7754));
  jand g07495(.dina(asqrt[26] ), .dinb(n7360), .dout(n7755));
  jand g07496(.dina(n7755), .dinb(n7754), .dout(n7756));
  jor  g07497(.dina(n7756), .dinb(n7753), .dout(n7757));
  jnot g07498(.din(n7367), .dout(n7758));
  jand g07499(.dina(n7755), .dinb(n7758), .dout(n7759));
  jnot g07500(.din(n7759), .dout(n7760));
  jand g07501(.dina(n7760), .dinb(n7757), .dout(n7761));
  jand g07502(.dina(n7761), .dinb(n7752), .dout(n7762));
  jor  g07503(.dina(n7762), .dinb(n7750), .dout(n7763));
  jand g07504(.dina(n7763), .dinb(asqrt[39] ), .dout(n7764));
  jor  g07505(.dina(n7763), .dinb(asqrt[39] ), .dout(n7765));
  jnot g07506(.din(n7372), .dout(n7766));
  jnot g07507(.din(n7373), .dout(n7767));
  jand g07508(.dina(asqrt[26] ), .dinb(n7369), .dout(n7768));
  jand g07509(.dina(n7768), .dinb(n7767), .dout(n7769));
  jor  g07510(.dina(n7769), .dinb(n7766), .dout(n7770));
  jnot g07511(.din(n7374), .dout(n7771));
  jand g07512(.dina(n7768), .dinb(n7771), .dout(n7772));
  jnot g07513(.din(n7772), .dout(n7773));
  jand g07514(.dina(n7773), .dinb(n7770), .dout(n7774));
  jand g07515(.dina(n7774), .dinb(n7765), .dout(n7775));
  jor  g07516(.dina(n7775), .dinb(n7764), .dout(n7776));
  jand g07517(.dina(n7776), .dinb(asqrt[40] ), .dout(n7777));
  jor  g07518(.dina(n7764), .dinb(asqrt[40] ), .dout(n7778));
  jor  g07519(.dina(n7778), .dinb(n7775), .dout(n7779));
  jnot g07520(.din(n7380), .dout(n7780));
  jnot g07521(.din(n7382), .dout(n7781));
  jand g07522(.dina(asqrt[26] ), .dinb(n7376), .dout(n7782));
  jand g07523(.dina(n7782), .dinb(n7781), .dout(n7783));
  jor  g07524(.dina(n7783), .dinb(n7780), .dout(n7784));
  jnot g07525(.din(n7383), .dout(n7785));
  jand g07526(.dina(n7782), .dinb(n7785), .dout(n7786));
  jnot g07527(.din(n7786), .dout(n7787));
  jand g07528(.dina(n7787), .dinb(n7784), .dout(n7788));
  jand g07529(.dina(n7788), .dinb(n7779), .dout(n7789));
  jor  g07530(.dina(n7789), .dinb(n7777), .dout(n7790));
  jand g07531(.dina(n7790), .dinb(asqrt[41] ), .dout(n7791));
  jxor g07532(.dina(n7384), .dinb(n3371), .dout(n7792));
  jand g07533(.dina(n7792), .dinb(asqrt[26] ), .dout(n7793));
  jxor g07534(.dina(n7793), .dinb(n7394), .dout(n7794));
  jnot g07535(.din(n7794), .dout(n7795));
  jor  g07536(.dina(n7790), .dinb(asqrt[41] ), .dout(n7796));
  jand g07537(.dina(n7796), .dinb(n7795), .dout(n7797));
  jor  g07538(.dina(n7797), .dinb(n7791), .dout(n7798));
  jand g07539(.dina(n7798), .dinb(asqrt[42] ), .dout(n7799));
  jnot g07540(.din(n7399), .dout(n7800));
  jand g07541(.dina(n7800), .dinb(n7397), .dout(n7801));
  jand g07542(.dina(n7801), .dinb(asqrt[26] ), .dout(n7802));
  jxor g07543(.dina(n7802), .dinb(n7407), .dout(n7803));
  jnot g07544(.din(n7803), .dout(n7804));
  jor  g07545(.dina(n7791), .dinb(asqrt[42] ), .dout(n7805));
  jor  g07546(.dina(n7805), .dinb(n7797), .dout(n7806));
  jand g07547(.dina(n7806), .dinb(n7804), .dout(n7807));
  jor  g07548(.dina(n7807), .dinb(n7799), .dout(n7808));
  jand g07549(.dina(n7808), .dinb(asqrt[43] ), .dout(n7809));
  jor  g07550(.dina(n7808), .dinb(asqrt[43] ), .dout(n7810));
  jnot g07551(.din(n7413), .dout(n7811));
  jnot g07552(.din(n7414), .dout(n7812));
  jand g07553(.dina(asqrt[26] ), .dinb(n7410), .dout(n7813));
  jand g07554(.dina(n7813), .dinb(n7812), .dout(n7814));
  jor  g07555(.dina(n7814), .dinb(n7811), .dout(n7815));
  jnot g07556(.din(n7415), .dout(n7816));
  jand g07557(.dina(n7813), .dinb(n7816), .dout(n7817));
  jnot g07558(.din(n7817), .dout(n7818));
  jand g07559(.dina(n7818), .dinb(n7815), .dout(n7819));
  jand g07560(.dina(n7819), .dinb(n7810), .dout(n7820));
  jor  g07561(.dina(n7820), .dinb(n7809), .dout(n7821));
  jand g07562(.dina(n7821), .dinb(asqrt[44] ), .dout(n7822));
  jor  g07563(.dina(n7809), .dinb(asqrt[44] ), .dout(n7823));
  jor  g07564(.dina(n7823), .dinb(n7820), .dout(n7824));
  jnot g07565(.din(n7421), .dout(n7825));
  jnot g07566(.din(n7423), .dout(n7826));
  jand g07567(.dina(asqrt[26] ), .dinb(n7417), .dout(n7827));
  jand g07568(.dina(n7827), .dinb(n7826), .dout(n7828));
  jor  g07569(.dina(n7828), .dinb(n7825), .dout(n7829));
  jnot g07570(.din(n7424), .dout(n7830));
  jand g07571(.dina(n7827), .dinb(n7830), .dout(n7831));
  jnot g07572(.din(n7831), .dout(n7832));
  jand g07573(.dina(n7832), .dinb(n7829), .dout(n7833));
  jand g07574(.dina(n7833), .dinb(n7824), .dout(n7834));
  jor  g07575(.dina(n7834), .dinb(n7822), .dout(n7835));
  jand g07576(.dina(n7835), .dinb(asqrt[45] ), .dout(n7836));
  jxor g07577(.dina(n7425), .dinb(n2420), .dout(n7837));
  jand g07578(.dina(n7837), .dinb(asqrt[26] ), .dout(n7838));
  jxor g07579(.dina(n7838), .dinb(n7435), .dout(n7839));
  jnot g07580(.din(n7839), .dout(n7840));
  jor  g07581(.dina(n7835), .dinb(asqrt[45] ), .dout(n7841));
  jand g07582(.dina(n7841), .dinb(n7840), .dout(n7842));
  jor  g07583(.dina(n7842), .dinb(n7836), .dout(n7843));
  jand g07584(.dina(n7843), .dinb(asqrt[46] ), .dout(n7844));
  jnot g07585(.din(n7440), .dout(n7845));
  jand g07586(.dina(n7845), .dinb(n7438), .dout(n7846));
  jand g07587(.dina(n7846), .dinb(asqrt[26] ), .dout(n7847));
  jxor g07588(.dina(n7847), .dinb(n7448), .dout(n7848));
  jnot g07589(.din(n7848), .dout(n7849));
  jor  g07590(.dina(n7836), .dinb(asqrt[46] ), .dout(n7850));
  jor  g07591(.dina(n7850), .dinb(n7842), .dout(n7851));
  jand g07592(.dina(n7851), .dinb(n7849), .dout(n7852));
  jor  g07593(.dina(n7852), .dinb(n7844), .dout(n7853));
  jand g07594(.dina(n7853), .dinb(asqrt[47] ), .dout(n7854));
  jor  g07595(.dina(n7853), .dinb(asqrt[47] ), .dout(n7855));
  jnot g07596(.din(n7454), .dout(n7856));
  jnot g07597(.din(n7455), .dout(n7857));
  jand g07598(.dina(asqrt[26] ), .dinb(n7451), .dout(n7858));
  jand g07599(.dina(n7858), .dinb(n7857), .dout(n7859));
  jor  g07600(.dina(n7859), .dinb(n7856), .dout(n7860));
  jnot g07601(.din(n7456), .dout(n7861));
  jand g07602(.dina(n7858), .dinb(n7861), .dout(n7862));
  jnot g07603(.din(n7862), .dout(n7863));
  jand g07604(.dina(n7863), .dinb(n7860), .dout(n7864));
  jand g07605(.dina(n7864), .dinb(n7855), .dout(n7865));
  jor  g07606(.dina(n7865), .dinb(n7854), .dout(n7866));
  jand g07607(.dina(n7866), .dinb(asqrt[48] ), .dout(n7867));
  jor  g07608(.dina(n7854), .dinb(asqrt[48] ), .dout(n7868));
  jor  g07609(.dina(n7868), .dinb(n7865), .dout(n7869));
  jnot g07610(.din(n7462), .dout(n7870));
  jnot g07611(.din(n7464), .dout(n7871));
  jand g07612(.dina(asqrt[26] ), .dinb(n7458), .dout(n7872));
  jand g07613(.dina(n7872), .dinb(n7871), .dout(n7873));
  jor  g07614(.dina(n7873), .dinb(n7870), .dout(n7874));
  jnot g07615(.din(n7465), .dout(n7875));
  jand g07616(.dina(n7872), .dinb(n7875), .dout(n7876));
  jnot g07617(.din(n7876), .dout(n7877));
  jand g07618(.dina(n7877), .dinb(n7874), .dout(n7878));
  jand g07619(.dina(n7878), .dinb(n7869), .dout(n7879));
  jor  g07620(.dina(n7879), .dinb(n7867), .dout(n7880));
  jand g07621(.dina(n7880), .dinb(asqrt[49] ), .dout(n7881));
  jxor g07622(.dina(n7466), .dinb(n1641), .dout(n7882));
  jand g07623(.dina(n7882), .dinb(asqrt[26] ), .dout(n7883));
  jxor g07624(.dina(n7883), .dinb(n7476), .dout(n7884));
  jnot g07625(.din(n7884), .dout(n7885));
  jor  g07626(.dina(n7880), .dinb(asqrt[49] ), .dout(n7886));
  jand g07627(.dina(n7886), .dinb(n7885), .dout(n7887));
  jor  g07628(.dina(n7887), .dinb(n7881), .dout(n7888));
  jand g07629(.dina(n7888), .dinb(asqrt[50] ), .dout(n7889));
  jnot g07630(.din(n7481), .dout(n7890));
  jand g07631(.dina(n7890), .dinb(n7479), .dout(n7891));
  jand g07632(.dina(n7891), .dinb(asqrt[26] ), .dout(n7892));
  jxor g07633(.dina(n7892), .dinb(n7489), .dout(n7893));
  jnot g07634(.din(n7893), .dout(n7894));
  jor  g07635(.dina(n7881), .dinb(asqrt[50] ), .dout(n7895));
  jor  g07636(.dina(n7895), .dinb(n7887), .dout(n7896));
  jand g07637(.dina(n7896), .dinb(n7894), .dout(n7897));
  jor  g07638(.dina(n7897), .dinb(n7889), .dout(n7898));
  jand g07639(.dina(n7898), .dinb(asqrt[51] ), .dout(n7899));
  jor  g07640(.dina(n7898), .dinb(asqrt[51] ), .dout(n7900));
  jnot g07641(.din(n7495), .dout(n7901));
  jnot g07642(.din(n7496), .dout(n7902));
  jand g07643(.dina(asqrt[26] ), .dinb(n7492), .dout(n7903));
  jand g07644(.dina(n7903), .dinb(n7902), .dout(n7904));
  jor  g07645(.dina(n7904), .dinb(n7901), .dout(n7905));
  jnot g07646(.din(n7497), .dout(n7906));
  jand g07647(.dina(n7903), .dinb(n7906), .dout(n7907));
  jnot g07648(.din(n7907), .dout(n7908));
  jand g07649(.dina(n7908), .dinb(n7905), .dout(n7909));
  jand g07650(.dina(n7909), .dinb(n7900), .dout(n7910));
  jor  g07651(.dina(n7910), .dinb(n7899), .dout(n7911));
  jand g07652(.dina(n7911), .dinb(asqrt[52] ), .dout(n7912));
  jor  g07653(.dina(n7899), .dinb(asqrt[52] ), .dout(n7913));
  jor  g07654(.dina(n7913), .dinb(n7910), .dout(n7914));
  jnot g07655(.din(n7503), .dout(n7915));
  jnot g07656(.din(n7505), .dout(n7916));
  jand g07657(.dina(asqrt[26] ), .dinb(n7499), .dout(n7917));
  jand g07658(.dina(n7917), .dinb(n7916), .dout(n7918));
  jor  g07659(.dina(n7918), .dinb(n7915), .dout(n7919));
  jnot g07660(.din(n7506), .dout(n7920));
  jand g07661(.dina(n7917), .dinb(n7920), .dout(n7921));
  jnot g07662(.din(n7921), .dout(n7922));
  jand g07663(.dina(n7922), .dinb(n7919), .dout(n7923));
  jand g07664(.dina(n7923), .dinb(n7914), .dout(n7924));
  jor  g07665(.dina(n7924), .dinb(n7912), .dout(n7925));
  jand g07666(.dina(n7925), .dinb(asqrt[53] ), .dout(n7926));
  jxor g07667(.dina(n7507), .dinb(n1034), .dout(n7927));
  jand g07668(.dina(n7927), .dinb(asqrt[26] ), .dout(n7928));
  jxor g07669(.dina(n7928), .dinb(n7517), .dout(n7929));
  jnot g07670(.din(n7929), .dout(n7930));
  jor  g07671(.dina(n7925), .dinb(asqrt[53] ), .dout(n7931));
  jand g07672(.dina(n7931), .dinb(n7930), .dout(n7932));
  jor  g07673(.dina(n7932), .dinb(n7926), .dout(n7933));
  jand g07674(.dina(n7933), .dinb(asqrt[54] ), .dout(n7934));
  jnot g07675(.din(n7522), .dout(n7935));
  jand g07676(.dina(n7935), .dinb(n7520), .dout(n7936));
  jand g07677(.dina(n7936), .dinb(asqrt[26] ), .dout(n7937));
  jxor g07678(.dina(n7937), .dinb(n7530), .dout(n7938));
  jnot g07679(.din(n7938), .dout(n7939));
  jor  g07680(.dina(n7926), .dinb(asqrt[54] ), .dout(n7940));
  jor  g07681(.dina(n7940), .dinb(n7932), .dout(n7941));
  jand g07682(.dina(n7941), .dinb(n7939), .dout(n7942));
  jor  g07683(.dina(n7942), .dinb(n7934), .dout(n7943));
  jand g07684(.dina(n7943), .dinb(asqrt[55] ), .dout(n7944));
  jor  g07685(.dina(n7943), .dinb(asqrt[55] ), .dout(n7945));
  jnot g07686(.din(n7536), .dout(n7946));
  jnot g07687(.din(n7537), .dout(n7947));
  jand g07688(.dina(asqrt[26] ), .dinb(n7533), .dout(n7948));
  jand g07689(.dina(n7948), .dinb(n7947), .dout(n7949));
  jor  g07690(.dina(n7949), .dinb(n7946), .dout(n7950));
  jnot g07691(.din(n7538), .dout(n7951));
  jand g07692(.dina(n7948), .dinb(n7951), .dout(n7952));
  jnot g07693(.din(n7952), .dout(n7953));
  jand g07694(.dina(n7953), .dinb(n7950), .dout(n7954));
  jand g07695(.dina(n7954), .dinb(n7945), .dout(n7955));
  jor  g07696(.dina(n7955), .dinb(n7944), .dout(n7956));
  jand g07697(.dina(n7956), .dinb(asqrt[56] ), .dout(n7957));
  jor  g07698(.dina(n7944), .dinb(asqrt[56] ), .dout(n7958));
  jor  g07699(.dina(n7958), .dinb(n7955), .dout(n7959));
  jnot g07700(.din(n7544), .dout(n7960));
  jnot g07701(.din(n7546), .dout(n7961));
  jand g07702(.dina(asqrt[26] ), .dinb(n7540), .dout(n7962));
  jand g07703(.dina(n7962), .dinb(n7961), .dout(n7963));
  jor  g07704(.dina(n7963), .dinb(n7960), .dout(n7964));
  jnot g07705(.din(n7547), .dout(n7965));
  jand g07706(.dina(n7962), .dinb(n7965), .dout(n7966));
  jnot g07707(.din(n7966), .dout(n7967));
  jand g07708(.dina(n7967), .dinb(n7964), .dout(n7968));
  jand g07709(.dina(n7968), .dinb(n7959), .dout(n7969));
  jor  g07710(.dina(n7969), .dinb(n7957), .dout(n7970));
  jand g07711(.dina(n7970), .dinb(asqrt[57] ), .dout(n7971));
  jxor g07712(.dina(n7548), .dinb(n590), .dout(n7972));
  jand g07713(.dina(n7972), .dinb(asqrt[26] ), .dout(n7973));
  jxor g07714(.dina(n7973), .dinb(n7558), .dout(n7974));
  jnot g07715(.din(n7974), .dout(n7975));
  jor  g07716(.dina(n7970), .dinb(asqrt[57] ), .dout(n7976));
  jand g07717(.dina(n7976), .dinb(n7975), .dout(n7977));
  jor  g07718(.dina(n7977), .dinb(n7971), .dout(n7978));
  jand g07719(.dina(n7978), .dinb(asqrt[58] ), .dout(n7979));
  jnot g07720(.din(n7563), .dout(n7980));
  jand g07721(.dina(n7980), .dinb(n7561), .dout(n7981));
  jand g07722(.dina(n7981), .dinb(asqrt[26] ), .dout(n7982));
  jxor g07723(.dina(n7982), .dinb(n7571), .dout(n7983));
  jnot g07724(.din(n7983), .dout(n7984));
  jor  g07725(.dina(n7971), .dinb(asqrt[58] ), .dout(n7985));
  jor  g07726(.dina(n7985), .dinb(n7977), .dout(n7986));
  jand g07727(.dina(n7986), .dinb(n7984), .dout(n7987));
  jor  g07728(.dina(n7987), .dinb(n7979), .dout(n7988));
  jand g07729(.dina(n7988), .dinb(asqrt[59] ), .dout(n7989));
  jor  g07730(.dina(n7988), .dinb(asqrt[59] ), .dout(n7990));
  jnot g07731(.din(n7577), .dout(n7991));
  jnot g07732(.din(n7578), .dout(n7992));
  jand g07733(.dina(asqrt[26] ), .dinb(n7574), .dout(n7993));
  jand g07734(.dina(n7993), .dinb(n7992), .dout(n7994));
  jor  g07735(.dina(n7994), .dinb(n7991), .dout(n7995));
  jnot g07736(.din(n7579), .dout(n7996));
  jand g07737(.dina(n7993), .dinb(n7996), .dout(n7997));
  jnot g07738(.din(n7997), .dout(n7998));
  jand g07739(.dina(n7998), .dinb(n7995), .dout(n7999));
  jand g07740(.dina(n7999), .dinb(n7990), .dout(n8000));
  jor  g07741(.dina(n8000), .dinb(n7989), .dout(n8001));
  jand g07742(.dina(n8001), .dinb(asqrt[60] ), .dout(n8002));
  jor  g07743(.dina(n7989), .dinb(asqrt[60] ), .dout(n8003));
  jor  g07744(.dina(n8003), .dinb(n8000), .dout(n8004));
  jnot g07745(.din(n7585), .dout(n8005));
  jnot g07746(.din(n7587), .dout(n8006));
  jand g07747(.dina(asqrt[26] ), .dinb(n7581), .dout(n8007));
  jand g07748(.dina(n8007), .dinb(n8006), .dout(n8008));
  jor  g07749(.dina(n8008), .dinb(n8005), .dout(n8009));
  jnot g07750(.din(n7588), .dout(n8010));
  jand g07751(.dina(n8007), .dinb(n8010), .dout(n8011));
  jnot g07752(.din(n8011), .dout(n8012));
  jand g07753(.dina(n8012), .dinb(n8009), .dout(n8013));
  jand g07754(.dina(n8013), .dinb(n8004), .dout(n8014));
  jor  g07755(.dina(n8014), .dinb(n8002), .dout(n8015));
  jand g07756(.dina(n8015), .dinb(asqrt[61] ), .dout(n8016));
  jxor g07757(.dina(n7589), .dinb(n290), .dout(n8017));
  jand g07758(.dina(n8017), .dinb(asqrt[26] ), .dout(n8018));
  jxor g07759(.dina(n8018), .dinb(n7599), .dout(n8019));
  jnot g07760(.din(n8019), .dout(n8020));
  jor  g07761(.dina(n8015), .dinb(asqrt[61] ), .dout(n8021));
  jand g07762(.dina(n8021), .dinb(n8020), .dout(n8022));
  jor  g07763(.dina(n8022), .dinb(n8016), .dout(n8023));
  jand g07764(.dina(n8023), .dinb(asqrt[62] ), .dout(n8024));
  jnot g07765(.din(n7604), .dout(n8025));
  jand g07766(.dina(n8025), .dinb(n7602), .dout(n8026));
  jand g07767(.dina(n8026), .dinb(asqrt[26] ), .dout(n8027));
  jxor g07768(.dina(n8027), .dinb(n7612), .dout(n8028));
  jnot g07769(.din(n8028), .dout(n8029));
  jor  g07770(.dina(n8016), .dinb(asqrt[62] ), .dout(n8030));
  jor  g07771(.dina(n8030), .dinb(n8022), .dout(n8031));
  jand g07772(.dina(n8031), .dinb(n8029), .dout(n8032));
  jor  g07773(.dina(n8032), .dinb(n8024), .dout(n8033));
  jxor g07774(.dina(n7614), .dinb(n199), .dout(n8034));
  jand g07775(.dina(n8034), .dinb(asqrt[26] ), .dout(n8035));
  jxor g07776(.dina(n8035), .dinb(n7619), .dout(n8036));
  jnot g07777(.din(n7621), .dout(n8037));
  jnot g07778(.din(n7625), .dout(n8038));
  jand g07779(.dina(asqrt[26] ), .dinb(n8038), .dout(n8039));
  jand g07780(.dina(n8039), .dinb(n8037), .dout(n8040));
  jor  g07781(.dina(n8040), .dinb(n7632), .dout(n8041));
  jor  g07782(.dina(n8041), .dinb(n8036), .dout(n8042));
  jnot g07783(.din(n8042), .dout(n8043));
  jand g07784(.dina(n8043), .dinb(n8033), .dout(n8044));
  jor  g07785(.dina(n8044), .dinb(asqrt[63] ), .dout(n8045));
  jnot g07786(.din(n8036), .dout(n8046));
  jor  g07787(.dina(n8046), .dinb(n8033), .dout(n8047));
  jor  g07788(.dina(n8039), .dinb(n8037), .dout(n8048));
  jand g07789(.dina(n8038), .dinb(n8037), .dout(n8049));
  jor  g07790(.dina(n8049), .dinb(n194), .dout(n8050));
  jnot g07791(.din(n8050), .dout(n8051));
  jand g07792(.dina(n8051), .dinb(n8048), .dout(n8052));
  jnot g07793(.din(asqrt[26] ), .dout(n8053));
  jnot g07794(.din(n8052), .dout(n8056));
  jand g07795(.dina(n8056), .dinb(n8047), .dout(n8057));
  jand g07796(.dina(n8057), .dinb(n8045), .dout(n8058));
  jxor g07797(.dina(n7745), .dinb(n3912), .dout(n8059));
  jor  g07798(.dina(n8059), .dinb(n8058), .dout(n8060));
  jxor g07799(.dina(n8060), .dinb(n7645), .dout(n8061));
  jor  g07800(.dina(n8058), .dinb(n7647), .dout(n8062));
  jnot g07801(.din(a[48] ), .dout(n8063));
  jnot g07802(.din(a[49] ), .dout(n8064));
  jand g07803(.dina(n7647), .dinb(n8064), .dout(n8065));
  jand g07804(.dina(n8065), .dinb(n8063), .dout(n8066));
  jnot g07805(.din(n8066), .dout(n8067));
  jand g07806(.dina(n8067), .dinb(n8062), .dout(n8068));
  jor  g07807(.dina(n8068), .dinb(n8053), .dout(n8069));
  jor  g07808(.dina(n8058), .dinb(a[50] ), .dout(n8070));
  jxor g07809(.dina(n8070), .dinb(n7648), .dout(n8071));
  jand g07810(.dina(n8068), .dinb(n8053), .dout(n8072));
  jor  g07811(.dina(n8072), .dinb(n8071), .dout(n8073));
  jand g07812(.dina(n8073), .dinb(n8069), .dout(n8074));
  jor  g07813(.dina(n8074), .dinb(n7265), .dout(n8075));
  jand g07814(.dina(n8069), .dinb(n7265), .dout(n8076));
  jand g07815(.dina(n8076), .dinb(n8073), .dout(n8077));
  jor  g07816(.dina(n8070), .dinb(a[51] ), .dout(n8078));
  jnot g07817(.din(n8045), .dout(n8079));
  jnot g07818(.din(n8047), .dout(n8080));
  jor  g07819(.dina(n8052), .dinb(n8053), .dout(n8081));
  jor  g07820(.dina(n8081), .dinb(n8080), .dout(n8082));
  jor  g07821(.dina(n8082), .dinb(n8079), .dout(n8083));
  jand g07822(.dina(n8083), .dinb(n8078), .dout(n8084));
  jxor g07823(.dina(n8084), .dinb(n7271), .dout(n8085));
  jor  g07824(.dina(n8085), .dinb(n8077), .dout(n8086));
  jand g07825(.dina(n8086), .dinb(n8075), .dout(n8087));
  jor  g07826(.dina(n8087), .dinb(n7260), .dout(n8088));
  jand g07827(.dina(n8087), .dinb(n7260), .dout(n8089));
  jxor g07828(.dina(n7651), .dinb(n7265), .dout(n8090));
  jor  g07829(.dina(n8090), .dinb(n8058), .dout(n8091));
  jxor g07830(.dina(n8091), .dinb(n7654), .dout(n8092));
  jor  g07831(.dina(n8092), .dinb(n8089), .dout(n8093));
  jand g07832(.dina(n8093), .dinb(n8088), .dout(n8094));
  jor  g07833(.dina(n8094), .dinb(n6505), .dout(n8095));
  jnot g07834(.din(n7660), .dout(n8096));
  jor  g07835(.dina(n8096), .dinb(n7658), .dout(n8097));
  jor  g07836(.dina(n8097), .dinb(n8058), .dout(n8098));
  jxor g07837(.dina(n8098), .dinb(n7669), .dout(n8099));
  jand g07838(.dina(n8088), .dinb(n6505), .dout(n8100));
  jand g07839(.dina(n8100), .dinb(n8093), .dout(n8101));
  jor  g07840(.dina(n8101), .dinb(n8099), .dout(n8102));
  jand g07841(.dina(n8102), .dinb(n8095), .dout(n8103));
  jor  g07842(.dina(n8103), .dinb(n6500), .dout(n8104));
  jand g07843(.dina(n8103), .dinb(n6500), .dout(n8105));
  jxor g07844(.dina(n7671), .dinb(n6505), .dout(n8106));
  jor  g07845(.dina(n8106), .dinb(n8058), .dout(n8107));
  jxor g07846(.dina(n8107), .dinb(n7676), .dout(n8108));
  jnot g07847(.din(n8108), .dout(n8109));
  jor  g07848(.dina(n8109), .dinb(n8105), .dout(n8110));
  jand g07849(.dina(n8110), .dinb(n8104), .dout(n8111));
  jor  g07850(.dina(n8111), .dinb(n5793), .dout(n8112));
  jand g07851(.dina(n8104), .dinb(n5793), .dout(n8113));
  jand g07852(.dina(n8113), .dinb(n8110), .dout(n8114));
  jnot g07853(.din(n7680), .dout(n8115));
  jnot g07854(.din(n8058), .dout(asqrt[25] ));
  jand g07855(.dina(asqrt[25] ), .dinb(n8115), .dout(n8117));
  jand g07856(.dina(n8117), .dinb(n7687), .dout(n8118));
  jor  g07857(.dina(n8118), .dinb(n7685), .dout(n8119));
  jand g07858(.dina(n8117), .dinb(n7688), .dout(n8120));
  jnot g07859(.din(n8120), .dout(n8121));
  jand g07860(.dina(n8121), .dinb(n8119), .dout(n8122));
  jnot g07861(.din(n8122), .dout(n8123));
  jor  g07862(.dina(n8123), .dinb(n8114), .dout(n8124));
  jand g07863(.dina(n8124), .dinb(n8112), .dout(n8125));
  jor  g07864(.dina(n8125), .dinb(n5788), .dout(n8126));
  jand g07865(.dina(n8125), .dinb(n5788), .dout(n8127));
  jnot g07866(.din(n7695), .dout(n8128));
  jxor g07867(.dina(n7689), .dinb(n5793), .dout(n8129));
  jor  g07868(.dina(n8129), .dinb(n8058), .dout(n8130));
  jxor g07869(.dina(n8130), .dinb(n8128), .dout(n8131));
  jnot g07870(.din(n8131), .dout(n8132));
  jor  g07871(.dina(n8132), .dinb(n8127), .dout(n8133));
  jand g07872(.dina(n8133), .dinb(n8126), .dout(n8134));
  jor  g07873(.dina(n8134), .dinb(n5121), .dout(n8135));
  jnot g07874(.din(n7700), .dout(n8136));
  jor  g07875(.dina(n8136), .dinb(n7698), .dout(n8137));
  jor  g07876(.dina(n8137), .dinb(n8058), .dout(n8138));
  jxor g07877(.dina(n8138), .dinb(n7709), .dout(n8139));
  jand g07878(.dina(n8126), .dinb(n5121), .dout(n8140));
  jand g07879(.dina(n8140), .dinb(n8133), .dout(n8141));
  jor  g07880(.dina(n8141), .dinb(n8139), .dout(n8142));
  jand g07881(.dina(n8142), .dinb(n8135), .dout(n8143));
  jor  g07882(.dina(n8143), .dinb(n5116), .dout(n8144));
  jand g07883(.dina(n8143), .dinb(n5116), .dout(n8145));
  jnot g07884(.din(n7716), .dout(n8146));
  jxor g07885(.dina(n7711), .dinb(n5121), .dout(n8147));
  jor  g07886(.dina(n8147), .dinb(n8058), .dout(n8148));
  jxor g07887(.dina(n8148), .dinb(n8146), .dout(n8149));
  jnot g07888(.din(n8149), .dout(n8150));
  jor  g07889(.dina(n8150), .dinb(n8145), .dout(n8151));
  jand g07890(.dina(n8151), .dinb(n8144), .dout(n8152));
  jor  g07891(.dina(n8152), .dinb(n4499), .dout(n8153));
  jand g07892(.dina(n8144), .dinb(n4499), .dout(n8154));
  jand g07893(.dina(n8154), .dinb(n8151), .dout(n8155));
  jnot g07894(.din(n7719), .dout(n8156));
  jand g07895(.dina(asqrt[25] ), .dinb(n8156), .dout(n8157));
  jand g07896(.dina(n8157), .dinb(n7726), .dout(n8158));
  jor  g07897(.dina(n8158), .dinb(n7724), .dout(n8159));
  jand g07898(.dina(n8157), .dinb(n7727), .dout(n8160));
  jnot g07899(.din(n8160), .dout(n8161));
  jand g07900(.dina(n8161), .dinb(n8159), .dout(n8162));
  jnot g07901(.din(n8162), .dout(n8163));
  jor  g07902(.dina(n8163), .dinb(n8155), .dout(n8164));
  jand g07903(.dina(n8164), .dinb(n8153), .dout(n8165));
  jor  g07904(.dina(n8165), .dinb(n4494), .dout(n8166));
  jxor g07905(.dina(n7728), .dinb(n4499), .dout(n8167));
  jor  g07906(.dina(n8167), .dinb(n8058), .dout(n8168));
  jxor g07907(.dina(n8168), .dinb(n7733), .dout(n8169));
  jand g07908(.dina(n8165), .dinb(n4494), .dout(n8170));
  jor  g07909(.dina(n8170), .dinb(n8169), .dout(n8171));
  jand g07910(.dina(n8171), .dinb(n8166), .dout(n8172));
  jor  g07911(.dina(n8172), .dinb(n3912), .dout(n8173));
  jand g07912(.dina(n8166), .dinb(n3912), .dout(n8174));
  jand g07913(.dina(n8174), .dinb(n8171), .dout(n8175));
  jnot g07914(.din(n7736), .dout(n8176));
  jand g07915(.dina(asqrt[25] ), .dinb(n8176), .dout(n8177));
  jand g07916(.dina(n8177), .dinb(n7743), .dout(n8178));
  jor  g07917(.dina(n8178), .dinb(n7741), .dout(n8179));
  jand g07918(.dina(n8177), .dinb(n7744), .dout(n8180));
  jnot g07919(.din(n8180), .dout(n8181));
  jand g07920(.dina(n8181), .dinb(n8179), .dout(n8182));
  jnot g07921(.din(n8182), .dout(n8183));
  jor  g07922(.dina(n8183), .dinb(n8175), .dout(n8184));
  jand g07923(.dina(n8184), .dinb(n8173), .dout(n8185));
  jor  g07924(.dina(n8185), .dinb(n3907), .dout(n8186));
  jand g07925(.dina(n8185), .dinb(n3907), .dout(n8187));
  jor  g07926(.dina(n8187), .dinb(n8061), .dout(n8188));
  jand g07927(.dina(n8188), .dinb(n8186), .dout(n8189));
  jor  g07928(.dina(n8189), .dinb(n3376), .dout(n8190));
  jnot g07929(.din(n7752), .dout(n8191));
  jor  g07930(.dina(n8191), .dinb(n7750), .dout(n8192));
  jor  g07931(.dina(n8192), .dinb(n8058), .dout(n8193));
  jxor g07932(.dina(n8193), .dinb(n7761), .dout(n8194));
  jand g07933(.dina(n8186), .dinb(n3376), .dout(n8195));
  jand g07934(.dina(n8195), .dinb(n8188), .dout(n8196));
  jor  g07935(.dina(n8196), .dinb(n8194), .dout(n8197));
  jand g07936(.dina(n8197), .dinb(n8190), .dout(n8198));
  jor  g07937(.dina(n8198), .dinb(n3371), .dout(n8199));
  jxor g07938(.dina(n7763), .dinb(n3376), .dout(n8200));
  jor  g07939(.dina(n8200), .dinb(n8058), .dout(n8201));
  jxor g07940(.dina(n8201), .dinb(n7774), .dout(n8202));
  jand g07941(.dina(n8198), .dinb(n3371), .dout(n8203));
  jor  g07942(.dina(n8203), .dinb(n8202), .dout(n8204));
  jand g07943(.dina(n8204), .dinb(n8199), .dout(n8205));
  jor  g07944(.dina(n8205), .dinb(n2875), .dout(n8206));
  jnot g07945(.din(n7779), .dout(n8207));
  jor  g07946(.dina(n8207), .dinb(n7777), .dout(n8208));
  jor  g07947(.dina(n8208), .dinb(n8058), .dout(n8209));
  jxor g07948(.dina(n8209), .dinb(n7788), .dout(n8210));
  jand g07949(.dina(n8199), .dinb(n2875), .dout(n8211));
  jand g07950(.dina(n8211), .dinb(n8204), .dout(n8212));
  jor  g07951(.dina(n8212), .dinb(n8210), .dout(n8213));
  jand g07952(.dina(n8213), .dinb(n8206), .dout(n8214));
  jor  g07953(.dina(n8214), .dinb(n2870), .dout(n8215));
  jand g07954(.dina(n8214), .dinb(n2870), .dout(n8216));
  jnot g07955(.din(n7791), .dout(n8217));
  jand g07956(.dina(asqrt[25] ), .dinb(n8217), .dout(n8218));
  jand g07957(.dina(n8218), .dinb(n7796), .dout(n8219));
  jor  g07958(.dina(n8219), .dinb(n7795), .dout(n8220));
  jand g07959(.dina(n8218), .dinb(n7797), .dout(n8221));
  jnot g07960(.din(n8221), .dout(n8222));
  jand g07961(.dina(n8222), .dinb(n8220), .dout(n8223));
  jnot g07962(.din(n8223), .dout(n8224));
  jor  g07963(.dina(n8224), .dinb(n8216), .dout(n8225));
  jand g07964(.dina(n8225), .dinb(n8215), .dout(n8226));
  jor  g07965(.dina(n8226), .dinb(n2425), .dout(n8227));
  jand g07966(.dina(n8215), .dinb(n2425), .dout(n8228));
  jand g07967(.dina(n8228), .dinb(n8225), .dout(n8229));
  jnot g07968(.din(n7799), .dout(n8230));
  jand g07969(.dina(asqrt[25] ), .dinb(n8230), .dout(n8231));
  jand g07970(.dina(n8231), .dinb(n7806), .dout(n8232));
  jor  g07971(.dina(n8232), .dinb(n7804), .dout(n8233));
  jand g07972(.dina(n8231), .dinb(n7807), .dout(n8234));
  jnot g07973(.din(n8234), .dout(n8235));
  jand g07974(.dina(n8235), .dinb(n8233), .dout(n8236));
  jnot g07975(.din(n8236), .dout(n8237));
  jor  g07976(.dina(n8237), .dinb(n8229), .dout(n8238));
  jand g07977(.dina(n8238), .dinb(n8227), .dout(n8239));
  jor  g07978(.dina(n8239), .dinb(n2420), .dout(n8240));
  jxor g07979(.dina(n7808), .dinb(n2425), .dout(n8241));
  jor  g07980(.dina(n8241), .dinb(n8058), .dout(n8242));
  jxor g07981(.dina(n8242), .dinb(n7819), .dout(n8243));
  jand g07982(.dina(n8239), .dinb(n2420), .dout(n8244));
  jor  g07983(.dina(n8244), .dinb(n8243), .dout(n8245));
  jand g07984(.dina(n8245), .dinb(n8240), .dout(n8246));
  jor  g07985(.dina(n8246), .dinb(n2010), .dout(n8247));
  jnot g07986(.din(n7824), .dout(n8248));
  jor  g07987(.dina(n8248), .dinb(n7822), .dout(n8249));
  jor  g07988(.dina(n8249), .dinb(n8058), .dout(n8250));
  jxor g07989(.dina(n8250), .dinb(n7833), .dout(n8251));
  jand g07990(.dina(n8240), .dinb(n2010), .dout(n8252));
  jand g07991(.dina(n8252), .dinb(n8245), .dout(n8253));
  jor  g07992(.dina(n8253), .dinb(n8251), .dout(n8254));
  jand g07993(.dina(n8254), .dinb(n8247), .dout(n8255));
  jor  g07994(.dina(n8255), .dinb(n2005), .dout(n8256));
  jand g07995(.dina(n8255), .dinb(n2005), .dout(n8257));
  jnot g07996(.din(n7836), .dout(n8258));
  jand g07997(.dina(asqrt[25] ), .dinb(n8258), .dout(n8259));
  jand g07998(.dina(n8259), .dinb(n7841), .dout(n8260));
  jor  g07999(.dina(n8260), .dinb(n7840), .dout(n8261));
  jand g08000(.dina(n8259), .dinb(n7842), .dout(n8262));
  jnot g08001(.din(n8262), .dout(n8263));
  jand g08002(.dina(n8263), .dinb(n8261), .dout(n8264));
  jnot g08003(.din(n8264), .dout(n8265));
  jor  g08004(.dina(n8265), .dinb(n8257), .dout(n8266));
  jand g08005(.dina(n8266), .dinb(n8256), .dout(n8267));
  jor  g08006(.dina(n8267), .dinb(n1646), .dout(n8268));
  jand g08007(.dina(n8256), .dinb(n1646), .dout(n8269));
  jand g08008(.dina(n8269), .dinb(n8266), .dout(n8270));
  jnot g08009(.din(n7844), .dout(n8271));
  jand g08010(.dina(asqrt[25] ), .dinb(n8271), .dout(n8272));
  jand g08011(.dina(n8272), .dinb(n7851), .dout(n8273));
  jor  g08012(.dina(n8273), .dinb(n7849), .dout(n8274));
  jand g08013(.dina(n8272), .dinb(n7852), .dout(n8275));
  jnot g08014(.din(n8275), .dout(n8276));
  jand g08015(.dina(n8276), .dinb(n8274), .dout(n8277));
  jnot g08016(.din(n8277), .dout(n8278));
  jor  g08017(.dina(n8278), .dinb(n8270), .dout(n8279));
  jand g08018(.dina(n8279), .dinb(n8268), .dout(n8280));
  jor  g08019(.dina(n8280), .dinb(n1641), .dout(n8281));
  jxor g08020(.dina(n7853), .dinb(n1646), .dout(n8282));
  jor  g08021(.dina(n8282), .dinb(n8058), .dout(n8283));
  jxor g08022(.dina(n8283), .dinb(n7864), .dout(n8284));
  jand g08023(.dina(n8280), .dinb(n1641), .dout(n8285));
  jor  g08024(.dina(n8285), .dinb(n8284), .dout(n8286));
  jand g08025(.dina(n8286), .dinb(n8281), .dout(n8287));
  jor  g08026(.dina(n8287), .dinb(n1317), .dout(n8288));
  jnot g08027(.din(n7869), .dout(n8289));
  jor  g08028(.dina(n8289), .dinb(n7867), .dout(n8290));
  jor  g08029(.dina(n8290), .dinb(n8058), .dout(n8291));
  jxor g08030(.dina(n8291), .dinb(n7878), .dout(n8292));
  jand g08031(.dina(n8281), .dinb(n1317), .dout(n8293));
  jand g08032(.dina(n8293), .dinb(n8286), .dout(n8294));
  jor  g08033(.dina(n8294), .dinb(n8292), .dout(n8295));
  jand g08034(.dina(n8295), .dinb(n8288), .dout(n8296));
  jor  g08035(.dina(n8296), .dinb(n1312), .dout(n8297));
  jand g08036(.dina(n8296), .dinb(n1312), .dout(n8298));
  jnot g08037(.din(n7881), .dout(n8299));
  jand g08038(.dina(asqrt[25] ), .dinb(n8299), .dout(n8300));
  jand g08039(.dina(n8300), .dinb(n7886), .dout(n8301));
  jor  g08040(.dina(n8301), .dinb(n7885), .dout(n8302));
  jand g08041(.dina(n8300), .dinb(n7887), .dout(n8303));
  jnot g08042(.din(n8303), .dout(n8304));
  jand g08043(.dina(n8304), .dinb(n8302), .dout(n8305));
  jnot g08044(.din(n8305), .dout(n8306));
  jor  g08045(.dina(n8306), .dinb(n8298), .dout(n8307));
  jand g08046(.dina(n8307), .dinb(n8297), .dout(n8308));
  jor  g08047(.dina(n8308), .dinb(n1039), .dout(n8309));
  jand g08048(.dina(n8297), .dinb(n1039), .dout(n8310));
  jand g08049(.dina(n8310), .dinb(n8307), .dout(n8311));
  jnot g08050(.din(n7889), .dout(n8312));
  jand g08051(.dina(asqrt[25] ), .dinb(n8312), .dout(n8313));
  jand g08052(.dina(n8313), .dinb(n7896), .dout(n8314));
  jor  g08053(.dina(n8314), .dinb(n7894), .dout(n8315));
  jand g08054(.dina(n8313), .dinb(n7897), .dout(n8316));
  jnot g08055(.din(n8316), .dout(n8317));
  jand g08056(.dina(n8317), .dinb(n8315), .dout(n8318));
  jnot g08057(.din(n8318), .dout(n8319));
  jor  g08058(.dina(n8319), .dinb(n8311), .dout(n8320));
  jand g08059(.dina(n8320), .dinb(n8309), .dout(n8321));
  jor  g08060(.dina(n8321), .dinb(n1034), .dout(n8322));
  jxor g08061(.dina(n7898), .dinb(n1039), .dout(n8323));
  jor  g08062(.dina(n8323), .dinb(n8058), .dout(n8324));
  jxor g08063(.dina(n8324), .dinb(n7909), .dout(n8325));
  jand g08064(.dina(n8321), .dinb(n1034), .dout(n8326));
  jor  g08065(.dina(n8326), .dinb(n8325), .dout(n8327));
  jand g08066(.dina(n8327), .dinb(n8322), .dout(n8328));
  jor  g08067(.dina(n8328), .dinb(n796), .dout(n8329));
  jnot g08068(.din(n7914), .dout(n8330));
  jor  g08069(.dina(n8330), .dinb(n7912), .dout(n8331));
  jor  g08070(.dina(n8331), .dinb(n8058), .dout(n8332));
  jxor g08071(.dina(n8332), .dinb(n7923), .dout(n8333));
  jand g08072(.dina(n8322), .dinb(n796), .dout(n8334));
  jand g08073(.dina(n8334), .dinb(n8327), .dout(n8335));
  jor  g08074(.dina(n8335), .dinb(n8333), .dout(n8336));
  jand g08075(.dina(n8336), .dinb(n8329), .dout(n8337));
  jor  g08076(.dina(n8337), .dinb(n791), .dout(n8338));
  jand g08077(.dina(n8337), .dinb(n791), .dout(n8339));
  jnot g08078(.din(n7926), .dout(n8340));
  jand g08079(.dina(asqrt[25] ), .dinb(n8340), .dout(n8341));
  jand g08080(.dina(n8341), .dinb(n7931), .dout(n8342));
  jor  g08081(.dina(n8342), .dinb(n7930), .dout(n8343));
  jand g08082(.dina(n8341), .dinb(n7932), .dout(n8344));
  jnot g08083(.din(n8344), .dout(n8345));
  jand g08084(.dina(n8345), .dinb(n8343), .dout(n8346));
  jnot g08085(.din(n8346), .dout(n8347));
  jor  g08086(.dina(n8347), .dinb(n8339), .dout(n8348));
  jand g08087(.dina(n8348), .dinb(n8338), .dout(n8349));
  jor  g08088(.dina(n8349), .dinb(n595), .dout(n8350));
  jand g08089(.dina(n8338), .dinb(n595), .dout(n8351));
  jand g08090(.dina(n8351), .dinb(n8348), .dout(n8352));
  jnot g08091(.din(n7934), .dout(n8353));
  jand g08092(.dina(asqrt[25] ), .dinb(n8353), .dout(n8354));
  jand g08093(.dina(n8354), .dinb(n7941), .dout(n8355));
  jor  g08094(.dina(n8355), .dinb(n7939), .dout(n8356));
  jand g08095(.dina(n8354), .dinb(n7942), .dout(n8357));
  jnot g08096(.din(n8357), .dout(n8358));
  jand g08097(.dina(n8358), .dinb(n8356), .dout(n8359));
  jnot g08098(.din(n8359), .dout(n8360));
  jor  g08099(.dina(n8360), .dinb(n8352), .dout(n8361));
  jand g08100(.dina(n8361), .dinb(n8350), .dout(n8362));
  jor  g08101(.dina(n8362), .dinb(n590), .dout(n8363));
  jxor g08102(.dina(n7943), .dinb(n595), .dout(n8364));
  jor  g08103(.dina(n8364), .dinb(n8058), .dout(n8365));
  jxor g08104(.dina(n8365), .dinb(n7954), .dout(n8366));
  jand g08105(.dina(n8362), .dinb(n590), .dout(n8367));
  jor  g08106(.dina(n8367), .dinb(n8366), .dout(n8368));
  jand g08107(.dina(n8368), .dinb(n8363), .dout(n8369));
  jor  g08108(.dina(n8369), .dinb(n430), .dout(n8370));
  jnot g08109(.din(n7959), .dout(n8371));
  jor  g08110(.dina(n8371), .dinb(n7957), .dout(n8372));
  jor  g08111(.dina(n8372), .dinb(n8058), .dout(n8373));
  jxor g08112(.dina(n8373), .dinb(n7968), .dout(n8374));
  jand g08113(.dina(n8363), .dinb(n430), .dout(n8375));
  jand g08114(.dina(n8375), .dinb(n8368), .dout(n8376));
  jor  g08115(.dina(n8376), .dinb(n8374), .dout(n8377));
  jand g08116(.dina(n8377), .dinb(n8370), .dout(n8378));
  jor  g08117(.dina(n8378), .dinb(n425), .dout(n8379));
  jand g08118(.dina(n8378), .dinb(n425), .dout(n8380));
  jnot g08119(.din(n7971), .dout(n8381));
  jand g08120(.dina(asqrt[25] ), .dinb(n8381), .dout(n8382));
  jand g08121(.dina(n8382), .dinb(n7976), .dout(n8383));
  jor  g08122(.dina(n8383), .dinb(n7975), .dout(n8384));
  jand g08123(.dina(n8382), .dinb(n7977), .dout(n8385));
  jnot g08124(.din(n8385), .dout(n8386));
  jand g08125(.dina(n8386), .dinb(n8384), .dout(n8387));
  jnot g08126(.din(n8387), .dout(n8388));
  jor  g08127(.dina(n8388), .dinb(n8380), .dout(n8389));
  jand g08128(.dina(n8389), .dinb(n8379), .dout(n8390));
  jor  g08129(.dina(n8390), .dinb(n305), .dout(n8391));
  jand g08130(.dina(n8379), .dinb(n305), .dout(n8392));
  jand g08131(.dina(n8392), .dinb(n8389), .dout(n8393));
  jnot g08132(.din(n7979), .dout(n8394));
  jand g08133(.dina(asqrt[25] ), .dinb(n8394), .dout(n8395));
  jand g08134(.dina(n8395), .dinb(n7986), .dout(n8396));
  jor  g08135(.dina(n8396), .dinb(n7984), .dout(n8397));
  jand g08136(.dina(n8395), .dinb(n7987), .dout(n8398));
  jnot g08137(.din(n8398), .dout(n8399));
  jand g08138(.dina(n8399), .dinb(n8397), .dout(n8400));
  jnot g08139(.din(n8400), .dout(n8401));
  jor  g08140(.dina(n8401), .dinb(n8393), .dout(n8402));
  jand g08141(.dina(n8402), .dinb(n8391), .dout(n8403));
  jor  g08142(.dina(n8403), .dinb(n290), .dout(n8404));
  jxor g08143(.dina(n7988), .dinb(n305), .dout(n8405));
  jor  g08144(.dina(n8405), .dinb(n8058), .dout(n8406));
  jxor g08145(.dina(n8406), .dinb(n7999), .dout(n8407));
  jand g08146(.dina(n8403), .dinb(n290), .dout(n8408));
  jor  g08147(.dina(n8408), .dinb(n8407), .dout(n8409));
  jand g08148(.dina(n8409), .dinb(n8404), .dout(n8410));
  jor  g08149(.dina(n8410), .dinb(n223), .dout(n8411));
  jnot g08150(.din(n8004), .dout(n8412));
  jor  g08151(.dina(n8412), .dinb(n8002), .dout(n8413));
  jor  g08152(.dina(n8413), .dinb(n8058), .dout(n8414));
  jxor g08153(.dina(n8414), .dinb(n8013), .dout(n8415));
  jand g08154(.dina(n8404), .dinb(n223), .dout(n8416));
  jand g08155(.dina(n8416), .dinb(n8409), .dout(n8417));
  jor  g08156(.dina(n8417), .dinb(n8415), .dout(n8418));
  jand g08157(.dina(n8418), .dinb(n8411), .dout(n8419));
  jor  g08158(.dina(n8419), .dinb(n199), .dout(n8420));
  jand g08159(.dina(n8419), .dinb(n199), .dout(n8421));
  jnot g08160(.din(n8016), .dout(n8422));
  jand g08161(.dina(asqrt[25] ), .dinb(n8422), .dout(n8423));
  jand g08162(.dina(n8423), .dinb(n8021), .dout(n8424));
  jor  g08163(.dina(n8424), .dinb(n8020), .dout(n8425));
  jand g08164(.dina(n8423), .dinb(n8022), .dout(n8426));
  jnot g08165(.din(n8426), .dout(n8427));
  jand g08166(.dina(n8427), .dinb(n8425), .dout(n8428));
  jnot g08167(.din(n8428), .dout(n8429));
  jor  g08168(.dina(n8429), .dinb(n8421), .dout(n8430));
  jand g08169(.dina(n8430), .dinb(n8420), .dout(n8431));
  jnot g08170(.din(n8024), .dout(n8432));
  jand g08171(.dina(asqrt[25] ), .dinb(n8432), .dout(n8433));
  jand g08172(.dina(n8433), .dinb(n8031), .dout(n8434));
  jor  g08173(.dina(n8434), .dinb(n8029), .dout(n8435));
  jand g08174(.dina(n8433), .dinb(n8032), .dout(n8436));
  jnot g08175(.din(n8436), .dout(n8437));
  jand g08176(.dina(n8437), .dinb(n8435), .dout(n8438));
  jnot g08177(.din(n8438), .dout(n8439));
  jand g08178(.dina(asqrt[25] ), .dinb(n8046), .dout(n8440));
  jand g08179(.dina(n8440), .dinb(n8033), .dout(n8441));
  jor  g08180(.dina(n8441), .dinb(n8080), .dout(n8442));
  jor  g08181(.dina(n8442), .dinb(n8439), .dout(n8443));
  jor  g08182(.dina(n8443), .dinb(n8431), .dout(n8444));
  jand g08183(.dina(n8444), .dinb(n194), .dout(n8445));
  jand g08184(.dina(n8439), .dinb(n8431), .dout(n8446));
  jor  g08185(.dina(n8440), .dinb(n8033), .dout(n8447));
  jand g08186(.dina(n8046), .dinb(n8033), .dout(n8448));
  jor  g08187(.dina(n8448), .dinb(n194), .dout(n8449));
  jnot g08188(.din(n8449), .dout(n8450));
  jand g08189(.dina(n8450), .dinb(n8447), .dout(n8451));
  jor  g08190(.dina(n8451), .dinb(n8446), .dout(n8454));
  jor  g08191(.dina(n8454), .dinb(n8445), .dout(asqrt[24] ));
  jxor g08192(.dina(n8185), .dinb(n3907), .dout(n8456));
  jand g08193(.dina(n8456), .dinb(asqrt[24] ), .dout(n8457));
  jxor g08194(.dina(n8457), .dinb(n8061), .dout(n8458));
  jand g08195(.dina(asqrt[24] ), .dinb(a[48] ), .dout(n8459));
  jnot g08196(.din(a[46] ), .dout(n8460));
  jnot g08197(.din(a[47] ), .dout(n8461));
  jand g08198(.dina(n8063), .dinb(n8461), .dout(n8462));
  jand g08199(.dina(n8462), .dinb(n8460), .dout(n8463));
  jor  g08200(.dina(n8463), .dinb(n8459), .dout(n8464));
  jand g08201(.dina(n8464), .dinb(asqrt[25] ), .dout(n8465));
  jand g08202(.dina(asqrt[24] ), .dinb(n8063), .dout(n8466));
  jxor g08203(.dina(n8466), .dinb(n8064), .dout(n8467));
  jor  g08204(.dina(n8464), .dinb(asqrt[25] ), .dout(n8468));
  jand g08205(.dina(n8468), .dinb(n8467), .dout(n8469));
  jor  g08206(.dina(n8469), .dinb(n8465), .dout(n8470));
  jand g08207(.dina(n8470), .dinb(asqrt[26] ), .dout(n8471));
  jor  g08208(.dina(n8465), .dinb(asqrt[26] ), .dout(n8472));
  jor  g08209(.dina(n8472), .dinb(n8469), .dout(n8473));
  jand g08210(.dina(n8466), .dinb(n8064), .dout(n8474));
  jnot g08211(.din(n8445), .dout(n8475));
  jnot g08212(.din(n8446), .dout(n8476));
  jnot g08213(.din(n8451), .dout(n8477));
  jand g08214(.dina(n8477), .dinb(asqrt[25] ), .dout(n8478));
  jand g08215(.dina(n8478), .dinb(n8476), .dout(n8479));
  jand g08216(.dina(n8479), .dinb(n8475), .dout(n8480));
  jor  g08217(.dina(n8480), .dinb(n8474), .dout(n8481));
  jxor g08218(.dina(n8481), .dinb(n7647), .dout(n8482));
  jand g08219(.dina(n8482), .dinb(n8473), .dout(n8483));
  jor  g08220(.dina(n8483), .dinb(n8471), .dout(n8484));
  jand g08221(.dina(n8484), .dinb(asqrt[27] ), .dout(n8485));
  jor  g08222(.dina(n8484), .dinb(asqrt[27] ), .dout(n8486));
  jxor g08223(.dina(n8068), .dinb(n8053), .dout(n8487));
  jand g08224(.dina(n8487), .dinb(asqrt[24] ), .dout(n8488));
  jxor g08225(.dina(n8488), .dinb(n8071), .dout(n8489));
  jnot g08226(.din(n8489), .dout(n8490));
  jand g08227(.dina(n8490), .dinb(n8486), .dout(n8491));
  jor  g08228(.dina(n8491), .dinb(n8485), .dout(n8492));
  jand g08229(.dina(n8492), .dinb(asqrt[28] ), .dout(n8493));
  jnot g08230(.din(n8077), .dout(n8494));
  jand g08231(.dina(n8494), .dinb(n8075), .dout(n8495));
  jand g08232(.dina(n8495), .dinb(asqrt[24] ), .dout(n8496));
  jxor g08233(.dina(n8496), .dinb(n8085), .dout(n8497));
  jnot g08234(.din(n8497), .dout(n8498));
  jor  g08235(.dina(n8485), .dinb(asqrt[28] ), .dout(n8499));
  jor  g08236(.dina(n8499), .dinb(n8491), .dout(n8500));
  jand g08237(.dina(n8500), .dinb(n8498), .dout(n8501));
  jor  g08238(.dina(n8501), .dinb(n8493), .dout(n8502));
  jand g08239(.dina(n8502), .dinb(asqrt[29] ), .dout(n8503));
  jor  g08240(.dina(n8502), .dinb(asqrt[29] ), .dout(n8504));
  jnot g08241(.din(n8092), .dout(n8505));
  jxor g08242(.dina(n8087), .dinb(n7260), .dout(n8506));
  jand g08243(.dina(n8506), .dinb(asqrt[24] ), .dout(n8507));
  jxor g08244(.dina(n8507), .dinb(n8505), .dout(n8508));
  jand g08245(.dina(n8508), .dinb(n8504), .dout(n8509));
  jor  g08246(.dina(n8509), .dinb(n8503), .dout(n8510));
  jand g08247(.dina(n8510), .dinb(asqrt[30] ), .dout(n8511));
  jor  g08248(.dina(n8503), .dinb(asqrt[30] ), .dout(n8512));
  jor  g08249(.dina(n8512), .dinb(n8509), .dout(n8513));
  jnot g08250(.din(n8099), .dout(n8514));
  jnot g08251(.din(n8101), .dout(n8515));
  jand g08252(.dina(asqrt[24] ), .dinb(n8095), .dout(n8516));
  jand g08253(.dina(n8516), .dinb(n8515), .dout(n8517));
  jor  g08254(.dina(n8517), .dinb(n8514), .dout(n8518));
  jnot g08255(.din(n8102), .dout(n8519));
  jand g08256(.dina(n8516), .dinb(n8519), .dout(n8520));
  jnot g08257(.din(n8520), .dout(n8521));
  jand g08258(.dina(n8521), .dinb(n8518), .dout(n8522));
  jand g08259(.dina(n8522), .dinb(n8513), .dout(n8523));
  jor  g08260(.dina(n8523), .dinb(n8511), .dout(n8524));
  jand g08261(.dina(n8524), .dinb(asqrt[31] ), .dout(n8525));
  jor  g08262(.dina(n8524), .dinb(asqrt[31] ), .dout(n8526));
  jxor g08263(.dina(n8103), .dinb(n6500), .dout(n8527));
  jand g08264(.dina(n8527), .dinb(asqrt[24] ), .dout(n8528));
  jxor g08265(.dina(n8528), .dinb(n8108), .dout(n8529));
  jand g08266(.dina(n8529), .dinb(n8526), .dout(n8530));
  jor  g08267(.dina(n8530), .dinb(n8525), .dout(n8531));
  jand g08268(.dina(n8531), .dinb(asqrt[32] ), .dout(n8532));
  jnot g08269(.din(n8114), .dout(n8533));
  jand g08270(.dina(n8533), .dinb(n8112), .dout(n8534));
  jand g08271(.dina(n8534), .dinb(asqrt[24] ), .dout(n8535));
  jxor g08272(.dina(n8535), .dinb(n8123), .dout(n8536));
  jnot g08273(.din(n8536), .dout(n8537));
  jor  g08274(.dina(n8525), .dinb(asqrt[32] ), .dout(n8538));
  jor  g08275(.dina(n8538), .dinb(n8530), .dout(n8539));
  jand g08276(.dina(n8539), .dinb(n8537), .dout(n8540));
  jor  g08277(.dina(n8540), .dinb(n8532), .dout(n8541));
  jand g08278(.dina(n8541), .dinb(asqrt[33] ), .dout(n8542));
  jor  g08279(.dina(n8541), .dinb(asqrt[33] ), .dout(n8543));
  jxor g08280(.dina(n8125), .dinb(n5788), .dout(n8544));
  jand g08281(.dina(n8544), .dinb(asqrt[24] ), .dout(n8545));
  jxor g08282(.dina(n8545), .dinb(n8131), .dout(n8546));
  jand g08283(.dina(n8546), .dinb(n8543), .dout(n8547));
  jor  g08284(.dina(n8547), .dinb(n8542), .dout(n8548));
  jand g08285(.dina(n8548), .dinb(asqrt[34] ), .dout(n8549));
  jor  g08286(.dina(n8542), .dinb(asqrt[34] ), .dout(n8550));
  jor  g08287(.dina(n8550), .dinb(n8547), .dout(n8551));
  jnot g08288(.din(n8139), .dout(n8552));
  jnot g08289(.din(n8141), .dout(n8553));
  jand g08290(.dina(asqrt[24] ), .dinb(n8135), .dout(n8554));
  jand g08291(.dina(n8554), .dinb(n8553), .dout(n8555));
  jor  g08292(.dina(n8555), .dinb(n8552), .dout(n8556));
  jnot g08293(.din(n8142), .dout(n8557));
  jand g08294(.dina(n8554), .dinb(n8557), .dout(n8558));
  jnot g08295(.din(n8558), .dout(n8559));
  jand g08296(.dina(n8559), .dinb(n8556), .dout(n8560));
  jand g08297(.dina(n8560), .dinb(n8551), .dout(n8561));
  jor  g08298(.dina(n8561), .dinb(n8549), .dout(n8562));
  jand g08299(.dina(n8562), .dinb(asqrt[35] ), .dout(n8563));
  jxor g08300(.dina(n8143), .dinb(n5116), .dout(n8564));
  jand g08301(.dina(n8564), .dinb(asqrt[24] ), .dout(n8565));
  jxor g08302(.dina(n8565), .dinb(n8150), .dout(n8566));
  jnot g08303(.din(n8566), .dout(n8567));
  jor  g08304(.dina(n8562), .dinb(asqrt[35] ), .dout(n8568));
  jand g08305(.dina(n8568), .dinb(n8567), .dout(n8569));
  jor  g08306(.dina(n8569), .dinb(n8563), .dout(n8570));
  jand g08307(.dina(n8570), .dinb(asqrt[36] ), .dout(n8571));
  jnot g08308(.din(n8155), .dout(n8572));
  jand g08309(.dina(n8572), .dinb(n8153), .dout(n8573));
  jand g08310(.dina(n8573), .dinb(asqrt[24] ), .dout(n8574));
  jxor g08311(.dina(n8574), .dinb(n8163), .dout(n8575));
  jnot g08312(.din(n8575), .dout(n8576));
  jor  g08313(.dina(n8563), .dinb(asqrt[36] ), .dout(n8577));
  jor  g08314(.dina(n8577), .dinb(n8569), .dout(n8578));
  jand g08315(.dina(n8578), .dinb(n8576), .dout(n8579));
  jor  g08316(.dina(n8579), .dinb(n8571), .dout(n8580));
  jand g08317(.dina(n8580), .dinb(asqrt[37] ), .dout(n8581));
  jor  g08318(.dina(n8580), .dinb(asqrt[37] ), .dout(n8582));
  jnot g08319(.din(n8169), .dout(n8583));
  jnot g08320(.din(n8170), .dout(n8584));
  jand g08321(.dina(asqrt[24] ), .dinb(n8166), .dout(n8585));
  jand g08322(.dina(n8585), .dinb(n8584), .dout(n8586));
  jor  g08323(.dina(n8586), .dinb(n8583), .dout(n8587));
  jnot g08324(.din(n8171), .dout(n8588));
  jand g08325(.dina(n8585), .dinb(n8588), .dout(n8589));
  jnot g08326(.din(n8589), .dout(n8590));
  jand g08327(.dina(n8590), .dinb(n8587), .dout(n8591));
  jand g08328(.dina(n8591), .dinb(n8582), .dout(n8592));
  jor  g08329(.dina(n8592), .dinb(n8581), .dout(n8593));
  jand g08330(.dina(n8593), .dinb(asqrt[38] ), .dout(n8594));
  jnot g08331(.din(n8175), .dout(n8595));
  jand g08332(.dina(n8595), .dinb(n8173), .dout(n8596));
  jand g08333(.dina(n8596), .dinb(asqrt[24] ), .dout(n8597));
  jxor g08334(.dina(n8597), .dinb(n8183), .dout(n8598));
  jnot g08335(.din(n8598), .dout(n8599));
  jor  g08336(.dina(n8581), .dinb(asqrt[38] ), .dout(n8600));
  jor  g08337(.dina(n8600), .dinb(n8592), .dout(n8601));
  jand g08338(.dina(n8601), .dinb(n8599), .dout(n8602));
  jor  g08339(.dina(n8602), .dinb(n8594), .dout(n8603));
  jand g08340(.dina(n8603), .dinb(asqrt[39] ), .dout(n8604));
  jnot g08341(.din(n8458), .dout(n8605));
  jor  g08342(.dina(n8603), .dinb(asqrt[39] ), .dout(n8606));
  jand g08343(.dina(n8606), .dinb(n8605), .dout(n8607));
  jor  g08344(.dina(n8607), .dinb(n8604), .dout(n8608));
  jand g08345(.dina(n8608), .dinb(asqrt[40] ), .dout(n8609));
  jor  g08346(.dina(n8604), .dinb(asqrt[40] ), .dout(n8610));
  jor  g08347(.dina(n8610), .dinb(n8607), .dout(n8611));
  jnot g08348(.din(n8194), .dout(n8612));
  jnot g08349(.din(n8196), .dout(n8613));
  jand g08350(.dina(asqrt[24] ), .dinb(n8190), .dout(n8614));
  jand g08351(.dina(n8614), .dinb(n8613), .dout(n8615));
  jor  g08352(.dina(n8615), .dinb(n8612), .dout(n8616));
  jnot g08353(.din(n8197), .dout(n8617));
  jand g08354(.dina(n8614), .dinb(n8617), .dout(n8618));
  jnot g08355(.din(n8618), .dout(n8619));
  jand g08356(.dina(n8619), .dinb(n8616), .dout(n8620));
  jand g08357(.dina(n8620), .dinb(n8611), .dout(n8621));
  jor  g08358(.dina(n8621), .dinb(n8609), .dout(n8622));
  jand g08359(.dina(n8622), .dinb(asqrt[41] ), .dout(n8623));
  jor  g08360(.dina(n8622), .dinb(asqrt[41] ), .dout(n8624));
  jnot g08361(.din(n8202), .dout(n8625));
  jnot g08362(.din(n8203), .dout(n8626));
  jand g08363(.dina(asqrt[24] ), .dinb(n8199), .dout(n8627));
  jand g08364(.dina(n8627), .dinb(n8626), .dout(n8628));
  jor  g08365(.dina(n8628), .dinb(n8625), .dout(n8629));
  jnot g08366(.din(n8204), .dout(n8630));
  jand g08367(.dina(n8627), .dinb(n8630), .dout(n8631));
  jnot g08368(.din(n8631), .dout(n8632));
  jand g08369(.dina(n8632), .dinb(n8629), .dout(n8633));
  jand g08370(.dina(n8633), .dinb(n8624), .dout(n8634));
  jor  g08371(.dina(n8634), .dinb(n8623), .dout(n8635));
  jand g08372(.dina(n8635), .dinb(asqrt[42] ), .dout(n8636));
  jor  g08373(.dina(n8623), .dinb(asqrt[42] ), .dout(n8637));
  jor  g08374(.dina(n8637), .dinb(n8634), .dout(n8638));
  jnot g08375(.din(n8210), .dout(n8639));
  jnot g08376(.din(n8212), .dout(n8640));
  jand g08377(.dina(asqrt[24] ), .dinb(n8206), .dout(n8641));
  jand g08378(.dina(n8641), .dinb(n8640), .dout(n8642));
  jor  g08379(.dina(n8642), .dinb(n8639), .dout(n8643));
  jnot g08380(.din(n8213), .dout(n8644));
  jand g08381(.dina(n8641), .dinb(n8644), .dout(n8645));
  jnot g08382(.din(n8645), .dout(n8646));
  jand g08383(.dina(n8646), .dinb(n8643), .dout(n8647));
  jand g08384(.dina(n8647), .dinb(n8638), .dout(n8648));
  jor  g08385(.dina(n8648), .dinb(n8636), .dout(n8649));
  jand g08386(.dina(n8649), .dinb(asqrt[43] ), .dout(n8650));
  jxor g08387(.dina(n8214), .dinb(n2870), .dout(n8651));
  jand g08388(.dina(n8651), .dinb(asqrt[24] ), .dout(n8652));
  jxor g08389(.dina(n8652), .dinb(n8224), .dout(n8653));
  jnot g08390(.din(n8653), .dout(n8654));
  jor  g08391(.dina(n8649), .dinb(asqrt[43] ), .dout(n8655));
  jand g08392(.dina(n8655), .dinb(n8654), .dout(n8656));
  jor  g08393(.dina(n8656), .dinb(n8650), .dout(n8657));
  jand g08394(.dina(n8657), .dinb(asqrt[44] ), .dout(n8658));
  jnot g08395(.din(n8229), .dout(n8659));
  jand g08396(.dina(n8659), .dinb(n8227), .dout(n8660));
  jand g08397(.dina(n8660), .dinb(asqrt[24] ), .dout(n8661));
  jxor g08398(.dina(n8661), .dinb(n8237), .dout(n8662));
  jnot g08399(.din(n8662), .dout(n8663));
  jor  g08400(.dina(n8650), .dinb(asqrt[44] ), .dout(n8664));
  jor  g08401(.dina(n8664), .dinb(n8656), .dout(n8665));
  jand g08402(.dina(n8665), .dinb(n8663), .dout(n8666));
  jor  g08403(.dina(n8666), .dinb(n8658), .dout(n8667));
  jand g08404(.dina(n8667), .dinb(asqrt[45] ), .dout(n8668));
  jor  g08405(.dina(n8667), .dinb(asqrt[45] ), .dout(n8669));
  jnot g08406(.din(n8243), .dout(n8670));
  jnot g08407(.din(n8244), .dout(n8671));
  jand g08408(.dina(asqrt[24] ), .dinb(n8240), .dout(n8672));
  jand g08409(.dina(n8672), .dinb(n8671), .dout(n8673));
  jor  g08410(.dina(n8673), .dinb(n8670), .dout(n8674));
  jnot g08411(.din(n8245), .dout(n8675));
  jand g08412(.dina(n8672), .dinb(n8675), .dout(n8676));
  jnot g08413(.din(n8676), .dout(n8677));
  jand g08414(.dina(n8677), .dinb(n8674), .dout(n8678));
  jand g08415(.dina(n8678), .dinb(n8669), .dout(n8679));
  jor  g08416(.dina(n8679), .dinb(n8668), .dout(n8680));
  jand g08417(.dina(n8680), .dinb(asqrt[46] ), .dout(n8681));
  jor  g08418(.dina(n8668), .dinb(asqrt[46] ), .dout(n8682));
  jor  g08419(.dina(n8682), .dinb(n8679), .dout(n8683));
  jnot g08420(.din(n8251), .dout(n8684));
  jnot g08421(.din(n8253), .dout(n8685));
  jand g08422(.dina(asqrt[24] ), .dinb(n8247), .dout(n8686));
  jand g08423(.dina(n8686), .dinb(n8685), .dout(n8687));
  jor  g08424(.dina(n8687), .dinb(n8684), .dout(n8688));
  jnot g08425(.din(n8254), .dout(n8689));
  jand g08426(.dina(n8686), .dinb(n8689), .dout(n8690));
  jnot g08427(.din(n8690), .dout(n8691));
  jand g08428(.dina(n8691), .dinb(n8688), .dout(n8692));
  jand g08429(.dina(n8692), .dinb(n8683), .dout(n8693));
  jor  g08430(.dina(n8693), .dinb(n8681), .dout(n8694));
  jand g08431(.dina(n8694), .dinb(asqrt[47] ), .dout(n8695));
  jxor g08432(.dina(n8255), .dinb(n2005), .dout(n8696));
  jand g08433(.dina(n8696), .dinb(asqrt[24] ), .dout(n8697));
  jxor g08434(.dina(n8697), .dinb(n8265), .dout(n8698));
  jnot g08435(.din(n8698), .dout(n8699));
  jor  g08436(.dina(n8694), .dinb(asqrt[47] ), .dout(n8700));
  jand g08437(.dina(n8700), .dinb(n8699), .dout(n8701));
  jor  g08438(.dina(n8701), .dinb(n8695), .dout(n8702));
  jand g08439(.dina(n8702), .dinb(asqrt[48] ), .dout(n8703));
  jnot g08440(.din(n8270), .dout(n8704));
  jand g08441(.dina(n8704), .dinb(n8268), .dout(n8705));
  jand g08442(.dina(n8705), .dinb(asqrt[24] ), .dout(n8706));
  jxor g08443(.dina(n8706), .dinb(n8278), .dout(n8707));
  jnot g08444(.din(n8707), .dout(n8708));
  jor  g08445(.dina(n8695), .dinb(asqrt[48] ), .dout(n8709));
  jor  g08446(.dina(n8709), .dinb(n8701), .dout(n8710));
  jand g08447(.dina(n8710), .dinb(n8708), .dout(n8711));
  jor  g08448(.dina(n8711), .dinb(n8703), .dout(n8712));
  jand g08449(.dina(n8712), .dinb(asqrt[49] ), .dout(n8713));
  jor  g08450(.dina(n8712), .dinb(asqrt[49] ), .dout(n8714));
  jnot g08451(.din(n8284), .dout(n8715));
  jnot g08452(.din(n8285), .dout(n8716));
  jand g08453(.dina(asqrt[24] ), .dinb(n8281), .dout(n8717));
  jand g08454(.dina(n8717), .dinb(n8716), .dout(n8718));
  jor  g08455(.dina(n8718), .dinb(n8715), .dout(n8719));
  jnot g08456(.din(n8286), .dout(n8720));
  jand g08457(.dina(n8717), .dinb(n8720), .dout(n8721));
  jnot g08458(.din(n8721), .dout(n8722));
  jand g08459(.dina(n8722), .dinb(n8719), .dout(n8723));
  jand g08460(.dina(n8723), .dinb(n8714), .dout(n8724));
  jor  g08461(.dina(n8724), .dinb(n8713), .dout(n8725));
  jand g08462(.dina(n8725), .dinb(asqrt[50] ), .dout(n8726));
  jor  g08463(.dina(n8713), .dinb(asqrt[50] ), .dout(n8727));
  jor  g08464(.dina(n8727), .dinb(n8724), .dout(n8728));
  jnot g08465(.din(n8292), .dout(n8729));
  jnot g08466(.din(n8294), .dout(n8730));
  jand g08467(.dina(asqrt[24] ), .dinb(n8288), .dout(n8731));
  jand g08468(.dina(n8731), .dinb(n8730), .dout(n8732));
  jor  g08469(.dina(n8732), .dinb(n8729), .dout(n8733));
  jnot g08470(.din(n8295), .dout(n8734));
  jand g08471(.dina(n8731), .dinb(n8734), .dout(n8735));
  jnot g08472(.din(n8735), .dout(n8736));
  jand g08473(.dina(n8736), .dinb(n8733), .dout(n8737));
  jand g08474(.dina(n8737), .dinb(n8728), .dout(n8738));
  jor  g08475(.dina(n8738), .dinb(n8726), .dout(n8739));
  jand g08476(.dina(n8739), .dinb(asqrt[51] ), .dout(n8740));
  jxor g08477(.dina(n8296), .dinb(n1312), .dout(n8741));
  jand g08478(.dina(n8741), .dinb(asqrt[24] ), .dout(n8742));
  jxor g08479(.dina(n8742), .dinb(n8306), .dout(n8743));
  jnot g08480(.din(n8743), .dout(n8744));
  jor  g08481(.dina(n8739), .dinb(asqrt[51] ), .dout(n8745));
  jand g08482(.dina(n8745), .dinb(n8744), .dout(n8746));
  jor  g08483(.dina(n8746), .dinb(n8740), .dout(n8747));
  jand g08484(.dina(n8747), .dinb(asqrt[52] ), .dout(n8748));
  jnot g08485(.din(n8311), .dout(n8749));
  jand g08486(.dina(n8749), .dinb(n8309), .dout(n8750));
  jand g08487(.dina(n8750), .dinb(asqrt[24] ), .dout(n8751));
  jxor g08488(.dina(n8751), .dinb(n8319), .dout(n8752));
  jnot g08489(.din(n8752), .dout(n8753));
  jor  g08490(.dina(n8740), .dinb(asqrt[52] ), .dout(n8754));
  jor  g08491(.dina(n8754), .dinb(n8746), .dout(n8755));
  jand g08492(.dina(n8755), .dinb(n8753), .dout(n8756));
  jor  g08493(.dina(n8756), .dinb(n8748), .dout(n8757));
  jand g08494(.dina(n8757), .dinb(asqrt[53] ), .dout(n8758));
  jor  g08495(.dina(n8757), .dinb(asqrt[53] ), .dout(n8759));
  jnot g08496(.din(n8325), .dout(n8760));
  jnot g08497(.din(n8326), .dout(n8761));
  jand g08498(.dina(asqrt[24] ), .dinb(n8322), .dout(n8762));
  jand g08499(.dina(n8762), .dinb(n8761), .dout(n8763));
  jor  g08500(.dina(n8763), .dinb(n8760), .dout(n8764));
  jnot g08501(.din(n8327), .dout(n8765));
  jand g08502(.dina(n8762), .dinb(n8765), .dout(n8766));
  jnot g08503(.din(n8766), .dout(n8767));
  jand g08504(.dina(n8767), .dinb(n8764), .dout(n8768));
  jand g08505(.dina(n8768), .dinb(n8759), .dout(n8769));
  jor  g08506(.dina(n8769), .dinb(n8758), .dout(n8770));
  jand g08507(.dina(n8770), .dinb(asqrt[54] ), .dout(n8771));
  jor  g08508(.dina(n8758), .dinb(asqrt[54] ), .dout(n8772));
  jor  g08509(.dina(n8772), .dinb(n8769), .dout(n8773));
  jnot g08510(.din(n8333), .dout(n8774));
  jnot g08511(.din(n8335), .dout(n8775));
  jand g08512(.dina(asqrt[24] ), .dinb(n8329), .dout(n8776));
  jand g08513(.dina(n8776), .dinb(n8775), .dout(n8777));
  jor  g08514(.dina(n8777), .dinb(n8774), .dout(n8778));
  jnot g08515(.din(n8336), .dout(n8779));
  jand g08516(.dina(n8776), .dinb(n8779), .dout(n8780));
  jnot g08517(.din(n8780), .dout(n8781));
  jand g08518(.dina(n8781), .dinb(n8778), .dout(n8782));
  jand g08519(.dina(n8782), .dinb(n8773), .dout(n8783));
  jor  g08520(.dina(n8783), .dinb(n8771), .dout(n8784));
  jand g08521(.dina(n8784), .dinb(asqrt[55] ), .dout(n8785));
  jxor g08522(.dina(n8337), .dinb(n791), .dout(n8786));
  jand g08523(.dina(n8786), .dinb(asqrt[24] ), .dout(n8787));
  jxor g08524(.dina(n8787), .dinb(n8347), .dout(n8788));
  jnot g08525(.din(n8788), .dout(n8789));
  jor  g08526(.dina(n8784), .dinb(asqrt[55] ), .dout(n8790));
  jand g08527(.dina(n8790), .dinb(n8789), .dout(n8791));
  jor  g08528(.dina(n8791), .dinb(n8785), .dout(n8792));
  jand g08529(.dina(n8792), .dinb(asqrt[56] ), .dout(n8793));
  jnot g08530(.din(n8352), .dout(n8794));
  jand g08531(.dina(n8794), .dinb(n8350), .dout(n8795));
  jand g08532(.dina(n8795), .dinb(asqrt[24] ), .dout(n8796));
  jxor g08533(.dina(n8796), .dinb(n8360), .dout(n8797));
  jnot g08534(.din(n8797), .dout(n8798));
  jor  g08535(.dina(n8785), .dinb(asqrt[56] ), .dout(n8799));
  jor  g08536(.dina(n8799), .dinb(n8791), .dout(n8800));
  jand g08537(.dina(n8800), .dinb(n8798), .dout(n8801));
  jor  g08538(.dina(n8801), .dinb(n8793), .dout(n8802));
  jand g08539(.dina(n8802), .dinb(asqrt[57] ), .dout(n8803));
  jor  g08540(.dina(n8802), .dinb(asqrt[57] ), .dout(n8804));
  jnot g08541(.din(n8366), .dout(n8805));
  jnot g08542(.din(n8367), .dout(n8806));
  jand g08543(.dina(asqrt[24] ), .dinb(n8363), .dout(n8807));
  jand g08544(.dina(n8807), .dinb(n8806), .dout(n8808));
  jor  g08545(.dina(n8808), .dinb(n8805), .dout(n8809));
  jnot g08546(.din(n8368), .dout(n8810));
  jand g08547(.dina(n8807), .dinb(n8810), .dout(n8811));
  jnot g08548(.din(n8811), .dout(n8812));
  jand g08549(.dina(n8812), .dinb(n8809), .dout(n8813));
  jand g08550(.dina(n8813), .dinb(n8804), .dout(n8814));
  jor  g08551(.dina(n8814), .dinb(n8803), .dout(n8815));
  jand g08552(.dina(n8815), .dinb(asqrt[58] ), .dout(n8816));
  jor  g08553(.dina(n8803), .dinb(asqrt[58] ), .dout(n8817));
  jor  g08554(.dina(n8817), .dinb(n8814), .dout(n8818));
  jnot g08555(.din(n8374), .dout(n8819));
  jnot g08556(.din(n8376), .dout(n8820));
  jand g08557(.dina(asqrt[24] ), .dinb(n8370), .dout(n8821));
  jand g08558(.dina(n8821), .dinb(n8820), .dout(n8822));
  jor  g08559(.dina(n8822), .dinb(n8819), .dout(n8823));
  jnot g08560(.din(n8377), .dout(n8824));
  jand g08561(.dina(n8821), .dinb(n8824), .dout(n8825));
  jnot g08562(.din(n8825), .dout(n8826));
  jand g08563(.dina(n8826), .dinb(n8823), .dout(n8827));
  jand g08564(.dina(n8827), .dinb(n8818), .dout(n8828));
  jor  g08565(.dina(n8828), .dinb(n8816), .dout(n8829));
  jand g08566(.dina(n8829), .dinb(asqrt[59] ), .dout(n8830));
  jxor g08567(.dina(n8378), .dinb(n425), .dout(n8831));
  jand g08568(.dina(n8831), .dinb(asqrt[24] ), .dout(n8832));
  jxor g08569(.dina(n8832), .dinb(n8388), .dout(n8833));
  jnot g08570(.din(n8833), .dout(n8834));
  jor  g08571(.dina(n8829), .dinb(asqrt[59] ), .dout(n8835));
  jand g08572(.dina(n8835), .dinb(n8834), .dout(n8836));
  jor  g08573(.dina(n8836), .dinb(n8830), .dout(n8837));
  jand g08574(.dina(n8837), .dinb(asqrt[60] ), .dout(n8838));
  jnot g08575(.din(n8393), .dout(n8839));
  jand g08576(.dina(n8839), .dinb(n8391), .dout(n8840));
  jand g08577(.dina(n8840), .dinb(asqrt[24] ), .dout(n8841));
  jxor g08578(.dina(n8841), .dinb(n8401), .dout(n8842));
  jnot g08579(.din(n8842), .dout(n8843));
  jor  g08580(.dina(n8830), .dinb(asqrt[60] ), .dout(n8844));
  jor  g08581(.dina(n8844), .dinb(n8836), .dout(n8845));
  jand g08582(.dina(n8845), .dinb(n8843), .dout(n8846));
  jor  g08583(.dina(n8846), .dinb(n8838), .dout(n8847));
  jand g08584(.dina(n8847), .dinb(asqrt[61] ), .dout(n8848));
  jor  g08585(.dina(n8847), .dinb(asqrt[61] ), .dout(n8849));
  jnot g08586(.din(n8407), .dout(n8850));
  jnot g08587(.din(n8408), .dout(n8851));
  jand g08588(.dina(asqrt[24] ), .dinb(n8404), .dout(n8852));
  jand g08589(.dina(n8852), .dinb(n8851), .dout(n8853));
  jor  g08590(.dina(n8853), .dinb(n8850), .dout(n8854));
  jnot g08591(.din(n8409), .dout(n8855));
  jand g08592(.dina(n8852), .dinb(n8855), .dout(n8856));
  jnot g08593(.din(n8856), .dout(n8857));
  jand g08594(.dina(n8857), .dinb(n8854), .dout(n8858));
  jand g08595(.dina(n8858), .dinb(n8849), .dout(n8859));
  jor  g08596(.dina(n8859), .dinb(n8848), .dout(n8860));
  jand g08597(.dina(n8860), .dinb(asqrt[62] ), .dout(n8861));
  jor  g08598(.dina(n8848), .dinb(asqrt[62] ), .dout(n8862));
  jor  g08599(.dina(n8862), .dinb(n8859), .dout(n8863));
  jnot g08600(.din(n8415), .dout(n8864));
  jnot g08601(.din(n8417), .dout(n8865));
  jand g08602(.dina(asqrt[24] ), .dinb(n8411), .dout(n8866));
  jand g08603(.dina(n8866), .dinb(n8865), .dout(n8867));
  jor  g08604(.dina(n8867), .dinb(n8864), .dout(n8868));
  jnot g08605(.din(n8418), .dout(n8869));
  jand g08606(.dina(n8866), .dinb(n8869), .dout(n8870));
  jnot g08607(.din(n8870), .dout(n8871));
  jand g08608(.dina(n8871), .dinb(n8868), .dout(n8872));
  jand g08609(.dina(n8872), .dinb(n8863), .dout(n8873));
  jor  g08610(.dina(n8873), .dinb(n8861), .dout(n8874));
  jxor g08611(.dina(n8419), .dinb(n199), .dout(n8875));
  jand g08612(.dina(n8875), .dinb(asqrt[24] ), .dout(n8876));
  jxor g08613(.dina(n8876), .dinb(n8429), .dout(n8877));
  jnot g08614(.din(n8431), .dout(n8878));
  jand g08615(.dina(asqrt[24] ), .dinb(n8438), .dout(n8879));
  jand g08616(.dina(n8879), .dinb(n8878), .dout(n8880));
  jor  g08617(.dina(n8880), .dinb(n8446), .dout(n8881));
  jor  g08618(.dina(n8881), .dinb(n8877), .dout(n8882));
  jnot g08619(.din(n8882), .dout(n8883));
  jand g08620(.dina(n8883), .dinb(n8874), .dout(n8884));
  jor  g08621(.dina(n8884), .dinb(asqrt[63] ), .dout(n8885));
  jnot g08622(.din(n8877), .dout(n8886));
  jor  g08623(.dina(n8886), .dinb(n8874), .dout(n8887));
  jor  g08624(.dina(n8879), .dinb(n8878), .dout(n8888));
  jand g08625(.dina(n8438), .dinb(n8878), .dout(n8889));
  jor  g08626(.dina(n8889), .dinb(n194), .dout(n8890));
  jnot g08627(.din(n8890), .dout(n8891));
  jand g08628(.dina(n8891), .dinb(n8888), .dout(n8892));
  jnot g08629(.din(asqrt[24] ), .dout(n8893));
  jnot g08630(.din(n8892), .dout(n8896));
  jand g08631(.dina(n8896), .dinb(n8887), .dout(n8897));
  jand g08632(.dina(n8897), .dinb(n8885), .dout(n8898));
  jxor g08633(.dina(n8603), .dinb(n3376), .dout(n8899));
  jor  g08634(.dina(n8899), .dinb(n8898), .dout(n8900));
  jxor g08635(.dina(n8900), .dinb(n8458), .dout(n8901));
  jor  g08636(.dina(n8898), .dinb(n8460), .dout(n8902));
  jnot g08637(.din(a[44] ), .dout(n8903));
  jnot g08638(.din(a[45] ), .dout(n8904));
  jand g08639(.dina(n8460), .dinb(n8904), .dout(n8905));
  jand g08640(.dina(n8905), .dinb(n8903), .dout(n8906));
  jnot g08641(.din(n8906), .dout(n8907));
  jand g08642(.dina(n8907), .dinb(n8902), .dout(n8908));
  jor  g08643(.dina(n8908), .dinb(n8893), .dout(n8909));
  jor  g08644(.dina(n8898), .dinb(a[46] ), .dout(n8910));
  jxor g08645(.dina(n8910), .dinb(n8461), .dout(n8911));
  jand g08646(.dina(n8908), .dinb(n8893), .dout(n8912));
  jor  g08647(.dina(n8912), .dinb(n8911), .dout(n8913));
  jand g08648(.dina(n8913), .dinb(n8909), .dout(n8914));
  jor  g08649(.dina(n8914), .dinb(n8058), .dout(n8915));
  jand g08650(.dina(n8909), .dinb(n8058), .dout(n8916));
  jand g08651(.dina(n8916), .dinb(n8913), .dout(n8917));
  jor  g08652(.dina(n8910), .dinb(a[47] ), .dout(n8918));
  jnot g08653(.din(n8885), .dout(n8919));
  jnot g08654(.din(n8887), .dout(n8920));
  jor  g08655(.dina(n8892), .dinb(n8893), .dout(n8921));
  jor  g08656(.dina(n8921), .dinb(n8920), .dout(n8922));
  jor  g08657(.dina(n8922), .dinb(n8919), .dout(n8923));
  jand g08658(.dina(n8923), .dinb(n8918), .dout(n8924));
  jxor g08659(.dina(n8924), .dinb(n8063), .dout(n8925));
  jor  g08660(.dina(n8925), .dinb(n8917), .dout(n8926));
  jand g08661(.dina(n8926), .dinb(n8915), .dout(n8927));
  jor  g08662(.dina(n8927), .dinb(n8053), .dout(n8928));
  jand g08663(.dina(n8927), .dinb(n8053), .dout(n8929));
  jxor g08664(.dina(n8464), .dinb(n8058), .dout(n8930));
  jor  g08665(.dina(n8930), .dinb(n8898), .dout(n8931));
  jxor g08666(.dina(n8931), .dinb(n8467), .dout(n8932));
  jor  g08667(.dina(n8932), .dinb(n8929), .dout(n8933));
  jand g08668(.dina(n8933), .dinb(n8928), .dout(n8934));
  jor  g08669(.dina(n8934), .dinb(n7265), .dout(n8935));
  jnot g08670(.din(n8473), .dout(n8936));
  jor  g08671(.dina(n8936), .dinb(n8471), .dout(n8937));
  jor  g08672(.dina(n8937), .dinb(n8898), .dout(n8938));
  jxor g08673(.dina(n8938), .dinb(n8482), .dout(n8939));
  jand g08674(.dina(n8928), .dinb(n7265), .dout(n8940));
  jand g08675(.dina(n8940), .dinb(n8933), .dout(n8941));
  jor  g08676(.dina(n8941), .dinb(n8939), .dout(n8942));
  jand g08677(.dina(n8942), .dinb(n8935), .dout(n8943));
  jor  g08678(.dina(n8943), .dinb(n7260), .dout(n8944));
  jand g08679(.dina(n8943), .dinb(n7260), .dout(n8945));
  jxor g08680(.dina(n8484), .dinb(n7265), .dout(n8946));
  jor  g08681(.dina(n8946), .dinb(n8898), .dout(n8947));
  jxor g08682(.dina(n8947), .dinb(n8489), .dout(n8948));
  jnot g08683(.din(n8948), .dout(n8949));
  jor  g08684(.dina(n8949), .dinb(n8945), .dout(n8950));
  jand g08685(.dina(n8950), .dinb(n8944), .dout(n8951));
  jor  g08686(.dina(n8951), .dinb(n6505), .dout(n8952));
  jand g08687(.dina(n8944), .dinb(n6505), .dout(n8953));
  jand g08688(.dina(n8953), .dinb(n8950), .dout(n8954));
  jnot g08689(.din(n8493), .dout(n8955));
  jnot g08690(.din(n8898), .dout(asqrt[23] ));
  jand g08691(.dina(asqrt[23] ), .dinb(n8955), .dout(n8957));
  jand g08692(.dina(n8957), .dinb(n8500), .dout(n8958));
  jor  g08693(.dina(n8958), .dinb(n8498), .dout(n8959));
  jand g08694(.dina(n8957), .dinb(n8501), .dout(n8960));
  jnot g08695(.din(n8960), .dout(n8961));
  jand g08696(.dina(n8961), .dinb(n8959), .dout(n8962));
  jnot g08697(.din(n8962), .dout(n8963));
  jor  g08698(.dina(n8963), .dinb(n8954), .dout(n8964));
  jand g08699(.dina(n8964), .dinb(n8952), .dout(n8965));
  jor  g08700(.dina(n8965), .dinb(n6500), .dout(n8966));
  jand g08701(.dina(n8965), .dinb(n6500), .dout(n8967));
  jnot g08702(.din(n8508), .dout(n8968));
  jxor g08703(.dina(n8502), .dinb(n6505), .dout(n8969));
  jor  g08704(.dina(n8969), .dinb(n8898), .dout(n8970));
  jxor g08705(.dina(n8970), .dinb(n8968), .dout(n8971));
  jnot g08706(.din(n8971), .dout(n8972));
  jor  g08707(.dina(n8972), .dinb(n8967), .dout(n8973));
  jand g08708(.dina(n8973), .dinb(n8966), .dout(n8974));
  jor  g08709(.dina(n8974), .dinb(n5793), .dout(n8975));
  jnot g08710(.din(n8513), .dout(n8976));
  jor  g08711(.dina(n8976), .dinb(n8511), .dout(n8977));
  jor  g08712(.dina(n8977), .dinb(n8898), .dout(n8978));
  jxor g08713(.dina(n8978), .dinb(n8522), .dout(n8979));
  jand g08714(.dina(n8966), .dinb(n5793), .dout(n8980));
  jand g08715(.dina(n8980), .dinb(n8973), .dout(n8981));
  jor  g08716(.dina(n8981), .dinb(n8979), .dout(n8982));
  jand g08717(.dina(n8982), .dinb(n8975), .dout(n8983));
  jor  g08718(.dina(n8983), .dinb(n5788), .dout(n8984));
  jand g08719(.dina(n8983), .dinb(n5788), .dout(n8985));
  jnot g08720(.din(n8529), .dout(n8986));
  jxor g08721(.dina(n8524), .dinb(n5793), .dout(n8987));
  jor  g08722(.dina(n8987), .dinb(n8898), .dout(n8988));
  jxor g08723(.dina(n8988), .dinb(n8986), .dout(n8989));
  jnot g08724(.din(n8989), .dout(n8990));
  jor  g08725(.dina(n8990), .dinb(n8985), .dout(n8991));
  jand g08726(.dina(n8991), .dinb(n8984), .dout(n8992));
  jor  g08727(.dina(n8992), .dinb(n5121), .dout(n8993));
  jand g08728(.dina(n8984), .dinb(n5121), .dout(n8994));
  jand g08729(.dina(n8994), .dinb(n8991), .dout(n8995));
  jnot g08730(.din(n8532), .dout(n8996));
  jand g08731(.dina(asqrt[23] ), .dinb(n8996), .dout(n8997));
  jand g08732(.dina(n8997), .dinb(n8539), .dout(n8998));
  jor  g08733(.dina(n8998), .dinb(n8537), .dout(n8999));
  jand g08734(.dina(n8997), .dinb(n8540), .dout(n9000));
  jnot g08735(.din(n9000), .dout(n9001));
  jand g08736(.dina(n9001), .dinb(n8999), .dout(n9002));
  jnot g08737(.din(n9002), .dout(n9003));
  jor  g08738(.dina(n9003), .dinb(n8995), .dout(n9004));
  jand g08739(.dina(n9004), .dinb(n8993), .dout(n9005));
  jor  g08740(.dina(n9005), .dinb(n5116), .dout(n9006));
  jxor g08741(.dina(n8541), .dinb(n5121), .dout(n9007));
  jor  g08742(.dina(n9007), .dinb(n8898), .dout(n9008));
  jxor g08743(.dina(n9008), .dinb(n8546), .dout(n9009));
  jand g08744(.dina(n9005), .dinb(n5116), .dout(n9010));
  jor  g08745(.dina(n9010), .dinb(n9009), .dout(n9011));
  jand g08746(.dina(n9011), .dinb(n9006), .dout(n9012));
  jor  g08747(.dina(n9012), .dinb(n4499), .dout(n9013));
  jnot g08748(.din(n8551), .dout(n9014));
  jor  g08749(.dina(n9014), .dinb(n8549), .dout(n9015));
  jor  g08750(.dina(n9015), .dinb(n8898), .dout(n9016));
  jxor g08751(.dina(n9016), .dinb(n8560), .dout(n9017));
  jand g08752(.dina(n9006), .dinb(n4499), .dout(n9018));
  jand g08753(.dina(n9018), .dinb(n9011), .dout(n9019));
  jor  g08754(.dina(n9019), .dinb(n9017), .dout(n9020));
  jand g08755(.dina(n9020), .dinb(n9013), .dout(n9021));
  jor  g08756(.dina(n9021), .dinb(n4494), .dout(n9022));
  jand g08757(.dina(n9021), .dinb(n4494), .dout(n9023));
  jnot g08758(.din(n8563), .dout(n9024));
  jand g08759(.dina(asqrt[23] ), .dinb(n9024), .dout(n9025));
  jand g08760(.dina(n9025), .dinb(n8568), .dout(n9026));
  jor  g08761(.dina(n9026), .dinb(n8567), .dout(n9027));
  jand g08762(.dina(n9025), .dinb(n8569), .dout(n9028));
  jnot g08763(.din(n9028), .dout(n9029));
  jand g08764(.dina(n9029), .dinb(n9027), .dout(n9030));
  jnot g08765(.din(n9030), .dout(n9031));
  jor  g08766(.dina(n9031), .dinb(n9023), .dout(n9032));
  jand g08767(.dina(n9032), .dinb(n9022), .dout(n9033));
  jor  g08768(.dina(n9033), .dinb(n3912), .dout(n9034));
  jand g08769(.dina(n9022), .dinb(n3912), .dout(n9035));
  jand g08770(.dina(n9035), .dinb(n9032), .dout(n9036));
  jnot g08771(.din(n8571), .dout(n9037));
  jand g08772(.dina(asqrt[23] ), .dinb(n9037), .dout(n9038));
  jand g08773(.dina(n9038), .dinb(n8578), .dout(n9039));
  jor  g08774(.dina(n9039), .dinb(n8576), .dout(n9040));
  jand g08775(.dina(n9038), .dinb(n8579), .dout(n9041));
  jnot g08776(.din(n9041), .dout(n9042));
  jand g08777(.dina(n9042), .dinb(n9040), .dout(n9043));
  jnot g08778(.din(n9043), .dout(n9044));
  jor  g08779(.dina(n9044), .dinb(n9036), .dout(n9045));
  jand g08780(.dina(n9045), .dinb(n9034), .dout(n9046));
  jor  g08781(.dina(n9046), .dinb(n3907), .dout(n9047));
  jxor g08782(.dina(n8580), .dinb(n3912), .dout(n9048));
  jor  g08783(.dina(n9048), .dinb(n8898), .dout(n9049));
  jxor g08784(.dina(n9049), .dinb(n8591), .dout(n9050));
  jand g08785(.dina(n9046), .dinb(n3907), .dout(n9051));
  jor  g08786(.dina(n9051), .dinb(n9050), .dout(n9052));
  jand g08787(.dina(n9052), .dinb(n9047), .dout(n9053));
  jor  g08788(.dina(n9053), .dinb(n3376), .dout(n9054));
  jand g08789(.dina(n9047), .dinb(n3376), .dout(n9055));
  jand g08790(.dina(n9055), .dinb(n9052), .dout(n9056));
  jnot g08791(.din(n8594), .dout(n9057));
  jand g08792(.dina(asqrt[23] ), .dinb(n9057), .dout(n9058));
  jand g08793(.dina(n9058), .dinb(n8601), .dout(n9059));
  jor  g08794(.dina(n9059), .dinb(n8599), .dout(n9060));
  jand g08795(.dina(n9058), .dinb(n8602), .dout(n9061));
  jnot g08796(.din(n9061), .dout(n9062));
  jand g08797(.dina(n9062), .dinb(n9060), .dout(n9063));
  jnot g08798(.din(n9063), .dout(n9064));
  jor  g08799(.dina(n9064), .dinb(n9056), .dout(n9065));
  jand g08800(.dina(n9065), .dinb(n9054), .dout(n9066));
  jor  g08801(.dina(n9066), .dinb(n3371), .dout(n9067));
  jnot g08802(.din(n8901), .dout(n9068));
  jand g08803(.dina(n9066), .dinb(n3371), .dout(n9069));
  jor  g08804(.dina(n9069), .dinb(n9068), .dout(n9070));
  jand g08805(.dina(n9070), .dinb(n9067), .dout(n9071));
  jor  g08806(.dina(n9071), .dinb(n2875), .dout(n9072));
  jnot g08807(.din(n8611), .dout(n9073));
  jor  g08808(.dina(n9073), .dinb(n8609), .dout(n9074));
  jor  g08809(.dina(n9074), .dinb(n8898), .dout(n9075));
  jxor g08810(.dina(n9075), .dinb(n8620), .dout(n9076));
  jand g08811(.dina(n9067), .dinb(n2875), .dout(n9077));
  jand g08812(.dina(n9077), .dinb(n9070), .dout(n9078));
  jor  g08813(.dina(n9078), .dinb(n9076), .dout(n9079));
  jand g08814(.dina(n9079), .dinb(n9072), .dout(n9080));
  jor  g08815(.dina(n9080), .dinb(n2870), .dout(n9081));
  jxor g08816(.dina(n8622), .dinb(n2875), .dout(n9082));
  jor  g08817(.dina(n9082), .dinb(n8898), .dout(n9083));
  jxor g08818(.dina(n9083), .dinb(n8633), .dout(n9084));
  jand g08819(.dina(n9080), .dinb(n2870), .dout(n9085));
  jor  g08820(.dina(n9085), .dinb(n9084), .dout(n9086));
  jand g08821(.dina(n9086), .dinb(n9081), .dout(n9087));
  jor  g08822(.dina(n9087), .dinb(n2425), .dout(n9088));
  jnot g08823(.din(n8638), .dout(n9089));
  jor  g08824(.dina(n9089), .dinb(n8636), .dout(n9090));
  jor  g08825(.dina(n9090), .dinb(n8898), .dout(n9091));
  jxor g08826(.dina(n9091), .dinb(n8647), .dout(n9092));
  jand g08827(.dina(n9081), .dinb(n2425), .dout(n9093));
  jand g08828(.dina(n9093), .dinb(n9086), .dout(n9094));
  jor  g08829(.dina(n9094), .dinb(n9092), .dout(n9095));
  jand g08830(.dina(n9095), .dinb(n9088), .dout(n9096));
  jor  g08831(.dina(n9096), .dinb(n2420), .dout(n9097));
  jand g08832(.dina(n9096), .dinb(n2420), .dout(n9098));
  jnot g08833(.din(n8650), .dout(n9099));
  jand g08834(.dina(asqrt[23] ), .dinb(n9099), .dout(n9100));
  jand g08835(.dina(n9100), .dinb(n8655), .dout(n9101));
  jor  g08836(.dina(n9101), .dinb(n8654), .dout(n9102));
  jand g08837(.dina(n9100), .dinb(n8656), .dout(n9103));
  jnot g08838(.din(n9103), .dout(n9104));
  jand g08839(.dina(n9104), .dinb(n9102), .dout(n9105));
  jnot g08840(.din(n9105), .dout(n9106));
  jor  g08841(.dina(n9106), .dinb(n9098), .dout(n9107));
  jand g08842(.dina(n9107), .dinb(n9097), .dout(n9108));
  jor  g08843(.dina(n9108), .dinb(n2010), .dout(n9109));
  jand g08844(.dina(n9097), .dinb(n2010), .dout(n9110));
  jand g08845(.dina(n9110), .dinb(n9107), .dout(n9111));
  jnot g08846(.din(n8658), .dout(n9112));
  jand g08847(.dina(asqrt[23] ), .dinb(n9112), .dout(n9113));
  jand g08848(.dina(n9113), .dinb(n8665), .dout(n9114));
  jor  g08849(.dina(n9114), .dinb(n8663), .dout(n9115));
  jand g08850(.dina(n9113), .dinb(n8666), .dout(n9116));
  jnot g08851(.din(n9116), .dout(n9117));
  jand g08852(.dina(n9117), .dinb(n9115), .dout(n9118));
  jnot g08853(.din(n9118), .dout(n9119));
  jor  g08854(.dina(n9119), .dinb(n9111), .dout(n9120));
  jand g08855(.dina(n9120), .dinb(n9109), .dout(n9121));
  jor  g08856(.dina(n9121), .dinb(n2005), .dout(n9122));
  jxor g08857(.dina(n8667), .dinb(n2010), .dout(n9123));
  jor  g08858(.dina(n9123), .dinb(n8898), .dout(n9124));
  jxor g08859(.dina(n9124), .dinb(n8678), .dout(n9125));
  jand g08860(.dina(n9121), .dinb(n2005), .dout(n9126));
  jor  g08861(.dina(n9126), .dinb(n9125), .dout(n9127));
  jand g08862(.dina(n9127), .dinb(n9122), .dout(n9128));
  jor  g08863(.dina(n9128), .dinb(n1646), .dout(n9129));
  jnot g08864(.din(n8683), .dout(n9130));
  jor  g08865(.dina(n9130), .dinb(n8681), .dout(n9131));
  jor  g08866(.dina(n9131), .dinb(n8898), .dout(n9132));
  jxor g08867(.dina(n9132), .dinb(n8692), .dout(n9133));
  jand g08868(.dina(n9122), .dinb(n1646), .dout(n9134));
  jand g08869(.dina(n9134), .dinb(n9127), .dout(n9135));
  jor  g08870(.dina(n9135), .dinb(n9133), .dout(n9136));
  jand g08871(.dina(n9136), .dinb(n9129), .dout(n9137));
  jor  g08872(.dina(n9137), .dinb(n1641), .dout(n9138));
  jand g08873(.dina(n9137), .dinb(n1641), .dout(n9139));
  jnot g08874(.din(n8695), .dout(n9140));
  jand g08875(.dina(asqrt[23] ), .dinb(n9140), .dout(n9141));
  jand g08876(.dina(n9141), .dinb(n8700), .dout(n9142));
  jor  g08877(.dina(n9142), .dinb(n8699), .dout(n9143));
  jand g08878(.dina(n9141), .dinb(n8701), .dout(n9144));
  jnot g08879(.din(n9144), .dout(n9145));
  jand g08880(.dina(n9145), .dinb(n9143), .dout(n9146));
  jnot g08881(.din(n9146), .dout(n9147));
  jor  g08882(.dina(n9147), .dinb(n9139), .dout(n9148));
  jand g08883(.dina(n9148), .dinb(n9138), .dout(n9149));
  jor  g08884(.dina(n9149), .dinb(n1317), .dout(n9150));
  jand g08885(.dina(n9138), .dinb(n1317), .dout(n9151));
  jand g08886(.dina(n9151), .dinb(n9148), .dout(n9152));
  jnot g08887(.din(n8703), .dout(n9153));
  jand g08888(.dina(asqrt[23] ), .dinb(n9153), .dout(n9154));
  jand g08889(.dina(n9154), .dinb(n8710), .dout(n9155));
  jor  g08890(.dina(n9155), .dinb(n8708), .dout(n9156));
  jand g08891(.dina(n9154), .dinb(n8711), .dout(n9157));
  jnot g08892(.din(n9157), .dout(n9158));
  jand g08893(.dina(n9158), .dinb(n9156), .dout(n9159));
  jnot g08894(.din(n9159), .dout(n9160));
  jor  g08895(.dina(n9160), .dinb(n9152), .dout(n9161));
  jand g08896(.dina(n9161), .dinb(n9150), .dout(n9162));
  jor  g08897(.dina(n9162), .dinb(n1312), .dout(n9163));
  jxor g08898(.dina(n8712), .dinb(n1317), .dout(n9164));
  jor  g08899(.dina(n9164), .dinb(n8898), .dout(n9165));
  jxor g08900(.dina(n9165), .dinb(n8723), .dout(n9166));
  jand g08901(.dina(n9162), .dinb(n1312), .dout(n9167));
  jor  g08902(.dina(n9167), .dinb(n9166), .dout(n9168));
  jand g08903(.dina(n9168), .dinb(n9163), .dout(n9169));
  jor  g08904(.dina(n9169), .dinb(n1039), .dout(n9170));
  jnot g08905(.din(n8728), .dout(n9171));
  jor  g08906(.dina(n9171), .dinb(n8726), .dout(n9172));
  jor  g08907(.dina(n9172), .dinb(n8898), .dout(n9173));
  jxor g08908(.dina(n9173), .dinb(n8737), .dout(n9174));
  jand g08909(.dina(n9163), .dinb(n1039), .dout(n9175));
  jand g08910(.dina(n9175), .dinb(n9168), .dout(n9176));
  jor  g08911(.dina(n9176), .dinb(n9174), .dout(n9177));
  jand g08912(.dina(n9177), .dinb(n9170), .dout(n9178));
  jor  g08913(.dina(n9178), .dinb(n1034), .dout(n9179));
  jand g08914(.dina(n9178), .dinb(n1034), .dout(n9180));
  jnot g08915(.din(n8740), .dout(n9181));
  jand g08916(.dina(asqrt[23] ), .dinb(n9181), .dout(n9182));
  jand g08917(.dina(n9182), .dinb(n8745), .dout(n9183));
  jor  g08918(.dina(n9183), .dinb(n8744), .dout(n9184));
  jand g08919(.dina(n9182), .dinb(n8746), .dout(n9185));
  jnot g08920(.din(n9185), .dout(n9186));
  jand g08921(.dina(n9186), .dinb(n9184), .dout(n9187));
  jnot g08922(.din(n9187), .dout(n9188));
  jor  g08923(.dina(n9188), .dinb(n9180), .dout(n9189));
  jand g08924(.dina(n9189), .dinb(n9179), .dout(n9190));
  jor  g08925(.dina(n9190), .dinb(n796), .dout(n9191));
  jand g08926(.dina(n9179), .dinb(n796), .dout(n9192));
  jand g08927(.dina(n9192), .dinb(n9189), .dout(n9193));
  jnot g08928(.din(n8748), .dout(n9194));
  jand g08929(.dina(asqrt[23] ), .dinb(n9194), .dout(n9195));
  jand g08930(.dina(n9195), .dinb(n8755), .dout(n9196));
  jor  g08931(.dina(n9196), .dinb(n8753), .dout(n9197));
  jand g08932(.dina(n9195), .dinb(n8756), .dout(n9198));
  jnot g08933(.din(n9198), .dout(n9199));
  jand g08934(.dina(n9199), .dinb(n9197), .dout(n9200));
  jnot g08935(.din(n9200), .dout(n9201));
  jor  g08936(.dina(n9201), .dinb(n9193), .dout(n9202));
  jand g08937(.dina(n9202), .dinb(n9191), .dout(n9203));
  jor  g08938(.dina(n9203), .dinb(n791), .dout(n9204));
  jxor g08939(.dina(n8757), .dinb(n796), .dout(n9205));
  jor  g08940(.dina(n9205), .dinb(n8898), .dout(n9206));
  jxor g08941(.dina(n9206), .dinb(n8768), .dout(n9207));
  jand g08942(.dina(n9203), .dinb(n791), .dout(n9208));
  jor  g08943(.dina(n9208), .dinb(n9207), .dout(n9209));
  jand g08944(.dina(n9209), .dinb(n9204), .dout(n9210));
  jor  g08945(.dina(n9210), .dinb(n595), .dout(n9211));
  jnot g08946(.din(n8773), .dout(n9212));
  jor  g08947(.dina(n9212), .dinb(n8771), .dout(n9213));
  jor  g08948(.dina(n9213), .dinb(n8898), .dout(n9214));
  jxor g08949(.dina(n9214), .dinb(n8782), .dout(n9215));
  jand g08950(.dina(n9204), .dinb(n595), .dout(n9216));
  jand g08951(.dina(n9216), .dinb(n9209), .dout(n9217));
  jor  g08952(.dina(n9217), .dinb(n9215), .dout(n9218));
  jand g08953(.dina(n9218), .dinb(n9211), .dout(n9219));
  jor  g08954(.dina(n9219), .dinb(n590), .dout(n9220));
  jand g08955(.dina(n9219), .dinb(n590), .dout(n9221));
  jnot g08956(.din(n8785), .dout(n9222));
  jand g08957(.dina(asqrt[23] ), .dinb(n9222), .dout(n9223));
  jand g08958(.dina(n9223), .dinb(n8790), .dout(n9224));
  jor  g08959(.dina(n9224), .dinb(n8789), .dout(n9225));
  jand g08960(.dina(n9223), .dinb(n8791), .dout(n9226));
  jnot g08961(.din(n9226), .dout(n9227));
  jand g08962(.dina(n9227), .dinb(n9225), .dout(n9228));
  jnot g08963(.din(n9228), .dout(n9229));
  jor  g08964(.dina(n9229), .dinb(n9221), .dout(n9230));
  jand g08965(.dina(n9230), .dinb(n9220), .dout(n9231));
  jor  g08966(.dina(n9231), .dinb(n430), .dout(n9232));
  jand g08967(.dina(n9220), .dinb(n430), .dout(n9233));
  jand g08968(.dina(n9233), .dinb(n9230), .dout(n9234));
  jnot g08969(.din(n8793), .dout(n9235));
  jand g08970(.dina(asqrt[23] ), .dinb(n9235), .dout(n9236));
  jand g08971(.dina(n9236), .dinb(n8800), .dout(n9237));
  jor  g08972(.dina(n9237), .dinb(n8798), .dout(n9238));
  jand g08973(.dina(n9236), .dinb(n8801), .dout(n9239));
  jnot g08974(.din(n9239), .dout(n9240));
  jand g08975(.dina(n9240), .dinb(n9238), .dout(n9241));
  jnot g08976(.din(n9241), .dout(n9242));
  jor  g08977(.dina(n9242), .dinb(n9234), .dout(n9243));
  jand g08978(.dina(n9243), .dinb(n9232), .dout(n9244));
  jor  g08979(.dina(n9244), .dinb(n425), .dout(n9245));
  jxor g08980(.dina(n8802), .dinb(n430), .dout(n9246));
  jor  g08981(.dina(n9246), .dinb(n8898), .dout(n9247));
  jxor g08982(.dina(n9247), .dinb(n8813), .dout(n9248));
  jand g08983(.dina(n9244), .dinb(n425), .dout(n9249));
  jor  g08984(.dina(n9249), .dinb(n9248), .dout(n9250));
  jand g08985(.dina(n9250), .dinb(n9245), .dout(n9251));
  jor  g08986(.dina(n9251), .dinb(n305), .dout(n9252));
  jnot g08987(.din(n8818), .dout(n9253));
  jor  g08988(.dina(n9253), .dinb(n8816), .dout(n9254));
  jor  g08989(.dina(n9254), .dinb(n8898), .dout(n9255));
  jxor g08990(.dina(n9255), .dinb(n8827), .dout(n9256));
  jand g08991(.dina(n9245), .dinb(n305), .dout(n9257));
  jand g08992(.dina(n9257), .dinb(n9250), .dout(n9258));
  jor  g08993(.dina(n9258), .dinb(n9256), .dout(n9259));
  jand g08994(.dina(n9259), .dinb(n9252), .dout(n9260));
  jor  g08995(.dina(n9260), .dinb(n290), .dout(n9261));
  jand g08996(.dina(n9260), .dinb(n290), .dout(n9262));
  jnot g08997(.din(n8830), .dout(n9263));
  jand g08998(.dina(asqrt[23] ), .dinb(n9263), .dout(n9264));
  jand g08999(.dina(n9264), .dinb(n8835), .dout(n9265));
  jor  g09000(.dina(n9265), .dinb(n8834), .dout(n9266));
  jand g09001(.dina(n9264), .dinb(n8836), .dout(n9267));
  jnot g09002(.din(n9267), .dout(n9268));
  jand g09003(.dina(n9268), .dinb(n9266), .dout(n9269));
  jnot g09004(.din(n9269), .dout(n9270));
  jor  g09005(.dina(n9270), .dinb(n9262), .dout(n9271));
  jand g09006(.dina(n9271), .dinb(n9261), .dout(n9272));
  jor  g09007(.dina(n9272), .dinb(n223), .dout(n9273));
  jand g09008(.dina(n9261), .dinb(n223), .dout(n9274));
  jand g09009(.dina(n9274), .dinb(n9271), .dout(n9275));
  jnot g09010(.din(n8838), .dout(n9276));
  jand g09011(.dina(asqrt[23] ), .dinb(n9276), .dout(n9277));
  jand g09012(.dina(n9277), .dinb(n8845), .dout(n9278));
  jor  g09013(.dina(n9278), .dinb(n8843), .dout(n9279));
  jand g09014(.dina(n9277), .dinb(n8846), .dout(n9280));
  jnot g09015(.din(n9280), .dout(n9281));
  jand g09016(.dina(n9281), .dinb(n9279), .dout(n9282));
  jnot g09017(.din(n9282), .dout(n9283));
  jor  g09018(.dina(n9283), .dinb(n9275), .dout(n9284));
  jand g09019(.dina(n9284), .dinb(n9273), .dout(n9285));
  jor  g09020(.dina(n9285), .dinb(n199), .dout(n9286));
  jand g09021(.dina(n9285), .dinb(n199), .dout(n9287));
  jxor g09022(.dina(n8847), .dinb(n223), .dout(n9288));
  jor  g09023(.dina(n9288), .dinb(n8898), .dout(n9289));
  jxor g09024(.dina(n9289), .dinb(n8858), .dout(n9290));
  jor  g09025(.dina(n9290), .dinb(n9287), .dout(n9291));
  jand g09026(.dina(n9291), .dinb(n9286), .dout(n9292));
  jnot g09027(.din(n8863), .dout(n9293));
  jor  g09028(.dina(n9293), .dinb(n8861), .dout(n9294));
  jor  g09029(.dina(n9294), .dinb(n8898), .dout(n9295));
  jxor g09030(.dina(n9295), .dinb(n8872), .dout(n9296));
  jand g09031(.dina(asqrt[23] ), .dinb(n8886), .dout(n9297));
  jand g09032(.dina(n9297), .dinb(n8874), .dout(n9298));
  jor  g09033(.dina(n9298), .dinb(n8920), .dout(n9299));
  jor  g09034(.dina(n9299), .dinb(n9296), .dout(n9300));
  jor  g09035(.dina(n9300), .dinb(n9292), .dout(n9301));
  jand g09036(.dina(n9301), .dinb(n194), .dout(n9302));
  jand g09037(.dina(n9296), .dinb(n9292), .dout(n9303));
  jor  g09038(.dina(n9297), .dinb(n8874), .dout(n9304));
  jand g09039(.dina(n8886), .dinb(n8874), .dout(n9305));
  jor  g09040(.dina(n9305), .dinb(n194), .dout(n9306));
  jnot g09041(.din(n9306), .dout(n9307));
  jand g09042(.dina(n9307), .dinb(n9304), .dout(n9308));
  jor  g09043(.dina(n9308), .dinb(n9303), .dout(n9311));
  jor  g09044(.dina(n9311), .dinb(n9302), .dout(asqrt[22] ));
  jxor g09045(.dina(n9066), .dinb(n3371), .dout(n9313));
  jand g09046(.dina(n9313), .dinb(asqrt[22] ), .dout(n9314));
  jxor g09047(.dina(n9314), .dinb(n8901), .dout(n9315));
  jnot g09048(.din(n9315), .dout(n9316));
  jand g09049(.dina(asqrt[22] ), .dinb(a[44] ), .dout(n9317));
  jnot g09050(.din(a[42] ), .dout(n9318));
  jnot g09051(.din(a[43] ), .dout(n9319));
  jand g09052(.dina(n8903), .dinb(n9319), .dout(n9320));
  jand g09053(.dina(n9320), .dinb(n9318), .dout(n9321));
  jor  g09054(.dina(n9321), .dinb(n9317), .dout(n9322));
  jand g09055(.dina(n9322), .dinb(asqrt[23] ), .dout(n9323));
  jand g09056(.dina(asqrt[22] ), .dinb(n8903), .dout(n9324));
  jxor g09057(.dina(n9324), .dinb(n8904), .dout(n9325));
  jor  g09058(.dina(n9322), .dinb(asqrt[23] ), .dout(n9326));
  jand g09059(.dina(n9326), .dinb(n9325), .dout(n9327));
  jor  g09060(.dina(n9327), .dinb(n9323), .dout(n9328));
  jand g09061(.dina(n9328), .dinb(asqrt[24] ), .dout(n9329));
  jor  g09062(.dina(n9323), .dinb(asqrt[24] ), .dout(n9330));
  jor  g09063(.dina(n9330), .dinb(n9327), .dout(n9331));
  jand g09064(.dina(n9324), .dinb(n8904), .dout(n9332));
  jnot g09065(.din(n9302), .dout(n9333));
  jnot g09066(.din(n9303), .dout(n9334));
  jnot g09067(.din(n9308), .dout(n9335));
  jand g09068(.dina(n9335), .dinb(asqrt[23] ), .dout(n9336));
  jand g09069(.dina(n9336), .dinb(n9334), .dout(n9337));
  jand g09070(.dina(n9337), .dinb(n9333), .dout(n9338));
  jor  g09071(.dina(n9338), .dinb(n9332), .dout(n9339));
  jxor g09072(.dina(n9339), .dinb(n8460), .dout(n9340));
  jand g09073(.dina(n9340), .dinb(n9331), .dout(n9341));
  jor  g09074(.dina(n9341), .dinb(n9329), .dout(n9342));
  jand g09075(.dina(n9342), .dinb(asqrt[25] ), .dout(n9343));
  jor  g09076(.dina(n9342), .dinb(asqrt[25] ), .dout(n9344));
  jxor g09077(.dina(n8908), .dinb(n8893), .dout(n9345));
  jand g09078(.dina(n9345), .dinb(asqrt[22] ), .dout(n9346));
  jxor g09079(.dina(n9346), .dinb(n8911), .dout(n9347));
  jnot g09080(.din(n9347), .dout(n9348));
  jand g09081(.dina(n9348), .dinb(n9344), .dout(n9349));
  jor  g09082(.dina(n9349), .dinb(n9343), .dout(n9350));
  jand g09083(.dina(n9350), .dinb(asqrt[26] ), .dout(n9351));
  jnot g09084(.din(n8917), .dout(n9352));
  jand g09085(.dina(n9352), .dinb(n8915), .dout(n9353));
  jand g09086(.dina(n9353), .dinb(asqrt[22] ), .dout(n9354));
  jxor g09087(.dina(n9354), .dinb(n8925), .dout(n9355));
  jnot g09088(.din(n9355), .dout(n9356));
  jor  g09089(.dina(n9343), .dinb(asqrt[26] ), .dout(n9357));
  jor  g09090(.dina(n9357), .dinb(n9349), .dout(n9358));
  jand g09091(.dina(n9358), .dinb(n9356), .dout(n9359));
  jor  g09092(.dina(n9359), .dinb(n9351), .dout(n9360));
  jand g09093(.dina(n9360), .dinb(asqrt[27] ), .dout(n9361));
  jor  g09094(.dina(n9360), .dinb(asqrt[27] ), .dout(n9362));
  jnot g09095(.din(n8932), .dout(n9363));
  jxor g09096(.dina(n8927), .dinb(n8053), .dout(n9364));
  jand g09097(.dina(n9364), .dinb(asqrt[22] ), .dout(n9365));
  jxor g09098(.dina(n9365), .dinb(n9363), .dout(n9366));
  jand g09099(.dina(n9366), .dinb(n9362), .dout(n9367));
  jor  g09100(.dina(n9367), .dinb(n9361), .dout(n9368));
  jand g09101(.dina(n9368), .dinb(asqrt[28] ), .dout(n9369));
  jor  g09102(.dina(n9361), .dinb(asqrt[28] ), .dout(n9370));
  jor  g09103(.dina(n9370), .dinb(n9367), .dout(n9371));
  jnot g09104(.din(n8939), .dout(n9372));
  jnot g09105(.din(n8941), .dout(n9373));
  jand g09106(.dina(asqrt[22] ), .dinb(n8935), .dout(n9374));
  jand g09107(.dina(n9374), .dinb(n9373), .dout(n9375));
  jor  g09108(.dina(n9375), .dinb(n9372), .dout(n9376));
  jnot g09109(.din(n8942), .dout(n9377));
  jand g09110(.dina(n9374), .dinb(n9377), .dout(n9378));
  jnot g09111(.din(n9378), .dout(n9379));
  jand g09112(.dina(n9379), .dinb(n9376), .dout(n9380));
  jand g09113(.dina(n9380), .dinb(n9371), .dout(n9381));
  jor  g09114(.dina(n9381), .dinb(n9369), .dout(n9382));
  jand g09115(.dina(n9382), .dinb(asqrt[29] ), .dout(n9383));
  jor  g09116(.dina(n9382), .dinb(asqrt[29] ), .dout(n9384));
  jxor g09117(.dina(n8943), .dinb(n7260), .dout(n9385));
  jand g09118(.dina(n9385), .dinb(asqrt[22] ), .dout(n9386));
  jxor g09119(.dina(n9386), .dinb(n8948), .dout(n9387));
  jand g09120(.dina(n9387), .dinb(n9384), .dout(n9388));
  jor  g09121(.dina(n9388), .dinb(n9383), .dout(n9389));
  jand g09122(.dina(n9389), .dinb(asqrt[30] ), .dout(n9390));
  jnot g09123(.din(n8954), .dout(n9391));
  jand g09124(.dina(n9391), .dinb(n8952), .dout(n9392));
  jand g09125(.dina(n9392), .dinb(asqrt[22] ), .dout(n9393));
  jxor g09126(.dina(n9393), .dinb(n8963), .dout(n9394));
  jnot g09127(.din(n9394), .dout(n9395));
  jor  g09128(.dina(n9383), .dinb(asqrt[30] ), .dout(n9396));
  jor  g09129(.dina(n9396), .dinb(n9388), .dout(n9397));
  jand g09130(.dina(n9397), .dinb(n9395), .dout(n9398));
  jor  g09131(.dina(n9398), .dinb(n9390), .dout(n9399));
  jand g09132(.dina(n9399), .dinb(asqrt[31] ), .dout(n9400));
  jor  g09133(.dina(n9399), .dinb(asqrt[31] ), .dout(n9401));
  jxor g09134(.dina(n8965), .dinb(n6500), .dout(n9402));
  jand g09135(.dina(n9402), .dinb(asqrt[22] ), .dout(n9403));
  jxor g09136(.dina(n9403), .dinb(n8971), .dout(n9404));
  jand g09137(.dina(n9404), .dinb(n9401), .dout(n9405));
  jor  g09138(.dina(n9405), .dinb(n9400), .dout(n9406));
  jand g09139(.dina(n9406), .dinb(asqrt[32] ), .dout(n9407));
  jor  g09140(.dina(n9400), .dinb(asqrt[32] ), .dout(n9408));
  jor  g09141(.dina(n9408), .dinb(n9405), .dout(n9409));
  jnot g09142(.din(n8979), .dout(n9410));
  jnot g09143(.din(n8981), .dout(n9411));
  jand g09144(.dina(asqrt[22] ), .dinb(n8975), .dout(n9412));
  jand g09145(.dina(n9412), .dinb(n9411), .dout(n9413));
  jor  g09146(.dina(n9413), .dinb(n9410), .dout(n9414));
  jnot g09147(.din(n8982), .dout(n9415));
  jand g09148(.dina(n9412), .dinb(n9415), .dout(n9416));
  jnot g09149(.din(n9416), .dout(n9417));
  jand g09150(.dina(n9417), .dinb(n9414), .dout(n9418));
  jand g09151(.dina(n9418), .dinb(n9409), .dout(n9419));
  jor  g09152(.dina(n9419), .dinb(n9407), .dout(n9420));
  jand g09153(.dina(n9420), .dinb(asqrt[33] ), .dout(n9421));
  jxor g09154(.dina(n8983), .dinb(n5788), .dout(n9422));
  jand g09155(.dina(n9422), .dinb(asqrt[22] ), .dout(n9423));
  jxor g09156(.dina(n9423), .dinb(n8990), .dout(n9424));
  jnot g09157(.din(n9424), .dout(n9425));
  jor  g09158(.dina(n9420), .dinb(asqrt[33] ), .dout(n9426));
  jand g09159(.dina(n9426), .dinb(n9425), .dout(n9427));
  jor  g09160(.dina(n9427), .dinb(n9421), .dout(n9428));
  jand g09161(.dina(n9428), .dinb(asqrt[34] ), .dout(n9429));
  jnot g09162(.din(n8995), .dout(n9430));
  jand g09163(.dina(n9430), .dinb(n8993), .dout(n9431));
  jand g09164(.dina(n9431), .dinb(asqrt[22] ), .dout(n9432));
  jxor g09165(.dina(n9432), .dinb(n9003), .dout(n9433));
  jnot g09166(.din(n9433), .dout(n9434));
  jor  g09167(.dina(n9421), .dinb(asqrt[34] ), .dout(n9435));
  jor  g09168(.dina(n9435), .dinb(n9427), .dout(n9436));
  jand g09169(.dina(n9436), .dinb(n9434), .dout(n9437));
  jor  g09170(.dina(n9437), .dinb(n9429), .dout(n9438));
  jand g09171(.dina(n9438), .dinb(asqrt[35] ), .dout(n9439));
  jor  g09172(.dina(n9438), .dinb(asqrt[35] ), .dout(n9440));
  jnot g09173(.din(n9009), .dout(n9441));
  jnot g09174(.din(n9010), .dout(n9442));
  jand g09175(.dina(asqrt[22] ), .dinb(n9006), .dout(n9443));
  jand g09176(.dina(n9443), .dinb(n9442), .dout(n9444));
  jor  g09177(.dina(n9444), .dinb(n9441), .dout(n9445));
  jnot g09178(.din(n9011), .dout(n9446));
  jand g09179(.dina(n9443), .dinb(n9446), .dout(n9447));
  jnot g09180(.din(n9447), .dout(n9448));
  jand g09181(.dina(n9448), .dinb(n9445), .dout(n9449));
  jand g09182(.dina(n9449), .dinb(n9440), .dout(n9450));
  jor  g09183(.dina(n9450), .dinb(n9439), .dout(n9451));
  jand g09184(.dina(n9451), .dinb(asqrt[36] ), .dout(n9452));
  jor  g09185(.dina(n9439), .dinb(asqrt[36] ), .dout(n9453));
  jor  g09186(.dina(n9453), .dinb(n9450), .dout(n9454));
  jnot g09187(.din(n9017), .dout(n9455));
  jnot g09188(.din(n9019), .dout(n9456));
  jand g09189(.dina(asqrt[22] ), .dinb(n9013), .dout(n9457));
  jand g09190(.dina(n9457), .dinb(n9456), .dout(n9458));
  jor  g09191(.dina(n9458), .dinb(n9455), .dout(n9459));
  jnot g09192(.din(n9020), .dout(n9460));
  jand g09193(.dina(n9457), .dinb(n9460), .dout(n9461));
  jnot g09194(.din(n9461), .dout(n9462));
  jand g09195(.dina(n9462), .dinb(n9459), .dout(n9463));
  jand g09196(.dina(n9463), .dinb(n9454), .dout(n9464));
  jor  g09197(.dina(n9464), .dinb(n9452), .dout(n9465));
  jand g09198(.dina(n9465), .dinb(asqrt[37] ), .dout(n9466));
  jxor g09199(.dina(n9021), .dinb(n4494), .dout(n9467));
  jand g09200(.dina(n9467), .dinb(asqrt[22] ), .dout(n9468));
  jxor g09201(.dina(n9468), .dinb(n9031), .dout(n9469));
  jnot g09202(.din(n9469), .dout(n9470));
  jor  g09203(.dina(n9465), .dinb(asqrt[37] ), .dout(n9471));
  jand g09204(.dina(n9471), .dinb(n9470), .dout(n9472));
  jor  g09205(.dina(n9472), .dinb(n9466), .dout(n9473));
  jand g09206(.dina(n9473), .dinb(asqrt[38] ), .dout(n9474));
  jnot g09207(.din(n9036), .dout(n9475));
  jand g09208(.dina(n9475), .dinb(n9034), .dout(n9476));
  jand g09209(.dina(n9476), .dinb(asqrt[22] ), .dout(n9477));
  jxor g09210(.dina(n9477), .dinb(n9044), .dout(n9478));
  jnot g09211(.din(n9478), .dout(n9479));
  jor  g09212(.dina(n9466), .dinb(asqrt[38] ), .dout(n9480));
  jor  g09213(.dina(n9480), .dinb(n9472), .dout(n9481));
  jand g09214(.dina(n9481), .dinb(n9479), .dout(n9482));
  jor  g09215(.dina(n9482), .dinb(n9474), .dout(n9483));
  jand g09216(.dina(n9483), .dinb(asqrt[39] ), .dout(n9484));
  jor  g09217(.dina(n9483), .dinb(asqrt[39] ), .dout(n9485));
  jnot g09218(.din(n9050), .dout(n9486));
  jnot g09219(.din(n9051), .dout(n9487));
  jand g09220(.dina(asqrt[22] ), .dinb(n9047), .dout(n9488));
  jand g09221(.dina(n9488), .dinb(n9487), .dout(n9489));
  jor  g09222(.dina(n9489), .dinb(n9486), .dout(n9490));
  jnot g09223(.din(n9052), .dout(n9491));
  jand g09224(.dina(n9488), .dinb(n9491), .dout(n9492));
  jnot g09225(.din(n9492), .dout(n9493));
  jand g09226(.dina(n9493), .dinb(n9490), .dout(n9494));
  jand g09227(.dina(n9494), .dinb(n9485), .dout(n9495));
  jor  g09228(.dina(n9495), .dinb(n9484), .dout(n9496));
  jand g09229(.dina(n9496), .dinb(asqrt[40] ), .dout(n9497));
  jnot g09230(.din(n9056), .dout(n9498));
  jand g09231(.dina(n9498), .dinb(n9054), .dout(n9499));
  jand g09232(.dina(n9499), .dinb(asqrt[22] ), .dout(n9500));
  jxor g09233(.dina(n9500), .dinb(n9064), .dout(n9501));
  jnot g09234(.din(n9501), .dout(n9502));
  jor  g09235(.dina(n9484), .dinb(asqrt[40] ), .dout(n9503));
  jor  g09236(.dina(n9503), .dinb(n9495), .dout(n9504));
  jand g09237(.dina(n9504), .dinb(n9502), .dout(n9505));
  jor  g09238(.dina(n9505), .dinb(n9497), .dout(n9506));
  jand g09239(.dina(n9506), .dinb(asqrt[41] ), .dout(n9507));
  jor  g09240(.dina(n9506), .dinb(asqrt[41] ), .dout(n9508));
  jand g09241(.dina(n9508), .dinb(n9315), .dout(n9509));
  jor  g09242(.dina(n9509), .dinb(n9507), .dout(n9510));
  jand g09243(.dina(n9510), .dinb(asqrt[42] ), .dout(n9511));
  jor  g09244(.dina(n9507), .dinb(asqrt[42] ), .dout(n9512));
  jor  g09245(.dina(n9512), .dinb(n9509), .dout(n9513));
  jnot g09246(.din(n9076), .dout(n9514));
  jnot g09247(.din(n9078), .dout(n9515));
  jand g09248(.dina(asqrt[22] ), .dinb(n9072), .dout(n9516));
  jand g09249(.dina(n9516), .dinb(n9515), .dout(n9517));
  jor  g09250(.dina(n9517), .dinb(n9514), .dout(n9518));
  jnot g09251(.din(n9079), .dout(n9519));
  jand g09252(.dina(n9516), .dinb(n9519), .dout(n9520));
  jnot g09253(.din(n9520), .dout(n9521));
  jand g09254(.dina(n9521), .dinb(n9518), .dout(n9522));
  jand g09255(.dina(n9522), .dinb(n9513), .dout(n9523));
  jor  g09256(.dina(n9523), .dinb(n9511), .dout(n9524));
  jand g09257(.dina(n9524), .dinb(asqrt[43] ), .dout(n9525));
  jor  g09258(.dina(n9524), .dinb(asqrt[43] ), .dout(n9526));
  jnot g09259(.din(n9084), .dout(n9527));
  jnot g09260(.din(n9085), .dout(n9528));
  jand g09261(.dina(asqrt[22] ), .dinb(n9081), .dout(n9529));
  jand g09262(.dina(n9529), .dinb(n9528), .dout(n9530));
  jor  g09263(.dina(n9530), .dinb(n9527), .dout(n9531));
  jnot g09264(.din(n9086), .dout(n9532));
  jand g09265(.dina(n9529), .dinb(n9532), .dout(n9533));
  jnot g09266(.din(n9533), .dout(n9534));
  jand g09267(.dina(n9534), .dinb(n9531), .dout(n9535));
  jand g09268(.dina(n9535), .dinb(n9526), .dout(n9536));
  jor  g09269(.dina(n9536), .dinb(n9525), .dout(n9537));
  jand g09270(.dina(n9537), .dinb(asqrt[44] ), .dout(n9538));
  jor  g09271(.dina(n9525), .dinb(asqrt[44] ), .dout(n9539));
  jor  g09272(.dina(n9539), .dinb(n9536), .dout(n9540));
  jnot g09273(.din(n9092), .dout(n9541));
  jnot g09274(.din(n9094), .dout(n9542));
  jand g09275(.dina(asqrt[22] ), .dinb(n9088), .dout(n9543));
  jand g09276(.dina(n9543), .dinb(n9542), .dout(n9544));
  jor  g09277(.dina(n9544), .dinb(n9541), .dout(n9545));
  jnot g09278(.din(n9095), .dout(n9546));
  jand g09279(.dina(n9543), .dinb(n9546), .dout(n9547));
  jnot g09280(.din(n9547), .dout(n9548));
  jand g09281(.dina(n9548), .dinb(n9545), .dout(n9549));
  jand g09282(.dina(n9549), .dinb(n9540), .dout(n9550));
  jor  g09283(.dina(n9550), .dinb(n9538), .dout(n9551));
  jand g09284(.dina(n9551), .dinb(asqrt[45] ), .dout(n9552));
  jxor g09285(.dina(n9096), .dinb(n2420), .dout(n9553));
  jand g09286(.dina(n9553), .dinb(asqrt[22] ), .dout(n9554));
  jxor g09287(.dina(n9554), .dinb(n9106), .dout(n9555));
  jnot g09288(.din(n9555), .dout(n9556));
  jor  g09289(.dina(n9551), .dinb(asqrt[45] ), .dout(n9557));
  jand g09290(.dina(n9557), .dinb(n9556), .dout(n9558));
  jor  g09291(.dina(n9558), .dinb(n9552), .dout(n9559));
  jand g09292(.dina(n9559), .dinb(asqrt[46] ), .dout(n9560));
  jnot g09293(.din(n9111), .dout(n9561));
  jand g09294(.dina(n9561), .dinb(n9109), .dout(n9562));
  jand g09295(.dina(n9562), .dinb(asqrt[22] ), .dout(n9563));
  jxor g09296(.dina(n9563), .dinb(n9119), .dout(n9564));
  jnot g09297(.din(n9564), .dout(n9565));
  jor  g09298(.dina(n9552), .dinb(asqrt[46] ), .dout(n9566));
  jor  g09299(.dina(n9566), .dinb(n9558), .dout(n9567));
  jand g09300(.dina(n9567), .dinb(n9565), .dout(n9568));
  jor  g09301(.dina(n9568), .dinb(n9560), .dout(n9569));
  jand g09302(.dina(n9569), .dinb(asqrt[47] ), .dout(n9570));
  jor  g09303(.dina(n9569), .dinb(asqrt[47] ), .dout(n9571));
  jnot g09304(.din(n9125), .dout(n9572));
  jnot g09305(.din(n9126), .dout(n9573));
  jand g09306(.dina(asqrt[22] ), .dinb(n9122), .dout(n9574));
  jand g09307(.dina(n9574), .dinb(n9573), .dout(n9575));
  jor  g09308(.dina(n9575), .dinb(n9572), .dout(n9576));
  jnot g09309(.din(n9127), .dout(n9577));
  jand g09310(.dina(n9574), .dinb(n9577), .dout(n9578));
  jnot g09311(.din(n9578), .dout(n9579));
  jand g09312(.dina(n9579), .dinb(n9576), .dout(n9580));
  jand g09313(.dina(n9580), .dinb(n9571), .dout(n9581));
  jor  g09314(.dina(n9581), .dinb(n9570), .dout(n9582));
  jand g09315(.dina(n9582), .dinb(asqrt[48] ), .dout(n9583));
  jor  g09316(.dina(n9570), .dinb(asqrt[48] ), .dout(n9584));
  jor  g09317(.dina(n9584), .dinb(n9581), .dout(n9585));
  jnot g09318(.din(n9133), .dout(n9586));
  jnot g09319(.din(n9135), .dout(n9587));
  jand g09320(.dina(asqrt[22] ), .dinb(n9129), .dout(n9588));
  jand g09321(.dina(n9588), .dinb(n9587), .dout(n9589));
  jor  g09322(.dina(n9589), .dinb(n9586), .dout(n9590));
  jnot g09323(.din(n9136), .dout(n9591));
  jand g09324(.dina(n9588), .dinb(n9591), .dout(n9592));
  jnot g09325(.din(n9592), .dout(n9593));
  jand g09326(.dina(n9593), .dinb(n9590), .dout(n9594));
  jand g09327(.dina(n9594), .dinb(n9585), .dout(n9595));
  jor  g09328(.dina(n9595), .dinb(n9583), .dout(n9596));
  jand g09329(.dina(n9596), .dinb(asqrt[49] ), .dout(n9597));
  jxor g09330(.dina(n9137), .dinb(n1641), .dout(n9598));
  jand g09331(.dina(n9598), .dinb(asqrt[22] ), .dout(n9599));
  jxor g09332(.dina(n9599), .dinb(n9147), .dout(n9600));
  jnot g09333(.din(n9600), .dout(n9601));
  jor  g09334(.dina(n9596), .dinb(asqrt[49] ), .dout(n9602));
  jand g09335(.dina(n9602), .dinb(n9601), .dout(n9603));
  jor  g09336(.dina(n9603), .dinb(n9597), .dout(n9604));
  jand g09337(.dina(n9604), .dinb(asqrt[50] ), .dout(n9605));
  jnot g09338(.din(n9152), .dout(n9606));
  jand g09339(.dina(n9606), .dinb(n9150), .dout(n9607));
  jand g09340(.dina(n9607), .dinb(asqrt[22] ), .dout(n9608));
  jxor g09341(.dina(n9608), .dinb(n9160), .dout(n9609));
  jnot g09342(.din(n9609), .dout(n9610));
  jor  g09343(.dina(n9597), .dinb(asqrt[50] ), .dout(n9611));
  jor  g09344(.dina(n9611), .dinb(n9603), .dout(n9612));
  jand g09345(.dina(n9612), .dinb(n9610), .dout(n9613));
  jor  g09346(.dina(n9613), .dinb(n9605), .dout(n9614));
  jand g09347(.dina(n9614), .dinb(asqrt[51] ), .dout(n9615));
  jor  g09348(.dina(n9614), .dinb(asqrt[51] ), .dout(n9616));
  jnot g09349(.din(n9166), .dout(n9617));
  jnot g09350(.din(n9167), .dout(n9618));
  jand g09351(.dina(asqrt[22] ), .dinb(n9163), .dout(n9619));
  jand g09352(.dina(n9619), .dinb(n9618), .dout(n9620));
  jor  g09353(.dina(n9620), .dinb(n9617), .dout(n9621));
  jnot g09354(.din(n9168), .dout(n9622));
  jand g09355(.dina(n9619), .dinb(n9622), .dout(n9623));
  jnot g09356(.din(n9623), .dout(n9624));
  jand g09357(.dina(n9624), .dinb(n9621), .dout(n9625));
  jand g09358(.dina(n9625), .dinb(n9616), .dout(n9626));
  jor  g09359(.dina(n9626), .dinb(n9615), .dout(n9627));
  jand g09360(.dina(n9627), .dinb(asqrt[52] ), .dout(n9628));
  jor  g09361(.dina(n9615), .dinb(asqrt[52] ), .dout(n9629));
  jor  g09362(.dina(n9629), .dinb(n9626), .dout(n9630));
  jnot g09363(.din(n9174), .dout(n9631));
  jnot g09364(.din(n9176), .dout(n9632));
  jand g09365(.dina(asqrt[22] ), .dinb(n9170), .dout(n9633));
  jand g09366(.dina(n9633), .dinb(n9632), .dout(n9634));
  jor  g09367(.dina(n9634), .dinb(n9631), .dout(n9635));
  jnot g09368(.din(n9177), .dout(n9636));
  jand g09369(.dina(n9633), .dinb(n9636), .dout(n9637));
  jnot g09370(.din(n9637), .dout(n9638));
  jand g09371(.dina(n9638), .dinb(n9635), .dout(n9639));
  jand g09372(.dina(n9639), .dinb(n9630), .dout(n9640));
  jor  g09373(.dina(n9640), .dinb(n9628), .dout(n9641));
  jand g09374(.dina(n9641), .dinb(asqrt[53] ), .dout(n9642));
  jxor g09375(.dina(n9178), .dinb(n1034), .dout(n9643));
  jand g09376(.dina(n9643), .dinb(asqrt[22] ), .dout(n9644));
  jxor g09377(.dina(n9644), .dinb(n9188), .dout(n9645));
  jnot g09378(.din(n9645), .dout(n9646));
  jor  g09379(.dina(n9641), .dinb(asqrt[53] ), .dout(n9647));
  jand g09380(.dina(n9647), .dinb(n9646), .dout(n9648));
  jor  g09381(.dina(n9648), .dinb(n9642), .dout(n9649));
  jand g09382(.dina(n9649), .dinb(asqrt[54] ), .dout(n9650));
  jnot g09383(.din(n9193), .dout(n9651));
  jand g09384(.dina(n9651), .dinb(n9191), .dout(n9652));
  jand g09385(.dina(n9652), .dinb(asqrt[22] ), .dout(n9653));
  jxor g09386(.dina(n9653), .dinb(n9201), .dout(n9654));
  jnot g09387(.din(n9654), .dout(n9655));
  jor  g09388(.dina(n9642), .dinb(asqrt[54] ), .dout(n9656));
  jor  g09389(.dina(n9656), .dinb(n9648), .dout(n9657));
  jand g09390(.dina(n9657), .dinb(n9655), .dout(n9658));
  jor  g09391(.dina(n9658), .dinb(n9650), .dout(n9659));
  jand g09392(.dina(n9659), .dinb(asqrt[55] ), .dout(n9660));
  jor  g09393(.dina(n9659), .dinb(asqrt[55] ), .dout(n9661));
  jnot g09394(.din(n9207), .dout(n9662));
  jnot g09395(.din(n9208), .dout(n9663));
  jand g09396(.dina(asqrt[22] ), .dinb(n9204), .dout(n9664));
  jand g09397(.dina(n9664), .dinb(n9663), .dout(n9665));
  jor  g09398(.dina(n9665), .dinb(n9662), .dout(n9666));
  jnot g09399(.din(n9209), .dout(n9667));
  jand g09400(.dina(n9664), .dinb(n9667), .dout(n9668));
  jnot g09401(.din(n9668), .dout(n9669));
  jand g09402(.dina(n9669), .dinb(n9666), .dout(n9670));
  jand g09403(.dina(n9670), .dinb(n9661), .dout(n9671));
  jor  g09404(.dina(n9671), .dinb(n9660), .dout(n9672));
  jand g09405(.dina(n9672), .dinb(asqrt[56] ), .dout(n9673));
  jor  g09406(.dina(n9660), .dinb(asqrt[56] ), .dout(n9674));
  jor  g09407(.dina(n9674), .dinb(n9671), .dout(n9675));
  jnot g09408(.din(n9215), .dout(n9676));
  jnot g09409(.din(n9217), .dout(n9677));
  jand g09410(.dina(asqrt[22] ), .dinb(n9211), .dout(n9678));
  jand g09411(.dina(n9678), .dinb(n9677), .dout(n9679));
  jor  g09412(.dina(n9679), .dinb(n9676), .dout(n9680));
  jnot g09413(.din(n9218), .dout(n9681));
  jand g09414(.dina(n9678), .dinb(n9681), .dout(n9682));
  jnot g09415(.din(n9682), .dout(n9683));
  jand g09416(.dina(n9683), .dinb(n9680), .dout(n9684));
  jand g09417(.dina(n9684), .dinb(n9675), .dout(n9685));
  jor  g09418(.dina(n9685), .dinb(n9673), .dout(n9686));
  jand g09419(.dina(n9686), .dinb(asqrt[57] ), .dout(n9687));
  jxor g09420(.dina(n9219), .dinb(n590), .dout(n9688));
  jand g09421(.dina(n9688), .dinb(asqrt[22] ), .dout(n9689));
  jxor g09422(.dina(n9689), .dinb(n9229), .dout(n9690));
  jnot g09423(.din(n9690), .dout(n9691));
  jor  g09424(.dina(n9686), .dinb(asqrt[57] ), .dout(n9692));
  jand g09425(.dina(n9692), .dinb(n9691), .dout(n9693));
  jor  g09426(.dina(n9693), .dinb(n9687), .dout(n9694));
  jand g09427(.dina(n9694), .dinb(asqrt[58] ), .dout(n9695));
  jnot g09428(.din(n9234), .dout(n9696));
  jand g09429(.dina(n9696), .dinb(n9232), .dout(n9697));
  jand g09430(.dina(n9697), .dinb(asqrt[22] ), .dout(n9698));
  jxor g09431(.dina(n9698), .dinb(n9242), .dout(n9699));
  jnot g09432(.din(n9699), .dout(n9700));
  jor  g09433(.dina(n9687), .dinb(asqrt[58] ), .dout(n9701));
  jor  g09434(.dina(n9701), .dinb(n9693), .dout(n9702));
  jand g09435(.dina(n9702), .dinb(n9700), .dout(n9703));
  jor  g09436(.dina(n9703), .dinb(n9695), .dout(n9704));
  jand g09437(.dina(n9704), .dinb(asqrt[59] ), .dout(n9705));
  jor  g09438(.dina(n9704), .dinb(asqrt[59] ), .dout(n9706));
  jnot g09439(.din(n9248), .dout(n9707));
  jnot g09440(.din(n9249), .dout(n9708));
  jand g09441(.dina(asqrt[22] ), .dinb(n9245), .dout(n9709));
  jand g09442(.dina(n9709), .dinb(n9708), .dout(n9710));
  jor  g09443(.dina(n9710), .dinb(n9707), .dout(n9711));
  jnot g09444(.din(n9250), .dout(n9712));
  jand g09445(.dina(n9709), .dinb(n9712), .dout(n9713));
  jnot g09446(.din(n9713), .dout(n9714));
  jand g09447(.dina(n9714), .dinb(n9711), .dout(n9715));
  jand g09448(.dina(n9715), .dinb(n9706), .dout(n9716));
  jor  g09449(.dina(n9716), .dinb(n9705), .dout(n9717));
  jand g09450(.dina(n9717), .dinb(asqrt[60] ), .dout(n9718));
  jor  g09451(.dina(n9705), .dinb(asqrt[60] ), .dout(n9719));
  jor  g09452(.dina(n9719), .dinb(n9716), .dout(n9720));
  jnot g09453(.din(n9256), .dout(n9721));
  jnot g09454(.din(n9258), .dout(n9722));
  jand g09455(.dina(asqrt[22] ), .dinb(n9252), .dout(n9723));
  jand g09456(.dina(n9723), .dinb(n9722), .dout(n9724));
  jor  g09457(.dina(n9724), .dinb(n9721), .dout(n9725));
  jnot g09458(.din(n9259), .dout(n9726));
  jand g09459(.dina(n9723), .dinb(n9726), .dout(n9727));
  jnot g09460(.din(n9727), .dout(n9728));
  jand g09461(.dina(n9728), .dinb(n9725), .dout(n9729));
  jand g09462(.dina(n9729), .dinb(n9720), .dout(n9730));
  jor  g09463(.dina(n9730), .dinb(n9718), .dout(n9731));
  jand g09464(.dina(n9731), .dinb(asqrt[61] ), .dout(n9732));
  jxor g09465(.dina(n9260), .dinb(n290), .dout(n9733));
  jand g09466(.dina(n9733), .dinb(asqrt[22] ), .dout(n9734));
  jxor g09467(.dina(n9734), .dinb(n9270), .dout(n9735));
  jnot g09468(.din(n9735), .dout(n9736));
  jor  g09469(.dina(n9731), .dinb(asqrt[61] ), .dout(n9737));
  jand g09470(.dina(n9737), .dinb(n9736), .dout(n9738));
  jor  g09471(.dina(n9738), .dinb(n9732), .dout(n9739));
  jand g09472(.dina(n9739), .dinb(asqrt[62] ), .dout(n9740));
  jnot g09473(.din(n9275), .dout(n9741));
  jand g09474(.dina(n9741), .dinb(n9273), .dout(n9742));
  jand g09475(.dina(n9742), .dinb(asqrt[22] ), .dout(n9743));
  jxor g09476(.dina(n9743), .dinb(n9283), .dout(n9744));
  jnot g09477(.din(n9744), .dout(n9745));
  jor  g09478(.dina(n9732), .dinb(asqrt[62] ), .dout(n9746));
  jor  g09479(.dina(n9746), .dinb(n9738), .dout(n9747));
  jand g09480(.dina(n9747), .dinb(n9745), .dout(n9748));
  jor  g09481(.dina(n9748), .dinb(n9740), .dout(n9749));
  jxor g09482(.dina(n9285), .dinb(n199), .dout(n9750));
  jand g09483(.dina(n9750), .dinb(asqrt[22] ), .dout(n9751));
  jxor g09484(.dina(n9751), .dinb(n9290), .dout(n9752));
  jnot g09485(.din(n9292), .dout(n9753));
  jnot g09486(.din(n9296), .dout(n9754));
  jand g09487(.dina(asqrt[22] ), .dinb(n9754), .dout(n9755));
  jand g09488(.dina(n9755), .dinb(n9753), .dout(n9756));
  jor  g09489(.dina(n9756), .dinb(n9303), .dout(n9757));
  jor  g09490(.dina(n9757), .dinb(n9752), .dout(n9758));
  jnot g09491(.din(n9758), .dout(n9759));
  jand g09492(.dina(n9759), .dinb(n9749), .dout(n9760));
  jor  g09493(.dina(n9760), .dinb(asqrt[63] ), .dout(n9761));
  jnot g09494(.din(n9752), .dout(n9762));
  jor  g09495(.dina(n9762), .dinb(n9749), .dout(n9763));
  jor  g09496(.dina(n9755), .dinb(n9753), .dout(n9764));
  jand g09497(.dina(n9754), .dinb(n9753), .dout(n9765));
  jor  g09498(.dina(n9765), .dinb(n194), .dout(n9766));
  jnot g09499(.din(n9766), .dout(n9767));
  jand g09500(.dina(n9767), .dinb(n9764), .dout(n9768));
  jnot g09501(.din(asqrt[22] ), .dout(n9769));
  jnot g09502(.din(n9768), .dout(n9772));
  jand g09503(.dina(n9772), .dinb(n9763), .dout(n9773));
  jand g09504(.dina(n9773), .dinb(n9761), .dout(n9774));
  jxor g09505(.dina(n9506), .dinb(n2875), .dout(n9775));
  jor  g09506(.dina(n9775), .dinb(n9774), .dout(n9776));
  jxor g09507(.dina(n9776), .dinb(n9316), .dout(n9777));
  jnot g09508(.din(n9777), .dout(n9778));
  jor  g09509(.dina(n9774), .dinb(n9318), .dout(n9779));
  jnot g09510(.din(a[40] ), .dout(n9780));
  jnot g09511(.din(a[41] ), .dout(n9781));
  jand g09512(.dina(n9318), .dinb(n9781), .dout(n9782));
  jand g09513(.dina(n9782), .dinb(n9780), .dout(n9783));
  jnot g09514(.din(n9783), .dout(n9784));
  jand g09515(.dina(n9784), .dinb(n9779), .dout(n9785));
  jor  g09516(.dina(n9785), .dinb(n9769), .dout(n9786));
  jor  g09517(.dina(n9774), .dinb(a[42] ), .dout(n9787));
  jxor g09518(.dina(n9787), .dinb(n9319), .dout(n9788));
  jand g09519(.dina(n9785), .dinb(n9769), .dout(n9789));
  jor  g09520(.dina(n9789), .dinb(n9788), .dout(n9790));
  jand g09521(.dina(n9790), .dinb(n9786), .dout(n9791));
  jor  g09522(.dina(n9791), .dinb(n8898), .dout(n9792));
  jand g09523(.dina(n9786), .dinb(n8898), .dout(n9793));
  jand g09524(.dina(n9793), .dinb(n9790), .dout(n9794));
  jor  g09525(.dina(n9787), .dinb(a[43] ), .dout(n9795));
  jnot g09526(.din(n9761), .dout(n9796));
  jnot g09527(.din(n9763), .dout(n9797));
  jor  g09528(.dina(n9768), .dinb(n9769), .dout(n9798));
  jor  g09529(.dina(n9798), .dinb(n9797), .dout(n9799));
  jor  g09530(.dina(n9799), .dinb(n9796), .dout(n9800));
  jand g09531(.dina(n9800), .dinb(n9795), .dout(n9801));
  jxor g09532(.dina(n9801), .dinb(n8903), .dout(n9802));
  jor  g09533(.dina(n9802), .dinb(n9794), .dout(n9803));
  jand g09534(.dina(n9803), .dinb(n9792), .dout(n9804));
  jor  g09535(.dina(n9804), .dinb(n8893), .dout(n9805));
  jand g09536(.dina(n9804), .dinb(n8893), .dout(n9806));
  jxor g09537(.dina(n9322), .dinb(n8898), .dout(n9807));
  jor  g09538(.dina(n9807), .dinb(n9774), .dout(n9808));
  jxor g09539(.dina(n9808), .dinb(n9325), .dout(n9809));
  jor  g09540(.dina(n9809), .dinb(n9806), .dout(n9810));
  jand g09541(.dina(n9810), .dinb(n9805), .dout(n9811));
  jor  g09542(.dina(n9811), .dinb(n8058), .dout(n9812));
  jnot g09543(.din(n9331), .dout(n9813));
  jor  g09544(.dina(n9813), .dinb(n9329), .dout(n9814));
  jor  g09545(.dina(n9814), .dinb(n9774), .dout(n9815));
  jxor g09546(.dina(n9815), .dinb(n9340), .dout(n9816));
  jand g09547(.dina(n9805), .dinb(n8058), .dout(n9817));
  jand g09548(.dina(n9817), .dinb(n9810), .dout(n9818));
  jor  g09549(.dina(n9818), .dinb(n9816), .dout(n9819));
  jand g09550(.dina(n9819), .dinb(n9812), .dout(n9820));
  jor  g09551(.dina(n9820), .dinb(n8053), .dout(n9821));
  jand g09552(.dina(n9820), .dinb(n8053), .dout(n9822));
  jxor g09553(.dina(n9342), .dinb(n8058), .dout(n9823));
  jor  g09554(.dina(n9823), .dinb(n9774), .dout(n9824));
  jxor g09555(.dina(n9824), .dinb(n9347), .dout(n9825));
  jnot g09556(.din(n9825), .dout(n9826));
  jor  g09557(.dina(n9826), .dinb(n9822), .dout(n9827));
  jand g09558(.dina(n9827), .dinb(n9821), .dout(n9828));
  jor  g09559(.dina(n9828), .dinb(n7265), .dout(n9829));
  jand g09560(.dina(n9821), .dinb(n7265), .dout(n9830));
  jand g09561(.dina(n9830), .dinb(n9827), .dout(n9831));
  jnot g09562(.din(n9351), .dout(n9832));
  jnot g09563(.din(n9774), .dout(asqrt[21] ));
  jand g09564(.dina(asqrt[21] ), .dinb(n9832), .dout(n9834));
  jand g09565(.dina(n9834), .dinb(n9358), .dout(n9835));
  jor  g09566(.dina(n9835), .dinb(n9356), .dout(n9836));
  jand g09567(.dina(n9834), .dinb(n9359), .dout(n9837));
  jnot g09568(.din(n9837), .dout(n9838));
  jand g09569(.dina(n9838), .dinb(n9836), .dout(n9839));
  jnot g09570(.din(n9839), .dout(n9840));
  jor  g09571(.dina(n9840), .dinb(n9831), .dout(n9841));
  jand g09572(.dina(n9841), .dinb(n9829), .dout(n9842));
  jor  g09573(.dina(n9842), .dinb(n7260), .dout(n9843));
  jand g09574(.dina(n9842), .dinb(n7260), .dout(n9844));
  jnot g09575(.din(n9366), .dout(n9845));
  jxor g09576(.dina(n9360), .dinb(n7265), .dout(n9846));
  jor  g09577(.dina(n9846), .dinb(n9774), .dout(n9847));
  jxor g09578(.dina(n9847), .dinb(n9845), .dout(n9848));
  jnot g09579(.din(n9848), .dout(n9849));
  jor  g09580(.dina(n9849), .dinb(n9844), .dout(n9850));
  jand g09581(.dina(n9850), .dinb(n9843), .dout(n9851));
  jor  g09582(.dina(n9851), .dinb(n6505), .dout(n9852));
  jnot g09583(.din(n9371), .dout(n9853));
  jor  g09584(.dina(n9853), .dinb(n9369), .dout(n9854));
  jor  g09585(.dina(n9854), .dinb(n9774), .dout(n9855));
  jxor g09586(.dina(n9855), .dinb(n9380), .dout(n9856));
  jand g09587(.dina(n9843), .dinb(n6505), .dout(n9857));
  jand g09588(.dina(n9857), .dinb(n9850), .dout(n9858));
  jor  g09589(.dina(n9858), .dinb(n9856), .dout(n9859));
  jand g09590(.dina(n9859), .dinb(n9852), .dout(n9860));
  jor  g09591(.dina(n9860), .dinb(n6500), .dout(n9861));
  jand g09592(.dina(n9860), .dinb(n6500), .dout(n9862));
  jnot g09593(.din(n9387), .dout(n9863));
  jxor g09594(.dina(n9382), .dinb(n6505), .dout(n9864));
  jor  g09595(.dina(n9864), .dinb(n9774), .dout(n9865));
  jxor g09596(.dina(n9865), .dinb(n9863), .dout(n9866));
  jnot g09597(.din(n9866), .dout(n9867));
  jor  g09598(.dina(n9867), .dinb(n9862), .dout(n9868));
  jand g09599(.dina(n9868), .dinb(n9861), .dout(n9869));
  jor  g09600(.dina(n9869), .dinb(n5793), .dout(n9870));
  jand g09601(.dina(n9861), .dinb(n5793), .dout(n9871));
  jand g09602(.dina(n9871), .dinb(n9868), .dout(n9872));
  jnot g09603(.din(n9390), .dout(n9873));
  jand g09604(.dina(asqrt[21] ), .dinb(n9873), .dout(n9874));
  jand g09605(.dina(n9874), .dinb(n9397), .dout(n9875));
  jor  g09606(.dina(n9875), .dinb(n9395), .dout(n9876));
  jand g09607(.dina(n9874), .dinb(n9398), .dout(n9877));
  jnot g09608(.din(n9877), .dout(n9878));
  jand g09609(.dina(n9878), .dinb(n9876), .dout(n9879));
  jnot g09610(.din(n9879), .dout(n9880));
  jor  g09611(.dina(n9880), .dinb(n9872), .dout(n9881));
  jand g09612(.dina(n9881), .dinb(n9870), .dout(n9882));
  jor  g09613(.dina(n9882), .dinb(n5788), .dout(n9883));
  jxor g09614(.dina(n9399), .dinb(n5793), .dout(n9884));
  jor  g09615(.dina(n9884), .dinb(n9774), .dout(n9885));
  jxor g09616(.dina(n9885), .dinb(n9404), .dout(n9886));
  jand g09617(.dina(n9882), .dinb(n5788), .dout(n9887));
  jor  g09618(.dina(n9887), .dinb(n9886), .dout(n9888));
  jand g09619(.dina(n9888), .dinb(n9883), .dout(n9889));
  jor  g09620(.dina(n9889), .dinb(n5121), .dout(n9890));
  jnot g09621(.din(n9409), .dout(n9891));
  jor  g09622(.dina(n9891), .dinb(n9407), .dout(n9892));
  jor  g09623(.dina(n9892), .dinb(n9774), .dout(n9893));
  jxor g09624(.dina(n9893), .dinb(n9418), .dout(n9894));
  jand g09625(.dina(n9883), .dinb(n5121), .dout(n9895));
  jand g09626(.dina(n9895), .dinb(n9888), .dout(n9896));
  jor  g09627(.dina(n9896), .dinb(n9894), .dout(n9897));
  jand g09628(.dina(n9897), .dinb(n9890), .dout(n9898));
  jor  g09629(.dina(n9898), .dinb(n5116), .dout(n9899));
  jand g09630(.dina(n9898), .dinb(n5116), .dout(n9900));
  jnot g09631(.din(n9421), .dout(n9901));
  jand g09632(.dina(asqrt[21] ), .dinb(n9901), .dout(n9902));
  jand g09633(.dina(n9902), .dinb(n9426), .dout(n9903));
  jor  g09634(.dina(n9903), .dinb(n9425), .dout(n9904));
  jand g09635(.dina(n9902), .dinb(n9427), .dout(n9905));
  jnot g09636(.din(n9905), .dout(n9906));
  jand g09637(.dina(n9906), .dinb(n9904), .dout(n9907));
  jnot g09638(.din(n9907), .dout(n9908));
  jor  g09639(.dina(n9908), .dinb(n9900), .dout(n9909));
  jand g09640(.dina(n9909), .dinb(n9899), .dout(n9910));
  jor  g09641(.dina(n9910), .dinb(n4499), .dout(n9911));
  jand g09642(.dina(n9899), .dinb(n4499), .dout(n9912));
  jand g09643(.dina(n9912), .dinb(n9909), .dout(n9913));
  jnot g09644(.din(n9429), .dout(n9914));
  jand g09645(.dina(asqrt[21] ), .dinb(n9914), .dout(n9915));
  jand g09646(.dina(n9915), .dinb(n9436), .dout(n9916));
  jor  g09647(.dina(n9916), .dinb(n9434), .dout(n9917));
  jand g09648(.dina(n9915), .dinb(n9437), .dout(n9918));
  jnot g09649(.din(n9918), .dout(n9919));
  jand g09650(.dina(n9919), .dinb(n9917), .dout(n9920));
  jnot g09651(.din(n9920), .dout(n9921));
  jor  g09652(.dina(n9921), .dinb(n9913), .dout(n9922));
  jand g09653(.dina(n9922), .dinb(n9911), .dout(n9923));
  jor  g09654(.dina(n9923), .dinb(n4494), .dout(n9924));
  jxor g09655(.dina(n9438), .dinb(n4499), .dout(n9925));
  jor  g09656(.dina(n9925), .dinb(n9774), .dout(n9926));
  jxor g09657(.dina(n9926), .dinb(n9449), .dout(n9927));
  jand g09658(.dina(n9923), .dinb(n4494), .dout(n9928));
  jor  g09659(.dina(n9928), .dinb(n9927), .dout(n9929));
  jand g09660(.dina(n9929), .dinb(n9924), .dout(n9930));
  jor  g09661(.dina(n9930), .dinb(n3912), .dout(n9931));
  jnot g09662(.din(n9454), .dout(n9932));
  jor  g09663(.dina(n9932), .dinb(n9452), .dout(n9933));
  jor  g09664(.dina(n9933), .dinb(n9774), .dout(n9934));
  jxor g09665(.dina(n9934), .dinb(n9463), .dout(n9935));
  jand g09666(.dina(n9924), .dinb(n3912), .dout(n9936));
  jand g09667(.dina(n9936), .dinb(n9929), .dout(n9937));
  jor  g09668(.dina(n9937), .dinb(n9935), .dout(n9938));
  jand g09669(.dina(n9938), .dinb(n9931), .dout(n9939));
  jor  g09670(.dina(n9939), .dinb(n3907), .dout(n9940));
  jand g09671(.dina(n9939), .dinb(n3907), .dout(n9941));
  jnot g09672(.din(n9466), .dout(n9942));
  jand g09673(.dina(asqrt[21] ), .dinb(n9942), .dout(n9943));
  jand g09674(.dina(n9943), .dinb(n9471), .dout(n9944));
  jor  g09675(.dina(n9944), .dinb(n9470), .dout(n9945));
  jand g09676(.dina(n9943), .dinb(n9472), .dout(n9946));
  jnot g09677(.din(n9946), .dout(n9947));
  jand g09678(.dina(n9947), .dinb(n9945), .dout(n9948));
  jnot g09679(.din(n9948), .dout(n9949));
  jor  g09680(.dina(n9949), .dinb(n9941), .dout(n9950));
  jand g09681(.dina(n9950), .dinb(n9940), .dout(n9951));
  jor  g09682(.dina(n9951), .dinb(n3376), .dout(n9952));
  jand g09683(.dina(n9940), .dinb(n3376), .dout(n9953));
  jand g09684(.dina(n9953), .dinb(n9950), .dout(n9954));
  jnot g09685(.din(n9474), .dout(n9955));
  jand g09686(.dina(asqrt[21] ), .dinb(n9955), .dout(n9956));
  jand g09687(.dina(n9956), .dinb(n9481), .dout(n9957));
  jor  g09688(.dina(n9957), .dinb(n9479), .dout(n9958));
  jand g09689(.dina(n9956), .dinb(n9482), .dout(n9959));
  jnot g09690(.din(n9959), .dout(n9960));
  jand g09691(.dina(n9960), .dinb(n9958), .dout(n9961));
  jnot g09692(.din(n9961), .dout(n9962));
  jor  g09693(.dina(n9962), .dinb(n9954), .dout(n9963));
  jand g09694(.dina(n9963), .dinb(n9952), .dout(n9964));
  jor  g09695(.dina(n9964), .dinb(n3371), .dout(n9965));
  jxor g09696(.dina(n9483), .dinb(n3376), .dout(n9966));
  jor  g09697(.dina(n9966), .dinb(n9774), .dout(n9967));
  jxor g09698(.dina(n9967), .dinb(n9494), .dout(n9968));
  jand g09699(.dina(n9964), .dinb(n3371), .dout(n9969));
  jor  g09700(.dina(n9969), .dinb(n9968), .dout(n9970));
  jand g09701(.dina(n9970), .dinb(n9965), .dout(n9971));
  jor  g09702(.dina(n9971), .dinb(n2875), .dout(n9972));
  jand g09703(.dina(n9965), .dinb(n2875), .dout(n9973));
  jand g09704(.dina(n9973), .dinb(n9970), .dout(n9974));
  jnot g09705(.din(n9497), .dout(n9975));
  jand g09706(.dina(asqrt[21] ), .dinb(n9975), .dout(n9976));
  jand g09707(.dina(n9976), .dinb(n9504), .dout(n9977));
  jor  g09708(.dina(n9977), .dinb(n9502), .dout(n9978));
  jand g09709(.dina(n9976), .dinb(n9505), .dout(n9979));
  jnot g09710(.din(n9979), .dout(n9980));
  jand g09711(.dina(n9980), .dinb(n9978), .dout(n9981));
  jnot g09712(.din(n9981), .dout(n9982));
  jor  g09713(.dina(n9982), .dinb(n9974), .dout(n9983));
  jand g09714(.dina(n9983), .dinb(n9972), .dout(n9984));
  jor  g09715(.dina(n9984), .dinb(n2870), .dout(n9985));
  jand g09716(.dina(n9984), .dinb(n2870), .dout(n9986));
  jor  g09717(.dina(n9986), .dinb(n9778), .dout(n9987));
  jand g09718(.dina(n9987), .dinb(n9985), .dout(n9988));
  jor  g09719(.dina(n9988), .dinb(n2425), .dout(n9989));
  jnot g09720(.din(n9513), .dout(n9990));
  jor  g09721(.dina(n9990), .dinb(n9511), .dout(n9991));
  jor  g09722(.dina(n9991), .dinb(n9774), .dout(n9992));
  jxor g09723(.dina(n9992), .dinb(n9522), .dout(n9993));
  jand g09724(.dina(n9985), .dinb(n2425), .dout(n9994));
  jand g09725(.dina(n9994), .dinb(n9987), .dout(n9995));
  jor  g09726(.dina(n9995), .dinb(n9993), .dout(n9996));
  jand g09727(.dina(n9996), .dinb(n9989), .dout(n9997));
  jor  g09728(.dina(n9997), .dinb(n2420), .dout(n9998));
  jxor g09729(.dina(n9524), .dinb(n2425), .dout(n9999));
  jor  g09730(.dina(n9999), .dinb(n9774), .dout(n10000));
  jxor g09731(.dina(n10000), .dinb(n9535), .dout(n10001));
  jand g09732(.dina(n9997), .dinb(n2420), .dout(n10002));
  jor  g09733(.dina(n10002), .dinb(n10001), .dout(n10003));
  jand g09734(.dina(n10003), .dinb(n9998), .dout(n10004));
  jor  g09735(.dina(n10004), .dinb(n2010), .dout(n10005));
  jnot g09736(.din(n9540), .dout(n10006));
  jor  g09737(.dina(n10006), .dinb(n9538), .dout(n10007));
  jor  g09738(.dina(n10007), .dinb(n9774), .dout(n10008));
  jxor g09739(.dina(n10008), .dinb(n9549), .dout(n10009));
  jand g09740(.dina(n9998), .dinb(n2010), .dout(n10010));
  jand g09741(.dina(n10010), .dinb(n10003), .dout(n10011));
  jor  g09742(.dina(n10011), .dinb(n10009), .dout(n10012));
  jand g09743(.dina(n10012), .dinb(n10005), .dout(n10013));
  jor  g09744(.dina(n10013), .dinb(n2005), .dout(n10014));
  jand g09745(.dina(n10013), .dinb(n2005), .dout(n10015));
  jnot g09746(.din(n9552), .dout(n10016));
  jand g09747(.dina(asqrt[21] ), .dinb(n10016), .dout(n10017));
  jand g09748(.dina(n10017), .dinb(n9557), .dout(n10018));
  jor  g09749(.dina(n10018), .dinb(n9556), .dout(n10019));
  jand g09750(.dina(n10017), .dinb(n9558), .dout(n10020));
  jnot g09751(.din(n10020), .dout(n10021));
  jand g09752(.dina(n10021), .dinb(n10019), .dout(n10022));
  jnot g09753(.din(n10022), .dout(n10023));
  jor  g09754(.dina(n10023), .dinb(n10015), .dout(n10024));
  jand g09755(.dina(n10024), .dinb(n10014), .dout(n10025));
  jor  g09756(.dina(n10025), .dinb(n1646), .dout(n10026));
  jand g09757(.dina(n10014), .dinb(n1646), .dout(n10027));
  jand g09758(.dina(n10027), .dinb(n10024), .dout(n10028));
  jnot g09759(.din(n9560), .dout(n10029));
  jand g09760(.dina(asqrt[21] ), .dinb(n10029), .dout(n10030));
  jand g09761(.dina(n10030), .dinb(n9567), .dout(n10031));
  jor  g09762(.dina(n10031), .dinb(n9565), .dout(n10032));
  jand g09763(.dina(n10030), .dinb(n9568), .dout(n10033));
  jnot g09764(.din(n10033), .dout(n10034));
  jand g09765(.dina(n10034), .dinb(n10032), .dout(n10035));
  jnot g09766(.din(n10035), .dout(n10036));
  jor  g09767(.dina(n10036), .dinb(n10028), .dout(n10037));
  jand g09768(.dina(n10037), .dinb(n10026), .dout(n10038));
  jor  g09769(.dina(n10038), .dinb(n1641), .dout(n10039));
  jxor g09770(.dina(n9569), .dinb(n1646), .dout(n10040));
  jor  g09771(.dina(n10040), .dinb(n9774), .dout(n10041));
  jxor g09772(.dina(n10041), .dinb(n9580), .dout(n10042));
  jand g09773(.dina(n10038), .dinb(n1641), .dout(n10043));
  jor  g09774(.dina(n10043), .dinb(n10042), .dout(n10044));
  jand g09775(.dina(n10044), .dinb(n10039), .dout(n10045));
  jor  g09776(.dina(n10045), .dinb(n1317), .dout(n10046));
  jnot g09777(.din(n9585), .dout(n10047));
  jor  g09778(.dina(n10047), .dinb(n9583), .dout(n10048));
  jor  g09779(.dina(n10048), .dinb(n9774), .dout(n10049));
  jxor g09780(.dina(n10049), .dinb(n9594), .dout(n10050));
  jand g09781(.dina(n10039), .dinb(n1317), .dout(n10051));
  jand g09782(.dina(n10051), .dinb(n10044), .dout(n10052));
  jor  g09783(.dina(n10052), .dinb(n10050), .dout(n10053));
  jand g09784(.dina(n10053), .dinb(n10046), .dout(n10054));
  jor  g09785(.dina(n10054), .dinb(n1312), .dout(n10055));
  jand g09786(.dina(n10054), .dinb(n1312), .dout(n10056));
  jnot g09787(.din(n9597), .dout(n10057));
  jand g09788(.dina(asqrt[21] ), .dinb(n10057), .dout(n10058));
  jand g09789(.dina(n10058), .dinb(n9602), .dout(n10059));
  jor  g09790(.dina(n10059), .dinb(n9601), .dout(n10060));
  jand g09791(.dina(n10058), .dinb(n9603), .dout(n10061));
  jnot g09792(.din(n10061), .dout(n10062));
  jand g09793(.dina(n10062), .dinb(n10060), .dout(n10063));
  jnot g09794(.din(n10063), .dout(n10064));
  jor  g09795(.dina(n10064), .dinb(n10056), .dout(n10065));
  jand g09796(.dina(n10065), .dinb(n10055), .dout(n10066));
  jor  g09797(.dina(n10066), .dinb(n1039), .dout(n10067));
  jand g09798(.dina(n10055), .dinb(n1039), .dout(n10068));
  jand g09799(.dina(n10068), .dinb(n10065), .dout(n10069));
  jnot g09800(.din(n9605), .dout(n10070));
  jand g09801(.dina(asqrt[21] ), .dinb(n10070), .dout(n10071));
  jand g09802(.dina(n10071), .dinb(n9612), .dout(n10072));
  jor  g09803(.dina(n10072), .dinb(n9610), .dout(n10073));
  jand g09804(.dina(n10071), .dinb(n9613), .dout(n10074));
  jnot g09805(.din(n10074), .dout(n10075));
  jand g09806(.dina(n10075), .dinb(n10073), .dout(n10076));
  jnot g09807(.din(n10076), .dout(n10077));
  jor  g09808(.dina(n10077), .dinb(n10069), .dout(n10078));
  jand g09809(.dina(n10078), .dinb(n10067), .dout(n10079));
  jor  g09810(.dina(n10079), .dinb(n1034), .dout(n10080));
  jxor g09811(.dina(n9614), .dinb(n1039), .dout(n10081));
  jor  g09812(.dina(n10081), .dinb(n9774), .dout(n10082));
  jxor g09813(.dina(n10082), .dinb(n9625), .dout(n10083));
  jand g09814(.dina(n10079), .dinb(n1034), .dout(n10084));
  jor  g09815(.dina(n10084), .dinb(n10083), .dout(n10085));
  jand g09816(.dina(n10085), .dinb(n10080), .dout(n10086));
  jor  g09817(.dina(n10086), .dinb(n796), .dout(n10087));
  jnot g09818(.din(n9630), .dout(n10088));
  jor  g09819(.dina(n10088), .dinb(n9628), .dout(n10089));
  jor  g09820(.dina(n10089), .dinb(n9774), .dout(n10090));
  jxor g09821(.dina(n10090), .dinb(n9639), .dout(n10091));
  jand g09822(.dina(n10080), .dinb(n796), .dout(n10092));
  jand g09823(.dina(n10092), .dinb(n10085), .dout(n10093));
  jor  g09824(.dina(n10093), .dinb(n10091), .dout(n10094));
  jand g09825(.dina(n10094), .dinb(n10087), .dout(n10095));
  jor  g09826(.dina(n10095), .dinb(n791), .dout(n10096));
  jand g09827(.dina(n10095), .dinb(n791), .dout(n10097));
  jnot g09828(.din(n9642), .dout(n10098));
  jand g09829(.dina(asqrt[21] ), .dinb(n10098), .dout(n10099));
  jand g09830(.dina(n10099), .dinb(n9647), .dout(n10100));
  jor  g09831(.dina(n10100), .dinb(n9646), .dout(n10101));
  jand g09832(.dina(n10099), .dinb(n9648), .dout(n10102));
  jnot g09833(.din(n10102), .dout(n10103));
  jand g09834(.dina(n10103), .dinb(n10101), .dout(n10104));
  jnot g09835(.din(n10104), .dout(n10105));
  jor  g09836(.dina(n10105), .dinb(n10097), .dout(n10106));
  jand g09837(.dina(n10106), .dinb(n10096), .dout(n10107));
  jor  g09838(.dina(n10107), .dinb(n595), .dout(n10108));
  jand g09839(.dina(n10096), .dinb(n595), .dout(n10109));
  jand g09840(.dina(n10109), .dinb(n10106), .dout(n10110));
  jnot g09841(.din(n9650), .dout(n10111));
  jand g09842(.dina(asqrt[21] ), .dinb(n10111), .dout(n10112));
  jand g09843(.dina(n10112), .dinb(n9657), .dout(n10113));
  jor  g09844(.dina(n10113), .dinb(n9655), .dout(n10114));
  jand g09845(.dina(n10112), .dinb(n9658), .dout(n10115));
  jnot g09846(.din(n10115), .dout(n10116));
  jand g09847(.dina(n10116), .dinb(n10114), .dout(n10117));
  jnot g09848(.din(n10117), .dout(n10118));
  jor  g09849(.dina(n10118), .dinb(n10110), .dout(n10119));
  jand g09850(.dina(n10119), .dinb(n10108), .dout(n10120));
  jor  g09851(.dina(n10120), .dinb(n590), .dout(n10121));
  jxor g09852(.dina(n9659), .dinb(n595), .dout(n10122));
  jor  g09853(.dina(n10122), .dinb(n9774), .dout(n10123));
  jxor g09854(.dina(n10123), .dinb(n9670), .dout(n10124));
  jand g09855(.dina(n10120), .dinb(n590), .dout(n10125));
  jor  g09856(.dina(n10125), .dinb(n10124), .dout(n10126));
  jand g09857(.dina(n10126), .dinb(n10121), .dout(n10127));
  jor  g09858(.dina(n10127), .dinb(n430), .dout(n10128));
  jnot g09859(.din(n9675), .dout(n10129));
  jor  g09860(.dina(n10129), .dinb(n9673), .dout(n10130));
  jor  g09861(.dina(n10130), .dinb(n9774), .dout(n10131));
  jxor g09862(.dina(n10131), .dinb(n9684), .dout(n10132));
  jand g09863(.dina(n10121), .dinb(n430), .dout(n10133));
  jand g09864(.dina(n10133), .dinb(n10126), .dout(n10134));
  jor  g09865(.dina(n10134), .dinb(n10132), .dout(n10135));
  jand g09866(.dina(n10135), .dinb(n10128), .dout(n10136));
  jor  g09867(.dina(n10136), .dinb(n425), .dout(n10137));
  jand g09868(.dina(n10136), .dinb(n425), .dout(n10138));
  jnot g09869(.din(n9687), .dout(n10139));
  jand g09870(.dina(asqrt[21] ), .dinb(n10139), .dout(n10140));
  jand g09871(.dina(n10140), .dinb(n9692), .dout(n10141));
  jor  g09872(.dina(n10141), .dinb(n9691), .dout(n10142));
  jand g09873(.dina(n10140), .dinb(n9693), .dout(n10143));
  jnot g09874(.din(n10143), .dout(n10144));
  jand g09875(.dina(n10144), .dinb(n10142), .dout(n10145));
  jnot g09876(.din(n10145), .dout(n10146));
  jor  g09877(.dina(n10146), .dinb(n10138), .dout(n10147));
  jand g09878(.dina(n10147), .dinb(n10137), .dout(n10148));
  jor  g09879(.dina(n10148), .dinb(n305), .dout(n10149));
  jand g09880(.dina(n10137), .dinb(n305), .dout(n10150));
  jand g09881(.dina(n10150), .dinb(n10147), .dout(n10151));
  jnot g09882(.din(n9695), .dout(n10152));
  jand g09883(.dina(asqrt[21] ), .dinb(n10152), .dout(n10153));
  jand g09884(.dina(n10153), .dinb(n9702), .dout(n10154));
  jor  g09885(.dina(n10154), .dinb(n9700), .dout(n10155));
  jand g09886(.dina(n10153), .dinb(n9703), .dout(n10156));
  jnot g09887(.din(n10156), .dout(n10157));
  jand g09888(.dina(n10157), .dinb(n10155), .dout(n10158));
  jnot g09889(.din(n10158), .dout(n10159));
  jor  g09890(.dina(n10159), .dinb(n10151), .dout(n10160));
  jand g09891(.dina(n10160), .dinb(n10149), .dout(n10161));
  jor  g09892(.dina(n10161), .dinb(n290), .dout(n10162));
  jxor g09893(.dina(n9704), .dinb(n305), .dout(n10163));
  jor  g09894(.dina(n10163), .dinb(n9774), .dout(n10164));
  jxor g09895(.dina(n10164), .dinb(n9715), .dout(n10165));
  jand g09896(.dina(n10161), .dinb(n290), .dout(n10166));
  jor  g09897(.dina(n10166), .dinb(n10165), .dout(n10167));
  jand g09898(.dina(n10167), .dinb(n10162), .dout(n10168));
  jor  g09899(.dina(n10168), .dinb(n223), .dout(n10169));
  jnot g09900(.din(n9720), .dout(n10170));
  jor  g09901(.dina(n10170), .dinb(n9718), .dout(n10171));
  jor  g09902(.dina(n10171), .dinb(n9774), .dout(n10172));
  jxor g09903(.dina(n10172), .dinb(n9729), .dout(n10173));
  jand g09904(.dina(n10162), .dinb(n223), .dout(n10174));
  jand g09905(.dina(n10174), .dinb(n10167), .dout(n10175));
  jor  g09906(.dina(n10175), .dinb(n10173), .dout(n10176));
  jand g09907(.dina(n10176), .dinb(n10169), .dout(n10177));
  jor  g09908(.dina(n10177), .dinb(n199), .dout(n10178));
  jand g09909(.dina(n10177), .dinb(n199), .dout(n10179));
  jnot g09910(.din(n9732), .dout(n10180));
  jand g09911(.dina(asqrt[21] ), .dinb(n10180), .dout(n10181));
  jand g09912(.dina(n10181), .dinb(n9737), .dout(n10182));
  jor  g09913(.dina(n10182), .dinb(n9736), .dout(n10183));
  jand g09914(.dina(n10181), .dinb(n9738), .dout(n10184));
  jnot g09915(.din(n10184), .dout(n10185));
  jand g09916(.dina(n10185), .dinb(n10183), .dout(n10186));
  jnot g09917(.din(n10186), .dout(n10187));
  jor  g09918(.dina(n10187), .dinb(n10179), .dout(n10188));
  jand g09919(.dina(n10188), .dinb(n10178), .dout(n10189));
  jnot g09920(.din(n9740), .dout(n10190));
  jand g09921(.dina(asqrt[21] ), .dinb(n10190), .dout(n10191));
  jand g09922(.dina(n10191), .dinb(n9747), .dout(n10192));
  jor  g09923(.dina(n10192), .dinb(n9745), .dout(n10193));
  jand g09924(.dina(n10191), .dinb(n9748), .dout(n10194));
  jnot g09925(.din(n10194), .dout(n10195));
  jand g09926(.dina(n10195), .dinb(n10193), .dout(n10196));
  jnot g09927(.din(n10196), .dout(n10197));
  jand g09928(.dina(asqrt[21] ), .dinb(n9762), .dout(n10198));
  jand g09929(.dina(n10198), .dinb(n9749), .dout(n10199));
  jor  g09930(.dina(n10199), .dinb(n9797), .dout(n10200));
  jor  g09931(.dina(n10200), .dinb(n10197), .dout(n10201));
  jor  g09932(.dina(n10201), .dinb(n10189), .dout(n10202));
  jand g09933(.dina(n10202), .dinb(n194), .dout(n10203));
  jand g09934(.dina(n10197), .dinb(n10189), .dout(n10204));
  jor  g09935(.dina(n10198), .dinb(n9749), .dout(n10205));
  jand g09936(.dina(n9762), .dinb(n9749), .dout(n10206));
  jor  g09937(.dina(n10206), .dinb(n194), .dout(n10207));
  jnot g09938(.din(n10207), .dout(n10208));
  jand g09939(.dina(n10208), .dinb(n10205), .dout(n10209));
  jor  g09940(.dina(n10209), .dinb(n10204), .dout(n10212));
  jor  g09941(.dina(n10212), .dinb(n10203), .dout(asqrt[20] ));
  jxor g09942(.dina(n9984), .dinb(n2870), .dout(n10214));
  jand g09943(.dina(n10214), .dinb(asqrt[20] ), .dout(n10215));
  jxor g09944(.dina(n10215), .dinb(n9778), .dout(n10216));
  jnot g09945(.din(n10216), .dout(n10217));
  jand g09946(.dina(asqrt[20] ), .dinb(a[40] ), .dout(n10218));
  jnot g09947(.din(a[38] ), .dout(n10219));
  jnot g09948(.din(a[39] ), .dout(n10220));
  jand g09949(.dina(n9780), .dinb(n10220), .dout(n10221));
  jand g09950(.dina(n10221), .dinb(n10219), .dout(n10222));
  jor  g09951(.dina(n10222), .dinb(n10218), .dout(n10223));
  jand g09952(.dina(n10223), .dinb(asqrt[21] ), .dout(n10224));
  jand g09953(.dina(asqrt[20] ), .dinb(n9780), .dout(n10225));
  jxor g09954(.dina(n10225), .dinb(n9781), .dout(n10226));
  jor  g09955(.dina(n10223), .dinb(asqrt[21] ), .dout(n10227));
  jand g09956(.dina(n10227), .dinb(n10226), .dout(n10228));
  jor  g09957(.dina(n10228), .dinb(n10224), .dout(n10229));
  jand g09958(.dina(n10229), .dinb(asqrt[22] ), .dout(n10230));
  jor  g09959(.dina(n10224), .dinb(asqrt[22] ), .dout(n10231));
  jor  g09960(.dina(n10231), .dinb(n10228), .dout(n10232));
  jand g09961(.dina(n10225), .dinb(n9781), .dout(n10233));
  jnot g09962(.din(n10203), .dout(n10234));
  jnot g09963(.din(n10204), .dout(n10235));
  jnot g09964(.din(n10209), .dout(n10236));
  jand g09965(.dina(n10236), .dinb(asqrt[21] ), .dout(n10237));
  jand g09966(.dina(n10237), .dinb(n10235), .dout(n10238));
  jand g09967(.dina(n10238), .dinb(n10234), .dout(n10239));
  jor  g09968(.dina(n10239), .dinb(n10233), .dout(n10240));
  jxor g09969(.dina(n10240), .dinb(n9318), .dout(n10241));
  jand g09970(.dina(n10241), .dinb(n10232), .dout(n10242));
  jor  g09971(.dina(n10242), .dinb(n10230), .dout(n10243));
  jand g09972(.dina(n10243), .dinb(asqrt[23] ), .dout(n10244));
  jor  g09973(.dina(n10243), .dinb(asqrt[23] ), .dout(n10245));
  jxor g09974(.dina(n9785), .dinb(n9769), .dout(n10246));
  jand g09975(.dina(n10246), .dinb(asqrt[20] ), .dout(n10247));
  jxor g09976(.dina(n10247), .dinb(n9788), .dout(n10248));
  jnot g09977(.din(n10248), .dout(n10249));
  jand g09978(.dina(n10249), .dinb(n10245), .dout(n10250));
  jor  g09979(.dina(n10250), .dinb(n10244), .dout(n10251));
  jand g09980(.dina(n10251), .dinb(asqrt[24] ), .dout(n10252));
  jnot g09981(.din(n9794), .dout(n10253));
  jand g09982(.dina(n10253), .dinb(n9792), .dout(n10254));
  jand g09983(.dina(n10254), .dinb(asqrt[20] ), .dout(n10255));
  jxor g09984(.dina(n10255), .dinb(n9802), .dout(n10256));
  jnot g09985(.din(n10256), .dout(n10257));
  jor  g09986(.dina(n10244), .dinb(asqrt[24] ), .dout(n10258));
  jor  g09987(.dina(n10258), .dinb(n10250), .dout(n10259));
  jand g09988(.dina(n10259), .dinb(n10257), .dout(n10260));
  jor  g09989(.dina(n10260), .dinb(n10252), .dout(n10261));
  jand g09990(.dina(n10261), .dinb(asqrt[25] ), .dout(n10262));
  jor  g09991(.dina(n10261), .dinb(asqrt[25] ), .dout(n10263));
  jnot g09992(.din(n9809), .dout(n10264));
  jxor g09993(.dina(n9804), .dinb(n8893), .dout(n10265));
  jand g09994(.dina(n10265), .dinb(asqrt[20] ), .dout(n10266));
  jxor g09995(.dina(n10266), .dinb(n10264), .dout(n10267));
  jand g09996(.dina(n10267), .dinb(n10263), .dout(n10268));
  jor  g09997(.dina(n10268), .dinb(n10262), .dout(n10269));
  jand g09998(.dina(n10269), .dinb(asqrt[26] ), .dout(n10270));
  jor  g09999(.dina(n10262), .dinb(asqrt[26] ), .dout(n10271));
  jor  g10000(.dina(n10271), .dinb(n10268), .dout(n10272));
  jnot g10001(.din(n9816), .dout(n10273));
  jnot g10002(.din(n9818), .dout(n10274));
  jand g10003(.dina(asqrt[20] ), .dinb(n9812), .dout(n10275));
  jand g10004(.dina(n10275), .dinb(n10274), .dout(n10276));
  jor  g10005(.dina(n10276), .dinb(n10273), .dout(n10277));
  jnot g10006(.din(n9819), .dout(n10278));
  jand g10007(.dina(n10275), .dinb(n10278), .dout(n10279));
  jnot g10008(.din(n10279), .dout(n10280));
  jand g10009(.dina(n10280), .dinb(n10277), .dout(n10281));
  jand g10010(.dina(n10281), .dinb(n10272), .dout(n10282));
  jor  g10011(.dina(n10282), .dinb(n10270), .dout(n10283));
  jand g10012(.dina(n10283), .dinb(asqrt[27] ), .dout(n10284));
  jor  g10013(.dina(n10283), .dinb(asqrt[27] ), .dout(n10285));
  jxor g10014(.dina(n9820), .dinb(n8053), .dout(n10286));
  jand g10015(.dina(n10286), .dinb(asqrt[20] ), .dout(n10287));
  jxor g10016(.dina(n10287), .dinb(n9825), .dout(n10288));
  jand g10017(.dina(n10288), .dinb(n10285), .dout(n10289));
  jor  g10018(.dina(n10289), .dinb(n10284), .dout(n10290));
  jand g10019(.dina(n10290), .dinb(asqrt[28] ), .dout(n10291));
  jnot g10020(.din(n9831), .dout(n10292));
  jand g10021(.dina(n10292), .dinb(n9829), .dout(n10293));
  jand g10022(.dina(n10293), .dinb(asqrt[20] ), .dout(n10294));
  jxor g10023(.dina(n10294), .dinb(n9840), .dout(n10295));
  jnot g10024(.din(n10295), .dout(n10296));
  jor  g10025(.dina(n10284), .dinb(asqrt[28] ), .dout(n10297));
  jor  g10026(.dina(n10297), .dinb(n10289), .dout(n10298));
  jand g10027(.dina(n10298), .dinb(n10296), .dout(n10299));
  jor  g10028(.dina(n10299), .dinb(n10291), .dout(n10300));
  jand g10029(.dina(n10300), .dinb(asqrt[29] ), .dout(n10301));
  jor  g10030(.dina(n10300), .dinb(asqrt[29] ), .dout(n10302));
  jxor g10031(.dina(n9842), .dinb(n7260), .dout(n10303));
  jand g10032(.dina(n10303), .dinb(asqrt[20] ), .dout(n10304));
  jxor g10033(.dina(n10304), .dinb(n9848), .dout(n10305));
  jand g10034(.dina(n10305), .dinb(n10302), .dout(n10306));
  jor  g10035(.dina(n10306), .dinb(n10301), .dout(n10307));
  jand g10036(.dina(n10307), .dinb(asqrt[30] ), .dout(n10308));
  jor  g10037(.dina(n10301), .dinb(asqrt[30] ), .dout(n10309));
  jor  g10038(.dina(n10309), .dinb(n10306), .dout(n10310));
  jnot g10039(.din(n9856), .dout(n10311));
  jnot g10040(.din(n9858), .dout(n10312));
  jand g10041(.dina(asqrt[20] ), .dinb(n9852), .dout(n10313));
  jand g10042(.dina(n10313), .dinb(n10312), .dout(n10314));
  jor  g10043(.dina(n10314), .dinb(n10311), .dout(n10315));
  jnot g10044(.din(n9859), .dout(n10316));
  jand g10045(.dina(n10313), .dinb(n10316), .dout(n10317));
  jnot g10046(.din(n10317), .dout(n10318));
  jand g10047(.dina(n10318), .dinb(n10315), .dout(n10319));
  jand g10048(.dina(n10319), .dinb(n10310), .dout(n10320));
  jor  g10049(.dina(n10320), .dinb(n10308), .dout(n10321));
  jand g10050(.dina(n10321), .dinb(asqrt[31] ), .dout(n10322));
  jxor g10051(.dina(n9860), .dinb(n6500), .dout(n10323));
  jand g10052(.dina(n10323), .dinb(asqrt[20] ), .dout(n10324));
  jxor g10053(.dina(n10324), .dinb(n9867), .dout(n10325));
  jnot g10054(.din(n10325), .dout(n10326));
  jor  g10055(.dina(n10321), .dinb(asqrt[31] ), .dout(n10327));
  jand g10056(.dina(n10327), .dinb(n10326), .dout(n10328));
  jor  g10057(.dina(n10328), .dinb(n10322), .dout(n10329));
  jand g10058(.dina(n10329), .dinb(asqrt[32] ), .dout(n10330));
  jnot g10059(.din(n9872), .dout(n10331));
  jand g10060(.dina(n10331), .dinb(n9870), .dout(n10332));
  jand g10061(.dina(n10332), .dinb(asqrt[20] ), .dout(n10333));
  jxor g10062(.dina(n10333), .dinb(n9880), .dout(n10334));
  jnot g10063(.din(n10334), .dout(n10335));
  jor  g10064(.dina(n10322), .dinb(asqrt[32] ), .dout(n10336));
  jor  g10065(.dina(n10336), .dinb(n10328), .dout(n10337));
  jand g10066(.dina(n10337), .dinb(n10335), .dout(n10338));
  jor  g10067(.dina(n10338), .dinb(n10330), .dout(n10339));
  jand g10068(.dina(n10339), .dinb(asqrt[33] ), .dout(n10340));
  jor  g10069(.dina(n10339), .dinb(asqrt[33] ), .dout(n10341));
  jnot g10070(.din(n9886), .dout(n10342));
  jnot g10071(.din(n9887), .dout(n10343));
  jand g10072(.dina(asqrt[20] ), .dinb(n9883), .dout(n10344));
  jand g10073(.dina(n10344), .dinb(n10343), .dout(n10345));
  jor  g10074(.dina(n10345), .dinb(n10342), .dout(n10346));
  jnot g10075(.din(n9888), .dout(n10347));
  jand g10076(.dina(n10344), .dinb(n10347), .dout(n10348));
  jnot g10077(.din(n10348), .dout(n10349));
  jand g10078(.dina(n10349), .dinb(n10346), .dout(n10350));
  jand g10079(.dina(n10350), .dinb(n10341), .dout(n10351));
  jor  g10080(.dina(n10351), .dinb(n10340), .dout(n10352));
  jand g10081(.dina(n10352), .dinb(asqrt[34] ), .dout(n10353));
  jor  g10082(.dina(n10340), .dinb(asqrt[34] ), .dout(n10354));
  jor  g10083(.dina(n10354), .dinb(n10351), .dout(n10355));
  jnot g10084(.din(n9894), .dout(n10356));
  jnot g10085(.din(n9896), .dout(n10357));
  jand g10086(.dina(asqrt[20] ), .dinb(n9890), .dout(n10358));
  jand g10087(.dina(n10358), .dinb(n10357), .dout(n10359));
  jor  g10088(.dina(n10359), .dinb(n10356), .dout(n10360));
  jnot g10089(.din(n9897), .dout(n10361));
  jand g10090(.dina(n10358), .dinb(n10361), .dout(n10362));
  jnot g10091(.din(n10362), .dout(n10363));
  jand g10092(.dina(n10363), .dinb(n10360), .dout(n10364));
  jand g10093(.dina(n10364), .dinb(n10355), .dout(n10365));
  jor  g10094(.dina(n10365), .dinb(n10353), .dout(n10366));
  jand g10095(.dina(n10366), .dinb(asqrt[35] ), .dout(n10367));
  jxor g10096(.dina(n9898), .dinb(n5116), .dout(n10368));
  jand g10097(.dina(n10368), .dinb(asqrt[20] ), .dout(n10369));
  jxor g10098(.dina(n10369), .dinb(n9908), .dout(n10370));
  jnot g10099(.din(n10370), .dout(n10371));
  jor  g10100(.dina(n10366), .dinb(asqrt[35] ), .dout(n10372));
  jand g10101(.dina(n10372), .dinb(n10371), .dout(n10373));
  jor  g10102(.dina(n10373), .dinb(n10367), .dout(n10374));
  jand g10103(.dina(n10374), .dinb(asqrt[36] ), .dout(n10375));
  jnot g10104(.din(n9913), .dout(n10376));
  jand g10105(.dina(n10376), .dinb(n9911), .dout(n10377));
  jand g10106(.dina(n10377), .dinb(asqrt[20] ), .dout(n10378));
  jxor g10107(.dina(n10378), .dinb(n9921), .dout(n10379));
  jnot g10108(.din(n10379), .dout(n10380));
  jor  g10109(.dina(n10367), .dinb(asqrt[36] ), .dout(n10381));
  jor  g10110(.dina(n10381), .dinb(n10373), .dout(n10382));
  jand g10111(.dina(n10382), .dinb(n10380), .dout(n10383));
  jor  g10112(.dina(n10383), .dinb(n10375), .dout(n10384));
  jand g10113(.dina(n10384), .dinb(asqrt[37] ), .dout(n10385));
  jor  g10114(.dina(n10384), .dinb(asqrt[37] ), .dout(n10386));
  jnot g10115(.din(n9927), .dout(n10387));
  jnot g10116(.din(n9928), .dout(n10388));
  jand g10117(.dina(asqrt[20] ), .dinb(n9924), .dout(n10389));
  jand g10118(.dina(n10389), .dinb(n10388), .dout(n10390));
  jor  g10119(.dina(n10390), .dinb(n10387), .dout(n10391));
  jnot g10120(.din(n9929), .dout(n10392));
  jand g10121(.dina(n10389), .dinb(n10392), .dout(n10393));
  jnot g10122(.din(n10393), .dout(n10394));
  jand g10123(.dina(n10394), .dinb(n10391), .dout(n10395));
  jand g10124(.dina(n10395), .dinb(n10386), .dout(n10396));
  jor  g10125(.dina(n10396), .dinb(n10385), .dout(n10397));
  jand g10126(.dina(n10397), .dinb(asqrt[38] ), .dout(n10398));
  jor  g10127(.dina(n10385), .dinb(asqrt[38] ), .dout(n10399));
  jor  g10128(.dina(n10399), .dinb(n10396), .dout(n10400));
  jnot g10129(.din(n9935), .dout(n10401));
  jnot g10130(.din(n9937), .dout(n10402));
  jand g10131(.dina(asqrt[20] ), .dinb(n9931), .dout(n10403));
  jand g10132(.dina(n10403), .dinb(n10402), .dout(n10404));
  jor  g10133(.dina(n10404), .dinb(n10401), .dout(n10405));
  jnot g10134(.din(n9938), .dout(n10406));
  jand g10135(.dina(n10403), .dinb(n10406), .dout(n10407));
  jnot g10136(.din(n10407), .dout(n10408));
  jand g10137(.dina(n10408), .dinb(n10405), .dout(n10409));
  jand g10138(.dina(n10409), .dinb(n10400), .dout(n10410));
  jor  g10139(.dina(n10410), .dinb(n10398), .dout(n10411));
  jand g10140(.dina(n10411), .dinb(asqrt[39] ), .dout(n10412));
  jxor g10141(.dina(n9939), .dinb(n3907), .dout(n10413));
  jand g10142(.dina(n10413), .dinb(asqrt[20] ), .dout(n10414));
  jxor g10143(.dina(n10414), .dinb(n9949), .dout(n10415));
  jnot g10144(.din(n10415), .dout(n10416));
  jor  g10145(.dina(n10411), .dinb(asqrt[39] ), .dout(n10417));
  jand g10146(.dina(n10417), .dinb(n10416), .dout(n10418));
  jor  g10147(.dina(n10418), .dinb(n10412), .dout(n10419));
  jand g10148(.dina(n10419), .dinb(asqrt[40] ), .dout(n10420));
  jnot g10149(.din(n9954), .dout(n10421));
  jand g10150(.dina(n10421), .dinb(n9952), .dout(n10422));
  jand g10151(.dina(n10422), .dinb(asqrt[20] ), .dout(n10423));
  jxor g10152(.dina(n10423), .dinb(n9962), .dout(n10424));
  jnot g10153(.din(n10424), .dout(n10425));
  jor  g10154(.dina(n10412), .dinb(asqrt[40] ), .dout(n10426));
  jor  g10155(.dina(n10426), .dinb(n10418), .dout(n10427));
  jand g10156(.dina(n10427), .dinb(n10425), .dout(n10428));
  jor  g10157(.dina(n10428), .dinb(n10420), .dout(n10429));
  jand g10158(.dina(n10429), .dinb(asqrt[41] ), .dout(n10430));
  jor  g10159(.dina(n10429), .dinb(asqrt[41] ), .dout(n10431));
  jnot g10160(.din(n9968), .dout(n10432));
  jnot g10161(.din(n9969), .dout(n10433));
  jand g10162(.dina(asqrt[20] ), .dinb(n9965), .dout(n10434));
  jand g10163(.dina(n10434), .dinb(n10433), .dout(n10435));
  jor  g10164(.dina(n10435), .dinb(n10432), .dout(n10436));
  jnot g10165(.din(n9970), .dout(n10437));
  jand g10166(.dina(n10434), .dinb(n10437), .dout(n10438));
  jnot g10167(.din(n10438), .dout(n10439));
  jand g10168(.dina(n10439), .dinb(n10436), .dout(n10440));
  jand g10169(.dina(n10440), .dinb(n10431), .dout(n10441));
  jor  g10170(.dina(n10441), .dinb(n10430), .dout(n10442));
  jand g10171(.dina(n10442), .dinb(asqrt[42] ), .dout(n10443));
  jnot g10172(.din(n9974), .dout(n10444));
  jand g10173(.dina(n10444), .dinb(n9972), .dout(n10445));
  jand g10174(.dina(n10445), .dinb(asqrt[20] ), .dout(n10446));
  jxor g10175(.dina(n10446), .dinb(n9982), .dout(n10447));
  jnot g10176(.din(n10447), .dout(n10448));
  jor  g10177(.dina(n10430), .dinb(asqrt[42] ), .dout(n10449));
  jor  g10178(.dina(n10449), .dinb(n10441), .dout(n10450));
  jand g10179(.dina(n10450), .dinb(n10448), .dout(n10451));
  jor  g10180(.dina(n10451), .dinb(n10443), .dout(n10452));
  jand g10181(.dina(n10452), .dinb(asqrt[43] ), .dout(n10453));
  jor  g10182(.dina(n10452), .dinb(asqrt[43] ), .dout(n10454));
  jand g10183(.dina(n10454), .dinb(n10217), .dout(n10455));
  jor  g10184(.dina(n10455), .dinb(n10453), .dout(n10456));
  jand g10185(.dina(n10456), .dinb(asqrt[44] ), .dout(n10457));
  jor  g10186(.dina(n10453), .dinb(asqrt[44] ), .dout(n10458));
  jor  g10187(.dina(n10458), .dinb(n10455), .dout(n10459));
  jnot g10188(.din(n9993), .dout(n10460));
  jnot g10189(.din(n9995), .dout(n10461));
  jand g10190(.dina(asqrt[20] ), .dinb(n9989), .dout(n10462));
  jand g10191(.dina(n10462), .dinb(n10461), .dout(n10463));
  jor  g10192(.dina(n10463), .dinb(n10460), .dout(n10464));
  jnot g10193(.din(n9996), .dout(n10465));
  jand g10194(.dina(n10462), .dinb(n10465), .dout(n10466));
  jnot g10195(.din(n10466), .dout(n10467));
  jand g10196(.dina(n10467), .dinb(n10464), .dout(n10468));
  jand g10197(.dina(n10468), .dinb(n10459), .dout(n10469));
  jor  g10198(.dina(n10469), .dinb(n10457), .dout(n10470));
  jand g10199(.dina(n10470), .dinb(asqrt[45] ), .dout(n10471));
  jor  g10200(.dina(n10470), .dinb(asqrt[45] ), .dout(n10472));
  jnot g10201(.din(n10001), .dout(n10473));
  jnot g10202(.din(n10002), .dout(n10474));
  jand g10203(.dina(asqrt[20] ), .dinb(n9998), .dout(n10475));
  jand g10204(.dina(n10475), .dinb(n10474), .dout(n10476));
  jor  g10205(.dina(n10476), .dinb(n10473), .dout(n10477));
  jnot g10206(.din(n10003), .dout(n10478));
  jand g10207(.dina(n10475), .dinb(n10478), .dout(n10479));
  jnot g10208(.din(n10479), .dout(n10480));
  jand g10209(.dina(n10480), .dinb(n10477), .dout(n10481));
  jand g10210(.dina(n10481), .dinb(n10472), .dout(n10482));
  jor  g10211(.dina(n10482), .dinb(n10471), .dout(n10483));
  jand g10212(.dina(n10483), .dinb(asqrt[46] ), .dout(n10484));
  jor  g10213(.dina(n10471), .dinb(asqrt[46] ), .dout(n10485));
  jor  g10214(.dina(n10485), .dinb(n10482), .dout(n10486));
  jnot g10215(.din(n10009), .dout(n10487));
  jnot g10216(.din(n10011), .dout(n10488));
  jand g10217(.dina(asqrt[20] ), .dinb(n10005), .dout(n10489));
  jand g10218(.dina(n10489), .dinb(n10488), .dout(n10490));
  jor  g10219(.dina(n10490), .dinb(n10487), .dout(n10491));
  jnot g10220(.din(n10012), .dout(n10492));
  jand g10221(.dina(n10489), .dinb(n10492), .dout(n10493));
  jnot g10222(.din(n10493), .dout(n10494));
  jand g10223(.dina(n10494), .dinb(n10491), .dout(n10495));
  jand g10224(.dina(n10495), .dinb(n10486), .dout(n10496));
  jor  g10225(.dina(n10496), .dinb(n10484), .dout(n10497));
  jand g10226(.dina(n10497), .dinb(asqrt[47] ), .dout(n10498));
  jxor g10227(.dina(n10013), .dinb(n2005), .dout(n10499));
  jand g10228(.dina(n10499), .dinb(asqrt[20] ), .dout(n10500));
  jxor g10229(.dina(n10500), .dinb(n10023), .dout(n10501));
  jnot g10230(.din(n10501), .dout(n10502));
  jor  g10231(.dina(n10497), .dinb(asqrt[47] ), .dout(n10503));
  jand g10232(.dina(n10503), .dinb(n10502), .dout(n10504));
  jor  g10233(.dina(n10504), .dinb(n10498), .dout(n10505));
  jand g10234(.dina(n10505), .dinb(asqrt[48] ), .dout(n10506));
  jnot g10235(.din(n10028), .dout(n10507));
  jand g10236(.dina(n10507), .dinb(n10026), .dout(n10508));
  jand g10237(.dina(n10508), .dinb(asqrt[20] ), .dout(n10509));
  jxor g10238(.dina(n10509), .dinb(n10036), .dout(n10510));
  jnot g10239(.din(n10510), .dout(n10511));
  jor  g10240(.dina(n10498), .dinb(asqrt[48] ), .dout(n10512));
  jor  g10241(.dina(n10512), .dinb(n10504), .dout(n10513));
  jand g10242(.dina(n10513), .dinb(n10511), .dout(n10514));
  jor  g10243(.dina(n10514), .dinb(n10506), .dout(n10515));
  jand g10244(.dina(n10515), .dinb(asqrt[49] ), .dout(n10516));
  jor  g10245(.dina(n10515), .dinb(asqrt[49] ), .dout(n10517));
  jnot g10246(.din(n10042), .dout(n10518));
  jnot g10247(.din(n10043), .dout(n10519));
  jand g10248(.dina(asqrt[20] ), .dinb(n10039), .dout(n10520));
  jand g10249(.dina(n10520), .dinb(n10519), .dout(n10521));
  jor  g10250(.dina(n10521), .dinb(n10518), .dout(n10522));
  jnot g10251(.din(n10044), .dout(n10523));
  jand g10252(.dina(n10520), .dinb(n10523), .dout(n10524));
  jnot g10253(.din(n10524), .dout(n10525));
  jand g10254(.dina(n10525), .dinb(n10522), .dout(n10526));
  jand g10255(.dina(n10526), .dinb(n10517), .dout(n10527));
  jor  g10256(.dina(n10527), .dinb(n10516), .dout(n10528));
  jand g10257(.dina(n10528), .dinb(asqrt[50] ), .dout(n10529));
  jor  g10258(.dina(n10516), .dinb(asqrt[50] ), .dout(n10530));
  jor  g10259(.dina(n10530), .dinb(n10527), .dout(n10531));
  jnot g10260(.din(n10050), .dout(n10532));
  jnot g10261(.din(n10052), .dout(n10533));
  jand g10262(.dina(asqrt[20] ), .dinb(n10046), .dout(n10534));
  jand g10263(.dina(n10534), .dinb(n10533), .dout(n10535));
  jor  g10264(.dina(n10535), .dinb(n10532), .dout(n10536));
  jnot g10265(.din(n10053), .dout(n10537));
  jand g10266(.dina(n10534), .dinb(n10537), .dout(n10538));
  jnot g10267(.din(n10538), .dout(n10539));
  jand g10268(.dina(n10539), .dinb(n10536), .dout(n10540));
  jand g10269(.dina(n10540), .dinb(n10531), .dout(n10541));
  jor  g10270(.dina(n10541), .dinb(n10529), .dout(n10542));
  jand g10271(.dina(n10542), .dinb(asqrt[51] ), .dout(n10543));
  jxor g10272(.dina(n10054), .dinb(n1312), .dout(n10544));
  jand g10273(.dina(n10544), .dinb(asqrt[20] ), .dout(n10545));
  jxor g10274(.dina(n10545), .dinb(n10064), .dout(n10546));
  jnot g10275(.din(n10546), .dout(n10547));
  jor  g10276(.dina(n10542), .dinb(asqrt[51] ), .dout(n10548));
  jand g10277(.dina(n10548), .dinb(n10547), .dout(n10549));
  jor  g10278(.dina(n10549), .dinb(n10543), .dout(n10550));
  jand g10279(.dina(n10550), .dinb(asqrt[52] ), .dout(n10551));
  jnot g10280(.din(n10069), .dout(n10552));
  jand g10281(.dina(n10552), .dinb(n10067), .dout(n10553));
  jand g10282(.dina(n10553), .dinb(asqrt[20] ), .dout(n10554));
  jxor g10283(.dina(n10554), .dinb(n10077), .dout(n10555));
  jnot g10284(.din(n10555), .dout(n10556));
  jor  g10285(.dina(n10543), .dinb(asqrt[52] ), .dout(n10557));
  jor  g10286(.dina(n10557), .dinb(n10549), .dout(n10558));
  jand g10287(.dina(n10558), .dinb(n10556), .dout(n10559));
  jor  g10288(.dina(n10559), .dinb(n10551), .dout(n10560));
  jand g10289(.dina(n10560), .dinb(asqrt[53] ), .dout(n10561));
  jor  g10290(.dina(n10560), .dinb(asqrt[53] ), .dout(n10562));
  jnot g10291(.din(n10083), .dout(n10563));
  jnot g10292(.din(n10084), .dout(n10564));
  jand g10293(.dina(asqrt[20] ), .dinb(n10080), .dout(n10565));
  jand g10294(.dina(n10565), .dinb(n10564), .dout(n10566));
  jor  g10295(.dina(n10566), .dinb(n10563), .dout(n10567));
  jnot g10296(.din(n10085), .dout(n10568));
  jand g10297(.dina(n10565), .dinb(n10568), .dout(n10569));
  jnot g10298(.din(n10569), .dout(n10570));
  jand g10299(.dina(n10570), .dinb(n10567), .dout(n10571));
  jand g10300(.dina(n10571), .dinb(n10562), .dout(n10572));
  jor  g10301(.dina(n10572), .dinb(n10561), .dout(n10573));
  jand g10302(.dina(n10573), .dinb(asqrt[54] ), .dout(n10574));
  jor  g10303(.dina(n10561), .dinb(asqrt[54] ), .dout(n10575));
  jor  g10304(.dina(n10575), .dinb(n10572), .dout(n10576));
  jnot g10305(.din(n10091), .dout(n10577));
  jnot g10306(.din(n10093), .dout(n10578));
  jand g10307(.dina(asqrt[20] ), .dinb(n10087), .dout(n10579));
  jand g10308(.dina(n10579), .dinb(n10578), .dout(n10580));
  jor  g10309(.dina(n10580), .dinb(n10577), .dout(n10581));
  jnot g10310(.din(n10094), .dout(n10582));
  jand g10311(.dina(n10579), .dinb(n10582), .dout(n10583));
  jnot g10312(.din(n10583), .dout(n10584));
  jand g10313(.dina(n10584), .dinb(n10581), .dout(n10585));
  jand g10314(.dina(n10585), .dinb(n10576), .dout(n10586));
  jor  g10315(.dina(n10586), .dinb(n10574), .dout(n10587));
  jand g10316(.dina(n10587), .dinb(asqrt[55] ), .dout(n10588));
  jxor g10317(.dina(n10095), .dinb(n791), .dout(n10589));
  jand g10318(.dina(n10589), .dinb(asqrt[20] ), .dout(n10590));
  jxor g10319(.dina(n10590), .dinb(n10105), .dout(n10591));
  jnot g10320(.din(n10591), .dout(n10592));
  jor  g10321(.dina(n10587), .dinb(asqrt[55] ), .dout(n10593));
  jand g10322(.dina(n10593), .dinb(n10592), .dout(n10594));
  jor  g10323(.dina(n10594), .dinb(n10588), .dout(n10595));
  jand g10324(.dina(n10595), .dinb(asqrt[56] ), .dout(n10596));
  jnot g10325(.din(n10110), .dout(n10597));
  jand g10326(.dina(n10597), .dinb(n10108), .dout(n10598));
  jand g10327(.dina(n10598), .dinb(asqrt[20] ), .dout(n10599));
  jxor g10328(.dina(n10599), .dinb(n10118), .dout(n10600));
  jnot g10329(.din(n10600), .dout(n10601));
  jor  g10330(.dina(n10588), .dinb(asqrt[56] ), .dout(n10602));
  jor  g10331(.dina(n10602), .dinb(n10594), .dout(n10603));
  jand g10332(.dina(n10603), .dinb(n10601), .dout(n10604));
  jor  g10333(.dina(n10604), .dinb(n10596), .dout(n10605));
  jand g10334(.dina(n10605), .dinb(asqrt[57] ), .dout(n10606));
  jor  g10335(.dina(n10605), .dinb(asqrt[57] ), .dout(n10607));
  jnot g10336(.din(n10124), .dout(n10608));
  jnot g10337(.din(n10125), .dout(n10609));
  jand g10338(.dina(asqrt[20] ), .dinb(n10121), .dout(n10610));
  jand g10339(.dina(n10610), .dinb(n10609), .dout(n10611));
  jor  g10340(.dina(n10611), .dinb(n10608), .dout(n10612));
  jnot g10341(.din(n10126), .dout(n10613));
  jand g10342(.dina(n10610), .dinb(n10613), .dout(n10614));
  jnot g10343(.din(n10614), .dout(n10615));
  jand g10344(.dina(n10615), .dinb(n10612), .dout(n10616));
  jand g10345(.dina(n10616), .dinb(n10607), .dout(n10617));
  jor  g10346(.dina(n10617), .dinb(n10606), .dout(n10618));
  jand g10347(.dina(n10618), .dinb(asqrt[58] ), .dout(n10619));
  jor  g10348(.dina(n10606), .dinb(asqrt[58] ), .dout(n10620));
  jor  g10349(.dina(n10620), .dinb(n10617), .dout(n10621));
  jnot g10350(.din(n10132), .dout(n10622));
  jnot g10351(.din(n10134), .dout(n10623));
  jand g10352(.dina(asqrt[20] ), .dinb(n10128), .dout(n10624));
  jand g10353(.dina(n10624), .dinb(n10623), .dout(n10625));
  jor  g10354(.dina(n10625), .dinb(n10622), .dout(n10626));
  jnot g10355(.din(n10135), .dout(n10627));
  jand g10356(.dina(n10624), .dinb(n10627), .dout(n10628));
  jnot g10357(.din(n10628), .dout(n10629));
  jand g10358(.dina(n10629), .dinb(n10626), .dout(n10630));
  jand g10359(.dina(n10630), .dinb(n10621), .dout(n10631));
  jor  g10360(.dina(n10631), .dinb(n10619), .dout(n10632));
  jand g10361(.dina(n10632), .dinb(asqrt[59] ), .dout(n10633));
  jxor g10362(.dina(n10136), .dinb(n425), .dout(n10634));
  jand g10363(.dina(n10634), .dinb(asqrt[20] ), .dout(n10635));
  jxor g10364(.dina(n10635), .dinb(n10146), .dout(n10636));
  jnot g10365(.din(n10636), .dout(n10637));
  jor  g10366(.dina(n10632), .dinb(asqrt[59] ), .dout(n10638));
  jand g10367(.dina(n10638), .dinb(n10637), .dout(n10639));
  jor  g10368(.dina(n10639), .dinb(n10633), .dout(n10640));
  jand g10369(.dina(n10640), .dinb(asqrt[60] ), .dout(n10641));
  jnot g10370(.din(n10151), .dout(n10642));
  jand g10371(.dina(n10642), .dinb(n10149), .dout(n10643));
  jand g10372(.dina(n10643), .dinb(asqrt[20] ), .dout(n10644));
  jxor g10373(.dina(n10644), .dinb(n10159), .dout(n10645));
  jnot g10374(.din(n10645), .dout(n10646));
  jor  g10375(.dina(n10633), .dinb(asqrt[60] ), .dout(n10647));
  jor  g10376(.dina(n10647), .dinb(n10639), .dout(n10648));
  jand g10377(.dina(n10648), .dinb(n10646), .dout(n10649));
  jor  g10378(.dina(n10649), .dinb(n10641), .dout(n10650));
  jand g10379(.dina(n10650), .dinb(asqrt[61] ), .dout(n10651));
  jor  g10380(.dina(n10650), .dinb(asqrt[61] ), .dout(n10652));
  jnot g10381(.din(n10165), .dout(n10653));
  jnot g10382(.din(n10166), .dout(n10654));
  jand g10383(.dina(asqrt[20] ), .dinb(n10162), .dout(n10655));
  jand g10384(.dina(n10655), .dinb(n10654), .dout(n10656));
  jor  g10385(.dina(n10656), .dinb(n10653), .dout(n10657));
  jnot g10386(.din(n10167), .dout(n10658));
  jand g10387(.dina(n10655), .dinb(n10658), .dout(n10659));
  jnot g10388(.din(n10659), .dout(n10660));
  jand g10389(.dina(n10660), .dinb(n10657), .dout(n10661));
  jand g10390(.dina(n10661), .dinb(n10652), .dout(n10662));
  jor  g10391(.dina(n10662), .dinb(n10651), .dout(n10663));
  jand g10392(.dina(n10663), .dinb(asqrt[62] ), .dout(n10664));
  jor  g10393(.dina(n10651), .dinb(asqrt[62] ), .dout(n10665));
  jor  g10394(.dina(n10665), .dinb(n10662), .dout(n10666));
  jnot g10395(.din(n10173), .dout(n10667));
  jnot g10396(.din(n10175), .dout(n10668));
  jand g10397(.dina(asqrt[20] ), .dinb(n10169), .dout(n10669));
  jand g10398(.dina(n10669), .dinb(n10668), .dout(n10670));
  jor  g10399(.dina(n10670), .dinb(n10667), .dout(n10671));
  jnot g10400(.din(n10176), .dout(n10672));
  jand g10401(.dina(n10669), .dinb(n10672), .dout(n10673));
  jnot g10402(.din(n10673), .dout(n10674));
  jand g10403(.dina(n10674), .dinb(n10671), .dout(n10675));
  jand g10404(.dina(n10675), .dinb(n10666), .dout(n10676));
  jor  g10405(.dina(n10676), .dinb(n10664), .dout(n10677));
  jxor g10406(.dina(n10177), .dinb(n199), .dout(n10678));
  jand g10407(.dina(n10678), .dinb(asqrt[20] ), .dout(n10679));
  jxor g10408(.dina(n10679), .dinb(n10187), .dout(n10680));
  jnot g10409(.din(n10189), .dout(n10681));
  jand g10410(.dina(asqrt[20] ), .dinb(n10196), .dout(n10682));
  jand g10411(.dina(n10682), .dinb(n10681), .dout(n10683));
  jor  g10412(.dina(n10683), .dinb(n10204), .dout(n10684));
  jor  g10413(.dina(n10684), .dinb(n10680), .dout(n10685));
  jnot g10414(.din(n10685), .dout(n10686));
  jand g10415(.dina(n10686), .dinb(n10677), .dout(n10687));
  jor  g10416(.dina(n10687), .dinb(asqrt[63] ), .dout(n10688));
  jnot g10417(.din(n10680), .dout(n10689));
  jor  g10418(.dina(n10689), .dinb(n10677), .dout(n10690));
  jor  g10419(.dina(n10682), .dinb(n10681), .dout(n10691));
  jand g10420(.dina(n10196), .dinb(n10681), .dout(n10692));
  jor  g10421(.dina(n10692), .dinb(n194), .dout(n10693));
  jnot g10422(.din(n10693), .dout(n10694));
  jand g10423(.dina(n10694), .dinb(n10691), .dout(n10695));
  jnot g10424(.din(asqrt[20] ), .dout(n10696));
  jnot g10425(.din(n10695), .dout(n10699));
  jand g10426(.dina(n10699), .dinb(n10690), .dout(n10700));
  jand g10427(.dina(n10700), .dinb(n10688), .dout(n10701));
  jxor g10428(.dina(n10452), .dinb(n2425), .dout(n10702));
  jor  g10429(.dina(n10702), .dinb(n10701), .dout(n10703));
  jxor g10430(.dina(n10703), .dinb(n10217), .dout(n10704));
  jor  g10431(.dina(n10701), .dinb(n10219), .dout(n10705));
  jnot g10432(.din(a[36] ), .dout(n10706));
  jnot g10433(.din(a[37] ), .dout(n10707));
  jand g10434(.dina(n10219), .dinb(n10707), .dout(n10708));
  jand g10435(.dina(n10708), .dinb(n10706), .dout(n10709));
  jnot g10436(.din(n10709), .dout(n10710));
  jand g10437(.dina(n10710), .dinb(n10705), .dout(n10711));
  jor  g10438(.dina(n10711), .dinb(n10696), .dout(n10712));
  jor  g10439(.dina(n10701), .dinb(a[38] ), .dout(n10713));
  jxor g10440(.dina(n10713), .dinb(n10220), .dout(n10714));
  jand g10441(.dina(n10711), .dinb(n10696), .dout(n10715));
  jor  g10442(.dina(n10715), .dinb(n10714), .dout(n10716));
  jand g10443(.dina(n10716), .dinb(n10712), .dout(n10717));
  jor  g10444(.dina(n10717), .dinb(n9774), .dout(n10718));
  jand g10445(.dina(n10712), .dinb(n9774), .dout(n10719));
  jand g10446(.dina(n10719), .dinb(n10716), .dout(n10720));
  jor  g10447(.dina(n10713), .dinb(a[39] ), .dout(n10721));
  jnot g10448(.din(n10688), .dout(n10722));
  jnot g10449(.din(n10690), .dout(n10723));
  jor  g10450(.dina(n10695), .dinb(n10696), .dout(n10724));
  jor  g10451(.dina(n10724), .dinb(n10723), .dout(n10725));
  jor  g10452(.dina(n10725), .dinb(n10722), .dout(n10726));
  jand g10453(.dina(n10726), .dinb(n10721), .dout(n10727));
  jxor g10454(.dina(n10727), .dinb(n9780), .dout(n10728));
  jor  g10455(.dina(n10728), .dinb(n10720), .dout(n10729));
  jand g10456(.dina(n10729), .dinb(n10718), .dout(n10730));
  jor  g10457(.dina(n10730), .dinb(n9769), .dout(n10731));
  jand g10458(.dina(n10730), .dinb(n9769), .dout(n10732));
  jxor g10459(.dina(n10223), .dinb(n9774), .dout(n10733));
  jor  g10460(.dina(n10733), .dinb(n10701), .dout(n10734));
  jxor g10461(.dina(n10734), .dinb(n10226), .dout(n10735));
  jor  g10462(.dina(n10735), .dinb(n10732), .dout(n10736));
  jand g10463(.dina(n10736), .dinb(n10731), .dout(n10737));
  jor  g10464(.dina(n10737), .dinb(n8898), .dout(n10738));
  jnot g10465(.din(n10232), .dout(n10739));
  jor  g10466(.dina(n10739), .dinb(n10230), .dout(n10740));
  jor  g10467(.dina(n10740), .dinb(n10701), .dout(n10741));
  jxor g10468(.dina(n10741), .dinb(n10241), .dout(n10742));
  jand g10469(.dina(n10731), .dinb(n8898), .dout(n10743));
  jand g10470(.dina(n10743), .dinb(n10736), .dout(n10744));
  jor  g10471(.dina(n10744), .dinb(n10742), .dout(n10745));
  jand g10472(.dina(n10745), .dinb(n10738), .dout(n10746));
  jor  g10473(.dina(n10746), .dinb(n8893), .dout(n10747));
  jand g10474(.dina(n10746), .dinb(n8893), .dout(n10748));
  jxor g10475(.dina(n10243), .dinb(n8898), .dout(n10749));
  jor  g10476(.dina(n10749), .dinb(n10701), .dout(n10750));
  jxor g10477(.dina(n10750), .dinb(n10248), .dout(n10751));
  jnot g10478(.din(n10751), .dout(n10752));
  jor  g10479(.dina(n10752), .dinb(n10748), .dout(n10753));
  jand g10480(.dina(n10753), .dinb(n10747), .dout(n10754));
  jor  g10481(.dina(n10754), .dinb(n8058), .dout(n10755));
  jand g10482(.dina(n10747), .dinb(n8058), .dout(n10756));
  jand g10483(.dina(n10756), .dinb(n10753), .dout(n10757));
  jnot g10484(.din(n10252), .dout(n10758));
  jnot g10485(.din(n10701), .dout(asqrt[19] ));
  jand g10486(.dina(asqrt[19] ), .dinb(n10758), .dout(n10760));
  jand g10487(.dina(n10760), .dinb(n10259), .dout(n10761));
  jor  g10488(.dina(n10761), .dinb(n10257), .dout(n10762));
  jand g10489(.dina(n10760), .dinb(n10260), .dout(n10763));
  jnot g10490(.din(n10763), .dout(n10764));
  jand g10491(.dina(n10764), .dinb(n10762), .dout(n10765));
  jnot g10492(.din(n10765), .dout(n10766));
  jor  g10493(.dina(n10766), .dinb(n10757), .dout(n10767));
  jand g10494(.dina(n10767), .dinb(n10755), .dout(n10768));
  jor  g10495(.dina(n10768), .dinb(n8053), .dout(n10769));
  jand g10496(.dina(n10768), .dinb(n8053), .dout(n10770));
  jnot g10497(.din(n10267), .dout(n10771));
  jxor g10498(.dina(n10261), .dinb(n8058), .dout(n10772));
  jor  g10499(.dina(n10772), .dinb(n10701), .dout(n10773));
  jxor g10500(.dina(n10773), .dinb(n10771), .dout(n10774));
  jnot g10501(.din(n10774), .dout(n10775));
  jor  g10502(.dina(n10775), .dinb(n10770), .dout(n10776));
  jand g10503(.dina(n10776), .dinb(n10769), .dout(n10777));
  jor  g10504(.dina(n10777), .dinb(n7265), .dout(n10778));
  jnot g10505(.din(n10272), .dout(n10779));
  jor  g10506(.dina(n10779), .dinb(n10270), .dout(n10780));
  jor  g10507(.dina(n10780), .dinb(n10701), .dout(n10781));
  jxor g10508(.dina(n10781), .dinb(n10281), .dout(n10782));
  jand g10509(.dina(n10769), .dinb(n7265), .dout(n10783));
  jand g10510(.dina(n10783), .dinb(n10776), .dout(n10784));
  jor  g10511(.dina(n10784), .dinb(n10782), .dout(n10785));
  jand g10512(.dina(n10785), .dinb(n10778), .dout(n10786));
  jor  g10513(.dina(n10786), .dinb(n7260), .dout(n10787));
  jand g10514(.dina(n10786), .dinb(n7260), .dout(n10788));
  jnot g10515(.din(n10288), .dout(n10789));
  jxor g10516(.dina(n10283), .dinb(n7265), .dout(n10790));
  jor  g10517(.dina(n10790), .dinb(n10701), .dout(n10791));
  jxor g10518(.dina(n10791), .dinb(n10789), .dout(n10792));
  jnot g10519(.din(n10792), .dout(n10793));
  jor  g10520(.dina(n10793), .dinb(n10788), .dout(n10794));
  jand g10521(.dina(n10794), .dinb(n10787), .dout(n10795));
  jor  g10522(.dina(n10795), .dinb(n6505), .dout(n10796));
  jand g10523(.dina(n10787), .dinb(n6505), .dout(n10797));
  jand g10524(.dina(n10797), .dinb(n10794), .dout(n10798));
  jnot g10525(.din(n10291), .dout(n10799));
  jand g10526(.dina(asqrt[19] ), .dinb(n10799), .dout(n10800));
  jand g10527(.dina(n10800), .dinb(n10298), .dout(n10801));
  jor  g10528(.dina(n10801), .dinb(n10296), .dout(n10802));
  jand g10529(.dina(n10800), .dinb(n10299), .dout(n10803));
  jnot g10530(.din(n10803), .dout(n10804));
  jand g10531(.dina(n10804), .dinb(n10802), .dout(n10805));
  jnot g10532(.din(n10805), .dout(n10806));
  jor  g10533(.dina(n10806), .dinb(n10798), .dout(n10807));
  jand g10534(.dina(n10807), .dinb(n10796), .dout(n10808));
  jor  g10535(.dina(n10808), .dinb(n6500), .dout(n10809));
  jxor g10536(.dina(n10300), .dinb(n6505), .dout(n10810));
  jor  g10537(.dina(n10810), .dinb(n10701), .dout(n10811));
  jxor g10538(.dina(n10811), .dinb(n10305), .dout(n10812));
  jand g10539(.dina(n10808), .dinb(n6500), .dout(n10813));
  jor  g10540(.dina(n10813), .dinb(n10812), .dout(n10814));
  jand g10541(.dina(n10814), .dinb(n10809), .dout(n10815));
  jor  g10542(.dina(n10815), .dinb(n5793), .dout(n10816));
  jnot g10543(.din(n10310), .dout(n10817));
  jor  g10544(.dina(n10817), .dinb(n10308), .dout(n10818));
  jor  g10545(.dina(n10818), .dinb(n10701), .dout(n10819));
  jxor g10546(.dina(n10819), .dinb(n10319), .dout(n10820));
  jand g10547(.dina(n10809), .dinb(n5793), .dout(n10821));
  jand g10548(.dina(n10821), .dinb(n10814), .dout(n10822));
  jor  g10549(.dina(n10822), .dinb(n10820), .dout(n10823));
  jand g10550(.dina(n10823), .dinb(n10816), .dout(n10824));
  jor  g10551(.dina(n10824), .dinb(n5788), .dout(n10825));
  jand g10552(.dina(n10824), .dinb(n5788), .dout(n10826));
  jnot g10553(.din(n10322), .dout(n10827));
  jand g10554(.dina(asqrt[19] ), .dinb(n10827), .dout(n10828));
  jand g10555(.dina(n10828), .dinb(n10327), .dout(n10829));
  jor  g10556(.dina(n10829), .dinb(n10326), .dout(n10830));
  jand g10557(.dina(n10828), .dinb(n10328), .dout(n10831));
  jnot g10558(.din(n10831), .dout(n10832));
  jand g10559(.dina(n10832), .dinb(n10830), .dout(n10833));
  jnot g10560(.din(n10833), .dout(n10834));
  jor  g10561(.dina(n10834), .dinb(n10826), .dout(n10835));
  jand g10562(.dina(n10835), .dinb(n10825), .dout(n10836));
  jor  g10563(.dina(n10836), .dinb(n5121), .dout(n10837));
  jand g10564(.dina(n10825), .dinb(n5121), .dout(n10838));
  jand g10565(.dina(n10838), .dinb(n10835), .dout(n10839));
  jnot g10566(.din(n10330), .dout(n10840));
  jand g10567(.dina(asqrt[19] ), .dinb(n10840), .dout(n10841));
  jand g10568(.dina(n10841), .dinb(n10337), .dout(n10842));
  jor  g10569(.dina(n10842), .dinb(n10335), .dout(n10843));
  jand g10570(.dina(n10841), .dinb(n10338), .dout(n10844));
  jnot g10571(.din(n10844), .dout(n10845));
  jand g10572(.dina(n10845), .dinb(n10843), .dout(n10846));
  jnot g10573(.din(n10846), .dout(n10847));
  jor  g10574(.dina(n10847), .dinb(n10839), .dout(n10848));
  jand g10575(.dina(n10848), .dinb(n10837), .dout(n10849));
  jor  g10576(.dina(n10849), .dinb(n5116), .dout(n10850));
  jxor g10577(.dina(n10339), .dinb(n5121), .dout(n10851));
  jor  g10578(.dina(n10851), .dinb(n10701), .dout(n10852));
  jxor g10579(.dina(n10852), .dinb(n10350), .dout(n10853));
  jand g10580(.dina(n10849), .dinb(n5116), .dout(n10854));
  jor  g10581(.dina(n10854), .dinb(n10853), .dout(n10855));
  jand g10582(.dina(n10855), .dinb(n10850), .dout(n10856));
  jor  g10583(.dina(n10856), .dinb(n4499), .dout(n10857));
  jnot g10584(.din(n10355), .dout(n10858));
  jor  g10585(.dina(n10858), .dinb(n10353), .dout(n10859));
  jor  g10586(.dina(n10859), .dinb(n10701), .dout(n10860));
  jxor g10587(.dina(n10860), .dinb(n10364), .dout(n10861));
  jand g10588(.dina(n10850), .dinb(n4499), .dout(n10862));
  jand g10589(.dina(n10862), .dinb(n10855), .dout(n10863));
  jor  g10590(.dina(n10863), .dinb(n10861), .dout(n10864));
  jand g10591(.dina(n10864), .dinb(n10857), .dout(n10865));
  jor  g10592(.dina(n10865), .dinb(n4494), .dout(n10866));
  jand g10593(.dina(n10865), .dinb(n4494), .dout(n10867));
  jnot g10594(.din(n10367), .dout(n10868));
  jand g10595(.dina(asqrt[19] ), .dinb(n10868), .dout(n10869));
  jand g10596(.dina(n10869), .dinb(n10372), .dout(n10870));
  jor  g10597(.dina(n10870), .dinb(n10371), .dout(n10871));
  jand g10598(.dina(n10869), .dinb(n10373), .dout(n10872));
  jnot g10599(.din(n10872), .dout(n10873));
  jand g10600(.dina(n10873), .dinb(n10871), .dout(n10874));
  jnot g10601(.din(n10874), .dout(n10875));
  jor  g10602(.dina(n10875), .dinb(n10867), .dout(n10876));
  jand g10603(.dina(n10876), .dinb(n10866), .dout(n10877));
  jor  g10604(.dina(n10877), .dinb(n3912), .dout(n10878));
  jand g10605(.dina(n10866), .dinb(n3912), .dout(n10879));
  jand g10606(.dina(n10879), .dinb(n10876), .dout(n10880));
  jnot g10607(.din(n10375), .dout(n10881));
  jand g10608(.dina(asqrt[19] ), .dinb(n10881), .dout(n10882));
  jand g10609(.dina(n10882), .dinb(n10382), .dout(n10883));
  jor  g10610(.dina(n10883), .dinb(n10380), .dout(n10884));
  jand g10611(.dina(n10882), .dinb(n10383), .dout(n10885));
  jnot g10612(.din(n10885), .dout(n10886));
  jand g10613(.dina(n10886), .dinb(n10884), .dout(n10887));
  jnot g10614(.din(n10887), .dout(n10888));
  jor  g10615(.dina(n10888), .dinb(n10880), .dout(n10889));
  jand g10616(.dina(n10889), .dinb(n10878), .dout(n10890));
  jor  g10617(.dina(n10890), .dinb(n3907), .dout(n10891));
  jxor g10618(.dina(n10384), .dinb(n3912), .dout(n10892));
  jor  g10619(.dina(n10892), .dinb(n10701), .dout(n10893));
  jxor g10620(.dina(n10893), .dinb(n10395), .dout(n10894));
  jand g10621(.dina(n10890), .dinb(n3907), .dout(n10895));
  jor  g10622(.dina(n10895), .dinb(n10894), .dout(n10896));
  jand g10623(.dina(n10896), .dinb(n10891), .dout(n10897));
  jor  g10624(.dina(n10897), .dinb(n3376), .dout(n10898));
  jnot g10625(.din(n10400), .dout(n10899));
  jor  g10626(.dina(n10899), .dinb(n10398), .dout(n10900));
  jor  g10627(.dina(n10900), .dinb(n10701), .dout(n10901));
  jxor g10628(.dina(n10901), .dinb(n10409), .dout(n10902));
  jand g10629(.dina(n10891), .dinb(n3376), .dout(n10903));
  jand g10630(.dina(n10903), .dinb(n10896), .dout(n10904));
  jor  g10631(.dina(n10904), .dinb(n10902), .dout(n10905));
  jand g10632(.dina(n10905), .dinb(n10898), .dout(n10906));
  jor  g10633(.dina(n10906), .dinb(n3371), .dout(n10907));
  jand g10634(.dina(n10906), .dinb(n3371), .dout(n10908));
  jnot g10635(.din(n10412), .dout(n10909));
  jand g10636(.dina(asqrt[19] ), .dinb(n10909), .dout(n10910));
  jand g10637(.dina(n10910), .dinb(n10417), .dout(n10911));
  jor  g10638(.dina(n10911), .dinb(n10416), .dout(n10912));
  jand g10639(.dina(n10910), .dinb(n10418), .dout(n10913));
  jnot g10640(.din(n10913), .dout(n10914));
  jand g10641(.dina(n10914), .dinb(n10912), .dout(n10915));
  jnot g10642(.din(n10915), .dout(n10916));
  jor  g10643(.dina(n10916), .dinb(n10908), .dout(n10917));
  jand g10644(.dina(n10917), .dinb(n10907), .dout(n10918));
  jor  g10645(.dina(n10918), .dinb(n2875), .dout(n10919));
  jand g10646(.dina(n10907), .dinb(n2875), .dout(n10920));
  jand g10647(.dina(n10920), .dinb(n10917), .dout(n10921));
  jnot g10648(.din(n10420), .dout(n10922));
  jand g10649(.dina(asqrt[19] ), .dinb(n10922), .dout(n10923));
  jand g10650(.dina(n10923), .dinb(n10427), .dout(n10924));
  jor  g10651(.dina(n10924), .dinb(n10425), .dout(n10925));
  jand g10652(.dina(n10923), .dinb(n10428), .dout(n10926));
  jnot g10653(.din(n10926), .dout(n10927));
  jand g10654(.dina(n10927), .dinb(n10925), .dout(n10928));
  jnot g10655(.din(n10928), .dout(n10929));
  jor  g10656(.dina(n10929), .dinb(n10921), .dout(n10930));
  jand g10657(.dina(n10930), .dinb(n10919), .dout(n10931));
  jor  g10658(.dina(n10931), .dinb(n2870), .dout(n10932));
  jxor g10659(.dina(n10429), .dinb(n2875), .dout(n10933));
  jor  g10660(.dina(n10933), .dinb(n10701), .dout(n10934));
  jxor g10661(.dina(n10934), .dinb(n10440), .dout(n10935));
  jand g10662(.dina(n10931), .dinb(n2870), .dout(n10936));
  jor  g10663(.dina(n10936), .dinb(n10935), .dout(n10937));
  jand g10664(.dina(n10937), .dinb(n10932), .dout(n10938));
  jor  g10665(.dina(n10938), .dinb(n2425), .dout(n10939));
  jand g10666(.dina(n10932), .dinb(n2425), .dout(n10940));
  jand g10667(.dina(n10940), .dinb(n10937), .dout(n10941));
  jnot g10668(.din(n10443), .dout(n10942));
  jand g10669(.dina(asqrt[19] ), .dinb(n10942), .dout(n10943));
  jand g10670(.dina(n10943), .dinb(n10450), .dout(n10944));
  jor  g10671(.dina(n10944), .dinb(n10448), .dout(n10945));
  jand g10672(.dina(n10943), .dinb(n10451), .dout(n10946));
  jnot g10673(.din(n10946), .dout(n10947));
  jand g10674(.dina(n10947), .dinb(n10945), .dout(n10948));
  jnot g10675(.din(n10948), .dout(n10949));
  jor  g10676(.dina(n10949), .dinb(n10941), .dout(n10950));
  jand g10677(.dina(n10950), .dinb(n10939), .dout(n10951));
  jor  g10678(.dina(n10951), .dinb(n2420), .dout(n10952));
  jand g10679(.dina(n10951), .dinb(n2420), .dout(n10953));
  jor  g10680(.dina(n10953), .dinb(n10704), .dout(n10954));
  jand g10681(.dina(n10954), .dinb(n10952), .dout(n10955));
  jor  g10682(.dina(n10955), .dinb(n2010), .dout(n10956));
  jnot g10683(.din(n10459), .dout(n10957));
  jor  g10684(.dina(n10957), .dinb(n10457), .dout(n10958));
  jor  g10685(.dina(n10958), .dinb(n10701), .dout(n10959));
  jxor g10686(.dina(n10959), .dinb(n10468), .dout(n10960));
  jand g10687(.dina(n10952), .dinb(n2010), .dout(n10961));
  jand g10688(.dina(n10961), .dinb(n10954), .dout(n10962));
  jor  g10689(.dina(n10962), .dinb(n10960), .dout(n10963));
  jand g10690(.dina(n10963), .dinb(n10956), .dout(n10964));
  jor  g10691(.dina(n10964), .dinb(n2005), .dout(n10965));
  jxor g10692(.dina(n10470), .dinb(n2010), .dout(n10966));
  jor  g10693(.dina(n10966), .dinb(n10701), .dout(n10967));
  jxor g10694(.dina(n10967), .dinb(n10481), .dout(n10968));
  jand g10695(.dina(n10964), .dinb(n2005), .dout(n10969));
  jor  g10696(.dina(n10969), .dinb(n10968), .dout(n10970));
  jand g10697(.dina(n10970), .dinb(n10965), .dout(n10971));
  jor  g10698(.dina(n10971), .dinb(n1646), .dout(n10972));
  jnot g10699(.din(n10486), .dout(n10973));
  jor  g10700(.dina(n10973), .dinb(n10484), .dout(n10974));
  jor  g10701(.dina(n10974), .dinb(n10701), .dout(n10975));
  jxor g10702(.dina(n10975), .dinb(n10495), .dout(n10976));
  jand g10703(.dina(n10965), .dinb(n1646), .dout(n10977));
  jand g10704(.dina(n10977), .dinb(n10970), .dout(n10978));
  jor  g10705(.dina(n10978), .dinb(n10976), .dout(n10979));
  jand g10706(.dina(n10979), .dinb(n10972), .dout(n10980));
  jor  g10707(.dina(n10980), .dinb(n1641), .dout(n10981));
  jand g10708(.dina(n10980), .dinb(n1641), .dout(n10982));
  jnot g10709(.din(n10498), .dout(n10983));
  jand g10710(.dina(asqrt[19] ), .dinb(n10983), .dout(n10984));
  jand g10711(.dina(n10984), .dinb(n10503), .dout(n10985));
  jor  g10712(.dina(n10985), .dinb(n10502), .dout(n10986));
  jand g10713(.dina(n10984), .dinb(n10504), .dout(n10987));
  jnot g10714(.din(n10987), .dout(n10988));
  jand g10715(.dina(n10988), .dinb(n10986), .dout(n10989));
  jnot g10716(.din(n10989), .dout(n10990));
  jor  g10717(.dina(n10990), .dinb(n10982), .dout(n10991));
  jand g10718(.dina(n10991), .dinb(n10981), .dout(n10992));
  jor  g10719(.dina(n10992), .dinb(n1317), .dout(n10993));
  jand g10720(.dina(n10981), .dinb(n1317), .dout(n10994));
  jand g10721(.dina(n10994), .dinb(n10991), .dout(n10995));
  jnot g10722(.din(n10506), .dout(n10996));
  jand g10723(.dina(asqrt[19] ), .dinb(n10996), .dout(n10997));
  jand g10724(.dina(n10997), .dinb(n10513), .dout(n10998));
  jor  g10725(.dina(n10998), .dinb(n10511), .dout(n10999));
  jand g10726(.dina(n10997), .dinb(n10514), .dout(n11000));
  jnot g10727(.din(n11000), .dout(n11001));
  jand g10728(.dina(n11001), .dinb(n10999), .dout(n11002));
  jnot g10729(.din(n11002), .dout(n11003));
  jor  g10730(.dina(n11003), .dinb(n10995), .dout(n11004));
  jand g10731(.dina(n11004), .dinb(n10993), .dout(n11005));
  jor  g10732(.dina(n11005), .dinb(n1312), .dout(n11006));
  jxor g10733(.dina(n10515), .dinb(n1317), .dout(n11007));
  jor  g10734(.dina(n11007), .dinb(n10701), .dout(n11008));
  jxor g10735(.dina(n11008), .dinb(n10526), .dout(n11009));
  jand g10736(.dina(n11005), .dinb(n1312), .dout(n11010));
  jor  g10737(.dina(n11010), .dinb(n11009), .dout(n11011));
  jand g10738(.dina(n11011), .dinb(n11006), .dout(n11012));
  jor  g10739(.dina(n11012), .dinb(n1039), .dout(n11013));
  jnot g10740(.din(n10531), .dout(n11014));
  jor  g10741(.dina(n11014), .dinb(n10529), .dout(n11015));
  jor  g10742(.dina(n11015), .dinb(n10701), .dout(n11016));
  jxor g10743(.dina(n11016), .dinb(n10540), .dout(n11017));
  jand g10744(.dina(n11006), .dinb(n1039), .dout(n11018));
  jand g10745(.dina(n11018), .dinb(n11011), .dout(n11019));
  jor  g10746(.dina(n11019), .dinb(n11017), .dout(n11020));
  jand g10747(.dina(n11020), .dinb(n11013), .dout(n11021));
  jor  g10748(.dina(n11021), .dinb(n1034), .dout(n11022));
  jand g10749(.dina(n11021), .dinb(n1034), .dout(n11023));
  jnot g10750(.din(n10543), .dout(n11024));
  jand g10751(.dina(asqrt[19] ), .dinb(n11024), .dout(n11025));
  jand g10752(.dina(n11025), .dinb(n10548), .dout(n11026));
  jor  g10753(.dina(n11026), .dinb(n10547), .dout(n11027));
  jand g10754(.dina(n11025), .dinb(n10549), .dout(n11028));
  jnot g10755(.din(n11028), .dout(n11029));
  jand g10756(.dina(n11029), .dinb(n11027), .dout(n11030));
  jnot g10757(.din(n11030), .dout(n11031));
  jor  g10758(.dina(n11031), .dinb(n11023), .dout(n11032));
  jand g10759(.dina(n11032), .dinb(n11022), .dout(n11033));
  jor  g10760(.dina(n11033), .dinb(n796), .dout(n11034));
  jand g10761(.dina(n11022), .dinb(n796), .dout(n11035));
  jand g10762(.dina(n11035), .dinb(n11032), .dout(n11036));
  jnot g10763(.din(n10551), .dout(n11037));
  jand g10764(.dina(asqrt[19] ), .dinb(n11037), .dout(n11038));
  jand g10765(.dina(n11038), .dinb(n10558), .dout(n11039));
  jor  g10766(.dina(n11039), .dinb(n10556), .dout(n11040));
  jand g10767(.dina(n11038), .dinb(n10559), .dout(n11041));
  jnot g10768(.din(n11041), .dout(n11042));
  jand g10769(.dina(n11042), .dinb(n11040), .dout(n11043));
  jnot g10770(.din(n11043), .dout(n11044));
  jor  g10771(.dina(n11044), .dinb(n11036), .dout(n11045));
  jand g10772(.dina(n11045), .dinb(n11034), .dout(n11046));
  jor  g10773(.dina(n11046), .dinb(n791), .dout(n11047));
  jxor g10774(.dina(n10560), .dinb(n796), .dout(n11048));
  jor  g10775(.dina(n11048), .dinb(n10701), .dout(n11049));
  jxor g10776(.dina(n11049), .dinb(n10571), .dout(n11050));
  jand g10777(.dina(n11046), .dinb(n791), .dout(n11051));
  jor  g10778(.dina(n11051), .dinb(n11050), .dout(n11052));
  jand g10779(.dina(n11052), .dinb(n11047), .dout(n11053));
  jor  g10780(.dina(n11053), .dinb(n595), .dout(n11054));
  jnot g10781(.din(n10576), .dout(n11055));
  jor  g10782(.dina(n11055), .dinb(n10574), .dout(n11056));
  jor  g10783(.dina(n11056), .dinb(n10701), .dout(n11057));
  jxor g10784(.dina(n11057), .dinb(n10585), .dout(n11058));
  jand g10785(.dina(n11047), .dinb(n595), .dout(n11059));
  jand g10786(.dina(n11059), .dinb(n11052), .dout(n11060));
  jor  g10787(.dina(n11060), .dinb(n11058), .dout(n11061));
  jand g10788(.dina(n11061), .dinb(n11054), .dout(n11062));
  jor  g10789(.dina(n11062), .dinb(n590), .dout(n11063));
  jand g10790(.dina(n11062), .dinb(n590), .dout(n11064));
  jnot g10791(.din(n10588), .dout(n11065));
  jand g10792(.dina(asqrt[19] ), .dinb(n11065), .dout(n11066));
  jand g10793(.dina(n11066), .dinb(n10593), .dout(n11067));
  jor  g10794(.dina(n11067), .dinb(n10592), .dout(n11068));
  jand g10795(.dina(n11066), .dinb(n10594), .dout(n11069));
  jnot g10796(.din(n11069), .dout(n11070));
  jand g10797(.dina(n11070), .dinb(n11068), .dout(n11071));
  jnot g10798(.din(n11071), .dout(n11072));
  jor  g10799(.dina(n11072), .dinb(n11064), .dout(n11073));
  jand g10800(.dina(n11073), .dinb(n11063), .dout(n11074));
  jor  g10801(.dina(n11074), .dinb(n430), .dout(n11075));
  jand g10802(.dina(n11063), .dinb(n430), .dout(n11076));
  jand g10803(.dina(n11076), .dinb(n11073), .dout(n11077));
  jnot g10804(.din(n10596), .dout(n11078));
  jand g10805(.dina(asqrt[19] ), .dinb(n11078), .dout(n11079));
  jand g10806(.dina(n11079), .dinb(n10603), .dout(n11080));
  jor  g10807(.dina(n11080), .dinb(n10601), .dout(n11081));
  jand g10808(.dina(n11079), .dinb(n10604), .dout(n11082));
  jnot g10809(.din(n11082), .dout(n11083));
  jand g10810(.dina(n11083), .dinb(n11081), .dout(n11084));
  jnot g10811(.din(n11084), .dout(n11085));
  jor  g10812(.dina(n11085), .dinb(n11077), .dout(n11086));
  jand g10813(.dina(n11086), .dinb(n11075), .dout(n11087));
  jor  g10814(.dina(n11087), .dinb(n425), .dout(n11088));
  jxor g10815(.dina(n10605), .dinb(n430), .dout(n11089));
  jor  g10816(.dina(n11089), .dinb(n10701), .dout(n11090));
  jxor g10817(.dina(n11090), .dinb(n10616), .dout(n11091));
  jand g10818(.dina(n11087), .dinb(n425), .dout(n11092));
  jor  g10819(.dina(n11092), .dinb(n11091), .dout(n11093));
  jand g10820(.dina(n11093), .dinb(n11088), .dout(n11094));
  jor  g10821(.dina(n11094), .dinb(n305), .dout(n11095));
  jnot g10822(.din(n10621), .dout(n11096));
  jor  g10823(.dina(n11096), .dinb(n10619), .dout(n11097));
  jor  g10824(.dina(n11097), .dinb(n10701), .dout(n11098));
  jxor g10825(.dina(n11098), .dinb(n10630), .dout(n11099));
  jand g10826(.dina(n11088), .dinb(n305), .dout(n11100));
  jand g10827(.dina(n11100), .dinb(n11093), .dout(n11101));
  jor  g10828(.dina(n11101), .dinb(n11099), .dout(n11102));
  jand g10829(.dina(n11102), .dinb(n11095), .dout(n11103));
  jor  g10830(.dina(n11103), .dinb(n290), .dout(n11104));
  jand g10831(.dina(n11103), .dinb(n290), .dout(n11105));
  jnot g10832(.din(n10633), .dout(n11106));
  jand g10833(.dina(asqrt[19] ), .dinb(n11106), .dout(n11107));
  jand g10834(.dina(n11107), .dinb(n10638), .dout(n11108));
  jor  g10835(.dina(n11108), .dinb(n10637), .dout(n11109));
  jand g10836(.dina(n11107), .dinb(n10639), .dout(n11110));
  jnot g10837(.din(n11110), .dout(n11111));
  jand g10838(.dina(n11111), .dinb(n11109), .dout(n11112));
  jnot g10839(.din(n11112), .dout(n11113));
  jor  g10840(.dina(n11113), .dinb(n11105), .dout(n11114));
  jand g10841(.dina(n11114), .dinb(n11104), .dout(n11115));
  jor  g10842(.dina(n11115), .dinb(n223), .dout(n11116));
  jand g10843(.dina(n11104), .dinb(n223), .dout(n11117));
  jand g10844(.dina(n11117), .dinb(n11114), .dout(n11118));
  jnot g10845(.din(n10641), .dout(n11119));
  jand g10846(.dina(asqrt[19] ), .dinb(n11119), .dout(n11120));
  jand g10847(.dina(n11120), .dinb(n10648), .dout(n11121));
  jor  g10848(.dina(n11121), .dinb(n10646), .dout(n11122));
  jand g10849(.dina(n11120), .dinb(n10649), .dout(n11123));
  jnot g10850(.din(n11123), .dout(n11124));
  jand g10851(.dina(n11124), .dinb(n11122), .dout(n11125));
  jnot g10852(.din(n11125), .dout(n11126));
  jor  g10853(.dina(n11126), .dinb(n11118), .dout(n11127));
  jand g10854(.dina(n11127), .dinb(n11116), .dout(n11128));
  jor  g10855(.dina(n11128), .dinb(n199), .dout(n11129));
  jand g10856(.dina(n11128), .dinb(n199), .dout(n11130));
  jxor g10857(.dina(n10650), .dinb(n223), .dout(n11131));
  jor  g10858(.dina(n11131), .dinb(n10701), .dout(n11132));
  jxor g10859(.dina(n11132), .dinb(n10661), .dout(n11133));
  jor  g10860(.dina(n11133), .dinb(n11130), .dout(n11134));
  jand g10861(.dina(n11134), .dinb(n11129), .dout(n11135));
  jnot g10862(.din(n10666), .dout(n11136));
  jor  g10863(.dina(n11136), .dinb(n10664), .dout(n11137));
  jor  g10864(.dina(n11137), .dinb(n10701), .dout(n11138));
  jxor g10865(.dina(n11138), .dinb(n10675), .dout(n11139));
  jand g10866(.dina(asqrt[19] ), .dinb(n10689), .dout(n11140));
  jand g10867(.dina(n11140), .dinb(n10677), .dout(n11141));
  jor  g10868(.dina(n11141), .dinb(n10723), .dout(n11142));
  jor  g10869(.dina(n11142), .dinb(n11139), .dout(n11143));
  jor  g10870(.dina(n11143), .dinb(n11135), .dout(n11144));
  jand g10871(.dina(n11144), .dinb(n194), .dout(n11145));
  jand g10872(.dina(n11139), .dinb(n11135), .dout(n11146));
  jor  g10873(.dina(n11140), .dinb(n10677), .dout(n11147));
  jand g10874(.dina(n10689), .dinb(n10677), .dout(n11148));
  jor  g10875(.dina(n11148), .dinb(n194), .dout(n11149));
  jnot g10876(.din(n11149), .dout(n11150));
  jand g10877(.dina(n11150), .dinb(n11147), .dout(n11151));
  jor  g10878(.dina(n11151), .dinb(n11146), .dout(n11154));
  jor  g10879(.dina(n11154), .dinb(n11145), .dout(asqrt[18] ));
  jxor g10880(.dina(n10951), .dinb(n2420), .dout(n11156));
  jand g10881(.dina(n11156), .dinb(asqrt[18] ), .dout(n11157));
  jxor g10882(.dina(n11157), .dinb(n10704), .dout(n11158));
  jand g10883(.dina(asqrt[18] ), .dinb(a[36] ), .dout(n11159));
  jnot g10884(.din(a[34] ), .dout(n11160));
  jnot g10885(.din(a[35] ), .dout(n11161));
  jand g10886(.dina(n10706), .dinb(n11161), .dout(n11162));
  jand g10887(.dina(n11162), .dinb(n11160), .dout(n11163));
  jor  g10888(.dina(n11163), .dinb(n11159), .dout(n11164));
  jand g10889(.dina(n11164), .dinb(asqrt[19] ), .dout(n11165));
  jand g10890(.dina(asqrt[18] ), .dinb(n10706), .dout(n11166));
  jxor g10891(.dina(n11166), .dinb(n10707), .dout(n11167));
  jor  g10892(.dina(n11164), .dinb(asqrt[19] ), .dout(n11168));
  jand g10893(.dina(n11168), .dinb(n11167), .dout(n11169));
  jor  g10894(.dina(n11169), .dinb(n11165), .dout(n11170));
  jand g10895(.dina(n11170), .dinb(asqrt[20] ), .dout(n11171));
  jor  g10896(.dina(n11165), .dinb(asqrt[20] ), .dout(n11172));
  jor  g10897(.dina(n11172), .dinb(n11169), .dout(n11173));
  jand g10898(.dina(n11166), .dinb(n10707), .dout(n11174));
  jnot g10899(.din(n11145), .dout(n11175));
  jnot g10900(.din(n11146), .dout(n11176));
  jnot g10901(.din(n11151), .dout(n11177));
  jand g10902(.dina(n11177), .dinb(asqrt[19] ), .dout(n11178));
  jand g10903(.dina(n11178), .dinb(n11176), .dout(n11179));
  jand g10904(.dina(n11179), .dinb(n11175), .dout(n11180));
  jor  g10905(.dina(n11180), .dinb(n11174), .dout(n11181));
  jxor g10906(.dina(n11181), .dinb(n10219), .dout(n11182));
  jand g10907(.dina(n11182), .dinb(n11173), .dout(n11183));
  jor  g10908(.dina(n11183), .dinb(n11171), .dout(n11184));
  jand g10909(.dina(n11184), .dinb(asqrt[21] ), .dout(n11185));
  jor  g10910(.dina(n11184), .dinb(asqrt[21] ), .dout(n11186));
  jxor g10911(.dina(n10711), .dinb(n10696), .dout(n11187));
  jand g10912(.dina(n11187), .dinb(asqrt[18] ), .dout(n11188));
  jxor g10913(.dina(n11188), .dinb(n10714), .dout(n11189));
  jnot g10914(.din(n11189), .dout(n11190));
  jand g10915(.dina(n11190), .dinb(n11186), .dout(n11191));
  jor  g10916(.dina(n11191), .dinb(n11185), .dout(n11192));
  jand g10917(.dina(n11192), .dinb(asqrt[22] ), .dout(n11193));
  jnot g10918(.din(n10720), .dout(n11194));
  jand g10919(.dina(n11194), .dinb(n10718), .dout(n11195));
  jand g10920(.dina(n11195), .dinb(asqrt[18] ), .dout(n11196));
  jxor g10921(.dina(n11196), .dinb(n10728), .dout(n11197));
  jnot g10922(.din(n11197), .dout(n11198));
  jor  g10923(.dina(n11185), .dinb(asqrt[22] ), .dout(n11199));
  jor  g10924(.dina(n11199), .dinb(n11191), .dout(n11200));
  jand g10925(.dina(n11200), .dinb(n11198), .dout(n11201));
  jor  g10926(.dina(n11201), .dinb(n11193), .dout(n11202));
  jand g10927(.dina(n11202), .dinb(asqrt[23] ), .dout(n11203));
  jor  g10928(.dina(n11202), .dinb(asqrt[23] ), .dout(n11204));
  jnot g10929(.din(n10735), .dout(n11205));
  jxor g10930(.dina(n10730), .dinb(n9769), .dout(n11206));
  jand g10931(.dina(n11206), .dinb(asqrt[18] ), .dout(n11207));
  jxor g10932(.dina(n11207), .dinb(n11205), .dout(n11208));
  jand g10933(.dina(n11208), .dinb(n11204), .dout(n11209));
  jor  g10934(.dina(n11209), .dinb(n11203), .dout(n11210));
  jand g10935(.dina(n11210), .dinb(asqrt[24] ), .dout(n11211));
  jor  g10936(.dina(n11203), .dinb(asqrt[24] ), .dout(n11212));
  jor  g10937(.dina(n11212), .dinb(n11209), .dout(n11213));
  jnot g10938(.din(n10742), .dout(n11214));
  jnot g10939(.din(n10744), .dout(n11215));
  jand g10940(.dina(asqrt[18] ), .dinb(n10738), .dout(n11216));
  jand g10941(.dina(n11216), .dinb(n11215), .dout(n11217));
  jor  g10942(.dina(n11217), .dinb(n11214), .dout(n11218));
  jnot g10943(.din(n10745), .dout(n11219));
  jand g10944(.dina(n11216), .dinb(n11219), .dout(n11220));
  jnot g10945(.din(n11220), .dout(n11221));
  jand g10946(.dina(n11221), .dinb(n11218), .dout(n11222));
  jand g10947(.dina(n11222), .dinb(n11213), .dout(n11223));
  jor  g10948(.dina(n11223), .dinb(n11211), .dout(n11224));
  jand g10949(.dina(n11224), .dinb(asqrt[25] ), .dout(n11225));
  jor  g10950(.dina(n11224), .dinb(asqrt[25] ), .dout(n11226));
  jxor g10951(.dina(n10746), .dinb(n8893), .dout(n11227));
  jand g10952(.dina(n11227), .dinb(asqrt[18] ), .dout(n11228));
  jxor g10953(.dina(n11228), .dinb(n10751), .dout(n11229));
  jand g10954(.dina(n11229), .dinb(n11226), .dout(n11230));
  jor  g10955(.dina(n11230), .dinb(n11225), .dout(n11231));
  jand g10956(.dina(n11231), .dinb(asqrt[26] ), .dout(n11232));
  jnot g10957(.din(n10757), .dout(n11233));
  jand g10958(.dina(n11233), .dinb(n10755), .dout(n11234));
  jand g10959(.dina(n11234), .dinb(asqrt[18] ), .dout(n11235));
  jxor g10960(.dina(n11235), .dinb(n10766), .dout(n11236));
  jnot g10961(.din(n11236), .dout(n11237));
  jor  g10962(.dina(n11225), .dinb(asqrt[26] ), .dout(n11238));
  jor  g10963(.dina(n11238), .dinb(n11230), .dout(n11239));
  jand g10964(.dina(n11239), .dinb(n11237), .dout(n11240));
  jor  g10965(.dina(n11240), .dinb(n11232), .dout(n11241));
  jand g10966(.dina(n11241), .dinb(asqrt[27] ), .dout(n11242));
  jor  g10967(.dina(n11241), .dinb(asqrt[27] ), .dout(n11243));
  jxor g10968(.dina(n10768), .dinb(n8053), .dout(n11244));
  jand g10969(.dina(n11244), .dinb(asqrt[18] ), .dout(n11245));
  jxor g10970(.dina(n11245), .dinb(n10774), .dout(n11246));
  jand g10971(.dina(n11246), .dinb(n11243), .dout(n11247));
  jor  g10972(.dina(n11247), .dinb(n11242), .dout(n11248));
  jand g10973(.dina(n11248), .dinb(asqrt[28] ), .dout(n11249));
  jor  g10974(.dina(n11242), .dinb(asqrt[28] ), .dout(n11250));
  jor  g10975(.dina(n11250), .dinb(n11247), .dout(n11251));
  jnot g10976(.din(n10782), .dout(n11252));
  jnot g10977(.din(n10784), .dout(n11253));
  jand g10978(.dina(asqrt[18] ), .dinb(n10778), .dout(n11254));
  jand g10979(.dina(n11254), .dinb(n11253), .dout(n11255));
  jor  g10980(.dina(n11255), .dinb(n11252), .dout(n11256));
  jnot g10981(.din(n10785), .dout(n11257));
  jand g10982(.dina(n11254), .dinb(n11257), .dout(n11258));
  jnot g10983(.din(n11258), .dout(n11259));
  jand g10984(.dina(n11259), .dinb(n11256), .dout(n11260));
  jand g10985(.dina(n11260), .dinb(n11251), .dout(n11261));
  jor  g10986(.dina(n11261), .dinb(n11249), .dout(n11262));
  jand g10987(.dina(n11262), .dinb(asqrt[29] ), .dout(n11263));
  jxor g10988(.dina(n10786), .dinb(n7260), .dout(n11264));
  jand g10989(.dina(n11264), .dinb(asqrt[18] ), .dout(n11265));
  jxor g10990(.dina(n11265), .dinb(n10793), .dout(n11266));
  jnot g10991(.din(n11266), .dout(n11267));
  jor  g10992(.dina(n11262), .dinb(asqrt[29] ), .dout(n11268));
  jand g10993(.dina(n11268), .dinb(n11267), .dout(n11269));
  jor  g10994(.dina(n11269), .dinb(n11263), .dout(n11270));
  jand g10995(.dina(n11270), .dinb(asqrt[30] ), .dout(n11271));
  jnot g10996(.din(n10798), .dout(n11272));
  jand g10997(.dina(n11272), .dinb(n10796), .dout(n11273));
  jand g10998(.dina(n11273), .dinb(asqrt[18] ), .dout(n11274));
  jxor g10999(.dina(n11274), .dinb(n10806), .dout(n11275));
  jnot g11000(.din(n11275), .dout(n11276));
  jor  g11001(.dina(n11263), .dinb(asqrt[30] ), .dout(n11277));
  jor  g11002(.dina(n11277), .dinb(n11269), .dout(n11278));
  jand g11003(.dina(n11278), .dinb(n11276), .dout(n11279));
  jor  g11004(.dina(n11279), .dinb(n11271), .dout(n11280));
  jand g11005(.dina(n11280), .dinb(asqrt[31] ), .dout(n11281));
  jor  g11006(.dina(n11280), .dinb(asqrt[31] ), .dout(n11282));
  jnot g11007(.din(n10812), .dout(n11283));
  jnot g11008(.din(n10813), .dout(n11284));
  jand g11009(.dina(asqrt[18] ), .dinb(n10809), .dout(n11285));
  jand g11010(.dina(n11285), .dinb(n11284), .dout(n11286));
  jor  g11011(.dina(n11286), .dinb(n11283), .dout(n11287));
  jnot g11012(.din(n10814), .dout(n11288));
  jand g11013(.dina(n11285), .dinb(n11288), .dout(n11289));
  jnot g11014(.din(n11289), .dout(n11290));
  jand g11015(.dina(n11290), .dinb(n11287), .dout(n11291));
  jand g11016(.dina(n11291), .dinb(n11282), .dout(n11292));
  jor  g11017(.dina(n11292), .dinb(n11281), .dout(n11293));
  jand g11018(.dina(n11293), .dinb(asqrt[32] ), .dout(n11294));
  jor  g11019(.dina(n11281), .dinb(asqrt[32] ), .dout(n11295));
  jor  g11020(.dina(n11295), .dinb(n11292), .dout(n11296));
  jnot g11021(.din(n10820), .dout(n11297));
  jnot g11022(.din(n10822), .dout(n11298));
  jand g11023(.dina(asqrt[18] ), .dinb(n10816), .dout(n11299));
  jand g11024(.dina(n11299), .dinb(n11298), .dout(n11300));
  jor  g11025(.dina(n11300), .dinb(n11297), .dout(n11301));
  jnot g11026(.din(n10823), .dout(n11302));
  jand g11027(.dina(n11299), .dinb(n11302), .dout(n11303));
  jnot g11028(.din(n11303), .dout(n11304));
  jand g11029(.dina(n11304), .dinb(n11301), .dout(n11305));
  jand g11030(.dina(n11305), .dinb(n11296), .dout(n11306));
  jor  g11031(.dina(n11306), .dinb(n11294), .dout(n11307));
  jand g11032(.dina(n11307), .dinb(asqrt[33] ), .dout(n11308));
  jxor g11033(.dina(n10824), .dinb(n5788), .dout(n11309));
  jand g11034(.dina(n11309), .dinb(asqrt[18] ), .dout(n11310));
  jxor g11035(.dina(n11310), .dinb(n10834), .dout(n11311));
  jnot g11036(.din(n11311), .dout(n11312));
  jor  g11037(.dina(n11307), .dinb(asqrt[33] ), .dout(n11313));
  jand g11038(.dina(n11313), .dinb(n11312), .dout(n11314));
  jor  g11039(.dina(n11314), .dinb(n11308), .dout(n11315));
  jand g11040(.dina(n11315), .dinb(asqrt[34] ), .dout(n11316));
  jnot g11041(.din(n10839), .dout(n11317));
  jand g11042(.dina(n11317), .dinb(n10837), .dout(n11318));
  jand g11043(.dina(n11318), .dinb(asqrt[18] ), .dout(n11319));
  jxor g11044(.dina(n11319), .dinb(n10847), .dout(n11320));
  jnot g11045(.din(n11320), .dout(n11321));
  jor  g11046(.dina(n11308), .dinb(asqrt[34] ), .dout(n11322));
  jor  g11047(.dina(n11322), .dinb(n11314), .dout(n11323));
  jand g11048(.dina(n11323), .dinb(n11321), .dout(n11324));
  jor  g11049(.dina(n11324), .dinb(n11316), .dout(n11325));
  jand g11050(.dina(n11325), .dinb(asqrt[35] ), .dout(n11326));
  jor  g11051(.dina(n11325), .dinb(asqrt[35] ), .dout(n11327));
  jnot g11052(.din(n10853), .dout(n11328));
  jnot g11053(.din(n10854), .dout(n11329));
  jand g11054(.dina(asqrt[18] ), .dinb(n10850), .dout(n11330));
  jand g11055(.dina(n11330), .dinb(n11329), .dout(n11331));
  jor  g11056(.dina(n11331), .dinb(n11328), .dout(n11332));
  jnot g11057(.din(n10855), .dout(n11333));
  jand g11058(.dina(n11330), .dinb(n11333), .dout(n11334));
  jnot g11059(.din(n11334), .dout(n11335));
  jand g11060(.dina(n11335), .dinb(n11332), .dout(n11336));
  jand g11061(.dina(n11336), .dinb(n11327), .dout(n11337));
  jor  g11062(.dina(n11337), .dinb(n11326), .dout(n11338));
  jand g11063(.dina(n11338), .dinb(asqrt[36] ), .dout(n11339));
  jor  g11064(.dina(n11326), .dinb(asqrt[36] ), .dout(n11340));
  jor  g11065(.dina(n11340), .dinb(n11337), .dout(n11341));
  jnot g11066(.din(n10861), .dout(n11342));
  jnot g11067(.din(n10863), .dout(n11343));
  jand g11068(.dina(asqrt[18] ), .dinb(n10857), .dout(n11344));
  jand g11069(.dina(n11344), .dinb(n11343), .dout(n11345));
  jor  g11070(.dina(n11345), .dinb(n11342), .dout(n11346));
  jnot g11071(.din(n10864), .dout(n11347));
  jand g11072(.dina(n11344), .dinb(n11347), .dout(n11348));
  jnot g11073(.din(n11348), .dout(n11349));
  jand g11074(.dina(n11349), .dinb(n11346), .dout(n11350));
  jand g11075(.dina(n11350), .dinb(n11341), .dout(n11351));
  jor  g11076(.dina(n11351), .dinb(n11339), .dout(n11352));
  jand g11077(.dina(n11352), .dinb(asqrt[37] ), .dout(n11353));
  jxor g11078(.dina(n10865), .dinb(n4494), .dout(n11354));
  jand g11079(.dina(n11354), .dinb(asqrt[18] ), .dout(n11355));
  jxor g11080(.dina(n11355), .dinb(n10875), .dout(n11356));
  jnot g11081(.din(n11356), .dout(n11357));
  jor  g11082(.dina(n11352), .dinb(asqrt[37] ), .dout(n11358));
  jand g11083(.dina(n11358), .dinb(n11357), .dout(n11359));
  jor  g11084(.dina(n11359), .dinb(n11353), .dout(n11360));
  jand g11085(.dina(n11360), .dinb(asqrt[38] ), .dout(n11361));
  jnot g11086(.din(n10880), .dout(n11362));
  jand g11087(.dina(n11362), .dinb(n10878), .dout(n11363));
  jand g11088(.dina(n11363), .dinb(asqrt[18] ), .dout(n11364));
  jxor g11089(.dina(n11364), .dinb(n10888), .dout(n11365));
  jnot g11090(.din(n11365), .dout(n11366));
  jor  g11091(.dina(n11353), .dinb(asqrt[38] ), .dout(n11367));
  jor  g11092(.dina(n11367), .dinb(n11359), .dout(n11368));
  jand g11093(.dina(n11368), .dinb(n11366), .dout(n11369));
  jor  g11094(.dina(n11369), .dinb(n11361), .dout(n11370));
  jand g11095(.dina(n11370), .dinb(asqrt[39] ), .dout(n11371));
  jor  g11096(.dina(n11370), .dinb(asqrt[39] ), .dout(n11372));
  jnot g11097(.din(n10894), .dout(n11373));
  jnot g11098(.din(n10895), .dout(n11374));
  jand g11099(.dina(asqrt[18] ), .dinb(n10891), .dout(n11375));
  jand g11100(.dina(n11375), .dinb(n11374), .dout(n11376));
  jor  g11101(.dina(n11376), .dinb(n11373), .dout(n11377));
  jnot g11102(.din(n10896), .dout(n11378));
  jand g11103(.dina(n11375), .dinb(n11378), .dout(n11379));
  jnot g11104(.din(n11379), .dout(n11380));
  jand g11105(.dina(n11380), .dinb(n11377), .dout(n11381));
  jand g11106(.dina(n11381), .dinb(n11372), .dout(n11382));
  jor  g11107(.dina(n11382), .dinb(n11371), .dout(n11383));
  jand g11108(.dina(n11383), .dinb(asqrt[40] ), .dout(n11384));
  jor  g11109(.dina(n11371), .dinb(asqrt[40] ), .dout(n11385));
  jor  g11110(.dina(n11385), .dinb(n11382), .dout(n11386));
  jnot g11111(.din(n10902), .dout(n11387));
  jnot g11112(.din(n10904), .dout(n11388));
  jand g11113(.dina(asqrt[18] ), .dinb(n10898), .dout(n11389));
  jand g11114(.dina(n11389), .dinb(n11388), .dout(n11390));
  jor  g11115(.dina(n11390), .dinb(n11387), .dout(n11391));
  jnot g11116(.din(n10905), .dout(n11392));
  jand g11117(.dina(n11389), .dinb(n11392), .dout(n11393));
  jnot g11118(.din(n11393), .dout(n11394));
  jand g11119(.dina(n11394), .dinb(n11391), .dout(n11395));
  jand g11120(.dina(n11395), .dinb(n11386), .dout(n11396));
  jor  g11121(.dina(n11396), .dinb(n11384), .dout(n11397));
  jand g11122(.dina(n11397), .dinb(asqrt[41] ), .dout(n11398));
  jxor g11123(.dina(n10906), .dinb(n3371), .dout(n11399));
  jand g11124(.dina(n11399), .dinb(asqrt[18] ), .dout(n11400));
  jxor g11125(.dina(n11400), .dinb(n10916), .dout(n11401));
  jnot g11126(.din(n11401), .dout(n11402));
  jor  g11127(.dina(n11397), .dinb(asqrt[41] ), .dout(n11403));
  jand g11128(.dina(n11403), .dinb(n11402), .dout(n11404));
  jor  g11129(.dina(n11404), .dinb(n11398), .dout(n11405));
  jand g11130(.dina(n11405), .dinb(asqrt[42] ), .dout(n11406));
  jnot g11131(.din(n10921), .dout(n11407));
  jand g11132(.dina(n11407), .dinb(n10919), .dout(n11408));
  jand g11133(.dina(n11408), .dinb(asqrt[18] ), .dout(n11409));
  jxor g11134(.dina(n11409), .dinb(n10929), .dout(n11410));
  jnot g11135(.din(n11410), .dout(n11411));
  jor  g11136(.dina(n11398), .dinb(asqrt[42] ), .dout(n11412));
  jor  g11137(.dina(n11412), .dinb(n11404), .dout(n11413));
  jand g11138(.dina(n11413), .dinb(n11411), .dout(n11414));
  jor  g11139(.dina(n11414), .dinb(n11406), .dout(n11415));
  jand g11140(.dina(n11415), .dinb(asqrt[43] ), .dout(n11416));
  jor  g11141(.dina(n11415), .dinb(asqrt[43] ), .dout(n11417));
  jnot g11142(.din(n10935), .dout(n11418));
  jnot g11143(.din(n10936), .dout(n11419));
  jand g11144(.dina(asqrt[18] ), .dinb(n10932), .dout(n11420));
  jand g11145(.dina(n11420), .dinb(n11419), .dout(n11421));
  jor  g11146(.dina(n11421), .dinb(n11418), .dout(n11422));
  jnot g11147(.din(n10937), .dout(n11423));
  jand g11148(.dina(n11420), .dinb(n11423), .dout(n11424));
  jnot g11149(.din(n11424), .dout(n11425));
  jand g11150(.dina(n11425), .dinb(n11422), .dout(n11426));
  jand g11151(.dina(n11426), .dinb(n11417), .dout(n11427));
  jor  g11152(.dina(n11427), .dinb(n11416), .dout(n11428));
  jand g11153(.dina(n11428), .dinb(asqrt[44] ), .dout(n11429));
  jnot g11154(.din(n10941), .dout(n11430));
  jand g11155(.dina(n11430), .dinb(n10939), .dout(n11431));
  jand g11156(.dina(n11431), .dinb(asqrt[18] ), .dout(n11432));
  jxor g11157(.dina(n11432), .dinb(n10949), .dout(n11433));
  jnot g11158(.din(n11433), .dout(n11434));
  jor  g11159(.dina(n11416), .dinb(asqrt[44] ), .dout(n11435));
  jor  g11160(.dina(n11435), .dinb(n11427), .dout(n11436));
  jand g11161(.dina(n11436), .dinb(n11434), .dout(n11437));
  jor  g11162(.dina(n11437), .dinb(n11429), .dout(n11438));
  jand g11163(.dina(n11438), .dinb(asqrt[45] ), .dout(n11439));
  jnot g11164(.din(n11158), .dout(n11440));
  jor  g11165(.dina(n11438), .dinb(asqrt[45] ), .dout(n11441));
  jand g11166(.dina(n11441), .dinb(n11440), .dout(n11442));
  jor  g11167(.dina(n11442), .dinb(n11439), .dout(n11443));
  jand g11168(.dina(n11443), .dinb(asqrt[46] ), .dout(n11444));
  jor  g11169(.dina(n11439), .dinb(asqrt[46] ), .dout(n11445));
  jor  g11170(.dina(n11445), .dinb(n11442), .dout(n11446));
  jnot g11171(.din(n10960), .dout(n11447));
  jnot g11172(.din(n10962), .dout(n11448));
  jand g11173(.dina(asqrt[18] ), .dinb(n10956), .dout(n11449));
  jand g11174(.dina(n11449), .dinb(n11448), .dout(n11450));
  jor  g11175(.dina(n11450), .dinb(n11447), .dout(n11451));
  jnot g11176(.din(n10963), .dout(n11452));
  jand g11177(.dina(n11449), .dinb(n11452), .dout(n11453));
  jnot g11178(.din(n11453), .dout(n11454));
  jand g11179(.dina(n11454), .dinb(n11451), .dout(n11455));
  jand g11180(.dina(n11455), .dinb(n11446), .dout(n11456));
  jor  g11181(.dina(n11456), .dinb(n11444), .dout(n11457));
  jand g11182(.dina(n11457), .dinb(asqrt[47] ), .dout(n11458));
  jor  g11183(.dina(n11457), .dinb(asqrt[47] ), .dout(n11459));
  jnot g11184(.din(n10968), .dout(n11460));
  jnot g11185(.din(n10969), .dout(n11461));
  jand g11186(.dina(asqrt[18] ), .dinb(n10965), .dout(n11462));
  jand g11187(.dina(n11462), .dinb(n11461), .dout(n11463));
  jor  g11188(.dina(n11463), .dinb(n11460), .dout(n11464));
  jnot g11189(.din(n10970), .dout(n11465));
  jand g11190(.dina(n11462), .dinb(n11465), .dout(n11466));
  jnot g11191(.din(n11466), .dout(n11467));
  jand g11192(.dina(n11467), .dinb(n11464), .dout(n11468));
  jand g11193(.dina(n11468), .dinb(n11459), .dout(n11469));
  jor  g11194(.dina(n11469), .dinb(n11458), .dout(n11470));
  jand g11195(.dina(n11470), .dinb(asqrt[48] ), .dout(n11471));
  jor  g11196(.dina(n11458), .dinb(asqrt[48] ), .dout(n11472));
  jor  g11197(.dina(n11472), .dinb(n11469), .dout(n11473));
  jnot g11198(.din(n10976), .dout(n11474));
  jnot g11199(.din(n10978), .dout(n11475));
  jand g11200(.dina(asqrt[18] ), .dinb(n10972), .dout(n11476));
  jand g11201(.dina(n11476), .dinb(n11475), .dout(n11477));
  jor  g11202(.dina(n11477), .dinb(n11474), .dout(n11478));
  jnot g11203(.din(n10979), .dout(n11479));
  jand g11204(.dina(n11476), .dinb(n11479), .dout(n11480));
  jnot g11205(.din(n11480), .dout(n11481));
  jand g11206(.dina(n11481), .dinb(n11478), .dout(n11482));
  jand g11207(.dina(n11482), .dinb(n11473), .dout(n11483));
  jor  g11208(.dina(n11483), .dinb(n11471), .dout(n11484));
  jand g11209(.dina(n11484), .dinb(asqrt[49] ), .dout(n11485));
  jxor g11210(.dina(n10980), .dinb(n1641), .dout(n11486));
  jand g11211(.dina(n11486), .dinb(asqrt[18] ), .dout(n11487));
  jxor g11212(.dina(n11487), .dinb(n10990), .dout(n11488));
  jnot g11213(.din(n11488), .dout(n11489));
  jor  g11214(.dina(n11484), .dinb(asqrt[49] ), .dout(n11490));
  jand g11215(.dina(n11490), .dinb(n11489), .dout(n11491));
  jor  g11216(.dina(n11491), .dinb(n11485), .dout(n11492));
  jand g11217(.dina(n11492), .dinb(asqrt[50] ), .dout(n11493));
  jnot g11218(.din(n10995), .dout(n11494));
  jand g11219(.dina(n11494), .dinb(n10993), .dout(n11495));
  jand g11220(.dina(n11495), .dinb(asqrt[18] ), .dout(n11496));
  jxor g11221(.dina(n11496), .dinb(n11003), .dout(n11497));
  jnot g11222(.din(n11497), .dout(n11498));
  jor  g11223(.dina(n11485), .dinb(asqrt[50] ), .dout(n11499));
  jor  g11224(.dina(n11499), .dinb(n11491), .dout(n11500));
  jand g11225(.dina(n11500), .dinb(n11498), .dout(n11501));
  jor  g11226(.dina(n11501), .dinb(n11493), .dout(n11502));
  jand g11227(.dina(n11502), .dinb(asqrt[51] ), .dout(n11503));
  jor  g11228(.dina(n11502), .dinb(asqrt[51] ), .dout(n11504));
  jnot g11229(.din(n11009), .dout(n11505));
  jnot g11230(.din(n11010), .dout(n11506));
  jand g11231(.dina(asqrt[18] ), .dinb(n11006), .dout(n11507));
  jand g11232(.dina(n11507), .dinb(n11506), .dout(n11508));
  jor  g11233(.dina(n11508), .dinb(n11505), .dout(n11509));
  jnot g11234(.din(n11011), .dout(n11510));
  jand g11235(.dina(n11507), .dinb(n11510), .dout(n11511));
  jnot g11236(.din(n11511), .dout(n11512));
  jand g11237(.dina(n11512), .dinb(n11509), .dout(n11513));
  jand g11238(.dina(n11513), .dinb(n11504), .dout(n11514));
  jor  g11239(.dina(n11514), .dinb(n11503), .dout(n11515));
  jand g11240(.dina(n11515), .dinb(asqrt[52] ), .dout(n11516));
  jor  g11241(.dina(n11503), .dinb(asqrt[52] ), .dout(n11517));
  jor  g11242(.dina(n11517), .dinb(n11514), .dout(n11518));
  jnot g11243(.din(n11017), .dout(n11519));
  jnot g11244(.din(n11019), .dout(n11520));
  jand g11245(.dina(asqrt[18] ), .dinb(n11013), .dout(n11521));
  jand g11246(.dina(n11521), .dinb(n11520), .dout(n11522));
  jor  g11247(.dina(n11522), .dinb(n11519), .dout(n11523));
  jnot g11248(.din(n11020), .dout(n11524));
  jand g11249(.dina(n11521), .dinb(n11524), .dout(n11525));
  jnot g11250(.din(n11525), .dout(n11526));
  jand g11251(.dina(n11526), .dinb(n11523), .dout(n11527));
  jand g11252(.dina(n11527), .dinb(n11518), .dout(n11528));
  jor  g11253(.dina(n11528), .dinb(n11516), .dout(n11529));
  jand g11254(.dina(n11529), .dinb(asqrt[53] ), .dout(n11530));
  jxor g11255(.dina(n11021), .dinb(n1034), .dout(n11531));
  jand g11256(.dina(n11531), .dinb(asqrt[18] ), .dout(n11532));
  jxor g11257(.dina(n11532), .dinb(n11031), .dout(n11533));
  jnot g11258(.din(n11533), .dout(n11534));
  jor  g11259(.dina(n11529), .dinb(asqrt[53] ), .dout(n11535));
  jand g11260(.dina(n11535), .dinb(n11534), .dout(n11536));
  jor  g11261(.dina(n11536), .dinb(n11530), .dout(n11537));
  jand g11262(.dina(n11537), .dinb(asqrt[54] ), .dout(n11538));
  jnot g11263(.din(n11036), .dout(n11539));
  jand g11264(.dina(n11539), .dinb(n11034), .dout(n11540));
  jand g11265(.dina(n11540), .dinb(asqrt[18] ), .dout(n11541));
  jxor g11266(.dina(n11541), .dinb(n11044), .dout(n11542));
  jnot g11267(.din(n11542), .dout(n11543));
  jor  g11268(.dina(n11530), .dinb(asqrt[54] ), .dout(n11544));
  jor  g11269(.dina(n11544), .dinb(n11536), .dout(n11545));
  jand g11270(.dina(n11545), .dinb(n11543), .dout(n11546));
  jor  g11271(.dina(n11546), .dinb(n11538), .dout(n11547));
  jand g11272(.dina(n11547), .dinb(asqrt[55] ), .dout(n11548));
  jor  g11273(.dina(n11547), .dinb(asqrt[55] ), .dout(n11549));
  jnot g11274(.din(n11050), .dout(n11550));
  jnot g11275(.din(n11051), .dout(n11551));
  jand g11276(.dina(asqrt[18] ), .dinb(n11047), .dout(n11552));
  jand g11277(.dina(n11552), .dinb(n11551), .dout(n11553));
  jor  g11278(.dina(n11553), .dinb(n11550), .dout(n11554));
  jnot g11279(.din(n11052), .dout(n11555));
  jand g11280(.dina(n11552), .dinb(n11555), .dout(n11556));
  jnot g11281(.din(n11556), .dout(n11557));
  jand g11282(.dina(n11557), .dinb(n11554), .dout(n11558));
  jand g11283(.dina(n11558), .dinb(n11549), .dout(n11559));
  jor  g11284(.dina(n11559), .dinb(n11548), .dout(n11560));
  jand g11285(.dina(n11560), .dinb(asqrt[56] ), .dout(n11561));
  jor  g11286(.dina(n11548), .dinb(asqrt[56] ), .dout(n11562));
  jor  g11287(.dina(n11562), .dinb(n11559), .dout(n11563));
  jnot g11288(.din(n11058), .dout(n11564));
  jnot g11289(.din(n11060), .dout(n11565));
  jand g11290(.dina(asqrt[18] ), .dinb(n11054), .dout(n11566));
  jand g11291(.dina(n11566), .dinb(n11565), .dout(n11567));
  jor  g11292(.dina(n11567), .dinb(n11564), .dout(n11568));
  jnot g11293(.din(n11061), .dout(n11569));
  jand g11294(.dina(n11566), .dinb(n11569), .dout(n11570));
  jnot g11295(.din(n11570), .dout(n11571));
  jand g11296(.dina(n11571), .dinb(n11568), .dout(n11572));
  jand g11297(.dina(n11572), .dinb(n11563), .dout(n11573));
  jor  g11298(.dina(n11573), .dinb(n11561), .dout(n11574));
  jand g11299(.dina(n11574), .dinb(asqrt[57] ), .dout(n11575));
  jxor g11300(.dina(n11062), .dinb(n590), .dout(n11576));
  jand g11301(.dina(n11576), .dinb(asqrt[18] ), .dout(n11577));
  jxor g11302(.dina(n11577), .dinb(n11072), .dout(n11578));
  jnot g11303(.din(n11578), .dout(n11579));
  jor  g11304(.dina(n11574), .dinb(asqrt[57] ), .dout(n11580));
  jand g11305(.dina(n11580), .dinb(n11579), .dout(n11581));
  jor  g11306(.dina(n11581), .dinb(n11575), .dout(n11582));
  jand g11307(.dina(n11582), .dinb(asqrt[58] ), .dout(n11583));
  jnot g11308(.din(n11077), .dout(n11584));
  jand g11309(.dina(n11584), .dinb(n11075), .dout(n11585));
  jand g11310(.dina(n11585), .dinb(asqrt[18] ), .dout(n11586));
  jxor g11311(.dina(n11586), .dinb(n11085), .dout(n11587));
  jnot g11312(.din(n11587), .dout(n11588));
  jor  g11313(.dina(n11575), .dinb(asqrt[58] ), .dout(n11589));
  jor  g11314(.dina(n11589), .dinb(n11581), .dout(n11590));
  jand g11315(.dina(n11590), .dinb(n11588), .dout(n11591));
  jor  g11316(.dina(n11591), .dinb(n11583), .dout(n11592));
  jand g11317(.dina(n11592), .dinb(asqrt[59] ), .dout(n11593));
  jor  g11318(.dina(n11592), .dinb(asqrt[59] ), .dout(n11594));
  jnot g11319(.din(n11091), .dout(n11595));
  jnot g11320(.din(n11092), .dout(n11596));
  jand g11321(.dina(asqrt[18] ), .dinb(n11088), .dout(n11597));
  jand g11322(.dina(n11597), .dinb(n11596), .dout(n11598));
  jor  g11323(.dina(n11598), .dinb(n11595), .dout(n11599));
  jnot g11324(.din(n11093), .dout(n11600));
  jand g11325(.dina(n11597), .dinb(n11600), .dout(n11601));
  jnot g11326(.din(n11601), .dout(n11602));
  jand g11327(.dina(n11602), .dinb(n11599), .dout(n11603));
  jand g11328(.dina(n11603), .dinb(n11594), .dout(n11604));
  jor  g11329(.dina(n11604), .dinb(n11593), .dout(n11605));
  jand g11330(.dina(n11605), .dinb(asqrt[60] ), .dout(n11606));
  jor  g11331(.dina(n11593), .dinb(asqrt[60] ), .dout(n11607));
  jor  g11332(.dina(n11607), .dinb(n11604), .dout(n11608));
  jnot g11333(.din(n11099), .dout(n11609));
  jnot g11334(.din(n11101), .dout(n11610));
  jand g11335(.dina(asqrt[18] ), .dinb(n11095), .dout(n11611));
  jand g11336(.dina(n11611), .dinb(n11610), .dout(n11612));
  jor  g11337(.dina(n11612), .dinb(n11609), .dout(n11613));
  jnot g11338(.din(n11102), .dout(n11614));
  jand g11339(.dina(n11611), .dinb(n11614), .dout(n11615));
  jnot g11340(.din(n11615), .dout(n11616));
  jand g11341(.dina(n11616), .dinb(n11613), .dout(n11617));
  jand g11342(.dina(n11617), .dinb(n11608), .dout(n11618));
  jor  g11343(.dina(n11618), .dinb(n11606), .dout(n11619));
  jand g11344(.dina(n11619), .dinb(asqrt[61] ), .dout(n11620));
  jxor g11345(.dina(n11103), .dinb(n290), .dout(n11621));
  jand g11346(.dina(n11621), .dinb(asqrt[18] ), .dout(n11622));
  jxor g11347(.dina(n11622), .dinb(n11113), .dout(n11623));
  jnot g11348(.din(n11623), .dout(n11624));
  jor  g11349(.dina(n11619), .dinb(asqrt[61] ), .dout(n11625));
  jand g11350(.dina(n11625), .dinb(n11624), .dout(n11626));
  jor  g11351(.dina(n11626), .dinb(n11620), .dout(n11627));
  jand g11352(.dina(n11627), .dinb(asqrt[62] ), .dout(n11628));
  jnot g11353(.din(n11118), .dout(n11629));
  jand g11354(.dina(n11629), .dinb(n11116), .dout(n11630));
  jand g11355(.dina(n11630), .dinb(asqrt[18] ), .dout(n11631));
  jxor g11356(.dina(n11631), .dinb(n11126), .dout(n11632));
  jnot g11357(.din(n11632), .dout(n11633));
  jor  g11358(.dina(n11620), .dinb(asqrt[62] ), .dout(n11634));
  jor  g11359(.dina(n11634), .dinb(n11626), .dout(n11635));
  jand g11360(.dina(n11635), .dinb(n11633), .dout(n11636));
  jor  g11361(.dina(n11636), .dinb(n11628), .dout(n11637));
  jxor g11362(.dina(n11128), .dinb(n199), .dout(n11638));
  jand g11363(.dina(n11638), .dinb(asqrt[18] ), .dout(n11639));
  jxor g11364(.dina(n11639), .dinb(n11133), .dout(n11640));
  jnot g11365(.din(n11135), .dout(n11641));
  jnot g11366(.din(n11139), .dout(n11642));
  jand g11367(.dina(asqrt[18] ), .dinb(n11642), .dout(n11643));
  jand g11368(.dina(n11643), .dinb(n11641), .dout(n11644));
  jor  g11369(.dina(n11644), .dinb(n11146), .dout(n11645));
  jor  g11370(.dina(n11645), .dinb(n11640), .dout(n11646));
  jnot g11371(.din(n11646), .dout(n11647));
  jand g11372(.dina(n11647), .dinb(n11637), .dout(n11648));
  jor  g11373(.dina(n11648), .dinb(asqrt[63] ), .dout(n11649));
  jnot g11374(.din(n11640), .dout(n11650));
  jor  g11375(.dina(n11650), .dinb(n11637), .dout(n11651));
  jor  g11376(.dina(n11643), .dinb(n11641), .dout(n11652));
  jand g11377(.dina(n11642), .dinb(n11641), .dout(n11653));
  jor  g11378(.dina(n11653), .dinb(n194), .dout(n11654));
  jnot g11379(.din(n11654), .dout(n11655));
  jand g11380(.dina(n11655), .dinb(n11652), .dout(n11656));
  jnot g11381(.din(asqrt[18] ), .dout(n11657));
  jnot g11382(.din(n11656), .dout(n11660));
  jand g11383(.dina(n11660), .dinb(n11651), .dout(n11661));
  jand g11384(.dina(n11661), .dinb(n11649), .dout(n11662));
  jxor g11385(.dina(n11438), .dinb(n2010), .dout(n11663));
  jor  g11386(.dina(n11663), .dinb(n11662), .dout(n11664));
  jxor g11387(.dina(n11664), .dinb(n11158), .dout(n11665));
  jor  g11388(.dina(n11662), .dinb(n11160), .dout(n11666));
  jnot g11389(.din(a[32] ), .dout(n11667));
  jnot g11390(.din(a[33] ), .dout(n11668));
  jand g11391(.dina(n11160), .dinb(n11668), .dout(n11669));
  jand g11392(.dina(n11669), .dinb(n11667), .dout(n11670));
  jnot g11393(.din(n11670), .dout(n11671));
  jand g11394(.dina(n11671), .dinb(n11666), .dout(n11672));
  jor  g11395(.dina(n11672), .dinb(n11657), .dout(n11673));
  jor  g11396(.dina(n11662), .dinb(a[34] ), .dout(n11674));
  jxor g11397(.dina(n11674), .dinb(n11161), .dout(n11675));
  jand g11398(.dina(n11672), .dinb(n11657), .dout(n11676));
  jor  g11399(.dina(n11676), .dinb(n11675), .dout(n11677));
  jand g11400(.dina(n11677), .dinb(n11673), .dout(n11678));
  jor  g11401(.dina(n11678), .dinb(n10701), .dout(n11679));
  jand g11402(.dina(n11673), .dinb(n10701), .dout(n11680));
  jand g11403(.dina(n11680), .dinb(n11677), .dout(n11681));
  jor  g11404(.dina(n11674), .dinb(a[35] ), .dout(n11682));
  jnot g11405(.din(n11649), .dout(n11683));
  jnot g11406(.din(n11651), .dout(n11684));
  jor  g11407(.dina(n11656), .dinb(n11657), .dout(n11685));
  jor  g11408(.dina(n11685), .dinb(n11684), .dout(n11686));
  jor  g11409(.dina(n11686), .dinb(n11683), .dout(n11687));
  jand g11410(.dina(n11687), .dinb(n11682), .dout(n11688));
  jxor g11411(.dina(n11688), .dinb(n10706), .dout(n11689));
  jor  g11412(.dina(n11689), .dinb(n11681), .dout(n11690));
  jand g11413(.dina(n11690), .dinb(n11679), .dout(n11691));
  jor  g11414(.dina(n11691), .dinb(n10696), .dout(n11692));
  jand g11415(.dina(n11691), .dinb(n10696), .dout(n11693));
  jxor g11416(.dina(n11164), .dinb(n10701), .dout(n11694));
  jor  g11417(.dina(n11694), .dinb(n11662), .dout(n11695));
  jxor g11418(.dina(n11695), .dinb(n11167), .dout(n11696));
  jor  g11419(.dina(n11696), .dinb(n11693), .dout(n11697));
  jand g11420(.dina(n11697), .dinb(n11692), .dout(n11698));
  jor  g11421(.dina(n11698), .dinb(n9774), .dout(n11699));
  jnot g11422(.din(n11173), .dout(n11700));
  jor  g11423(.dina(n11700), .dinb(n11171), .dout(n11701));
  jor  g11424(.dina(n11701), .dinb(n11662), .dout(n11702));
  jxor g11425(.dina(n11702), .dinb(n11182), .dout(n11703));
  jand g11426(.dina(n11692), .dinb(n9774), .dout(n11704));
  jand g11427(.dina(n11704), .dinb(n11697), .dout(n11705));
  jor  g11428(.dina(n11705), .dinb(n11703), .dout(n11706));
  jand g11429(.dina(n11706), .dinb(n11699), .dout(n11707));
  jor  g11430(.dina(n11707), .dinb(n9769), .dout(n11708));
  jand g11431(.dina(n11707), .dinb(n9769), .dout(n11709));
  jxor g11432(.dina(n11184), .dinb(n9774), .dout(n11710));
  jor  g11433(.dina(n11710), .dinb(n11662), .dout(n11711));
  jxor g11434(.dina(n11711), .dinb(n11189), .dout(n11712));
  jnot g11435(.din(n11712), .dout(n11713));
  jor  g11436(.dina(n11713), .dinb(n11709), .dout(n11714));
  jand g11437(.dina(n11714), .dinb(n11708), .dout(n11715));
  jor  g11438(.dina(n11715), .dinb(n8898), .dout(n11716));
  jand g11439(.dina(n11708), .dinb(n8898), .dout(n11717));
  jand g11440(.dina(n11717), .dinb(n11714), .dout(n11718));
  jnot g11441(.din(n11193), .dout(n11719));
  jnot g11442(.din(n11662), .dout(asqrt[17] ));
  jand g11443(.dina(asqrt[17] ), .dinb(n11719), .dout(n11721));
  jand g11444(.dina(n11721), .dinb(n11200), .dout(n11722));
  jor  g11445(.dina(n11722), .dinb(n11198), .dout(n11723));
  jand g11446(.dina(n11721), .dinb(n11201), .dout(n11724));
  jnot g11447(.din(n11724), .dout(n11725));
  jand g11448(.dina(n11725), .dinb(n11723), .dout(n11726));
  jnot g11449(.din(n11726), .dout(n11727));
  jor  g11450(.dina(n11727), .dinb(n11718), .dout(n11728));
  jand g11451(.dina(n11728), .dinb(n11716), .dout(n11729));
  jor  g11452(.dina(n11729), .dinb(n8893), .dout(n11730));
  jand g11453(.dina(n11729), .dinb(n8893), .dout(n11731));
  jnot g11454(.din(n11208), .dout(n11732));
  jxor g11455(.dina(n11202), .dinb(n8898), .dout(n11733));
  jor  g11456(.dina(n11733), .dinb(n11662), .dout(n11734));
  jxor g11457(.dina(n11734), .dinb(n11732), .dout(n11735));
  jnot g11458(.din(n11735), .dout(n11736));
  jor  g11459(.dina(n11736), .dinb(n11731), .dout(n11737));
  jand g11460(.dina(n11737), .dinb(n11730), .dout(n11738));
  jor  g11461(.dina(n11738), .dinb(n8058), .dout(n11739));
  jnot g11462(.din(n11213), .dout(n11740));
  jor  g11463(.dina(n11740), .dinb(n11211), .dout(n11741));
  jor  g11464(.dina(n11741), .dinb(n11662), .dout(n11742));
  jxor g11465(.dina(n11742), .dinb(n11222), .dout(n11743));
  jand g11466(.dina(n11730), .dinb(n8058), .dout(n11744));
  jand g11467(.dina(n11744), .dinb(n11737), .dout(n11745));
  jor  g11468(.dina(n11745), .dinb(n11743), .dout(n11746));
  jand g11469(.dina(n11746), .dinb(n11739), .dout(n11747));
  jor  g11470(.dina(n11747), .dinb(n8053), .dout(n11748));
  jand g11471(.dina(n11747), .dinb(n8053), .dout(n11749));
  jnot g11472(.din(n11229), .dout(n11750));
  jxor g11473(.dina(n11224), .dinb(n8058), .dout(n11751));
  jor  g11474(.dina(n11751), .dinb(n11662), .dout(n11752));
  jxor g11475(.dina(n11752), .dinb(n11750), .dout(n11753));
  jnot g11476(.din(n11753), .dout(n11754));
  jor  g11477(.dina(n11754), .dinb(n11749), .dout(n11755));
  jand g11478(.dina(n11755), .dinb(n11748), .dout(n11756));
  jor  g11479(.dina(n11756), .dinb(n7265), .dout(n11757));
  jand g11480(.dina(n11748), .dinb(n7265), .dout(n11758));
  jand g11481(.dina(n11758), .dinb(n11755), .dout(n11759));
  jnot g11482(.din(n11232), .dout(n11760));
  jand g11483(.dina(asqrt[17] ), .dinb(n11760), .dout(n11761));
  jand g11484(.dina(n11761), .dinb(n11239), .dout(n11762));
  jor  g11485(.dina(n11762), .dinb(n11237), .dout(n11763));
  jand g11486(.dina(n11761), .dinb(n11240), .dout(n11764));
  jnot g11487(.din(n11764), .dout(n11765));
  jand g11488(.dina(n11765), .dinb(n11763), .dout(n11766));
  jnot g11489(.din(n11766), .dout(n11767));
  jor  g11490(.dina(n11767), .dinb(n11759), .dout(n11768));
  jand g11491(.dina(n11768), .dinb(n11757), .dout(n11769));
  jor  g11492(.dina(n11769), .dinb(n7260), .dout(n11770));
  jxor g11493(.dina(n11241), .dinb(n7265), .dout(n11771));
  jor  g11494(.dina(n11771), .dinb(n11662), .dout(n11772));
  jxor g11495(.dina(n11772), .dinb(n11246), .dout(n11773));
  jand g11496(.dina(n11769), .dinb(n7260), .dout(n11774));
  jor  g11497(.dina(n11774), .dinb(n11773), .dout(n11775));
  jand g11498(.dina(n11775), .dinb(n11770), .dout(n11776));
  jor  g11499(.dina(n11776), .dinb(n6505), .dout(n11777));
  jnot g11500(.din(n11251), .dout(n11778));
  jor  g11501(.dina(n11778), .dinb(n11249), .dout(n11779));
  jor  g11502(.dina(n11779), .dinb(n11662), .dout(n11780));
  jxor g11503(.dina(n11780), .dinb(n11260), .dout(n11781));
  jand g11504(.dina(n11770), .dinb(n6505), .dout(n11782));
  jand g11505(.dina(n11782), .dinb(n11775), .dout(n11783));
  jor  g11506(.dina(n11783), .dinb(n11781), .dout(n11784));
  jand g11507(.dina(n11784), .dinb(n11777), .dout(n11785));
  jor  g11508(.dina(n11785), .dinb(n6500), .dout(n11786));
  jand g11509(.dina(n11785), .dinb(n6500), .dout(n11787));
  jnot g11510(.din(n11263), .dout(n11788));
  jand g11511(.dina(asqrt[17] ), .dinb(n11788), .dout(n11789));
  jand g11512(.dina(n11789), .dinb(n11268), .dout(n11790));
  jor  g11513(.dina(n11790), .dinb(n11267), .dout(n11791));
  jand g11514(.dina(n11789), .dinb(n11269), .dout(n11792));
  jnot g11515(.din(n11792), .dout(n11793));
  jand g11516(.dina(n11793), .dinb(n11791), .dout(n11794));
  jnot g11517(.din(n11794), .dout(n11795));
  jor  g11518(.dina(n11795), .dinb(n11787), .dout(n11796));
  jand g11519(.dina(n11796), .dinb(n11786), .dout(n11797));
  jor  g11520(.dina(n11797), .dinb(n5793), .dout(n11798));
  jand g11521(.dina(n11786), .dinb(n5793), .dout(n11799));
  jand g11522(.dina(n11799), .dinb(n11796), .dout(n11800));
  jnot g11523(.din(n11271), .dout(n11801));
  jand g11524(.dina(asqrt[17] ), .dinb(n11801), .dout(n11802));
  jand g11525(.dina(n11802), .dinb(n11278), .dout(n11803));
  jor  g11526(.dina(n11803), .dinb(n11276), .dout(n11804));
  jand g11527(.dina(n11802), .dinb(n11279), .dout(n11805));
  jnot g11528(.din(n11805), .dout(n11806));
  jand g11529(.dina(n11806), .dinb(n11804), .dout(n11807));
  jnot g11530(.din(n11807), .dout(n11808));
  jor  g11531(.dina(n11808), .dinb(n11800), .dout(n11809));
  jand g11532(.dina(n11809), .dinb(n11798), .dout(n11810));
  jor  g11533(.dina(n11810), .dinb(n5788), .dout(n11811));
  jxor g11534(.dina(n11280), .dinb(n5793), .dout(n11812));
  jor  g11535(.dina(n11812), .dinb(n11662), .dout(n11813));
  jxor g11536(.dina(n11813), .dinb(n11291), .dout(n11814));
  jand g11537(.dina(n11810), .dinb(n5788), .dout(n11815));
  jor  g11538(.dina(n11815), .dinb(n11814), .dout(n11816));
  jand g11539(.dina(n11816), .dinb(n11811), .dout(n11817));
  jor  g11540(.dina(n11817), .dinb(n5121), .dout(n11818));
  jnot g11541(.din(n11296), .dout(n11819));
  jor  g11542(.dina(n11819), .dinb(n11294), .dout(n11820));
  jor  g11543(.dina(n11820), .dinb(n11662), .dout(n11821));
  jxor g11544(.dina(n11821), .dinb(n11305), .dout(n11822));
  jand g11545(.dina(n11811), .dinb(n5121), .dout(n11823));
  jand g11546(.dina(n11823), .dinb(n11816), .dout(n11824));
  jor  g11547(.dina(n11824), .dinb(n11822), .dout(n11825));
  jand g11548(.dina(n11825), .dinb(n11818), .dout(n11826));
  jor  g11549(.dina(n11826), .dinb(n5116), .dout(n11827));
  jand g11550(.dina(n11826), .dinb(n5116), .dout(n11828));
  jnot g11551(.din(n11308), .dout(n11829));
  jand g11552(.dina(asqrt[17] ), .dinb(n11829), .dout(n11830));
  jand g11553(.dina(n11830), .dinb(n11313), .dout(n11831));
  jor  g11554(.dina(n11831), .dinb(n11312), .dout(n11832));
  jand g11555(.dina(n11830), .dinb(n11314), .dout(n11833));
  jnot g11556(.din(n11833), .dout(n11834));
  jand g11557(.dina(n11834), .dinb(n11832), .dout(n11835));
  jnot g11558(.din(n11835), .dout(n11836));
  jor  g11559(.dina(n11836), .dinb(n11828), .dout(n11837));
  jand g11560(.dina(n11837), .dinb(n11827), .dout(n11838));
  jor  g11561(.dina(n11838), .dinb(n4499), .dout(n11839));
  jand g11562(.dina(n11827), .dinb(n4499), .dout(n11840));
  jand g11563(.dina(n11840), .dinb(n11837), .dout(n11841));
  jnot g11564(.din(n11316), .dout(n11842));
  jand g11565(.dina(asqrt[17] ), .dinb(n11842), .dout(n11843));
  jand g11566(.dina(n11843), .dinb(n11323), .dout(n11844));
  jor  g11567(.dina(n11844), .dinb(n11321), .dout(n11845));
  jand g11568(.dina(n11843), .dinb(n11324), .dout(n11846));
  jnot g11569(.din(n11846), .dout(n11847));
  jand g11570(.dina(n11847), .dinb(n11845), .dout(n11848));
  jnot g11571(.din(n11848), .dout(n11849));
  jor  g11572(.dina(n11849), .dinb(n11841), .dout(n11850));
  jand g11573(.dina(n11850), .dinb(n11839), .dout(n11851));
  jor  g11574(.dina(n11851), .dinb(n4494), .dout(n11852));
  jxor g11575(.dina(n11325), .dinb(n4499), .dout(n11853));
  jor  g11576(.dina(n11853), .dinb(n11662), .dout(n11854));
  jxor g11577(.dina(n11854), .dinb(n11336), .dout(n11855));
  jand g11578(.dina(n11851), .dinb(n4494), .dout(n11856));
  jor  g11579(.dina(n11856), .dinb(n11855), .dout(n11857));
  jand g11580(.dina(n11857), .dinb(n11852), .dout(n11858));
  jor  g11581(.dina(n11858), .dinb(n3912), .dout(n11859));
  jnot g11582(.din(n11341), .dout(n11860));
  jor  g11583(.dina(n11860), .dinb(n11339), .dout(n11861));
  jor  g11584(.dina(n11861), .dinb(n11662), .dout(n11862));
  jxor g11585(.dina(n11862), .dinb(n11350), .dout(n11863));
  jand g11586(.dina(n11852), .dinb(n3912), .dout(n11864));
  jand g11587(.dina(n11864), .dinb(n11857), .dout(n11865));
  jor  g11588(.dina(n11865), .dinb(n11863), .dout(n11866));
  jand g11589(.dina(n11866), .dinb(n11859), .dout(n11867));
  jor  g11590(.dina(n11867), .dinb(n3907), .dout(n11868));
  jand g11591(.dina(n11867), .dinb(n3907), .dout(n11869));
  jnot g11592(.din(n11353), .dout(n11870));
  jand g11593(.dina(asqrt[17] ), .dinb(n11870), .dout(n11871));
  jand g11594(.dina(n11871), .dinb(n11358), .dout(n11872));
  jor  g11595(.dina(n11872), .dinb(n11357), .dout(n11873));
  jand g11596(.dina(n11871), .dinb(n11359), .dout(n11874));
  jnot g11597(.din(n11874), .dout(n11875));
  jand g11598(.dina(n11875), .dinb(n11873), .dout(n11876));
  jnot g11599(.din(n11876), .dout(n11877));
  jor  g11600(.dina(n11877), .dinb(n11869), .dout(n11878));
  jand g11601(.dina(n11878), .dinb(n11868), .dout(n11879));
  jor  g11602(.dina(n11879), .dinb(n3376), .dout(n11880));
  jand g11603(.dina(n11868), .dinb(n3376), .dout(n11881));
  jand g11604(.dina(n11881), .dinb(n11878), .dout(n11882));
  jnot g11605(.din(n11361), .dout(n11883));
  jand g11606(.dina(asqrt[17] ), .dinb(n11883), .dout(n11884));
  jand g11607(.dina(n11884), .dinb(n11368), .dout(n11885));
  jor  g11608(.dina(n11885), .dinb(n11366), .dout(n11886));
  jand g11609(.dina(n11884), .dinb(n11369), .dout(n11887));
  jnot g11610(.din(n11887), .dout(n11888));
  jand g11611(.dina(n11888), .dinb(n11886), .dout(n11889));
  jnot g11612(.din(n11889), .dout(n11890));
  jor  g11613(.dina(n11890), .dinb(n11882), .dout(n11891));
  jand g11614(.dina(n11891), .dinb(n11880), .dout(n11892));
  jor  g11615(.dina(n11892), .dinb(n3371), .dout(n11893));
  jxor g11616(.dina(n11370), .dinb(n3376), .dout(n11894));
  jor  g11617(.dina(n11894), .dinb(n11662), .dout(n11895));
  jxor g11618(.dina(n11895), .dinb(n11381), .dout(n11896));
  jand g11619(.dina(n11892), .dinb(n3371), .dout(n11897));
  jor  g11620(.dina(n11897), .dinb(n11896), .dout(n11898));
  jand g11621(.dina(n11898), .dinb(n11893), .dout(n11899));
  jor  g11622(.dina(n11899), .dinb(n2875), .dout(n11900));
  jnot g11623(.din(n11386), .dout(n11901));
  jor  g11624(.dina(n11901), .dinb(n11384), .dout(n11902));
  jor  g11625(.dina(n11902), .dinb(n11662), .dout(n11903));
  jxor g11626(.dina(n11903), .dinb(n11395), .dout(n11904));
  jand g11627(.dina(n11893), .dinb(n2875), .dout(n11905));
  jand g11628(.dina(n11905), .dinb(n11898), .dout(n11906));
  jor  g11629(.dina(n11906), .dinb(n11904), .dout(n11907));
  jand g11630(.dina(n11907), .dinb(n11900), .dout(n11908));
  jor  g11631(.dina(n11908), .dinb(n2870), .dout(n11909));
  jand g11632(.dina(n11908), .dinb(n2870), .dout(n11910));
  jnot g11633(.din(n11398), .dout(n11911));
  jand g11634(.dina(asqrt[17] ), .dinb(n11911), .dout(n11912));
  jand g11635(.dina(n11912), .dinb(n11403), .dout(n11913));
  jor  g11636(.dina(n11913), .dinb(n11402), .dout(n11914));
  jand g11637(.dina(n11912), .dinb(n11404), .dout(n11915));
  jnot g11638(.din(n11915), .dout(n11916));
  jand g11639(.dina(n11916), .dinb(n11914), .dout(n11917));
  jnot g11640(.din(n11917), .dout(n11918));
  jor  g11641(.dina(n11918), .dinb(n11910), .dout(n11919));
  jand g11642(.dina(n11919), .dinb(n11909), .dout(n11920));
  jor  g11643(.dina(n11920), .dinb(n2425), .dout(n11921));
  jand g11644(.dina(n11909), .dinb(n2425), .dout(n11922));
  jand g11645(.dina(n11922), .dinb(n11919), .dout(n11923));
  jnot g11646(.din(n11406), .dout(n11924));
  jand g11647(.dina(asqrt[17] ), .dinb(n11924), .dout(n11925));
  jand g11648(.dina(n11925), .dinb(n11413), .dout(n11926));
  jor  g11649(.dina(n11926), .dinb(n11411), .dout(n11927));
  jand g11650(.dina(n11925), .dinb(n11414), .dout(n11928));
  jnot g11651(.din(n11928), .dout(n11929));
  jand g11652(.dina(n11929), .dinb(n11927), .dout(n11930));
  jnot g11653(.din(n11930), .dout(n11931));
  jor  g11654(.dina(n11931), .dinb(n11923), .dout(n11932));
  jand g11655(.dina(n11932), .dinb(n11921), .dout(n11933));
  jor  g11656(.dina(n11933), .dinb(n2420), .dout(n11934));
  jxor g11657(.dina(n11415), .dinb(n2425), .dout(n11935));
  jor  g11658(.dina(n11935), .dinb(n11662), .dout(n11936));
  jxor g11659(.dina(n11936), .dinb(n11426), .dout(n11937));
  jand g11660(.dina(n11933), .dinb(n2420), .dout(n11938));
  jor  g11661(.dina(n11938), .dinb(n11937), .dout(n11939));
  jand g11662(.dina(n11939), .dinb(n11934), .dout(n11940));
  jor  g11663(.dina(n11940), .dinb(n2010), .dout(n11941));
  jand g11664(.dina(n11934), .dinb(n2010), .dout(n11942));
  jand g11665(.dina(n11942), .dinb(n11939), .dout(n11943));
  jnot g11666(.din(n11429), .dout(n11944));
  jand g11667(.dina(asqrt[17] ), .dinb(n11944), .dout(n11945));
  jand g11668(.dina(n11945), .dinb(n11436), .dout(n11946));
  jor  g11669(.dina(n11946), .dinb(n11434), .dout(n11947));
  jand g11670(.dina(n11945), .dinb(n11437), .dout(n11948));
  jnot g11671(.din(n11948), .dout(n11949));
  jand g11672(.dina(n11949), .dinb(n11947), .dout(n11950));
  jnot g11673(.din(n11950), .dout(n11951));
  jor  g11674(.dina(n11951), .dinb(n11943), .dout(n11952));
  jand g11675(.dina(n11952), .dinb(n11941), .dout(n11953));
  jor  g11676(.dina(n11953), .dinb(n2005), .dout(n11954));
  jnot g11677(.din(n11665), .dout(n11955));
  jand g11678(.dina(n11953), .dinb(n2005), .dout(n11956));
  jor  g11679(.dina(n11956), .dinb(n11955), .dout(n11957));
  jand g11680(.dina(n11957), .dinb(n11954), .dout(n11958));
  jor  g11681(.dina(n11958), .dinb(n1646), .dout(n11959));
  jnot g11682(.din(n11446), .dout(n11960));
  jor  g11683(.dina(n11960), .dinb(n11444), .dout(n11961));
  jor  g11684(.dina(n11961), .dinb(n11662), .dout(n11962));
  jxor g11685(.dina(n11962), .dinb(n11455), .dout(n11963));
  jand g11686(.dina(n11954), .dinb(n1646), .dout(n11964));
  jand g11687(.dina(n11964), .dinb(n11957), .dout(n11965));
  jor  g11688(.dina(n11965), .dinb(n11963), .dout(n11966));
  jand g11689(.dina(n11966), .dinb(n11959), .dout(n11967));
  jor  g11690(.dina(n11967), .dinb(n1641), .dout(n11968));
  jxor g11691(.dina(n11457), .dinb(n1646), .dout(n11969));
  jor  g11692(.dina(n11969), .dinb(n11662), .dout(n11970));
  jxor g11693(.dina(n11970), .dinb(n11468), .dout(n11971));
  jand g11694(.dina(n11967), .dinb(n1641), .dout(n11972));
  jor  g11695(.dina(n11972), .dinb(n11971), .dout(n11973));
  jand g11696(.dina(n11973), .dinb(n11968), .dout(n11974));
  jor  g11697(.dina(n11974), .dinb(n1317), .dout(n11975));
  jnot g11698(.din(n11473), .dout(n11976));
  jor  g11699(.dina(n11976), .dinb(n11471), .dout(n11977));
  jor  g11700(.dina(n11977), .dinb(n11662), .dout(n11978));
  jxor g11701(.dina(n11978), .dinb(n11482), .dout(n11979));
  jand g11702(.dina(n11968), .dinb(n1317), .dout(n11980));
  jand g11703(.dina(n11980), .dinb(n11973), .dout(n11981));
  jor  g11704(.dina(n11981), .dinb(n11979), .dout(n11982));
  jand g11705(.dina(n11982), .dinb(n11975), .dout(n11983));
  jor  g11706(.dina(n11983), .dinb(n1312), .dout(n11984));
  jand g11707(.dina(n11983), .dinb(n1312), .dout(n11985));
  jnot g11708(.din(n11485), .dout(n11986));
  jand g11709(.dina(asqrt[17] ), .dinb(n11986), .dout(n11987));
  jand g11710(.dina(n11987), .dinb(n11490), .dout(n11988));
  jor  g11711(.dina(n11988), .dinb(n11489), .dout(n11989));
  jand g11712(.dina(n11987), .dinb(n11491), .dout(n11990));
  jnot g11713(.din(n11990), .dout(n11991));
  jand g11714(.dina(n11991), .dinb(n11989), .dout(n11992));
  jnot g11715(.din(n11992), .dout(n11993));
  jor  g11716(.dina(n11993), .dinb(n11985), .dout(n11994));
  jand g11717(.dina(n11994), .dinb(n11984), .dout(n11995));
  jor  g11718(.dina(n11995), .dinb(n1039), .dout(n11996));
  jand g11719(.dina(n11984), .dinb(n1039), .dout(n11997));
  jand g11720(.dina(n11997), .dinb(n11994), .dout(n11998));
  jnot g11721(.din(n11493), .dout(n11999));
  jand g11722(.dina(asqrt[17] ), .dinb(n11999), .dout(n12000));
  jand g11723(.dina(n12000), .dinb(n11500), .dout(n12001));
  jor  g11724(.dina(n12001), .dinb(n11498), .dout(n12002));
  jand g11725(.dina(n12000), .dinb(n11501), .dout(n12003));
  jnot g11726(.din(n12003), .dout(n12004));
  jand g11727(.dina(n12004), .dinb(n12002), .dout(n12005));
  jnot g11728(.din(n12005), .dout(n12006));
  jor  g11729(.dina(n12006), .dinb(n11998), .dout(n12007));
  jand g11730(.dina(n12007), .dinb(n11996), .dout(n12008));
  jor  g11731(.dina(n12008), .dinb(n1034), .dout(n12009));
  jxor g11732(.dina(n11502), .dinb(n1039), .dout(n12010));
  jor  g11733(.dina(n12010), .dinb(n11662), .dout(n12011));
  jxor g11734(.dina(n12011), .dinb(n11513), .dout(n12012));
  jand g11735(.dina(n12008), .dinb(n1034), .dout(n12013));
  jor  g11736(.dina(n12013), .dinb(n12012), .dout(n12014));
  jand g11737(.dina(n12014), .dinb(n12009), .dout(n12015));
  jor  g11738(.dina(n12015), .dinb(n796), .dout(n12016));
  jnot g11739(.din(n11518), .dout(n12017));
  jor  g11740(.dina(n12017), .dinb(n11516), .dout(n12018));
  jor  g11741(.dina(n12018), .dinb(n11662), .dout(n12019));
  jxor g11742(.dina(n12019), .dinb(n11527), .dout(n12020));
  jand g11743(.dina(n12009), .dinb(n796), .dout(n12021));
  jand g11744(.dina(n12021), .dinb(n12014), .dout(n12022));
  jor  g11745(.dina(n12022), .dinb(n12020), .dout(n12023));
  jand g11746(.dina(n12023), .dinb(n12016), .dout(n12024));
  jor  g11747(.dina(n12024), .dinb(n791), .dout(n12025));
  jand g11748(.dina(n12024), .dinb(n791), .dout(n12026));
  jnot g11749(.din(n11530), .dout(n12027));
  jand g11750(.dina(asqrt[17] ), .dinb(n12027), .dout(n12028));
  jand g11751(.dina(n12028), .dinb(n11535), .dout(n12029));
  jor  g11752(.dina(n12029), .dinb(n11534), .dout(n12030));
  jand g11753(.dina(n12028), .dinb(n11536), .dout(n12031));
  jnot g11754(.din(n12031), .dout(n12032));
  jand g11755(.dina(n12032), .dinb(n12030), .dout(n12033));
  jnot g11756(.din(n12033), .dout(n12034));
  jor  g11757(.dina(n12034), .dinb(n12026), .dout(n12035));
  jand g11758(.dina(n12035), .dinb(n12025), .dout(n12036));
  jor  g11759(.dina(n12036), .dinb(n595), .dout(n12037));
  jand g11760(.dina(n12025), .dinb(n595), .dout(n12038));
  jand g11761(.dina(n12038), .dinb(n12035), .dout(n12039));
  jnot g11762(.din(n11538), .dout(n12040));
  jand g11763(.dina(asqrt[17] ), .dinb(n12040), .dout(n12041));
  jand g11764(.dina(n12041), .dinb(n11545), .dout(n12042));
  jor  g11765(.dina(n12042), .dinb(n11543), .dout(n12043));
  jand g11766(.dina(n12041), .dinb(n11546), .dout(n12044));
  jnot g11767(.din(n12044), .dout(n12045));
  jand g11768(.dina(n12045), .dinb(n12043), .dout(n12046));
  jnot g11769(.din(n12046), .dout(n12047));
  jor  g11770(.dina(n12047), .dinb(n12039), .dout(n12048));
  jand g11771(.dina(n12048), .dinb(n12037), .dout(n12049));
  jor  g11772(.dina(n12049), .dinb(n590), .dout(n12050));
  jxor g11773(.dina(n11547), .dinb(n595), .dout(n12051));
  jor  g11774(.dina(n12051), .dinb(n11662), .dout(n12052));
  jxor g11775(.dina(n12052), .dinb(n11558), .dout(n12053));
  jand g11776(.dina(n12049), .dinb(n590), .dout(n12054));
  jor  g11777(.dina(n12054), .dinb(n12053), .dout(n12055));
  jand g11778(.dina(n12055), .dinb(n12050), .dout(n12056));
  jor  g11779(.dina(n12056), .dinb(n430), .dout(n12057));
  jnot g11780(.din(n11563), .dout(n12058));
  jor  g11781(.dina(n12058), .dinb(n11561), .dout(n12059));
  jor  g11782(.dina(n12059), .dinb(n11662), .dout(n12060));
  jxor g11783(.dina(n12060), .dinb(n11572), .dout(n12061));
  jand g11784(.dina(n12050), .dinb(n430), .dout(n12062));
  jand g11785(.dina(n12062), .dinb(n12055), .dout(n12063));
  jor  g11786(.dina(n12063), .dinb(n12061), .dout(n12064));
  jand g11787(.dina(n12064), .dinb(n12057), .dout(n12065));
  jor  g11788(.dina(n12065), .dinb(n425), .dout(n12066));
  jand g11789(.dina(n12065), .dinb(n425), .dout(n12067));
  jnot g11790(.din(n11575), .dout(n12068));
  jand g11791(.dina(asqrt[17] ), .dinb(n12068), .dout(n12069));
  jand g11792(.dina(n12069), .dinb(n11580), .dout(n12070));
  jor  g11793(.dina(n12070), .dinb(n11579), .dout(n12071));
  jand g11794(.dina(n12069), .dinb(n11581), .dout(n12072));
  jnot g11795(.din(n12072), .dout(n12073));
  jand g11796(.dina(n12073), .dinb(n12071), .dout(n12074));
  jnot g11797(.din(n12074), .dout(n12075));
  jor  g11798(.dina(n12075), .dinb(n12067), .dout(n12076));
  jand g11799(.dina(n12076), .dinb(n12066), .dout(n12077));
  jor  g11800(.dina(n12077), .dinb(n305), .dout(n12078));
  jand g11801(.dina(n12066), .dinb(n305), .dout(n12079));
  jand g11802(.dina(n12079), .dinb(n12076), .dout(n12080));
  jnot g11803(.din(n11583), .dout(n12081));
  jand g11804(.dina(asqrt[17] ), .dinb(n12081), .dout(n12082));
  jand g11805(.dina(n12082), .dinb(n11590), .dout(n12083));
  jor  g11806(.dina(n12083), .dinb(n11588), .dout(n12084));
  jand g11807(.dina(n12082), .dinb(n11591), .dout(n12085));
  jnot g11808(.din(n12085), .dout(n12086));
  jand g11809(.dina(n12086), .dinb(n12084), .dout(n12087));
  jnot g11810(.din(n12087), .dout(n12088));
  jor  g11811(.dina(n12088), .dinb(n12080), .dout(n12089));
  jand g11812(.dina(n12089), .dinb(n12078), .dout(n12090));
  jor  g11813(.dina(n12090), .dinb(n290), .dout(n12091));
  jxor g11814(.dina(n11592), .dinb(n305), .dout(n12092));
  jor  g11815(.dina(n12092), .dinb(n11662), .dout(n12093));
  jxor g11816(.dina(n12093), .dinb(n11603), .dout(n12094));
  jand g11817(.dina(n12090), .dinb(n290), .dout(n12095));
  jor  g11818(.dina(n12095), .dinb(n12094), .dout(n12096));
  jand g11819(.dina(n12096), .dinb(n12091), .dout(n12097));
  jor  g11820(.dina(n12097), .dinb(n223), .dout(n12098));
  jnot g11821(.din(n11608), .dout(n12099));
  jor  g11822(.dina(n12099), .dinb(n11606), .dout(n12100));
  jor  g11823(.dina(n12100), .dinb(n11662), .dout(n12101));
  jxor g11824(.dina(n12101), .dinb(n11617), .dout(n12102));
  jand g11825(.dina(n12091), .dinb(n223), .dout(n12103));
  jand g11826(.dina(n12103), .dinb(n12096), .dout(n12104));
  jor  g11827(.dina(n12104), .dinb(n12102), .dout(n12105));
  jand g11828(.dina(n12105), .dinb(n12098), .dout(n12106));
  jor  g11829(.dina(n12106), .dinb(n199), .dout(n12107));
  jand g11830(.dina(n12106), .dinb(n199), .dout(n12108));
  jnot g11831(.din(n11620), .dout(n12109));
  jand g11832(.dina(asqrt[17] ), .dinb(n12109), .dout(n12110));
  jand g11833(.dina(n12110), .dinb(n11625), .dout(n12111));
  jor  g11834(.dina(n12111), .dinb(n11624), .dout(n12112));
  jand g11835(.dina(n12110), .dinb(n11626), .dout(n12113));
  jnot g11836(.din(n12113), .dout(n12114));
  jand g11837(.dina(n12114), .dinb(n12112), .dout(n12115));
  jnot g11838(.din(n12115), .dout(n12116));
  jor  g11839(.dina(n12116), .dinb(n12108), .dout(n12117));
  jand g11840(.dina(n12117), .dinb(n12107), .dout(n12118));
  jnot g11841(.din(n11628), .dout(n12119));
  jand g11842(.dina(asqrt[17] ), .dinb(n12119), .dout(n12120));
  jand g11843(.dina(n12120), .dinb(n11635), .dout(n12121));
  jor  g11844(.dina(n12121), .dinb(n11633), .dout(n12122));
  jand g11845(.dina(n12120), .dinb(n11636), .dout(n12123));
  jnot g11846(.din(n12123), .dout(n12124));
  jand g11847(.dina(n12124), .dinb(n12122), .dout(n12125));
  jnot g11848(.din(n12125), .dout(n12126));
  jand g11849(.dina(asqrt[17] ), .dinb(n11650), .dout(n12127));
  jand g11850(.dina(n12127), .dinb(n11637), .dout(n12128));
  jor  g11851(.dina(n12128), .dinb(n11684), .dout(n12129));
  jor  g11852(.dina(n12129), .dinb(n12126), .dout(n12130));
  jor  g11853(.dina(n12130), .dinb(n12118), .dout(n12131));
  jand g11854(.dina(n12131), .dinb(n194), .dout(n12132));
  jand g11855(.dina(n12126), .dinb(n12118), .dout(n12133));
  jor  g11856(.dina(n12127), .dinb(n11637), .dout(n12134));
  jand g11857(.dina(n11650), .dinb(n11637), .dout(n12135));
  jor  g11858(.dina(n12135), .dinb(n194), .dout(n12136));
  jnot g11859(.din(n12136), .dout(n12137));
  jand g11860(.dina(n12137), .dinb(n12134), .dout(n12138));
  jor  g11861(.dina(n12138), .dinb(n12133), .dout(n12141));
  jor  g11862(.dina(n12141), .dinb(n12132), .dout(asqrt[16] ));
  jxor g11863(.dina(n11953), .dinb(n2005), .dout(n12143));
  jand g11864(.dina(n12143), .dinb(asqrt[16] ), .dout(n12144));
  jxor g11865(.dina(n12144), .dinb(n11665), .dout(n12145));
  jnot g11866(.din(n12145), .dout(n12146));
  jand g11867(.dina(asqrt[16] ), .dinb(a[32] ), .dout(n12147));
  jnot g11868(.din(a[30] ), .dout(n12148));
  jnot g11869(.din(a[31] ), .dout(n12149));
  jand g11870(.dina(n11667), .dinb(n12149), .dout(n12150));
  jand g11871(.dina(n12150), .dinb(n12148), .dout(n12151));
  jor  g11872(.dina(n12151), .dinb(n12147), .dout(n12152));
  jand g11873(.dina(n12152), .dinb(asqrt[17] ), .dout(n12153));
  jand g11874(.dina(asqrt[16] ), .dinb(n11667), .dout(n12154));
  jxor g11875(.dina(n12154), .dinb(n11668), .dout(n12155));
  jor  g11876(.dina(n12152), .dinb(asqrt[17] ), .dout(n12156));
  jand g11877(.dina(n12156), .dinb(n12155), .dout(n12157));
  jor  g11878(.dina(n12157), .dinb(n12153), .dout(n12158));
  jand g11879(.dina(n12158), .dinb(asqrt[18] ), .dout(n12159));
  jor  g11880(.dina(n12153), .dinb(asqrt[18] ), .dout(n12160));
  jor  g11881(.dina(n12160), .dinb(n12157), .dout(n12161));
  jand g11882(.dina(n12154), .dinb(n11668), .dout(n12162));
  jnot g11883(.din(n12132), .dout(n12163));
  jnot g11884(.din(n12133), .dout(n12164));
  jnot g11885(.din(n12138), .dout(n12165));
  jand g11886(.dina(n12165), .dinb(asqrt[17] ), .dout(n12166));
  jand g11887(.dina(n12166), .dinb(n12164), .dout(n12167));
  jand g11888(.dina(n12167), .dinb(n12163), .dout(n12168));
  jor  g11889(.dina(n12168), .dinb(n12162), .dout(n12169));
  jxor g11890(.dina(n12169), .dinb(n11160), .dout(n12170));
  jand g11891(.dina(n12170), .dinb(n12161), .dout(n12171));
  jor  g11892(.dina(n12171), .dinb(n12159), .dout(n12172));
  jand g11893(.dina(n12172), .dinb(asqrt[19] ), .dout(n12173));
  jor  g11894(.dina(n12172), .dinb(asqrt[19] ), .dout(n12174));
  jxor g11895(.dina(n11672), .dinb(n11657), .dout(n12175));
  jand g11896(.dina(n12175), .dinb(asqrt[16] ), .dout(n12176));
  jxor g11897(.dina(n12176), .dinb(n11675), .dout(n12177));
  jnot g11898(.din(n12177), .dout(n12178));
  jand g11899(.dina(n12178), .dinb(n12174), .dout(n12179));
  jor  g11900(.dina(n12179), .dinb(n12173), .dout(n12180));
  jand g11901(.dina(n12180), .dinb(asqrt[20] ), .dout(n12181));
  jnot g11902(.din(n11681), .dout(n12182));
  jand g11903(.dina(n12182), .dinb(n11679), .dout(n12183));
  jand g11904(.dina(n12183), .dinb(asqrt[16] ), .dout(n12184));
  jxor g11905(.dina(n12184), .dinb(n11689), .dout(n12185));
  jnot g11906(.din(n12185), .dout(n12186));
  jor  g11907(.dina(n12173), .dinb(asqrt[20] ), .dout(n12187));
  jor  g11908(.dina(n12187), .dinb(n12179), .dout(n12188));
  jand g11909(.dina(n12188), .dinb(n12186), .dout(n12189));
  jor  g11910(.dina(n12189), .dinb(n12181), .dout(n12190));
  jand g11911(.dina(n12190), .dinb(asqrt[21] ), .dout(n12191));
  jor  g11912(.dina(n12190), .dinb(asqrt[21] ), .dout(n12192));
  jnot g11913(.din(n11696), .dout(n12193));
  jxor g11914(.dina(n11691), .dinb(n10696), .dout(n12194));
  jand g11915(.dina(n12194), .dinb(asqrt[16] ), .dout(n12195));
  jxor g11916(.dina(n12195), .dinb(n12193), .dout(n12196));
  jand g11917(.dina(n12196), .dinb(n12192), .dout(n12197));
  jor  g11918(.dina(n12197), .dinb(n12191), .dout(n12198));
  jand g11919(.dina(n12198), .dinb(asqrt[22] ), .dout(n12199));
  jor  g11920(.dina(n12191), .dinb(asqrt[22] ), .dout(n12200));
  jor  g11921(.dina(n12200), .dinb(n12197), .dout(n12201));
  jnot g11922(.din(n11703), .dout(n12202));
  jnot g11923(.din(n11705), .dout(n12203));
  jand g11924(.dina(asqrt[16] ), .dinb(n11699), .dout(n12204));
  jand g11925(.dina(n12204), .dinb(n12203), .dout(n12205));
  jor  g11926(.dina(n12205), .dinb(n12202), .dout(n12206));
  jnot g11927(.din(n11706), .dout(n12207));
  jand g11928(.dina(n12204), .dinb(n12207), .dout(n12208));
  jnot g11929(.din(n12208), .dout(n12209));
  jand g11930(.dina(n12209), .dinb(n12206), .dout(n12210));
  jand g11931(.dina(n12210), .dinb(n12201), .dout(n12211));
  jor  g11932(.dina(n12211), .dinb(n12199), .dout(n12212));
  jand g11933(.dina(n12212), .dinb(asqrt[23] ), .dout(n12213));
  jor  g11934(.dina(n12212), .dinb(asqrt[23] ), .dout(n12214));
  jxor g11935(.dina(n11707), .dinb(n9769), .dout(n12215));
  jand g11936(.dina(n12215), .dinb(asqrt[16] ), .dout(n12216));
  jxor g11937(.dina(n12216), .dinb(n11712), .dout(n12217));
  jand g11938(.dina(n12217), .dinb(n12214), .dout(n12218));
  jor  g11939(.dina(n12218), .dinb(n12213), .dout(n12219));
  jand g11940(.dina(n12219), .dinb(asqrt[24] ), .dout(n12220));
  jnot g11941(.din(n11718), .dout(n12221));
  jand g11942(.dina(n12221), .dinb(n11716), .dout(n12222));
  jand g11943(.dina(n12222), .dinb(asqrt[16] ), .dout(n12223));
  jxor g11944(.dina(n12223), .dinb(n11727), .dout(n12224));
  jnot g11945(.din(n12224), .dout(n12225));
  jor  g11946(.dina(n12213), .dinb(asqrt[24] ), .dout(n12226));
  jor  g11947(.dina(n12226), .dinb(n12218), .dout(n12227));
  jand g11948(.dina(n12227), .dinb(n12225), .dout(n12228));
  jor  g11949(.dina(n12228), .dinb(n12220), .dout(n12229));
  jand g11950(.dina(n12229), .dinb(asqrt[25] ), .dout(n12230));
  jor  g11951(.dina(n12229), .dinb(asqrt[25] ), .dout(n12231));
  jxor g11952(.dina(n11729), .dinb(n8893), .dout(n12232));
  jand g11953(.dina(n12232), .dinb(asqrt[16] ), .dout(n12233));
  jxor g11954(.dina(n12233), .dinb(n11735), .dout(n12234));
  jand g11955(.dina(n12234), .dinb(n12231), .dout(n12235));
  jor  g11956(.dina(n12235), .dinb(n12230), .dout(n12236));
  jand g11957(.dina(n12236), .dinb(asqrt[26] ), .dout(n12237));
  jor  g11958(.dina(n12230), .dinb(asqrt[26] ), .dout(n12238));
  jor  g11959(.dina(n12238), .dinb(n12235), .dout(n12239));
  jnot g11960(.din(n11743), .dout(n12240));
  jnot g11961(.din(n11745), .dout(n12241));
  jand g11962(.dina(asqrt[16] ), .dinb(n11739), .dout(n12242));
  jand g11963(.dina(n12242), .dinb(n12241), .dout(n12243));
  jor  g11964(.dina(n12243), .dinb(n12240), .dout(n12244));
  jnot g11965(.din(n11746), .dout(n12245));
  jand g11966(.dina(n12242), .dinb(n12245), .dout(n12246));
  jnot g11967(.din(n12246), .dout(n12247));
  jand g11968(.dina(n12247), .dinb(n12244), .dout(n12248));
  jand g11969(.dina(n12248), .dinb(n12239), .dout(n12249));
  jor  g11970(.dina(n12249), .dinb(n12237), .dout(n12250));
  jand g11971(.dina(n12250), .dinb(asqrt[27] ), .dout(n12251));
  jxor g11972(.dina(n11747), .dinb(n8053), .dout(n12252));
  jand g11973(.dina(n12252), .dinb(asqrt[16] ), .dout(n12253));
  jxor g11974(.dina(n12253), .dinb(n11754), .dout(n12254));
  jnot g11975(.din(n12254), .dout(n12255));
  jor  g11976(.dina(n12250), .dinb(asqrt[27] ), .dout(n12256));
  jand g11977(.dina(n12256), .dinb(n12255), .dout(n12257));
  jor  g11978(.dina(n12257), .dinb(n12251), .dout(n12258));
  jand g11979(.dina(n12258), .dinb(asqrt[28] ), .dout(n12259));
  jnot g11980(.din(n11759), .dout(n12260));
  jand g11981(.dina(n12260), .dinb(n11757), .dout(n12261));
  jand g11982(.dina(n12261), .dinb(asqrt[16] ), .dout(n12262));
  jxor g11983(.dina(n12262), .dinb(n11767), .dout(n12263));
  jnot g11984(.din(n12263), .dout(n12264));
  jor  g11985(.dina(n12251), .dinb(asqrt[28] ), .dout(n12265));
  jor  g11986(.dina(n12265), .dinb(n12257), .dout(n12266));
  jand g11987(.dina(n12266), .dinb(n12264), .dout(n12267));
  jor  g11988(.dina(n12267), .dinb(n12259), .dout(n12268));
  jand g11989(.dina(n12268), .dinb(asqrt[29] ), .dout(n12269));
  jor  g11990(.dina(n12268), .dinb(asqrt[29] ), .dout(n12270));
  jnot g11991(.din(n11773), .dout(n12271));
  jnot g11992(.din(n11774), .dout(n12272));
  jand g11993(.dina(asqrt[16] ), .dinb(n11770), .dout(n12273));
  jand g11994(.dina(n12273), .dinb(n12272), .dout(n12274));
  jor  g11995(.dina(n12274), .dinb(n12271), .dout(n12275));
  jnot g11996(.din(n11775), .dout(n12276));
  jand g11997(.dina(n12273), .dinb(n12276), .dout(n12277));
  jnot g11998(.din(n12277), .dout(n12278));
  jand g11999(.dina(n12278), .dinb(n12275), .dout(n12279));
  jand g12000(.dina(n12279), .dinb(n12270), .dout(n12280));
  jor  g12001(.dina(n12280), .dinb(n12269), .dout(n12281));
  jand g12002(.dina(n12281), .dinb(asqrt[30] ), .dout(n12282));
  jor  g12003(.dina(n12269), .dinb(asqrt[30] ), .dout(n12283));
  jor  g12004(.dina(n12283), .dinb(n12280), .dout(n12284));
  jnot g12005(.din(n11781), .dout(n12285));
  jnot g12006(.din(n11783), .dout(n12286));
  jand g12007(.dina(asqrt[16] ), .dinb(n11777), .dout(n12287));
  jand g12008(.dina(n12287), .dinb(n12286), .dout(n12288));
  jor  g12009(.dina(n12288), .dinb(n12285), .dout(n12289));
  jnot g12010(.din(n11784), .dout(n12290));
  jand g12011(.dina(n12287), .dinb(n12290), .dout(n12291));
  jnot g12012(.din(n12291), .dout(n12292));
  jand g12013(.dina(n12292), .dinb(n12289), .dout(n12293));
  jand g12014(.dina(n12293), .dinb(n12284), .dout(n12294));
  jor  g12015(.dina(n12294), .dinb(n12282), .dout(n12295));
  jand g12016(.dina(n12295), .dinb(asqrt[31] ), .dout(n12296));
  jxor g12017(.dina(n11785), .dinb(n6500), .dout(n12297));
  jand g12018(.dina(n12297), .dinb(asqrt[16] ), .dout(n12298));
  jxor g12019(.dina(n12298), .dinb(n11795), .dout(n12299));
  jnot g12020(.din(n12299), .dout(n12300));
  jor  g12021(.dina(n12295), .dinb(asqrt[31] ), .dout(n12301));
  jand g12022(.dina(n12301), .dinb(n12300), .dout(n12302));
  jor  g12023(.dina(n12302), .dinb(n12296), .dout(n12303));
  jand g12024(.dina(n12303), .dinb(asqrt[32] ), .dout(n12304));
  jnot g12025(.din(n11800), .dout(n12305));
  jand g12026(.dina(n12305), .dinb(n11798), .dout(n12306));
  jand g12027(.dina(n12306), .dinb(asqrt[16] ), .dout(n12307));
  jxor g12028(.dina(n12307), .dinb(n11808), .dout(n12308));
  jnot g12029(.din(n12308), .dout(n12309));
  jor  g12030(.dina(n12296), .dinb(asqrt[32] ), .dout(n12310));
  jor  g12031(.dina(n12310), .dinb(n12302), .dout(n12311));
  jand g12032(.dina(n12311), .dinb(n12309), .dout(n12312));
  jor  g12033(.dina(n12312), .dinb(n12304), .dout(n12313));
  jand g12034(.dina(n12313), .dinb(asqrt[33] ), .dout(n12314));
  jor  g12035(.dina(n12313), .dinb(asqrt[33] ), .dout(n12315));
  jnot g12036(.din(n11814), .dout(n12316));
  jnot g12037(.din(n11815), .dout(n12317));
  jand g12038(.dina(asqrt[16] ), .dinb(n11811), .dout(n12318));
  jand g12039(.dina(n12318), .dinb(n12317), .dout(n12319));
  jor  g12040(.dina(n12319), .dinb(n12316), .dout(n12320));
  jnot g12041(.din(n11816), .dout(n12321));
  jand g12042(.dina(n12318), .dinb(n12321), .dout(n12322));
  jnot g12043(.din(n12322), .dout(n12323));
  jand g12044(.dina(n12323), .dinb(n12320), .dout(n12324));
  jand g12045(.dina(n12324), .dinb(n12315), .dout(n12325));
  jor  g12046(.dina(n12325), .dinb(n12314), .dout(n12326));
  jand g12047(.dina(n12326), .dinb(asqrt[34] ), .dout(n12327));
  jor  g12048(.dina(n12314), .dinb(asqrt[34] ), .dout(n12328));
  jor  g12049(.dina(n12328), .dinb(n12325), .dout(n12329));
  jnot g12050(.din(n11822), .dout(n12330));
  jnot g12051(.din(n11824), .dout(n12331));
  jand g12052(.dina(asqrt[16] ), .dinb(n11818), .dout(n12332));
  jand g12053(.dina(n12332), .dinb(n12331), .dout(n12333));
  jor  g12054(.dina(n12333), .dinb(n12330), .dout(n12334));
  jnot g12055(.din(n11825), .dout(n12335));
  jand g12056(.dina(n12332), .dinb(n12335), .dout(n12336));
  jnot g12057(.din(n12336), .dout(n12337));
  jand g12058(.dina(n12337), .dinb(n12334), .dout(n12338));
  jand g12059(.dina(n12338), .dinb(n12329), .dout(n12339));
  jor  g12060(.dina(n12339), .dinb(n12327), .dout(n12340));
  jand g12061(.dina(n12340), .dinb(asqrt[35] ), .dout(n12341));
  jxor g12062(.dina(n11826), .dinb(n5116), .dout(n12342));
  jand g12063(.dina(n12342), .dinb(asqrt[16] ), .dout(n12343));
  jxor g12064(.dina(n12343), .dinb(n11836), .dout(n12344));
  jnot g12065(.din(n12344), .dout(n12345));
  jor  g12066(.dina(n12340), .dinb(asqrt[35] ), .dout(n12346));
  jand g12067(.dina(n12346), .dinb(n12345), .dout(n12347));
  jor  g12068(.dina(n12347), .dinb(n12341), .dout(n12348));
  jand g12069(.dina(n12348), .dinb(asqrt[36] ), .dout(n12349));
  jnot g12070(.din(n11841), .dout(n12350));
  jand g12071(.dina(n12350), .dinb(n11839), .dout(n12351));
  jand g12072(.dina(n12351), .dinb(asqrt[16] ), .dout(n12352));
  jxor g12073(.dina(n12352), .dinb(n11849), .dout(n12353));
  jnot g12074(.din(n12353), .dout(n12354));
  jor  g12075(.dina(n12341), .dinb(asqrt[36] ), .dout(n12355));
  jor  g12076(.dina(n12355), .dinb(n12347), .dout(n12356));
  jand g12077(.dina(n12356), .dinb(n12354), .dout(n12357));
  jor  g12078(.dina(n12357), .dinb(n12349), .dout(n12358));
  jand g12079(.dina(n12358), .dinb(asqrt[37] ), .dout(n12359));
  jor  g12080(.dina(n12358), .dinb(asqrt[37] ), .dout(n12360));
  jnot g12081(.din(n11855), .dout(n12361));
  jnot g12082(.din(n11856), .dout(n12362));
  jand g12083(.dina(asqrt[16] ), .dinb(n11852), .dout(n12363));
  jand g12084(.dina(n12363), .dinb(n12362), .dout(n12364));
  jor  g12085(.dina(n12364), .dinb(n12361), .dout(n12365));
  jnot g12086(.din(n11857), .dout(n12366));
  jand g12087(.dina(n12363), .dinb(n12366), .dout(n12367));
  jnot g12088(.din(n12367), .dout(n12368));
  jand g12089(.dina(n12368), .dinb(n12365), .dout(n12369));
  jand g12090(.dina(n12369), .dinb(n12360), .dout(n12370));
  jor  g12091(.dina(n12370), .dinb(n12359), .dout(n12371));
  jand g12092(.dina(n12371), .dinb(asqrt[38] ), .dout(n12372));
  jor  g12093(.dina(n12359), .dinb(asqrt[38] ), .dout(n12373));
  jor  g12094(.dina(n12373), .dinb(n12370), .dout(n12374));
  jnot g12095(.din(n11863), .dout(n12375));
  jnot g12096(.din(n11865), .dout(n12376));
  jand g12097(.dina(asqrt[16] ), .dinb(n11859), .dout(n12377));
  jand g12098(.dina(n12377), .dinb(n12376), .dout(n12378));
  jor  g12099(.dina(n12378), .dinb(n12375), .dout(n12379));
  jnot g12100(.din(n11866), .dout(n12380));
  jand g12101(.dina(n12377), .dinb(n12380), .dout(n12381));
  jnot g12102(.din(n12381), .dout(n12382));
  jand g12103(.dina(n12382), .dinb(n12379), .dout(n12383));
  jand g12104(.dina(n12383), .dinb(n12374), .dout(n12384));
  jor  g12105(.dina(n12384), .dinb(n12372), .dout(n12385));
  jand g12106(.dina(n12385), .dinb(asqrt[39] ), .dout(n12386));
  jxor g12107(.dina(n11867), .dinb(n3907), .dout(n12387));
  jand g12108(.dina(n12387), .dinb(asqrt[16] ), .dout(n12388));
  jxor g12109(.dina(n12388), .dinb(n11877), .dout(n12389));
  jnot g12110(.din(n12389), .dout(n12390));
  jor  g12111(.dina(n12385), .dinb(asqrt[39] ), .dout(n12391));
  jand g12112(.dina(n12391), .dinb(n12390), .dout(n12392));
  jor  g12113(.dina(n12392), .dinb(n12386), .dout(n12393));
  jand g12114(.dina(n12393), .dinb(asqrt[40] ), .dout(n12394));
  jnot g12115(.din(n11882), .dout(n12395));
  jand g12116(.dina(n12395), .dinb(n11880), .dout(n12396));
  jand g12117(.dina(n12396), .dinb(asqrt[16] ), .dout(n12397));
  jxor g12118(.dina(n12397), .dinb(n11890), .dout(n12398));
  jnot g12119(.din(n12398), .dout(n12399));
  jor  g12120(.dina(n12386), .dinb(asqrt[40] ), .dout(n12400));
  jor  g12121(.dina(n12400), .dinb(n12392), .dout(n12401));
  jand g12122(.dina(n12401), .dinb(n12399), .dout(n12402));
  jor  g12123(.dina(n12402), .dinb(n12394), .dout(n12403));
  jand g12124(.dina(n12403), .dinb(asqrt[41] ), .dout(n12404));
  jor  g12125(.dina(n12403), .dinb(asqrt[41] ), .dout(n12405));
  jnot g12126(.din(n11896), .dout(n12406));
  jnot g12127(.din(n11897), .dout(n12407));
  jand g12128(.dina(asqrt[16] ), .dinb(n11893), .dout(n12408));
  jand g12129(.dina(n12408), .dinb(n12407), .dout(n12409));
  jor  g12130(.dina(n12409), .dinb(n12406), .dout(n12410));
  jnot g12131(.din(n11898), .dout(n12411));
  jand g12132(.dina(n12408), .dinb(n12411), .dout(n12412));
  jnot g12133(.din(n12412), .dout(n12413));
  jand g12134(.dina(n12413), .dinb(n12410), .dout(n12414));
  jand g12135(.dina(n12414), .dinb(n12405), .dout(n12415));
  jor  g12136(.dina(n12415), .dinb(n12404), .dout(n12416));
  jand g12137(.dina(n12416), .dinb(asqrt[42] ), .dout(n12417));
  jor  g12138(.dina(n12404), .dinb(asqrt[42] ), .dout(n12418));
  jor  g12139(.dina(n12418), .dinb(n12415), .dout(n12419));
  jnot g12140(.din(n11904), .dout(n12420));
  jnot g12141(.din(n11906), .dout(n12421));
  jand g12142(.dina(asqrt[16] ), .dinb(n11900), .dout(n12422));
  jand g12143(.dina(n12422), .dinb(n12421), .dout(n12423));
  jor  g12144(.dina(n12423), .dinb(n12420), .dout(n12424));
  jnot g12145(.din(n11907), .dout(n12425));
  jand g12146(.dina(n12422), .dinb(n12425), .dout(n12426));
  jnot g12147(.din(n12426), .dout(n12427));
  jand g12148(.dina(n12427), .dinb(n12424), .dout(n12428));
  jand g12149(.dina(n12428), .dinb(n12419), .dout(n12429));
  jor  g12150(.dina(n12429), .dinb(n12417), .dout(n12430));
  jand g12151(.dina(n12430), .dinb(asqrt[43] ), .dout(n12431));
  jxor g12152(.dina(n11908), .dinb(n2870), .dout(n12432));
  jand g12153(.dina(n12432), .dinb(asqrt[16] ), .dout(n12433));
  jxor g12154(.dina(n12433), .dinb(n11918), .dout(n12434));
  jnot g12155(.din(n12434), .dout(n12435));
  jor  g12156(.dina(n12430), .dinb(asqrt[43] ), .dout(n12436));
  jand g12157(.dina(n12436), .dinb(n12435), .dout(n12437));
  jor  g12158(.dina(n12437), .dinb(n12431), .dout(n12438));
  jand g12159(.dina(n12438), .dinb(asqrt[44] ), .dout(n12439));
  jnot g12160(.din(n11923), .dout(n12440));
  jand g12161(.dina(n12440), .dinb(n11921), .dout(n12441));
  jand g12162(.dina(n12441), .dinb(asqrt[16] ), .dout(n12442));
  jxor g12163(.dina(n12442), .dinb(n11931), .dout(n12443));
  jnot g12164(.din(n12443), .dout(n12444));
  jor  g12165(.dina(n12431), .dinb(asqrt[44] ), .dout(n12445));
  jor  g12166(.dina(n12445), .dinb(n12437), .dout(n12446));
  jand g12167(.dina(n12446), .dinb(n12444), .dout(n12447));
  jor  g12168(.dina(n12447), .dinb(n12439), .dout(n12448));
  jand g12169(.dina(n12448), .dinb(asqrt[45] ), .dout(n12449));
  jor  g12170(.dina(n12448), .dinb(asqrt[45] ), .dout(n12450));
  jnot g12171(.din(n11937), .dout(n12451));
  jnot g12172(.din(n11938), .dout(n12452));
  jand g12173(.dina(asqrt[16] ), .dinb(n11934), .dout(n12453));
  jand g12174(.dina(n12453), .dinb(n12452), .dout(n12454));
  jor  g12175(.dina(n12454), .dinb(n12451), .dout(n12455));
  jnot g12176(.din(n11939), .dout(n12456));
  jand g12177(.dina(n12453), .dinb(n12456), .dout(n12457));
  jnot g12178(.din(n12457), .dout(n12458));
  jand g12179(.dina(n12458), .dinb(n12455), .dout(n12459));
  jand g12180(.dina(n12459), .dinb(n12450), .dout(n12460));
  jor  g12181(.dina(n12460), .dinb(n12449), .dout(n12461));
  jand g12182(.dina(n12461), .dinb(asqrt[46] ), .dout(n12462));
  jnot g12183(.din(n11943), .dout(n12463));
  jand g12184(.dina(n12463), .dinb(n11941), .dout(n12464));
  jand g12185(.dina(n12464), .dinb(asqrt[16] ), .dout(n12465));
  jxor g12186(.dina(n12465), .dinb(n11951), .dout(n12466));
  jnot g12187(.din(n12466), .dout(n12467));
  jor  g12188(.dina(n12449), .dinb(asqrt[46] ), .dout(n12468));
  jor  g12189(.dina(n12468), .dinb(n12460), .dout(n12469));
  jand g12190(.dina(n12469), .dinb(n12467), .dout(n12470));
  jor  g12191(.dina(n12470), .dinb(n12462), .dout(n12471));
  jand g12192(.dina(n12471), .dinb(asqrt[47] ), .dout(n12472));
  jor  g12193(.dina(n12471), .dinb(asqrt[47] ), .dout(n12473));
  jand g12194(.dina(n12473), .dinb(n12145), .dout(n12474));
  jor  g12195(.dina(n12474), .dinb(n12472), .dout(n12475));
  jand g12196(.dina(n12475), .dinb(asqrt[48] ), .dout(n12476));
  jor  g12197(.dina(n12472), .dinb(asqrt[48] ), .dout(n12477));
  jor  g12198(.dina(n12477), .dinb(n12474), .dout(n12478));
  jnot g12199(.din(n11963), .dout(n12479));
  jnot g12200(.din(n11965), .dout(n12480));
  jand g12201(.dina(asqrt[16] ), .dinb(n11959), .dout(n12481));
  jand g12202(.dina(n12481), .dinb(n12480), .dout(n12482));
  jor  g12203(.dina(n12482), .dinb(n12479), .dout(n12483));
  jnot g12204(.din(n11966), .dout(n12484));
  jand g12205(.dina(n12481), .dinb(n12484), .dout(n12485));
  jnot g12206(.din(n12485), .dout(n12486));
  jand g12207(.dina(n12486), .dinb(n12483), .dout(n12487));
  jand g12208(.dina(n12487), .dinb(n12478), .dout(n12488));
  jor  g12209(.dina(n12488), .dinb(n12476), .dout(n12489));
  jand g12210(.dina(n12489), .dinb(asqrt[49] ), .dout(n12490));
  jor  g12211(.dina(n12489), .dinb(asqrt[49] ), .dout(n12491));
  jnot g12212(.din(n11971), .dout(n12492));
  jnot g12213(.din(n11972), .dout(n12493));
  jand g12214(.dina(asqrt[16] ), .dinb(n11968), .dout(n12494));
  jand g12215(.dina(n12494), .dinb(n12493), .dout(n12495));
  jor  g12216(.dina(n12495), .dinb(n12492), .dout(n12496));
  jnot g12217(.din(n11973), .dout(n12497));
  jand g12218(.dina(n12494), .dinb(n12497), .dout(n12498));
  jnot g12219(.din(n12498), .dout(n12499));
  jand g12220(.dina(n12499), .dinb(n12496), .dout(n12500));
  jand g12221(.dina(n12500), .dinb(n12491), .dout(n12501));
  jor  g12222(.dina(n12501), .dinb(n12490), .dout(n12502));
  jand g12223(.dina(n12502), .dinb(asqrt[50] ), .dout(n12503));
  jor  g12224(.dina(n12490), .dinb(asqrt[50] ), .dout(n12504));
  jor  g12225(.dina(n12504), .dinb(n12501), .dout(n12505));
  jnot g12226(.din(n11979), .dout(n12506));
  jnot g12227(.din(n11981), .dout(n12507));
  jand g12228(.dina(asqrt[16] ), .dinb(n11975), .dout(n12508));
  jand g12229(.dina(n12508), .dinb(n12507), .dout(n12509));
  jor  g12230(.dina(n12509), .dinb(n12506), .dout(n12510));
  jnot g12231(.din(n11982), .dout(n12511));
  jand g12232(.dina(n12508), .dinb(n12511), .dout(n12512));
  jnot g12233(.din(n12512), .dout(n12513));
  jand g12234(.dina(n12513), .dinb(n12510), .dout(n12514));
  jand g12235(.dina(n12514), .dinb(n12505), .dout(n12515));
  jor  g12236(.dina(n12515), .dinb(n12503), .dout(n12516));
  jand g12237(.dina(n12516), .dinb(asqrt[51] ), .dout(n12517));
  jxor g12238(.dina(n11983), .dinb(n1312), .dout(n12518));
  jand g12239(.dina(n12518), .dinb(asqrt[16] ), .dout(n12519));
  jxor g12240(.dina(n12519), .dinb(n11993), .dout(n12520));
  jnot g12241(.din(n12520), .dout(n12521));
  jor  g12242(.dina(n12516), .dinb(asqrt[51] ), .dout(n12522));
  jand g12243(.dina(n12522), .dinb(n12521), .dout(n12523));
  jor  g12244(.dina(n12523), .dinb(n12517), .dout(n12524));
  jand g12245(.dina(n12524), .dinb(asqrt[52] ), .dout(n12525));
  jnot g12246(.din(n11998), .dout(n12526));
  jand g12247(.dina(n12526), .dinb(n11996), .dout(n12527));
  jand g12248(.dina(n12527), .dinb(asqrt[16] ), .dout(n12528));
  jxor g12249(.dina(n12528), .dinb(n12006), .dout(n12529));
  jnot g12250(.din(n12529), .dout(n12530));
  jor  g12251(.dina(n12517), .dinb(asqrt[52] ), .dout(n12531));
  jor  g12252(.dina(n12531), .dinb(n12523), .dout(n12532));
  jand g12253(.dina(n12532), .dinb(n12530), .dout(n12533));
  jor  g12254(.dina(n12533), .dinb(n12525), .dout(n12534));
  jand g12255(.dina(n12534), .dinb(asqrt[53] ), .dout(n12535));
  jor  g12256(.dina(n12534), .dinb(asqrt[53] ), .dout(n12536));
  jnot g12257(.din(n12012), .dout(n12537));
  jnot g12258(.din(n12013), .dout(n12538));
  jand g12259(.dina(asqrt[16] ), .dinb(n12009), .dout(n12539));
  jand g12260(.dina(n12539), .dinb(n12538), .dout(n12540));
  jor  g12261(.dina(n12540), .dinb(n12537), .dout(n12541));
  jnot g12262(.din(n12014), .dout(n12542));
  jand g12263(.dina(n12539), .dinb(n12542), .dout(n12543));
  jnot g12264(.din(n12543), .dout(n12544));
  jand g12265(.dina(n12544), .dinb(n12541), .dout(n12545));
  jand g12266(.dina(n12545), .dinb(n12536), .dout(n12546));
  jor  g12267(.dina(n12546), .dinb(n12535), .dout(n12547));
  jand g12268(.dina(n12547), .dinb(asqrt[54] ), .dout(n12548));
  jor  g12269(.dina(n12535), .dinb(asqrt[54] ), .dout(n12549));
  jor  g12270(.dina(n12549), .dinb(n12546), .dout(n12550));
  jnot g12271(.din(n12020), .dout(n12551));
  jnot g12272(.din(n12022), .dout(n12552));
  jand g12273(.dina(asqrt[16] ), .dinb(n12016), .dout(n12553));
  jand g12274(.dina(n12553), .dinb(n12552), .dout(n12554));
  jor  g12275(.dina(n12554), .dinb(n12551), .dout(n12555));
  jnot g12276(.din(n12023), .dout(n12556));
  jand g12277(.dina(n12553), .dinb(n12556), .dout(n12557));
  jnot g12278(.din(n12557), .dout(n12558));
  jand g12279(.dina(n12558), .dinb(n12555), .dout(n12559));
  jand g12280(.dina(n12559), .dinb(n12550), .dout(n12560));
  jor  g12281(.dina(n12560), .dinb(n12548), .dout(n12561));
  jand g12282(.dina(n12561), .dinb(asqrt[55] ), .dout(n12562));
  jxor g12283(.dina(n12024), .dinb(n791), .dout(n12563));
  jand g12284(.dina(n12563), .dinb(asqrt[16] ), .dout(n12564));
  jxor g12285(.dina(n12564), .dinb(n12034), .dout(n12565));
  jnot g12286(.din(n12565), .dout(n12566));
  jor  g12287(.dina(n12561), .dinb(asqrt[55] ), .dout(n12567));
  jand g12288(.dina(n12567), .dinb(n12566), .dout(n12568));
  jor  g12289(.dina(n12568), .dinb(n12562), .dout(n12569));
  jand g12290(.dina(n12569), .dinb(asqrt[56] ), .dout(n12570));
  jnot g12291(.din(n12039), .dout(n12571));
  jand g12292(.dina(n12571), .dinb(n12037), .dout(n12572));
  jand g12293(.dina(n12572), .dinb(asqrt[16] ), .dout(n12573));
  jxor g12294(.dina(n12573), .dinb(n12047), .dout(n12574));
  jnot g12295(.din(n12574), .dout(n12575));
  jor  g12296(.dina(n12562), .dinb(asqrt[56] ), .dout(n12576));
  jor  g12297(.dina(n12576), .dinb(n12568), .dout(n12577));
  jand g12298(.dina(n12577), .dinb(n12575), .dout(n12578));
  jor  g12299(.dina(n12578), .dinb(n12570), .dout(n12579));
  jand g12300(.dina(n12579), .dinb(asqrt[57] ), .dout(n12580));
  jor  g12301(.dina(n12579), .dinb(asqrt[57] ), .dout(n12581));
  jnot g12302(.din(n12053), .dout(n12582));
  jnot g12303(.din(n12054), .dout(n12583));
  jand g12304(.dina(asqrt[16] ), .dinb(n12050), .dout(n12584));
  jand g12305(.dina(n12584), .dinb(n12583), .dout(n12585));
  jor  g12306(.dina(n12585), .dinb(n12582), .dout(n12586));
  jnot g12307(.din(n12055), .dout(n12587));
  jand g12308(.dina(n12584), .dinb(n12587), .dout(n12588));
  jnot g12309(.din(n12588), .dout(n12589));
  jand g12310(.dina(n12589), .dinb(n12586), .dout(n12590));
  jand g12311(.dina(n12590), .dinb(n12581), .dout(n12591));
  jor  g12312(.dina(n12591), .dinb(n12580), .dout(n12592));
  jand g12313(.dina(n12592), .dinb(asqrt[58] ), .dout(n12593));
  jor  g12314(.dina(n12580), .dinb(asqrt[58] ), .dout(n12594));
  jor  g12315(.dina(n12594), .dinb(n12591), .dout(n12595));
  jnot g12316(.din(n12061), .dout(n12596));
  jnot g12317(.din(n12063), .dout(n12597));
  jand g12318(.dina(asqrt[16] ), .dinb(n12057), .dout(n12598));
  jand g12319(.dina(n12598), .dinb(n12597), .dout(n12599));
  jor  g12320(.dina(n12599), .dinb(n12596), .dout(n12600));
  jnot g12321(.din(n12064), .dout(n12601));
  jand g12322(.dina(n12598), .dinb(n12601), .dout(n12602));
  jnot g12323(.din(n12602), .dout(n12603));
  jand g12324(.dina(n12603), .dinb(n12600), .dout(n12604));
  jand g12325(.dina(n12604), .dinb(n12595), .dout(n12605));
  jor  g12326(.dina(n12605), .dinb(n12593), .dout(n12606));
  jand g12327(.dina(n12606), .dinb(asqrt[59] ), .dout(n12607));
  jxor g12328(.dina(n12065), .dinb(n425), .dout(n12608));
  jand g12329(.dina(n12608), .dinb(asqrt[16] ), .dout(n12609));
  jxor g12330(.dina(n12609), .dinb(n12075), .dout(n12610));
  jnot g12331(.din(n12610), .dout(n12611));
  jor  g12332(.dina(n12606), .dinb(asqrt[59] ), .dout(n12612));
  jand g12333(.dina(n12612), .dinb(n12611), .dout(n12613));
  jor  g12334(.dina(n12613), .dinb(n12607), .dout(n12614));
  jand g12335(.dina(n12614), .dinb(asqrt[60] ), .dout(n12615));
  jnot g12336(.din(n12080), .dout(n12616));
  jand g12337(.dina(n12616), .dinb(n12078), .dout(n12617));
  jand g12338(.dina(n12617), .dinb(asqrt[16] ), .dout(n12618));
  jxor g12339(.dina(n12618), .dinb(n12088), .dout(n12619));
  jnot g12340(.din(n12619), .dout(n12620));
  jor  g12341(.dina(n12607), .dinb(asqrt[60] ), .dout(n12621));
  jor  g12342(.dina(n12621), .dinb(n12613), .dout(n12622));
  jand g12343(.dina(n12622), .dinb(n12620), .dout(n12623));
  jor  g12344(.dina(n12623), .dinb(n12615), .dout(n12624));
  jand g12345(.dina(n12624), .dinb(asqrt[61] ), .dout(n12625));
  jor  g12346(.dina(n12624), .dinb(asqrt[61] ), .dout(n12626));
  jnot g12347(.din(n12094), .dout(n12627));
  jnot g12348(.din(n12095), .dout(n12628));
  jand g12349(.dina(asqrt[16] ), .dinb(n12091), .dout(n12629));
  jand g12350(.dina(n12629), .dinb(n12628), .dout(n12630));
  jor  g12351(.dina(n12630), .dinb(n12627), .dout(n12631));
  jnot g12352(.din(n12096), .dout(n12632));
  jand g12353(.dina(n12629), .dinb(n12632), .dout(n12633));
  jnot g12354(.din(n12633), .dout(n12634));
  jand g12355(.dina(n12634), .dinb(n12631), .dout(n12635));
  jand g12356(.dina(n12635), .dinb(n12626), .dout(n12636));
  jor  g12357(.dina(n12636), .dinb(n12625), .dout(n12637));
  jand g12358(.dina(n12637), .dinb(asqrt[62] ), .dout(n12638));
  jor  g12359(.dina(n12625), .dinb(asqrt[62] ), .dout(n12639));
  jor  g12360(.dina(n12639), .dinb(n12636), .dout(n12640));
  jnot g12361(.din(n12102), .dout(n12641));
  jnot g12362(.din(n12104), .dout(n12642));
  jand g12363(.dina(asqrt[16] ), .dinb(n12098), .dout(n12643));
  jand g12364(.dina(n12643), .dinb(n12642), .dout(n12644));
  jor  g12365(.dina(n12644), .dinb(n12641), .dout(n12645));
  jnot g12366(.din(n12105), .dout(n12646));
  jand g12367(.dina(n12643), .dinb(n12646), .dout(n12647));
  jnot g12368(.din(n12647), .dout(n12648));
  jand g12369(.dina(n12648), .dinb(n12645), .dout(n12649));
  jand g12370(.dina(n12649), .dinb(n12640), .dout(n12650));
  jor  g12371(.dina(n12650), .dinb(n12638), .dout(n12651));
  jxor g12372(.dina(n12106), .dinb(n199), .dout(n12652));
  jand g12373(.dina(n12652), .dinb(asqrt[16] ), .dout(n12653));
  jxor g12374(.dina(n12653), .dinb(n12116), .dout(n12654));
  jnot g12375(.din(n12118), .dout(n12655));
  jand g12376(.dina(asqrt[16] ), .dinb(n12125), .dout(n12656));
  jand g12377(.dina(n12656), .dinb(n12655), .dout(n12657));
  jor  g12378(.dina(n12657), .dinb(n12133), .dout(n12658));
  jor  g12379(.dina(n12658), .dinb(n12654), .dout(n12659));
  jnot g12380(.din(n12659), .dout(n12660));
  jand g12381(.dina(n12660), .dinb(n12651), .dout(n12661));
  jor  g12382(.dina(n12661), .dinb(asqrt[63] ), .dout(n12662));
  jnot g12383(.din(n12654), .dout(n12663));
  jor  g12384(.dina(n12663), .dinb(n12651), .dout(n12664));
  jor  g12385(.dina(n12656), .dinb(n12655), .dout(n12665));
  jand g12386(.dina(n12125), .dinb(n12655), .dout(n12666));
  jor  g12387(.dina(n12666), .dinb(n194), .dout(n12667));
  jnot g12388(.din(n12667), .dout(n12668));
  jand g12389(.dina(n12668), .dinb(n12665), .dout(n12669));
  jnot g12390(.din(asqrt[16] ), .dout(n12670));
  jnot g12391(.din(n12669), .dout(n12673));
  jand g12392(.dina(n12673), .dinb(n12664), .dout(n12674));
  jand g12393(.dina(n12674), .dinb(n12662), .dout(n12675));
  jxor g12394(.dina(n12471), .dinb(n1646), .dout(n12676));
  jor  g12395(.dina(n12676), .dinb(n12675), .dout(n12677));
  jxor g12396(.dina(n12677), .dinb(n12146), .dout(n12678));
  jnot g12397(.din(n12678), .dout(n12679));
  jor  g12398(.dina(n12675), .dinb(n12148), .dout(n12680));
  jnot g12399(.din(a[28] ), .dout(n12681));
  jnot g12400(.din(a[29] ), .dout(n12682));
  jand g12401(.dina(n12148), .dinb(n12682), .dout(n12683));
  jand g12402(.dina(n12683), .dinb(n12681), .dout(n12684));
  jnot g12403(.din(n12684), .dout(n12685));
  jand g12404(.dina(n12685), .dinb(n12680), .dout(n12686));
  jor  g12405(.dina(n12686), .dinb(n12670), .dout(n12687));
  jor  g12406(.dina(n12675), .dinb(a[30] ), .dout(n12688));
  jxor g12407(.dina(n12688), .dinb(n12149), .dout(n12689));
  jand g12408(.dina(n12686), .dinb(n12670), .dout(n12690));
  jor  g12409(.dina(n12690), .dinb(n12689), .dout(n12691));
  jand g12410(.dina(n12691), .dinb(n12687), .dout(n12692));
  jor  g12411(.dina(n12692), .dinb(n11662), .dout(n12693));
  jand g12412(.dina(n12687), .dinb(n11662), .dout(n12694));
  jand g12413(.dina(n12694), .dinb(n12691), .dout(n12695));
  jor  g12414(.dina(n12688), .dinb(a[31] ), .dout(n12696));
  jnot g12415(.din(n12662), .dout(n12697));
  jnot g12416(.din(n12664), .dout(n12698));
  jor  g12417(.dina(n12669), .dinb(n12670), .dout(n12699));
  jor  g12418(.dina(n12699), .dinb(n12698), .dout(n12700));
  jor  g12419(.dina(n12700), .dinb(n12697), .dout(n12701));
  jand g12420(.dina(n12701), .dinb(n12696), .dout(n12702));
  jxor g12421(.dina(n12702), .dinb(n11667), .dout(n12703));
  jor  g12422(.dina(n12703), .dinb(n12695), .dout(n12704));
  jand g12423(.dina(n12704), .dinb(n12693), .dout(n12705));
  jor  g12424(.dina(n12705), .dinb(n11657), .dout(n12706));
  jand g12425(.dina(n12705), .dinb(n11657), .dout(n12707));
  jxor g12426(.dina(n12152), .dinb(n11662), .dout(n12708));
  jor  g12427(.dina(n12708), .dinb(n12675), .dout(n12709));
  jxor g12428(.dina(n12709), .dinb(n12155), .dout(n12710));
  jor  g12429(.dina(n12710), .dinb(n12707), .dout(n12711));
  jand g12430(.dina(n12711), .dinb(n12706), .dout(n12712));
  jor  g12431(.dina(n12712), .dinb(n10701), .dout(n12713));
  jnot g12432(.din(n12161), .dout(n12714));
  jor  g12433(.dina(n12714), .dinb(n12159), .dout(n12715));
  jor  g12434(.dina(n12715), .dinb(n12675), .dout(n12716));
  jxor g12435(.dina(n12716), .dinb(n12170), .dout(n12717));
  jand g12436(.dina(n12706), .dinb(n10701), .dout(n12718));
  jand g12437(.dina(n12718), .dinb(n12711), .dout(n12719));
  jor  g12438(.dina(n12719), .dinb(n12717), .dout(n12720));
  jand g12439(.dina(n12720), .dinb(n12713), .dout(n12721));
  jor  g12440(.dina(n12721), .dinb(n10696), .dout(n12722));
  jand g12441(.dina(n12721), .dinb(n10696), .dout(n12723));
  jxor g12442(.dina(n12172), .dinb(n10701), .dout(n12724));
  jor  g12443(.dina(n12724), .dinb(n12675), .dout(n12725));
  jxor g12444(.dina(n12725), .dinb(n12177), .dout(n12726));
  jnot g12445(.din(n12726), .dout(n12727));
  jor  g12446(.dina(n12727), .dinb(n12723), .dout(n12728));
  jand g12447(.dina(n12728), .dinb(n12722), .dout(n12729));
  jor  g12448(.dina(n12729), .dinb(n9774), .dout(n12730));
  jand g12449(.dina(n12722), .dinb(n9774), .dout(n12731));
  jand g12450(.dina(n12731), .dinb(n12728), .dout(n12732));
  jnot g12451(.din(n12181), .dout(n12733));
  jnot g12452(.din(n12675), .dout(asqrt[15] ));
  jand g12453(.dina(asqrt[15] ), .dinb(n12733), .dout(n12735));
  jand g12454(.dina(n12735), .dinb(n12188), .dout(n12736));
  jor  g12455(.dina(n12736), .dinb(n12186), .dout(n12737));
  jand g12456(.dina(n12735), .dinb(n12189), .dout(n12738));
  jnot g12457(.din(n12738), .dout(n12739));
  jand g12458(.dina(n12739), .dinb(n12737), .dout(n12740));
  jnot g12459(.din(n12740), .dout(n12741));
  jor  g12460(.dina(n12741), .dinb(n12732), .dout(n12742));
  jand g12461(.dina(n12742), .dinb(n12730), .dout(n12743));
  jor  g12462(.dina(n12743), .dinb(n9769), .dout(n12744));
  jand g12463(.dina(n12743), .dinb(n9769), .dout(n12745));
  jnot g12464(.din(n12196), .dout(n12746));
  jxor g12465(.dina(n12190), .dinb(n9774), .dout(n12747));
  jor  g12466(.dina(n12747), .dinb(n12675), .dout(n12748));
  jxor g12467(.dina(n12748), .dinb(n12746), .dout(n12749));
  jnot g12468(.din(n12749), .dout(n12750));
  jor  g12469(.dina(n12750), .dinb(n12745), .dout(n12751));
  jand g12470(.dina(n12751), .dinb(n12744), .dout(n12752));
  jor  g12471(.dina(n12752), .dinb(n8898), .dout(n12753));
  jnot g12472(.din(n12201), .dout(n12754));
  jor  g12473(.dina(n12754), .dinb(n12199), .dout(n12755));
  jor  g12474(.dina(n12755), .dinb(n12675), .dout(n12756));
  jxor g12475(.dina(n12756), .dinb(n12210), .dout(n12757));
  jand g12476(.dina(n12744), .dinb(n8898), .dout(n12758));
  jand g12477(.dina(n12758), .dinb(n12751), .dout(n12759));
  jor  g12478(.dina(n12759), .dinb(n12757), .dout(n12760));
  jand g12479(.dina(n12760), .dinb(n12753), .dout(n12761));
  jor  g12480(.dina(n12761), .dinb(n8893), .dout(n12762));
  jand g12481(.dina(n12761), .dinb(n8893), .dout(n12763));
  jnot g12482(.din(n12217), .dout(n12764));
  jxor g12483(.dina(n12212), .dinb(n8898), .dout(n12765));
  jor  g12484(.dina(n12765), .dinb(n12675), .dout(n12766));
  jxor g12485(.dina(n12766), .dinb(n12764), .dout(n12767));
  jnot g12486(.din(n12767), .dout(n12768));
  jor  g12487(.dina(n12768), .dinb(n12763), .dout(n12769));
  jand g12488(.dina(n12769), .dinb(n12762), .dout(n12770));
  jor  g12489(.dina(n12770), .dinb(n8058), .dout(n12771));
  jand g12490(.dina(n12762), .dinb(n8058), .dout(n12772));
  jand g12491(.dina(n12772), .dinb(n12769), .dout(n12773));
  jnot g12492(.din(n12220), .dout(n12774));
  jand g12493(.dina(asqrt[15] ), .dinb(n12774), .dout(n12775));
  jand g12494(.dina(n12775), .dinb(n12227), .dout(n12776));
  jor  g12495(.dina(n12776), .dinb(n12225), .dout(n12777));
  jand g12496(.dina(n12775), .dinb(n12228), .dout(n12778));
  jnot g12497(.din(n12778), .dout(n12779));
  jand g12498(.dina(n12779), .dinb(n12777), .dout(n12780));
  jnot g12499(.din(n12780), .dout(n12781));
  jor  g12500(.dina(n12781), .dinb(n12773), .dout(n12782));
  jand g12501(.dina(n12782), .dinb(n12771), .dout(n12783));
  jor  g12502(.dina(n12783), .dinb(n8053), .dout(n12784));
  jxor g12503(.dina(n12229), .dinb(n8058), .dout(n12785));
  jor  g12504(.dina(n12785), .dinb(n12675), .dout(n12786));
  jxor g12505(.dina(n12786), .dinb(n12234), .dout(n12787));
  jand g12506(.dina(n12783), .dinb(n8053), .dout(n12788));
  jor  g12507(.dina(n12788), .dinb(n12787), .dout(n12789));
  jand g12508(.dina(n12789), .dinb(n12784), .dout(n12790));
  jor  g12509(.dina(n12790), .dinb(n7265), .dout(n12791));
  jnot g12510(.din(n12239), .dout(n12792));
  jor  g12511(.dina(n12792), .dinb(n12237), .dout(n12793));
  jor  g12512(.dina(n12793), .dinb(n12675), .dout(n12794));
  jxor g12513(.dina(n12794), .dinb(n12248), .dout(n12795));
  jand g12514(.dina(n12784), .dinb(n7265), .dout(n12796));
  jand g12515(.dina(n12796), .dinb(n12789), .dout(n12797));
  jor  g12516(.dina(n12797), .dinb(n12795), .dout(n12798));
  jand g12517(.dina(n12798), .dinb(n12791), .dout(n12799));
  jor  g12518(.dina(n12799), .dinb(n7260), .dout(n12800));
  jand g12519(.dina(n12799), .dinb(n7260), .dout(n12801));
  jnot g12520(.din(n12251), .dout(n12802));
  jand g12521(.dina(asqrt[15] ), .dinb(n12802), .dout(n12803));
  jand g12522(.dina(n12803), .dinb(n12256), .dout(n12804));
  jor  g12523(.dina(n12804), .dinb(n12255), .dout(n12805));
  jand g12524(.dina(n12803), .dinb(n12257), .dout(n12806));
  jnot g12525(.din(n12806), .dout(n12807));
  jand g12526(.dina(n12807), .dinb(n12805), .dout(n12808));
  jnot g12527(.din(n12808), .dout(n12809));
  jor  g12528(.dina(n12809), .dinb(n12801), .dout(n12810));
  jand g12529(.dina(n12810), .dinb(n12800), .dout(n12811));
  jor  g12530(.dina(n12811), .dinb(n6505), .dout(n12812));
  jand g12531(.dina(n12800), .dinb(n6505), .dout(n12813));
  jand g12532(.dina(n12813), .dinb(n12810), .dout(n12814));
  jnot g12533(.din(n12259), .dout(n12815));
  jand g12534(.dina(asqrt[15] ), .dinb(n12815), .dout(n12816));
  jand g12535(.dina(n12816), .dinb(n12266), .dout(n12817));
  jor  g12536(.dina(n12817), .dinb(n12264), .dout(n12818));
  jand g12537(.dina(n12816), .dinb(n12267), .dout(n12819));
  jnot g12538(.din(n12819), .dout(n12820));
  jand g12539(.dina(n12820), .dinb(n12818), .dout(n12821));
  jnot g12540(.din(n12821), .dout(n12822));
  jor  g12541(.dina(n12822), .dinb(n12814), .dout(n12823));
  jand g12542(.dina(n12823), .dinb(n12812), .dout(n12824));
  jor  g12543(.dina(n12824), .dinb(n6500), .dout(n12825));
  jxor g12544(.dina(n12268), .dinb(n6505), .dout(n12826));
  jor  g12545(.dina(n12826), .dinb(n12675), .dout(n12827));
  jxor g12546(.dina(n12827), .dinb(n12279), .dout(n12828));
  jand g12547(.dina(n12824), .dinb(n6500), .dout(n12829));
  jor  g12548(.dina(n12829), .dinb(n12828), .dout(n12830));
  jand g12549(.dina(n12830), .dinb(n12825), .dout(n12831));
  jor  g12550(.dina(n12831), .dinb(n5793), .dout(n12832));
  jnot g12551(.din(n12284), .dout(n12833));
  jor  g12552(.dina(n12833), .dinb(n12282), .dout(n12834));
  jor  g12553(.dina(n12834), .dinb(n12675), .dout(n12835));
  jxor g12554(.dina(n12835), .dinb(n12293), .dout(n12836));
  jand g12555(.dina(n12825), .dinb(n5793), .dout(n12837));
  jand g12556(.dina(n12837), .dinb(n12830), .dout(n12838));
  jor  g12557(.dina(n12838), .dinb(n12836), .dout(n12839));
  jand g12558(.dina(n12839), .dinb(n12832), .dout(n12840));
  jor  g12559(.dina(n12840), .dinb(n5788), .dout(n12841));
  jand g12560(.dina(n12840), .dinb(n5788), .dout(n12842));
  jnot g12561(.din(n12296), .dout(n12843));
  jand g12562(.dina(asqrt[15] ), .dinb(n12843), .dout(n12844));
  jand g12563(.dina(n12844), .dinb(n12301), .dout(n12845));
  jor  g12564(.dina(n12845), .dinb(n12300), .dout(n12846));
  jand g12565(.dina(n12844), .dinb(n12302), .dout(n12847));
  jnot g12566(.din(n12847), .dout(n12848));
  jand g12567(.dina(n12848), .dinb(n12846), .dout(n12849));
  jnot g12568(.din(n12849), .dout(n12850));
  jor  g12569(.dina(n12850), .dinb(n12842), .dout(n12851));
  jand g12570(.dina(n12851), .dinb(n12841), .dout(n12852));
  jor  g12571(.dina(n12852), .dinb(n5121), .dout(n12853));
  jand g12572(.dina(n12841), .dinb(n5121), .dout(n12854));
  jand g12573(.dina(n12854), .dinb(n12851), .dout(n12855));
  jnot g12574(.din(n12304), .dout(n12856));
  jand g12575(.dina(asqrt[15] ), .dinb(n12856), .dout(n12857));
  jand g12576(.dina(n12857), .dinb(n12311), .dout(n12858));
  jor  g12577(.dina(n12858), .dinb(n12309), .dout(n12859));
  jand g12578(.dina(n12857), .dinb(n12312), .dout(n12860));
  jnot g12579(.din(n12860), .dout(n12861));
  jand g12580(.dina(n12861), .dinb(n12859), .dout(n12862));
  jnot g12581(.din(n12862), .dout(n12863));
  jor  g12582(.dina(n12863), .dinb(n12855), .dout(n12864));
  jand g12583(.dina(n12864), .dinb(n12853), .dout(n12865));
  jor  g12584(.dina(n12865), .dinb(n5116), .dout(n12866));
  jxor g12585(.dina(n12313), .dinb(n5121), .dout(n12867));
  jor  g12586(.dina(n12867), .dinb(n12675), .dout(n12868));
  jxor g12587(.dina(n12868), .dinb(n12324), .dout(n12869));
  jand g12588(.dina(n12865), .dinb(n5116), .dout(n12870));
  jor  g12589(.dina(n12870), .dinb(n12869), .dout(n12871));
  jand g12590(.dina(n12871), .dinb(n12866), .dout(n12872));
  jor  g12591(.dina(n12872), .dinb(n4499), .dout(n12873));
  jnot g12592(.din(n12329), .dout(n12874));
  jor  g12593(.dina(n12874), .dinb(n12327), .dout(n12875));
  jor  g12594(.dina(n12875), .dinb(n12675), .dout(n12876));
  jxor g12595(.dina(n12876), .dinb(n12338), .dout(n12877));
  jand g12596(.dina(n12866), .dinb(n4499), .dout(n12878));
  jand g12597(.dina(n12878), .dinb(n12871), .dout(n12879));
  jor  g12598(.dina(n12879), .dinb(n12877), .dout(n12880));
  jand g12599(.dina(n12880), .dinb(n12873), .dout(n12881));
  jor  g12600(.dina(n12881), .dinb(n4494), .dout(n12882));
  jand g12601(.dina(n12881), .dinb(n4494), .dout(n12883));
  jnot g12602(.din(n12341), .dout(n12884));
  jand g12603(.dina(asqrt[15] ), .dinb(n12884), .dout(n12885));
  jand g12604(.dina(n12885), .dinb(n12346), .dout(n12886));
  jor  g12605(.dina(n12886), .dinb(n12345), .dout(n12887));
  jand g12606(.dina(n12885), .dinb(n12347), .dout(n12888));
  jnot g12607(.din(n12888), .dout(n12889));
  jand g12608(.dina(n12889), .dinb(n12887), .dout(n12890));
  jnot g12609(.din(n12890), .dout(n12891));
  jor  g12610(.dina(n12891), .dinb(n12883), .dout(n12892));
  jand g12611(.dina(n12892), .dinb(n12882), .dout(n12893));
  jor  g12612(.dina(n12893), .dinb(n3912), .dout(n12894));
  jand g12613(.dina(n12882), .dinb(n3912), .dout(n12895));
  jand g12614(.dina(n12895), .dinb(n12892), .dout(n12896));
  jnot g12615(.din(n12349), .dout(n12897));
  jand g12616(.dina(asqrt[15] ), .dinb(n12897), .dout(n12898));
  jand g12617(.dina(n12898), .dinb(n12356), .dout(n12899));
  jor  g12618(.dina(n12899), .dinb(n12354), .dout(n12900));
  jand g12619(.dina(n12898), .dinb(n12357), .dout(n12901));
  jnot g12620(.din(n12901), .dout(n12902));
  jand g12621(.dina(n12902), .dinb(n12900), .dout(n12903));
  jnot g12622(.din(n12903), .dout(n12904));
  jor  g12623(.dina(n12904), .dinb(n12896), .dout(n12905));
  jand g12624(.dina(n12905), .dinb(n12894), .dout(n12906));
  jor  g12625(.dina(n12906), .dinb(n3907), .dout(n12907));
  jxor g12626(.dina(n12358), .dinb(n3912), .dout(n12908));
  jor  g12627(.dina(n12908), .dinb(n12675), .dout(n12909));
  jxor g12628(.dina(n12909), .dinb(n12369), .dout(n12910));
  jand g12629(.dina(n12906), .dinb(n3907), .dout(n12911));
  jor  g12630(.dina(n12911), .dinb(n12910), .dout(n12912));
  jand g12631(.dina(n12912), .dinb(n12907), .dout(n12913));
  jor  g12632(.dina(n12913), .dinb(n3376), .dout(n12914));
  jnot g12633(.din(n12374), .dout(n12915));
  jor  g12634(.dina(n12915), .dinb(n12372), .dout(n12916));
  jor  g12635(.dina(n12916), .dinb(n12675), .dout(n12917));
  jxor g12636(.dina(n12917), .dinb(n12383), .dout(n12918));
  jand g12637(.dina(n12907), .dinb(n3376), .dout(n12919));
  jand g12638(.dina(n12919), .dinb(n12912), .dout(n12920));
  jor  g12639(.dina(n12920), .dinb(n12918), .dout(n12921));
  jand g12640(.dina(n12921), .dinb(n12914), .dout(n12922));
  jor  g12641(.dina(n12922), .dinb(n3371), .dout(n12923));
  jand g12642(.dina(n12922), .dinb(n3371), .dout(n12924));
  jnot g12643(.din(n12386), .dout(n12925));
  jand g12644(.dina(asqrt[15] ), .dinb(n12925), .dout(n12926));
  jand g12645(.dina(n12926), .dinb(n12391), .dout(n12927));
  jor  g12646(.dina(n12927), .dinb(n12390), .dout(n12928));
  jand g12647(.dina(n12926), .dinb(n12392), .dout(n12929));
  jnot g12648(.din(n12929), .dout(n12930));
  jand g12649(.dina(n12930), .dinb(n12928), .dout(n12931));
  jnot g12650(.din(n12931), .dout(n12932));
  jor  g12651(.dina(n12932), .dinb(n12924), .dout(n12933));
  jand g12652(.dina(n12933), .dinb(n12923), .dout(n12934));
  jor  g12653(.dina(n12934), .dinb(n2875), .dout(n12935));
  jand g12654(.dina(n12923), .dinb(n2875), .dout(n12936));
  jand g12655(.dina(n12936), .dinb(n12933), .dout(n12937));
  jnot g12656(.din(n12394), .dout(n12938));
  jand g12657(.dina(asqrt[15] ), .dinb(n12938), .dout(n12939));
  jand g12658(.dina(n12939), .dinb(n12401), .dout(n12940));
  jor  g12659(.dina(n12940), .dinb(n12399), .dout(n12941));
  jand g12660(.dina(n12939), .dinb(n12402), .dout(n12942));
  jnot g12661(.din(n12942), .dout(n12943));
  jand g12662(.dina(n12943), .dinb(n12941), .dout(n12944));
  jnot g12663(.din(n12944), .dout(n12945));
  jor  g12664(.dina(n12945), .dinb(n12937), .dout(n12946));
  jand g12665(.dina(n12946), .dinb(n12935), .dout(n12947));
  jor  g12666(.dina(n12947), .dinb(n2870), .dout(n12948));
  jxor g12667(.dina(n12403), .dinb(n2875), .dout(n12949));
  jor  g12668(.dina(n12949), .dinb(n12675), .dout(n12950));
  jxor g12669(.dina(n12950), .dinb(n12414), .dout(n12951));
  jand g12670(.dina(n12947), .dinb(n2870), .dout(n12952));
  jor  g12671(.dina(n12952), .dinb(n12951), .dout(n12953));
  jand g12672(.dina(n12953), .dinb(n12948), .dout(n12954));
  jor  g12673(.dina(n12954), .dinb(n2425), .dout(n12955));
  jnot g12674(.din(n12419), .dout(n12956));
  jor  g12675(.dina(n12956), .dinb(n12417), .dout(n12957));
  jor  g12676(.dina(n12957), .dinb(n12675), .dout(n12958));
  jxor g12677(.dina(n12958), .dinb(n12428), .dout(n12959));
  jand g12678(.dina(n12948), .dinb(n2425), .dout(n12960));
  jand g12679(.dina(n12960), .dinb(n12953), .dout(n12961));
  jor  g12680(.dina(n12961), .dinb(n12959), .dout(n12962));
  jand g12681(.dina(n12962), .dinb(n12955), .dout(n12963));
  jor  g12682(.dina(n12963), .dinb(n2420), .dout(n12964));
  jand g12683(.dina(n12963), .dinb(n2420), .dout(n12965));
  jnot g12684(.din(n12431), .dout(n12966));
  jand g12685(.dina(asqrt[15] ), .dinb(n12966), .dout(n12967));
  jand g12686(.dina(n12967), .dinb(n12436), .dout(n12968));
  jor  g12687(.dina(n12968), .dinb(n12435), .dout(n12969));
  jand g12688(.dina(n12967), .dinb(n12437), .dout(n12970));
  jnot g12689(.din(n12970), .dout(n12971));
  jand g12690(.dina(n12971), .dinb(n12969), .dout(n12972));
  jnot g12691(.din(n12972), .dout(n12973));
  jor  g12692(.dina(n12973), .dinb(n12965), .dout(n12974));
  jand g12693(.dina(n12974), .dinb(n12964), .dout(n12975));
  jor  g12694(.dina(n12975), .dinb(n2010), .dout(n12976));
  jand g12695(.dina(n12964), .dinb(n2010), .dout(n12977));
  jand g12696(.dina(n12977), .dinb(n12974), .dout(n12978));
  jnot g12697(.din(n12439), .dout(n12979));
  jand g12698(.dina(asqrt[15] ), .dinb(n12979), .dout(n12980));
  jand g12699(.dina(n12980), .dinb(n12446), .dout(n12981));
  jor  g12700(.dina(n12981), .dinb(n12444), .dout(n12982));
  jand g12701(.dina(n12980), .dinb(n12447), .dout(n12983));
  jnot g12702(.din(n12983), .dout(n12984));
  jand g12703(.dina(n12984), .dinb(n12982), .dout(n12985));
  jnot g12704(.din(n12985), .dout(n12986));
  jor  g12705(.dina(n12986), .dinb(n12978), .dout(n12987));
  jand g12706(.dina(n12987), .dinb(n12976), .dout(n12988));
  jor  g12707(.dina(n12988), .dinb(n2005), .dout(n12989));
  jxor g12708(.dina(n12448), .dinb(n2010), .dout(n12990));
  jor  g12709(.dina(n12990), .dinb(n12675), .dout(n12991));
  jxor g12710(.dina(n12991), .dinb(n12459), .dout(n12992));
  jand g12711(.dina(n12988), .dinb(n2005), .dout(n12993));
  jor  g12712(.dina(n12993), .dinb(n12992), .dout(n12994));
  jand g12713(.dina(n12994), .dinb(n12989), .dout(n12995));
  jor  g12714(.dina(n12995), .dinb(n1646), .dout(n12996));
  jand g12715(.dina(n12989), .dinb(n1646), .dout(n12997));
  jand g12716(.dina(n12997), .dinb(n12994), .dout(n12998));
  jnot g12717(.din(n12462), .dout(n12999));
  jand g12718(.dina(asqrt[15] ), .dinb(n12999), .dout(n13000));
  jand g12719(.dina(n13000), .dinb(n12469), .dout(n13001));
  jor  g12720(.dina(n13001), .dinb(n12467), .dout(n13002));
  jand g12721(.dina(n13000), .dinb(n12470), .dout(n13003));
  jnot g12722(.din(n13003), .dout(n13004));
  jand g12723(.dina(n13004), .dinb(n13002), .dout(n13005));
  jnot g12724(.din(n13005), .dout(n13006));
  jor  g12725(.dina(n13006), .dinb(n12998), .dout(n13007));
  jand g12726(.dina(n13007), .dinb(n12996), .dout(n13008));
  jor  g12727(.dina(n13008), .dinb(n1641), .dout(n13009));
  jand g12728(.dina(n13008), .dinb(n1641), .dout(n13010));
  jor  g12729(.dina(n13010), .dinb(n12679), .dout(n13011));
  jand g12730(.dina(n13011), .dinb(n13009), .dout(n13012));
  jor  g12731(.dina(n13012), .dinb(n1317), .dout(n13013));
  jnot g12732(.din(n12478), .dout(n13014));
  jor  g12733(.dina(n13014), .dinb(n12476), .dout(n13015));
  jor  g12734(.dina(n13015), .dinb(n12675), .dout(n13016));
  jxor g12735(.dina(n13016), .dinb(n12487), .dout(n13017));
  jand g12736(.dina(n13009), .dinb(n1317), .dout(n13018));
  jand g12737(.dina(n13018), .dinb(n13011), .dout(n13019));
  jor  g12738(.dina(n13019), .dinb(n13017), .dout(n13020));
  jand g12739(.dina(n13020), .dinb(n13013), .dout(n13021));
  jor  g12740(.dina(n13021), .dinb(n1312), .dout(n13022));
  jxor g12741(.dina(n12489), .dinb(n1317), .dout(n13023));
  jor  g12742(.dina(n13023), .dinb(n12675), .dout(n13024));
  jxor g12743(.dina(n13024), .dinb(n12500), .dout(n13025));
  jand g12744(.dina(n13021), .dinb(n1312), .dout(n13026));
  jor  g12745(.dina(n13026), .dinb(n13025), .dout(n13027));
  jand g12746(.dina(n13027), .dinb(n13022), .dout(n13028));
  jor  g12747(.dina(n13028), .dinb(n1039), .dout(n13029));
  jnot g12748(.din(n12505), .dout(n13030));
  jor  g12749(.dina(n13030), .dinb(n12503), .dout(n13031));
  jor  g12750(.dina(n13031), .dinb(n12675), .dout(n13032));
  jxor g12751(.dina(n13032), .dinb(n12514), .dout(n13033));
  jand g12752(.dina(n13022), .dinb(n1039), .dout(n13034));
  jand g12753(.dina(n13034), .dinb(n13027), .dout(n13035));
  jor  g12754(.dina(n13035), .dinb(n13033), .dout(n13036));
  jand g12755(.dina(n13036), .dinb(n13029), .dout(n13037));
  jor  g12756(.dina(n13037), .dinb(n1034), .dout(n13038));
  jand g12757(.dina(n13037), .dinb(n1034), .dout(n13039));
  jnot g12758(.din(n12517), .dout(n13040));
  jand g12759(.dina(asqrt[15] ), .dinb(n13040), .dout(n13041));
  jand g12760(.dina(n13041), .dinb(n12522), .dout(n13042));
  jor  g12761(.dina(n13042), .dinb(n12521), .dout(n13043));
  jand g12762(.dina(n13041), .dinb(n12523), .dout(n13044));
  jnot g12763(.din(n13044), .dout(n13045));
  jand g12764(.dina(n13045), .dinb(n13043), .dout(n13046));
  jnot g12765(.din(n13046), .dout(n13047));
  jor  g12766(.dina(n13047), .dinb(n13039), .dout(n13048));
  jand g12767(.dina(n13048), .dinb(n13038), .dout(n13049));
  jor  g12768(.dina(n13049), .dinb(n796), .dout(n13050));
  jand g12769(.dina(n13038), .dinb(n796), .dout(n13051));
  jand g12770(.dina(n13051), .dinb(n13048), .dout(n13052));
  jnot g12771(.din(n12525), .dout(n13053));
  jand g12772(.dina(asqrt[15] ), .dinb(n13053), .dout(n13054));
  jand g12773(.dina(n13054), .dinb(n12532), .dout(n13055));
  jor  g12774(.dina(n13055), .dinb(n12530), .dout(n13056));
  jand g12775(.dina(n13054), .dinb(n12533), .dout(n13057));
  jnot g12776(.din(n13057), .dout(n13058));
  jand g12777(.dina(n13058), .dinb(n13056), .dout(n13059));
  jnot g12778(.din(n13059), .dout(n13060));
  jor  g12779(.dina(n13060), .dinb(n13052), .dout(n13061));
  jand g12780(.dina(n13061), .dinb(n13050), .dout(n13062));
  jor  g12781(.dina(n13062), .dinb(n791), .dout(n13063));
  jxor g12782(.dina(n12534), .dinb(n796), .dout(n13064));
  jor  g12783(.dina(n13064), .dinb(n12675), .dout(n13065));
  jxor g12784(.dina(n13065), .dinb(n12545), .dout(n13066));
  jand g12785(.dina(n13062), .dinb(n791), .dout(n13067));
  jor  g12786(.dina(n13067), .dinb(n13066), .dout(n13068));
  jand g12787(.dina(n13068), .dinb(n13063), .dout(n13069));
  jor  g12788(.dina(n13069), .dinb(n595), .dout(n13070));
  jnot g12789(.din(n12550), .dout(n13071));
  jor  g12790(.dina(n13071), .dinb(n12548), .dout(n13072));
  jor  g12791(.dina(n13072), .dinb(n12675), .dout(n13073));
  jxor g12792(.dina(n13073), .dinb(n12559), .dout(n13074));
  jand g12793(.dina(n13063), .dinb(n595), .dout(n13075));
  jand g12794(.dina(n13075), .dinb(n13068), .dout(n13076));
  jor  g12795(.dina(n13076), .dinb(n13074), .dout(n13077));
  jand g12796(.dina(n13077), .dinb(n13070), .dout(n13078));
  jor  g12797(.dina(n13078), .dinb(n590), .dout(n13079));
  jand g12798(.dina(n13078), .dinb(n590), .dout(n13080));
  jnot g12799(.din(n12562), .dout(n13081));
  jand g12800(.dina(asqrt[15] ), .dinb(n13081), .dout(n13082));
  jand g12801(.dina(n13082), .dinb(n12567), .dout(n13083));
  jor  g12802(.dina(n13083), .dinb(n12566), .dout(n13084));
  jand g12803(.dina(n13082), .dinb(n12568), .dout(n13085));
  jnot g12804(.din(n13085), .dout(n13086));
  jand g12805(.dina(n13086), .dinb(n13084), .dout(n13087));
  jnot g12806(.din(n13087), .dout(n13088));
  jor  g12807(.dina(n13088), .dinb(n13080), .dout(n13089));
  jand g12808(.dina(n13089), .dinb(n13079), .dout(n13090));
  jor  g12809(.dina(n13090), .dinb(n430), .dout(n13091));
  jand g12810(.dina(n13079), .dinb(n430), .dout(n13092));
  jand g12811(.dina(n13092), .dinb(n13089), .dout(n13093));
  jnot g12812(.din(n12570), .dout(n13094));
  jand g12813(.dina(asqrt[15] ), .dinb(n13094), .dout(n13095));
  jand g12814(.dina(n13095), .dinb(n12577), .dout(n13096));
  jor  g12815(.dina(n13096), .dinb(n12575), .dout(n13097));
  jand g12816(.dina(n13095), .dinb(n12578), .dout(n13098));
  jnot g12817(.din(n13098), .dout(n13099));
  jand g12818(.dina(n13099), .dinb(n13097), .dout(n13100));
  jnot g12819(.din(n13100), .dout(n13101));
  jor  g12820(.dina(n13101), .dinb(n13093), .dout(n13102));
  jand g12821(.dina(n13102), .dinb(n13091), .dout(n13103));
  jor  g12822(.dina(n13103), .dinb(n425), .dout(n13104));
  jxor g12823(.dina(n12579), .dinb(n430), .dout(n13105));
  jor  g12824(.dina(n13105), .dinb(n12675), .dout(n13106));
  jxor g12825(.dina(n13106), .dinb(n12590), .dout(n13107));
  jand g12826(.dina(n13103), .dinb(n425), .dout(n13108));
  jor  g12827(.dina(n13108), .dinb(n13107), .dout(n13109));
  jand g12828(.dina(n13109), .dinb(n13104), .dout(n13110));
  jor  g12829(.dina(n13110), .dinb(n305), .dout(n13111));
  jnot g12830(.din(n12595), .dout(n13112));
  jor  g12831(.dina(n13112), .dinb(n12593), .dout(n13113));
  jor  g12832(.dina(n13113), .dinb(n12675), .dout(n13114));
  jxor g12833(.dina(n13114), .dinb(n12604), .dout(n13115));
  jand g12834(.dina(n13104), .dinb(n305), .dout(n13116));
  jand g12835(.dina(n13116), .dinb(n13109), .dout(n13117));
  jor  g12836(.dina(n13117), .dinb(n13115), .dout(n13118));
  jand g12837(.dina(n13118), .dinb(n13111), .dout(n13119));
  jor  g12838(.dina(n13119), .dinb(n290), .dout(n13120));
  jand g12839(.dina(n13119), .dinb(n290), .dout(n13121));
  jnot g12840(.din(n12607), .dout(n13122));
  jand g12841(.dina(asqrt[15] ), .dinb(n13122), .dout(n13123));
  jand g12842(.dina(n13123), .dinb(n12612), .dout(n13124));
  jor  g12843(.dina(n13124), .dinb(n12611), .dout(n13125));
  jand g12844(.dina(n13123), .dinb(n12613), .dout(n13126));
  jnot g12845(.din(n13126), .dout(n13127));
  jand g12846(.dina(n13127), .dinb(n13125), .dout(n13128));
  jnot g12847(.din(n13128), .dout(n13129));
  jor  g12848(.dina(n13129), .dinb(n13121), .dout(n13130));
  jand g12849(.dina(n13130), .dinb(n13120), .dout(n13131));
  jor  g12850(.dina(n13131), .dinb(n223), .dout(n13132));
  jand g12851(.dina(n13120), .dinb(n223), .dout(n13133));
  jand g12852(.dina(n13133), .dinb(n13130), .dout(n13134));
  jnot g12853(.din(n12615), .dout(n13135));
  jand g12854(.dina(asqrt[15] ), .dinb(n13135), .dout(n13136));
  jand g12855(.dina(n13136), .dinb(n12622), .dout(n13137));
  jor  g12856(.dina(n13137), .dinb(n12620), .dout(n13138));
  jand g12857(.dina(n13136), .dinb(n12623), .dout(n13139));
  jnot g12858(.din(n13139), .dout(n13140));
  jand g12859(.dina(n13140), .dinb(n13138), .dout(n13141));
  jnot g12860(.din(n13141), .dout(n13142));
  jor  g12861(.dina(n13142), .dinb(n13134), .dout(n13143));
  jand g12862(.dina(n13143), .dinb(n13132), .dout(n13144));
  jor  g12863(.dina(n13144), .dinb(n199), .dout(n13145));
  jand g12864(.dina(n13144), .dinb(n199), .dout(n13146));
  jxor g12865(.dina(n12624), .dinb(n223), .dout(n13147));
  jor  g12866(.dina(n13147), .dinb(n12675), .dout(n13148));
  jxor g12867(.dina(n13148), .dinb(n12635), .dout(n13149));
  jor  g12868(.dina(n13149), .dinb(n13146), .dout(n13150));
  jand g12869(.dina(n13150), .dinb(n13145), .dout(n13151));
  jnot g12870(.din(n12640), .dout(n13152));
  jor  g12871(.dina(n13152), .dinb(n12638), .dout(n13153));
  jor  g12872(.dina(n13153), .dinb(n12675), .dout(n13154));
  jxor g12873(.dina(n13154), .dinb(n12649), .dout(n13155));
  jand g12874(.dina(asqrt[15] ), .dinb(n12663), .dout(n13156));
  jand g12875(.dina(n13156), .dinb(n12651), .dout(n13157));
  jor  g12876(.dina(n13157), .dinb(n12698), .dout(n13158));
  jor  g12877(.dina(n13158), .dinb(n13155), .dout(n13159));
  jor  g12878(.dina(n13159), .dinb(n13151), .dout(n13160));
  jand g12879(.dina(n13160), .dinb(n194), .dout(n13161));
  jand g12880(.dina(n13155), .dinb(n13151), .dout(n13162));
  jor  g12881(.dina(n13156), .dinb(n12651), .dout(n13163));
  jand g12882(.dina(n12663), .dinb(n12651), .dout(n13164));
  jor  g12883(.dina(n13164), .dinb(n194), .dout(n13165));
  jnot g12884(.din(n13165), .dout(n13166));
  jand g12885(.dina(n13166), .dinb(n13163), .dout(n13167));
  jor  g12886(.dina(n13167), .dinb(n13162), .dout(n13170));
  jor  g12887(.dina(n13170), .dinb(n13161), .dout(asqrt[14] ));
  jxor g12888(.dina(n13008), .dinb(n1641), .dout(n13172));
  jand g12889(.dina(n13172), .dinb(asqrt[14] ), .dout(n13173));
  jxor g12890(.dina(n13173), .dinb(n12679), .dout(n13174));
  jnot g12891(.din(n13174), .dout(n13175));
  jand g12892(.dina(asqrt[14] ), .dinb(a[28] ), .dout(n13176));
  jnot g12893(.din(a[26] ), .dout(n13177));
  jnot g12894(.din(a[27] ), .dout(n13178));
  jand g12895(.dina(n12681), .dinb(n13178), .dout(n13179));
  jand g12896(.dina(n13179), .dinb(n13177), .dout(n13180));
  jor  g12897(.dina(n13180), .dinb(n13176), .dout(n13181));
  jand g12898(.dina(n13181), .dinb(asqrt[15] ), .dout(n13182));
  jand g12899(.dina(asqrt[14] ), .dinb(n12681), .dout(n13183));
  jxor g12900(.dina(n13183), .dinb(n12682), .dout(n13184));
  jor  g12901(.dina(n13181), .dinb(asqrt[15] ), .dout(n13185));
  jand g12902(.dina(n13185), .dinb(n13184), .dout(n13186));
  jor  g12903(.dina(n13186), .dinb(n13182), .dout(n13187));
  jand g12904(.dina(n13187), .dinb(asqrt[16] ), .dout(n13188));
  jor  g12905(.dina(n13182), .dinb(asqrt[16] ), .dout(n13189));
  jor  g12906(.dina(n13189), .dinb(n13186), .dout(n13190));
  jand g12907(.dina(n13183), .dinb(n12682), .dout(n13191));
  jnot g12908(.din(n13161), .dout(n13192));
  jnot g12909(.din(n13162), .dout(n13193));
  jnot g12910(.din(n13167), .dout(n13194));
  jand g12911(.dina(n13194), .dinb(asqrt[15] ), .dout(n13195));
  jand g12912(.dina(n13195), .dinb(n13193), .dout(n13196));
  jand g12913(.dina(n13196), .dinb(n13192), .dout(n13197));
  jor  g12914(.dina(n13197), .dinb(n13191), .dout(n13198));
  jxor g12915(.dina(n13198), .dinb(n12148), .dout(n13199));
  jand g12916(.dina(n13199), .dinb(n13190), .dout(n13200));
  jor  g12917(.dina(n13200), .dinb(n13188), .dout(n13201));
  jand g12918(.dina(n13201), .dinb(asqrt[17] ), .dout(n13202));
  jor  g12919(.dina(n13201), .dinb(asqrt[17] ), .dout(n13203));
  jxor g12920(.dina(n12686), .dinb(n12670), .dout(n13204));
  jand g12921(.dina(n13204), .dinb(asqrt[14] ), .dout(n13205));
  jxor g12922(.dina(n13205), .dinb(n12689), .dout(n13206));
  jnot g12923(.din(n13206), .dout(n13207));
  jand g12924(.dina(n13207), .dinb(n13203), .dout(n13208));
  jor  g12925(.dina(n13208), .dinb(n13202), .dout(n13209));
  jand g12926(.dina(n13209), .dinb(asqrt[18] ), .dout(n13210));
  jnot g12927(.din(n12695), .dout(n13211));
  jand g12928(.dina(n13211), .dinb(n12693), .dout(n13212));
  jand g12929(.dina(n13212), .dinb(asqrt[14] ), .dout(n13213));
  jxor g12930(.dina(n13213), .dinb(n12703), .dout(n13214));
  jnot g12931(.din(n13214), .dout(n13215));
  jor  g12932(.dina(n13202), .dinb(asqrt[18] ), .dout(n13216));
  jor  g12933(.dina(n13216), .dinb(n13208), .dout(n13217));
  jand g12934(.dina(n13217), .dinb(n13215), .dout(n13218));
  jor  g12935(.dina(n13218), .dinb(n13210), .dout(n13219));
  jand g12936(.dina(n13219), .dinb(asqrt[19] ), .dout(n13220));
  jor  g12937(.dina(n13219), .dinb(asqrt[19] ), .dout(n13221));
  jnot g12938(.din(n12710), .dout(n13222));
  jxor g12939(.dina(n12705), .dinb(n11657), .dout(n13223));
  jand g12940(.dina(n13223), .dinb(asqrt[14] ), .dout(n13224));
  jxor g12941(.dina(n13224), .dinb(n13222), .dout(n13225));
  jand g12942(.dina(n13225), .dinb(n13221), .dout(n13226));
  jor  g12943(.dina(n13226), .dinb(n13220), .dout(n13227));
  jand g12944(.dina(n13227), .dinb(asqrt[20] ), .dout(n13228));
  jor  g12945(.dina(n13220), .dinb(asqrt[20] ), .dout(n13229));
  jor  g12946(.dina(n13229), .dinb(n13226), .dout(n13230));
  jnot g12947(.din(n12717), .dout(n13231));
  jnot g12948(.din(n12719), .dout(n13232));
  jand g12949(.dina(asqrt[14] ), .dinb(n12713), .dout(n13233));
  jand g12950(.dina(n13233), .dinb(n13232), .dout(n13234));
  jor  g12951(.dina(n13234), .dinb(n13231), .dout(n13235));
  jnot g12952(.din(n12720), .dout(n13236));
  jand g12953(.dina(n13233), .dinb(n13236), .dout(n13237));
  jnot g12954(.din(n13237), .dout(n13238));
  jand g12955(.dina(n13238), .dinb(n13235), .dout(n13239));
  jand g12956(.dina(n13239), .dinb(n13230), .dout(n13240));
  jor  g12957(.dina(n13240), .dinb(n13228), .dout(n13241));
  jand g12958(.dina(n13241), .dinb(asqrt[21] ), .dout(n13242));
  jor  g12959(.dina(n13241), .dinb(asqrt[21] ), .dout(n13243));
  jxor g12960(.dina(n12721), .dinb(n10696), .dout(n13244));
  jand g12961(.dina(n13244), .dinb(asqrt[14] ), .dout(n13245));
  jxor g12962(.dina(n13245), .dinb(n12726), .dout(n13246));
  jand g12963(.dina(n13246), .dinb(n13243), .dout(n13247));
  jor  g12964(.dina(n13247), .dinb(n13242), .dout(n13248));
  jand g12965(.dina(n13248), .dinb(asqrt[22] ), .dout(n13249));
  jnot g12966(.din(n12732), .dout(n13250));
  jand g12967(.dina(n13250), .dinb(n12730), .dout(n13251));
  jand g12968(.dina(n13251), .dinb(asqrt[14] ), .dout(n13252));
  jxor g12969(.dina(n13252), .dinb(n12741), .dout(n13253));
  jnot g12970(.din(n13253), .dout(n13254));
  jor  g12971(.dina(n13242), .dinb(asqrt[22] ), .dout(n13255));
  jor  g12972(.dina(n13255), .dinb(n13247), .dout(n13256));
  jand g12973(.dina(n13256), .dinb(n13254), .dout(n13257));
  jor  g12974(.dina(n13257), .dinb(n13249), .dout(n13258));
  jand g12975(.dina(n13258), .dinb(asqrt[23] ), .dout(n13259));
  jor  g12976(.dina(n13258), .dinb(asqrt[23] ), .dout(n13260));
  jxor g12977(.dina(n12743), .dinb(n9769), .dout(n13261));
  jand g12978(.dina(n13261), .dinb(asqrt[14] ), .dout(n13262));
  jxor g12979(.dina(n13262), .dinb(n12749), .dout(n13263));
  jand g12980(.dina(n13263), .dinb(n13260), .dout(n13264));
  jor  g12981(.dina(n13264), .dinb(n13259), .dout(n13265));
  jand g12982(.dina(n13265), .dinb(asqrt[24] ), .dout(n13266));
  jor  g12983(.dina(n13259), .dinb(asqrt[24] ), .dout(n13267));
  jor  g12984(.dina(n13267), .dinb(n13264), .dout(n13268));
  jnot g12985(.din(n12757), .dout(n13269));
  jnot g12986(.din(n12759), .dout(n13270));
  jand g12987(.dina(asqrt[14] ), .dinb(n12753), .dout(n13271));
  jand g12988(.dina(n13271), .dinb(n13270), .dout(n13272));
  jor  g12989(.dina(n13272), .dinb(n13269), .dout(n13273));
  jnot g12990(.din(n12760), .dout(n13274));
  jand g12991(.dina(n13271), .dinb(n13274), .dout(n13275));
  jnot g12992(.din(n13275), .dout(n13276));
  jand g12993(.dina(n13276), .dinb(n13273), .dout(n13277));
  jand g12994(.dina(n13277), .dinb(n13268), .dout(n13278));
  jor  g12995(.dina(n13278), .dinb(n13266), .dout(n13279));
  jand g12996(.dina(n13279), .dinb(asqrt[25] ), .dout(n13280));
  jxor g12997(.dina(n12761), .dinb(n8893), .dout(n13281));
  jand g12998(.dina(n13281), .dinb(asqrt[14] ), .dout(n13282));
  jxor g12999(.dina(n13282), .dinb(n12768), .dout(n13283));
  jnot g13000(.din(n13283), .dout(n13284));
  jor  g13001(.dina(n13279), .dinb(asqrt[25] ), .dout(n13285));
  jand g13002(.dina(n13285), .dinb(n13284), .dout(n13286));
  jor  g13003(.dina(n13286), .dinb(n13280), .dout(n13287));
  jand g13004(.dina(n13287), .dinb(asqrt[26] ), .dout(n13288));
  jnot g13005(.din(n12773), .dout(n13289));
  jand g13006(.dina(n13289), .dinb(n12771), .dout(n13290));
  jand g13007(.dina(n13290), .dinb(asqrt[14] ), .dout(n13291));
  jxor g13008(.dina(n13291), .dinb(n12781), .dout(n13292));
  jnot g13009(.din(n13292), .dout(n13293));
  jor  g13010(.dina(n13280), .dinb(asqrt[26] ), .dout(n13294));
  jor  g13011(.dina(n13294), .dinb(n13286), .dout(n13295));
  jand g13012(.dina(n13295), .dinb(n13293), .dout(n13296));
  jor  g13013(.dina(n13296), .dinb(n13288), .dout(n13297));
  jand g13014(.dina(n13297), .dinb(asqrt[27] ), .dout(n13298));
  jor  g13015(.dina(n13297), .dinb(asqrt[27] ), .dout(n13299));
  jnot g13016(.din(n12787), .dout(n13300));
  jnot g13017(.din(n12788), .dout(n13301));
  jand g13018(.dina(asqrt[14] ), .dinb(n12784), .dout(n13302));
  jand g13019(.dina(n13302), .dinb(n13301), .dout(n13303));
  jor  g13020(.dina(n13303), .dinb(n13300), .dout(n13304));
  jnot g13021(.din(n12789), .dout(n13305));
  jand g13022(.dina(n13302), .dinb(n13305), .dout(n13306));
  jnot g13023(.din(n13306), .dout(n13307));
  jand g13024(.dina(n13307), .dinb(n13304), .dout(n13308));
  jand g13025(.dina(n13308), .dinb(n13299), .dout(n13309));
  jor  g13026(.dina(n13309), .dinb(n13298), .dout(n13310));
  jand g13027(.dina(n13310), .dinb(asqrt[28] ), .dout(n13311));
  jor  g13028(.dina(n13298), .dinb(asqrt[28] ), .dout(n13312));
  jor  g13029(.dina(n13312), .dinb(n13309), .dout(n13313));
  jnot g13030(.din(n12795), .dout(n13314));
  jnot g13031(.din(n12797), .dout(n13315));
  jand g13032(.dina(asqrt[14] ), .dinb(n12791), .dout(n13316));
  jand g13033(.dina(n13316), .dinb(n13315), .dout(n13317));
  jor  g13034(.dina(n13317), .dinb(n13314), .dout(n13318));
  jnot g13035(.din(n12798), .dout(n13319));
  jand g13036(.dina(n13316), .dinb(n13319), .dout(n13320));
  jnot g13037(.din(n13320), .dout(n13321));
  jand g13038(.dina(n13321), .dinb(n13318), .dout(n13322));
  jand g13039(.dina(n13322), .dinb(n13313), .dout(n13323));
  jor  g13040(.dina(n13323), .dinb(n13311), .dout(n13324));
  jand g13041(.dina(n13324), .dinb(asqrt[29] ), .dout(n13325));
  jxor g13042(.dina(n12799), .dinb(n7260), .dout(n13326));
  jand g13043(.dina(n13326), .dinb(asqrt[14] ), .dout(n13327));
  jxor g13044(.dina(n13327), .dinb(n12809), .dout(n13328));
  jnot g13045(.din(n13328), .dout(n13329));
  jor  g13046(.dina(n13324), .dinb(asqrt[29] ), .dout(n13330));
  jand g13047(.dina(n13330), .dinb(n13329), .dout(n13331));
  jor  g13048(.dina(n13331), .dinb(n13325), .dout(n13332));
  jand g13049(.dina(n13332), .dinb(asqrt[30] ), .dout(n13333));
  jnot g13050(.din(n12814), .dout(n13334));
  jand g13051(.dina(n13334), .dinb(n12812), .dout(n13335));
  jand g13052(.dina(n13335), .dinb(asqrt[14] ), .dout(n13336));
  jxor g13053(.dina(n13336), .dinb(n12822), .dout(n13337));
  jnot g13054(.din(n13337), .dout(n13338));
  jor  g13055(.dina(n13325), .dinb(asqrt[30] ), .dout(n13339));
  jor  g13056(.dina(n13339), .dinb(n13331), .dout(n13340));
  jand g13057(.dina(n13340), .dinb(n13338), .dout(n13341));
  jor  g13058(.dina(n13341), .dinb(n13333), .dout(n13342));
  jand g13059(.dina(n13342), .dinb(asqrt[31] ), .dout(n13343));
  jor  g13060(.dina(n13342), .dinb(asqrt[31] ), .dout(n13344));
  jnot g13061(.din(n12828), .dout(n13345));
  jnot g13062(.din(n12829), .dout(n13346));
  jand g13063(.dina(asqrt[14] ), .dinb(n12825), .dout(n13347));
  jand g13064(.dina(n13347), .dinb(n13346), .dout(n13348));
  jor  g13065(.dina(n13348), .dinb(n13345), .dout(n13349));
  jnot g13066(.din(n12830), .dout(n13350));
  jand g13067(.dina(n13347), .dinb(n13350), .dout(n13351));
  jnot g13068(.din(n13351), .dout(n13352));
  jand g13069(.dina(n13352), .dinb(n13349), .dout(n13353));
  jand g13070(.dina(n13353), .dinb(n13344), .dout(n13354));
  jor  g13071(.dina(n13354), .dinb(n13343), .dout(n13355));
  jand g13072(.dina(n13355), .dinb(asqrt[32] ), .dout(n13356));
  jor  g13073(.dina(n13343), .dinb(asqrt[32] ), .dout(n13357));
  jor  g13074(.dina(n13357), .dinb(n13354), .dout(n13358));
  jnot g13075(.din(n12836), .dout(n13359));
  jnot g13076(.din(n12838), .dout(n13360));
  jand g13077(.dina(asqrt[14] ), .dinb(n12832), .dout(n13361));
  jand g13078(.dina(n13361), .dinb(n13360), .dout(n13362));
  jor  g13079(.dina(n13362), .dinb(n13359), .dout(n13363));
  jnot g13080(.din(n12839), .dout(n13364));
  jand g13081(.dina(n13361), .dinb(n13364), .dout(n13365));
  jnot g13082(.din(n13365), .dout(n13366));
  jand g13083(.dina(n13366), .dinb(n13363), .dout(n13367));
  jand g13084(.dina(n13367), .dinb(n13358), .dout(n13368));
  jor  g13085(.dina(n13368), .dinb(n13356), .dout(n13369));
  jand g13086(.dina(n13369), .dinb(asqrt[33] ), .dout(n13370));
  jxor g13087(.dina(n12840), .dinb(n5788), .dout(n13371));
  jand g13088(.dina(n13371), .dinb(asqrt[14] ), .dout(n13372));
  jxor g13089(.dina(n13372), .dinb(n12850), .dout(n13373));
  jnot g13090(.din(n13373), .dout(n13374));
  jor  g13091(.dina(n13369), .dinb(asqrt[33] ), .dout(n13375));
  jand g13092(.dina(n13375), .dinb(n13374), .dout(n13376));
  jor  g13093(.dina(n13376), .dinb(n13370), .dout(n13377));
  jand g13094(.dina(n13377), .dinb(asqrt[34] ), .dout(n13378));
  jnot g13095(.din(n12855), .dout(n13379));
  jand g13096(.dina(n13379), .dinb(n12853), .dout(n13380));
  jand g13097(.dina(n13380), .dinb(asqrt[14] ), .dout(n13381));
  jxor g13098(.dina(n13381), .dinb(n12863), .dout(n13382));
  jnot g13099(.din(n13382), .dout(n13383));
  jor  g13100(.dina(n13370), .dinb(asqrt[34] ), .dout(n13384));
  jor  g13101(.dina(n13384), .dinb(n13376), .dout(n13385));
  jand g13102(.dina(n13385), .dinb(n13383), .dout(n13386));
  jor  g13103(.dina(n13386), .dinb(n13378), .dout(n13387));
  jand g13104(.dina(n13387), .dinb(asqrt[35] ), .dout(n13388));
  jor  g13105(.dina(n13387), .dinb(asqrt[35] ), .dout(n13389));
  jnot g13106(.din(n12869), .dout(n13390));
  jnot g13107(.din(n12870), .dout(n13391));
  jand g13108(.dina(asqrt[14] ), .dinb(n12866), .dout(n13392));
  jand g13109(.dina(n13392), .dinb(n13391), .dout(n13393));
  jor  g13110(.dina(n13393), .dinb(n13390), .dout(n13394));
  jnot g13111(.din(n12871), .dout(n13395));
  jand g13112(.dina(n13392), .dinb(n13395), .dout(n13396));
  jnot g13113(.din(n13396), .dout(n13397));
  jand g13114(.dina(n13397), .dinb(n13394), .dout(n13398));
  jand g13115(.dina(n13398), .dinb(n13389), .dout(n13399));
  jor  g13116(.dina(n13399), .dinb(n13388), .dout(n13400));
  jand g13117(.dina(n13400), .dinb(asqrt[36] ), .dout(n13401));
  jor  g13118(.dina(n13388), .dinb(asqrt[36] ), .dout(n13402));
  jor  g13119(.dina(n13402), .dinb(n13399), .dout(n13403));
  jnot g13120(.din(n12877), .dout(n13404));
  jnot g13121(.din(n12879), .dout(n13405));
  jand g13122(.dina(asqrt[14] ), .dinb(n12873), .dout(n13406));
  jand g13123(.dina(n13406), .dinb(n13405), .dout(n13407));
  jor  g13124(.dina(n13407), .dinb(n13404), .dout(n13408));
  jnot g13125(.din(n12880), .dout(n13409));
  jand g13126(.dina(n13406), .dinb(n13409), .dout(n13410));
  jnot g13127(.din(n13410), .dout(n13411));
  jand g13128(.dina(n13411), .dinb(n13408), .dout(n13412));
  jand g13129(.dina(n13412), .dinb(n13403), .dout(n13413));
  jor  g13130(.dina(n13413), .dinb(n13401), .dout(n13414));
  jand g13131(.dina(n13414), .dinb(asqrt[37] ), .dout(n13415));
  jxor g13132(.dina(n12881), .dinb(n4494), .dout(n13416));
  jand g13133(.dina(n13416), .dinb(asqrt[14] ), .dout(n13417));
  jxor g13134(.dina(n13417), .dinb(n12891), .dout(n13418));
  jnot g13135(.din(n13418), .dout(n13419));
  jor  g13136(.dina(n13414), .dinb(asqrt[37] ), .dout(n13420));
  jand g13137(.dina(n13420), .dinb(n13419), .dout(n13421));
  jor  g13138(.dina(n13421), .dinb(n13415), .dout(n13422));
  jand g13139(.dina(n13422), .dinb(asqrt[38] ), .dout(n13423));
  jnot g13140(.din(n12896), .dout(n13424));
  jand g13141(.dina(n13424), .dinb(n12894), .dout(n13425));
  jand g13142(.dina(n13425), .dinb(asqrt[14] ), .dout(n13426));
  jxor g13143(.dina(n13426), .dinb(n12904), .dout(n13427));
  jnot g13144(.din(n13427), .dout(n13428));
  jor  g13145(.dina(n13415), .dinb(asqrt[38] ), .dout(n13429));
  jor  g13146(.dina(n13429), .dinb(n13421), .dout(n13430));
  jand g13147(.dina(n13430), .dinb(n13428), .dout(n13431));
  jor  g13148(.dina(n13431), .dinb(n13423), .dout(n13432));
  jand g13149(.dina(n13432), .dinb(asqrt[39] ), .dout(n13433));
  jor  g13150(.dina(n13432), .dinb(asqrt[39] ), .dout(n13434));
  jnot g13151(.din(n12910), .dout(n13435));
  jnot g13152(.din(n12911), .dout(n13436));
  jand g13153(.dina(asqrt[14] ), .dinb(n12907), .dout(n13437));
  jand g13154(.dina(n13437), .dinb(n13436), .dout(n13438));
  jor  g13155(.dina(n13438), .dinb(n13435), .dout(n13439));
  jnot g13156(.din(n12912), .dout(n13440));
  jand g13157(.dina(n13437), .dinb(n13440), .dout(n13441));
  jnot g13158(.din(n13441), .dout(n13442));
  jand g13159(.dina(n13442), .dinb(n13439), .dout(n13443));
  jand g13160(.dina(n13443), .dinb(n13434), .dout(n13444));
  jor  g13161(.dina(n13444), .dinb(n13433), .dout(n13445));
  jand g13162(.dina(n13445), .dinb(asqrt[40] ), .dout(n13446));
  jor  g13163(.dina(n13433), .dinb(asqrt[40] ), .dout(n13447));
  jor  g13164(.dina(n13447), .dinb(n13444), .dout(n13448));
  jnot g13165(.din(n12918), .dout(n13449));
  jnot g13166(.din(n12920), .dout(n13450));
  jand g13167(.dina(asqrt[14] ), .dinb(n12914), .dout(n13451));
  jand g13168(.dina(n13451), .dinb(n13450), .dout(n13452));
  jor  g13169(.dina(n13452), .dinb(n13449), .dout(n13453));
  jnot g13170(.din(n12921), .dout(n13454));
  jand g13171(.dina(n13451), .dinb(n13454), .dout(n13455));
  jnot g13172(.din(n13455), .dout(n13456));
  jand g13173(.dina(n13456), .dinb(n13453), .dout(n13457));
  jand g13174(.dina(n13457), .dinb(n13448), .dout(n13458));
  jor  g13175(.dina(n13458), .dinb(n13446), .dout(n13459));
  jand g13176(.dina(n13459), .dinb(asqrt[41] ), .dout(n13460));
  jxor g13177(.dina(n12922), .dinb(n3371), .dout(n13461));
  jand g13178(.dina(n13461), .dinb(asqrt[14] ), .dout(n13462));
  jxor g13179(.dina(n13462), .dinb(n12932), .dout(n13463));
  jnot g13180(.din(n13463), .dout(n13464));
  jor  g13181(.dina(n13459), .dinb(asqrt[41] ), .dout(n13465));
  jand g13182(.dina(n13465), .dinb(n13464), .dout(n13466));
  jor  g13183(.dina(n13466), .dinb(n13460), .dout(n13467));
  jand g13184(.dina(n13467), .dinb(asqrt[42] ), .dout(n13468));
  jnot g13185(.din(n12937), .dout(n13469));
  jand g13186(.dina(n13469), .dinb(n12935), .dout(n13470));
  jand g13187(.dina(n13470), .dinb(asqrt[14] ), .dout(n13471));
  jxor g13188(.dina(n13471), .dinb(n12945), .dout(n13472));
  jnot g13189(.din(n13472), .dout(n13473));
  jor  g13190(.dina(n13460), .dinb(asqrt[42] ), .dout(n13474));
  jor  g13191(.dina(n13474), .dinb(n13466), .dout(n13475));
  jand g13192(.dina(n13475), .dinb(n13473), .dout(n13476));
  jor  g13193(.dina(n13476), .dinb(n13468), .dout(n13477));
  jand g13194(.dina(n13477), .dinb(asqrt[43] ), .dout(n13478));
  jor  g13195(.dina(n13477), .dinb(asqrt[43] ), .dout(n13479));
  jnot g13196(.din(n12951), .dout(n13480));
  jnot g13197(.din(n12952), .dout(n13481));
  jand g13198(.dina(asqrt[14] ), .dinb(n12948), .dout(n13482));
  jand g13199(.dina(n13482), .dinb(n13481), .dout(n13483));
  jor  g13200(.dina(n13483), .dinb(n13480), .dout(n13484));
  jnot g13201(.din(n12953), .dout(n13485));
  jand g13202(.dina(n13482), .dinb(n13485), .dout(n13486));
  jnot g13203(.din(n13486), .dout(n13487));
  jand g13204(.dina(n13487), .dinb(n13484), .dout(n13488));
  jand g13205(.dina(n13488), .dinb(n13479), .dout(n13489));
  jor  g13206(.dina(n13489), .dinb(n13478), .dout(n13490));
  jand g13207(.dina(n13490), .dinb(asqrt[44] ), .dout(n13491));
  jor  g13208(.dina(n13478), .dinb(asqrt[44] ), .dout(n13492));
  jor  g13209(.dina(n13492), .dinb(n13489), .dout(n13493));
  jnot g13210(.din(n12959), .dout(n13494));
  jnot g13211(.din(n12961), .dout(n13495));
  jand g13212(.dina(asqrt[14] ), .dinb(n12955), .dout(n13496));
  jand g13213(.dina(n13496), .dinb(n13495), .dout(n13497));
  jor  g13214(.dina(n13497), .dinb(n13494), .dout(n13498));
  jnot g13215(.din(n12962), .dout(n13499));
  jand g13216(.dina(n13496), .dinb(n13499), .dout(n13500));
  jnot g13217(.din(n13500), .dout(n13501));
  jand g13218(.dina(n13501), .dinb(n13498), .dout(n13502));
  jand g13219(.dina(n13502), .dinb(n13493), .dout(n13503));
  jor  g13220(.dina(n13503), .dinb(n13491), .dout(n13504));
  jand g13221(.dina(n13504), .dinb(asqrt[45] ), .dout(n13505));
  jxor g13222(.dina(n12963), .dinb(n2420), .dout(n13506));
  jand g13223(.dina(n13506), .dinb(asqrt[14] ), .dout(n13507));
  jxor g13224(.dina(n13507), .dinb(n12973), .dout(n13508));
  jnot g13225(.din(n13508), .dout(n13509));
  jor  g13226(.dina(n13504), .dinb(asqrt[45] ), .dout(n13510));
  jand g13227(.dina(n13510), .dinb(n13509), .dout(n13511));
  jor  g13228(.dina(n13511), .dinb(n13505), .dout(n13512));
  jand g13229(.dina(n13512), .dinb(asqrt[46] ), .dout(n13513));
  jnot g13230(.din(n12978), .dout(n13514));
  jand g13231(.dina(n13514), .dinb(n12976), .dout(n13515));
  jand g13232(.dina(n13515), .dinb(asqrt[14] ), .dout(n13516));
  jxor g13233(.dina(n13516), .dinb(n12986), .dout(n13517));
  jnot g13234(.din(n13517), .dout(n13518));
  jor  g13235(.dina(n13505), .dinb(asqrt[46] ), .dout(n13519));
  jor  g13236(.dina(n13519), .dinb(n13511), .dout(n13520));
  jand g13237(.dina(n13520), .dinb(n13518), .dout(n13521));
  jor  g13238(.dina(n13521), .dinb(n13513), .dout(n13522));
  jand g13239(.dina(n13522), .dinb(asqrt[47] ), .dout(n13523));
  jor  g13240(.dina(n13522), .dinb(asqrt[47] ), .dout(n13524));
  jnot g13241(.din(n12992), .dout(n13525));
  jnot g13242(.din(n12993), .dout(n13526));
  jand g13243(.dina(asqrt[14] ), .dinb(n12989), .dout(n13527));
  jand g13244(.dina(n13527), .dinb(n13526), .dout(n13528));
  jor  g13245(.dina(n13528), .dinb(n13525), .dout(n13529));
  jnot g13246(.din(n12994), .dout(n13530));
  jand g13247(.dina(n13527), .dinb(n13530), .dout(n13531));
  jnot g13248(.din(n13531), .dout(n13532));
  jand g13249(.dina(n13532), .dinb(n13529), .dout(n13533));
  jand g13250(.dina(n13533), .dinb(n13524), .dout(n13534));
  jor  g13251(.dina(n13534), .dinb(n13523), .dout(n13535));
  jand g13252(.dina(n13535), .dinb(asqrt[48] ), .dout(n13536));
  jnot g13253(.din(n12998), .dout(n13537));
  jand g13254(.dina(n13537), .dinb(n12996), .dout(n13538));
  jand g13255(.dina(n13538), .dinb(asqrt[14] ), .dout(n13539));
  jxor g13256(.dina(n13539), .dinb(n13006), .dout(n13540));
  jnot g13257(.din(n13540), .dout(n13541));
  jor  g13258(.dina(n13523), .dinb(asqrt[48] ), .dout(n13542));
  jor  g13259(.dina(n13542), .dinb(n13534), .dout(n13543));
  jand g13260(.dina(n13543), .dinb(n13541), .dout(n13544));
  jor  g13261(.dina(n13544), .dinb(n13536), .dout(n13545));
  jand g13262(.dina(n13545), .dinb(asqrt[49] ), .dout(n13546));
  jor  g13263(.dina(n13545), .dinb(asqrt[49] ), .dout(n13547));
  jand g13264(.dina(n13547), .dinb(n13175), .dout(n13548));
  jor  g13265(.dina(n13548), .dinb(n13546), .dout(n13549));
  jand g13266(.dina(n13549), .dinb(asqrt[50] ), .dout(n13550));
  jor  g13267(.dina(n13546), .dinb(asqrt[50] ), .dout(n13551));
  jor  g13268(.dina(n13551), .dinb(n13548), .dout(n13552));
  jnot g13269(.din(n13017), .dout(n13553));
  jnot g13270(.din(n13019), .dout(n13554));
  jand g13271(.dina(asqrt[14] ), .dinb(n13013), .dout(n13555));
  jand g13272(.dina(n13555), .dinb(n13554), .dout(n13556));
  jor  g13273(.dina(n13556), .dinb(n13553), .dout(n13557));
  jnot g13274(.din(n13020), .dout(n13558));
  jand g13275(.dina(n13555), .dinb(n13558), .dout(n13559));
  jnot g13276(.din(n13559), .dout(n13560));
  jand g13277(.dina(n13560), .dinb(n13557), .dout(n13561));
  jand g13278(.dina(n13561), .dinb(n13552), .dout(n13562));
  jor  g13279(.dina(n13562), .dinb(n13550), .dout(n13563));
  jand g13280(.dina(n13563), .dinb(asqrt[51] ), .dout(n13564));
  jor  g13281(.dina(n13563), .dinb(asqrt[51] ), .dout(n13565));
  jnot g13282(.din(n13025), .dout(n13566));
  jnot g13283(.din(n13026), .dout(n13567));
  jand g13284(.dina(asqrt[14] ), .dinb(n13022), .dout(n13568));
  jand g13285(.dina(n13568), .dinb(n13567), .dout(n13569));
  jor  g13286(.dina(n13569), .dinb(n13566), .dout(n13570));
  jnot g13287(.din(n13027), .dout(n13571));
  jand g13288(.dina(n13568), .dinb(n13571), .dout(n13572));
  jnot g13289(.din(n13572), .dout(n13573));
  jand g13290(.dina(n13573), .dinb(n13570), .dout(n13574));
  jand g13291(.dina(n13574), .dinb(n13565), .dout(n13575));
  jor  g13292(.dina(n13575), .dinb(n13564), .dout(n13576));
  jand g13293(.dina(n13576), .dinb(asqrt[52] ), .dout(n13577));
  jor  g13294(.dina(n13564), .dinb(asqrt[52] ), .dout(n13578));
  jor  g13295(.dina(n13578), .dinb(n13575), .dout(n13579));
  jnot g13296(.din(n13033), .dout(n13580));
  jnot g13297(.din(n13035), .dout(n13581));
  jand g13298(.dina(asqrt[14] ), .dinb(n13029), .dout(n13582));
  jand g13299(.dina(n13582), .dinb(n13581), .dout(n13583));
  jor  g13300(.dina(n13583), .dinb(n13580), .dout(n13584));
  jnot g13301(.din(n13036), .dout(n13585));
  jand g13302(.dina(n13582), .dinb(n13585), .dout(n13586));
  jnot g13303(.din(n13586), .dout(n13587));
  jand g13304(.dina(n13587), .dinb(n13584), .dout(n13588));
  jand g13305(.dina(n13588), .dinb(n13579), .dout(n13589));
  jor  g13306(.dina(n13589), .dinb(n13577), .dout(n13590));
  jand g13307(.dina(n13590), .dinb(asqrt[53] ), .dout(n13591));
  jxor g13308(.dina(n13037), .dinb(n1034), .dout(n13592));
  jand g13309(.dina(n13592), .dinb(asqrt[14] ), .dout(n13593));
  jxor g13310(.dina(n13593), .dinb(n13047), .dout(n13594));
  jnot g13311(.din(n13594), .dout(n13595));
  jor  g13312(.dina(n13590), .dinb(asqrt[53] ), .dout(n13596));
  jand g13313(.dina(n13596), .dinb(n13595), .dout(n13597));
  jor  g13314(.dina(n13597), .dinb(n13591), .dout(n13598));
  jand g13315(.dina(n13598), .dinb(asqrt[54] ), .dout(n13599));
  jnot g13316(.din(n13052), .dout(n13600));
  jand g13317(.dina(n13600), .dinb(n13050), .dout(n13601));
  jand g13318(.dina(n13601), .dinb(asqrt[14] ), .dout(n13602));
  jxor g13319(.dina(n13602), .dinb(n13060), .dout(n13603));
  jnot g13320(.din(n13603), .dout(n13604));
  jor  g13321(.dina(n13591), .dinb(asqrt[54] ), .dout(n13605));
  jor  g13322(.dina(n13605), .dinb(n13597), .dout(n13606));
  jand g13323(.dina(n13606), .dinb(n13604), .dout(n13607));
  jor  g13324(.dina(n13607), .dinb(n13599), .dout(n13608));
  jand g13325(.dina(n13608), .dinb(asqrt[55] ), .dout(n13609));
  jor  g13326(.dina(n13608), .dinb(asqrt[55] ), .dout(n13610));
  jnot g13327(.din(n13066), .dout(n13611));
  jnot g13328(.din(n13067), .dout(n13612));
  jand g13329(.dina(asqrt[14] ), .dinb(n13063), .dout(n13613));
  jand g13330(.dina(n13613), .dinb(n13612), .dout(n13614));
  jor  g13331(.dina(n13614), .dinb(n13611), .dout(n13615));
  jnot g13332(.din(n13068), .dout(n13616));
  jand g13333(.dina(n13613), .dinb(n13616), .dout(n13617));
  jnot g13334(.din(n13617), .dout(n13618));
  jand g13335(.dina(n13618), .dinb(n13615), .dout(n13619));
  jand g13336(.dina(n13619), .dinb(n13610), .dout(n13620));
  jor  g13337(.dina(n13620), .dinb(n13609), .dout(n13621));
  jand g13338(.dina(n13621), .dinb(asqrt[56] ), .dout(n13622));
  jor  g13339(.dina(n13609), .dinb(asqrt[56] ), .dout(n13623));
  jor  g13340(.dina(n13623), .dinb(n13620), .dout(n13624));
  jnot g13341(.din(n13074), .dout(n13625));
  jnot g13342(.din(n13076), .dout(n13626));
  jand g13343(.dina(asqrt[14] ), .dinb(n13070), .dout(n13627));
  jand g13344(.dina(n13627), .dinb(n13626), .dout(n13628));
  jor  g13345(.dina(n13628), .dinb(n13625), .dout(n13629));
  jnot g13346(.din(n13077), .dout(n13630));
  jand g13347(.dina(n13627), .dinb(n13630), .dout(n13631));
  jnot g13348(.din(n13631), .dout(n13632));
  jand g13349(.dina(n13632), .dinb(n13629), .dout(n13633));
  jand g13350(.dina(n13633), .dinb(n13624), .dout(n13634));
  jor  g13351(.dina(n13634), .dinb(n13622), .dout(n13635));
  jand g13352(.dina(n13635), .dinb(asqrt[57] ), .dout(n13636));
  jxor g13353(.dina(n13078), .dinb(n590), .dout(n13637));
  jand g13354(.dina(n13637), .dinb(asqrt[14] ), .dout(n13638));
  jxor g13355(.dina(n13638), .dinb(n13088), .dout(n13639));
  jnot g13356(.din(n13639), .dout(n13640));
  jor  g13357(.dina(n13635), .dinb(asqrt[57] ), .dout(n13641));
  jand g13358(.dina(n13641), .dinb(n13640), .dout(n13642));
  jor  g13359(.dina(n13642), .dinb(n13636), .dout(n13643));
  jand g13360(.dina(n13643), .dinb(asqrt[58] ), .dout(n13644));
  jnot g13361(.din(n13093), .dout(n13645));
  jand g13362(.dina(n13645), .dinb(n13091), .dout(n13646));
  jand g13363(.dina(n13646), .dinb(asqrt[14] ), .dout(n13647));
  jxor g13364(.dina(n13647), .dinb(n13101), .dout(n13648));
  jnot g13365(.din(n13648), .dout(n13649));
  jor  g13366(.dina(n13636), .dinb(asqrt[58] ), .dout(n13650));
  jor  g13367(.dina(n13650), .dinb(n13642), .dout(n13651));
  jand g13368(.dina(n13651), .dinb(n13649), .dout(n13652));
  jor  g13369(.dina(n13652), .dinb(n13644), .dout(n13653));
  jand g13370(.dina(n13653), .dinb(asqrt[59] ), .dout(n13654));
  jor  g13371(.dina(n13653), .dinb(asqrt[59] ), .dout(n13655));
  jnot g13372(.din(n13107), .dout(n13656));
  jnot g13373(.din(n13108), .dout(n13657));
  jand g13374(.dina(asqrt[14] ), .dinb(n13104), .dout(n13658));
  jand g13375(.dina(n13658), .dinb(n13657), .dout(n13659));
  jor  g13376(.dina(n13659), .dinb(n13656), .dout(n13660));
  jnot g13377(.din(n13109), .dout(n13661));
  jand g13378(.dina(n13658), .dinb(n13661), .dout(n13662));
  jnot g13379(.din(n13662), .dout(n13663));
  jand g13380(.dina(n13663), .dinb(n13660), .dout(n13664));
  jand g13381(.dina(n13664), .dinb(n13655), .dout(n13665));
  jor  g13382(.dina(n13665), .dinb(n13654), .dout(n13666));
  jand g13383(.dina(n13666), .dinb(asqrt[60] ), .dout(n13667));
  jor  g13384(.dina(n13654), .dinb(asqrt[60] ), .dout(n13668));
  jor  g13385(.dina(n13668), .dinb(n13665), .dout(n13669));
  jnot g13386(.din(n13115), .dout(n13670));
  jnot g13387(.din(n13117), .dout(n13671));
  jand g13388(.dina(asqrt[14] ), .dinb(n13111), .dout(n13672));
  jand g13389(.dina(n13672), .dinb(n13671), .dout(n13673));
  jor  g13390(.dina(n13673), .dinb(n13670), .dout(n13674));
  jnot g13391(.din(n13118), .dout(n13675));
  jand g13392(.dina(n13672), .dinb(n13675), .dout(n13676));
  jnot g13393(.din(n13676), .dout(n13677));
  jand g13394(.dina(n13677), .dinb(n13674), .dout(n13678));
  jand g13395(.dina(n13678), .dinb(n13669), .dout(n13679));
  jor  g13396(.dina(n13679), .dinb(n13667), .dout(n13680));
  jand g13397(.dina(n13680), .dinb(asqrt[61] ), .dout(n13681));
  jxor g13398(.dina(n13119), .dinb(n290), .dout(n13682));
  jand g13399(.dina(n13682), .dinb(asqrt[14] ), .dout(n13683));
  jxor g13400(.dina(n13683), .dinb(n13129), .dout(n13684));
  jnot g13401(.din(n13684), .dout(n13685));
  jor  g13402(.dina(n13680), .dinb(asqrt[61] ), .dout(n13686));
  jand g13403(.dina(n13686), .dinb(n13685), .dout(n13687));
  jor  g13404(.dina(n13687), .dinb(n13681), .dout(n13688));
  jand g13405(.dina(n13688), .dinb(asqrt[62] ), .dout(n13689));
  jnot g13406(.din(n13134), .dout(n13690));
  jand g13407(.dina(n13690), .dinb(n13132), .dout(n13691));
  jand g13408(.dina(n13691), .dinb(asqrt[14] ), .dout(n13692));
  jxor g13409(.dina(n13692), .dinb(n13142), .dout(n13693));
  jnot g13410(.din(n13693), .dout(n13694));
  jor  g13411(.dina(n13681), .dinb(asqrt[62] ), .dout(n13695));
  jor  g13412(.dina(n13695), .dinb(n13687), .dout(n13696));
  jand g13413(.dina(n13696), .dinb(n13694), .dout(n13697));
  jor  g13414(.dina(n13697), .dinb(n13689), .dout(n13698));
  jxor g13415(.dina(n13144), .dinb(n199), .dout(n13699));
  jand g13416(.dina(n13699), .dinb(asqrt[14] ), .dout(n13700));
  jxor g13417(.dina(n13700), .dinb(n13149), .dout(n13701));
  jnot g13418(.din(n13151), .dout(n13702));
  jnot g13419(.din(n13155), .dout(n13703));
  jand g13420(.dina(asqrt[14] ), .dinb(n13703), .dout(n13704));
  jand g13421(.dina(n13704), .dinb(n13702), .dout(n13705));
  jor  g13422(.dina(n13705), .dinb(n13162), .dout(n13706));
  jor  g13423(.dina(n13706), .dinb(n13701), .dout(n13707));
  jnot g13424(.din(n13707), .dout(n13708));
  jand g13425(.dina(n13708), .dinb(n13698), .dout(n13709));
  jor  g13426(.dina(n13709), .dinb(asqrt[63] ), .dout(n13710));
  jnot g13427(.din(n13701), .dout(n13711));
  jor  g13428(.dina(n13711), .dinb(n13698), .dout(n13712));
  jor  g13429(.dina(n13704), .dinb(n13702), .dout(n13713));
  jand g13430(.dina(n13703), .dinb(n13702), .dout(n13714));
  jor  g13431(.dina(n13714), .dinb(n194), .dout(n13715));
  jnot g13432(.din(n13715), .dout(n13716));
  jand g13433(.dina(n13716), .dinb(n13713), .dout(n13717));
  jnot g13434(.din(asqrt[14] ), .dout(n13718));
  jnot g13435(.din(n13717), .dout(n13721));
  jand g13436(.dina(n13721), .dinb(n13712), .dout(n13722));
  jand g13437(.dina(n13722), .dinb(n13710), .dout(n13723));
  jxor g13438(.dina(n13545), .dinb(n1317), .dout(n13724));
  jor  g13439(.dina(n13724), .dinb(n13723), .dout(n13725));
  jxor g13440(.dina(n13725), .dinb(n13175), .dout(n13726));
  jor  g13441(.dina(n13723), .dinb(n13177), .dout(n13727));
  jnot g13442(.din(a[24] ), .dout(n13728));
  jnot g13443(.din(a[25] ), .dout(n13729));
  jand g13444(.dina(n13177), .dinb(n13729), .dout(n13730));
  jand g13445(.dina(n13730), .dinb(n13728), .dout(n13731));
  jnot g13446(.din(n13731), .dout(n13732));
  jand g13447(.dina(n13732), .dinb(n13727), .dout(n13733));
  jor  g13448(.dina(n13733), .dinb(n13718), .dout(n13734));
  jor  g13449(.dina(n13723), .dinb(a[26] ), .dout(n13735));
  jxor g13450(.dina(n13735), .dinb(n13178), .dout(n13736));
  jand g13451(.dina(n13733), .dinb(n13718), .dout(n13737));
  jor  g13452(.dina(n13737), .dinb(n13736), .dout(n13738));
  jand g13453(.dina(n13738), .dinb(n13734), .dout(n13739));
  jor  g13454(.dina(n13739), .dinb(n12675), .dout(n13740));
  jand g13455(.dina(n13734), .dinb(n12675), .dout(n13741));
  jand g13456(.dina(n13741), .dinb(n13738), .dout(n13742));
  jor  g13457(.dina(n13735), .dinb(a[27] ), .dout(n13743));
  jnot g13458(.din(n13710), .dout(n13744));
  jnot g13459(.din(n13712), .dout(n13745));
  jor  g13460(.dina(n13717), .dinb(n13718), .dout(n13746));
  jor  g13461(.dina(n13746), .dinb(n13745), .dout(n13747));
  jor  g13462(.dina(n13747), .dinb(n13744), .dout(n13748));
  jand g13463(.dina(n13748), .dinb(n13743), .dout(n13749));
  jxor g13464(.dina(n13749), .dinb(n12681), .dout(n13750));
  jor  g13465(.dina(n13750), .dinb(n13742), .dout(n13751));
  jand g13466(.dina(n13751), .dinb(n13740), .dout(n13752));
  jor  g13467(.dina(n13752), .dinb(n12670), .dout(n13753));
  jand g13468(.dina(n13752), .dinb(n12670), .dout(n13754));
  jxor g13469(.dina(n13181), .dinb(n12675), .dout(n13755));
  jor  g13470(.dina(n13755), .dinb(n13723), .dout(n13756));
  jxor g13471(.dina(n13756), .dinb(n13184), .dout(n13757));
  jor  g13472(.dina(n13757), .dinb(n13754), .dout(n13758));
  jand g13473(.dina(n13758), .dinb(n13753), .dout(n13759));
  jor  g13474(.dina(n13759), .dinb(n11662), .dout(n13760));
  jnot g13475(.din(n13190), .dout(n13761));
  jor  g13476(.dina(n13761), .dinb(n13188), .dout(n13762));
  jor  g13477(.dina(n13762), .dinb(n13723), .dout(n13763));
  jxor g13478(.dina(n13763), .dinb(n13199), .dout(n13764));
  jand g13479(.dina(n13753), .dinb(n11662), .dout(n13765));
  jand g13480(.dina(n13765), .dinb(n13758), .dout(n13766));
  jor  g13481(.dina(n13766), .dinb(n13764), .dout(n13767));
  jand g13482(.dina(n13767), .dinb(n13760), .dout(n13768));
  jor  g13483(.dina(n13768), .dinb(n11657), .dout(n13769));
  jand g13484(.dina(n13768), .dinb(n11657), .dout(n13770));
  jxor g13485(.dina(n13201), .dinb(n11662), .dout(n13771));
  jor  g13486(.dina(n13771), .dinb(n13723), .dout(n13772));
  jxor g13487(.dina(n13772), .dinb(n13206), .dout(n13773));
  jnot g13488(.din(n13773), .dout(n13774));
  jor  g13489(.dina(n13774), .dinb(n13770), .dout(n13775));
  jand g13490(.dina(n13775), .dinb(n13769), .dout(n13776));
  jor  g13491(.dina(n13776), .dinb(n10701), .dout(n13777));
  jand g13492(.dina(n13769), .dinb(n10701), .dout(n13778));
  jand g13493(.dina(n13778), .dinb(n13775), .dout(n13779));
  jnot g13494(.din(n13210), .dout(n13780));
  jnot g13495(.din(n13723), .dout(asqrt[13] ));
  jand g13496(.dina(asqrt[13] ), .dinb(n13780), .dout(n13782));
  jand g13497(.dina(n13782), .dinb(n13217), .dout(n13783));
  jor  g13498(.dina(n13783), .dinb(n13215), .dout(n13784));
  jand g13499(.dina(n13782), .dinb(n13218), .dout(n13785));
  jnot g13500(.din(n13785), .dout(n13786));
  jand g13501(.dina(n13786), .dinb(n13784), .dout(n13787));
  jnot g13502(.din(n13787), .dout(n13788));
  jor  g13503(.dina(n13788), .dinb(n13779), .dout(n13789));
  jand g13504(.dina(n13789), .dinb(n13777), .dout(n13790));
  jor  g13505(.dina(n13790), .dinb(n10696), .dout(n13791));
  jand g13506(.dina(n13790), .dinb(n10696), .dout(n13792));
  jnot g13507(.din(n13225), .dout(n13793));
  jxor g13508(.dina(n13219), .dinb(n10701), .dout(n13794));
  jor  g13509(.dina(n13794), .dinb(n13723), .dout(n13795));
  jxor g13510(.dina(n13795), .dinb(n13793), .dout(n13796));
  jnot g13511(.din(n13796), .dout(n13797));
  jor  g13512(.dina(n13797), .dinb(n13792), .dout(n13798));
  jand g13513(.dina(n13798), .dinb(n13791), .dout(n13799));
  jor  g13514(.dina(n13799), .dinb(n9774), .dout(n13800));
  jnot g13515(.din(n13230), .dout(n13801));
  jor  g13516(.dina(n13801), .dinb(n13228), .dout(n13802));
  jor  g13517(.dina(n13802), .dinb(n13723), .dout(n13803));
  jxor g13518(.dina(n13803), .dinb(n13239), .dout(n13804));
  jand g13519(.dina(n13791), .dinb(n9774), .dout(n13805));
  jand g13520(.dina(n13805), .dinb(n13798), .dout(n13806));
  jor  g13521(.dina(n13806), .dinb(n13804), .dout(n13807));
  jand g13522(.dina(n13807), .dinb(n13800), .dout(n13808));
  jor  g13523(.dina(n13808), .dinb(n9769), .dout(n13809));
  jand g13524(.dina(n13808), .dinb(n9769), .dout(n13810));
  jnot g13525(.din(n13246), .dout(n13811));
  jxor g13526(.dina(n13241), .dinb(n9774), .dout(n13812));
  jor  g13527(.dina(n13812), .dinb(n13723), .dout(n13813));
  jxor g13528(.dina(n13813), .dinb(n13811), .dout(n13814));
  jnot g13529(.din(n13814), .dout(n13815));
  jor  g13530(.dina(n13815), .dinb(n13810), .dout(n13816));
  jand g13531(.dina(n13816), .dinb(n13809), .dout(n13817));
  jor  g13532(.dina(n13817), .dinb(n8898), .dout(n13818));
  jand g13533(.dina(n13809), .dinb(n8898), .dout(n13819));
  jand g13534(.dina(n13819), .dinb(n13816), .dout(n13820));
  jnot g13535(.din(n13249), .dout(n13821));
  jand g13536(.dina(asqrt[13] ), .dinb(n13821), .dout(n13822));
  jand g13537(.dina(n13822), .dinb(n13256), .dout(n13823));
  jor  g13538(.dina(n13823), .dinb(n13254), .dout(n13824));
  jand g13539(.dina(n13822), .dinb(n13257), .dout(n13825));
  jnot g13540(.din(n13825), .dout(n13826));
  jand g13541(.dina(n13826), .dinb(n13824), .dout(n13827));
  jnot g13542(.din(n13827), .dout(n13828));
  jor  g13543(.dina(n13828), .dinb(n13820), .dout(n13829));
  jand g13544(.dina(n13829), .dinb(n13818), .dout(n13830));
  jor  g13545(.dina(n13830), .dinb(n8893), .dout(n13831));
  jxor g13546(.dina(n13258), .dinb(n8898), .dout(n13832));
  jor  g13547(.dina(n13832), .dinb(n13723), .dout(n13833));
  jxor g13548(.dina(n13833), .dinb(n13263), .dout(n13834));
  jand g13549(.dina(n13830), .dinb(n8893), .dout(n13835));
  jor  g13550(.dina(n13835), .dinb(n13834), .dout(n13836));
  jand g13551(.dina(n13836), .dinb(n13831), .dout(n13837));
  jor  g13552(.dina(n13837), .dinb(n8058), .dout(n13838));
  jnot g13553(.din(n13268), .dout(n13839));
  jor  g13554(.dina(n13839), .dinb(n13266), .dout(n13840));
  jor  g13555(.dina(n13840), .dinb(n13723), .dout(n13841));
  jxor g13556(.dina(n13841), .dinb(n13277), .dout(n13842));
  jand g13557(.dina(n13831), .dinb(n8058), .dout(n13843));
  jand g13558(.dina(n13843), .dinb(n13836), .dout(n13844));
  jor  g13559(.dina(n13844), .dinb(n13842), .dout(n13845));
  jand g13560(.dina(n13845), .dinb(n13838), .dout(n13846));
  jor  g13561(.dina(n13846), .dinb(n8053), .dout(n13847));
  jand g13562(.dina(n13846), .dinb(n8053), .dout(n13848));
  jnot g13563(.din(n13280), .dout(n13849));
  jand g13564(.dina(asqrt[13] ), .dinb(n13849), .dout(n13850));
  jand g13565(.dina(n13850), .dinb(n13285), .dout(n13851));
  jor  g13566(.dina(n13851), .dinb(n13284), .dout(n13852));
  jand g13567(.dina(n13850), .dinb(n13286), .dout(n13853));
  jnot g13568(.din(n13853), .dout(n13854));
  jand g13569(.dina(n13854), .dinb(n13852), .dout(n13855));
  jnot g13570(.din(n13855), .dout(n13856));
  jor  g13571(.dina(n13856), .dinb(n13848), .dout(n13857));
  jand g13572(.dina(n13857), .dinb(n13847), .dout(n13858));
  jor  g13573(.dina(n13858), .dinb(n7265), .dout(n13859));
  jand g13574(.dina(n13847), .dinb(n7265), .dout(n13860));
  jand g13575(.dina(n13860), .dinb(n13857), .dout(n13861));
  jnot g13576(.din(n13288), .dout(n13862));
  jand g13577(.dina(asqrt[13] ), .dinb(n13862), .dout(n13863));
  jand g13578(.dina(n13863), .dinb(n13295), .dout(n13864));
  jor  g13579(.dina(n13864), .dinb(n13293), .dout(n13865));
  jand g13580(.dina(n13863), .dinb(n13296), .dout(n13866));
  jnot g13581(.din(n13866), .dout(n13867));
  jand g13582(.dina(n13867), .dinb(n13865), .dout(n13868));
  jnot g13583(.din(n13868), .dout(n13869));
  jor  g13584(.dina(n13869), .dinb(n13861), .dout(n13870));
  jand g13585(.dina(n13870), .dinb(n13859), .dout(n13871));
  jor  g13586(.dina(n13871), .dinb(n7260), .dout(n13872));
  jxor g13587(.dina(n13297), .dinb(n7265), .dout(n13873));
  jor  g13588(.dina(n13873), .dinb(n13723), .dout(n13874));
  jxor g13589(.dina(n13874), .dinb(n13308), .dout(n13875));
  jand g13590(.dina(n13871), .dinb(n7260), .dout(n13876));
  jor  g13591(.dina(n13876), .dinb(n13875), .dout(n13877));
  jand g13592(.dina(n13877), .dinb(n13872), .dout(n13878));
  jor  g13593(.dina(n13878), .dinb(n6505), .dout(n13879));
  jnot g13594(.din(n13313), .dout(n13880));
  jor  g13595(.dina(n13880), .dinb(n13311), .dout(n13881));
  jor  g13596(.dina(n13881), .dinb(n13723), .dout(n13882));
  jxor g13597(.dina(n13882), .dinb(n13322), .dout(n13883));
  jand g13598(.dina(n13872), .dinb(n6505), .dout(n13884));
  jand g13599(.dina(n13884), .dinb(n13877), .dout(n13885));
  jor  g13600(.dina(n13885), .dinb(n13883), .dout(n13886));
  jand g13601(.dina(n13886), .dinb(n13879), .dout(n13887));
  jor  g13602(.dina(n13887), .dinb(n6500), .dout(n13888));
  jand g13603(.dina(n13887), .dinb(n6500), .dout(n13889));
  jnot g13604(.din(n13325), .dout(n13890));
  jand g13605(.dina(asqrt[13] ), .dinb(n13890), .dout(n13891));
  jand g13606(.dina(n13891), .dinb(n13330), .dout(n13892));
  jor  g13607(.dina(n13892), .dinb(n13329), .dout(n13893));
  jand g13608(.dina(n13891), .dinb(n13331), .dout(n13894));
  jnot g13609(.din(n13894), .dout(n13895));
  jand g13610(.dina(n13895), .dinb(n13893), .dout(n13896));
  jnot g13611(.din(n13896), .dout(n13897));
  jor  g13612(.dina(n13897), .dinb(n13889), .dout(n13898));
  jand g13613(.dina(n13898), .dinb(n13888), .dout(n13899));
  jor  g13614(.dina(n13899), .dinb(n5793), .dout(n13900));
  jand g13615(.dina(n13888), .dinb(n5793), .dout(n13901));
  jand g13616(.dina(n13901), .dinb(n13898), .dout(n13902));
  jnot g13617(.din(n13333), .dout(n13903));
  jand g13618(.dina(asqrt[13] ), .dinb(n13903), .dout(n13904));
  jand g13619(.dina(n13904), .dinb(n13340), .dout(n13905));
  jor  g13620(.dina(n13905), .dinb(n13338), .dout(n13906));
  jand g13621(.dina(n13904), .dinb(n13341), .dout(n13907));
  jnot g13622(.din(n13907), .dout(n13908));
  jand g13623(.dina(n13908), .dinb(n13906), .dout(n13909));
  jnot g13624(.din(n13909), .dout(n13910));
  jor  g13625(.dina(n13910), .dinb(n13902), .dout(n13911));
  jand g13626(.dina(n13911), .dinb(n13900), .dout(n13912));
  jor  g13627(.dina(n13912), .dinb(n5788), .dout(n13913));
  jxor g13628(.dina(n13342), .dinb(n5793), .dout(n13914));
  jor  g13629(.dina(n13914), .dinb(n13723), .dout(n13915));
  jxor g13630(.dina(n13915), .dinb(n13353), .dout(n13916));
  jand g13631(.dina(n13912), .dinb(n5788), .dout(n13917));
  jor  g13632(.dina(n13917), .dinb(n13916), .dout(n13918));
  jand g13633(.dina(n13918), .dinb(n13913), .dout(n13919));
  jor  g13634(.dina(n13919), .dinb(n5121), .dout(n13920));
  jnot g13635(.din(n13358), .dout(n13921));
  jor  g13636(.dina(n13921), .dinb(n13356), .dout(n13922));
  jor  g13637(.dina(n13922), .dinb(n13723), .dout(n13923));
  jxor g13638(.dina(n13923), .dinb(n13367), .dout(n13924));
  jand g13639(.dina(n13913), .dinb(n5121), .dout(n13925));
  jand g13640(.dina(n13925), .dinb(n13918), .dout(n13926));
  jor  g13641(.dina(n13926), .dinb(n13924), .dout(n13927));
  jand g13642(.dina(n13927), .dinb(n13920), .dout(n13928));
  jor  g13643(.dina(n13928), .dinb(n5116), .dout(n13929));
  jand g13644(.dina(n13928), .dinb(n5116), .dout(n13930));
  jnot g13645(.din(n13370), .dout(n13931));
  jand g13646(.dina(asqrt[13] ), .dinb(n13931), .dout(n13932));
  jand g13647(.dina(n13932), .dinb(n13375), .dout(n13933));
  jor  g13648(.dina(n13933), .dinb(n13374), .dout(n13934));
  jand g13649(.dina(n13932), .dinb(n13376), .dout(n13935));
  jnot g13650(.din(n13935), .dout(n13936));
  jand g13651(.dina(n13936), .dinb(n13934), .dout(n13937));
  jnot g13652(.din(n13937), .dout(n13938));
  jor  g13653(.dina(n13938), .dinb(n13930), .dout(n13939));
  jand g13654(.dina(n13939), .dinb(n13929), .dout(n13940));
  jor  g13655(.dina(n13940), .dinb(n4499), .dout(n13941));
  jand g13656(.dina(n13929), .dinb(n4499), .dout(n13942));
  jand g13657(.dina(n13942), .dinb(n13939), .dout(n13943));
  jnot g13658(.din(n13378), .dout(n13944));
  jand g13659(.dina(asqrt[13] ), .dinb(n13944), .dout(n13945));
  jand g13660(.dina(n13945), .dinb(n13385), .dout(n13946));
  jor  g13661(.dina(n13946), .dinb(n13383), .dout(n13947));
  jand g13662(.dina(n13945), .dinb(n13386), .dout(n13948));
  jnot g13663(.din(n13948), .dout(n13949));
  jand g13664(.dina(n13949), .dinb(n13947), .dout(n13950));
  jnot g13665(.din(n13950), .dout(n13951));
  jor  g13666(.dina(n13951), .dinb(n13943), .dout(n13952));
  jand g13667(.dina(n13952), .dinb(n13941), .dout(n13953));
  jor  g13668(.dina(n13953), .dinb(n4494), .dout(n13954));
  jxor g13669(.dina(n13387), .dinb(n4499), .dout(n13955));
  jor  g13670(.dina(n13955), .dinb(n13723), .dout(n13956));
  jxor g13671(.dina(n13956), .dinb(n13398), .dout(n13957));
  jand g13672(.dina(n13953), .dinb(n4494), .dout(n13958));
  jor  g13673(.dina(n13958), .dinb(n13957), .dout(n13959));
  jand g13674(.dina(n13959), .dinb(n13954), .dout(n13960));
  jor  g13675(.dina(n13960), .dinb(n3912), .dout(n13961));
  jnot g13676(.din(n13403), .dout(n13962));
  jor  g13677(.dina(n13962), .dinb(n13401), .dout(n13963));
  jor  g13678(.dina(n13963), .dinb(n13723), .dout(n13964));
  jxor g13679(.dina(n13964), .dinb(n13412), .dout(n13965));
  jand g13680(.dina(n13954), .dinb(n3912), .dout(n13966));
  jand g13681(.dina(n13966), .dinb(n13959), .dout(n13967));
  jor  g13682(.dina(n13967), .dinb(n13965), .dout(n13968));
  jand g13683(.dina(n13968), .dinb(n13961), .dout(n13969));
  jor  g13684(.dina(n13969), .dinb(n3907), .dout(n13970));
  jand g13685(.dina(n13969), .dinb(n3907), .dout(n13971));
  jnot g13686(.din(n13415), .dout(n13972));
  jand g13687(.dina(asqrt[13] ), .dinb(n13972), .dout(n13973));
  jand g13688(.dina(n13973), .dinb(n13420), .dout(n13974));
  jor  g13689(.dina(n13974), .dinb(n13419), .dout(n13975));
  jand g13690(.dina(n13973), .dinb(n13421), .dout(n13976));
  jnot g13691(.din(n13976), .dout(n13977));
  jand g13692(.dina(n13977), .dinb(n13975), .dout(n13978));
  jnot g13693(.din(n13978), .dout(n13979));
  jor  g13694(.dina(n13979), .dinb(n13971), .dout(n13980));
  jand g13695(.dina(n13980), .dinb(n13970), .dout(n13981));
  jor  g13696(.dina(n13981), .dinb(n3376), .dout(n13982));
  jand g13697(.dina(n13970), .dinb(n3376), .dout(n13983));
  jand g13698(.dina(n13983), .dinb(n13980), .dout(n13984));
  jnot g13699(.din(n13423), .dout(n13985));
  jand g13700(.dina(asqrt[13] ), .dinb(n13985), .dout(n13986));
  jand g13701(.dina(n13986), .dinb(n13430), .dout(n13987));
  jor  g13702(.dina(n13987), .dinb(n13428), .dout(n13988));
  jand g13703(.dina(n13986), .dinb(n13431), .dout(n13989));
  jnot g13704(.din(n13989), .dout(n13990));
  jand g13705(.dina(n13990), .dinb(n13988), .dout(n13991));
  jnot g13706(.din(n13991), .dout(n13992));
  jor  g13707(.dina(n13992), .dinb(n13984), .dout(n13993));
  jand g13708(.dina(n13993), .dinb(n13982), .dout(n13994));
  jor  g13709(.dina(n13994), .dinb(n3371), .dout(n13995));
  jxor g13710(.dina(n13432), .dinb(n3376), .dout(n13996));
  jor  g13711(.dina(n13996), .dinb(n13723), .dout(n13997));
  jxor g13712(.dina(n13997), .dinb(n13443), .dout(n13998));
  jand g13713(.dina(n13994), .dinb(n3371), .dout(n13999));
  jor  g13714(.dina(n13999), .dinb(n13998), .dout(n14000));
  jand g13715(.dina(n14000), .dinb(n13995), .dout(n14001));
  jor  g13716(.dina(n14001), .dinb(n2875), .dout(n14002));
  jnot g13717(.din(n13448), .dout(n14003));
  jor  g13718(.dina(n14003), .dinb(n13446), .dout(n14004));
  jor  g13719(.dina(n14004), .dinb(n13723), .dout(n14005));
  jxor g13720(.dina(n14005), .dinb(n13457), .dout(n14006));
  jand g13721(.dina(n13995), .dinb(n2875), .dout(n14007));
  jand g13722(.dina(n14007), .dinb(n14000), .dout(n14008));
  jor  g13723(.dina(n14008), .dinb(n14006), .dout(n14009));
  jand g13724(.dina(n14009), .dinb(n14002), .dout(n14010));
  jor  g13725(.dina(n14010), .dinb(n2870), .dout(n14011));
  jand g13726(.dina(n14010), .dinb(n2870), .dout(n14012));
  jnot g13727(.din(n13460), .dout(n14013));
  jand g13728(.dina(asqrt[13] ), .dinb(n14013), .dout(n14014));
  jand g13729(.dina(n14014), .dinb(n13465), .dout(n14015));
  jor  g13730(.dina(n14015), .dinb(n13464), .dout(n14016));
  jand g13731(.dina(n14014), .dinb(n13466), .dout(n14017));
  jnot g13732(.din(n14017), .dout(n14018));
  jand g13733(.dina(n14018), .dinb(n14016), .dout(n14019));
  jnot g13734(.din(n14019), .dout(n14020));
  jor  g13735(.dina(n14020), .dinb(n14012), .dout(n14021));
  jand g13736(.dina(n14021), .dinb(n14011), .dout(n14022));
  jor  g13737(.dina(n14022), .dinb(n2425), .dout(n14023));
  jand g13738(.dina(n14011), .dinb(n2425), .dout(n14024));
  jand g13739(.dina(n14024), .dinb(n14021), .dout(n14025));
  jnot g13740(.din(n13468), .dout(n14026));
  jand g13741(.dina(asqrt[13] ), .dinb(n14026), .dout(n14027));
  jand g13742(.dina(n14027), .dinb(n13475), .dout(n14028));
  jor  g13743(.dina(n14028), .dinb(n13473), .dout(n14029));
  jand g13744(.dina(n14027), .dinb(n13476), .dout(n14030));
  jnot g13745(.din(n14030), .dout(n14031));
  jand g13746(.dina(n14031), .dinb(n14029), .dout(n14032));
  jnot g13747(.din(n14032), .dout(n14033));
  jor  g13748(.dina(n14033), .dinb(n14025), .dout(n14034));
  jand g13749(.dina(n14034), .dinb(n14023), .dout(n14035));
  jor  g13750(.dina(n14035), .dinb(n2420), .dout(n14036));
  jxor g13751(.dina(n13477), .dinb(n2425), .dout(n14037));
  jor  g13752(.dina(n14037), .dinb(n13723), .dout(n14038));
  jxor g13753(.dina(n14038), .dinb(n13488), .dout(n14039));
  jand g13754(.dina(n14035), .dinb(n2420), .dout(n14040));
  jor  g13755(.dina(n14040), .dinb(n14039), .dout(n14041));
  jand g13756(.dina(n14041), .dinb(n14036), .dout(n14042));
  jor  g13757(.dina(n14042), .dinb(n2010), .dout(n14043));
  jnot g13758(.din(n13493), .dout(n14044));
  jor  g13759(.dina(n14044), .dinb(n13491), .dout(n14045));
  jor  g13760(.dina(n14045), .dinb(n13723), .dout(n14046));
  jxor g13761(.dina(n14046), .dinb(n13502), .dout(n14047));
  jand g13762(.dina(n14036), .dinb(n2010), .dout(n14048));
  jand g13763(.dina(n14048), .dinb(n14041), .dout(n14049));
  jor  g13764(.dina(n14049), .dinb(n14047), .dout(n14050));
  jand g13765(.dina(n14050), .dinb(n14043), .dout(n14051));
  jor  g13766(.dina(n14051), .dinb(n2005), .dout(n14052));
  jand g13767(.dina(n14051), .dinb(n2005), .dout(n14053));
  jnot g13768(.din(n13505), .dout(n14054));
  jand g13769(.dina(asqrt[13] ), .dinb(n14054), .dout(n14055));
  jand g13770(.dina(n14055), .dinb(n13510), .dout(n14056));
  jor  g13771(.dina(n14056), .dinb(n13509), .dout(n14057));
  jand g13772(.dina(n14055), .dinb(n13511), .dout(n14058));
  jnot g13773(.din(n14058), .dout(n14059));
  jand g13774(.dina(n14059), .dinb(n14057), .dout(n14060));
  jnot g13775(.din(n14060), .dout(n14061));
  jor  g13776(.dina(n14061), .dinb(n14053), .dout(n14062));
  jand g13777(.dina(n14062), .dinb(n14052), .dout(n14063));
  jor  g13778(.dina(n14063), .dinb(n1646), .dout(n14064));
  jand g13779(.dina(n14052), .dinb(n1646), .dout(n14065));
  jand g13780(.dina(n14065), .dinb(n14062), .dout(n14066));
  jnot g13781(.din(n13513), .dout(n14067));
  jand g13782(.dina(asqrt[13] ), .dinb(n14067), .dout(n14068));
  jand g13783(.dina(n14068), .dinb(n13520), .dout(n14069));
  jor  g13784(.dina(n14069), .dinb(n13518), .dout(n14070));
  jand g13785(.dina(n14068), .dinb(n13521), .dout(n14071));
  jnot g13786(.din(n14071), .dout(n14072));
  jand g13787(.dina(n14072), .dinb(n14070), .dout(n14073));
  jnot g13788(.din(n14073), .dout(n14074));
  jor  g13789(.dina(n14074), .dinb(n14066), .dout(n14075));
  jand g13790(.dina(n14075), .dinb(n14064), .dout(n14076));
  jor  g13791(.dina(n14076), .dinb(n1641), .dout(n14077));
  jxor g13792(.dina(n13522), .dinb(n1646), .dout(n14078));
  jor  g13793(.dina(n14078), .dinb(n13723), .dout(n14079));
  jxor g13794(.dina(n14079), .dinb(n13533), .dout(n14080));
  jand g13795(.dina(n14076), .dinb(n1641), .dout(n14081));
  jor  g13796(.dina(n14081), .dinb(n14080), .dout(n14082));
  jand g13797(.dina(n14082), .dinb(n14077), .dout(n14083));
  jor  g13798(.dina(n14083), .dinb(n1317), .dout(n14084));
  jand g13799(.dina(n14077), .dinb(n1317), .dout(n14085));
  jand g13800(.dina(n14085), .dinb(n14082), .dout(n14086));
  jnot g13801(.din(n13536), .dout(n14087));
  jand g13802(.dina(asqrt[13] ), .dinb(n14087), .dout(n14088));
  jand g13803(.dina(n14088), .dinb(n13543), .dout(n14089));
  jor  g13804(.dina(n14089), .dinb(n13541), .dout(n14090));
  jand g13805(.dina(n14088), .dinb(n13544), .dout(n14091));
  jnot g13806(.din(n14091), .dout(n14092));
  jand g13807(.dina(n14092), .dinb(n14090), .dout(n14093));
  jnot g13808(.din(n14093), .dout(n14094));
  jor  g13809(.dina(n14094), .dinb(n14086), .dout(n14095));
  jand g13810(.dina(n14095), .dinb(n14084), .dout(n14096));
  jor  g13811(.dina(n14096), .dinb(n1312), .dout(n14097));
  jand g13812(.dina(n14096), .dinb(n1312), .dout(n14098));
  jor  g13813(.dina(n14098), .dinb(n13726), .dout(n14099));
  jand g13814(.dina(n14099), .dinb(n14097), .dout(n14100));
  jor  g13815(.dina(n14100), .dinb(n1039), .dout(n14101));
  jnot g13816(.din(n13552), .dout(n14102));
  jor  g13817(.dina(n14102), .dinb(n13550), .dout(n14103));
  jor  g13818(.dina(n14103), .dinb(n13723), .dout(n14104));
  jxor g13819(.dina(n14104), .dinb(n13561), .dout(n14105));
  jand g13820(.dina(n14097), .dinb(n1039), .dout(n14106));
  jand g13821(.dina(n14106), .dinb(n14099), .dout(n14107));
  jor  g13822(.dina(n14107), .dinb(n14105), .dout(n14108));
  jand g13823(.dina(n14108), .dinb(n14101), .dout(n14109));
  jor  g13824(.dina(n14109), .dinb(n1034), .dout(n14110));
  jxor g13825(.dina(n13563), .dinb(n1039), .dout(n14111));
  jor  g13826(.dina(n14111), .dinb(n13723), .dout(n14112));
  jxor g13827(.dina(n14112), .dinb(n13574), .dout(n14113));
  jand g13828(.dina(n14109), .dinb(n1034), .dout(n14114));
  jor  g13829(.dina(n14114), .dinb(n14113), .dout(n14115));
  jand g13830(.dina(n14115), .dinb(n14110), .dout(n14116));
  jor  g13831(.dina(n14116), .dinb(n796), .dout(n14117));
  jnot g13832(.din(n13579), .dout(n14118));
  jor  g13833(.dina(n14118), .dinb(n13577), .dout(n14119));
  jor  g13834(.dina(n14119), .dinb(n13723), .dout(n14120));
  jxor g13835(.dina(n14120), .dinb(n13588), .dout(n14121));
  jand g13836(.dina(n14110), .dinb(n796), .dout(n14122));
  jand g13837(.dina(n14122), .dinb(n14115), .dout(n14123));
  jor  g13838(.dina(n14123), .dinb(n14121), .dout(n14124));
  jand g13839(.dina(n14124), .dinb(n14117), .dout(n14125));
  jor  g13840(.dina(n14125), .dinb(n791), .dout(n14126));
  jand g13841(.dina(n14125), .dinb(n791), .dout(n14127));
  jnot g13842(.din(n13591), .dout(n14128));
  jand g13843(.dina(asqrt[13] ), .dinb(n14128), .dout(n14129));
  jand g13844(.dina(n14129), .dinb(n13596), .dout(n14130));
  jor  g13845(.dina(n14130), .dinb(n13595), .dout(n14131));
  jand g13846(.dina(n14129), .dinb(n13597), .dout(n14132));
  jnot g13847(.din(n14132), .dout(n14133));
  jand g13848(.dina(n14133), .dinb(n14131), .dout(n14134));
  jnot g13849(.din(n14134), .dout(n14135));
  jor  g13850(.dina(n14135), .dinb(n14127), .dout(n14136));
  jand g13851(.dina(n14136), .dinb(n14126), .dout(n14137));
  jor  g13852(.dina(n14137), .dinb(n595), .dout(n14138));
  jand g13853(.dina(n14126), .dinb(n595), .dout(n14139));
  jand g13854(.dina(n14139), .dinb(n14136), .dout(n14140));
  jnot g13855(.din(n13599), .dout(n14141));
  jand g13856(.dina(asqrt[13] ), .dinb(n14141), .dout(n14142));
  jand g13857(.dina(n14142), .dinb(n13606), .dout(n14143));
  jor  g13858(.dina(n14143), .dinb(n13604), .dout(n14144));
  jand g13859(.dina(n14142), .dinb(n13607), .dout(n14145));
  jnot g13860(.din(n14145), .dout(n14146));
  jand g13861(.dina(n14146), .dinb(n14144), .dout(n14147));
  jnot g13862(.din(n14147), .dout(n14148));
  jor  g13863(.dina(n14148), .dinb(n14140), .dout(n14149));
  jand g13864(.dina(n14149), .dinb(n14138), .dout(n14150));
  jor  g13865(.dina(n14150), .dinb(n590), .dout(n14151));
  jxor g13866(.dina(n13608), .dinb(n595), .dout(n14152));
  jor  g13867(.dina(n14152), .dinb(n13723), .dout(n14153));
  jxor g13868(.dina(n14153), .dinb(n13619), .dout(n14154));
  jand g13869(.dina(n14150), .dinb(n590), .dout(n14155));
  jor  g13870(.dina(n14155), .dinb(n14154), .dout(n14156));
  jand g13871(.dina(n14156), .dinb(n14151), .dout(n14157));
  jor  g13872(.dina(n14157), .dinb(n430), .dout(n14158));
  jnot g13873(.din(n13624), .dout(n14159));
  jor  g13874(.dina(n14159), .dinb(n13622), .dout(n14160));
  jor  g13875(.dina(n14160), .dinb(n13723), .dout(n14161));
  jxor g13876(.dina(n14161), .dinb(n13633), .dout(n14162));
  jand g13877(.dina(n14151), .dinb(n430), .dout(n14163));
  jand g13878(.dina(n14163), .dinb(n14156), .dout(n14164));
  jor  g13879(.dina(n14164), .dinb(n14162), .dout(n14165));
  jand g13880(.dina(n14165), .dinb(n14158), .dout(n14166));
  jor  g13881(.dina(n14166), .dinb(n425), .dout(n14167));
  jand g13882(.dina(n14166), .dinb(n425), .dout(n14168));
  jnot g13883(.din(n13636), .dout(n14169));
  jand g13884(.dina(asqrt[13] ), .dinb(n14169), .dout(n14170));
  jand g13885(.dina(n14170), .dinb(n13641), .dout(n14171));
  jor  g13886(.dina(n14171), .dinb(n13640), .dout(n14172));
  jand g13887(.dina(n14170), .dinb(n13642), .dout(n14173));
  jnot g13888(.din(n14173), .dout(n14174));
  jand g13889(.dina(n14174), .dinb(n14172), .dout(n14175));
  jnot g13890(.din(n14175), .dout(n14176));
  jor  g13891(.dina(n14176), .dinb(n14168), .dout(n14177));
  jand g13892(.dina(n14177), .dinb(n14167), .dout(n14178));
  jor  g13893(.dina(n14178), .dinb(n305), .dout(n14179));
  jand g13894(.dina(n14167), .dinb(n305), .dout(n14180));
  jand g13895(.dina(n14180), .dinb(n14177), .dout(n14181));
  jnot g13896(.din(n13644), .dout(n14182));
  jand g13897(.dina(asqrt[13] ), .dinb(n14182), .dout(n14183));
  jand g13898(.dina(n14183), .dinb(n13651), .dout(n14184));
  jor  g13899(.dina(n14184), .dinb(n13649), .dout(n14185));
  jand g13900(.dina(n14183), .dinb(n13652), .dout(n14186));
  jnot g13901(.din(n14186), .dout(n14187));
  jand g13902(.dina(n14187), .dinb(n14185), .dout(n14188));
  jnot g13903(.din(n14188), .dout(n14189));
  jor  g13904(.dina(n14189), .dinb(n14181), .dout(n14190));
  jand g13905(.dina(n14190), .dinb(n14179), .dout(n14191));
  jor  g13906(.dina(n14191), .dinb(n290), .dout(n14192));
  jxor g13907(.dina(n13653), .dinb(n305), .dout(n14193));
  jor  g13908(.dina(n14193), .dinb(n13723), .dout(n14194));
  jxor g13909(.dina(n14194), .dinb(n13664), .dout(n14195));
  jand g13910(.dina(n14191), .dinb(n290), .dout(n14196));
  jor  g13911(.dina(n14196), .dinb(n14195), .dout(n14197));
  jand g13912(.dina(n14197), .dinb(n14192), .dout(n14198));
  jor  g13913(.dina(n14198), .dinb(n223), .dout(n14199));
  jnot g13914(.din(n13669), .dout(n14200));
  jor  g13915(.dina(n14200), .dinb(n13667), .dout(n14201));
  jor  g13916(.dina(n14201), .dinb(n13723), .dout(n14202));
  jxor g13917(.dina(n14202), .dinb(n13678), .dout(n14203));
  jand g13918(.dina(n14192), .dinb(n223), .dout(n14204));
  jand g13919(.dina(n14204), .dinb(n14197), .dout(n14205));
  jor  g13920(.dina(n14205), .dinb(n14203), .dout(n14206));
  jand g13921(.dina(n14206), .dinb(n14199), .dout(n14207));
  jor  g13922(.dina(n14207), .dinb(n199), .dout(n14208));
  jand g13923(.dina(n14207), .dinb(n199), .dout(n14209));
  jnot g13924(.din(n13681), .dout(n14210));
  jand g13925(.dina(asqrt[13] ), .dinb(n14210), .dout(n14211));
  jand g13926(.dina(n14211), .dinb(n13686), .dout(n14212));
  jor  g13927(.dina(n14212), .dinb(n13685), .dout(n14213));
  jand g13928(.dina(n14211), .dinb(n13687), .dout(n14214));
  jnot g13929(.din(n14214), .dout(n14215));
  jand g13930(.dina(n14215), .dinb(n14213), .dout(n14216));
  jnot g13931(.din(n14216), .dout(n14217));
  jor  g13932(.dina(n14217), .dinb(n14209), .dout(n14218));
  jand g13933(.dina(n14218), .dinb(n14208), .dout(n14219));
  jnot g13934(.din(n13689), .dout(n14220));
  jand g13935(.dina(asqrt[13] ), .dinb(n14220), .dout(n14221));
  jand g13936(.dina(n14221), .dinb(n13696), .dout(n14222));
  jor  g13937(.dina(n14222), .dinb(n13694), .dout(n14223));
  jand g13938(.dina(n14221), .dinb(n13697), .dout(n14224));
  jnot g13939(.din(n14224), .dout(n14225));
  jand g13940(.dina(n14225), .dinb(n14223), .dout(n14226));
  jnot g13941(.din(n14226), .dout(n14227));
  jand g13942(.dina(asqrt[13] ), .dinb(n13711), .dout(n14228));
  jand g13943(.dina(n14228), .dinb(n13698), .dout(n14229));
  jor  g13944(.dina(n14229), .dinb(n13745), .dout(n14230));
  jor  g13945(.dina(n14230), .dinb(n14227), .dout(n14231));
  jor  g13946(.dina(n14231), .dinb(n14219), .dout(n14232));
  jand g13947(.dina(n14232), .dinb(n194), .dout(n14233));
  jand g13948(.dina(n14227), .dinb(n14219), .dout(n14234));
  jor  g13949(.dina(n14228), .dinb(n13698), .dout(n14235));
  jand g13950(.dina(n13711), .dinb(n13698), .dout(n14236));
  jor  g13951(.dina(n14236), .dinb(n194), .dout(n14237));
  jnot g13952(.din(n14237), .dout(n14238));
  jand g13953(.dina(n14238), .dinb(n14235), .dout(n14239));
  jor  g13954(.dina(n14239), .dinb(n14234), .dout(n14242));
  jor  g13955(.dina(n14242), .dinb(n14233), .dout(asqrt[12] ));
  jxor g13956(.dina(n14096), .dinb(n1312), .dout(n14244));
  jand g13957(.dina(n14244), .dinb(asqrt[12] ), .dout(n14245));
  jxor g13958(.dina(n14245), .dinb(n13726), .dout(n14246));
  jand g13959(.dina(asqrt[12] ), .dinb(a[24] ), .dout(n14247));
  jnot g13960(.din(a[22] ), .dout(n14248));
  jnot g13961(.din(a[23] ), .dout(n14249));
  jand g13962(.dina(n13728), .dinb(n14249), .dout(n14250));
  jand g13963(.dina(n14250), .dinb(n14248), .dout(n14251));
  jor  g13964(.dina(n14251), .dinb(n14247), .dout(n14252));
  jand g13965(.dina(n14252), .dinb(asqrt[13] ), .dout(n14253));
  jand g13966(.dina(asqrt[12] ), .dinb(n13728), .dout(n14254));
  jxor g13967(.dina(n14254), .dinb(n13729), .dout(n14255));
  jor  g13968(.dina(n14252), .dinb(asqrt[13] ), .dout(n14256));
  jand g13969(.dina(n14256), .dinb(n14255), .dout(n14257));
  jor  g13970(.dina(n14257), .dinb(n14253), .dout(n14258));
  jand g13971(.dina(n14258), .dinb(asqrt[14] ), .dout(n14259));
  jor  g13972(.dina(n14253), .dinb(asqrt[14] ), .dout(n14260));
  jor  g13973(.dina(n14260), .dinb(n14257), .dout(n14261));
  jand g13974(.dina(n14254), .dinb(n13729), .dout(n14262));
  jnot g13975(.din(n14233), .dout(n14263));
  jnot g13976(.din(n14234), .dout(n14264));
  jnot g13977(.din(n14239), .dout(n14265));
  jand g13978(.dina(n14265), .dinb(asqrt[13] ), .dout(n14266));
  jand g13979(.dina(n14266), .dinb(n14264), .dout(n14267));
  jand g13980(.dina(n14267), .dinb(n14263), .dout(n14268));
  jor  g13981(.dina(n14268), .dinb(n14262), .dout(n14269));
  jxor g13982(.dina(n14269), .dinb(n13177), .dout(n14270));
  jand g13983(.dina(n14270), .dinb(n14261), .dout(n14271));
  jor  g13984(.dina(n14271), .dinb(n14259), .dout(n14272));
  jand g13985(.dina(n14272), .dinb(asqrt[15] ), .dout(n14273));
  jor  g13986(.dina(n14272), .dinb(asqrt[15] ), .dout(n14274));
  jxor g13987(.dina(n13733), .dinb(n13718), .dout(n14275));
  jand g13988(.dina(n14275), .dinb(asqrt[12] ), .dout(n14276));
  jxor g13989(.dina(n14276), .dinb(n13736), .dout(n14277));
  jnot g13990(.din(n14277), .dout(n14278));
  jand g13991(.dina(n14278), .dinb(n14274), .dout(n14279));
  jor  g13992(.dina(n14279), .dinb(n14273), .dout(n14280));
  jand g13993(.dina(n14280), .dinb(asqrt[16] ), .dout(n14281));
  jnot g13994(.din(n13742), .dout(n14282));
  jand g13995(.dina(n14282), .dinb(n13740), .dout(n14283));
  jand g13996(.dina(n14283), .dinb(asqrt[12] ), .dout(n14284));
  jxor g13997(.dina(n14284), .dinb(n13750), .dout(n14285));
  jnot g13998(.din(n14285), .dout(n14286));
  jor  g13999(.dina(n14273), .dinb(asqrt[16] ), .dout(n14287));
  jor  g14000(.dina(n14287), .dinb(n14279), .dout(n14288));
  jand g14001(.dina(n14288), .dinb(n14286), .dout(n14289));
  jor  g14002(.dina(n14289), .dinb(n14281), .dout(n14290));
  jand g14003(.dina(n14290), .dinb(asqrt[17] ), .dout(n14291));
  jor  g14004(.dina(n14290), .dinb(asqrt[17] ), .dout(n14292));
  jnot g14005(.din(n13757), .dout(n14293));
  jxor g14006(.dina(n13752), .dinb(n12670), .dout(n14294));
  jand g14007(.dina(n14294), .dinb(asqrt[12] ), .dout(n14295));
  jxor g14008(.dina(n14295), .dinb(n14293), .dout(n14296));
  jand g14009(.dina(n14296), .dinb(n14292), .dout(n14297));
  jor  g14010(.dina(n14297), .dinb(n14291), .dout(n14298));
  jand g14011(.dina(n14298), .dinb(asqrt[18] ), .dout(n14299));
  jor  g14012(.dina(n14291), .dinb(asqrt[18] ), .dout(n14300));
  jor  g14013(.dina(n14300), .dinb(n14297), .dout(n14301));
  jnot g14014(.din(n13764), .dout(n14302));
  jnot g14015(.din(n13766), .dout(n14303));
  jand g14016(.dina(asqrt[12] ), .dinb(n13760), .dout(n14304));
  jand g14017(.dina(n14304), .dinb(n14303), .dout(n14305));
  jor  g14018(.dina(n14305), .dinb(n14302), .dout(n14306));
  jnot g14019(.din(n13767), .dout(n14307));
  jand g14020(.dina(n14304), .dinb(n14307), .dout(n14308));
  jnot g14021(.din(n14308), .dout(n14309));
  jand g14022(.dina(n14309), .dinb(n14306), .dout(n14310));
  jand g14023(.dina(n14310), .dinb(n14301), .dout(n14311));
  jor  g14024(.dina(n14311), .dinb(n14299), .dout(n14312));
  jand g14025(.dina(n14312), .dinb(asqrt[19] ), .dout(n14313));
  jor  g14026(.dina(n14312), .dinb(asqrt[19] ), .dout(n14314));
  jxor g14027(.dina(n13768), .dinb(n11657), .dout(n14315));
  jand g14028(.dina(n14315), .dinb(asqrt[12] ), .dout(n14316));
  jxor g14029(.dina(n14316), .dinb(n13773), .dout(n14317));
  jand g14030(.dina(n14317), .dinb(n14314), .dout(n14318));
  jor  g14031(.dina(n14318), .dinb(n14313), .dout(n14319));
  jand g14032(.dina(n14319), .dinb(asqrt[20] ), .dout(n14320));
  jnot g14033(.din(n13779), .dout(n14321));
  jand g14034(.dina(n14321), .dinb(n13777), .dout(n14322));
  jand g14035(.dina(n14322), .dinb(asqrt[12] ), .dout(n14323));
  jxor g14036(.dina(n14323), .dinb(n13788), .dout(n14324));
  jnot g14037(.din(n14324), .dout(n14325));
  jor  g14038(.dina(n14313), .dinb(asqrt[20] ), .dout(n14326));
  jor  g14039(.dina(n14326), .dinb(n14318), .dout(n14327));
  jand g14040(.dina(n14327), .dinb(n14325), .dout(n14328));
  jor  g14041(.dina(n14328), .dinb(n14320), .dout(n14329));
  jand g14042(.dina(n14329), .dinb(asqrt[21] ), .dout(n14330));
  jor  g14043(.dina(n14329), .dinb(asqrt[21] ), .dout(n14331));
  jxor g14044(.dina(n13790), .dinb(n10696), .dout(n14332));
  jand g14045(.dina(n14332), .dinb(asqrt[12] ), .dout(n14333));
  jxor g14046(.dina(n14333), .dinb(n13796), .dout(n14334));
  jand g14047(.dina(n14334), .dinb(n14331), .dout(n14335));
  jor  g14048(.dina(n14335), .dinb(n14330), .dout(n14336));
  jand g14049(.dina(n14336), .dinb(asqrt[22] ), .dout(n14337));
  jor  g14050(.dina(n14330), .dinb(asqrt[22] ), .dout(n14338));
  jor  g14051(.dina(n14338), .dinb(n14335), .dout(n14339));
  jnot g14052(.din(n13804), .dout(n14340));
  jnot g14053(.din(n13806), .dout(n14341));
  jand g14054(.dina(asqrt[12] ), .dinb(n13800), .dout(n14342));
  jand g14055(.dina(n14342), .dinb(n14341), .dout(n14343));
  jor  g14056(.dina(n14343), .dinb(n14340), .dout(n14344));
  jnot g14057(.din(n13807), .dout(n14345));
  jand g14058(.dina(n14342), .dinb(n14345), .dout(n14346));
  jnot g14059(.din(n14346), .dout(n14347));
  jand g14060(.dina(n14347), .dinb(n14344), .dout(n14348));
  jand g14061(.dina(n14348), .dinb(n14339), .dout(n14349));
  jor  g14062(.dina(n14349), .dinb(n14337), .dout(n14350));
  jand g14063(.dina(n14350), .dinb(asqrt[23] ), .dout(n14351));
  jxor g14064(.dina(n13808), .dinb(n9769), .dout(n14352));
  jand g14065(.dina(n14352), .dinb(asqrt[12] ), .dout(n14353));
  jxor g14066(.dina(n14353), .dinb(n13815), .dout(n14354));
  jnot g14067(.din(n14354), .dout(n14355));
  jor  g14068(.dina(n14350), .dinb(asqrt[23] ), .dout(n14356));
  jand g14069(.dina(n14356), .dinb(n14355), .dout(n14357));
  jor  g14070(.dina(n14357), .dinb(n14351), .dout(n14358));
  jand g14071(.dina(n14358), .dinb(asqrt[24] ), .dout(n14359));
  jnot g14072(.din(n13820), .dout(n14360));
  jand g14073(.dina(n14360), .dinb(n13818), .dout(n14361));
  jand g14074(.dina(n14361), .dinb(asqrt[12] ), .dout(n14362));
  jxor g14075(.dina(n14362), .dinb(n13828), .dout(n14363));
  jnot g14076(.din(n14363), .dout(n14364));
  jor  g14077(.dina(n14351), .dinb(asqrt[24] ), .dout(n14365));
  jor  g14078(.dina(n14365), .dinb(n14357), .dout(n14366));
  jand g14079(.dina(n14366), .dinb(n14364), .dout(n14367));
  jor  g14080(.dina(n14367), .dinb(n14359), .dout(n14368));
  jand g14081(.dina(n14368), .dinb(asqrt[25] ), .dout(n14369));
  jor  g14082(.dina(n14368), .dinb(asqrt[25] ), .dout(n14370));
  jnot g14083(.din(n13834), .dout(n14371));
  jnot g14084(.din(n13835), .dout(n14372));
  jand g14085(.dina(asqrt[12] ), .dinb(n13831), .dout(n14373));
  jand g14086(.dina(n14373), .dinb(n14372), .dout(n14374));
  jor  g14087(.dina(n14374), .dinb(n14371), .dout(n14375));
  jnot g14088(.din(n13836), .dout(n14376));
  jand g14089(.dina(n14373), .dinb(n14376), .dout(n14377));
  jnot g14090(.din(n14377), .dout(n14378));
  jand g14091(.dina(n14378), .dinb(n14375), .dout(n14379));
  jand g14092(.dina(n14379), .dinb(n14370), .dout(n14380));
  jor  g14093(.dina(n14380), .dinb(n14369), .dout(n14381));
  jand g14094(.dina(n14381), .dinb(asqrt[26] ), .dout(n14382));
  jor  g14095(.dina(n14369), .dinb(asqrt[26] ), .dout(n14383));
  jor  g14096(.dina(n14383), .dinb(n14380), .dout(n14384));
  jnot g14097(.din(n13842), .dout(n14385));
  jnot g14098(.din(n13844), .dout(n14386));
  jand g14099(.dina(asqrt[12] ), .dinb(n13838), .dout(n14387));
  jand g14100(.dina(n14387), .dinb(n14386), .dout(n14388));
  jor  g14101(.dina(n14388), .dinb(n14385), .dout(n14389));
  jnot g14102(.din(n13845), .dout(n14390));
  jand g14103(.dina(n14387), .dinb(n14390), .dout(n14391));
  jnot g14104(.din(n14391), .dout(n14392));
  jand g14105(.dina(n14392), .dinb(n14389), .dout(n14393));
  jand g14106(.dina(n14393), .dinb(n14384), .dout(n14394));
  jor  g14107(.dina(n14394), .dinb(n14382), .dout(n14395));
  jand g14108(.dina(n14395), .dinb(asqrt[27] ), .dout(n14396));
  jxor g14109(.dina(n13846), .dinb(n8053), .dout(n14397));
  jand g14110(.dina(n14397), .dinb(asqrt[12] ), .dout(n14398));
  jxor g14111(.dina(n14398), .dinb(n13856), .dout(n14399));
  jnot g14112(.din(n14399), .dout(n14400));
  jor  g14113(.dina(n14395), .dinb(asqrt[27] ), .dout(n14401));
  jand g14114(.dina(n14401), .dinb(n14400), .dout(n14402));
  jor  g14115(.dina(n14402), .dinb(n14396), .dout(n14403));
  jand g14116(.dina(n14403), .dinb(asqrt[28] ), .dout(n14404));
  jnot g14117(.din(n13861), .dout(n14405));
  jand g14118(.dina(n14405), .dinb(n13859), .dout(n14406));
  jand g14119(.dina(n14406), .dinb(asqrt[12] ), .dout(n14407));
  jxor g14120(.dina(n14407), .dinb(n13869), .dout(n14408));
  jnot g14121(.din(n14408), .dout(n14409));
  jor  g14122(.dina(n14396), .dinb(asqrt[28] ), .dout(n14410));
  jor  g14123(.dina(n14410), .dinb(n14402), .dout(n14411));
  jand g14124(.dina(n14411), .dinb(n14409), .dout(n14412));
  jor  g14125(.dina(n14412), .dinb(n14404), .dout(n14413));
  jand g14126(.dina(n14413), .dinb(asqrt[29] ), .dout(n14414));
  jor  g14127(.dina(n14413), .dinb(asqrt[29] ), .dout(n14415));
  jnot g14128(.din(n13875), .dout(n14416));
  jnot g14129(.din(n13876), .dout(n14417));
  jand g14130(.dina(asqrt[12] ), .dinb(n13872), .dout(n14418));
  jand g14131(.dina(n14418), .dinb(n14417), .dout(n14419));
  jor  g14132(.dina(n14419), .dinb(n14416), .dout(n14420));
  jnot g14133(.din(n13877), .dout(n14421));
  jand g14134(.dina(n14418), .dinb(n14421), .dout(n14422));
  jnot g14135(.din(n14422), .dout(n14423));
  jand g14136(.dina(n14423), .dinb(n14420), .dout(n14424));
  jand g14137(.dina(n14424), .dinb(n14415), .dout(n14425));
  jor  g14138(.dina(n14425), .dinb(n14414), .dout(n14426));
  jand g14139(.dina(n14426), .dinb(asqrt[30] ), .dout(n14427));
  jor  g14140(.dina(n14414), .dinb(asqrt[30] ), .dout(n14428));
  jor  g14141(.dina(n14428), .dinb(n14425), .dout(n14429));
  jnot g14142(.din(n13883), .dout(n14430));
  jnot g14143(.din(n13885), .dout(n14431));
  jand g14144(.dina(asqrt[12] ), .dinb(n13879), .dout(n14432));
  jand g14145(.dina(n14432), .dinb(n14431), .dout(n14433));
  jor  g14146(.dina(n14433), .dinb(n14430), .dout(n14434));
  jnot g14147(.din(n13886), .dout(n14435));
  jand g14148(.dina(n14432), .dinb(n14435), .dout(n14436));
  jnot g14149(.din(n14436), .dout(n14437));
  jand g14150(.dina(n14437), .dinb(n14434), .dout(n14438));
  jand g14151(.dina(n14438), .dinb(n14429), .dout(n14439));
  jor  g14152(.dina(n14439), .dinb(n14427), .dout(n14440));
  jand g14153(.dina(n14440), .dinb(asqrt[31] ), .dout(n14441));
  jxor g14154(.dina(n13887), .dinb(n6500), .dout(n14442));
  jand g14155(.dina(n14442), .dinb(asqrt[12] ), .dout(n14443));
  jxor g14156(.dina(n14443), .dinb(n13897), .dout(n14444));
  jnot g14157(.din(n14444), .dout(n14445));
  jor  g14158(.dina(n14440), .dinb(asqrt[31] ), .dout(n14446));
  jand g14159(.dina(n14446), .dinb(n14445), .dout(n14447));
  jor  g14160(.dina(n14447), .dinb(n14441), .dout(n14448));
  jand g14161(.dina(n14448), .dinb(asqrt[32] ), .dout(n14449));
  jnot g14162(.din(n13902), .dout(n14450));
  jand g14163(.dina(n14450), .dinb(n13900), .dout(n14451));
  jand g14164(.dina(n14451), .dinb(asqrt[12] ), .dout(n14452));
  jxor g14165(.dina(n14452), .dinb(n13910), .dout(n14453));
  jnot g14166(.din(n14453), .dout(n14454));
  jor  g14167(.dina(n14441), .dinb(asqrt[32] ), .dout(n14455));
  jor  g14168(.dina(n14455), .dinb(n14447), .dout(n14456));
  jand g14169(.dina(n14456), .dinb(n14454), .dout(n14457));
  jor  g14170(.dina(n14457), .dinb(n14449), .dout(n14458));
  jand g14171(.dina(n14458), .dinb(asqrt[33] ), .dout(n14459));
  jor  g14172(.dina(n14458), .dinb(asqrt[33] ), .dout(n14460));
  jnot g14173(.din(n13916), .dout(n14461));
  jnot g14174(.din(n13917), .dout(n14462));
  jand g14175(.dina(asqrt[12] ), .dinb(n13913), .dout(n14463));
  jand g14176(.dina(n14463), .dinb(n14462), .dout(n14464));
  jor  g14177(.dina(n14464), .dinb(n14461), .dout(n14465));
  jnot g14178(.din(n13918), .dout(n14466));
  jand g14179(.dina(n14463), .dinb(n14466), .dout(n14467));
  jnot g14180(.din(n14467), .dout(n14468));
  jand g14181(.dina(n14468), .dinb(n14465), .dout(n14469));
  jand g14182(.dina(n14469), .dinb(n14460), .dout(n14470));
  jor  g14183(.dina(n14470), .dinb(n14459), .dout(n14471));
  jand g14184(.dina(n14471), .dinb(asqrt[34] ), .dout(n14472));
  jor  g14185(.dina(n14459), .dinb(asqrt[34] ), .dout(n14473));
  jor  g14186(.dina(n14473), .dinb(n14470), .dout(n14474));
  jnot g14187(.din(n13924), .dout(n14475));
  jnot g14188(.din(n13926), .dout(n14476));
  jand g14189(.dina(asqrt[12] ), .dinb(n13920), .dout(n14477));
  jand g14190(.dina(n14477), .dinb(n14476), .dout(n14478));
  jor  g14191(.dina(n14478), .dinb(n14475), .dout(n14479));
  jnot g14192(.din(n13927), .dout(n14480));
  jand g14193(.dina(n14477), .dinb(n14480), .dout(n14481));
  jnot g14194(.din(n14481), .dout(n14482));
  jand g14195(.dina(n14482), .dinb(n14479), .dout(n14483));
  jand g14196(.dina(n14483), .dinb(n14474), .dout(n14484));
  jor  g14197(.dina(n14484), .dinb(n14472), .dout(n14485));
  jand g14198(.dina(n14485), .dinb(asqrt[35] ), .dout(n14486));
  jxor g14199(.dina(n13928), .dinb(n5116), .dout(n14487));
  jand g14200(.dina(n14487), .dinb(asqrt[12] ), .dout(n14488));
  jxor g14201(.dina(n14488), .dinb(n13938), .dout(n14489));
  jnot g14202(.din(n14489), .dout(n14490));
  jor  g14203(.dina(n14485), .dinb(asqrt[35] ), .dout(n14491));
  jand g14204(.dina(n14491), .dinb(n14490), .dout(n14492));
  jor  g14205(.dina(n14492), .dinb(n14486), .dout(n14493));
  jand g14206(.dina(n14493), .dinb(asqrt[36] ), .dout(n14494));
  jnot g14207(.din(n13943), .dout(n14495));
  jand g14208(.dina(n14495), .dinb(n13941), .dout(n14496));
  jand g14209(.dina(n14496), .dinb(asqrt[12] ), .dout(n14497));
  jxor g14210(.dina(n14497), .dinb(n13951), .dout(n14498));
  jnot g14211(.din(n14498), .dout(n14499));
  jor  g14212(.dina(n14486), .dinb(asqrt[36] ), .dout(n14500));
  jor  g14213(.dina(n14500), .dinb(n14492), .dout(n14501));
  jand g14214(.dina(n14501), .dinb(n14499), .dout(n14502));
  jor  g14215(.dina(n14502), .dinb(n14494), .dout(n14503));
  jand g14216(.dina(n14503), .dinb(asqrt[37] ), .dout(n14504));
  jor  g14217(.dina(n14503), .dinb(asqrt[37] ), .dout(n14505));
  jnot g14218(.din(n13957), .dout(n14506));
  jnot g14219(.din(n13958), .dout(n14507));
  jand g14220(.dina(asqrt[12] ), .dinb(n13954), .dout(n14508));
  jand g14221(.dina(n14508), .dinb(n14507), .dout(n14509));
  jor  g14222(.dina(n14509), .dinb(n14506), .dout(n14510));
  jnot g14223(.din(n13959), .dout(n14511));
  jand g14224(.dina(n14508), .dinb(n14511), .dout(n14512));
  jnot g14225(.din(n14512), .dout(n14513));
  jand g14226(.dina(n14513), .dinb(n14510), .dout(n14514));
  jand g14227(.dina(n14514), .dinb(n14505), .dout(n14515));
  jor  g14228(.dina(n14515), .dinb(n14504), .dout(n14516));
  jand g14229(.dina(n14516), .dinb(asqrt[38] ), .dout(n14517));
  jor  g14230(.dina(n14504), .dinb(asqrt[38] ), .dout(n14518));
  jor  g14231(.dina(n14518), .dinb(n14515), .dout(n14519));
  jnot g14232(.din(n13965), .dout(n14520));
  jnot g14233(.din(n13967), .dout(n14521));
  jand g14234(.dina(asqrt[12] ), .dinb(n13961), .dout(n14522));
  jand g14235(.dina(n14522), .dinb(n14521), .dout(n14523));
  jor  g14236(.dina(n14523), .dinb(n14520), .dout(n14524));
  jnot g14237(.din(n13968), .dout(n14525));
  jand g14238(.dina(n14522), .dinb(n14525), .dout(n14526));
  jnot g14239(.din(n14526), .dout(n14527));
  jand g14240(.dina(n14527), .dinb(n14524), .dout(n14528));
  jand g14241(.dina(n14528), .dinb(n14519), .dout(n14529));
  jor  g14242(.dina(n14529), .dinb(n14517), .dout(n14530));
  jand g14243(.dina(n14530), .dinb(asqrt[39] ), .dout(n14531));
  jxor g14244(.dina(n13969), .dinb(n3907), .dout(n14532));
  jand g14245(.dina(n14532), .dinb(asqrt[12] ), .dout(n14533));
  jxor g14246(.dina(n14533), .dinb(n13979), .dout(n14534));
  jnot g14247(.din(n14534), .dout(n14535));
  jor  g14248(.dina(n14530), .dinb(asqrt[39] ), .dout(n14536));
  jand g14249(.dina(n14536), .dinb(n14535), .dout(n14537));
  jor  g14250(.dina(n14537), .dinb(n14531), .dout(n14538));
  jand g14251(.dina(n14538), .dinb(asqrt[40] ), .dout(n14539));
  jnot g14252(.din(n13984), .dout(n14540));
  jand g14253(.dina(n14540), .dinb(n13982), .dout(n14541));
  jand g14254(.dina(n14541), .dinb(asqrt[12] ), .dout(n14542));
  jxor g14255(.dina(n14542), .dinb(n13992), .dout(n14543));
  jnot g14256(.din(n14543), .dout(n14544));
  jor  g14257(.dina(n14531), .dinb(asqrt[40] ), .dout(n14545));
  jor  g14258(.dina(n14545), .dinb(n14537), .dout(n14546));
  jand g14259(.dina(n14546), .dinb(n14544), .dout(n14547));
  jor  g14260(.dina(n14547), .dinb(n14539), .dout(n14548));
  jand g14261(.dina(n14548), .dinb(asqrt[41] ), .dout(n14549));
  jor  g14262(.dina(n14548), .dinb(asqrt[41] ), .dout(n14550));
  jnot g14263(.din(n13998), .dout(n14551));
  jnot g14264(.din(n13999), .dout(n14552));
  jand g14265(.dina(asqrt[12] ), .dinb(n13995), .dout(n14553));
  jand g14266(.dina(n14553), .dinb(n14552), .dout(n14554));
  jor  g14267(.dina(n14554), .dinb(n14551), .dout(n14555));
  jnot g14268(.din(n14000), .dout(n14556));
  jand g14269(.dina(n14553), .dinb(n14556), .dout(n14557));
  jnot g14270(.din(n14557), .dout(n14558));
  jand g14271(.dina(n14558), .dinb(n14555), .dout(n14559));
  jand g14272(.dina(n14559), .dinb(n14550), .dout(n14560));
  jor  g14273(.dina(n14560), .dinb(n14549), .dout(n14561));
  jand g14274(.dina(n14561), .dinb(asqrt[42] ), .dout(n14562));
  jor  g14275(.dina(n14549), .dinb(asqrt[42] ), .dout(n14563));
  jor  g14276(.dina(n14563), .dinb(n14560), .dout(n14564));
  jnot g14277(.din(n14006), .dout(n14565));
  jnot g14278(.din(n14008), .dout(n14566));
  jand g14279(.dina(asqrt[12] ), .dinb(n14002), .dout(n14567));
  jand g14280(.dina(n14567), .dinb(n14566), .dout(n14568));
  jor  g14281(.dina(n14568), .dinb(n14565), .dout(n14569));
  jnot g14282(.din(n14009), .dout(n14570));
  jand g14283(.dina(n14567), .dinb(n14570), .dout(n14571));
  jnot g14284(.din(n14571), .dout(n14572));
  jand g14285(.dina(n14572), .dinb(n14569), .dout(n14573));
  jand g14286(.dina(n14573), .dinb(n14564), .dout(n14574));
  jor  g14287(.dina(n14574), .dinb(n14562), .dout(n14575));
  jand g14288(.dina(n14575), .dinb(asqrt[43] ), .dout(n14576));
  jxor g14289(.dina(n14010), .dinb(n2870), .dout(n14577));
  jand g14290(.dina(n14577), .dinb(asqrt[12] ), .dout(n14578));
  jxor g14291(.dina(n14578), .dinb(n14020), .dout(n14579));
  jnot g14292(.din(n14579), .dout(n14580));
  jor  g14293(.dina(n14575), .dinb(asqrt[43] ), .dout(n14581));
  jand g14294(.dina(n14581), .dinb(n14580), .dout(n14582));
  jor  g14295(.dina(n14582), .dinb(n14576), .dout(n14583));
  jand g14296(.dina(n14583), .dinb(asqrt[44] ), .dout(n14584));
  jnot g14297(.din(n14025), .dout(n14585));
  jand g14298(.dina(n14585), .dinb(n14023), .dout(n14586));
  jand g14299(.dina(n14586), .dinb(asqrt[12] ), .dout(n14587));
  jxor g14300(.dina(n14587), .dinb(n14033), .dout(n14588));
  jnot g14301(.din(n14588), .dout(n14589));
  jor  g14302(.dina(n14576), .dinb(asqrt[44] ), .dout(n14590));
  jor  g14303(.dina(n14590), .dinb(n14582), .dout(n14591));
  jand g14304(.dina(n14591), .dinb(n14589), .dout(n14592));
  jor  g14305(.dina(n14592), .dinb(n14584), .dout(n14593));
  jand g14306(.dina(n14593), .dinb(asqrt[45] ), .dout(n14594));
  jor  g14307(.dina(n14593), .dinb(asqrt[45] ), .dout(n14595));
  jnot g14308(.din(n14039), .dout(n14596));
  jnot g14309(.din(n14040), .dout(n14597));
  jand g14310(.dina(asqrt[12] ), .dinb(n14036), .dout(n14598));
  jand g14311(.dina(n14598), .dinb(n14597), .dout(n14599));
  jor  g14312(.dina(n14599), .dinb(n14596), .dout(n14600));
  jnot g14313(.din(n14041), .dout(n14601));
  jand g14314(.dina(n14598), .dinb(n14601), .dout(n14602));
  jnot g14315(.din(n14602), .dout(n14603));
  jand g14316(.dina(n14603), .dinb(n14600), .dout(n14604));
  jand g14317(.dina(n14604), .dinb(n14595), .dout(n14605));
  jor  g14318(.dina(n14605), .dinb(n14594), .dout(n14606));
  jand g14319(.dina(n14606), .dinb(asqrt[46] ), .dout(n14607));
  jor  g14320(.dina(n14594), .dinb(asqrt[46] ), .dout(n14608));
  jor  g14321(.dina(n14608), .dinb(n14605), .dout(n14609));
  jnot g14322(.din(n14047), .dout(n14610));
  jnot g14323(.din(n14049), .dout(n14611));
  jand g14324(.dina(asqrt[12] ), .dinb(n14043), .dout(n14612));
  jand g14325(.dina(n14612), .dinb(n14611), .dout(n14613));
  jor  g14326(.dina(n14613), .dinb(n14610), .dout(n14614));
  jnot g14327(.din(n14050), .dout(n14615));
  jand g14328(.dina(n14612), .dinb(n14615), .dout(n14616));
  jnot g14329(.din(n14616), .dout(n14617));
  jand g14330(.dina(n14617), .dinb(n14614), .dout(n14618));
  jand g14331(.dina(n14618), .dinb(n14609), .dout(n14619));
  jor  g14332(.dina(n14619), .dinb(n14607), .dout(n14620));
  jand g14333(.dina(n14620), .dinb(asqrt[47] ), .dout(n14621));
  jxor g14334(.dina(n14051), .dinb(n2005), .dout(n14622));
  jand g14335(.dina(n14622), .dinb(asqrt[12] ), .dout(n14623));
  jxor g14336(.dina(n14623), .dinb(n14061), .dout(n14624));
  jnot g14337(.din(n14624), .dout(n14625));
  jor  g14338(.dina(n14620), .dinb(asqrt[47] ), .dout(n14626));
  jand g14339(.dina(n14626), .dinb(n14625), .dout(n14627));
  jor  g14340(.dina(n14627), .dinb(n14621), .dout(n14628));
  jand g14341(.dina(n14628), .dinb(asqrt[48] ), .dout(n14629));
  jnot g14342(.din(n14066), .dout(n14630));
  jand g14343(.dina(n14630), .dinb(n14064), .dout(n14631));
  jand g14344(.dina(n14631), .dinb(asqrt[12] ), .dout(n14632));
  jxor g14345(.dina(n14632), .dinb(n14074), .dout(n14633));
  jnot g14346(.din(n14633), .dout(n14634));
  jor  g14347(.dina(n14621), .dinb(asqrt[48] ), .dout(n14635));
  jor  g14348(.dina(n14635), .dinb(n14627), .dout(n14636));
  jand g14349(.dina(n14636), .dinb(n14634), .dout(n14637));
  jor  g14350(.dina(n14637), .dinb(n14629), .dout(n14638));
  jand g14351(.dina(n14638), .dinb(asqrt[49] ), .dout(n14639));
  jor  g14352(.dina(n14638), .dinb(asqrt[49] ), .dout(n14640));
  jnot g14353(.din(n14080), .dout(n14641));
  jnot g14354(.din(n14081), .dout(n14642));
  jand g14355(.dina(asqrt[12] ), .dinb(n14077), .dout(n14643));
  jand g14356(.dina(n14643), .dinb(n14642), .dout(n14644));
  jor  g14357(.dina(n14644), .dinb(n14641), .dout(n14645));
  jnot g14358(.din(n14082), .dout(n14646));
  jand g14359(.dina(n14643), .dinb(n14646), .dout(n14647));
  jnot g14360(.din(n14647), .dout(n14648));
  jand g14361(.dina(n14648), .dinb(n14645), .dout(n14649));
  jand g14362(.dina(n14649), .dinb(n14640), .dout(n14650));
  jor  g14363(.dina(n14650), .dinb(n14639), .dout(n14651));
  jand g14364(.dina(n14651), .dinb(asqrt[50] ), .dout(n14652));
  jnot g14365(.din(n14086), .dout(n14653));
  jand g14366(.dina(n14653), .dinb(n14084), .dout(n14654));
  jand g14367(.dina(n14654), .dinb(asqrt[12] ), .dout(n14655));
  jxor g14368(.dina(n14655), .dinb(n14094), .dout(n14656));
  jnot g14369(.din(n14656), .dout(n14657));
  jor  g14370(.dina(n14639), .dinb(asqrt[50] ), .dout(n14658));
  jor  g14371(.dina(n14658), .dinb(n14650), .dout(n14659));
  jand g14372(.dina(n14659), .dinb(n14657), .dout(n14660));
  jor  g14373(.dina(n14660), .dinb(n14652), .dout(n14661));
  jand g14374(.dina(n14661), .dinb(asqrt[51] ), .dout(n14662));
  jnot g14375(.din(n14246), .dout(n14663));
  jor  g14376(.dina(n14661), .dinb(asqrt[51] ), .dout(n14664));
  jand g14377(.dina(n14664), .dinb(n14663), .dout(n14665));
  jor  g14378(.dina(n14665), .dinb(n14662), .dout(n14666));
  jand g14379(.dina(n14666), .dinb(asqrt[52] ), .dout(n14667));
  jor  g14380(.dina(n14662), .dinb(asqrt[52] ), .dout(n14668));
  jor  g14381(.dina(n14668), .dinb(n14665), .dout(n14669));
  jnot g14382(.din(n14105), .dout(n14670));
  jnot g14383(.din(n14107), .dout(n14671));
  jand g14384(.dina(asqrt[12] ), .dinb(n14101), .dout(n14672));
  jand g14385(.dina(n14672), .dinb(n14671), .dout(n14673));
  jor  g14386(.dina(n14673), .dinb(n14670), .dout(n14674));
  jnot g14387(.din(n14108), .dout(n14675));
  jand g14388(.dina(n14672), .dinb(n14675), .dout(n14676));
  jnot g14389(.din(n14676), .dout(n14677));
  jand g14390(.dina(n14677), .dinb(n14674), .dout(n14678));
  jand g14391(.dina(n14678), .dinb(n14669), .dout(n14679));
  jor  g14392(.dina(n14679), .dinb(n14667), .dout(n14680));
  jand g14393(.dina(n14680), .dinb(asqrt[53] ), .dout(n14681));
  jor  g14394(.dina(n14680), .dinb(asqrt[53] ), .dout(n14682));
  jnot g14395(.din(n14113), .dout(n14683));
  jnot g14396(.din(n14114), .dout(n14684));
  jand g14397(.dina(asqrt[12] ), .dinb(n14110), .dout(n14685));
  jand g14398(.dina(n14685), .dinb(n14684), .dout(n14686));
  jor  g14399(.dina(n14686), .dinb(n14683), .dout(n14687));
  jnot g14400(.din(n14115), .dout(n14688));
  jand g14401(.dina(n14685), .dinb(n14688), .dout(n14689));
  jnot g14402(.din(n14689), .dout(n14690));
  jand g14403(.dina(n14690), .dinb(n14687), .dout(n14691));
  jand g14404(.dina(n14691), .dinb(n14682), .dout(n14692));
  jor  g14405(.dina(n14692), .dinb(n14681), .dout(n14693));
  jand g14406(.dina(n14693), .dinb(asqrt[54] ), .dout(n14694));
  jor  g14407(.dina(n14681), .dinb(asqrt[54] ), .dout(n14695));
  jor  g14408(.dina(n14695), .dinb(n14692), .dout(n14696));
  jnot g14409(.din(n14121), .dout(n14697));
  jnot g14410(.din(n14123), .dout(n14698));
  jand g14411(.dina(asqrt[12] ), .dinb(n14117), .dout(n14699));
  jand g14412(.dina(n14699), .dinb(n14698), .dout(n14700));
  jor  g14413(.dina(n14700), .dinb(n14697), .dout(n14701));
  jnot g14414(.din(n14124), .dout(n14702));
  jand g14415(.dina(n14699), .dinb(n14702), .dout(n14703));
  jnot g14416(.din(n14703), .dout(n14704));
  jand g14417(.dina(n14704), .dinb(n14701), .dout(n14705));
  jand g14418(.dina(n14705), .dinb(n14696), .dout(n14706));
  jor  g14419(.dina(n14706), .dinb(n14694), .dout(n14707));
  jand g14420(.dina(n14707), .dinb(asqrt[55] ), .dout(n14708));
  jxor g14421(.dina(n14125), .dinb(n791), .dout(n14709));
  jand g14422(.dina(n14709), .dinb(asqrt[12] ), .dout(n14710));
  jxor g14423(.dina(n14710), .dinb(n14135), .dout(n14711));
  jnot g14424(.din(n14711), .dout(n14712));
  jor  g14425(.dina(n14707), .dinb(asqrt[55] ), .dout(n14713));
  jand g14426(.dina(n14713), .dinb(n14712), .dout(n14714));
  jor  g14427(.dina(n14714), .dinb(n14708), .dout(n14715));
  jand g14428(.dina(n14715), .dinb(asqrt[56] ), .dout(n14716));
  jnot g14429(.din(n14140), .dout(n14717));
  jand g14430(.dina(n14717), .dinb(n14138), .dout(n14718));
  jand g14431(.dina(n14718), .dinb(asqrt[12] ), .dout(n14719));
  jxor g14432(.dina(n14719), .dinb(n14148), .dout(n14720));
  jnot g14433(.din(n14720), .dout(n14721));
  jor  g14434(.dina(n14708), .dinb(asqrt[56] ), .dout(n14722));
  jor  g14435(.dina(n14722), .dinb(n14714), .dout(n14723));
  jand g14436(.dina(n14723), .dinb(n14721), .dout(n14724));
  jor  g14437(.dina(n14724), .dinb(n14716), .dout(n14725));
  jand g14438(.dina(n14725), .dinb(asqrt[57] ), .dout(n14726));
  jor  g14439(.dina(n14725), .dinb(asqrt[57] ), .dout(n14727));
  jnot g14440(.din(n14154), .dout(n14728));
  jnot g14441(.din(n14155), .dout(n14729));
  jand g14442(.dina(asqrt[12] ), .dinb(n14151), .dout(n14730));
  jand g14443(.dina(n14730), .dinb(n14729), .dout(n14731));
  jor  g14444(.dina(n14731), .dinb(n14728), .dout(n14732));
  jnot g14445(.din(n14156), .dout(n14733));
  jand g14446(.dina(n14730), .dinb(n14733), .dout(n14734));
  jnot g14447(.din(n14734), .dout(n14735));
  jand g14448(.dina(n14735), .dinb(n14732), .dout(n14736));
  jand g14449(.dina(n14736), .dinb(n14727), .dout(n14737));
  jor  g14450(.dina(n14737), .dinb(n14726), .dout(n14738));
  jand g14451(.dina(n14738), .dinb(asqrt[58] ), .dout(n14739));
  jor  g14452(.dina(n14726), .dinb(asqrt[58] ), .dout(n14740));
  jor  g14453(.dina(n14740), .dinb(n14737), .dout(n14741));
  jnot g14454(.din(n14162), .dout(n14742));
  jnot g14455(.din(n14164), .dout(n14743));
  jand g14456(.dina(asqrt[12] ), .dinb(n14158), .dout(n14744));
  jand g14457(.dina(n14744), .dinb(n14743), .dout(n14745));
  jor  g14458(.dina(n14745), .dinb(n14742), .dout(n14746));
  jnot g14459(.din(n14165), .dout(n14747));
  jand g14460(.dina(n14744), .dinb(n14747), .dout(n14748));
  jnot g14461(.din(n14748), .dout(n14749));
  jand g14462(.dina(n14749), .dinb(n14746), .dout(n14750));
  jand g14463(.dina(n14750), .dinb(n14741), .dout(n14751));
  jor  g14464(.dina(n14751), .dinb(n14739), .dout(n14752));
  jand g14465(.dina(n14752), .dinb(asqrt[59] ), .dout(n14753));
  jxor g14466(.dina(n14166), .dinb(n425), .dout(n14754));
  jand g14467(.dina(n14754), .dinb(asqrt[12] ), .dout(n14755));
  jxor g14468(.dina(n14755), .dinb(n14176), .dout(n14756));
  jnot g14469(.din(n14756), .dout(n14757));
  jor  g14470(.dina(n14752), .dinb(asqrt[59] ), .dout(n14758));
  jand g14471(.dina(n14758), .dinb(n14757), .dout(n14759));
  jor  g14472(.dina(n14759), .dinb(n14753), .dout(n14760));
  jand g14473(.dina(n14760), .dinb(asqrt[60] ), .dout(n14761));
  jnot g14474(.din(n14181), .dout(n14762));
  jand g14475(.dina(n14762), .dinb(n14179), .dout(n14763));
  jand g14476(.dina(n14763), .dinb(asqrt[12] ), .dout(n14764));
  jxor g14477(.dina(n14764), .dinb(n14189), .dout(n14765));
  jnot g14478(.din(n14765), .dout(n14766));
  jor  g14479(.dina(n14753), .dinb(asqrt[60] ), .dout(n14767));
  jor  g14480(.dina(n14767), .dinb(n14759), .dout(n14768));
  jand g14481(.dina(n14768), .dinb(n14766), .dout(n14769));
  jor  g14482(.dina(n14769), .dinb(n14761), .dout(n14770));
  jand g14483(.dina(n14770), .dinb(asqrt[61] ), .dout(n14771));
  jor  g14484(.dina(n14770), .dinb(asqrt[61] ), .dout(n14772));
  jnot g14485(.din(n14195), .dout(n14773));
  jnot g14486(.din(n14196), .dout(n14774));
  jand g14487(.dina(asqrt[12] ), .dinb(n14192), .dout(n14775));
  jand g14488(.dina(n14775), .dinb(n14774), .dout(n14776));
  jor  g14489(.dina(n14776), .dinb(n14773), .dout(n14777));
  jnot g14490(.din(n14197), .dout(n14778));
  jand g14491(.dina(n14775), .dinb(n14778), .dout(n14779));
  jnot g14492(.din(n14779), .dout(n14780));
  jand g14493(.dina(n14780), .dinb(n14777), .dout(n14781));
  jand g14494(.dina(n14781), .dinb(n14772), .dout(n14782));
  jor  g14495(.dina(n14782), .dinb(n14771), .dout(n14783));
  jand g14496(.dina(n14783), .dinb(asqrt[62] ), .dout(n14784));
  jor  g14497(.dina(n14771), .dinb(asqrt[62] ), .dout(n14785));
  jor  g14498(.dina(n14785), .dinb(n14782), .dout(n14786));
  jnot g14499(.din(n14203), .dout(n14787));
  jnot g14500(.din(n14205), .dout(n14788));
  jand g14501(.dina(asqrt[12] ), .dinb(n14199), .dout(n14789));
  jand g14502(.dina(n14789), .dinb(n14788), .dout(n14790));
  jor  g14503(.dina(n14790), .dinb(n14787), .dout(n14791));
  jnot g14504(.din(n14206), .dout(n14792));
  jand g14505(.dina(n14789), .dinb(n14792), .dout(n14793));
  jnot g14506(.din(n14793), .dout(n14794));
  jand g14507(.dina(n14794), .dinb(n14791), .dout(n14795));
  jand g14508(.dina(n14795), .dinb(n14786), .dout(n14796));
  jor  g14509(.dina(n14796), .dinb(n14784), .dout(n14797));
  jxor g14510(.dina(n14207), .dinb(n199), .dout(n14798));
  jand g14511(.dina(n14798), .dinb(asqrt[12] ), .dout(n14799));
  jxor g14512(.dina(n14799), .dinb(n14217), .dout(n14800));
  jnot g14513(.din(n14219), .dout(n14801));
  jand g14514(.dina(asqrt[12] ), .dinb(n14226), .dout(n14802));
  jand g14515(.dina(n14802), .dinb(n14801), .dout(n14803));
  jor  g14516(.dina(n14803), .dinb(n14234), .dout(n14804));
  jor  g14517(.dina(n14804), .dinb(n14800), .dout(n14805));
  jnot g14518(.din(n14805), .dout(n14806));
  jand g14519(.dina(n14806), .dinb(n14797), .dout(n14807));
  jor  g14520(.dina(n14807), .dinb(asqrt[63] ), .dout(n14808));
  jnot g14521(.din(n14800), .dout(n14809));
  jor  g14522(.dina(n14809), .dinb(n14797), .dout(n14810));
  jor  g14523(.dina(n14802), .dinb(n14801), .dout(n14811));
  jand g14524(.dina(n14226), .dinb(n14801), .dout(n14812));
  jor  g14525(.dina(n14812), .dinb(n194), .dout(n14813));
  jnot g14526(.din(n14813), .dout(n14814));
  jand g14527(.dina(n14814), .dinb(n14811), .dout(n14815));
  jnot g14528(.din(asqrt[12] ), .dout(n14816));
  jnot g14529(.din(n14815), .dout(n14819));
  jand g14530(.dina(n14819), .dinb(n14810), .dout(n14820));
  jand g14531(.dina(n14820), .dinb(n14808), .dout(n14821));
  jxor g14532(.dina(n14661), .dinb(n1039), .dout(n14822));
  jor  g14533(.dina(n14822), .dinb(n14821), .dout(n14823));
  jxor g14534(.dina(n14823), .dinb(n14246), .dout(n14824));
  jor  g14535(.dina(n14821), .dinb(n14248), .dout(n14825));
  jnot g14536(.din(a[20] ), .dout(n14826));
  jnot g14537(.din(a[21] ), .dout(n14827));
  jand g14538(.dina(n14248), .dinb(n14827), .dout(n14828));
  jand g14539(.dina(n14828), .dinb(n14826), .dout(n14829));
  jnot g14540(.din(n14829), .dout(n14830));
  jand g14541(.dina(n14830), .dinb(n14825), .dout(n14831));
  jor  g14542(.dina(n14831), .dinb(n14816), .dout(n14832));
  jor  g14543(.dina(n14821), .dinb(a[22] ), .dout(n14833));
  jxor g14544(.dina(n14833), .dinb(n14249), .dout(n14834));
  jand g14545(.dina(n14831), .dinb(n14816), .dout(n14835));
  jor  g14546(.dina(n14835), .dinb(n14834), .dout(n14836));
  jand g14547(.dina(n14836), .dinb(n14832), .dout(n14837));
  jor  g14548(.dina(n14837), .dinb(n13723), .dout(n14838));
  jand g14549(.dina(n14832), .dinb(n13723), .dout(n14839));
  jand g14550(.dina(n14839), .dinb(n14836), .dout(n14840));
  jor  g14551(.dina(n14833), .dinb(a[23] ), .dout(n14841));
  jnot g14552(.din(n14808), .dout(n14842));
  jnot g14553(.din(n14810), .dout(n14843));
  jor  g14554(.dina(n14815), .dinb(n14816), .dout(n14844));
  jor  g14555(.dina(n14844), .dinb(n14843), .dout(n14845));
  jor  g14556(.dina(n14845), .dinb(n14842), .dout(n14846));
  jand g14557(.dina(n14846), .dinb(n14841), .dout(n14847));
  jxor g14558(.dina(n14847), .dinb(n13728), .dout(n14848));
  jor  g14559(.dina(n14848), .dinb(n14840), .dout(n14849));
  jand g14560(.dina(n14849), .dinb(n14838), .dout(n14850));
  jor  g14561(.dina(n14850), .dinb(n13718), .dout(n14851));
  jand g14562(.dina(n14850), .dinb(n13718), .dout(n14852));
  jxor g14563(.dina(n14252), .dinb(n13723), .dout(n14853));
  jor  g14564(.dina(n14853), .dinb(n14821), .dout(n14854));
  jxor g14565(.dina(n14854), .dinb(n14255), .dout(n14855));
  jor  g14566(.dina(n14855), .dinb(n14852), .dout(n14856));
  jand g14567(.dina(n14856), .dinb(n14851), .dout(n14857));
  jor  g14568(.dina(n14857), .dinb(n12675), .dout(n14858));
  jnot g14569(.din(n14261), .dout(n14859));
  jor  g14570(.dina(n14859), .dinb(n14259), .dout(n14860));
  jor  g14571(.dina(n14860), .dinb(n14821), .dout(n14861));
  jxor g14572(.dina(n14861), .dinb(n14270), .dout(n14862));
  jand g14573(.dina(n14851), .dinb(n12675), .dout(n14863));
  jand g14574(.dina(n14863), .dinb(n14856), .dout(n14864));
  jor  g14575(.dina(n14864), .dinb(n14862), .dout(n14865));
  jand g14576(.dina(n14865), .dinb(n14858), .dout(n14866));
  jor  g14577(.dina(n14866), .dinb(n12670), .dout(n14867));
  jand g14578(.dina(n14866), .dinb(n12670), .dout(n14868));
  jxor g14579(.dina(n14272), .dinb(n12675), .dout(n14869));
  jor  g14580(.dina(n14869), .dinb(n14821), .dout(n14870));
  jxor g14581(.dina(n14870), .dinb(n14277), .dout(n14871));
  jnot g14582(.din(n14871), .dout(n14872));
  jor  g14583(.dina(n14872), .dinb(n14868), .dout(n14873));
  jand g14584(.dina(n14873), .dinb(n14867), .dout(n14874));
  jor  g14585(.dina(n14874), .dinb(n11662), .dout(n14875));
  jand g14586(.dina(n14867), .dinb(n11662), .dout(n14876));
  jand g14587(.dina(n14876), .dinb(n14873), .dout(n14877));
  jnot g14588(.din(n14281), .dout(n14878));
  jnot g14589(.din(n14821), .dout(asqrt[11] ));
  jand g14590(.dina(asqrt[11] ), .dinb(n14878), .dout(n14880));
  jand g14591(.dina(n14880), .dinb(n14288), .dout(n14881));
  jor  g14592(.dina(n14881), .dinb(n14286), .dout(n14882));
  jand g14593(.dina(n14880), .dinb(n14289), .dout(n14883));
  jnot g14594(.din(n14883), .dout(n14884));
  jand g14595(.dina(n14884), .dinb(n14882), .dout(n14885));
  jnot g14596(.din(n14885), .dout(n14886));
  jor  g14597(.dina(n14886), .dinb(n14877), .dout(n14887));
  jand g14598(.dina(n14887), .dinb(n14875), .dout(n14888));
  jor  g14599(.dina(n14888), .dinb(n11657), .dout(n14889));
  jand g14600(.dina(n14888), .dinb(n11657), .dout(n14890));
  jnot g14601(.din(n14296), .dout(n14891));
  jxor g14602(.dina(n14290), .dinb(n11662), .dout(n14892));
  jor  g14603(.dina(n14892), .dinb(n14821), .dout(n14893));
  jxor g14604(.dina(n14893), .dinb(n14891), .dout(n14894));
  jnot g14605(.din(n14894), .dout(n14895));
  jor  g14606(.dina(n14895), .dinb(n14890), .dout(n14896));
  jand g14607(.dina(n14896), .dinb(n14889), .dout(n14897));
  jor  g14608(.dina(n14897), .dinb(n10701), .dout(n14898));
  jnot g14609(.din(n14301), .dout(n14899));
  jor  g14610(.dina(n14899), .dinb(n14299), .dout(n14900));
  jor  g14611(.dina(n14900), .dinb(n14821), .dout(n14901));
  jxor g14612(.dina(n14901), .dinb(n14310), .dout(n14902));
  jand g14613(.dina(n14889), .dinb(n10701), .dout(n14903));
  jand g14614(.dina(n14903), .dinb(n14896), .dout(n14904));
  jor  g14615(.dina(n14904), .dinb(n14902), .dout(n14905));
  jand g14616(.dina(n14905), .dinb(n14898), .dout(n14906));
  jor  g14617(.dina(n14906), .dinb(n10696), .dout(n14907));
  jand g14618(.dina(n14906), .dinb(n10696), .dout(n14908));
  jnot g14619(.din(n14317), .dout(n14909));
  jxor g14620(.dina(n14312), .dinb(n10701), .dout(n14910));
  jor  g14621(.dina(n14910), .dinb(n14821), .dout(n14911));
  jxor g14622(.dina(n14911), .dinb(n14909), .dout(n14912));
  jnot g14623(.din(n14912), .dout(n14913));
  jor  g14624(.dina(n14913), .dinb(n14908), .dout(n14914));
  jand g14625(.dina(n14914), .dinb(n14907), .dout(n14915));
  jor  g14626(.dina(n14915), .dinb(n9774), .dout(n14916));
  jand g14627(.dina(n14907), .dinb(n9774), .dout(n14917));
  jand g14628(.dina(n14917), .dinb(n14914), .dout(n14918));
  jnot g14629(.din(n14320), .dout(n14919));
  jand g14630(.dina(asqrt[11] ), .dinb(n14919), .dout(n14920));
  jand g14631(.dina(n14920), .dinb(n14327), .dout(n14921));
  jor  g14632(.dina(n14921), .dinb(n14325), .dout(n14922));
  jand g14633(.dina(n14920), .dinb(n14328), .dout(n14923));
  jnot g14634(.din(n14923), .dout(n14924));
  jand g14635(.dina(n14924), .dinb(n14922), .dout(n14925));
  jnot g14636(.din(n14925), .dout(n14926));
  jor  g14637(.dina(n14926), .dinb(n14918), .dout(n14927));
  jand g14638(.dina(n14927), .dinb(n14916), .dout(n14928));
  jor  g14639(.dina(n14928), .dinb(n9769), .dout(n14929));
  jxor g14640(.dina(n14329), .dinb(n9774), .dout(n14930));
  jor  g14641(.dina(n14930), .dinb(n14821), .dout(n14931));
  jxor g14642(.dina(n14931), .dinb(n14334), .dout(n14932));
  jand g14643(.dina(n14928), .dinb(n9769), .dout(n14933));
  jor  g14644(.dina(n14933), .dinb(n14932), .dout(n14934));
  jand g14645(.dina(n14934), .dinb(n14929), .dout(n14935));
  jor  g14646(.dina(n14935), .dinb(n8898), .dout(n14936));
  jnot g14647(.din(n14339), .dout(n14937));
  jor  g14648(.dina(n14937), .dinb(n14337), .dout(n14938));
  jor  g14649(.dina(n14938), .dinb(n14821), .dout(n14939));
  jxor g14650(.dina(n14939), .dinb(n14348), .dout(n14940));
  jand g14651(.dina(n14929), .dinb(n8898), .dout(n14941));
  jand g14652(.dina(n14941), .dinb(n14934), .dout(n14942));
  jor  g14653(.dina(n14942), .dinb(n14940), .dout(n14943));
  jand g14654(.dina(n14943), .dinb(n14936), .dout(n14944));
  jor  g14655(.dina(n14944), .dinb(n8893), .dout(n14945));
  jand g14656(.dina(n14944), .dinb(n8893), .dout(n14946));
  jnot g14657(.din(n14351), .dout(n14947));
  jand g14658(.dina(asqrt[11] ), .dinb(n14947), .dout(n14948));
  jand g14659(.dina(n14948), .dinb(n14356), .dout(n14949));
  jor  g14660(.dina(n14949), .dinb(n14355), .dout(n14950));
  jand g14661(.dina(n14948), .dinb(n14357), .dout(n14951));
  jnot g14662(.din(n14951), .dout(n14952));
  jand g14663(.dina(n14952), .dinb(n14950), .dout(n14953));
  jnot g14664(.din(n14953), .dout(n14954));
  jor  g14665(.dina(n14954), .dinb(n14946), .dout(n14955));
  jand g14666(.dina(n14955), .dinb(n14945), .dout(n14956));
  jor  g14667(.dina(n14956), .dinb(n8058), .dout(n14957));
  jand g14668(.dina(n14945), .dinb(n8058), .dout(n14958));
  jand g14669(.dina(n14958), .dinb(n14955), .dout(n14959));
  jnot g14670(.din(n14359), .dout(n14960));
  jand g14671(.dina(asqrt[11] ), .dinb(n14960), .dout(n14961));
  jand g14672(.dina(n14961), .dinb(n14366), .dout(n14962));
  jor  g14673(.dina(n14962), .dinb(n14364), .dout(n14963));
  jand g14674(.dina(n14961), .dinb(n14367), .dout(n14964));
  jnot g14675(.din(n14964), .dout(n14965));
  jand g14676(.dina(n14965), .dinb(n14963), .dout(n14966));
  jnot g14677(.din(n14966), .dout(n14967));
  jor  g14678(.dina(n14967), .dinb(n14959), .dout(n14968));
  jand g14679(.dina(n14968), .dinb(n14957), .dout(n14969));
  jor  g14680(.dina(n14969), .dinb(n8053), .dout(n14970));
  jxor g14681(.dina(n14368), .dinb(n8058), .dout(n14971));
  jor  g14682(.dina(n14971), .dinb(n14821), .dout(n14972));
  jxor g14683(.dina(n14972), .dinb(n14379), .dout(n14973));
  jand g14684(.dina(n14969), .dinb(n8053), .dout(n14974));
  jor  g14685(.dina(n14974), .dinb(n14973), .dout(n14975));
  jand g14686(.dina(n14975), .dinb(n14970), .dout(n14976));
  jor  g14687(.dina(n14976), .dinb(n7265), .dout(n14977));
  jnot g14688(.din(n14384), .dout(n14978));
  jor  g14689(.dina(n14978), .dinb(n14382), .dout(n14979));
  jor  g14690(.dina(n14979), .dinb(n14821), .dout(n14980));
  jxor g14691(.dina(n14980), .dinb(n14393), .dout(n14981));
  jand g14692(.dina(n14970), .dinb(n7265), .dout(n14982));
  jand g14693(.dina(n14982), .dinb(n14975), .dout(n14983));
  jor  g14694(.dina(n14983), .dinb(n14981), .dout(n14984));
  jand g14695(.dina(n14984), .dinb(n14977), .dout(n14985));
  jor  g14696(.dina(n14985), .dinb(n7260), .dout(n14986));
  jand g14697(.dina(n14985), .dinb(n7260), .dout(n14987));
  jnot g14698(.din(n14396), .dout(n14988));
  jand g14699(.dina(asqrt[11] ), .dinb(n14988), .dout(n14989));
  jand g14700(.dina(n14989), .dinb(n14401), .dout(n14990));
  jor  g14701(.dina(n14990), .dinb(n14400), .dout(n14991));
  jand g14702(.dina(n14989), .dinb(n14402), .dout(n14992));
  jnot g14703(.din(n14992), .dout(n14993));
  jand g14704(.dina(n14993), .dinb(n14991), .dout(n14994));
  jnot g14705(.din(n14994), .dout(n14995));
  jor  g14706(.dina(n14995), .dinb(n14987), .dout(n14996));
  jand g14707(.dina(n14996), .dinb(n14986), .dout(n14997));
  jor  g14708(.dina(n14997), .dinb(n6505), .dout(n14998));
  jand g14709(.dina(n14986), .dinb(n6505), .dout(n14999));
  jand g14710(.dina(n14999), .dinb(n14996), .dout(n15000));
  jnot g14711(.din(n14404), .dout(n15001));
  jand g14712(.dina(asqrt[11] ), .dinb(n15001), .dout(n15002));
  jand g14713(.dina(n15002), .dinb(n14411), .dout(n15003));
  jor  g14714(.dina(n15003), .dinb(n14409), .dout(n15004));
  jand g14715(.dina(n15002), .dinb(n14412), .dout(n15005));
  jnot g14716(.din(n15005), .dout(n15006));
  jand g14717(.dina(n15006), .dinb(n15004), .dout(n15007));
  jnot g14718(.din(n15007), .dout(n15008));
  jor  g14719(.dina(n15008), .dinb(n15000), .dout(n15009));
  jand g14720(.dina(n15009), .dinb(n14998), .dout(n15010));
  jor  g14721(.dina(n15010), .dinb(n6500), .dout(n15011));
  jxor g14722(.dina(n14413), .dinb(n6505), .dout(n15012));
  jor  g14723(.dina(n15012), .dinb(n14821), .dout(n15013));
  jxor g14724(.dina(n15013), .dinb(n14424), .dout(n15014));
  jand g14725(.dina(n15010), .dinb(n6500), .dout(n15015));
  jor  g14726(.dina(n15015), .dinb(n15014), .dout(n15016));
  jand g14727(.dina(n15016), .dinb(n15011), .dout(n15017));
  jor  g14728(.dina(n15017), .dinb(n5793), .dout(n15018));
  jnot g14729(.din(n14429), .dout(n15019));
  jor  g14730(.dina(n15019), .dinb(n14427), .dout(n15020));
  jor  g14731(.dina(n15020), .dinb(n14821), .dout(n15021));
  jxor g14732(.dina(n15021), .dinb(n14438), .dout(n15022));
  jand g14733(.dina(n15011), .dinb(n5793), .dout(n15023));
  jand g14734(.dina(n15023), .dinb(n15016), .dout(n15024));
  jor  g14735(.dina(n15024), .dinb(n15022), .dout(n15025));
  jand g14736(.dina(n15025), .dinb(n15018), .dout(n15026));
  jor  g14737(.dina(n15026), .dinb(n5788), .dout(n15027));
  jand g14738(.dina(n15026), .dinb(n5788), .dout(n15028));
  jnot g14739(.din(n14441), .dout(n15029));
  jand g14740(.dina(asqrt[11] ), .dinb(n15029), .dout(n15030));
  jand g14741(.dina(n15030), .dinb(n14446), .dout(n15031));
  jor  g14742(.dina(n15031), .dinb(n14445), .dout(n15032));
  jand g14743(.dina(n15030), .dinb(n14447), .dout(n15033));
  jnot g14744(.din(n15033), .dout(n15034));
  jand g14745(.dina(n15034), .dinb(n15032), .dout(n15035));
  jnot g14746(.din(n15035), .dout(n15036));
  jor  g14747(.dina(n15036), .dinb(n15028), .dout(n15037));
  jand g14748(.dina(n15037), .dinb(n15027), .dout(n15038));
  jor  g14749(.dina(n15038), .dinb(n5121), .dout(n15039));
  jand g14750(.dina(n15027), .dinb(n5121), .dout(n15040));
  jand g14751(.dina(n15040), .dinb(n15037), .dout(n15041));
  jnot g14752(.din(n14449), .dout(n15042));
  jand g14753(.dina(asqrt[11] ), .dinb(n15042), .dout(n15043));
  jand g14754(.dina(n15043), .dinb(n14456), .dout(n15044));
  jor  g14755(.dina(n15044), .dinb(n14454), .dout(n15045));
  jand g14756(.dina(n15043), .dinb(n14457), .dout(n15046));
  jnot g14757(.din(n15046), .dout(n15047));
  jand g14758(.dina(n15047), .dinb(n15045), .dout(n15048));
  jnot g14759(.din(n15048), .dout(n15049));
  jor  g14760(.dina(n15049), .dinb(n15041), .dout(n15050));
  jand g14761(.dina(n15050), .dinb(n15039), .dout(n15051));
  jor  g14762(.dina(n15051), .dinb(n5116), .dout(n15052));
  jxor g14763(.dina(n14458), .dinb(n5121), .dout(n15053));
  jor  g14764(.dina(n15053), .dinb(n14821), .dout(n15054));
  jxor g14765(.dina(n15054), .dinb(n14469), .dout(n15055));
  jand g14766(.dina(n15051), .dinb(n5116), .dout(n15056));
  jor  g14767(.dina(n15056), .dinb(n15055), .dout(n15057));
  jand g14768(.dina(n15057), .dinb(n15052), .dout(n15058));
  jor  g14769(.dina(n15058), .dinb(n4499), .dout(n15059));
  jnot g14770(.din(n14474), .dout(n15060));
  jor  g14771(.dina(n15060), .dinb(n14472), .dout(n15061));
  jor  g14772(.dina(n15061), .dinb(n14821), .dout(n15062));
  jxor g14773(.dina(n15062), .dinb(n14483), .dout(n15063));
  jand g14774(.dina(n15052), .dinb(n4499), .dout(n15064));
  jand g14775(.dina(n15064), .dinb(n15057), .dout(n15065));
  jor  g14776(.dina(n15065), .dinb(n15063), .dout(n15066));
  jand g14777(.dina(n15066), .dinb(n15059), .dout(n15067));
  jor  g14778(.dina(n15067), .dinb(n4494), .dout(n15068));
  jand g14779(.dina(n15067), .dinb(n4494), .dout(n15069));
  jnot g14780(.din(n14486), .dout(n15070));
  jand g14781(.dina(asqrt[11] ), .dinb(n15070), .dout(n15071));
  jand g14782(.dina(n15071), .dinb(n14491), .dout(n15072));
  jor  g14783(.dina(n15072), .dinb(n14490), .dout(n15073));
  jand g14784(.dina(n15071), .dinb(n14492), .dout(n15074));
  jnot g14785(.din(n15074), .dout(n15075));
  jand g14786(.dina(n15075), .dinb(n15073), .dout(n15076));
  jnot g14787(.din(n15076), .dout(n15077));
  jor  g14788(.dina(n15077), .dinb(n15069), .dout(n15078));
  jand g14789(.dina(n15078), .dinb(n15068), .dout(n15079));
  jor  g14790(.dina(n15079), .dinb(n3912), .dout(n15080));
  jand g14791(.dina(n15068), .dinb(n3912), .dout(n15081));
  jand g14792(.dina(n15081), .dinb(n15078), .dout(n15082));
  jnot g14793(.din(n14494), .dout(n15083));
  jand g14794(.dina(asqrt[11] ), .dinb(n15083), .dout(n15084));
  jand g14795(.dina(n15084), .dinb(n14501), .dout(n15085));
  jor  g14796(.dina(n15085), .dinb(n14499), .dout(n15086));
  jand g14797(.dina(n15084), .dinb(n14502), .dout(n15087));
  jnot g14798(.din(n15087), .dout(n15088));
  jand g14799(.dina(n15088), .dinb(n15086), .dout(n15089));
  jnot g14800(.din(n15089), .dout(n15090));
  jor  g14801(.dina(n15090), .dinb(n15082), .dout(n15091));
  jand g14802(.dina(n15091), .dinb(n15080), .dout(n15092));
  jor  g14803(.dina(n15092), .dinb(n3907), .dout(n15093));
  jxor g14804(.dina(n14503), .dinb(n3912), .dout(n15094));
  jor  g14805(.dina(n15094), .dinb(n14821), .dout(n15095));
  jxor g14806(.dina(n15095), .dinb(n14514), .dout(n15096));
  jand g14807(.dina(n15092), .dinb(n3907), .dout(n15097));
  jor  g14808(.dina(n15097), .dinb(n15096), .dout(n15098));
  jand g14809(.dina(n15098), .dinb(n15093), .dout(n15099));
  jor  g14810(.dina(n15099), .dinb(n3376), .dout(n15100));
  jnot g14811(.din(n14519), .dout(n15101));
  jor  g14812(.dina(n15101), .dinb(n14517), .dout(n15102));
  jor  g14813(.dina(n15102), .dinb(n14821), .dout(n15103));
  jxor g14814(.dina(n15103), .dinb(n14528), .dout(n15104));
  jand g14815(.dina(n15093), .dinb(n3376), .dout(n15105));
  jand g14816(.dina(n15105), .dinb(n15098), .dout(n15106));
  jor  g14817(.dina(n15106), .dinb(n15104), .dout(n15107));
  jand g14818(.dina(n15107), .dinb(n15100), .dout(n15108));
  jor  g14819(.dina(n15108), .dinb(n3371), .dout(n15109));
  jand g14820(.dina(n15108), .dinb(n3371), .dout(n15110));
  jnot g14821(.din(n14531), .dout(n15111));
  jand g14822(.dina(asqrt[11] ), .dinb(n15111), .dout(n15112));
  jand g14823(.dina(n15112), .dinb(n14536), .dout(n15113));
  jor  g14824(.dina(n15113), .dinb(n14535), .dout(n15114));
  jand g14825(.dina(n15112), .dinb(n14537), .dout(n15115));
  jnot g14826(.din(n15115), .dout(n15116));
  jand g14827(.dina(n15116), .dinb(n15114), .dout(n15117));
  jnot g14828(.din(n15117), .dout(n15118));
  jor  g14829(.dina(n15118), .dinb(n15110), .dout(n15119));
  jand g14830(.dina(n15119), .dinb(n15109), .dout(n15120));
  jor  g14831(.dina(n15120), .dinb(n2875), .dout(n15121));
  jand g14832(.dina(n15109), .dinb(n2875), .dout(n15122));
  jand g14833(.dina(n15122), .dinb(n15119), .dout(n15123));
  jnot g14834(.din(n14539), .dout(n15124));
  jand g14835(.dina(asqrt[11] ), .dinb(n15124), .dout(n15125));
  jand g14836(.dina(n15125), .dinb(n14546), .dout(n15126));
  jor  g14837(.dina(n15126), .dinb(n14544), .dout(n15127));
  jand g14838(.dina(n15125), .dinb(n14547), .dout(n15128));
  jnot g14839(.din(n15128), .dout(n15129));
  jand g14840(.dina(n15129), .dinb(n15127), .dout(n15130));
  jnot g14841(.din(n15130), .dout(n15131));
  jor  g14842(.dina(n15131), .dinb(n15123), .dout(n15132));
  jand g14843(.dina(n15132), .dinb(n15121), .dout(n15133));
  jor  g14844(.dina(n15133), .dinb(n2870), .dout(n15134));
  jxor g14845(.dina(n14548), .dinb(n2875), .dout(n15135));
  jor  g14846(.dina(n15135), .dinb(n14821), .dout(n15136));
  jxor g14847(.dina(n15136), .dinb(n14559), .dout(n15137));
  jand g14848(.dina(n15133), .dinb(n2870), .dout(n15138));
  jor  g14849(.dina(n15138), .dinb(n15137), .dout(n15139));
  jand g14850(.dina(n15139), .dinb(n15134), .dout(n15140));
  jor  g14851(.dina(n15140), .dinb(n2425), .dout(n15141));
  jnot g14852(.din(n14564), .dout(n15142));
  jor  g14853(.dina(n15142), .dinb(n14562), .dout(n15143));
  jor  g14854(.dina(n15143), .dinb(n14821), .dout(n15144));
  jxor g14855(.dina(n15144), .dinb(n14573), .dout(n15145));
  jand g14856(.dina(n15134), .dinb(n2425), .dout(n15146));
  jand g14857(.dina(n15146), .dinb(n15139), .dout(n15147));
  jor  g14858(.dina(n15147), .dinb(n15145), .dout(n15148));
  jand g14859(.dina(n15148), .dinb(n15141), .dout(n15149));
  jor  g14860(.dina(n15149), .dinb(n2420), .dout(n15150));
  jand g14861(.dina(n15149), .dinb(n2420), .dout(n15151));
  jnot g14862(.din(n14576), .dout(n15152));
  jand g14863(.dina(asqrt[11] ), .dinb(n15152), .dout(n15153));
  jand g14864(.dina(n15153), .dinb(n14581), .dout(n15154));
  jor  g14865(.dina(n15154), .dinb(n14580), .dout(n15155));
  jand g14866(.dina(n15153), .dinb(n14582), .dout(n15156));
  jnot g14867(.din(n15156), .dout(n15157));
  jand g14868(.dina(n15157), .dinb(n15155), .dout(n15158));
  jnot g14869(.din(n15158), .dout(n15159));
  jor  g14870(.dina(n15159), .dinb(n15151), .dout(n15160));
  jand g14871(.dina(n15160), .dinb(n15150), .dout(n15161));
  jor  g14872(.dina(n15161), .dinb(n2010), .dout(n15162));
  jand g14873(.dina(n15150), .dinb(n2010), .dout(n15163));
  jand g14874(.dina(n15163), .dinb(n15160), .dout(n15164));
  jnot g14875(.din(n14584), .dout(n15165));
  jand g14876(.dina(asqrt[11] ), .dinb(n15165), .dout(n15166));
  jand g14877(.dina(n15166), .dinb(n14591), .dout(n15167));
  jor  g14878(.dina(n15167), .dinb(n14589), .dout(n15168));
  jand g14879(.dina(n15166), .dinb(n14592), .dout(n15169));
  jnot g14880(.din(n15169), .dout(n15170));
  jand g14881(.dina(n15170), .dinb(n15168), .dout(n15171));
  jnot g14882(.din(n15171), .dout(n15172));
  jor  g14883(.dina(n15172), .dinb(n15164), .dout(n15173));
  jand g14884(.dina(n15173), .dinb(n15162), .dout(n15174));
  jor  g14885(.dina(n15174), .dinb(n2005), .dout(n15175));
  jxor g14886(.dina(n14593), .dinb(n2010), .dout(n15176));
  jor  g14887(.dina(n15176), .dinb(n14821), .dout(n15177));
  jxor g14888(.dina(n15177), .dinb(n14604), .dout(n15178));
  jand g14889(.dina(n15174), .dinb(n2005), .dout(n15179));
  jor  g14890(.dina(n15179), .dinb(n15178), .dout(n15180));
  jand g14891(.dina(n15180), .dinb(n15175), .dout(n15181));
  jor  g14892(.dina(n15181), .dinb(n1646), .dout(n15182));
  jnot g14893(.din(n14609), .dout(n15183));
  jor  g14894(.dina(n15183), .dinb(n14607), .dout(n15184));
  jor  g14895(.dina(n15184), .dinb(n14821), .dout(n15185));
  jxor g14896(.dina(n15185), .dinb(n14618), .dout(n15186));
  jand g14897(.dina(n15175), .dinb(n1646), .dout(n15187));
  jand g14898(.dina(n15187), .dinb(n15180), .dout(n15188));
  jor  g14899(.dina(n15188), .dinb(n15186), .dout(n15189));
  jand g14900(.dina(n15189), .dinb(n15182), .dout(n15190));
  jor  g14901(.dina(n15190), .dinb(n1641), .dout(n15191));
  jand g14902(.dina(n15190), .dinb(n1641), .dout(n15192));
  jnot g14903(.din(n14621), .dout(n15193));
  jand g14904(.dina(asqrt[11] ), .dinb(n15193), .dout(n15194));
  jand g14905(.dina(n15194), .dinb(n14626), .dout(n15195));
  jor  g14906(.dina(n15195), .dinb(n14625), .dout(n15196));
  jand g14907(.dina(n15194), .dinb(n14627), .dout(n15197));
  jnot g14908(.din(n15197), .dout(n15198));
  jand g14909(.dina(n15198), .dinb(n15196), .dout(n15199));
  jnot g14910(.din(n15199), .dout(n15200));
  jor  g14911(.dina(n15200), .dinb(n15192), .dout(n15201));
  jand g14912(.dina(n15201), .dinb(n15191), .dout(n15202));
  jor  g14913(.dina(n15202), .dinb(n1317), .dout(n15203));
  jand g14914(.dina(n15191), .dinb(n1317), .dout(n15204));
  jand g14915(.dina(n15204), .dinb(n15201), .dout(n15205));
  jnot g14916(.din(n14629), .dout(n15206));
  jand g14917(.dina(asqrt[11] ), .dinb(n15206), .dout(n15207));
  jand g14918(.dina(n15207), .dinb(n14636), .dout(n15208));
  jor  g14919(.dina(n15208), .dinb(n14634), .dout(n15209));
  jand g14920(.dina(n15207), .dinb(n14637), .dout(n15210));
  jnot g14921(.din(n15210), .dout(n15211));
  jand g14922(.dina(n15211), .dinb(n15209), .dout(n15212));
  jnot g14923(.din(n15212), .dout(n15213));
  jor  g14924(.dina(n15213), .dinb(n15205), .dout(n15214));
  jand g14925(.dina(n15214), .dinb(n15203), .dout(n15215));
  jor  g14926(.dina(n15215), .dinb(n1312), .dout(n15216));
  jxor g14927(.dina(n14638), .dinb(n1317), .dout(n15217));
  jor  g14928(.dina(n15217), .dinb(n14821), .dout(n15218));
  jxor g14929(.dina(n15218), .dinb(n14649), .dout(n15219));
  jand g14930(.dina(n15215), .dinb(n1312), .dout(n15220));
  jor  g14931(.dina(n15220), .dinb(n15219), .dout(n15221));
  jand g14932(.dina(n15221), .dinb(n15216), .dout(n15222));
  jor  g14933(.dina(n15222), .dinb(n1039), .dout(n15223));
  jand g14934(.dina(n15216), .dinb(n1039), .dout(n15224));
  jand g14935(.dina(n15224), .dinb(n15221), .dout(n15225));
  jnot g14936(.din(n14652), .dout(n15226));
  jand g14937(.dina(asqrt[11] ), .dinb(n15226), .dout(n15227));
  jand g14938(.dina(n15227), .dinb(n14659), .dout(n15228));
  jor  g14939(.dina(n15228), .dinb(n14657), .dout(n15229));
  jand g14940(.dina(n15227), .dinb(n14660), .dout(n15230));
  jnot g14941(.din(n15230), .dout(n15231));
  jand g14942(.dina(n15231), .dinb(n15229), .dout(n15232));
  jnot g14943(.din(n15232), .dout(n15233));
  jor  g14944(.dina(n15233), .dinb(n15225), .dout(n15234));
  jand g14945(.dina(n15234), .dinb(n15223), .dout(n15235));
  jor  g14946(.dina(n15235), .dinb(n1034), .dout(n15236));
  jnot g14947(.din(n14824), .dout(n15237));
  jand g14948(.dina(n15235), .dinb(n1034), .dout(n15238));
  jor  g14949(.dina(n15238), .dinb(n15237), .dout(n15239));
  jand g14950(.dina(n15239), .dinb(n15236), .dout(n15240));
  jor  g14951(.dina(n15240), .dinb(n796), .dout(n15241));
  jnot g14952(.din(n14669), .dout(n15242));
  jor  g14953(.dina(n15242), .dinb(n14667), .dout(n15243));
  jor  g14954(.dina(n15243), .dinb(n14821), .dout(n15244));
  jxor g14955(.dina(n15244), .dinb(n14678), .dout(n15245));
  jand g14956(.dina(n15236), .dinb(n796), .dout(n15246));
  jand g14957(.dina(n15246), .dinb(n15239), .dout(n15247));
  jor  g14958(.dina(n15247), .dinb(n15245), .dout(n15248));
  jand g14959(.dina(n15248), .dinb(n15241), .dout(n15249));
  jor  g14960(.dina(n15249), .dinb(n791), .dout(n15250));
  jxor g14961(.dina(n14680), .dinb(n796), .dout(n15251));
  jor  g14962(.dina(n15251), .dinb(n14821), .dout(n15252));
  jxor g14963(.dina(n15252), .dinb(n14691), .dout(n15253));
  jand g14964(.dina(n15249), .dinb(n791), .dout(n15254));
  jor  g14965(.dina(n15254), .dinb(n15253), .dout(n15255));
  jand g14966(.dina(n15255), .dinb(n15250), .dout(n15256));
  jor  g14967(.dina(n15256), .dinb(n595), .dout(n15257));
  jnot g14968(.din(n14696), .dout(n15258));
  jor  g14969(.dina(n15258), .dinb(n14694), .dout(n15259));
  jor  g14970(.dina(n15259), .dinb(n14821), .dout(n15260));
  jxor g14971(.dina(n15260), .dinb(n14705), .dout(n15261));
  jand g14972(.dina(n15250), .dinb(n595), .dout(n15262));
  jand g14973(.dina(n15262), .dinb(n15255), .dout(n15263));
  jor  g14974(.dina(n15263), .dinb(n15261), .dout(n15264));
  jand g14975(.dina(n15264), .dinb(n15257), .dout(n15265));
  jor  g14976(.dina(n15265), .dinb(n590), .dout(n15266));
  jand g14977(.dina(n15265), .dinb(n590), .dout(n15267));
  jnot g14978(.din(n14708), .dout(n15268));
  jand g14979(.dina(asqrt[11] ), .dinb(n15268), .dout(n15269));
  jand g14980(.dina(n15269), .dinb(n14713), .dout(n15270));
  jor  g14981(.dina(n15270), .dinb(n14712), .dout(n15271));
  jand g14982(.dina(n15269), .dinb(n14714), .dout(n15272));
  jnot g14983(.din(n15272), .dout(n15273));
  jand g14984(.dina(n15273), .dinb(n15271), .dout(n15274));
  jnot g14985(.din(n15274), .dout(n15275));
  jor  g14986(.dina(n15275), .dinb(n15267), .dout(n15276));
  jand g14987(.dina(n15276), .dinb(n15266), .dout(n15277));
  jor  g14988(.dina(n15277), .dinb(n430), .dout(n15278));
  jand g14989(.dina(n15266), .dinb(n430), .dout(n15279));
  jand g14990(.dina(n15279), .dinb(n15276), .dout(n15280));
  jnot g14991(.din(n14716), .dout(n15281));
  jand g14992(.dina(asqrt[11] ), .dinb(n15281), .dout(n15282));
  jand g14993(.dina(n15282), .dinb(n14723), .dout(n15283));
  jor  g14994(.dina(n15283), .dinb(n14721), .dout(n15284));
  jand g14995(.dina(n15282), .dinb(n14724), .dout(n15285));
  jnot g14996(.din(n15285), .dout(n15286));
  jand g14997(.dina(n15286), .dinb(n15284), .dout(n15287));
  jnot g14998(.din(n15287), .dout(n15288));
  jor  g14999(.dina(n15288), .dinb(n15280), .dout(n15289));
  jand g15000(.dina(n15289), .dinb(n15278), .dout(n15290));
  jor  g15001(.dina(n15290), .dinb(n425), .dout(n15291));
  jxor g15002(.dina(n14725), .dinb(n430), .dout(n15292));
  jor  g15003(.dina(n15292), .dinb(n14821), .dout(n15293));
  jxor g15004(.dina(n15293), .dinb(n14736), .dout(n15294));
  jand g15005(.dina(n15290), .dinb(n425), .dout(n15295));
  jor  g15006(.dina(n15295), .dinb(n15294), .dout(n15296));
  jand g15007(.dina(n15296), .dinb(n15291), .dout(n15297));
  jor  g15008(.dina(n15297), .dinb(n305), .dout(n15298));
  jnot g15009(.din(n14741), .dout(n15299));
  jor  g15010(.dina(n15299), .dinb(n14739), .dout(n15300));
  jor  g15011(.dina(n15300), .dinb(n14821), .dout(n15301));
  jxor g15012(.dina(n15301), .dinb(n14750), .dout(n15302));
  jand g15013(.dina(n15291), .dinb(n305), .dout(n15303));
  jand g15014(.dina(n15303), .dinb(n15296), .dout(n15304));
  jor  g15015(.dina(n15304), .dinb(n15302), .dout(n15305));
  jand g15016(.dina(n15305), .dinb(n15298), .dout(n15306));
  jor  g15017(.dina(n15306), .dinb(n290), .dout(n15307));
  jand g15018(.dina(n15306), .dinb(n290), .dout(n15308));
  jnot g15019(.din(n14753), .dout(n15309));
  jand g15020(.dina(asqrt[11] ), .dinb(n15309), .dout(n15310));
  jand g15021(.dina(n15310), .dinb(n14758), .dout(n15311));
  jor  g15022(.dina(n15311), .dinb(n14757), .dout(n15312));
  jand g15023(.dina(n15310), .dinb(n14759), .dout(n15313));
  jnot g15024(.din(n15313), .dout(n15314));
  jand g15025(.dina(n15314), .dinb(n15312), .dout(n15315));
  jnot g15026(.din(n15315), .dout(n15316));
  jor  g15027(.dina(n15316), .dinb(n15308), .dout(n15317));
  jand g15028(.dina(n15317), .dinb(n15307), .dout(n15318));
  jor  g15029(.dina(n15318), .dinb(n223), .dout(n15319));
  jand g15030(.dina(n15307), .dinb(n223), .dout(n15320));
  jand g15031(.dina(n15320), .dinb(n15317), .dout(n15321));
  jnot g15032(.din(n14761), .dout(n15322));
  jand g15033(.dina(asqrt[11] ), .dinb(n15322), .dout(n15323));
  jand g15034(.dina(n15323), .dinb(n14768), .dout(n15324));
  jor  g15035(.dina(n15324), .dinb(n14766), .dout(n15325));
  jand g15036(.dina(n15323), .dinb(n14769), .dout(n15326));
  jnot g15037(.din(n15326), .dout(n15327));
  jand g15038(.dina(n15327), .dinb(n15325), .dout(n15328));
  jnot g15039(.din(n15328), .dout(n15329));
  jor  g15040(.dina(n15329), .dinb(n15321), .dout(n15330));
  jand g15041(.dina(n15330), .dinb(n15319), .dout(n15331));
  jor  g15042(.dina(n15331), .dinb(n199), .dout(n15332));
  jand g15043(.dina(n15331), .dinb(n199), .dout(n15333));
  jxor g15044(.dina(n14770), .dinb(n223), .dout(n15334));
  jor  g15045(.dina(n15334), .dinb(n14821), .dout(n15335));
  jxor g15046(.dina(n15335), .dinb(n14781), .dout(n15336));
  jor  g15047(.dina(n15336), .dinb(n15333), .dout(n15337));
  jand g15048(.dina(n15337), .dinb(n15332), .dout(n15338));
  jnot g15049(.din(n14786), .dout(n15339));
  jor  g15050(.dina(n15339), .dinb(n14784), .dout(n15340));
  jor  g15051(.dina(n15340), .dinb(n14821), .dout(n15341));
  jxor g15052(.dina(n15341), .dinb(n14795), .dout(n15342));
  jand g15053(.dina(asqrt[11] ), .dinb(n14809), .dout(n15343));
  jand g15054(.dina(n15343), .dinb(n14797), .dout(n15344));
  jor  g15055(.dina(n15344), .dinb(n14843), .dout(n15345));
  jor  g15056(.dina(n15345), .dinb(n15342), .dout(n15346));
  jor  g15057(.dina(n15346), .dinb(n15338), .dout(n15347));
  jand g15058(.dina(n15347), .dinb(n194), .dout(n15348));
  jand g15059(.dina(n15342), .dinb(n15338), .dout(n15349));
  jor  g15060(.dina(n15343), .dinb(n14797), .dout(n15350));
  jand g15061(.dina(n14809), .dinb(n14797), .dout(n15351));
  jor  g15062(.dina(n15351), .dinb(n194), .dout(n15352));
  jnot g15063(.din(n15352), .dout(n15353));
  jand g15064(.dina(n15353), .dinb(n15350), .dout(n15354));
  jor  g15065(.dina(n15354), .dinb(n15349), .dout(n15357));
  jor  g15066(.dina(n15357), .dinb(n15348), .dout(asqrt[10] ));
  jxor g15067(.dina(n15235), .dinb(n1034), .dout(n15359));
  jand g15068(.dina(n15359), .dinb(asqrt[10] ), .dout(n15360));
  jxor g15069(.dina(n15360), .dinb(n14824), .dout(n15361));
  jnot g15070(.din(n15361), .dout(n15362));
  jand g15071(.dina(asqrt[10] ), .dinb(a[20] ), .dout(n15363));
  jnot g15072(.din(a[18] ), .dout(n15364));
  jnot g15073(.din(a[19] ), .dout(n15365));
  jand g15074(.dina(n14826), .dinb(n15365), .dout(n15366));
  jand g15075(.dina(n15366), .dinb(n15364), .dout(n15367));
  jor  g15076(.dina(n15367), .dinb(n15363), .dout(n15368));
  jand g15077(.dina(n15368), .dinb(asqrt[11] ), .dout(n15369));
  jand g15078(.dina(asqrt[10] ), .dinb(n14826), .dout(n15370));
  jxor g15079(.dina(n15370), .dinb(n14827), .dout(n15371));
  jor  g15080(.dina(n15368), .dinb(asqrt[11] ), .dout(n15372));
  jand g15081(.dina(n15372), .dinb(n15371), .dout(n15373));
  jor  g15082(.dina(n15373), .dinb(n15369), .dout(n15374));
  jand g15083(.dina(n15374), .dinb(asqrt[12] ), .dout(n15375));
  jor  g15084(.dina(n15369), .dinb(asqrt[12] ), .dout(n15376));
  jor  g15085(.dina(n15376), .dinb(n15373), .dout(n15377));
  jand g15086(.dina(n15370), .dinb(n14827), .dout(n15378));
  jnot g15087(.din(n15348), .dout(n15379));
  jnot g15088(.din(n15349), .dout(n15380));
  jnot g15089(.din(n15354), .dout(n15381));
  jand g15090(.dina(n15381), .dinb(asqrt[11] ), .dout(n15382));
  jand g15091(.dina(n15382), .dinb(n15380), .dout(n15383));
  jand g15092(.dina(n15383), .dinb(n15379), .dout(n15384));
  jor  g15093(.dina(n15384), .dinb(n15378), .dout(n15385));
  jxor g15094(.dina(n15385), .dinb(n14248), .dout(n15386));
  jand g15095(.dina(n15386), .dinb(n15377), .dout(n15387));
  jor  g15096(.dina(n15387), .dinb(n15375), .dout(n15388));
  jand g15097(.dina(n15388), .dinb(asqrt[13] ), .dout(n15389));
  jor  g15098(.dina(n15388), .dinb(asqrt[13] ), .dout(n15390));
  jxor g15099(.dina(n14831), .dinb(n14816), .dout(n15391));
  jand g15100(.dina(n15391), .dinb(asqrt[10] ), .dout(n15392));
  jxor g15101(.dina(n15392), .dinb(n14834), .dout(n15393));
  jnot g15102(.din(n15393), .dout(n15394));
  jand g15103(.dina(n15394), .dinb(n15390), .dout(n15395));
  jor  g15104(.dina(n15395), .dinb(n15389), .dout(n15396));
  jand g15105(.dina(n15396), .dinb(asqrt[14] ), .dout(n15397));
  jnot g15106(.din(n14840), .dout(n15398));
  jand g15107(.dina(n15398), .dinb(n14838), .dout(n15399));
  jand g15108(.dina(n15399), .dinb(asqrt[10] ), .dout(n15400));
  jxor g15109(.dina(n15400), .dinb(n14848), .dout(n15401));
  jnot g15110(.din(n15401), .dout(n15402));
  jor  g15111(.dina(n15389), .dinb(asqrt[14] ), .dout(n15403));
  jor  g15112(.dina(n15403), .dinb(n15395), .dout(n15404));
  jand g15113(.dina(n15404), .dinb(n15402), .dout(n15405));
  jor  g15114(.dina(n15405), .dinb(n15397), .dout(n15406));
  jand g15115(.dina(n15406), .dinb(asqrt[15] ), .dout(n15407));
  jor  g15116(.dina(n15406), .dinb(asqrt[15] ), .dout(n15408));
  jnot g15117(.din(n14855), .dout(n15409));
  jxor g15118(.dina(n14850), .dinb(n13718), .dout(n15410));
  jand g15119(.dina(n15410), .dinb(asqrt[10] ), .dout(n15411));
  jxor g15120(.dina(n15411), .dinb(n15409), .dout(n15412));
  jand g15121(.dina(n15412), .dinb(n15408), .dout(n15413));
  jor  g15122(.dina(n15413), .dinb(n15407), .dout(n15414));
  jand g15123(.dina(n15414), .dinb(asqrt[16] ), .dout(n15415));
  jor  g15124(.dina(n15407), .dinb(asqrt[16] ), .dout(n15416));
  jor  g15125(.dina(n15416), .dinb(n15413), .dout(n15417));
  jnot g15126(.din(n14862), .dout(n15418));
  jnot g15127(.din(n14864), .dout(n15419));
  jand g15128(.dina(asqrt[10] ), .dinb(n14858), .dout(n15420));
  jand g15129(.dina(n15420), .dinb(n15419), .dout(n15421));
  jor  g15130(.dina(n15421), .dinb(n15418), .dout(n15422));
  jnot g15131(.din(n14865), .dout(n15423));
  jand g15132(.dina(n15420), .dinb(n15423), .dout(n15424));
  jnot g15133(.din(n15424), .dout(n15425));
  jand g15134(.dina(n15425), .dinb(n15422), .dout(n15426));
  jand g15135(.dina(n15426), .dinb(n15417), .dout(n15427));
  jor  g15136(.dina(n15427), .dinb(n15415), .dout(n15428));
  jand g15137(.dina(n15428), .dinb(asqrt[17] ), .dout(n15429));
  jor  g15138(.dina(n15428), .dinb(asqrt[17] ), .dout(n15430));
  jxor g15139(.dina(n14866), .dinb(n12670), .dout(n15431));
  jand g15140(.dina(n15431), .dinb(asqrt[10] ), .dout(n15432));
  jxor g15141(.dina(n15432), .dinb(n14871), .dout(n15433));
  jand g15142(.dina(n15433), .dinb(n15430), .dout(n15434));
  jor  g15143(.dina(n15434), .dinb(n15429), .dout(n15435));
  jand g15144(.dina(n15435), .dinb(asqrt[18] ), .dout(n15436));
  jnot g15145(.din(n14877), .dout(n15437));
  jand g15146(.dina(n15437), .dinb(n14875), .dout(n15438));
  jand g15147(.dina(n15438), .dinb(asqrt[10] ), .dout(n15439));
  jxor g15148(.dina(n15439), .dinb(n14886), .dout(n15440));
  jnot g15149(.din(n15440), .dout(n15441));
  jor  g15150(.dina(n15429), .dinb(asqrt[18] ), .dout(n15442));
  jor  g15151(.dina(n15442), .dinb(n15434), .dout(n15443));
  jand g15152(.dina(n15443), .dinb(n15441), .dout(n15444));
  jor  g15153(.dina(n15444), .dinb(n15436), .dout(n15445));
  jand g15154(.dina(n15445), .dinb(asqrt[19] ), .dout(n15446));
  jor  g15155(.dina(n15445), .dinb(asqrt[19] ), .dout(n15447));
  jxor g15156(.dina(n14888), .dinb(n11657), .dout(n15448));
  jand g15157(.dina(n15448), .dinb(asqrt[10] ), .dout(n15449));
  jxor g15158(.dina(n15449), .dinb(n14894), .dout(n15450));
  jand g15159(.dina(n15450), .dinb(n15447), .dout(n15451));
  jor  g15160(.dina(n15451), .dinb(n15446), .dout(n15452));
  jand g15161(.dina(n15452), .dinb(asqrt[20] ), .dout(n15453));
  jor  g15162(.dina(n15446), .dinb(asqrt[20] ), .dout(n15454));
  jor  g15163(.dina(n15454), .dinb(n15451), .dout(n15455));
  jnot g15164(.din(n14902), .dout(n15456));
  jnot g15165(.din(n14904), .dout(n15457));
  jand g15166(.dina(asqrt[10] ), .dinb(n14898), .dout(n15458));
  jand g15167(.dina(n15458), .dinb(n15457), .dout(n15459));
  jor  g15168(.dina(n15459), .dinb(n15456), .dout(n15460));
  jnot g15169(.din(n14905), .dout(n15461));
  jand g15170(.dina(n15458), .dinb(n15461), .dout(n15462));
  jnot g15171(.din(n15462), .dout(n15463));
  jand g15172(.dina(n15463), .dinb(n15460), .dout(n15464));
  jand g15173(.dina(n15464), .dinb(n15455), .dout(n15465));
  jor  g15174(.dina(n15465), .dinb(n15453), .dout(n15466));
  jand g15175(.dina(n15466), .dinb(asqrt[21] ), .dout(n15467));
  jxor g15176(.dina(n14906), .dinb(n10696), .dout(n15468));
  jand g15177(.dina(n15468), .dinb(asqrt[10] ), .dout(n15469));
  jxor g15178(.dina(n15469), .dinb(n14913), .dout(n15470));
  jnot g15179(.din(n15470), .dout(n15471));
  jor  g15180(.dina(n15466), .dinb(asqrt[21] ), .dout(n15472));
  jand g15181(.dina(n15472), .dinb(n15471), .dout(n15473));
  jor  g15182(.dina(n15473), .dinb(n15467), .dout(n15474));
  jand g15183(.dina(n15474), .dinb(asqrt[22] ), .dout(n15475));
  jnot g15184(.din(n14918), .dout(n15476));
  jand g15185(.dina(n15476), .dinb(n14916), .dout(n15477));
  jand g15186(.dina(n15477), .dinb(asqrt[10] ), .dout(n15478));
  jxor g15187(.dina(n15478), .dinb(n14926), .dout(n15479));
  jnot g15188(.din(n15479), .dout(n15480));
  jor  g15189(.dina(n15467), .dinb(asqrt[22] ), .dout(n15481));
  jor  g15190(.dina(n15481), .dinb(n15473), .dout(n15482));
  jand g15191(.dina(n15482), .dinb(n15480), .dout(n15483));
  jor  g15192(.dina(n15483), .dinb(n15475), .dout(n15484));
  jand g15193(.dina(n15484), .dinb(asqrt[23] ), .dout(n15485));
  jor  g15194(.dina(n15484), .dinb(asqrt[23] ), .dout(n15486));
  jnot g15195(.din(n14932), .dout(n15487));
  jnot g15196(.din(n14933), .dout(n15488));
  jand g15197(.dina(asqrt[10] ), .dinb(n14929), .dout(n15489));
  jand g15198(.dina(n15489), .dinb(n15488), .dout(n15490));
  jor  g15199(.dina(n15490), .dinb(n15487), .dout(n15491));
  jnot g15200(.din(n14934), .dout(n15492));
  jand g15201(.dina(n15489), .dinb(n15492), .dout(n15493));
  jnot g15202(.din(n15493), .dout(n15494));
  jand g15203(.dina(n15494), .dinb(n15491), .dout(n15495));
  jand g15204(.dina(n15495), .dinb(n15486), .dout(n15496));
  jor  g15205(.dina(n15496), .dinb(n15485), .dout(n15497));
  jand g15206(.dina(n15497), .dinb(asqrt[24] ), .dout(n15498));
  jor  g15207(.dina(n15485), .dinb(asqrt[24] ), .dout(n15499));
  jor  g15208(.dina(n15499), .dinb(n15496), .dout(n15500));
  jnot g15209(.din(n14940), .dout(n15501));
  jnot g15210(.din(n14942), .dout(n15502));
  jand g15211(.dina(asqrt[10] ), .dinb(n14936), .dout(n15503));
  jand g15212(.dina(n15503), .dinb(n15502), .dout(n15504));
  jor  g15213(.dina(n15504), .dinb(n15501), .dout(n15505));
  jnot g15214(.din(n14943), .dout(n15506));
  jand g15215(.dina(n15503), .dinb(n15506), .dout(n15507));
  jnot g15216(.din(n15507), .dout(n15508));
  jand g15217(.dina(n15508), .dinb(n15505), .dout(n15509));
  jand g15218(.dina(n15509), .dinb(n15500), .dout(n15510));
  jor  g15219(.dina(n15510), .dinb(n15498), .dout(n15511));
  jand g15220(.dina(n15511), .dinb(asqrt[25] ), .dout(n15512));
  jxor g15221(.dina(n14944), .dinb(n8893), .dout(n15513));
  jand g15222(.dina(n15513), .dinb(asqrt[10] ), .dout(n15514));
  jxor g15223(.dina(n15514), .dinb(n14954), .dout(n15515));
  jnot g15224(.din(n15515), .dout(n15516));
  jor  g15225(.dina(n15511), .dinb(asqrt[25] ), .dout(n15517));
  jand g15226(.dina(n15517), .dinb(n15516), .dout(n15518));
  jor  g15227(.dina(n15518), .dinb(n15512), .dout(n15519));
  jand g15228(.dina(n15519), .dinb(asqrt[26] ), .dout(n15520));
  jnot g15229(.din(n14959), .dout(n15521));
  jand g15230(.dina(n15521), .dinb(n14957), .dout(n15522));
  jand g15231(.dina(n15522), .dinb(asqrt[10] ), .dout(n15523));
  jxor g15232(.dina(n15523), .dinb(n14967), .dout(n15524));
  jnot g15233(.din(n15524), .dout(n15525));
  jor  g15234(.dina(n15512), .dinb(asqrt[26] ), .dout(n15526));
  jor  g15235(.dina(n15526), .dinb(n15518), .dout(n15527));
  jand g15236(.dina(n15527), .dinb(n15525), .dout(n15528));
  jor  g15237(.dina(n15528), .dinb(n15520), .dout(n15529));
  jand g15238(.dina(n15529), .dinb(asqrt[27] ), .dout(n15530));
  jor  g15239(.dina(n15529), .dinb(asqrt[27] ), .dout(n15531));
  jnot g15240(.din(n14973), .dout(n15532));
  jnot g15241(.din(n14974), .dout(n15533));
  jand g15242(.dina(asqrt[10] ), .dinb(n14970), .dout(n15534));
  jand g15243(.dina(n15534), .dinb(n15533), .dout(n15535));
  jor  g15244(.dina(n15535), .dinb(n15532), .dout(n15536));
  jnot g15245(.din(n14975), .dout(n15537));
  jand g15246(.dina(n15534), .dinb(n15537), .dout(n15538));
  jnot g15247(.din(n15538), .dout(n15539));
  jand g15248(.dina(n15539), .dinb(n15536), .dout(n15540));
  jand g15249(.dina(n15540), .dinb(n15531), .dout(n15541));
  jor  g15250(.dina(n15541), .dinb(n15530), .dout(n15542));
  jand g15251(.dina(n15542), .dinb(asqrt[28] ), .dout(n15543));
  jor  g15252(.dina(n15530), .dinb(asqrt[28] ), .dout(n15544));
  jor  g15253(.dina(n15544), .dinb(n15541), .dout(n15545));
  jnot g15254(.din(n14981), .dout(n15546));
  jnot g15255(.din(n14983), .dout(n15547));
  jand g15256(.dina(asqrt[10] ), .dinb(n14977), .dout(n15548));
  jand g15257(.dina(n15548), .dinb(n15547), .dout(n15549));
  jor  g15258(.dina(n15549), .dinb(n15546), .dout(n15550));
  jnot g15259(.din(n14984), .dout(n15551));
  jand g15260(.dina(n15548), .dinb(n15551), .dout(n15552));
  jnot g15261(.din(n15552), .dout(n15553));
  jand g15262(.dina(n15553), .dinb(n15550), .dout(n15554));
  jand g15263(.dina(n15554), .dinb(n15545), .dout(n15555));
  jor  g15264(.dina(n15555), .dinb(n15543), .dout(n15556));
  jand g15265(.dina(n15556), .dinb(asqrt[29] ), .dout(n15557));
  jxor g15266(.dina(n14985), .dinb(n7260), .dout(n15558));
  jand g15267(.dina(n15558), .dinb(asqrt[10] ), .dout(n15559));
  jxor g15268(.dina(n15559), .dinb(n14995), .dout(n15560));
  jnot g15269(.din(n15560), .dout(n15561));
  jor  g15270(.dina(n15556), .dinb(asqrt[29] ), .dout(n15562));
  jand g15271(.dina(n15562), .dinb(n15561), .dout(n15563));
  jor  g15272(.dina(n15563), .dinb(n15557), .dout(n15564));
  jand g15273(.dina(n15564), .dinb(asqrt[30] ), .dout(n15565));
  jnot g15274(.din(n15000), .dout(n15566));
  jand g15275(.dina(n15566), .dinb(n14998), .dout(n15567));
  jand g15276(.dina(n15567), .dinb(asqrt[10] ), .dout(n15568));
  jxor g15277(.dina(n15568), .dinb(n15008), .dout(n15569));
  jnot g15278(.din(n15569), .dout(n15570));
  jor  g15279(.dina(n15557), .dinb(asqrt[30] ), .dout(n15571));
  jor  g15280(.dina(n15571), .dinb(n15563), .dout(n15572));
  jand g15281(.dina(n15572), .dinb(n15570), .dout(n15573));
  jor  g15282(.dina(n15573), .dinb(n15565), .dout(n15574));
  jand g15283(.dina(n15574), .dinb(asqrt[31] ), .dout(n15575));
  jor  g15284(.dina(n15574), .dinb(asqrt[31] ), .dout(n15576));
  jnot g15285(.din(n15014), .dout(n15577));
  jnot g15286(.din(n15015), .dout(n15578));
  jand g15287(.dina(asqrt[10] ), .dinb(n15011), .dout(n15579));
  jand g15288(.dina(n15579), .dinb(n15578), .dout(n15580));
  jor  g15289(.dina(n15580), .dinb(n15577), .dout(n15581));
  jnot g15290(.din(n15016), .dout(n15582));
  jand g15291(.dina(n15579), .dinb(n15582), .dout(n15583));
  jnot g15292(.din(n15583), .dout(n15584));
  jand g15293(.dina(n15584), .dinb(n15581), .dout(n15585));
  jand g15294(.dina(n15585), .dinb(n15576), .dout(n15586));
  jor  g15295(.dina(n15586), .dinb(n15575), .dout(n15587));
  jand g15296(.dina(n15587), .dinb(asqrt[32] ), .dout(n15588));
  jor  g15297(.dina(n15575), .dinb(asqrt[32] ), .dout(n15589));
  jor  g15298(.dina(n15589), .dinb(n15586), .dout(n15590));
  jnot g15299(.din(n15022), .dout(n15591));
  jnot g15300(.din(n15024), .dout(n15592));
  jand g15301(.dina(asqrt[10] ), .dinb(n15018), .dout(n15593));
  jand g15302(.dina(n15593), .dinb(n15592), .dout(n15594));
  jor  g15303(.dina(n15594), .dinb(n15591), .dout(n15595));
  jnot g15304(.din(n15025), .dout(n15596));
  jand g15305(.dina(n15593), .dinb(n15596), .dout(n15597));
  jnot g15306(.din(n15597), .dout(n15598));
  jand g15307(.dina(n15598), .dinb(n15595), .dout(n15599));
  jand g15308(.dina(n15599), .dinb(n15590), .dout(n15600));
  jor  g15309(.dina(n15600), .dinb(n15588), .dout(n15601));
  jand g15310(.dina(n15601), .dinb(asqrt[33] ), .dout(n15602));
  jxor g15311(.dina(n15026), .dinb(n5788), .dout(n15603));
  jand g15312(.dina(n15603), .dinb(asqrt[10] ), .dout(n15604));
  jxor g15313(.dina(n15604), .dinb(n15036), .dout(n15605));
  jnot g15314(.din(n15605), .dout(n15606));
  jor  g15315(.dina(n15601), .dinb(asqrt[33] ), .dout(n15607));
  jand g15316(.dina(n15607), .dinb(n15606), .dout(n15608));
  jor  g15317(.dina(n15608), .dinb(n15602), .dout(n15609));
  jand g15318(.dina(n15609), .dinb(asqrt[34] ), .dout(n15610));
  jnot g15319(.din(n15041), .dout(n15611));
  jand g15320(.dina(n15611), .dinb(n15039), .dout(n15612));
  jand g15321(.dina(n15612), .dinb(asqrt[10] ), .dout(n15613));
  jxor g15322(.dina(n15613), .dinb(n15049), .dout(n15614));
  jnot g15323(.din(n15614), .dout(n15615));
  jor  g15324(.dina(n15602), .dinb(asqrt[34] ), .dout(n15616));
  jor  g15325(.dina(n15616), .dinb(n15608), .dout(n15617));
  jand g15326(.dina(n15617), .dinb(n15615), .dout(n15618));
  jor  g15327(.dina(n15618), .dinb(n15610), .dout(n15619));
  jand g15328(.dina(n15619), .dinb(asqrt[35] ), .dout(n15620));
  jor  g15329(.dina(n15619), .dinb(asqrt[35] ), .dout(n15621));
  jnot g15330(.din(n15055), .dout(n15622));
  jnot g15331(.din(n15056), .dout(n15623));
  jand g15332(.dina(asqrt[10] ), .dinb(n15052), .dout(n15624));
  jand g15333(.dina(n15624), .dinb(n15623), .dout(n15625));
  jor  g15334(.dina(n15625), .dinb(n15622), .dout(n15626));
  jnot g15335(.din(n15057), .dout(n15627));
  jand g15336(.dina(n15624), .dinb(n15627), .dout(n15628));
  jnot g15337(.din(n15628), .dout(n15629));
  jand g15338(.dina(n15629), .dinb(n15626), .dout(n15630));
  jand g15339(.dina(n15630), .dinb(n15621), .dout(n15631));
  jor  g15340(.dina(n15631), .dinb(n15620), .dout(n15632));
  jand g15341(.dina(n15632), .dinb(asqrt[36] ), .dout(n15633));
  jor  g15342(.dina(n15620), .dinb(asqrt[36] ), .dout(n15634));
  jor  g15343(.dina(n15634), .dinb(n15631), .dout(n15635));
  jnot g15344(.din(n15063), .dout(n15636));
  jnot g15345(.din(n15065), .dout(n15637));
  jand g15346(.dina(asqrt[10] ), .dinb(n15059), .dout(n15638));
  jand g15347(.dina(n15638), .dinb(n15637), .dout(n15639));
  jor  g15348(.dina(n15639), .dinb(n15636), .dout(n15640));
  jnot g15349(.din(n15066), .dout(n15641));
  jand g15350(.dina(n15638), .dinb(n15641), .dout(n15642));
  jnot g15351(.din(n15642), .dout(n15643));
  jand g15352(.dina(n15643), .dinb(n15640), .dout(n15644));
  jand g15353(.dina(n15644), .dinb(n15635), .dout(n15645));
  jor  g15354(.dina(n15645), .dinb(n15633), .dout(n15646));
  jand g15355(.dina(n15646), .dinb(asqrt[37] ), .dout(n15647));
  jxor g15356(.dina(n15067), .dinb(n4494), .dout(n15648));
  jand g15357(.dina(n15648), .dinb(asqrt[10] ), .dout(n15649));
  jxor g15358(.dina(n15649), .dinb(n15077), .dout(n15650));
  jnot g15359(.din(n15650), .dout(n15651));
  jor  g15360(.dina(n15646), .dinb(asqrt[37] ), .dout(n15652));
  jand g15361(.dina(n15652), .dinb(n15651), .dout(n15653));
  jor  g15362(.dina(n15653), .dinb(n15647), .dout(n15654));
  jand g15363(.dina(n15654), .dinb(asqrt[38] ), .dout(n15655));
  jnot g15364(.din(n15082), .dout(n15656));
  jand g15365(.dina(n15656), .dinb(n15080), .dout(n15657));
  jand g15366(.dina(n15657), .dinb(asqrt[10] ), .dout(n15658));
  jxor g15367(.dina(n15658), .dinb(n15090), .dout(n15659));
  jnot g15368(.din(n15659), .dout(n15660));
  jor  g15369(.dina(n15647), .dinb(asqrt[38] ), .dout(n15661));
  jor  g15370(.dina(n15661), .dinb(n15653), .dout(n15662));
  jand g15371(.dina(n15662), .dinb(n15660), .dout(n15663));
  jor  g15372(.dina(n15663), .dinb(n15655), .dout(n15664));
  jand g15373(.dina(n15664), .dinb(asqrt[39] ), .dout(n15665));
  jor  g15374(.dina(n15664), .dinb(asqrt[39] ), .dout(n15666));
  jnot g15375(.din(n15096), .dout(n15667));
  jnot g15376(.din(n15097), .dout(n15668));
  jand g15377(.dina(asqrt[10] ), .dinb(n15093), .dout(n15669));
  jand g15378(.dina(n15669), .dinb(n15668), .dout(n15670));
  jor  g15379(.dina(n15670), .dinb(n15667), .dout(n15671));
  jnot g15380(.din(n15098), .dout(n15672));
  jand g15381(.dina(n15669), .dinb(n15672), .dout(n15673));
  jnot g15382(.din(n15673), .dout(n15674));
  jand g15383(.dina(n15674), .dinb(n15671), .dout(n15675));
  jand g15384(.dina(n15675), .dinb(n15666), .dout(n15676));
  jor  g15385(.dina(n15676), .dinb(n15665), .dout(n15677));
  jand g15386(.dina(n15677), .dinb(asqrt[40] ), .dout(n15678));
  jor  g15387(.dina(n15665), .dinb(asqrt[40] ), .dout(n15679));
  jor  g15388(.dina(n15679), .dinb(n15676), .dout(n15680));
  jnot g15389(.din(n15104), .dout(n15681));
  jnot g15390(.din(n15106), .dout(n15682));
  jand g15391(.dina(asqrt[10] ), .dinb(n15100), .dout(n15683));
  jand g15392(.dina(n15683), .dinb(n15682), .dout(n15684));
  jor  g15393(.dina(n15684), .dinb(n15681), .dout(n15685));
  jnot g15394(.din(n15107), .dout(n15686));
  jand g15395(.dina(n15683), .dinb(n15686), .dout(n15687));
  jnot g15396(.din(n15687), .dout(n15688));
  jand g15397(.dina(n15688), .dinb(n15685), .dout(n15689));
  jand g15398(.dina(n15689), .dinb(n15680), .dout(n15690));
  jor  g15399(.dina(n15690), .dinb(n15678), .dout(n15691));
  jand g15400(.dina(n15691), .dinb(asqrt[41] ), .dout(n15692));
  jxor g15401(.dina(n15108), .dinb(n3371), .dout(n15693));
  jand g15402(.dina(n15693), .dinb(asqrt[10] ), .dout(n15694));
  jxor g15403(.dina(n15694), .dinb(n15118), .dout(n15695));
  jnot g15404(.din(n15695), .dout(n15696));
  jor  g15405(.dina(n15691), .dinb(asqrt[41] ), .dout(n15697));
  jand g15406(.dina(n15697), .dinb(n15696), .dout(n15698));
  jor  g15407(.dina(n15698), .dinb(n15692), .dout(n15699));
  jand g15408(.dina(n15699), .dinb(asqrt[42] ), .dout(n15700));
  jnot g15409(.din(n15123), .dout(n15701));
  jand g15410(.dina(n15701), .dinb(n15121), .dout(n15702));
  jand g15411(.dina(n15702), .dinb(asqrt[10] ), .dout(n15703));
  jxor g15412(.dina(n15703), .dinb(n15131), .dout(n15704));
  jnot g15413(.din(n15704), .dout(n15705));
  jor  g15414(.dina(n15692), .dinb(asqrt[42] ), .dout(n15706));
  jor  g15415(.dina(n15706), .dinb(n15698), .dout(n15707));
  jand g15416(.dina(n15707), .dinb(n15705), .dout(n15708));
  jor  g15417(.dina(n15708), .dinb(n15700), .dout(n15709));
  jand g15418(.dina(n15709), .dinb(asqrt[43] ), .dout(n15710));
  jor  g15419(.dina(n15709), .dinb(asqrt[43] ), .dout(n15711));
  jnot g15420(.din(n15137), .dout(n15712));
  jnot g15421(.din(n15138), .dout(n15713));
  jand g15422(.dina(asqrt[10] ), .dinb(n15134), .dout(n15714));
  jand g15423(.dina(n15714), .dinb(n15713), .dout(n15715));
  jor  g15424(.dina(n15715), .dinb(n15712), .dout(n15716));
  jnot g15425(.din(n15139), .dout(n15717));
  jand g15426(.dina(n15714), .dinb(n15717), .dout(n15718));
  jnot g15427(.din(n15718), .dout(n15719));
  jand g15428(.dina(n15719), .dinb(n15716), .dout(n15720));
  jand g15429(.dina(n15720), .dinb(n15711), .dout(n15721));
  jor  g15430(.dina(n15721), .dinb(n15710), .dout(n15722));
  jand g15431(.dina(n15722), .dinb(asqrt[44] ), .dout(n15723));
  jor  g15432(.dina(n15710), .dinb(asqrt[44] ), .dout(n15724));
  jor  g15433(.dina(n15724), .dinb(n15721), .dout(n15725));
  jnot g15434(.din(n15145), .dout(n15726));
  jnot g15435(.din(n15147), .dout(n15727));
  jand g15436(.dina(asqrt[10] ), .dinb(n15141), .dout(n15728));
  jand g15437(.dina(n15728), .dinb(n15727), .dout(n15729));
  jor  g15438(.dina(n15729), .dinb(n15726), .dout(n15730));
  jnot g15439(.din(n15148), .dout(n15731));
  jand g15440(.dina(n15728), .dinb(n15731), .dout(n15732));
  jnot g15441(.din(n15732), .dout(n15733));
  jand g15442(.dina(n15733), .dinb(n15730), .dout(n15734));
  jand g15443(.dina(n15734), .dinb(n15725), .dout(n15735));
  jor  g15444(.dina(n15735), .dinb(n15723), .dout(n15736));
  jand g15445(.dina(n15736), .dinb(asqrt[45] ), .dout(n15737));
  jxor g15446(.dina(n15149), .dinb(n2420), .dout(n15738));
  jand g15447(.dina(n15738), .dinb(asqrt[10] ), .dout(n15739));
  jxor g15448(.dina(n15739), .dinb(n15159), .dout(n15740));
  jnot g15449(.din(n15740), .dout(n15741));
  jor  g15450(.dina(n15736), .dinb(asqrt[45] ), .dout(n15742));
  jand g15451(.dina(n15742), .dinb(n15741), .dout(n15743));
  jor  g15452(.dina(n15743), .dinb(n15737), .dout(n15744));
  jand g15453(.dina(n15744), .dinb(asqrt[46] ), .dout(n15745));
  jnot g15454(.din(n15164), .dout(n15746));
  jand g15455(.dina(n15746), .dinb(n15162), .dout(n15747));
  jand g15456(.dina(n15747), .dinb(asqrt[10] ), .dout(n15748));
  jxor g15457(.dina(n15748), .dinb(n15172), .dout(n15749));
  jnot g15458(.din(n15749), .dout(n15750));
  jor  g15459(.dina(n15737), .dinb(asqrt[46] ), .dout(n15751));
  jor  g15460(.dina(n15751), .dinb(n15743), .dout(n15752));
  jand g15461(.dina(n15752), .dinb(n15750), .dout(n15753));
  jor  g15462(.dina(n15753), .dinb(n15745), .dout(n15754));
  jand g15463(.dina(n15754), .dinb(asqrt[47] ), .dout(n15755));
  jor  g15464(.dina(n15754), .dinb(asqrt[47] ), .dout(n15756));
  jnot g15465(.din(n15178), .dout(n15757));
  jnot g15466(.din(n15179), .dout(n15758));
  jand g15467(.dina(asqrt[10] ), .dinb(n15175), .dout(n15759));
  jand g15468(.dina(n15759), .dinb(n15758), .dout(n15760));
  jor  g15469(.dina(n15760), .dinb(n15757), .dout(n15761));
  jnot g15470(.din(n15180), .dout(n15762));
  jand g15471(.dina(n15759), .dinb(n15762), .dout(n15763));
  jnot g15472(.din(n15763), .dout(n15764));
  jand g15473(.dina(n15764), .dinb(n15761), .dout(n15765));
  jand g15474(.dina(n15765), .dinb(n15756), .dout(n15766));
  jor  g15475(.dina(n15766), .dinb(n15755), .dout(n15767));
  jand g15476(.dina(n15767), .dinb(asqrt[48] ), .dout(n15768));
  jor  g15477(.dina(n15755), .dinb(asqrt[48] ), .dout(n15769));
  jor  g15478(.dina(n15769), .dinb(n15766), .dout(n15770));
  jnot g15479(.din(n15186), .dout(n15771));
  jnot g15480(.din(n15188), .dout(n15772));
  jand g15481(.dina(asqrt[10] ), .dinb(n15182), .dout(n15773));
  jand g15482(.dina(n15773), .dinb(n15772), .dout(n15774));
  jor  g15483(.dina(n15774), .dinb(n15771), .dout(n15775));
  jnot g15484(.din(n15189), .dout(n15776));
  jand g15485(.dina(n15773), .dinb(n15776), .dout(n15777));
  jnot g15486(.din(n15777), .dout(n15778));
  jand g15487(.dina(n15778), .dinb(n15775), .dout(n15779));
  jand g15488(.dina(n15779), .dinb(n15770), .dout(n15780));
  jor  g15489(.dina(n15780), .dinb(n15768), .dout(n15781));
  jand g15490(.dina(n15781), .dinb(asqrt[49] ), .dout(n15782));
  jxor g15491(.dina(n15190), .dinb(n1641), .dout(n15783));
  jand g15492(.dina(n15783), .dinb(asqrt[10] ), .dout(n15784));
  jxor g15493(.dina(n15784), .dinb(n15200), .dout(n15785));
  jnot g15494(.din(n15785), .dout(n15786));
  jor  g15495(.dina(n15781), .dinb(asqrt[49] ), .dout(n15787));
  jand g15496(.dina(n15787), .dinb(n15786), .dout(n15788));
  jor  g15497(.dina(n15788), .dinb(n15782), .dout(n15789));
  jand g15498(.dina(n15789), .dinb(asqrt[50] ), .dout(n15790));
  jnot g15499(.din(n15205), .dout(n15791));
  jand g15500(.dina(n15791), .dinb(n15203), .dout(n15792));
  jand g15501(.dina(n15792), .dinb(asqrt[10] ), .dout(n15793));
  jxor g15502(.dina(n15793), .dinb(n15213), .dout(n15794));
  jnot g15503(.din(n15794), .dout(n15795));
  jor  g15504(.dina(n15782), .dinb(asqrt[50] ), .dout(n15796));
  jor  g15505(.dina(n15796), .dinb(n15788), .dout(n15797));
  jand g15506(.dina(n15797), .dinb(n15795), .dout(n15798));
  jor  g15507(.dina(n15798), .dinb(n15790), .dout(n15799));
  jand g15508(.dina(n15799), .dinb(asqrt[51] ), .dout(n15800));
  jor  g15509(.dina(n15799), .dinb(asqrt[51] ), .dout(n15801));
  jnot g15510(.din(n15219), .dout(n15802));
  jnot g15511(.din(n15220), .dout(n15803));
  jand g15512(.dina(asqrt[10] ), .dinb(n15216), .dout(n15804));
  jand g15513(.dina(n15804), .dinb(n15803), .dout(n15805));
  jor  g15514(.dina(n15805), .dinb(n15802), .dout(n15806));
  jnot g15515(.din(n15221), .dout(n15807));
  jand g15516(.dina(n15804), .dinb(n15807), .dout(n15808));
  jnot g15517(.din(n15808), .dout(n15809));
  jand g15518(.dina(n15809), .dinb(n15806), .dout(n15810));
  jand g15519(.dina(n15810), .dinb(n15801), .dout(n15811));
  jor  g15520(.dina(n15811), .dinb(n15800), .dout(n15812));
  jand g15521(.dina(n15812), .dinb(asqrt[52] ), .dout(n15813));
  jnot g15522(.din(n15225), .dout(n15814));
  jand g15523(.dina(n15814), .dinb(n15223), .dout(n15815));
  jand g15524(.dina(n15815), .dinb(asqrt[10] ), .dout(n15816));
  jxor g15525(.dina(n15816), .dinb(n15233), .dout(n15817));
  jnot g15526(.din(n15817), .dout(n15818));
  jor  g15527(.dina(n15800), .dinb(asqrt[52] ), .dout(n15819));
  jor  g15528(.dina(n15819), .dinb(n15811), .dout(n15820));
  jand g15529(.dina(n15820), .dinb(n15818), .dout(n15821));
  jor  g15530(.dina(n15821), .dinb(n15813), .dout(n15822));
  jand g15531(.dina(n15822), .dinb(asqrt[53] ), .dout(n15823));
  jor  g15532(.dina(n15822), .dinb(asqrt[53] ), .dout(n15824));
  jand g15533(.dina(n15824), .dinb(n15361), .dout(n15825));
  jor  g15534(.dina(n15825), .dinb(n15823), .dout(n15826));
  jand g15535(.dina(n15826), .dinb(asqrt[54] ), .dout(n15827));
  jor  g15536(.dina(n15823), .dinb(asqrt[54] ), .dout(n15828));
  jor  g15537(.dina(n15828), .dinb(n15825), .dout(n15829));
  jnot g15538(.din(n15245), .dout(n15830));
  jnot g15539(.din(n15247), .dout(n15831));
  jand g15540(.dina(asqrt[10] ), .dinb(n15241), .dout(n15832));
  jand g15541(.dina(n15832), .dinb(n15831), .dout(n15833));
  jor  g15542(.dina(n15833), .dinb(n15830), .dout(n15834));
  jnot g15543(.din(n15248), .dout(n15835));
  jand g15544(.dina(n15832), .dinb(n15835), .dout(n15836));
  jnot g15545(.din(n15836), .dout(n15837));
  jand g15546(.dina(n15837), .dinb(n15834), .dout(n15838));
  jand g15547(.dina(n15838), .dinb(n15829), .dout(n15839));
  jor  g15548(.dina(n15839), .dinb(n15827), .dout(n15840));
  jand g15549(.dina(n15840), .dinb(asqrt[55] ), .dout(n15841));
  jor  g15550(.dina(n15840), .dinb(asqrt[55] ), .dout(n15842));
  jnot g15551(.din(n15253), .dout(n15843));
  jnot g15552(.din(n15254), .dout(n15844));
  jand g15553(.dina(asqrt[10] ), .dinb(n15250), .dout(n15845));
  jand g15554(.dina(n15845), .dinb(n15844), .dout(n15846));
  jor  g15555(.dina(n15846), .dinb(n15843), .dout(n15847));
  jnot g15556(.din(n15255), .dout(n15848));
  jand g15557(.dina(n15845), .dinb(n15848), .dout(n15849));
  jnot g15558(.din(n15849), .dout(n15850));
  jand g15559(.dina(n15850), .dinb(n15847), .dout(n15851));
  jand g15560(.dina(n15851), .dinb(n15842), .dout(n15852));
  jor  g15561(.dina(n15852), .dinb(n15841), .dout(n15853));
  jand g15562(.dina(n15853), .dinb(asqrt[56] ), .dout(n15854));
  jor  g15563(.dina(n15841), .dinb(asqrt[56] ), .dout(n15855));
  jor  g15564(.dina(n15855), .dinb(n15852), .dout(n15856));
  jnot g15565(.din(n15261), .dout(n15857));
  jnot g15566(.din(n15263), .dout(n15858));
  jand g15567(.dina(asqrt[10] ), .dinb(n15257), .dout(n15859));
  jand g15568(.dina(n15859), .dinb(n15858), .dout(n15860));
  jor  g15569(.dina(n15860), .dinb(n15857), .dout(n15861));
  jnot g15570(.din(n15264), .dout(n15862));
  jand g15571(.dina(n15859), .dinb(n15862), .dout(n15863));
  jnot g15572(.din(n15863), .dout(n15864));
  jand g15573(.dina(n15864), .dinb(n15861), .dout(n15865));
  jand g15574(.dina(n15865), .dinb(n15856), .dout(n15866));
  jor  g15575(.dina(n15866), .dinb(n15854), .dout(n15867));
  jand g15576(.dina(n15867), .dinb(asqrt[57] ), .dout(n15868));
  jxor g15577(.dina(n15265), .dinb(n590), .dout(n15869));
  jand g15578(.dina(n15869), .dinb(asqrt[10] ), .dout(n15870));
  jxor g15579(.dina(n15870), .dinb(n15275), .dout(n15871));
  jnot g15580(.din(n15871), .dout(n15872));
  jor  g15581(.dina(n15867), .dinb(asqrt[57] ), .dout(n15873));
  jand g15582(.dina(n15873), .dinb(n15872), .dout(n15874));
  jor  g15583(.dina(n15874), .dinb(n15868), .dout(n15875));
  jand g15584(.dina(n15875), .dinb(asqrt[58] ), .dout(n15876));
  jnot g15585(.din(n15280), .dout(n15877));
  jand g15586(.dina(n15877), .dinb(n15278), .dout(n15878));
  jand g15587(.dina(n15878), .dinb(asqrt[10] ), .dout(n15879));
  jxor g15588(.dina(n15879), .dinb(n15288), .dout(n15880));
  jnot g15589(.din(n15880), .dout(n15881));
  jor  g15590(.dina(n15868), .dinb(asqrt[58] ), .dout(n15882));
  jor  g15591(.dina(n15882), .dinb(n15874), .dout(n15883));
  jand g15592(.dina(n15883), .dinb(n15881), .dout(n15884));
  jor  g15593(.dina(n15884), .dinb(n15876), .dout(n15885));
  jand g15594(.dina(n15885), .dinb(asqrt[59] ), .dout(n15886));
  jor  g15595(.dina(n15885), .dinb(asqrt[59] ), .dout(n15887));
  jnot g15596(.din(n15294), .dout(n15888));
  jnot g15597(.din(n15295), .dout(n15889));
  jand g15598(.dina(asqrt[10] ), .dinb(n15291), .dout(n15890));
  jand g15599(.dina(n15890), .dinb(n15889), .dout(n15891));
  jor  g15600(.dina(n15891), .dinb(n15888), .dout(n15892));
  jnot g15601(.din(n15296), .dout(n15893));
  jand g15602(.dina(n15890), .dinb(n15893), .dout(n15894));
  jnot g15603(.din(n15894), .dout(n15895));
  jand g15604(.dina(n15895), .dinb(n15892), .dout(n15896));
  jand g15605(.dina(n15896), .dinb(n15887), .dout(n15897));
  jor  g15606(.dina(n15897), .dinb(n15886), .dout(n15898));
  jand g15607(.dina(n15898), .dinb(asqrt[60] ), .dout(n15899));
  jor  g15608(.dina(n15886), .dinb(asqrt[60] ), .dout(n15900));
  jor  g15609(.dina(n15900), .dinb(n15897), .dout(n15901));
  jnot g15610(.din(n15302), .dout(n15902));
  jnot g15611(.din(n15304), .dout(n15903));
  jand g15612(.dina(asqrt[10] ), .dinb(n15298), .dout(n15904));
  jand g15613(.dina(n15904), .dinb(n15903), .dout(n15905));
  jor  g15614(.dina(n15905), .dinb(n15902), .dout(n15906));
  jnot g15615(.din(n15305), .dout(n15907));
  jand g15616(.dina(n15904), .dinb(n15907), .dout(n15908));
  jnot g15617(.din(n15908), .dout(n15909));
  jand g15618(.dina(n15909), .dinb(n15906), .dout(n15910));
  jand g15619(.dina(n15910), .dinb(n15901), .dout(n15911));
  jor  g15620(.dina(n15911), .dinb(n15899), .dout(n15912));
  jand g15621(.dina(n15912), .dinb(asqrt[61] ), .dout(n15913));
  jxor g15622(.dina(n15306), .dinb(n290), .dout(n15914));
  jand g15623(.dina(n15914), .dinb(asqrt[10] ), .dout(n15915));
  jxor g15624(.dina(n15915), .dinb(n15316), .dout(n15916));
  jnot g15625(.din(n15916), .dout(n15917));
  jor  g15626(.dina(n15912), .dinb(asqrt[61] ), .dout(n15918));
  jand g15627(.dina(n15918), .dinb(n15917), .dout(n15919));
  jor  g15628(.dina(n15919), .dinb(n15913), .dout(n15920));
  jand g15629(.dina(n15920), .dinb(asqrt[62] ), .dout(n15921));
  jnot g15630(.din(n15321), .dout(n15922));
  jand g15631(.dina(n15922), .dinb(n15319), .dout(n15923));
  jand g15632(.dina(n15923), .dinb(asqrt[10] ), .dout(n15924));
  jxor g15633(.dina(n15924), .dinb(n15329), .dout(n15925));
  jnot g15634(.din(n15925), .dout(n15926));
  jor  g15635(.dina(n15913), .dinb(asqrt[62] ), .dout(n15927));
  jor  g15636(.dina(n15927), .dinb(n15919), .dout(n15928));
  jand g15637(.dina(n15928), .dinb(n15926), .dout(n15929));
  jor  g15638(.dina(n15929), .dinb(n15921), .dout(n15930));
  jxor g15639(.dina(n15331), .dinb(n199), .dout(n15931));
  jand g15640(.dina(n15931), .dinb(asqrt[10] ), .dout(n15932));
  jxor g15641(.dina(n15932), .dinb(n15336), .dout(n15933));
  jnot g15642(.din(n15338), .dout(n15934));
  jnot g15643(.din(n15342), .dout(n15935));
  jand g15644(.dina(asqrt[10] ), .dinb(n15935), .dout(n15936));
  jand g15645(.dina(n15936), .dinb(n15934), .dout(n15937));
  jor  g15646(.dina(n15937), .dinb(n15349), .dout(n15938));
  jor  g15647(.dina(n15938), .dinb(n15933), .dout(n15939));
  jnot g15648(.din(n15939), .dout(n15940));
  jand g15649(.dina(n15940), .dinb(n15930), .dout(n15941));
  jor  g15650(.dina(n15941), .dinb(asqrt[63] ), .dout(n15942));
  jnot g15651(.din(n15933), .dout(n15943));
  jor  g15652(.dina(n15943), .dinb(n15930), .dout(n15944));
  jor  g15653(.dina(n15936), .dinb(n15934), .dout(n15945));
  jand g15654(.dina(n15935), .dinb(n15934), .dout(n15946));
  jor  g15655(.dina(n15946), .dinb(n194), .dout(n15947));
  jnot g15656(.din(n15947), .dout(n15948));
  jand g15657(.dina(n15948), .dinb(n15945), .dout(n15949));
  jnot g15658(.din(asqrt[10] ), .dout(n15950));
  jnot g15659(.din(n15949), .dout(n15953));
  jand g15660(.dina(n15953), .dinb(n15944), .dout(n15954));
  jand g15661(.dina(n15954), .dinb(n15942), .dout(n15955));
  jxor g15662(.dina(n15822), .dinb(n796), .dout(n15956));
  jor  g15663(.dina(n15956), .dinb(n15955), .dout(n15957));
  jxor g15664(.dina(n15957), .dinb(n15362), .dout(n15958));
  jnot g15665(.din(n15958), .dout(n15959));
  jor  g15666(.dina(n15955), .dinb(n15364), .dout(n15960));
  jnot g15667(.din(a[16] ), .dout(n15961));
  jnot g15668(.din(a[17] ), .dout(n15962));
  jand g15669(.dina(n15364), .dinb(n15962), .dout(n15963));
  jand g15670(.dina(n15963), .dinb(n15961), .dout(n15964));
  jnot g15671(.din(n15964), .dout(n15965));
  jand g15672(.dina(n15965), .dinb(n15960), .dout(n15966));
  jor  g15673(.dina(n15966), .dinb(n15950), .dout(n15967));
  jor  g15674(.dina(n15955), .dinb(a[18] ), .dout(n15968));
  jxor g15675(.dina(n15968), .dinb(n15365), .dout(n15969));
  jand g15676(.dina(n15966), .dinb(n15950), .dout(n15970));
  jor  g15677(.dina(n15970), .dinb(n15969), .dout(n15971));
  jand g15678(.dina(n15971), .dinb(n15967), .dout(n15972));
  jor  g15679(.dina(n15972), .dinb(n14821), .dout(n15973));
  jand g15680(.dina(n15967), .dinb(n14821), .dout(n15974));
  jand g15681(.dina(n15974), .dinb(n15971), .dout(n15975));
  jor  g15682(.dina(n15968), .dinb(a[19] ), .dout(n15976));
  jnot g15683(.din(n15942), .dout(n15977));
  jnot g15684(.din(n15944), .dout(n15978));
  jor  g15685(.dina(n15949), .dinb(n15950), .dout(n15979));
  jor  g15686(.dina(n15979), .dinb(n15978), .dout(n15980));
  jor  g15687(.dina(n15980), .dinb(n15977), .dout(n15981));
  jand g15688(.dina(n15981), .dinb(n15976), .dout(n15982));
  jxor g15689(.dina(n15982), .dinb(n14826), .dout(n15983));
  jor  g15690(.dina(n15983), .dinb(n15975), .dout(n15984));
  jand g15691(.dina(n15984), .dinb(n15973), .dout(n15985));
  jor  g15692(.dina(n15985), .dinb(n14816), .dout(n15986));
  jand g15693(.dina(n15985), .dinb(n14816), .dout(n15987));
  jxor g15694(.dina(n15368), .dinb(n14821), .dout(n15988));
  jor  g15695(.dina(n15988), .dinb(n15955), .dout(n15989));
  jxor g15696(.dina(n15989), .dinb(n15371), .dout(n15990));
  jor  g15697(.dina(n15990), .dinb(n15987), .dout(n15991));
  jand g15698(.dina(n15991), .dinb(n15986), .dout(n15992));
  jor  g15699(.dina(n15992), .dinb(n13723), .dout(n15993));
  jnot g15700(.din(n15377), .dout(n15994));
  jor  g15701(.dina(n15994), .dinb(n15375), .dout(n15995));
  jor  g15702(.dina(n15995), .dinb(n15955), .dout(n15996));
  jxor g15703(.dina(n15996), .dinb(n15386), .dout(n15997));
  jand g15704(.dina(n15986), .dinb(n13723), .dout(n15998));
  jand g15705(.dina(n15998), .dinb(n15991), .dout(n15999));
  jor  g15706(.dina(n15999), .dinb(n15997), .dout(n16000));
  jand g15707(.dina(n16000), .dinb(n15993), .dout(n16001));
  jor  g15708(.dina(n16001), .dinb(n13718), .dout(n16002));
  jand g15709(.dina(n16001), .dinb(n13718), .dout(n16003));
  jxor g15710(.dina(n15388), .dinb(n13723), .dout(n16004));
  jor  g15711(.dina(n16004), .dinb(n15955), .dout(n16005));
  jxor g15712(.dina(n16005), .dinb(n15393), .dout(n16006));
  jnot g15713(.din(n16006), .dout(n16007));
  jor  g15714(.dina(n16007), .dinb(n16003), .dout(n16008));
  jand g15715(.dina(n16008), .dinb(n16002), .dout(n16009));
  jor  g15716(.dina(n16009), .dinb(n12675), .dout(n16010));
  jand g15717(.dina(n16002), .dinb(n12675), .dout(n16011));
  jand g15718(.dina(n16011), .dinb(n16008), .dout(n16012));
  jnot g15719(.din(n15397), .dout(n16013));
  jnot g15720(.din(n15955), .dout(asqrt[9] ));
  jand g15721(.dina(asqrt[9] ), .dinb(n16013), .dout(n16015));
  jand g15722(.dina(n16015), .dinb(n15404), .dout(n16016));
  jor  g15723(.dina(n16016), .dinb(n15402), .dout(n16017));
  jand g15724(.dina(n16015), .dinb(n15405), .dout(n16018));
  jnot g15725(.din(n16018), .dout(n16019));
  jand g15726(.dina(n16019), .dinb(n16017), .dout(n16020));
  jnot g15727(.din(n16020), .dout(n16021));
  jor  g15728(.dina(n16021), .dinb(n16012), .dout(n16022));
  jand g15729(.dina(n16022), .dinb(n16010), .dout(n16023));
  jor  g15730(.dina(n16023), .dinb(n12670), .dout(n16024));
  jand g15731(.dina(n16023), .dinb(n12670), .dout(n16025));
  jnot g15732(.din(n15412), .dout(n16026));
  jxor g15733(.dina(n15406), .dinb(n12675), .dout(n16027));
  jor  g15734(.dina(n16027), .dinb(n15955), .dout(n16028));
  jxor g15735(.dina(n16028), .dinb(n16026), .dout(n16029));
  jnot g15736(.din(n16029), .dout(n16030));
  jor  g15737(.dina(n16030), .dinb(n16025), .dout(n16031));
  jand g15738(.dina(n16031), .dinb(n16024), .dout(n16032));
  jor  g15739(.dina(n16032), .dinb(n11662), .dout(n16033));
  jnot g15740(.din(n15417), .dout(n16034));
  jor  g15741(.dina(n16034), .dinb(n15415), .dout(n16035));
  jor  g15742(.dina(n16035), .dinb(n15955), .dout(n16036));
  jxor g15743(.dina(n16036), .dinb(n15426), .dout(n16037));
  jand g15744(.dina(n16024), .dinb(n11662), .dout(n16038));
  jand g15745(.dina(n16038), .dinb(n16031), .dout(n16039));
  jor  g15746(.dina(n16039), .dinb(n16037), .dout(n16040));
  jand g15747(.dina(n16040), .dinb(n16033), .dout(n16041));
  jor  g15748(.dina(n16041), .dinb(n11657), .dout(n16042));
  jand g15749(.dina(n16041), .dinb(n11657), .dout(n16043));
  jnot g15750(.din(n15433), .dout(n16044));
  jxor g15751(.dina(n15428), .dinb(n11662), .dout(n16045));
  jor  g15752(.dina(n16045), .dinb(n15955), .dout(n16046));
  jxor g15753(.dina(n16046), .dinb(n16044), .dout(n16047));
  jnot g15754(.din(n16047), .dout(n16048));
  jor  g15755(.dina(n16048), .dinb(n16043), .dout(n16049));
  jand g15756(.dina(n16049), .dinb(n16042), .dout(n16050));
  jor  g15757(.dina(n16050), .dinb(n10701), .dout(n16051));
  jand g15758(.dina(n16042), .dinb(n10701), .dout(n16052));
  jand g15759(.dina(n16052), .dinb(n16049), .dout(n16053));
  jnot g15760(.din(n15436), .dout(n16054));
  jand g15761(.dina(asqrt[9] ), .dinb(n16054), .dout(n16055));
  jand g15762(.dina(n16055), .dinb(n15443), .dout(n16056));
  jor  g15763(.dina(n16056), .dinb(n15441), .dout(n16057));
  jand g15764(.dina(n16055), .dinb(n15444), .dout(n16058));
  jnot g15765(.din(n16058), .dout(n16059));
  jand g15766(.dina(n16059), .dinb(n16057), .dout(n16060));
  jnot g15767(.din(n16060), .dout(n16061));
  jor  g15768(.dina(n16061), .dinb(n16053), .dout(n16062));
  jand g15769(.dina(n16062), .dinb(n16051), .dout(n16063));
  jor  g15770(.dina(n16063), .dinb(n10696), .dout(n16064));
  jxor g15771(.dina(n15445), .dinb(n10701), .dout(n16065));
  jor  g15772(.dina(n16065), .dinb(n15955), .dout(n16066));
  jxor g15773(.dina(n16066), .dinb(n15450), .dout(n16067));
  jand g15774(.dina(n16063), .dinb(n10696), .dout(n16068));
  jor  g15775(.dina(n16068), .dinb(n16067), .dout(n16069));
  jand g15776(.dina(n16069), .dinb(n16064), .dout(n16070));
  jor  g15777(.dina(n16070), .dinb(n9774), .dout(n16071));
  jnot g15778(.din(n15455), .dout(n16072));
  jor  g15779(.dina(n16072), .dinb(n15453), .dout(n16073));
  jor  g15780(.dina(n16073), .dinb(n15955), .dout(n16074));
  jxor g15781(.dina(n16074), .dinb(n15464), .dout(n16075));
  jand g15782(.dina(n16064), .dinb(n9774), .dout(n16076));
  jand g15783(.dina(n16076), .dinb(n16069), .dout(n16077));
  jor  g15784(.dina(n16077), .dinb(n16075), .dout(n16078));
  jand g15785(.dina(n16078), .dinb(n16071), .dout(n16079));
  jor  g15786(.dina(n16079), .dinb(n9769), .dout(n16080));
  jand g15787(.dina(n16079), .dinb(n9769), .dout(n16081));
  jnot g15788(.din(n15467), .dout(n16082));
  jand g15789(.dina(asqrt[9] ), .dinb(n16082), .dout(n16083));
  jand g15790(.dina(n16083), .dinb(n15472), .dout(n16084));
  jor  g15791(.dina(n16084), .dinb(n15471), .dout(n16085));
  jand g15792(.dina(n16083), .dinb(n15473), .dout(n16086));
  jnot g15793(.din(n16086), .dout(n16087));
  jand g15794(.dina(n16087), .dinb(n16085), .dout(n16088));
  jnot g15795(.din(n16088), .dout(n16089));
  jor  g15796(.dina(n16089), .dinb(n16081), .dout(n16090));
  jand g15797(.dina(n16090), .dinb(n16080), .dout(n16091));
  jor  g15798(.dina(n16091), .dinb(n8898), .dout(n16092));
  jand g15799(.dina(n16080), .dinb(n8898), .dout(n16093));
  jand g15800(.dina(n16093), .dinb(n16090), .dout(n16094));
  jnot g15801(.din(n15475), .dout(n16095));
  jand g15802(.dina(asqrt[9] ), .dinb(n16095), .dout(n16096));
  jand g15803(.dina(n16096), .dinb(n15482), .dout(n16097));
  jor  g15804(.dina(n16097), .dinb(n15480), .dout(n16098));
  jand g15805(.dina(n16096), .dinb(n15483), .dout(n16099));
  jnot g15806(.din(n16099), .dout(n16100));
  jand g15807(.dina(n16100), .dinb(n16098), .dout(n16101));
  jnot g15808(.din(n16101), .dout(n16102));
  jor  g15809(.dina(n16102), .dinb(n16094), .dout(n16103));
  jand g15810(.dina(n16103), .dinb(n16092), .dout(n16104));
  jor  g15811(.dina(n16104), .dinb(n8893), .dout(n16105));
  jxor g15812(.dina(n15484), .dinb(n8898), .dout(n16106));
  jor  g15813(.dina(n16106), .dinb(n15955), .dout(n16107));
  jxor g15814(.dina(n16107), .dinb(n15495), .dout(n16108));
  jand g15815(.dina(n16104), .dinb(n8893), .dout(n16109));
  jor  g15816(.dina(n16109), .dinb(n16108), .dout(n16110));
  jand g15817(.dina(n16110), .dinb(n16105), .dout(n16111));
  jor  g15818(.dina(n16111), .dinb(n8058), .dout(n16112));
  jnot g15819(.din(n15500), .dout(n16113));
  jor  g15820(.dina(n16113), .dinb(n15498), .dout(n16114));
  jor  g15821(.dina(n16114), .dinb(n15955), .dout(n16115));
  jxor g15822(.dina(n16115), .dinb(n15509), .dout(n16116));
  jand g15823(.dina(n16105), .dinb(n8058), .dout(n16117));
  jand g15824(.dina(n16117), .dinb(n16110), .dout(n16118));
  jor  g15825(.dina(n16118), .dinb(n16116), .dout(n16119));
  jand g15826(.dina(n16119), .dinb(n16112), .dout(n16120));
  jor  g15827(.dina(n16120), .dinb(n8053), .dout(n16121));
  jand g15828(.dina(n16120), .dinb(n8053), .dout(n16122));
  jnot g15829(.din(n15512), .dout(n16123));
  jand g15830(.dina(asqrt[9] ), .dinb(n16123), .dout(n16124));
  jand g15831(.dina(n16124), .dinb(n15517), .dout(n16125));
  jor  g15832(.dina(n16125), .dinb(n15516), .dout(n16126));
  jand g15833(.dina(n16124), .dinb(n15518), .dout(n16127));
  jnot g15834(.din(n16127), .dout(n16128));
  jand g15835(.dina(n16128), .dinb(n16126), .dout(n16129));
  jnot g15836(.din(n16129), .dout(n16130));
  jor  g15837(.dina(n16130), .dinb(n16122), .dout(n16131));
  jand g15838(.dina(n16131), .dinb(n16121), .dout(n16132));
  jor  g15839(.dina(n16132), .dinb(n7265), .dout(n16133));
  jand g15840(.dina(n16121), .dinb(n7265), .dout(n16134));
  jand g15841(.dina(n16134), .dinb(n16131), .dout(n16135));
  jnot g15842(.din(n15520), .dout(n16136));
  jand g15843(.dina(asqrt[9] ), .dinb(n16136), .dout(n16137));
  jand g15844(.dina(n16137), .dinb(n15527), .dout(n16138));
  jor  g15845(.dina(n16138), .dinb(n15525), .dout(n16139));
  jand g15846(.dina(n16137), .dinb(n15528), .dout(n16140));
  jnot g15847(.din(n16140), .dout(n16141));
  jand g15848(.dina(n16141), .dinb(n16139), .dout(n16142));
  jnot g15849(.din(n16142), .dout(n16143));
  jor  g15850(.dina(n16143), .dinb(n16135), .dout(n16144));
  jand g15851(.dina(n16144), .dinb(n16133), .dout(n16145));
  jor  g15852(.dina(n16145), .dinb(n7260), .dout(n16146));
  jxor g15853(.dina(n15529), .dinb(n7265), .dout(n16147));
  jor  g15854(.dina(n16147), .dinb(n15955), .dout(n16148));
  jxor g15855(.dina(n16148), .dinb(n15540), .dout(n16149));
  jand g15856(.dina(n16145), .dinb(n7260), .dout(n16150));
  jor  g15857(.dina(n16150), .dinb(n16149), .dout(n16151));
  jand g15858(.dina(n16151), .dinb(n16146), .dout(n16152));
  jor  g15859(.dina(n16152), .dinb(n6505), .dout(n16153));
  jnot g15860(.din(n15545), .dout(n16154));
  jor  g15861(.dina(n16154), .dinb(n15543), .dout(n16155));
  jor  g15862(.dina(n16155), .dinb(n15955), .dout(n16156));
  jxor g15863(.dina(n16156), .dinb(n15554), .dout(n16157));
  jand g15864(.dina(n16146), .dinb(n6505), .dout(n16158));
  jand g15865(.dina(n16158), .dinb(n16151), .dout(n16159));
  jor  g15866(.dina(n16159), .dinb(n16157), .dout(n16160));
  jand g15867(.dina(n16160), .dinb(n16153), .dout(n16161));
  jor  g15868(.dina(n16161), .dinb(n6500), .dout(n16162));
  jand g15869(.dina(n16161), .dinb(n6500), .dout(n16163));
  jnot g15870(.din(n15557), .dout(n16164));
  jand g15871(.dina(asqrt[9] ), .dinb(n16164), .dout(n16165));
  jand g15872(.dina(n16165), .dinb(n15562), .dout(n16166));
  jor  g15873(.dina(n16166), .dinb(n15561), .dout(n16167));
  jand g15874(.dina(n16165), .dinb(n15563), .dout(n16168));
  jnot g15875(.din(n16168), .dout(n16169));
  jand g15876(.dina(n16169), .dinb(n16167), .dout(n16170));
  jnot g15877(.din(n16170), .dout(n16171));
  jor  g15878(.dina(n16171), .dinb(n16163), .dout(n16172));
  jand g15879(.dina(n16172), .dinb(n16162), .dout(n16173));
  jor  g15880(.dina(n16173), .dinb(n5793), .dout(n16174));
  jand g15881(.dina(n16162), .dinb(n5793), .dout(n16175));
  jand g15882(.dina(n16175), .dinb(n16172), .dout(n16176));
  jnot g15883(.din(n15565), .dout(n16177));
  jand g15884(.dina(asqrt[9] ), .dinb(n16177), .dout(n16178));
  jand g15885(.dina(n16178), .dinb(n15572), .dout(n16179));
  jor  g15886(.dina(n16179), .dinb(n15570), .dout(n16180));
  jand g15887(.dina(n16178), .dinb(n15573), .dout(n16181));
  jnot g15888(.din(n16181), .dout(n16182));
  jand g15889(.dina(n16182), .dinb(n16180), .dout(n16183));
  jnot g15890(.din(n16183), .dout(n16184));
  jor  g15891(.dina(n16184), .dinb(n16176), .dout(n16185));
  jand g15892(.dina(n16185), .dinb(n16174), .dout(n16186));
  jor  g15893(.dina(n16186), .dinb(n5788), .dout(n16187));
  jxor g15894(.dina(n15574), .dinb(n5793), .dout(n16188));
  jor  g15895(.dina(n16188), .dinb(n15955), .dout(n16189));
  jxor g15896(.dina(n16189), .dinb(n15585), .dout(n16190));
  jand g15897(.dina(n16186), .dinb(n5788), .dout(n16191));
  jor  g15898(.dina(n16191), .dinb(n16190), .dout(n16192));
  jand g15899(.dina(n16192), .dinb(n16187), .dout(n16193));
  jor  g15900(.dina(n16193), .dinb(n5121), .dout(n16194));
  jnot g15901(.din(n15590), .dout(n16195));
  jor  g15902(.dina(n16195), .dinb(n15588), .dout(n16196));
  jor  g15903(.dina(n16196), .dinb(n15955), .dout(n16197));
  jxor g15904(.dina(n16197), .dinb(n15599), .dout(n16198));
  jand g15905(.dina(n16187), .dinb(n5121), .dout(n16199));
  jand g15906(.dina(n16199), .dinb(n16192), .dout(n16200));
  jor  g15907(.dina(n16200), .dinb(n16198), .dout(n16201));
  jand g15908(.dina(n16201), .dinb(n16194), .dout(n16202));
  jor  g15909(.dina(n16202), .dinb(n5116), .dout(n16203));
  jand g15910(.dina(n16202), .dinb(n5116), .dout(n16204));
  jnot g15911(.din(n15602), .dout(n16205));
  jand g15912(.dina(asqrt[9] ), .dinb(n16205), .dout(n16206));
  jand g15913(.dina(n16206), .dinb(n15607), .dout(n16207));
  jor  g15914(.dina(n16207), .dinb(n15606), .dout(n16208));
  jand g15915(.dina(n16206), .dinb(n15608), .dout(n16209));
  jnot g15916(.din(n16209), .dout(n16210));
  jand g15917(.dina(n16210), .dinb(n16208), .dout(n16211));
  jnot g15918(.din(n16211), .dout(n16212));
  jor  g15919(.dina(n16212), .dinb(n16204), .dout(n16213));
  jand g15920(.dina(n16213), .dinb(n16203), .dout(n16214));
  jor  g15921(.dina(n16214), .dinb(n4499), .dout(n16215));
  jand g15922(.dina(n16203), .dinb(n4499), .dout(n16216));
  jand g15923(.dina(n16216), .dinb(n16213), .dout(n16217));
  jnot g15924(.din(n15610), .dout(n16218));
  jand g15925(.dina(asqrt[9] ), .dinb(n16218), .dout(n16219));
  jand g15926(.dina(n16219), .dinb(n15617), .dout(n16220));
  jor  g15927(.dina(n16220), .dinb(n15615), .dout(n16221));
  jand g15928(.dina(n16219), .dinb(n15618), .dout(n16222));
  jnot g15929(.din(n16222), .dout(n16223));
  jand g15930(.dina(n16223), .dinb(n16221), .dout(n16224));
  jnot g15931(.din(n16224), .dout(n16225));
  jor  g15932(.dina(n16225), .dinb(n16217), .dout(n16226));
  jand g15933(.dina(n16226), .dinb(n16215), .dout(n16227));
  jor  g15934(.dina(n16227), .dinb(n4494), .dout(n16228));
  jxor g15935(.dina(n15619), .dinb(n4499), .dout(n16229));
  jor  g15936(.dina(n16229), .dinb(n15955), .dout(n16230));
  jxor g15937(.dina(n16230), .dinb(n15630), .dout(n16231));
  jand g15938(.dina(n16227), .dinb(n4494), .dout(n16232));
  jor  g15939(.dina(n16232), .dinb(n16231), .dout(n16233));
  jand g15940(.dina(n16233), .dinb(n16228), .dout(n16234));
  jor  g15941(.dina(n16234), .dinb(n3912), .dout(n16235));
  jnot g15942(.din(n15635), .dout(n16236));
  jor  g15943(.dina(n16236), .dinb(n15633), .dout(n16237));
  jor  g15944(.dina(n16237), .dinb(n15955), .dout(n16238));
  jxor g15945(.dina(n16238), .dinb(n15644), .dout(n16239));
  jand g15946(.dina(n16228), .dinb(n3912), .dout(n16240));
  jand g15947(.dina(n16240), .dinb(n16233), .dout(n16241));
  jor  g15948(.dina(n16241), .dinb(n16239), .dout(n16242));
  jand g15949(.dina(n16242), .dinb(n16235), .dout(n16243));
  jor  g15950(.dina(n16243), .dinb(n3907), .dout(n16244));
  jand g15951(.dina(n16243), .dinb(n3907), .dout(n16245));
  jnot g15952(.din(n15647), .dout(n16246));
  jand g15953(.dina(asqrt[9] ), .dinb(n16246), .dout(n16247));
  jand g15954(.dina(n16247), .dinb(n15652), .dout(n16248));
  jor  g15955(.dina(n16248), .dinb(n15651), .dout(n16249));
  jand g15956(.dina(n16247), .dinb(n15653), .dout(n16250));
  jnot g15957(.din(n16250), .dout(n16251));
  jand g15958(.dina(n16251), .dinb(n16249), .dout(n16252));
  jnot g15959(.din(n16252), .dout(n16253));
  jor  g15960(.dina(n16253), .dinb(n16245), .dout(n16254));
  jand g15961(.dina(n16254), .dinb(n16244), .dout(n16255));
  jor  g15962(.dina(n16255), .dinb(n3376), .dout(n16256));
  jand g15963(.dina(n16244), .dinb(n3376), .dout(n16257));
  jand g15964(.dina(n16257), .dinb(n16254), .dout(n16258));
  jnot g15965(.din(n15655), .dout(n16259));
  jand g15966(.dina(asqrt[9] ), .dinb(n16259), .dout(n16260));
  jand g15967(.dina(n16260), .dinb(n15662), .dout(n16261));
  jor  g15968(.dina(n16261), .dinb(n15660), .dout(n16262));
  jand g15969(.dina(n16260), .dinb(n15663), .dout(n16263));
  jnot g15970(.din(n16263), .dout(n16264));
  jand g15971(.dina(n16264), .dinb(n16262), .dout(n16265));
  jnot g15972(.din(n16265), .dout(n16266));
  jor  g15973(.dina(n16266), .dinb(n16258), .dout(n16267));
  jand g15974(.dina(n16267), .dinb(n16256), .dout(n16268));
  jor  g15975(.dina(n16268), .dinb(n3371), .dout(n16269));
  jxor g15976(.dina(n15664), .dinb(n3376), .dout(n16270));
  jor  g15977(.dina(n16270), .dinb(n15955), .dout(n16271));
  jxor g15978(.dina(n16271), .dinb(n15675), .dout(n16272));
  jand g15979(.dina(n16268), .dinb(n3371), .dout(n16273));
  jor  g15980(.dina(n16273), .dinb(n16272), .dout(n16274));
  jand g15981(.dina(n16274), .dinb(n16269), .dout(n16275));
  jor  g15982(.dina(n16275), .dinb(n2875), .dout(n16276));
  jnot g15983(.din(n15680), .dout(n16277));
  jor  g15984(.dina(n16277), .dinb(n15678), .dout(n16278));
  jor  g15985(.dina(n16278), .dinb(n15955), .dout(n16279));
  jxor g15986(.dina(n16279), .dinb(n15689), .dout(n16280));
  jand g15987(.dina(n16269), .dinb(n2875), .dout(n16281));
  jand g15988(.dina(n16281), .dinb(n16274), .dout(n16282));
  jor  g15989(.dina(n16282), .dinb(n16280), .dout(n16283));
  jand g15990(.dina(n16283), .dinb(n16276), .dout(n16284));
  jor  g15991(.dina(n16284), .dinb(n2870), .dout(n16285));
  jand g15992(.dina(n16284), .dinb(n2870), .dout(n16286));
  jnot g15993(.din(n15692), .dout(n16287));
  jand g15994(.dina(asqrt[9] ), .dinb(n16287), .dout(n16288));
  jand g15995(.dina(n16288), .dinb(n15697), .dout(n16289));
  jor  g15996(.dina(n16289), .dinb(n15696), .dout(n16290));
  jand g15997(.dina(n16288), .dinb(n15698), .dout(n16291));
  jnot g15998(.din(n16291), .dout(n16292));
  jand g15999(.dina(n16292), .dinb(n16290), .dout(n16293));
  jnot g16000(.din(n16293), .dout(n16294));
  jor  g16001(.dina(n16294), .dinb(n16286), .dout(n16295));
  jand g16002(.dina(n16295), .dinb(n16285), .dout(n16296));
  jor  g16003(.dina(n16296), .dinb(n2425), .dout(n16297));
  jand g16004(.dina(n16285), .dinb(n2425), .dout(n16298));
  jand g16005(.dina(n16298), .dinb(n16295), .dout(n16299));
  jnot g16006(.din(n15700), .dout(n16300));
  jand g16007(.dina(asqrt[9] ), .dinb(n16300), .dout(n16301));
  jand g16008(.dina(n16301), .dinb(n15707), .dout(n16302));
  jor  g16009(.dina(n16302), .dinb(n15705), .dout(n16303));
  jand g16010(.dina(n16301), .dinb(n15708), .dout(n16304));
  jnot g16011(.din(n16304), .dout(n16305));
  jand g16012(.dina(n16305), .dinb(n16303), .dout(n16306));
  jnot g16013(.din(n16306), .dout(n16307));
  jor  g16014(.dina(n16307), .dinb(n16299), .dout(n16308));
  jand g16015(.dina(n16308), .dinb(n16297), .dout(n16309));
  jor  g16016(.dina(n16309), .dinb(n2420), .dout(n16310));
  jxor g16017(.dina(n15709), .dinb(n2425), .dout(n16311));
  jor  g16018(.dina(n16311), .dinb(n15955), .dout(n16312));
  jxor g16019(.dina(n16312), .dinb(n15720), .dout(n16313));
  jand g16020(.dina(n16309), .dinb(n2420), .dout(n16314));
  jor  g16021(.dina(n16314), .dinb(n16313), .dout(n16315));
  jand g16022(.dina(n16315), .dinb(n16310), .dout(n16316));
  jor  g16023(.dina(n16316), .dinb(n2010), .dout(n16317));
  jnot g16024(.din(n15725), .dout(n16318));
  jor  g16025(.dina(n16318), .dinb(n15723), .dout(n16319));
  jor  g16026(.dina(n16319), .dinb(n15955), .dout(n16320));
  jxor g16027(.dina(n16320), .dinb(n15734), .dout(n16321));
  jand g16028(.dina(n16310), .dinb(n2010), .dout(n16322));
  jand g16029(.dina(n16322), .dinb(n16315), .dout(n16323));
  jor  g16030(.dina(n16323), .dinb(n16321), .dout(n16324));
  jand g16031(.dina(n16324), .dinb(n16317), .dout(n16325));
  jor  g16032(.dina(n16325), .dinb(n2005), .dout(n16326));
  jand g16033(.dina(n16325), .dinb(n2005), .dout(n16327));
  jnot g16034(.din(n15737), .dout(n16328));
  jand g16035(.dina(asqrt[9] ), .dinb(n16328), .dout(n16329));
  jand g16036(.dina(n16329), .dinb(n15742), .dout(n16330));
  jor  g16037(.dina(n16330), .dinb(n15741), .dout(n16331));
  jand g16038(.dina(n16329), .dinb(n15743), .dout(n16332));
  jnot g16039(.din(n16332), .dout(n16333));
  jand g16040(.dina(n16333), .dinb(n16331), .dout(n16334));
  jnot g16041(.din(n16334), .dout(n16335));
  jor  g16042(.dina(n16335), .dinb(n16327), .dout(n16336));
  jand g16043(.dina(n16336), .dinb(n16326), .dout(n16337));
  jor  g16044(.dina(n16337), .dinb(n1646), .dout(n16338));
  jand g16045(.dina(n16326), .dinb(n1646), .dout(n16339));
  jand g16046(.dina(n16339), .dinb(n16336), .dout(n16340));
  jnot g16047(.din(n15745), .dout(n16341));
  jand g16048(.dina(asqrt[9] ), .dinb(n16341), .dout(n16342));
  jand g16049(.dina(n16342), .dinb(n15752), .dout(n16343));
  jor  g16050(.dina(n16343), .dinb(n15750), .dout(n16344));
  jand g16051(.dina(n16342), .dinb(n15753), .dout(n16345));
  jnot g16052(.din(n16345), .dout(n16346));
  jand g16053(.dina(n16346), .dinb(n16344), .dout(n16347));
  jnot g16054(.din(n16347), .dout(n16348));
  jor  g16055(.dina(n16348), .dinb(n16340), .dout(n16349));
  jand g16056(.dina(n16349), .dinb(n16338), .dout(n16350));
  jor  g16057(.dina(n16350), .dinb(n1641), .dout(n16351));
  jxor g16058(.dina(n15754), .dinb(n1646), .dout(n16352));
  jor  g16059(.dina(n16352), .dinb(n15955), .dout(n16353));
  jxor g16060(.dina(n16353), .dinb(n15765), .dout(n16354));
  jand g16061(.dina(n16350), .dinb(n1641), .dout(n16355));
  jor  g16062(.dina(n16355), .dinb(n16354), .dout(n16356));
  jand g16063(.dina(n16356), .dinb(n16351), .dout(n16357));
  jor  g16064(.dina(n16357), .dinb(n1317), .dout(n16358));
  jnot g16065(.din(n15770), .dout(n16359));
  jor  g16066(.dina(n16359), .dinb(n15768), .dout(n16360));
  jor  g16067(.dina(n16360), .dinb(n15955), .dout(n16361));
  jxor g16068(.dina(n16361), .dinb(n15779), .dout(n16362));
  jand g16069(.dina(n16351), .dinb(n1317), .dout(n16363));
  jand g16070(.dina(n16363), .dinb(n16356), .dout(n16364));
  jor  g16071(.dina(n16364), .dinb(n16362), .dout(n16365));
  jand g16072(.dina(n16365), .dinb(n16358), .dout(n16366));
  jor  g16073(.dina(n16366), .dinb(n1312), .dout(n16367));
  jand g16074(.dina(n16366), .dinb(n1312), .dout(n16368));
  jnot g16075(.din(n15782), .dout(n16369));
  jand g16076(.dina(asqrt[9] ), .dinb(n16369), .dout(n16370));
  jand g16077(.dina(n16370), .dinb(n15787), .dout(n16371));
  jor  g16078(.dina(n16371), .dinb(n15786), .dout(n16372));
  jand g16079(.dina(n16370), .dinb(n15788), .dout(n16373));
  jnot g16080(.din(n16373), .dout(n16374));
  jand g16081(.dina(n16374), .dinb(n16372), .dout(n16375));
  jnot g16082(.din(n16375), .dout(n16376));
  jor  g16083(.dina(n16376), .dinb(n16368), .dout(n16377));
  jand g16084(.dina(n16377), .dinb(n16367), .dout(n16378));
  jor  g16085(.dina(n16378), .dinb(n1039), .dout(n16379));
  jand g16086(.dina(n16367), .dinb(n1039), .dout(n16380));
  jand g16087(.dina(n16380), .dinb(n16377), .dout(n16381));
  jnot g16088(.din(n15790), .dout(n16382));
  jand g16089(.dina(asqrt[9] ), .dinb(n16382), .dout(n16383));
  jand g16090(.dina(n16383), .dinb(n15797), .dout(n16384));
  jor  g16091(.dina(n16384), .dinb(n15795), .dout(n16385));
  jand g16092(.dina(n16383), .dinb(n15798), .dout(n16386));
  jnot g16093(.din(n16386), .dout(n16387));
  jand g16094(.dina(n16387), .dinb(n16385), .dout(n16388));
  jnot g16095(.din(n16388), .dout(n16389));
  jor  g16096(.dina(n16389), .dinb(n16381), .dout(n16390));
  jand g16097(.dina(n16390), .dinb(n16379), .dout(n16391));
  jor  g16098(.dina(n16391), .dinb(n1034), .dout(n16392));
  jxor g16099(.dina(n15799), .dinb(n1039), .dout(n16393));
  jor  g16100(.dina(n16393), .dinb(n15955), .dout(n16394));
  jxor g16101(.dina(n16394), .dinb(n15810), .dout(n16395));
  jand g16102(.dina(n16391), .dinb(n1034), .dout(n16396));
  jor  g16103(.dina(n16396), .dinb(n16395), .dout(n16397));
  jand g16104(.dina(n16397), .dinb(n16392), .dout(n16398));
  jor  g16105(.dina(n16398), .dinb(n796), .dout(n16399));
  jand g16106(.dina(n16392), .dinb(n796), .dout(n16400));
  jand g16107(.dina(n16400), .dinb(n16397), .dout(n16401));
  jnot g16108(.din(n15813), .dout(n16402));
  jand g16109(.dina(asqrt[9] ), .dinb(n16402), .dout(n16403));
  jand g16110(.dina(n16403), .dinb(n15820), .dout(n16404));
  jor  g16111(.dina(n16404), .dinb(n15818), .dout(n16405));
  jand g16112(.dina(n16403), .dinb(n15821), .dout(n16406));
  jnot g16113(.din(n16406), .dout(n16407));
  jand g16114(.dina(n16407), .dinb(n16405), .dout(n16408));
  jnot g16115(.din(n16408), .dout(n16409));
  jor  g16116(.dina(n16409), .dinb(n16401), .dout(n16410));
  jand g16117(.dina(n16410), .dinb(n16399), .dout(n16411));
  jor  g16118(.dina(n16411), .dinb(n791), .dout(n16412));
  jand g16119(.dina(n16411), .dinb(n791), .dout(n16413));
  jor  g16120(.dina(n16413), .dinb(n15959), .dout(n16414));
  jand g16121(.dina(n16414), .dinb(n16412), .dout(n16415));
  jor  g16122(.dina(n16415), .dinb(n595), .dout(n16416));
  jnot g16123(.din(n15829), .dout(n16417));
  jor  g16124(.dina(n16417), .dinb(n15827), .dout(n16418));
  jor  g16125(.dina(n16418), .dinb(n15955), .dout(n16419));
  jxor g16126(.dina(n16419), .dinb(n15838), .dout(n16420));
  jand g16127(.dina(n16412), .dinb(n595), .dout(n16421));
  jand g16128(.dina(n16421), .dinb(n16414), .dout(n16422));
  jor  g16129(.dina(n16422), .dinb(n16420), .dout(n16423));
  jand g16130(.dina(n16423), .dinb(n16416), .dout(n16424));
  jor  g16131(.dina(n16424), .dinb(n590), .dout(n16425));
  jxor g16132(.dina(n15840), .dinb(n595), .dout(n16426));
  jor  g16133(.dina(n16426), .dinb(n15955), .dout(n16427));
  jxor g16134(.dina(n16427), .dinb(n15851), .dout(n16428));
  jand g16135(.dina(n16424), .dinb(n590), .dout(n16429));
  jor  g16136(.dina(n16429), .dinb(n16428), .dout(n16430));
  jand g16137(.dina(n16430), .dinb(n16425), .dout(n16431));
  jor  g16138(.dina(n16431), .dinb(n430), .dout(n16432));
  jnot g16139(.din(n15856), .dout(n16433));
  jor  g16140(.dina(n16433), .dinb(n15854), .dout(n16434));
  jor  g16141(.dina(n16434), .dinb(n15955), .dout(n16435));
  jxor g16142(.dina(n16435), .dinb(n15865), .dout(n16436));
  jand g16143(.dina(n16425), .dinb(n430), .dout(n16437));
  jand g16144(.dina(n16437), .dinb(n16430), .dout(n16438));
  jor  g16145(.dina(n16438), .dinb(n16436), .dout(n16439));
  jand g16146(.dina(n16439), .dinb(n16432), .dout(n16440));
  jor  g16147(.dina(n16440), .dinb(n425), .dout(n16441));
  jand g16148(.dina(n16440), .dinb(n425), .dout(n16442));
  jnot g16149(.din(n15868), .dout(n16443));
  jand g16150(.dina(asqrt[9] ), .dinb(n16443), .dout(n16444));
  jand g16151(.dina(n16444), .dinb(n15873), .dout(n16445));
  jor  g16152(.dina(n16445), .dinb(n15872), .dout(n16446));
  jand g16153(.dina(n16444), .dinb(n15874), .dout(n16447));
  jnot g16154(.din(n16447), .dout(n16448));
  jand g16155(.dina(n16448), .dinb(n16446), .dout(n16449));
  jnot g16156(.din(n16449), .dout(n16450));
  jor  g16157(.dina(n16450), .dinb(n16442), .dout(n16451));
  jand g16158(.dina(n16451), .dinb(n16441), .dout(n16452));
  jor  g16159(.dina(n16452), .dinb(n305), .dout(n16453));
  jand g16160(.dina(n16441), .dinb(n305), .dout(n16454));
  jand g16161(.dina(n16454), .dinb(n16451), .dout(n16455));
  jnot g16162(.din(n15876), .dout(n16456));
  jand g16163(.dina(asqrt[9] ), .dinb(n16456), .dout(n16457));
  jand g16164(.dina(n16457), .dinb(n15883), .dout(n16458));
  jor  g16165(.dina(n16458), .dinb(n15881), .dout(n16459));
  jand g16166(.dina(n16457), .dinb(n15884), .dout(n16460));
  jnot g16167(.din(n16460), .dout(n16461));
  jand g16168(.dina(n16461), .dinb(n16459), .dout(n16462));
  jnot g16169(.din(n16462), .dout(n16463));
  jor  g16170(.dina(n16463), .dinb(n16455), .dout(n16464));
  jand g16171(.dina(n16464), .dinb(n16453), .dout(n16465));
  jor  g16172(.dina(n16465), .dinb(n290), .dout(n16466));
  jxor g16173(.dina(n15885), .dinb(n305), .dout(n16467));
  jor  g16174(.dina(n16467), .dinb(n15955), .dout(n16468));
  jxor g16175(.dina(n16468), .dinb(n15896), .dout(n16469));
  jand g16176(.dina(n16465), .dinb(n290), .dout(n16470));
  jor  g16177(.dina(n16470), .dinb(n16469), .dout(n16471));
  jand g16178(.dina(n16471), .dinb(n16466), .dout(n16472));
  jor  g16179(.dina(n16472), .dinb(n223), .dout(n16473));
  jnot g16180(.din(n15901), .dout(n16474));
  jor  g16181(.dina(n16474), .dinb(n15899), .dout(n16475));
  jor  g16182(.dina(n16475), .dinb(n15955), .dout(n16476));
  jxor g16183(.dina(n16476), .dinb(n15910), .dout(n16477));
  jand g16184(.dina(n16466), .dinb(n223), .dout(n16478));
  jand g16185(.dina(n16478), .dinb(n16471), .dout(n16479));
  jor  g16186(.dina(n16479), .dinb(n16477), .dout(n16480));
  jand g16187(.dina(n16480), .dinb(n16473), .dout(n16481));
  jor  g16188(.dina(n16481), .dinb(n199), .dout(n16482));
  jand g16189(.dina(n16481), .dinb(n199), .dout(n16483));
  jnot g16190(.din(n15913), .dout(n16484));
  jand g16191(.dina(asqrt[9] ), .dinb(n16484), .dout(n16485));
  jand g16192(.dina(n16485), .dinb(n15918), .dout(n16486));
  jor  g16193(.dina(n16486), .dinb(n15917), .dout(n16487));
  jand g16194(.dina(n16485), .dinb(n15919), .dout(n16488));
  jnot g16195(.din(n16488), .dout(n16489));
  jand g16196(.dina(n16489), .dinb(n16487), .dout(n16490));
  jnot g16197(.din(n16490), .dout(n16491));
  jor  g16198(.dina(n16491), .dinb(n16483), .dout(n16492));
  jand g16199(.dina(n16492), .dinb(n16482), .dout(n16493));
  jnot g16200(.din(n15921), .dout(n16494));
  jand g16201(.dina(asqrt[9] ), .dinb(n16494), .dout(n16495));
  jand g16202(.dina(n16495), .dinb(n15928), .dout(n16496));
  jor  g16203(.dina(n16496), .dinb(n15926), .dout(n16497));
  jand g16204(.dina(n16495), .dinb(n15929), .dout(n16498));
  jnot g16205(.din(n16498), .dout(n16499));
  jand g16206(.dina(n16499), .dinb(n16497), .dout(n16500));
  jnot g16207(.din(n16500), .dout(n16501));
  jand g16208(.dina(asqrt[9] ), .dinb(n15943), .dout(n16502));
  jand g16209(.dina(n16502), .dinb(n15930), .dout(n16503));
  jor  g16210(.dina(n16503), .dinb(n15978), .dout(n16504));
  jor  g16211(.dina(n16504), .dinb(n16501), .dout(n16505));
  jor  g16212(.dina(n16505), .dinb(n16493), .dout(n16506));
  jand g16213(.dina(n16506), .dinb(n194), .dout(n16507));
  jand g16214(.dina(n16501), .dinb(n16493), .dout(n16508));
  jor  g16215(.dina(n16502), .dinb(n15930), .dout(n16509));
  jand g16216(.dina(n15943), .dinb(n15930), .dout(n16510));
  jor  g16217(.dina(n16510), .dinb(n194), .dout(n16511));
  jnot g16218(.din(n16511), .dout(n16512));
  jand g16219(.dina(n16512), .dinb(n16509), .dout(n16513));
  jor  g16220(.dina(n16513), .dinb(n16508), .dout(n16516));
  jor  g16221(.dina(n16516), .dinb(n16507), .dout(asqrt[8] ));
  jxor g16222(.dina(n16411), .dinb(n791), .dout(n16518));
  jand g16223(.dina(n16518), .dinb(asqrt[8] ), .dout(n16519));
  jxor g16224(.dina(n16519), .dinb(n15959), .dout(n16520));
  jnot g16225(.din(n16520), .dout(n16521));
  jand g16226(.dina(asqrt[8] ), .dinb(a[16] ), .dout(n16522));
  jnot g16227(.din(a[14] ), .dout(n16523));
  jnot g16228(.din(a[15] ), .dout(n16524));
  jand g16229(.dina(n15961), .dinb(n16524), .dout(n16525));
  jand g16230(.dina(n16525), .dinb(n16523), .dout(n16526));
  jor  g16231(.dina(n16526), .dinb(n16522), .dout(n16527));
  jand g16232(.dina(n16527), .dinb(asqrt[9] ), .dout(n16528));
  jand g16233(.dina(asqrt[8] ), .dinb(n15961), .dout(n16529));
  jxor g16234(.dina(n16529), .dinb(n15962), .dout(n16530));
  jor  g16235(.dina(n16527), .dinb(asqrt[9] ), .dout(n16531));
  jand g16236(.dina(n16531), .dinb(n16530), .dout(n16532));
  jor  g16237(.dina(n16532), .dinb(n16528), .dout(n16533));
  jand g16238(.dina(n16533), .dinb(asqrt[10] ), .dout(n16534));
  jor  g16239(.dina(n16528), .dinb(asqrt[10] ), .dout(n16535));
  jor  g16240(.dina(n16535), .dinb(n16532), .dout(n16536));
  jand g16241(.dina(n16529), .dinb(n15962), .dout(n16537));
  jnot g16242(.din(n16507), .dout(n16538));
  jnot g16243(.din(n16508), .dout(n16539));
  jnot g16244(.din(n16513), .dout(n16540));
  jand g16245(.dina(n16540), .dinb(asqrt[9] ), .dout(n16541));
  jand g16246(.dina(n16541), .dinb(n16539), .dout(n16542));
  jand g16247(.dina(n16542), .dinb(n16538), .dout(n16543));
  jor  g16248(.dina(n16543), .dinb(n16537), .dout(n16544));
  jxor g16249(.dina(n16544), .dinb(n15364), .dout(n16545));
  jand g16250(.dina(n16545), .dinb(n16536), .dout(n16546));
  jor  g16251(.dina(n16546), .dinb(n16534), .dout(n16547));
  jand g16252(.dina(n16547), .dinb(asqrt[11] ), .dout(n16548));
  jor  g16253(.dina(n16547), .dinb(asqrt[11] ), .dout(n16549));
  jxor g16254(.dina(n15966), .dinb(n15950), .dout(n16550));
  jand g16255(.dina(n16550), .dinb(asqrt[8] ), .dout(n16551));
  jxor g16256(.dina(n16551), .dinb(n15969), .dout(n16552));
  jnot g16257(.din(n16552), .dout(n16553));
  jand g16258(.dina(n16553), .dinb(n16549), .dout(n16554));
  jor  g16259(.dina(n16554), .dinb(n16548), .dout(n16555));
  jand g16260(.dina(n16555), .dinb(asqrt[12] ), .dout(n16556));
  jnot g16261(.din(n15975), .dout(n16557));
  jand g16262(.dina(n16557), .dinb(n15973), .dout(n16558));
  jand g16263(.dina(n16558), .dinb(asqrt[8] ), .dout(n16559));
  jxor g16264(.dina(n16559), .dinb(n15983), .dout(n16560));
  jnot g16265(.din(n16560), .dout(n16561));
  jor  g16266(.dina(n16548), .dinb(asqrt[12] ), .dout(n16562));
  jor  g16267(.dina(n16562), .dinb(n16554), .dout(n16563));
  jand g16268(.dina(n16563), .dinb(n16561), .dout(n16564));
  jor  g16269(.dina(n16564), .dinb(n16556), .dout(n16565));
  jand g16270(.dina(n16565), .dinb(asqrt[13] ), .dout(n16566));
  jor  g16271(.dina(n16565), .dinb(asqrt[13] ), .dout(n16567));
  jnot g16272(.din(n15990), .dout(n16568));
  jxor g16273(.dina(n15985), .dinb(n14816), .dout(n16569));
  jand g16274(.dina(n16569), .dinb(asqrt[8] ), .dout(n16570));
  jxor g16275(.dina(n16570), .dinb(n16568), .dout(n16571));
  jand g16276(.dina(n16571), .dinb(n16567), .dout(n16572));
  jor  g16277(.dina(n16572), .dinb(n16566), .dout(n16573));
  jand g16278(.dina(n16573), .dinb(asqrt[14] ), .dout(n16574));
  jor  g16279(.dina(n16566), .dinb(asqrt[14] ), .dout(n16575));
  jor  g16280(.dina(n16575), .dinb(n16572), .dout(n16576));
  jnot g16281(.din(n15997), .dout(n16577));
  jnot g16282(.din(n15999), .dout(n16578));
  jand g16283(.dina(asqrt[8] ), .dinb(n15993), .dout(n16579));
  jand g16284(.dina(n16579), .dinb(n16578), .dout(n16580));
  jor  g16285(.dina(n16580), .dinb(n16577), .dout(n16581));
  jnot g16286(.din(n16000), .dout(n16582));
  jand g16287(.dina(n16579), .dinb(n16582), .dout(n16583));
  jnot g16288(.din(n16583), .dout(n16584));
  jand g16289(.dina(n16584), .dinb(n16581), .dout(n16585));
  jand g16290(.dina(n16585), .dinb(n16576), .dout(n16586));
  jor  g16291(.dina(n16586), .dinb(n16574), .dout(n16587));
  jand g16292(.dina(n16587), .dinb(asqrt[15] ), .dout(n16588));
  jor  g16293(.dina(n16587), .dinb(asqrt[15] ), .dout(n16589));
  jxor g16294(.dina(n16001), .dinb(n13718), .dout(n16590));
  jand g16295(.dina(n16590), .dinb(asqrt[8] ), .dout(n16591));
  jxor g16296(.dina(n16591), .dinb(n16006), .dout(n16592));
  jand g16297(.dina(n16592), .dinb(n16589), .dout(n16593));
  jor  g16298(.dina(n16593), .dinb(n16588), .dout(n16594));
  jand g16299(.dina(n16594), .dinb(asqrt[16] ), .dout(n16595));
  jnot g16300(.din(n16012), .dout(n16596));
  jand g16301(.dina(n16596), .dinb(n16010), .dout(n16597));
  jand g16302(.dina(n16597), .dinb(asqrt[8] ), .dout(n16598));
  jxor g16303(.dina(n16598), .dinb(n16021), .dout(n16599));
  jnot g16304(.din(n16599), .dout(n16600));
  jor  g16305(.dina(n16588), .dinb(asqrt[16] ), .dout(n16601));
  jor  g16306(.dina(n16601), .dinb(n16593), .dout(n16602));
  jand g16307(.dina(n16602), .dinb(n16600), .dout(n16603));
  jor  g16308(.dina(n16603), .dinb(n16595), .dout(n16604));
  jand g16309(.dina(n16604), .dinb(asqrt[17] ), .dout(n16605));
  jor  g16310(.dina(n16604), .dinb(asqrt[17] ), .dout(n16606));
  jxor g16311(.dina(n16023), .dinb(n12670), .dout(n16607));
  jand g16312(.dina(n16607), .dinb(asqrt[8] ), .dout(n16608));
  jxor g16313(.dina(n16608), .dinb(n16029), .dout(n16609));
  jand g16314(.dina(n16609), .dinb(n16606), .dout(n16610));
  jor  g16315(.dina(n16610), .dinb(n16605), .dout(n16611));
  jand g16316(.dina(n16611), .dinb(asqrt[18] ), .dout(n16612));
  jor  g16317(.dina(n16605), .dinb(asqrt[18] ), .dout(n16613));
  jor  g16318(.dina(n16613), .dinb(n16610), .dout(n16614));
  jnot g16319(.din(n16037), .dout(n16615));
  jnot g16320(.din(n16039), .dout(n16616));
  jand g16321(.dina(asqrt[8] ), .dinb(n16033), .dout(n16617));
  jand g16322(.dina(n16617), .dinb(n16616), .dout(n16618));
  jor  g16323(.dina(n16618), .dinb(n16615), .dout(n16619));
  jnot g16324(.din(n16040), .dout(n16620));
  jand g16325(.dina(n16617), .dinb(n16620), .dout(n16621));
  jnot g16326(.din(n16621), .dout(n16622));
  jand g16327(.dina(n16622), .dinb(n16619), .dout(n16623));
  jand g16328(.dina(n16623), .dinb(n16614), .dout(n16624));
  jor  g16329(.dina(n16624), .dinb(n16612), .dout(n16625));
  jand g16330(.dina(n16625), .dinb(asqrt[19] ), .dout(n16626));
  jxor g16331(.dina(n16041), .dinb(n11657), .dout(n16627));
  jand g16332(.dina(n16627), .dinb(asqrt[8] ), .dout(n16628));
  jxor g16333(.dina(n16628), .dinb(n16048), .dout(n16629));
  jnot g16334(.din(n16629), .dout(n16630));
  jor  g16335(.dina(n16625), .dinb(asqrt[19] ), .dout(n16631));
  jand g16336(.dina(n16631), .dinb(n16630), .dout(n16632));
  jor  g16337(.dina(n16632), .dinb(n16626), .dout(n16633));
  jand g16338(.dina(n16633), .dinb(asqrt[20] ), .dout(n16634));
  jnot g16339(.din(n16053), .dout(n16635));
  jand g16340(.dina(n16635), .dinb(n16051), .dout(n16636));
  jand g16341(.dina(n16636), .dinb(asqrt[8] ), .dout(n16637));
  jxor g16342(.dina(n16637), .dinb(n16061), .dout(n16638));
  jnot g16343(.din(n16638), .dout(n16639));
  jor  g16344(.dina(n16626), .dinb(asqrt[20] ), .dout(n16640));
  jor  g16345(.dina(n16640), .dinb(n16632), .dout(n16641));
  jand g16346(.dina(n16641), .dinb(n16639), .dout(n16642));
  jor  g16347(.dina(n16642), .dinb(n16634), .dout(n16643));
  jand g16348(.dina(n16643), .dinb(asqrt[21] ), .dout(n16644));
  jor  g16349(.dina(n16643), .dinb(asqrt[21] ), .dout(n16645));
  jnot g16350(.din(n16067), .dout(n16646));
  jnot g16351(.din(n16068), .dout(n16647));
  jand g16352(.dina(asqrt[8] ), .dinb(n16064), .dout(n16648));
  jand g16353(.dina(n16648), .dinb(n16647), .dout(n16649));
  jor  g16354(.dina(n16649), .dinb(n16646), .dout(n16650));
  jnot g16355(.din(n16069), .dout(n16651));
  jand g16356(.dina(n16648), .dinb(n16651), .dout(n16652));
  jnot g16357(.din(n16652), .dout(n16653));
  jand g16358(.dina(n16653), .dinb(n16650), .dout(n16654));
  jand g16359(.dina(n16654), .dinb(n16645), .dout(n16655));
  jor  g16360(.dina(n16655), .dinb(n16644), .dout(n16656));
  jand g16361(.dina(n16656), .dinb(asqrt[22] ), .dout(n16657));
  jor  g16362(.dina(n16644), .dinb(asqrt[22] ), .dout(n16658));
  jor  g16363(.dina(n16658), .dinb(n16655), .dout(n16659));
  jnot g16364(.din(n16075), .dout(n16660));
  jnot g16365(.din(n16077), .dout(n16661));
  jand g16366(.dina(asqrt[8] ), .dinb(n16071), .dout(n16662));
  jand g16367(.dina(n16662), .dinb(n16661), .dout(n16663));
  jor  g16368(.dina(n16663), .dinb(n16660), .dout(n16664));
  jnot g16369(.din(n16078), .dout(n16665));
  jand g16370(.dina(n16662), .dinb(n16665), .dout(n16666));
  jnot g16371(.din(n16666), .dout(n16667));
  jand g16372(.dina(n16667), .dinb(n16664), .dout(n16668));
  jand g16373(.dina(n16668), .dinb(n16659), .dout(n16669));
  jor  g16374(.dina(n16669), .dinb(n16657), .dout(n16670));
  jand g16375(.dina(n16670), .dinb(asqrt[23] ), .dout(n16671));
  jxor g16376(.dina(n16079), .dinb(n9769), .dout(n16672));
  jand g16377(.dina(n16672), .dinb(asqrt[8] ), .dout(n16673));
  jxor g16378(.dina(n16673), .dinb(n16089), .dout(n16674));
  jnot g16379(.din(n16674), .dout(n16675));
  jor  g16380(.dina(n16670), .dinb(asqrt[23] ), .dout(n16676));
  jand g16381(.dina(n16676), .dinb(n16675), .dout(n16677));
  jor  g16382(.dina(n16677), .dinb(n16671), .dout(n16678));
  jand g16383(.dina(n16678), .dinb(asqrt[24] ), .dout(n16679));
  jnot g16384(.din(n16094), .dout(n16680));
  jand g16385(.dina(n16680), .dinb(n16092), .dout(n16681));
  jand g16386(.dina(n16681), .dinb(asqrt[8] ), .dout(n16682));
  jxor g16387(.dina(n16682), .dinb(n16102), .dout(n16683));
  jnot g16388(.din(n16683), .dout(n16684));
  jor  g16389(.dina(n16671), .dinb(asqrt[24] ), .dout(n16685));
  jor  g16390(.dina(n16685), .dinb(n16677), .dout(n16686));
  jand g16391(.dina(n16686), .dinb(n16684), .dout(n16687));
  jor  g16392(.dina(n16687), .dinb(n16679), .dout(n16688));
  jand g16393(.dina(n16688), .dinb(asqrt[25] ), .dout(n16689));
  jor  g16394(.dina(n16688), .dinb(asqrt[25] ), .dout(n16690));
  jnot g16395(.din(n16108), .dout(n16691));
  jnot g16396(.din(n16109), .dout(n16692));
  jand g16397(.dina(asqrt[8] ), .dinb(n16105), .dout(n16693));
  jand g16398(.dina(n16693), .dinb(n16692), .dout(n16694));
  jor  g16399(.dina(n16694), .dinb(n16691), .dout(n16695));
  jnot g16400(.din(n16110), .dout(n16696));
  jand g16401(.dina(n16693), .dinb(n16696), .dout(n16697));
  jnot g16402(.din(n16697), .dout(n16698));
  jand g16403(.dina(n16698), .dinb(n16695), .dout(n16699));
  jand g16404(.dina(n16699), .dinb(n16690), .dout(n16700));
  jor  g16405(.dina(n16700), .dinb(n16689), .dout(n16701));
  jand g16406(.dina(n16701), .dinb(asqrt[26] ), .dout(n16702));
  jor  g16407(.dina(n16689), .dinb(asqrt[26] ), .dout(n16703));
  jor  g16408(.dina(n16703), .dinb(n16700), .dout(n16704));
  jnot g16409(.din(n16116), .dout(n16705));
  jnot g16410(.din(n16118), .dout(n16706));
  jand g16411(.dina(asqrt[8] ), .dinb(n16112), .dout(n16707));
  jand g16412(.dina(n16707), .dinb(n16706), .dout(n16708));
  jor  g16413(.dina(n16708), .dinb(n16705), .dout(n16709));
  jnot g16414(.din(n16119), .dout(n16710));
  jand g16415(.dina(n16707), .dinb(n16710), .dout(n16711));
  jnot g16416(.din(n16711), .dout(n16712));
  jand g16417(.dina(n16712), .dinb(n16709), .dout(n16713));
  jand g16418(.dina(n16713), .dinb(n16704), .dout(n16714));
  jor  g16419(.dina(n16714), .dinb(n16702), .dout(n16715));
  jand g16420(.dina(n16715), .dinb(asqrt[27] ), .dout(n16716));
  jxor g16421(.dina(n16120), .dinb(n8053), .dout(n16717));
  jand g16422(.dina(n16717), .dinb(asqrt[8] ), .dout(n16718));
  jxor g16423(.dina(n16718), .dinb(n16130), .dout(n16719));
  jnot g16424(.din(n16719), .dout(n16720));
  jor  g16425(.dina(n16715), .dinb(asqrt[27] ), .dout(n16721));
  jand g16426(.dina(n16721), .dinb(n16720), .dout(n16722));
  jor  g16427(.dina(n16722), .dinb(n16716), .dout(n16723));
  jand g16428(.dina(n16723), .dinb(asqrt[28] ), .dout(n16724));
  jnot g16429(.din(n16135), .dout(n16725));
  jand g16430(.dina(n16725), .dinb(n16133), .dout(n16726));
  jand g16431(.dina(n16726), .dinb(asqrt[8] ), .dout(n16727));
  jxor g16432(.dina(n16727), .dinb(n16143), .dout(n16728));
  jnot g16433(.din(n16728), .dout(n16729));
  jor  g16434(.dina(n16716), .dinb(asqrt[28] ), .dout(n16730));
  jor  g16435(.dina(n16730), .dinb(n16722), .dout(n16731));
  jand g16436(.dina(n16731), .dinb(n16729), .dout(n16732));
  jor  g16437(.dina(n16732), .dinb(n16724), .dout(n16733));
  jand g16438(.dina(n16733), .dinb(asqrt[29] ), .dout(n16734));
  jor  g16439(.dina(n16733), .dinb(asqrt[29] ), .dout(n16735));
  jnot g16440(.din(n16149), .dout(n16736));
  jnot g16441(.din(n16150), .dout(n16737));
  jand g16442(.dina(asqrt[8] ), .dinb(n16146), .dout(n16738));
  jand g16443(.dina(n16738), .dinb(n16737), .dout(n16739));
  jor  g16444(.dina(n16739), .dinb(n16736), .dout(n16740));
  jnot g16445(.din(n16151), .dout(n16741));
  jand g16446(.dina(n16738), .dinb(n16741), .dout(n16742));
  jnot g16447(.din(n16742), .dout(n16743));
  jand g16448(.dina(n16743), .dinb(n16740), .dout(n16744));
  jand g16449(.dina(n16744), .dinb(n16735), .dout(n16745));
  jor  g16450(.dina(n16745), .dinb(n16734), .dout(n16746));
  jand g16451(.dina(n16746), .dinb(asqrt[30] ), .dout(n16747));
  jor  g16452(.dina(n16734), .dinb(asqrt[30] ), .dout(n16748));
  jor  g16453(.dina(n16748), .dinb(n16745), .dout(n16749));
  jnot g16454(.din(n16157), .dout(n16750));
  jnot g16455(.din(n16159), .dout(n16751));
  jand g16456(.dina(asqrt[8] ), .dinb(n16153), .dout(n16752));
  jand g16457(.dina(n16752), .dinb(n16751), .dout(n16753));
  jor  g16458(.dina(n16753), .dinb(n16750), .dout(n16754));
  jnot g16459(.din(n16160), .dout(n16755));
  jand g16460(.dina(n16752), .dinb(n16755), .dout(n16756));
  jnot g16461(.din(n16756), .dout(n16757));
  jand g16462(.dina(n16757), .dinb(n16754), .dout(n16758));
  jand g16463(.dina(n16758), .dinb(n16749), .dout(n16759));
  jor  g16464(.dina(n16759), .dinb(n16747), .dout(n16760));
  jand g16465(.dina(n16760), .dinb(asqrt[31] ), .dout(n16761));
  jxor g16466(.dina(n16161), .dinb(n6500), .dout(n16762));
  jand g16467(.dina(n16762), .dinb(asqrt[8] ), .dout(n16763));
  jxor g16468(.dina(n16763), .dinb(n16171), .dout(n16764));
  jnot g16469(.din(n16764), .dout(n16765));
  jor  g16470(.dina(n16760), .dinb(asqrt[31] ), .dout(n16766));
  jand g16471(.dina(n16766), .dinb(n16765), .dout(n16767));
  jor  g16472(.dina(n16767), .dinb(n16761), .dout(n16768));
  jand g16473(.dina(n16768), .dinb(asqrt[32] ), .dout(n16769));
  jnot g16474(.din(n16176), .dout(n16770));
  jand g16475(.dina(n16770), .dinb(n16174), .dout(n16771));
  jand g16476(.dina(n16771), .dinb(asqrt[8] ), .dout(n16772));
  jxor g16477(.dina(n16772), .dinb(n16184), .dout(n16773));
  jnot g16478(.din(n16773), .dout(n16774));
  jor  g16479(.dina(n16761), .dinb(asqrt[32] ), .dout(n16775));
  jor  g16480(.dina(n16775), .dinb(n16767), .dout(n16776));
  jand g16481(.dina(n16776), .dinb(n16774), .dout(n16777));
  jor  g16482(.dina(n16777), .dinb(n16769), .dout(n16778));
  jand g16483(.dina(n16778), .dinb(asqrt[33] ), .dout(n16779));
  jor  g16484(.dina(n16778), .dinb(asqrt[33] ), .dout(n16780));
  jnot g16485(.din(n16190), .dout(n16781));
  jnot g16486(.din(n16191), .dout(n16782));
  jand g16487(.dina(asqrt[8] ), .dinb(n16187), .dout(n16783));
  jand g16488(.dina(n16783), .dinb(n16782), .dout(n16784));
  jor  g16489(.dina(n16784), .dinb(n16781), .dout(n16785));
  jnot g16490(.din(n16192), .dout(n16786));
  jand g16491(.dina(n16783), .dinb(n16786), .dout(n16787));
  jnot g16492(.din(n16787), .dout(n16788));
  jand g16493(.dina(n16788), .dinb(n16785), .dout(n16789));
  jand g16494(.dina(n16789), .dinb(n16780), .dout(n16790));
  jor  g16495(.dina(n16790), .dinb(n16779), .dout(n16791));
  jand g16496(.dina(n16791), .dinb(asqrt[34] ), .dout(n16792));
  jor  g16497(.dina(n16779), .dinb(asqrt[34] ), .dout(n16793));
  jor  g16498(.dina(n16793), .dinb(n16790), .dout(n16794));
  jnot g16499(.din(n16198), .dout(n16795));
  jnot g16500(.din(n16200), .dout(n16796));
  jand g16501(.dina(asqrt[8] ), .dinb(n16194), .dout(n16797));
  jand g16502(.dina(n16797), .dinb(n16796), .dout(n16798));
  jor  g16503(.dina(n16798), .dinb(n16795), .dout(n16799));
  jnot g16504(.din(n16201), .dout(n16800));
  jand g16505(.dina(n16797), .dinb(n16800), .dout(n16801));
  jnot g16506(.din(n16801), .dout(n16802));
  jand g16507(.dina(n16802), .dinb(n16799), .dout(n16803));
  jand g16508(.dina(n16803), .dinb(n16794), .dout(n16804));
  jor  g16509(.dina(n16804), .dinb(n16792), .dout(n16805));
  jand g16510(.dina(n16805), .dinb(asqrt[35] ), .dout(n16806));
  jxor g16511(.dina(n16202), .dinb(n5116), .dout(n16807));
  jand g16512(.dina(n16807), .dinb(asqrt[8] ), .dout(n16808));
  jxor g16513(.dina(n16808), .dinb(n16212), .dout(n16809));
  jnot g16514(.din(n16809), .dout(n16810));
  jor  g16515(.dina(n16805), .dinb(asqrt[35] ), .dout(n16811));
  jand g16516(.dina(n16811), .dinb(n16810), .dout(n16812));
  jor  g16517(.dina(n16812), .dinb(n16806), .dout(n16813));
  jand g16518(.dina(n16813), .dinb(asqrt[36] ), .dout(n16814));
  jnot g16519(.din(n16217), .dout(n16815));
  jand g16520(.dina(n16815), .dinb(n16215), .dout(n16816));
  jand g16521(.dina(n16816), .dinb(asqrt[8] ), .dout(n16817));
  jxor g16522(.dina(n16817), .dinb(n16225), .dout(n16818));
  jnot g16523(.din(n16818), .dout(n16819));
  jor  g16524(.dina(n16806), .dinb(asqrt[36] ), .dout(n16820));
  jor  g16525(.dina(n16820), .dinb(n16812), .dout(n16821));
  jand g16526(.dina(n16821), .dinb(n16819), .dout(n16822));
  jor  g16527(.dina(n16822), .dinb(n16814), .dout(n16823));
  jand g16528(.dina(n16823), .dinb(asqrt[37] ), .dout(n16824));
  jor  g16529(.dina(n16823), .dinb(asqrt[37] ), .dout(n16825));
  jnot g16530(.din(n16231), .dout(n16826));
  jnot g16531(.din(n16232), .dout(n16827));
  jand g16532(.dina(asqrt[8] ), .dinb(n16228), .dout(n16828));
  jand g16533(.dina(n16828), .dinb(n16827), .dout(n16829));
  jor  g16534(.dina(n16829), .dinb(n16826), .dout(n16830));
  jnot g16535(.din(n16233), .dout(n16831));
  jand g16536(.dina(n16828), .dinb(n16831), .dout(n16832));
  jnot g16537(.din(n16832), .dout(n16833));
  jand g16538(.dina(n16833), .dinb(n16830), .dout(n16834));
  jand g16539(.dina(n16834), .dinb(n16825), .dout(n16835));
  jor  g16540(.dina(n16835), .dinb(n16824), .dout(n16836));
  jand g16541(.dina(n16836), .dinb(asqrt[38] ), .dout(n16837));
  jor  g16542(.dina(n16824), .dinb(asqrt[38] ), .dout(n16838));
  jor  g16543(.dina(n16838), .dinb(n16835), .dout(n16839));
  jnot g16544(.din(n16239), .dout(n16840));
  jnot g16545(.din(n16241), .dout(n16841));
  jand g16546(.dina(asqrt[8] ), .dinb(n16235), .dout(n16842));
  jand g16547(.dina(n16842), .dinb(n16841), .dout(n16843));
  jor  g16548(.dina(n16843), .dinb(n16840), .dout(n16844));
  jnot g16549(.din(n16242), .dout(n16845));
  jand g16550(.dina(n16842), .dinb(n16845), .dout(n16846));
  jnot g16551(.din(n16846), .dout(n16847));
  jand g16552(.dina(n16847), .dinb(n16844), .dout(n16848));
  jand g16553(.dina(n16848), .dinb(n16839), .dout(n16849));
  jor  g16554(.dina(n16849), .dinb(n16837), .dout(n16850));
  jand g16555(.dina(n16850), .dinb(asqrt[39] ), .dout(n16851));
  jxor g16556(.dina(n16243), .dinb(n3907), .dout(n16852));
  jand g16557(.dina(n16852), .dinb(asqrt[8] ), .dout(n16853));
  jxor g16558(.dina(n16853), .dinb(n16253), .dout(n16854));
  jnot g16559(.din(n16854), .dout(n16855));
  jor  g16560(.dina(n16850), .dinb(asqrt[39] ), .dout(n16856));
  jand g16561(.dina(n16856), .dinb(n16855), .dout(n16857));
  jor  g16562(.dina(n16857), .dinb(n16851), .dout(n16858));
  jand g16563(.dina(n16858), .dinb(asqrt[40] ), .dout(n16859));
  jnot g16564(.din(n16258), .dout(n16860));
  jand g16565(.dina(n16860), .dinb(n16256), .dout(n16861));
  jand g16566(.dina(n16861), .dinb(asqrt[8] ), .dout(n16862));
  jxor g16567(.dina(n16862), .dinb(n16266), .dout(n16863));
  jnot g16568(.din(n16863), .dout(n16864));
  jor  g16569(.dina(n16851), .dinb(asqrt[40] ), .dout(n16865));
  jor  g16570(.dina(n16865), .dinb(n16857), .dout(n16866));
  jand g16571(.dina(n16866), .dinb(n16864), .dout(n16867));
  jor  g16572(.dina(n16867), .dinb(n16859), .dout(n16868));
  jand g16573(.dina(n16868), .dinb(asqrt[41] ), .dout(n16869));
  jor  g16574(.dina(n16868), .dinb(asqrt[41] ), .dout(n16870));
  jnot g16575(.din(n16272), .dout(n16871));
  jnot g16576(.din(n16273), .dout(n16872));
  jand g16577(.dina(asqrt[8] ), .dinb(n16269), .dout(n16873));
  jand g16578(.dina(n16873), .dinb(n16872), .dout(n16874));
  jor  g16579(.dina(n16874), .dinb(n16871), .dout(n16875));
  jnot g16580(.din(n16274), .dout(n16876));
  jand g16581(.dina(n16873), .dinb(n16876), .dout(n16877));
  jnot g16582(.din(n16877), .dout(n16878));
  jand g16583(.dina(n16878), .dinb(n16875), .dout(n16879));
  jand g16584(.dina(n16879), .dinb(n16870), .dout(n16880));
  jor  g16585(.dina(n16880), .dinb(n16869), .dout(n16881));
  jand g16586(.dina(n16881), .dinb(asqrt[42] ), .dout(n16882));
  jor  g16587(.dina(n16869), .dinb(asqrt[42] ), .dout(n16883));
  jor  g16588(.dina(n16883), .dinb(n16880), .dout(n16884));
  jnot g16589(.din(n16280), .dout(n16885));
  jnot g16590(.din(n16282), .dout(n16886));
  jand g16591(.dina(asqrt[8] ), .dinb(n16276), .dout(n16887));
  jand g16592(.dina(n16887), .dinb(n16886), .dout(n16888));
  jor  g16593(.dina(n16888), .dinb(n16885), .dout(n16889));
  jnot g16594(.din(n16283), .dout(n16890));
  jand g16595(.dina(n16887), .dinb(n16890), .dout(n16891));
  jnot g16596(.din(n16891), .dout(n16892));
  jand g16597(.dina(n16892), .dinb(n16889), .dout(n16893));
  jand g16598(.dina(n16893), .dinb(n16884), .dout(n16894));
  jor  g16599(.dina(n16894), .dinb(n16882), .dout(n16895));
  jand g16600(.dina(n16895), .dinb(asqrt[43] ), .dout(n16896));
  jxor g16601(.dina(n16284), .dinb(n2870), .dout(n16897));
  jand g16602(.dina(n16897), .dinb(asqrt[8] ), .dout(n16898));
  jxor g16603(.dina(n16898), .dinb(n16294), .dout(n16899));
  jnot g16604(.din(n16899), .dout(n16900));
  jor  g16605(.dina(n16895), .dinb(asqrt[43] ), .dout(n16901));
  jand g16606(.dina(n16901), .dinb(n16900), .dout(n16902));
  jor  g16607(.dina(n16902), .dinb(n16896), .dout(n16903));
  jand g16608(.dina(n16903), .dinb(asqrt[44] ), .dout(n16904));
  jnot g16609(.din(n16299), .dout(n16905));
  jand g16610(.dina(n16905), .dinb(n16297), .dout(n16906));
  jand g16611(.dina(n16906), .dinb(asqrt[8] ), .dout(n16907));
  jxor g16612(.dina(n16907), .dinb(n16307), .dout(n16908));
  jnot g16613(.din(n16908), .dout(n16909));
  jor  g16614(.dina(n16896), .dinb(asqrt[44] ), .dout(n16910));
  jor  g16615(.dina(n16910), .dinb(n16902), .dout(n16911));
  jand g16616(.dina(n16911), .dinb(n16909), .dout(n16912));
  jor  g16617(.dina(n16912), .dinb(n16904), .dout(n16913));
  jand g16618(.dina(n16913), .dinb(asqrt[45] ), .dout(n16914));
  jor  g16619(.dina(n16913), .dinb(asqrt[45] ), .dout(n16915));
  jnot g16620(.din(n16313), .dout(n16916));
  jnot g16621(.din(n16314), .dout(n16917));
  jand g16622(.dina(asqrt[8] ), .dinb(n16310), .dout(n16918));
  jand g16623(.dina(n16918), .dinb(n16917), .dout(n16919));
  jor  g16624(.dina(n16919), .dinb(n16916), .dout(n16920));
  jnot g16625(.din(n16315), .dout(n16921));
  jand g16626(.dina(n16918), .dinb(n16921), .dout(n16922));
  jnot g16627(.din(n16922), .dout(n16923));
  jand g16628(.dina(n16923), .dinb(n16920), .dout(n16924));
  jand g16629(.dina(n16924), .dinb(n16915), .dout(n16925));
  jor  g16630(.dina(n16925), .dinb(n16914), .dout(n16926));
  jand g16631(.dina(n16926), .dinb(asqrt[46] ), .dout(n16927));
  jor  g16632(.dina(n16914), .dinb(asqrt[46] ), .dout(n16928));
  jor  g16633(.dina(n16928), .dinb(n16925), .dout(n16929));
  jnot g16634(.din(n16321), .dout(n16930));
  jnot g16635(.din(n16323), .dout(n16931));
  jand g16636(.dina(asqrt[8] ), .dinb(n16317), .dout(n16932));
  jand g16637(.dina(n16932), .dinb(n16931), .dout(n16933));
  jor  g16638(.dina(n16933), .dinb(n16930), .dout(n16934));
  jnot g16639(.din(n16324), .dout(n16935));
  jand g16640(.dina(n16932), .dinb(n16935), .dout(n16936));
  jnot g16641(.din(n16936), .dout(n16937));
  jand g16642(.dina(n16937), .dinb(n16934), .dout(n16938));
  jand g16643(.dina(n16938), .dinb(n16929), .dout(n16939));
  jor  g16644(.dina(n16939), .dinb(n16927), .dout(n16940));
  jand g16645(.dina(n16940), .dinb(asqrt[47] ), .dout(n16941));
  jxor g16646(.dina(n16325), .dinb(n2005), .dout(n16942));
  jand g16647(.dina(n16942), .dinb(asqrt[8] ), .dout(n16943));
  jxor g16648(.dina(n16943), .dinb(n16335), .dout(n16944));
  jnot g16649(.din(n16944), .dout(n16945));
  jor  g16650(.dina(n16940), .dinb(asqrt[47] ), .dout(n16946));
  jand g16651(.dina(n16946), .dinb(n16945), .dout(n16947));
  jor  g16652(.dina(n16947), .dinb(n16941), .dout(n16948));
  jand g16653(.dina(n16948), .dinb(asqrt[48] ), .dout(n16949));
  jnot g16654(.din(n16340), .dout(n16950));
  jand g16655(.dina(n16950), .dinb(n16338), .dout(n16951));
  jand g16656(.dina(n16951), .dinb(asqrt[8] ), .dout(n16952));
  jxor g16657(.dina(n16952), .dinb(n16348), .dout(n16953));
  jnot g16658(.din(n16953), .dout(n16954));
  jor  g16659(.dina(n16941), .dinb(asqrt[48] ), .dout(n16955));
  jor  g16660(.dina(n16955), .dinb(n16947), .dout(n16956));
  jand g16661(.dina(n16956), .dinb(n16954), .dout(n16957));
  jor  g16662(.dina(n16957), .dinb(n16949), .dout(n16958));
  jand g16663(.dina(n16958), .dinb(asqrt[49] ), .dout(n16959));
  jor  g16664(.dina(n16958), .dinb(asqrt[49] ), .dout(n16960));
  jnot g16665(.din(n16354), .dout(n16961));
  jnot g16666(.din(n16355), .dout(n16962));
  jand g16667(.dina(asqrt[8] ), .dinb(n16351), .dout(n16963));
  jand g16668(.dina(n16963), .dinb(n16962), .dout(n16964));
  jor  g16669(.dina(n16964), .dinb(n16961), .dout(n16965));
  jnot g16670(.din(n16356), .dout(n16966));
  jand g16671(.dina(n16963), .dinb(n16966), .dout(n16967));
  jnot g16672(.din(n16967), .dout(n16968));
  jand g16673(.dina(n16968), .dinb(n16965), .dout(n16969));
  jand g16674(.dina(n16969), .dinb(n16960), .dout(n16970));
  jor  g16675(.dina(n16970), .dinb(n16959), .dout(n16971));
  jand g16676(.dina(n16971), .dinb(asqrt[50] ), .dout(n16972));
  jor  g16677(.dina(n16959), .dinb(asqrt[50] ), .dout(n16973));
  jor  g16678(.dina(n16973), .dinb(n16970), .dout(n16974));
  jnot g16679(.din(n16362), .dout(n16975));
  jnot g16680(.din(n16364), .dout(n16976));
  jand g16681(.dina(asqrt[8] ), .dinb(n16358), .dout(n16977));
  jand g16682(.dina(n16977), .dinb(n16976), .dout(n16978));
  jor  g16683(.dina(n16978), .dinb(n16975), .dout(n16979));
  jnot g16684(.din(n16365), .dout(n16980));
  jand g16685(.dina(n16977), .dinb(n16980), .dout(n16981));
  jnot g16686(.din(n16981), .dout(n16982));
  jand g16687(.dina(n16982), .dinb(n16979), .dout(n16983));
  jand g16688(.dina(n16983), .dinb(n16974), .dout(n16984));
  jor  g16689(.dina(n16984), .dinb(n16972), .dout(n16985));
  jand g16690(.dina(n16985), .dinb(asqrt[51] ), .dout(n16986));
  jxor g16691(.dina(n16366), .dinb(n1312), .dout(n16987));
  jand g16692(.dina(n16987), .dinb(asqrt[8] ), .dout(n16988));
  jxor g16693(.dina(n16988), .dinb(n16376), .dout(n16989));
  jnot g16694(.din(n16989), .dout(n16990));
  jor  g16695(.dina(n16985), .dinb(asqrt[51] ), .dout(n16991));
  jand g16696(.dina(n16991), .dinb(n16990), .dout(n16992));
  jor  g16697(.dina(n16992), .dinb(n16986), .dout(n16993));
  jand g16698(.dina(n16993), .dinb(asqrt[52] ), .dout(n16994));
  jnot g16699(.din(n16381), .dout(n16995));
  jand g16700(.dina(n16995), .dinb(n16379), .dout(n16996));
  jand g16701(.dina(n16996), .dinb(asqrt[8] ), .dout(n16997));
  jxor g16702(.dina(n16997), .dinb(n16389), .dout(n16998));
  jnot g16703(.din(n16998), .dout(n16999));
  jor  g16704(.dina(n16986), .dinb(asqrt[52] ), .dout(n17000));
  jor  g16705(.dina(n17000), .dinb(n16992), .dout(n17001));
  jand g16706(.dina(n17001), .dinb(n16999), .dout(n17002));
  jor  g16707(.dina(n17002), .dinb(n16994), .dout(n17003));
  jand g16708(.dina(n17003), .dinb(asqrt[53] ), .dout(n17004));
  jor  g16709(.dina(n17003), .dinb(asqrt[53] ), .dout(n17005));
  jnot g16710(.din(n16395), .dout(n17006));
  jnot g16711(.din(n16396), .dout(n17007));
  jand g16712(.dina(asqrt[8] ), .dinb(n16392), .dout(n17008));
  jand g16713(.dina(n17008), .dinb(n17007), .dout(n17009));
  jor  g16714(.dina(n17009), .dinb(n17006), .dout(n17010));
  jnot g16715(.din(n16397), .dout(n17011));
  jand g16716(.dina(n17008), .dinb(n17011), .dout(n17012));
  jnot g16717(.din(n17012), .dout(n17013));
  jand g16718(.dina(n17013), .dinb(n17010), .dout(n17014));
  jand g16719(.dina(n17014), .dinb(n17005), .dout(n17015));
  jor  g16720(.dina(n17015), .dinb(n17004), .dout(n17016));
  jand g16721(.dina(n17016), .dinb(asqrt[54] ), .dout(n17017));
  jnot g16722(.din(n16401), .dout(n17018));
  jand g16723(.dina(n17018), .dinb(n16399), .dout(n17019));
  jand g16724(.dina(n17019), .dinb(asqrt[8] ), .dout(n17020));
  jxor g16725(.dina(n17020), .dinb(n16409), .dout(n17021));
  jnot g16726(.din(n17021), .dout(n17022));
  jor  g16727(.dina(n17004), .dinb(asqrt[54] ), .dout(n17023));
  jor  g16728(.dina(n17023), .dinb(n17015), .dout(n17024));
  jand g16729(.dina(n17024), .dinb(n17022), .dout(n17025));
  jor  g16730(.dina(n17025), .dinb(n17017), .dout(n17026));
  jand g16731(.dina(n17026), .dinb(asqrt[55] ), .dout(n17027));
  jor  g16732(.dina(n17026), .dinb(asqrt[55] ), .dout(n17028));
  jand g16733(.dina(n17028), .dinb(n16521), .dout(n17029));
  jor  g16734(.dina(n17029), .dinb(n17027), .dout(n17030));
  jand g16735(.dina(n17030), .dinb(asqrt[56] ), .dout(n17031));
  jor  g16736(.dina(n17027), .dinb(asqrt[56] ), .dout(n17032));
  jor  g16737(.dina(n17032), .dinb(n17029), .dout(n17033));
  jnot g16738(.din(n16420), .dout(n17034));
  jnot g16739(.din(n16422), .dout(n17035));
  jand g16740(.dina(asqrt[8] ), .dinb(n16416), .dout(n17036));
  jand g16741(.dina(n17036), .dinb(n17035), .dout(n17037));
  jor  g16742(.dina(n17037), .dinb(n17034), .dout(n17038));
  jnot g16743(.din(n16423), .dout(n17039));
  jand g16744(.dina(n17036), .dinb(n17039), .dout(n17040));
  jnot g16745(.din(n17040), .dout(n17041));
  jand g16746(.dina(n17041), .dinb(n17038), .dout(n17042));
  jand g16747(.dina(n17042), .dinb(n17033), .dout(n17043));
  jor  g16748(.dina(n17043), .dinb(n17031), .dout(n17044));
  jand g16749(.dina(n17044), .dinb(asqrt[57] ), .dout(n17045));
  jor  g16750(.dina(n17044), .dinb(asqrt[57] ), .dout(n17046));
  jnot g16751(.din(n16428), .dout(n17047));
  jnot g16752(.din(n16429), .dout(n17048));
  jand g16753(.dina(asqrt[8] ), .dinb(n16425), .dout(n17049));
  jand g16754(.dina(n17049), .dinb(n17048), .dout(n17050));
  jor  g16755(.dina(n17050), .dinb(n17047), .dout(n17051));
  jnot g16756(.din(n16430), .dout(n17052));
  jand g16757(.dina(n17049), .dinb(n17052), .dout(n17053));
  jnot g16758(.din(n17053), .dout(n17054));
  jand g16759(.dina(n17054), .dinb(n17051), .dout(n17055));
  jand g16760(.dina(n17055), .dinb(n17046), .dout(n17056));
  jor  g16761(.dina(n17056), .dinb(n17045), .dout(n17057));
  jand g16762(.dina(n17057), .dinb(asqrt[58] ), .dout(n17058));
  jor  g16763(.dina(n17045), .dinb(asqrt[58] ), .dout(n17059));
  jor  g16764(.dina(n17059), .dinb(n17056), .dout(n17060));
  jnot g16765(.din(n16436), .dout(n17061));
  jnot g16766(.din(n16438), .dout(n17062));
  jand g16767(.dina(asqrt[8] ), .dinb(n16432), .dout(n17063));
  jand g16768(.dina(n17063), .dinb(n17062), .dout(n17064));
  jor  g16769(.dina(n17064), .dinb(n17061), .dout(n17065));
  jnot g16770(.din(n16439), .dout(n17066));
  jand g16771(.dina(n17063), .dinb(n17066), .dout(n17067));
  jnot g16772(.din(n17067), .dout(n17068));
  jand g16773(.dina(n17068), .dinb(n17065), .dout(n17069));
  jand g16774(.dina(n17069), .dinb(n17060), .dout(n17070));
  jor  g16775(.dina(n17070), .dinb(n17058), .dout(n17071));
  jand g16776(.dina(n17071), .dinb(asqrt[59] ), .dout(n17072));
  jxor g16777(.dina(n16440), .dinb(n425), .dout(n17073));
  jand g16778(.dina(n17073), .dinb(asqrt[8] ), .dout(n17074));
  jxor g16779(.dina(n17074), .dinb(n16450), .dout(n17075));
  jnot g16780(.din(n17075), .dout(n17076));
  jor  g16781(.dina(n17071), .dinb(asqrt[59] ), .dout(n17077));
  jand g16782(.dina(n17077), .dinb(n17076), .dout(n17078));
  jor  g16783(.dina(n17078), .dinb(n17072), .dout(n17079));
  jand g16784(.dina(n17079), .dinb(asqrt[60] ), .dout(n17080));
  jnot g16785(.din(n16455), .dout(n17081));
  jand g16786(.dina(n17081), .dinb(n16453), .dout(n17082));
  jand g16787(.dina(n17082), .dinb(asqrt[8] ), .dout(n17083));
  jxor g16788(.dina(n17083), .dinb(n16463), .dout(n17084));
  jnot g16789(.din(n17084), .dout(n17085));
  jor  g16790(.dina(n17072), .dinb(asqrt[60] ), .dout(n17086));
  jor  g16791(.dina(n17086), .dinb(n17078), .dout(n17087));
  jand g16792(.dina(n17087), .dinb(n17085), .dout(n17088));
  jor  g16793(.dina(n17088), .dinb(n17080), .dout(n17089));
  jand g16794(.dina(n17089), .dinb(asqrt[61] ), .dout(n17090));
  jor  g16795(.dina(n17089), .dinb(asqrt[61] ), .dout(n17091));
  jnot g16796(.din(n16469), .dout(n17092));
  jnot g16797(.din(n16470), .dout(n17093));
  jand g16798(.dina(asqrt[8] ), .dinb(n16466), .dout(n17094));
  jand g16799(.dina(n17094), .dinb(n17093), .dout(n17095));
  jor  g16800(.dina(n17095), .dinb(n17092), .dout(n17096));
  jnot g16801(.din(n16471), .dout(n17097));
  jand g16802(.dina(n17094), .dinb(n17097), .dout(n17098));
  jnot g16803(.din(n17098), .dout(n17099));
  jand g16804(.dina(n17099), .dinb(n17096), .dout(n17100));
  jand g16805(.dina(n17100), .dinb(n17091), .dout(n17101));
  jor  g16806(.dina(n17101), .dinb(n17090), .dout(n17102));
  jand g16807(.dina(n17102), .dinb(asqrt[62] ), .dout(n17103));
  jor  g16808(.dina(n17090), .dinb(asqrt[62] ), .dout(n17104));
  jor  g16809(.dina(n17104), .dinb(n17101), .dout(n17105));
  jnot g16810(.din(n16477), .dout(n17106));
  jnot g16811(.din(n16479), .dout(n17107));
  jand g16812(.dina(asqrt[8] ), .dinb(n16473), .dout(n17108));
  jand g16813(.dina(n17108), .dinb(n17107), .dout(n17109));
  jor  g16814(.dina(n17109), .dinb(n17106), .dout(n17110));
  jnot g16815(.din(n16480), .dout(n17111));
  jand g16816(.dina(n17108), .dinb(n17111), .dout(n17112));
  jnot g16817(.din(n17112), .dout(n17113));
  jand g16818(.dina(n17113), .dinb(n17110), .dout(n17114));
  jand g16819(.dina(n17114), .dinb(n17105), .dout(n17115));
  jor  g16820(.dina(n17115), .dinb(n17103), .dout(n17116));
  jxor g16821(.dina(n16481), .dinb(n199), .dout(n17117));
  jand g16822(.dina(n17117), .dinb(asqrt[8] ), .dout(n17118));
  jxor g16823(.dina(n17118), .dinb(n16491), .dout(n17119));
  jnot g16824(.din(n16493), .dout(n17120));
  jand g16825(.dina(asqrt[8] ), .dinb(n16500), .dout(n17121));
  jand g16826(.dina(n17121), .dinb(n17120), .dout(n17122));
  jor  g16827(.dina(n17122), .dinb(n16508), .dout(n17123));
  jor  g16828(.dina(n17123), .dinb(n17119), .dout(n17124));
  jnot g16829(.din(n17124), .dout(n17125));
  jand g16830(.dina(n17125), .dinb(n17116), .dout(n17126));
  jor  g16831(.dina(n17126), .dinb(asqrt[63] ), .dout(n17127));
  jnot g16832(.din(n17119), .dout(n17128));
  jor  g16833(.dina(n17128), .dinb(n17116), .dout(n17129));
  jor  g16834(.dina(n17121), .dinb(n17120), .dout(n17130));
  jand g16835(.dina(n16500), .dinb(n17120), .dout(n17131));
  jor  g16836(.dina(n17131), .dinb(n194), .dout(n17132));
  jnot g16837(.din(n17132), .dout(n17133));
  jand g16838(.dina(n17133), .dinb(n17130), .dout(n17134));
  jnot g16839(.din(asqrt[8] ), .dout(n17135));
  jnot g16840(.din(n17134), .dout(n17138));
  jand g16841(.dina(n17138), .dinb(n17129), .dout(n17139));
  jand g16842(.dina(n17139), .dinb(n17127), .dout(n17140));
  jxor g16843(.dina(n17026), .dinb(n595), .dout(n17141));
  jor  g16844(.dina(n17141), .dinb(n17140), .dout(n17142));
  jxor g16845(.dina(n17142), .dinb(n16521), .dout(n17143));
  jor  g16846(.dina(n17140), .dinb(n16523), .dout(n17144));
  jnot g16847(.din(a[12] ), .dout(n17145));
  jnot g16848(.din(a[13] ), .dout(n17146));
  jand g16849(.dina(n16523), .dinb(n17146), .dout(n17147));
  jand g16850(.dina(n17147), .dinb(n17145), .dout(n17148));
  jnot g16851(.din(n17148), .dout(n17149));
  jand g16852(.dina(n17149), .dinb(n17144), .dout(n17150));
  jor  g16853(.dina(n17150), .dinb(n17135), .dout(n17151));
  jor  g16854(.dina(n17140), .dinb(a[14] ), .dout(n17152));
  jxor g16855(.dina(n17152), .dinb(n16524), .dout(n17153));
  jand g16856(.dina(n17150), .dinb(n17135), .dout(n17154));
  jor  g16857(.dina(n17154), .dinb(n17153), .dout(n17155));
  jand g16858(.dina(n17155), .dinb(n17151), .dout(n17156));
  jor  g16859(.dina(n17156), .dinb(n15955), .dout(n17157));
  jand g16860(.dina(n17151), .dinb(n15955), .dout(n17158));
  jand g16861(.dina(n17158), .dinb(n17155), .dout(n17159));
  jor  g16862(.dina(n17152), .dinb(a[15] ), .dout(n17160));
  jnot g16863(.din(n17127), .dout(n17161));
  jnot g16864(.din(n17129), .dout(n17162));
  jor  g16865(.dina(n17134), .dinb(n17135), .dout(n17163));
  jor  g16866(.dina(n17163), .dinb(n17162), .dout(n17164));
  jor  g16867(.dina(n17164), .dinb(n17161), .dout(n17165));
  jand g16868(.dina(n17165), .dinb(n17160), .dout(n17166));
  jxor g16869(.dina(n17166), .dinb(n15961), .dout(n17167));
  jor  g16870(.dina(n17167), .dinb(n17159), .dout(n17168));
  jand g16871(.dina(n17168), .dinb(n17157), .dout(n17169));
  jor  g16872(.dina(n17169), .dinb(n15950), .dout(n17170));
  jand g16873(.dina(n17169), .dinb(n15950), .dout(n17171));
  jxor g16874(.dina(n16527), .dinb(n15955), .dout(n17172));
  jor  g16875(.dina(n17172), .dinb(n17140), .dout(n17173));
  jxor g16876(.dina(n17173), .dinb(n16530), .dout(n17174));
  jor  g16877(.dina(n17174), .dinb(n17171), .dout(n17175));
  jand g16878(.dina(n17175), .dinb(n17170), .dout(n17176));
  jor  g16879(.dina(n17176), .dinb(n14821), .dout(n17177));
  jnot g16880(.din(n16536), .dout(n17178));
  jor  g16881(.dina(n17178), .dinb(n16534), .dout(n17179));
  jor  g16882(.dina(n17179), .dinb(n17140), .dout(n17180));
  jxor g16883(.dina(n17180), .dinb(n16545), .dout(n17181));
  jand g16884(.dina(n17170), .dinb(n14821), .dout(n17182));
  jand g16885(.dina(n17182), .dinb(n17175), .dout(n17183));
  jor  g16886(.dina(n17183), .dinb(n17181), .dout(n17184));
  jand g16887(.dina(n17184), .dinb(n17177), .dout(n17185));
  jor  g16888(.dina(n17185), .dinb(n14816), .dout(n17186));
  jand g16889(.dina(n17185), .dinb(n14816), .dout(n17187));
  jxor g16890(.dina(n16547), .dinb(n14821), .dout(n17188));
  jor  g16891(.dina(n17188), .dinb(n17140), .dout(n17189));
  jxor g16892(.dina(n17189), .dinb(n16552), .dout(n17190));
  jnot g16893(.din(n17190), .dout(n17191));
  jor  g16894(.dina(n17191), .dinb(n17187), .dout(n17192));
  jand g16895(.dina(n17192), .dinb(n17186), .dout(n17193));
  jor  g16896(.dina(n17193), .dinb(n13723), .dout(n17194));
  jand g16897(.dina(n17186), .dinb(n13723), .dout(n17195));
  jand g16898(.dina(n17195), .dinb(n17192), .dout(n17196));
  jnot g16899(.din(n16556), .dout(n17197));
  jnot g16900(.din(n17140), .dout(asqrt[7] ));
  jand g16901(.dina(asqrt[7] ), .dinb(n17197), .dout(n17199));
  jand g16902(.dina(n17199), .dinb(n16563), .dout(n17200));
  jor  g16903(.dina(n17200), .dinb(n16561), .dout(n17201));
  jand g16904(.dina(n17199), .dinb(n16564), .dout(n17202));
  jnot g16905(.din(n17202), .dout(n17203));
  jand g16906(.dina(n17203), .dinb(n17201), .dout(n17204));
  jnot g16907(.din(n17204), .dout(n17205));
  jor  g16908(.dina(n17205), .dinb(n17196), .dout(n17206));
  jand g16909(.dina(n17206), .dinb(n17194), .dout(n17207));
  jor  g16910(.dina(n17207), .dinb(n13718), .dout(n17208));
  jand g16911(.dina(n17207), .dinb(n13718), .dout(n17209));
  jnot g16912(.din(n16571), .dout(n17210));
  jxor g16913(.dina(n16565), .dinb(n13723), .dout(n17211));
  jor  g16914(.dina(n17211), .dinb(n17140), .dout(n17212));
  jxor g16915(.dina(n17212), .dinb(n17210), .dout(n17213));
  jnot g16916(.din(n17213), .dout(n17214));
  jor  g16917(.dina(n17214), .dinb(n17209), .dout(n17215));
  jand g16918(.dina(n17215), .dinb(n17208), .dout(n17216));
  jor  g16919(.dina(n17216), .dinb(n12675), .dout(n17217));
  jnot g16920(.din(n16576), .dout(n17218));
  jor  g16921(.dina(n17218), .dinb(n16574), .dout(n17219));
  jor  g16922(.dina(n17219), .dinb(n17140), .dout(n17220));
  jxor g16923(.dina(n17220), .dinb(n16585), .dout(n17221));
  jand g16924(.dina(n17208), .dinb(n12675), .dout(n17222));
  jand g16925(.dina(n17222), .dinb(n17215), .dout(n17223));
  jor  g16926(.dina(n17223), .dinb(n17221), .dout(n17224));
  jand g16927(.dina(n17224), .dinb(n17217), .dout(n17225));
  jor  g16928(.dina(n17225), .dinb(n12670), .dout(n17226));
  jand g16929(.dina(n17225), .dinb(n12670), .dout(n17227));
  jnot g16930(.din(n16592), .dout(n17228));
  jxor g16931(.dina(n16587), .dinb(n12675), .dout(n17229));
  jor  g16932(.dina(n17229), .dinb(n17140), .dout(n17230));
  jxor g16933(.dina(n17230), .dinb(n17228), .dout(n17231));
  jnot g16934(.din(n17231), .dout(n17232));
  jor  g16935(.dina(n17232), .dinb(n17227), .dout(n17233));
  jand g16936(.dina(n17233), .dinb(n17226), .dout(n17234));
  jor  g16937(.dina(n17234), .dinb(n11662), .dout(n17235));
  jand g16938(.dina(n17226), .dinb(n11662), .dout(n17236));
  jand g16939(.dina(n17236), .dinb(n17233), .dout(n17237));
  jnot g16940(.din(n16595), .dout(n17238));
  jand g16941(.dina(asqrt[7] ), .dinb(n17238), .dout(n17239));
  jand g16942(.dina(n17239), .dinb(n16602), .dout(n17240));
  jor  g16943(.dina(n17240), .dinb(n16600), .dout(n17241));
  jand g16944(.dina(n17239), .dinb(n16603), .dout(n17242));
  jnot g16945(.din(n17242), .dout(n17243));
  jand g16946(.dina(n17243), .dinb(n17241), .dout(n17244));
  jnot g16947(.din(n17244), .dout(n17245));
  jor  g16948(.dina(n17245), .dinb(n17237), .dout(n17246));
  jand g16949(.dina(n17246), .dinb(n17235), .dout(n17247));
  jor  g16950(.dina(n17247), .dinb(n11657), .dout(n17248));
  jxor g16951(.dina(n16604), .dinb(n11662), .dout(n17249));
  jor  g16952(.dina(n17249), .dinb(n17140), .dout(n17250));
  jxor g16953(.dina(n17250), .dinb(n16609), .dout(n17251));
  jand g16954(.dina(n17247), .dinb(n11657), .dout(n17252));
  jor  g16955(.dina(n17252), .dinb(n17251), .dout(n17253));
  jand g16956(.dina(n17253), .dinb(n17248), .dout(n17254));
  jor  g16957(.dina(n17254), .dinb(n10701), .dout(n17255));
  jnot g16958(.din(n16614), .dout(n17256));
  jor  g16959(.dina(n17256), .dinb(n16612), .dout(n17257));
  jor  g16960(.dina(n17257), .dinb(n17140), .dout(n17258));
  jxor g16961(.dina(n17258), .dinb(n16623), .dout(n17259));
  jand g16962(.dina(n17248), .dinb(n10701), .dout(n17260));
  jand g16963(.dina(n17260), .dinb(n17253), .dout(n17261));
  jor  g16964(.dina(n17261), .dinb(n17259), .dout(n17262));
  jand g16965(.dina(n17262), .dinb(n17255), .dout(n17263));
  jor  g16966(.dina(n17263), .dinb(n10696), .dout(n17264));
  jand g16967(.dina(n17263), .dinb(n10696), .dout(n17265));
  jnot g16968(.din(n16626), .dout(n17266));
  jand g16969(.dina(asqrt[7] ), .dinb(n17266), .dout(n17267));
  jand g16970(.dina(n17267), .dinb(n16631), .dout(n17268));
  jor  g16971(.dina(n17268), .dinb(n16630), .dout(n17269));
  jand g16972(.dina(n17267), .dinb(n16632), .dout(n17270));
  jnot g16973(.din(n17270), .dout(n17271));
  jand g16974(.dina(n17271), .dinb(n17269), .dout(n17272));
  jnot g16975(.din(n17272), .dout(n17273));
  jor  g16976(.dina(n17273), .dinb(n17265), .dout(n17274));
  jand g16977(.dina(n17274), .dinb(n17264), .dout(n17275));
  jor  g16978(.dina(n17275), .dinb(n9774), .dout(n17276));
  jand g16979(.dina(n17264), .dinb(n9774), .dout(n17277));
  jand g16980(.dina(n17277), .dinb(n17274), .dout(n17278));
  jnot g16981(.din(n16634), .dout(n17279));
  jand g16982(.dina(asqrt[7] ), .dinb(n17279), .dout(n17280));
  jand g16983(.dina(n17280), .dinb(n16641), .dout(n17281));
  jor  g16984(.dina(n17281), .dinb(n16639), .dout(n17282));
  jand g16985(.dina(n17280), .dinb(n16642), .dout(n17283));
  jnot g16986(.din(n17283), .dout(n17284));
  jand g16987(.dina(n17284), .dinb(n17282), .dout(n17285));
  jnot g16988(.din(n17285), .dout(n17286));
  jor  g16989(.dina(n17286), .dinb(n17278), .dout(n17287));
  jand g16990(.dina(n17287), .dinb(n17276), .dout(n17288));
  jor  g16991(.dina(n17288), .dinb(n9769), .dout(n17289));
  jxor g16992(.dina(n16643), .dinb(n9774), .dout(n17290));
  jor  g16993(.dina(n17290), .dinb(n17140), .dout(n17291));
  jxor g16994(.dina(n17291), .dinb(n16654), .dout(n17292));
  jand g16995(.dina(n17288), .dinb(n9769), .dout(n17293));
  jor  g16996(.dina(n17293), .dinb(n17292), .dout(n17294));
  jand g16997(.dina(n17294), .dinb(n17289), .dout(n17295));
  jor  g16998(.dina(n17295), .dinb(n8898), .dout(n17296));
  jnot g16999(.din(n16659), .dout(n17297));
  jor  g17000(.dina(n17297), .dinb(n16657), .dout(n17298));
  jor  g17001(.dina(n17298), .dinb(n17140), .dout(n17299));
  jxor g17002(.dina(n17299), .dinb(n16668), .dout(n17300));
  jand g17003(.dina(n17289), .dinb(n8898), .dout(n17301));
  jand g17004(.dina(n17301), .dinb(n17294), .dout(n17302));
  jor  g17005(.dina(n17302), .dinb(n17300), .dout(n17303));
  jand g17006(.dina(n17303), .dinb(n17296), .dout(n17304));
  jor  g17007(.dina(n17304), .dinb(n8893), .dout(n17305));
  jand g17008(.dina(n17304), .dinb(n8893), .dout(n17306));
  jnot g17009(.din(n16671), .dout(n17307));
  jand g17010(.dina(asqrt[7] ), .dinb(n17307), .dout(n17308));
  jand g17011(.dina(n17308), .dinb(n16676), .dout(n17309));
  jor  g17012(.dina(n17309), .dinb(n16675), .dout(n17310));
  jand g17013(.dina(n17308), .dinb(n16677), .dout(n17311));
  jnot g17014(.din(n17311), .dout(n17312));
  jand g17015(.dina(n17312), .dinb(n17310), .dout(n17313));
  jnot g17016(.din(n17313), .dout(n17314));
  jor  g17017(.dina(n17314), .dinb(n17306), .dout(n17315));
  jand g17018(.dina(n17315), .dinb(n17305), .dout(n17316));
  jor  g17019(.dina(n17316), .dinb(n8058), .dout(n17317));
  jand g17020(.dina(n17305), .dinb(n8058), .dout(n17318));
  jand g17021(.dina(n17318), .dinb(n17315), .dout(n17319));
  jnot g17022(.din(n16679), .dout(n17320));
  jand g17023(.dina(asqrt[7] ), .dinb(n17320), .dout(n17321));
  jand g17024(.dina(n17321), .dinb(n16686), .dout(n17322));
  jor  g17025(.dina(n17322), .dinb(n16684), .dout(n17323));
  jand g17026(.dina(n17321), .dinb(n16687), .dout(n17324));
  jnot g17027(.din(n17324), .dout(n17325));
  jand g17028(.dina(n17325), .dinb(n17323), .dout(n17326));
  jnot g17029(.din(n17326), .dout(n17327));
  jor  g17030(.dina(n17327), .dinb(n17319), .dout(n17328));
  jand g17031(.dina(n17328), .dinb(n17317), .dout(n17329));
  jor  g17032(.dina(n17329), .dinb(n8053), .dout(n17330));
  jxor g17033(.dina(n16688), .dinb(n8058), .dout(n17331));
  jor  g17034(.dina(n17331), .dinb(n17140), .dout(n17332));
  jxor g17035(.dina(n17332), .dinb(n16699), .dout(n17333));
  jand g17036(.dina(n17329), .dinb(n8053), .dout(n17334));
  jor  g17037(.dina(n17334), .dinb(n17333), .dout(n17335));
  jand g17038(.dina(n17335), .dinb(n17330), .dout(n17336));
  jor  g17039(.dina(n17336), .dinb(n7265), .dout(n17337));
  jnot g17040(.din(n16704), .dout(n17338));
  jor  g17041(.dina(n17338), .dinb(n16702), .dout(n17339));
  jor  g17042(.dina(n17339), .dinb(n17140), .dout(n17340));
  jxor g17043(.dina(n17340), .dinb(n16713), .dout(n17341));
  jand g17044(.dina(n17330), .dinb(n7265), .dout(n17342));
  jand g17045(.dina(n17342), .dinb(n17335), .dout(n17343));
  jor  g17046(.dina(n17343), .dinb(n17341), .dout(n17344));
  jand g17047(.dina(n17344), .dinb(n17337), .dout(n17345));
  jor  g17048(.dina(n17345), .dinb(n7260), .dout(n17346));
  jand g17049(.dina(n17345), .dinb(n7260), .dout(n17347));
  jnot g17050(.din(n16716), .dout(n17348));
  jand g17051(.dina(asqrt[7] ), .dinb(n17348), .dout(n17349));
  jand g17052(.dina(n17349), .dinb(n16721), .dout(n17350));
  jor  g17053(.dina(n17350), .dinb(n16720), .dout(n17351));
  jand g17054(.dina(n17349), .dinb(n16722), .dout(n17352));
  jnot g17055(.din(n17352), .dout(n17353));
  jand g17056(.dina(n17353), .dinb(n17351), .dout(n17354));
  jnot g17057(.din(n17354), .dout(n17355));
  jor  g17058(.dina(n17355), .dinb(n17347), .dout(n17356));
  jand g17059(.dina(n17356), .dinb(n17346), .dout(n17357));
  jor  g17060(.dina(n17357), .dinb(n6505), .dout(n17358));
  jand g17061(.dina(n17346), .dinb(n6505), .dout(n17359));
  jand g17062(.dina(n17359), .dinb(n17356), .dout(n17360));
  jnot g17063(.din(n16724), .dout(n17361));
  jand g17064(.dina(asqrt[7] ), .dinb(n17361), .dout(n17362));
  jand g17065(.dina(n17362), .dinb(n16731), .dout(n17363));
  jor  g17066(.dina(n17363), .dinb(n16729), .dout(n17364));
  jand g17067(.dina(n17362), .dinb(n16732), .dout(n17365));
  jnot g17068(.din(n17365), .dout(n17366));
  jand g17069(.dina(n17366), .dinb(n17364), .dout(n17367));
  jnot g17070(.din(n17367), .dout(n17368));
  jor  g17071(.dina(n17368), .dinb(n17360), .dout(n17369));
  jand g17072(.dina(n17369), .dinb(n17358), .dout(n17370));
  jor  g17073(.dina(n17370), .dinb(n6500), .dout(n17371));
  jxor g17074(.dina(n16733), .dinb(n6505), .dout(n17372));
  jor  g17075(.dina(n17372), .dinb(n17140), .dout(n17373));
  jxor g17076(.dina(n17373), .dinb(n16744), .dout(n17374));
  jand g17077(.dina(n17370), .dinb(n6500), .dout(n17375));
  jor  g17078(.dina(n17375), .dinb(n17374), .dout(n17376));
  jand g17079(.dina(n17376), .dinb(n17371), .dout(n17377));
  jor  g17080(.dina(n17377), .dinb(n5793), .dout(n17378));
  jnot g17081(.din(n16749), .dout(n17379));
  jor  g17082(.dina(n17379), .dinb(n16747), .dout(n17380));
  jor  g17083(.dina(n17380), .dinb(n17140), .dout(n17381));
  jxor g17084(.dina(n17381), .dinb(n16758), .dout(n17382));
  jand g17085(.dina(n17371), .dinb(n5793), .dout(n17383));
  jand g17086(.dina(n17383), .dinb(n17376), .dout(n17384));
  jor  g17087(.dina(n17384), .dinb(n17382), .dout(n17385));
  jand g17088(.dina(n17385), .dinb(n17378), .dout(n17386));
  jor  g17089(.dina(n17386), .dinb(n5788), .dout(n17387));
  jand g17090(.dina(n17386), .dinb(n5788), .dout(n17388));
  jnot g17091(.din(n16761), .dout(n17389));
  jand g17092(.dina(asqrt[7] ), .dinb(n17389), .dout(n17390));
  jand g17093(.dina(n17390), .dinb(n16766), .dout(n17391));
  jor  g17094(.dina(n17391), .dinb(n16765), .dout(n17392));
  jand g17095(.dina(n17390), .dinb(n16767), .dout(n17393));
  jnot g17096(.din(n17393), .dout(n17394));
  jand g17097(.dina(n17394), .dinb(n17392), .dout(n17395));
  jnot g17098(.din(n17395), .dout(n17396));
  jor  g17099(.dina(n17396), .dinb(n17388), .dout(n17397));
  jand g17100(.dina(n17397), .dinb(n17387), .dout(n17398));
  jor  g17101(.dina(n17398), .dinb(n5121), .dout(n17399));
  jand g17102(.dina(n17387), .dinb(n5121), .dout(n17400));
  jand g17103(.dina(n17400), .dinb(n17397), .dout(n17401));
  jnot g17104(.din(n16769), .dout(n17402));
  jand g17105(.dina(asqrt[7] ), .dinb(n17402), .dout(n17403));
  jand g17106(.dina(n17403), .dinb(n16776), .dout(n17404));
  jor  g17107(.dina(n17404), .dinb(n16774), .dout(n17405));
  jand g17108(.dina(n17403), .dinb(n16777), .dout(n17406));
  jnot g17109(.din(n17406), .dout(n17407));
  jand g17110(.dina(n17407), .dinb(n17405), .dout(n17408));
  jnot g17111(.din(n17408), .dout(n17409));
  jor  g17112(.dina(n17409), .dinb(n17401), .dout(n17410));
  jand g17113(.dina(n17410), .dinb(n17399), .dout(n17411));
  jor  g17114(.dina(n17411), .dinb(n5116), .dout(n17412));
  jxor g17115(.dina(n16778), .dinb(n5121), .dout(n17413));
  jor  g17116(.dina(n17413), .dinb(n17140), .dout(n17414));
  jxor g17117(.dina(n17414), .dinb(n16789), .dout(n17415));
  jand g17118(.dina(n17411), .dinb(n5116), .dout(n17416));
  jor  g17119(.dina(n17416), .dinb(n17415), .dout(n17417));
  jand g17120(.dina(n17417), .dinb(n17412), .dout(n17418));
  jor  g17121(.dina(n17418), .dinb(n4499), .dout(n17419));
  jnot g17122(.din(n16794), .dout(n17420));
  jor  g17123(.dina(n17420), .dinb(n16792), .dout(n17421));
  jor  g17124(.dina(n17421), .dinb(n17140), .dout(n17422));
  jxor g17125(.dina(n17422), .dinb(n16803), .dout(n17423));
  jand g17126(.dina(n17412), .dinb(n4499), .dout(n17424));
  jand g17127(.dina(n17424), .dinb(n17417), .dout(n17425));
  jor  g17128(.dina(n17425), .dinb(n17423), .dout(n17426));
  jand g17129(.dina(n17426), .dinb(n17419), .dout(n17427));
  jor  g17130(.dina(n17427), .dinb(n4494), .dout(n17428));
  jand g17131(.dina(n17427), .dinb(n4494), .dout(n17429));
  jnot g17132(.din(n16806), .dout(n17430));
  jand g17133(.dina(asqrt[7] ), .dinb(n17430), .dout(n17431));
  jand g17134(.dina(n17431), .dinb(n16811), .dout(n17432));
  jor  g17135(.dina(n17432), .dinb(n16810), .dout(n17433));
  jand g17136(.dina(n17431), .dinb(n16812), .dout(n17434));
  jnot g17137(.din(n17434), .dout(n17435));
  jand g17138(.dina(n17435), .dinb(n17433), .dout(n17436));
  jnot g17139(.din(n17436), .dout(n17437));
  jor  g17140(.dina(n17437), .dinb(n17429), .dout(n17438));
  jand g17141(.dina(n17438), .dinb(n17428), .dout(n17439));
  jor  g17142(.dina(n17439), .dinb(n3912), .dout(n17440));
  jand g17143(.dina(n17428), .dinb(n3912), .dout(n17441));
  jand g17144(.dina(n17441), .dinb(n17438), .dout(n17442));
  jnot g17145(.din(n16814), .dout(n17443));
  jand g17146(.dina(asqrt[7] ), .dinb(n17443), .dout(n17444));
  jand g17147(.dina(n17444), .dinb(n16821), .dout(n17445));
  jor  g17148(.dina(n17445), .dinb(n16819), .dout(n17446));
  jand g17149(.dina(n17444), .dinb(n16822), .dout(n17447));
  jnot g17150(.din(n17447), .dout(n17448));
  jand g17151(.dina(n17448), .dinb(n17446), .dout(n17449));
  jnot g17152(.din(n17449), .dout(n17450));
  jor  g17153(.dina(n17450), .dinb(n17442), .dout(n17451));
  jand g17154(.dina(n17451), .dinb(n17440), .dout(n17452));
  jor  g17155(.dina(n17452), .dinb(n3907), .dout(n17453));
  jxor g17156(.dina(n16823), .dinb(n3912), .dout(n17454));
  jor  g17157(.dina(n17454), .dinb(n17140), .dout(n17455));
  jxor g17158(.dina(n17455), .dinb(n16834), .dout(n17456));
  jand g17159(.dina(n17452), .dinb(n3907), .dout(n17457));
  jor  g17160(.dina(n17457), .dinb(n17456), .dout(n17458));
  jand g17161(.dina(n17458), .dinb(n17453), .dout(n17459));
  jor  g17162(.dina(n17459), .dinb(n3376), .dout(n17460));
  jnot g17163(.din(n16839), .dout(n17461));
  jor  g17164(.dina(n17461), .dinb(n16837), .dout(n17462));
  jor  g17165(.dina(n17462), .dinb(n17140), .dout(n17463));
  jxor g17166(.dina(n17463), .dinb(n16848), .dout(n17464));
  jand g17167(.dina(n17453), .dinb(n3376), .dout(n17465));
  jand g17168(.dina(n17465), .dinb(n17458), .dout(n17466));
  jor  g17169(.dina(n17466), .dinb(n17464), .dout(n17467));
  jand g17170(.dina(n17467), .dinb(n17460), .dout(n17468));
  jor  g17171(.dina(n17468), .dinb(n3371), .dout(n17469));
  jand g17172(.dina(n17468), .dinb(n3371), .dout(n17470));
  jnot g17173(.din(n16851), .dout(n17471));
  jand g17174(.dina(asqrt[7] ), .dinb(n17471), .dout(n17472));
  jand g17175(.dina(n17472), .dinb(n16856), .dout(n17473));
  jor  g17176(.dina(n17473), .dinb(n16855), .dout(n17474));
  jand g17177(.dina(n17472), .dinb(n16857), .dout(n17475));
  jnot g17178(.din(n17475), .dout(n17476));
  jand g17179(.dina(n17476), .dinb(n17474), .dout(n17477));
  jnot g17180(.din(n17477), .dout(n17478));
  jor  g17181(.dina(n17478), .dinb(n17470), .dout(n17479));
  jand g17182(.dina(n17479), .dinb(n17469), .dout(n17480));
  jor  g17183(.dina(n17480), .dinb(n2875), .dout(n17481));
  jand g17184(.dina(n17469), .dinb(n2875), .dout(n17482));
  jand g17185(.dina(n17482), .dinb(n17479), .dout(n17483));
  jnot g17186(.din(n16859), .dout(n17484));
  jand g17187(.dina(asqrt[7] ), .dinb(n17484), .dout(n17485));
  jand g17188(.dina(n17485), .dinb(n16866), .dout(n17486));
  jor  g17189(.dina(n17486), .dinb(n16864), .dout(n17487));
  jand g17190(.dina(n17485), .dinb(n16867), .dout(n17488));
  jnot g17191(.din(n17488), .dout(n17489));
  jand g17192(.dina(n17489), .dinb(n17487), .dout(n17490));
  jnot g17193(.din(n17490), .dout(n17491));
  jor  g17194(.dina(n17491), .dinb(n17483), .dout(n17492));
  jand g17195(.dina(n17492), .dinb(n17481), .dout(n17493));
  jor  g17196(.dina(n17493), .dinb(n2870), .dout(n17494));
  jxor g17197(.dina(n16868), .dinb(n2875), .dout(n17495));
  jor  g17198(.dina(n17495), .dinb(n17140), .dout(n17496));
  jxor g17199(.dina(n17496), .dinb(n16879), .dout(n17497));
  jand g17200(.dina(n17493), .dinb(n2870), .dout(n17498));
  jor  g17201(.dina(n17498), .dinb(n17497), .dout(n17499));
  jand g17202(.dina(n17499), .dinb(n17494), .dout(n17500));
  jor  g17203(.dina(n17500), .dinb(n2425), .dout(n17501));
  jnot g17204(.din(n16884), .dout(n17502));
  jor  g17205(.dina(n17502), .dinb(n16882), .dout(n17503));
  jor  g17206(.dina(n17503), .dinb(n17140), .dout(n17504));
  jxor g17207(.dina(n17504), .dinb(n16893), .dout(n17505));
  jand g17208(.dina(n17494), .dinb(n2425), .dout(n17506));
  jand g17209(.dina(n17506), .dinb(n17499), .dout(n17507));
  jor  g17210(.dina(n17507), .dinb(n17505), .dout(n17508));
  jand g17211(.dina(n17508), .dinb(n17501), .dout(n17509));
  jor  g17212(.dina(n17509), .dinb(n2420), .dout(n17510));
  jand g17213(.dina(n17509), .dinb(n2420), .dout(n17511));
  jnot g17214(.din(n16896), .dout(n17512));
  jand g17215(.dina(asqrt[7] ), .dinb(n17512), .dout(n17513));
  jand g17216(.dina(n17513), .dinb(n16901), .dout(n17514));
  jor  g17217(.dina(n17514), .dinb(n16900), .dout(n17515));
  jand g17218(.dina(n17513), .dinb(n16902), .dout(n17516));
  jnot g17219(.din(n17516), .dout(n17517));
  jand g17220(.dina(n17517), .dinb(n17515), .dout(n17518));
  jnot g17221(.din(n17518), .dout(n17519));
  jor  g17222(.dina(n17519), .dinb(n17511), .dout(n17520));
  jand g17223(.dina(n17520), .dinb(n17510), .dout(n17521));
  jor  g17224(.dina(n17521), .dinb(n2010), .dout(n17522));
  jand g17225(.dina(n17510), .dinb(n2010), .dout(n17523));
  jand g17226(.dina(n17523), .dinb(n17520), .dout(n17524));
  jnot g17227(.din(n16904), .dout(n17525));
  jand g17228(.dina(asqrt[7] ), .dinb(n17525), .dout(n17526));
  jand g17229(.dina(n17526), .dinb(n16911), .dout(n17527));
  jor  g17230(.dina(n17527), .dinb(n16909), .dout(n17528));
  jand g17231(.dina(n17526), .dinb(n16912), .dout(n17529));
  jnot g17232(.din(n17529), .dout(n17530));
  jand g17233(.dina(n17530), .dinb(n17528), .dout(n17531));
  jnot g17234(.din(n17531), .dout(n17532));
  jor  g17235(.dina(n17532), .dinb(n17524), .dout(n17533));
  jand g17236(.dina(n17533), .dinb(n17522), .dout(n17534));
  jor  g17237(.dina(n17534), .dinb(n2005), .dout(n17535));
  jxor g17238(.dina(n16913), .dinb(n2010), .dout(n17536));
  jor  g17239(.dina(n17536), .dinb(n17140), .dout(n17537));
  jxor g17240(.dina(n17537), .dinb(n16924), .dout(n17538));
  jand g17241(.dina(n17534), .dinb(n2005), .dout(n17539));
  jor  g17242(.dina(n17539), .dinb(n17538), .dout(n17540));
  jand g17243(.dina(n17540), .dinb(n17535), .dout(n17541));
  jor  g17244(.dina(n17541), .dinb(n1646), .dout(n17542));
  jnot g17245(.din(n16929), .dout(n17543));
  jor  g17246(.dina(n17543), .dinb(n16927), .dout(n17544));
  jor  g17247(.dina(n17544), .dinb(n17140), .dout(n17545));
  jxor g17248(.dina(n17545), .dinb(n16938), .dout(n17546));
  jand g17249(.dina(n17535), .dinb(n1646), .dout(n17547));
  jand g17250(.dina(n17547), .dinb(n17540), .dout(n17548));
  jor  g17251(.dina(n17548), .dinb(n17546), .dout(n17549));
  jand g17252(.dina(n17549), .dinb(n17542), .dout(n17550));
  jor  g17253(.dina(n17550), .dinb(n1641), .dout(n17551));
  jand g17254(.dina(n17550), .dinb(n1641), .dout(n17552));
  jnot g17255(.din(n16941), .dout(n17553));
  jand g17256(.dina(asqrt[7] ), .dinb(n17553), .dout(n17554));
  jand g17257(.dina(n17554), .dinb(n16946), .dout(n17555));
  jor  g17258(.dina(n17555), .dinb(n16945), .dout(n17556));
  jand g17259(.dina(n17554), .dinb(n16947), .dout(n17557));
  jnot g17260(.din(n17557), .dout(n17558));
  jand g17261(.dina(n17558), .dinb(n17556), .dout(n17559));
  jnot g17262(.din(n17559), .dout(n17560));
  jor  g17263(.dina(n17560), .dinb(n17552), .dout(n17561));
  jand g17264(.dina(n17561), .dinb(n17551), .dout(n17562));
  jor  g17265(.dina(n17562), .dinb(n1317), .dout(n17563));
  jand g17266(.dina(n17551), .dinb(n1317), .dout(n17564));
  jand g17267(.dina(n17564), .dinb(n17561), .dout(n17565));
  jnot g17268(.din(n16949), .dout(n17566));
  jand g17269(.dina(asqrt[7] ), .dinb(n17566), .dout(n17567));
  jand g17270(.dina(n17567), .dinb(n16956), .dout(n17568));
  jor  g17271(.dina(n17568), .dinb(n16954), .dout(n17569));
  jand g17272(.dina(n17567), .dinb(n16957), .dout(n17570));
  jnot g17273(.din(n17570), .dout(n17571));
  jand g17274(.dina(n17571), .dinb(n17569), .dout(n17572));
  jnot g17275(.din(n17572), .dout(n17573));
  jor  g17276(.dina(n17573), .dinb(n17565), .dout(n17574));
  jand g17277(.dina(n17574), .dinb(n17563), .dout(n17575));
  jor  g17278(.dina(n17575), .dinb(n1312), .dout(n17576));
  jxor g17279(.dina(n16958), .dinb(n1317), .dout(n17577));
  jor  g17280(.dina(n17577), .dinb(n17140), .dout(n17578));
  jxor g17281(.dina(n17578), .dinb(n16969), .dout(n17579));
  jand g17282(.dina(n17575), .dinb(n1312), .dout(n17580));
  jor  g17283(.dina(n17580), .dinb(n17579), .dout(n17581));
  jand g17284(.dina(n17581), .dinb(n17576), .dout(n17582));
  jor  g17285(.dina(n17582), .dinb(n1039), .dout(n17583));
  jnot g17286(.din(n16974), .dout(n17584));
  jor  g17287(.dina(n17584), .dinb(n16972), .dout(n17585));
  jor  g17288(.dina(n17585), .dinb(n17140), .dout(n17586));
  jxor g17289(.dina(n17586), .dinb(n16983), .dout(n17587));
  jand g17290(.dina(n17576), .dinb(n1039), .dout(n17588));
  jand g17291(.dina(n17588), .dinb(n17581), .dout(n17589));
  jor  g17292(.dina(n17589), .dinb(n17587), .dout(n17590));
  jand g17293(.dina(n17590), .dinb(n17583), .dout(n17591));
  jor  g17294(.dina(n17591), .dinb(n1034), .dout(n17592));
  jand g17295(.dina(n17591), .dinb(n1034), .dout(n17593));
  jnot g17296(.din(n16986), .dout(n17594));
  jand g17297(.dina(asqrt[7] ), .dinb(n17594), .dout(n17595));
  jand g17298(.dina(n17595), .dinb(n16991), .dout(n17596));
  jor  g17299(.dina(n17596), .dinb(n16990), .dout(n17597));
  jand g17300(.dina(n17595), .dinb(n16992), .dout(n17598));
  jnot g17301(.din(n17598), .dout(n17599));
  jand g17302(.dina(n17599), .dinb(n17597), .dout(n17600));
  jnot g17303(.din(n17600), .dout(n17601));
  jor  g17304(.dina(n17601), .dinb(n17593), .dout(n17602));
  jand g17305(.dina(n17602), .dinb(n17592), .dout(n17603));
  jor  g17306(.dina(n17603), .dinb(n796), .dout(n17604));
  jand g17307(.dina(n17592), .dinb(n796), .dout(n17605));
  jand g17308(.dina(n17605), .dinb(n17602), .dout(n17606));
  jnot g17309(.din(n16994), .dout(n17607));
  jand g17310(.dina(asqrt[7] ), .dinb(n17607), .dout(n17608));
  jand g17311(.dina(n17608), .dinb(n17001), .dout(n17609));
  jor  g17312(.dina(n17609), .dinb(n16999), .dout(n17610));
  jand g17313(.dina(n17608), .dinb(n17002), .dout(n17611));
  jnot g17314(.din(n17611), .dout(n17612));
  jand g17315(.dina(n17612), .dinb(n17610), .dout(n17613));
  jnot g17316(.din(n17613), .dout(n17614));
  jor  g17317(.dina(n17614), .dinb(n17606), .dout(n17615));
  jand g17318(.dina(n17615), .dinb(n17604), .dout(n17616));
  jor  g17319(.dina(n17616), .dinb(n791), .dout(n17617));
  jxor g17320(.dina(n17003), .dinb(n796), .dout(n17618));
  jor  g17321(.dina(n17618), .dinb(n17140), .dout(n17619));
  jxor g17322(.dina(n17619), .dinb(n17014), .dout(n17620));
  jand g17323(.dina(n17616), .dinb(n791), .dout(n17621));
  jor  g17324(.dina(n17621), .dinb(n17620), .dout(n17622));
  jand g17325(.dina(n17622), .dinb(n17617), .dout(n17623));
  jor  g17326(.dina(n17623), .dinb(n595), .dout(n17624));
  jand g17327(.dina(n17617), .dinb(n595), .dout(n17625));
  jand g17328(.dina(n17625), .dinb(n17622), .dout(n17626));
  jnot g17329(.din(n17017), .dout(n17627));
  jand g17330(.dina(asqrt[7] ), .dinb(n17627), .dout(n17628));
  jand g17331(.dina(n17628), .dinb(n17024), .dout(n17629));
  jor  g17332(.dina(n17629), .dinb(n17022), .dout(n17630));
  jand g17333(.dina(n17628), .dinb(n17025), .dout(n17631));
  jnot g17334(.din(n17631), .dout(n17632));
  jand g17335(.dina(n17632), .dinb(n17630), .dout(n17633));
  jnot g17336(.din(n17633), .dout(n17634));
  jor  g17337(.dina(n17634), .dinb(n17626), .dout(n17635));
  jand g17338(.dina(n17635), .dinb(n17624), .dout(n17636));
  jor  g17339(.dina(n17636), .dinb(n590), .dout(n17637));
  jand g17340(.dina(n17636), .dinb(n590), .dout(n17638));
  jor  g17341(.dina(n17638), .dinb(n17143), .dout(n17639));
  jand g17342(.dina(n17639), .dinb(n17637), .dout(n17640));
  jor  g17343(.dina(n17640), .dinb(n430), .dout(n17641));
  jnot g17344(.din(n17033), .dout(n17642));
  jor  g17345(.dina(n17642), .dinb(n17031), .dout(n17643));
  jor  g17346(.dina(n17643), .dinb(n17140), .dout(n17644));
  jxor g17347(.dina(n17644), .dinb(n17042), .dout(n17645));
  jand g17348(.dina(n17637), .dinb(n430), .dout(n17646));
  jand g17349(.dina(n17646), .dinb(n17639), .dout(n17647));
  jor  g17350(.dina(n17647), .dinb(n17645), .dout(n17648));
  jand g17351(.dina(n17648), .dinb(n17641), .dout(n17649));
  jor  g17352(.dina(n17649), .dinb(n425), .dout(n17650));
  jxor g17353(.dina(n17044), .dinb(n430), .dout(n17651));
  jor  g17354(.dina(n17651), .dinb(n17140), .dout(n17652));
  jxor g17355(.dina(n17652), .dinb(n17055), .dout(n17653));
  jand g17356(.dina(n17649), .dinb(n425), .dout(n17654));
  jor  g17357(.dina(n17654), .dinb(n17653), .dout(n17655));
  jand g17358(.dina(n17655), .dinb(n17650), .dout(n17656));
  jor  g17359(.dina(n17656), .dinb(n305), .dout(n17657));
  jnot g17360(.din(n17060), .dout(n17658));
  jor  g17361(.dina(n17658), .dinb(n17058), .dout(n17659));
  jor  g17362(.dina(n17659), .dinb(n17140), .dout(n17660));
  jxor g17363(.dina(n17660), .dinb(n17069), .dout(n17661));
  jand g17364(.dina(n17650), .dinb(n305), .dout(n17662));
  jand g17365(.dina(n17662), .dinb(n17655), .dout(n17663));
  jor  g17366(.dina(n17663), .dinb(n17661), .dout(n17664));
  jand g17367(.dina(n17664), .dinb(n17657), .dout(n17665));
  jor  g17368(.dina(n17665), .dinb(n290), .dout(n17666));
  jand g17369(.dina(n17665), .dinb(n290), .dout(n17667));
  jnot g17370(.din(n17072), .dout(n17668));
  jand g17371(.dina(asqrt[7] ), .dinb(n17668), .dout(n17669));
  jand g17372(.dina(n17669), .dinb(n17077), .dout(n17670));
  jor  g17373(.dina(n17670), .dinb(n17076), .dout(n17671));
  jand g17374(.dina(n17669), .dinb(n17078), .dout(n17672));
  jnot g17375(.din(n17672), .dout(n17673));
  jand g17376(.dina(n17673), .dinb(n17671), .dout(n17674));
  jnot g17377(.din(n17674), .dout(n17675));
  jor  g17378(.dina(n17675), .dinb(n17667), .dout(n17676));
  jand g17379(.dina(n17676), .dinb(n17666), .dout(n17677));
  jor  g17380(.dina(n17677), .dinb(n223), .dout(n17678));
  jand g17381(.dina(n17666), .dinb(n223), .dout(n17679));
  jand g17382(.dina(n17679), .dinb(n17676), .dout(n17680));
  jnot g17383(.din(n17080), .dout(n17681));
  jand g17384(.dina(asqrt[7] ), .dinb(n17681), .dout(n17682));
  jand g17385(.dina(n17682), .dinb(n17087), .dout(n17683));
  jor  g17386(.dina(n17683), .dinb(n17085), .dout(n17684));
  jand g17387(.dina(n17682), .dinb(n17088), .dout(n17685));
  jnot g17388(.din(n17685), .dout(n17686));
  jand g17389(.dina(n17686), .dinb(n17684), .dout(n17687));
  jnot g17390(.din(n17687), .dout(n17688));
  jor  g17391(.dina(n17688), .dinb(n17680), .dout(n17689));
  jand g17392(.dina(n17689), .dinb(n17678), .dout(n17690));
  jor  g17393(.dina(n17690), .dinb(n199), .dout(n17691));
  jand g17394(.dina(n17690), .dinb(n199), .dout(n17692));
  jxor g17395(.dina(n17089), .dinb(n223), .dout(n17693));
  jor  g17396(.dina(n17693), .dinb(n17140), .dout(n17694));
  jxor g17397(.dina(n17694), .dinb(n17100), .dout(n17695));
  jor  g17398(.dina(n17695), .dinb(n17692), .dout(n17696));
  jand g17399(.dina(n17696), .dinb(n17691), .dout(n17697));
  jnot g17400(.din(n17105), .dout(n17698));
  jor  g17401(.dina(n17698), .dinb(n17103), .dout(n17699));
  jor  g17402(.dina(n17699), .dinb(n17140), .dout(n17700));
  jxor g17403(.dina(n17700), .dinb(n17114), .dout(n17701));
  jand g17404(.dina(asqrt[7] ), .dinb(n17128), .dout(n17702));
  jand g17405(.dina(n17702), .dinb(n17116), .dout(n17703));
  jor  g17406(.dina(n17703), .dinb(n17162), .dout(n17704));
  jor  g17407(.dina(n17704), .dinb(n17701), .dout(n17705));
  jor  g17408(.dina(n17705), .dinb(n17697), .dout(n17706));
  jand g17409(.dina(n17706), .dinb(n194), .dout(n17707));
  jand g17410(.dina(n17701), .dinb(n17697), .dout(n17708));
  jor  g17411(.dina(n17702), .dinb(n17116), .dout(n17709));
  jand g17412(.dina(n17128), .dinb(n17116), .dout(n17710));
  jor  g17413(.dina(n17710), .dinb(n194), .dout(n17711));
  jnot g17414(.din(n17711), .dout(n17712));
  jand g17415(.dina(n17712), .dinb(n17709), .dout(n17713));
  jor  g17416(.dina(n17713), .dinb(n17708), .dout(n17716));
  jor  g17417(.dina(n17716), .dinb(n17707), .dout(asqrt[6] ));
  jxor g17418(.dina(n17636), .dinb(n590), .dout(n17718));
  jand g17419(.dina(n17718), .dinb(asqrt[6] ), .dout(n17719));
  jxor g17420(.dina(n17719), .dinb(n17143), .dout(n17720));
  jand g17421(.dina(asqrt[6] ), .dinb(a[12] ), .dout(n17721));
  jnot g17422(.din(a[10] ), .dout(n17722));
  jnot g17423(.din(a[11] ), .dout(n17723));
  jand g17424(.dina(n17145), .dinb(n17723), .dout(n17724));
  jand g17425(.dina(n17724), .dinb(n17722), .dout(n17725));
  jor  g17426(.dina(n17725), .dinb(n17721), .dout(n17726));
  jand g17427(.dina(n17726), .dinb(asqrt[7] ), .dout(n17727));
  jand g17428(.dina(asqrt[6] ), .dinb(n17145), .dout(n17728));
  jxor g17429(.dina(n17728), .dinb(n17146), .dout(n17729));
  jor  g17430(.dina(n17726), .dinb(asqrt[7] ), .dout(n17730));
  jand g17431(.dina(n17730), .dinb(n17729), .dout(n17731));
  jor  g17432(.dina(n17731), .dinb(n17727), .dout(n17732));
  jand g17433(.dina(n17732), .dinb(asqrt[8] ), .dout(n17733));
  jor  g17434(.dina(n17727), .dinb(asqrt[8] ), .dout(n17734));
  jor  g17435(.dina(n17734), .dinb(n17731), .dout(n17735));
  jand g17436(.dina(n17728), .dinb(n17146), .dout(n17736));
  jnot g17437(.din(n17707), .dout(n17737));
  jnot g17438(.din(n17708), .dout(n17738));
  jnot g17439(.din(n17713), .dout(n17739));
  jand g17440(.dina(n17739), .dinb(asqrt[7] ), .dout(n17740));
  jand g17441(.dina(n17740), .dinb(n17738), .dout(n17741));
  jand g17442(.dina(n17741), .dinb(n17737), .dout(n17742));
  jor  g17443(.dina(n17742), .dinb(n17736), .dout(n17743));
  jxor g17444(.dina(n17743), .dinb(n16523), .dout(n17744));
  jand g17445(.dina(n17744), .dinb(n17735), .dout(n17745));
  jor  g17446(.dina(n17745), .dinb(n17733), .dout(n17746));
  jand g17447(.dina(n17746), .dinb(asqrt[9] ), .dout(n17747));
  jor  g17448(.dina(n17746), .dinb(asqrt[9] ), .dout(n17748));
  jxor g17449(.dina(n17150), .dinb(n17135), .dout(n17749));
  jand g17450(.dina(n17749), .dinb(asqrt[6] ), .dout(n17750));
  jxor g17451(.dina(n17750), .dinb(n17153), .dout(n17751));
  jnot g17452(.din(n17751), .dout(n17752));
  jand g17453(.dina(n17752), .dinb(n17748), .dout(n17753));
  jor  g17454(.dina(n17753), .dinb(n17747), .dout(n17754));
  jand g17455(.dina(n17754), .dinb(asqrt[10] ), .dout(n17755));
  jnot g17456(.din(n17159), .dout(n17756));
  jand g17457(.dina(n17756), .dinb(n17157), .dout(n17757));
  jand g17458(.dina(n17757), .dinb(asqrt[6] ), .dout(n17758));
  jxor g17459(.dina(n17758), .dinb(n17167), .dout(n17759));
  jnot g17460(.din(n17759), .dout(n17760));
  jor  g17461(.dina(n17747), .dinb(asqrt[10] ), .dout(n17761));
  jor  g17462(.dina(n17761), .dinb(n17753), .dout(n17762));
  jand g17463(.dina(n17762), .dinb(n17760), .dout(n17763));
  jor  g17464(.dina(n17763), .dinb(n17755), .dout(n17764));
  jand g17465(.dina(n17764), .dinb(asqrt[11] ), .dout(n17765));
  jor  g17466(.dina(n17764), .dinb(asqrt[11] ), .dout(n17766));
  jnot g17467(.din(n17174), .dout(n17767));
  jxor g17468(.dina(n17169), .dinb(n15950), .dout(n17768));
  jand g17469(.dina(n17768), .dinb(asqrt[6] ), .dout(n17769));
  jxor g17470(.dina(n17769), .dinb(n17767), .dout(n17770));
  jand g17471(.dina(n17770), .dinb(n17766), .dout(n17771));
  jor  g17472(.dina(n17771), .dinb(n17765), .dout(n17772));
  jand g17473(.dina(n17772), .dinb(asqrt[12] ), .dout(n17773));
  jor  g17474(.dina(n17765), .dinb(asqrt[12] ), .dout(n17774));
  jor  g17475(.dina(n17774), .dinb(n17771), .dout(n17775));
  jnot g17476(.din(n17181), .dout(n17776));
  jnot g17477(.din(n17183), .dout(n17777));
  jand g17478(.dina(asqrt[6] ), .dinb(n17177), .dout(n17778));
  jand g17479(.dina(n17778), .dinb(n17777), .dout(n17779));
  jor  g17480(.dina(n17779), .dinb(n17776), .dout(n17780));
  jnot g17481(.din(n17184), .dout(n17781));
  jand g17482(.dina(n17778), .dinb(n17781), .dout(n17782));
  jnot g17483(.din(n17782), .dout(n17783));
  jand g17484(.dina(n17783), .dinb(n17780), .dout(n17784));
  jand g17485(.dina(n17784), .dinb(n17775), .dout(n17785));
  jor  g17486(.dina(n17785), .dinb(n17773), .dout(n17786));
  jand g17487(.dina(n17786), .dinb(asqrt[13] ), .dout(n17787));
  jor  g17488(.dina(n17786), .dinb(asqrt[13] ), .dout(n17788));
  jxor g17489(.dina(n17185), .dinb(n14816), .dout(n17789));
  jand g17490(.dina(n17789), .dinb(asqrt[6] ), .dout(n17790));
  jxor g17491(.dina(n17790), .dinb(n17190), .dout(n17791));
  jand g17492(.dina(n17791), .dinb(n17788), .dout(n17792));
  jor  g17493(.dina(n17792), .dinb(n17787), .dout(n17793));
  jand g17494(.dina(n17793), .dinb(asqrt[14] ), .dout(n17794));
  jnot g17495(.din(n17196), .dout(n17795));
  jand g17496(.dina(n17795), .dinb(n17194), .dout(n17796));
  jand g17497(.dina(n17796), .dinb(asqrt[6] ), .dout(n17797));
  jxor g17498(.dina(n17797), .dinb(n17205), .dout(n17798));
  jnot g17499(.din(n17798), .dout(n17799));
  jor  g17500(.dina(n17787), .dinb(asqrt[14] ), .dout(n17800));
  jor  g17501(.dina(n17800), .dinb(n17792), .dout(n17801));
  jand g17502(.dina(n17801), .dinb(n17799), .dout(n17802));
  jor  g17503(.dina(n17802), .dinb(n17794), .dout(n17803));
  jand g17504(.dina(n17803), .dinb(asqrt[15] ), .dout(n17804));
  jor  g17505(.dina(n17803), .dinb(asqrt[15] ), .dout(n17805));
  jxor g17506(.dina(n17207), .dinb(n13718), .dout(n17806));
  jand g17507(.dina(n17806), .dinb(asqrt[6] ), .dout(n17807));
  jxor g17508(.dina(n17807), .dinb(n17213), .dout(n17808));
  jand g17509(.dina(n17808), .dinb(n17805), .dout(n17809));
  jor  g17510(.dina(n17809), .dinb(n17804), .dout(n17810));
  jand g17511(.dina(n17810), .dinb(asqrt[16] ), .dout(n17811));
  jor  g17512(.dina(n17804), .dinb(asqrt[16] ), .dout(n17812));
  jor  g17513(.dina(n17812), .dinb(n17809), .dout(n17813));
  jnot g17514(.din(n17221), .dout(n17814));
  jnot g17515(.din(n17223), .dout(n17815));
  jand g17516(.dina(asqrt[6] ), .dinb(n17217), .dout(n17816));
  jand g17517(.dina(n17816), .dinb(n17815), .dout(n17817));
  jor  g17518(.dina(n17817), .dinb(n17814), .dout(n17818));
  jnot g17519(.din(n17224), .dout(n17819));
  jand g17520(.dina(n17816), .dinb(n17819), .dout(n17820));
  jnot g17521(.din(n17820), .dout(n17821));
  jand g17522(.dina(n17821), .dinb(n17818), .dout(n17822));
  jand g17523(.dina(n17822), .dinb(n17813), .dout(n17823));
  jor  g17524(.dina(n17823), .dinb(n17811), .dout(n17824));
  jand g17525(.dina(n17824), .dinb(asqrt[17] ), .dout(n17825));
  jxor g17526(.dina(n17225), .dinb(n12670), .dout(n17826));
  jand g17527(.dina(n17826), .dinb(asqrt[6] ), .dout(n17827));
  jxor g17528(.dina(n17827), .dinb(n17232), .dout(n17828));
  jnot g17529(.din(n17828), .dout(n17829));
  jor  g17530(.dina(n17824), .dinb(asqrt[17] ), .dout(n17830));
  jand g17531(.dina(n17830), .dinb(n17829), .dout(n17831));
  jor  g17532(.dina(n17831), .dinb(n17825), .dout(n17832));
  jand g17533(.dina(n17832), .dinb(asqrt[18] ), .dout(n17833));
  jnot g17534(.din(n17237), .dout(n17834));
  jand g17535(.dina(n17834), .dinb(n17235), .dout(n17835));
  jand g17536(.dina(n17835), .dinb(asqrt[6] ), .dout(n17836));
  jxor g17537(.dina(n17836), .dinb(n17245), .dout(n17837));
  jnot g17538(.din(n17837), .dout(n17838));
  jor  g17539(.dina(n17825), .dinb(asqrt[18] ), .dout(n17839));
  jor  g17540(.dina(n17839), .dinb(n17831), .dout(n17840));
  jand g17541(.dina(n17840), .dinb(n17838), .dout(n17841));
  jor  g17542(.dina(n17841), .dinb(n17833), .dout(n17842));
  jand g17543(.dina(n17842), .dinb(asqrt[19] ), .dout(n17843));
  jor  g17544(.dina(n17842), .dinb(asqrt[19] ), .dout(n17844));
  jnot g17545(.din(n17251), .dout(n17845));
  jnot g17546(.din(n17252), .dout(n17846));
  jand g17547(.dina(asqrt[6] ), .dinb(n17248), .dout(n17847));
  jand g17548(.dina(n17847), .dinb(n17846), .dout(n17848));
  jor  g17549(.dina(n17848), .dinb(n17845), .dout(n17849));
  jnot g17550(.din(n17253), .dout(n17850));
  jand g17551(.dina(n17847), .dinb(n17850), .dout(n17851));
  jnot g17552(.din(n17851), .dout(n17852));
  jand g17553(.dina(n17852), .dinb(n17849), .dout(n17853));
  jand g17554(.dina(n17853), .dinb(n17844), .dout(n17854));
  jor  g17555(.dina(n17854), .dinb(n17843), .dout(n17855));
  jand g17556(.dina(n17855), .dinb(asqrt[20] ), .dout(n17856));
  jor  g17557(.dina(n17843), .dinb(asqrt[20] ), .dout(n17857));
  jor  g17558(.dina(n17857), .dinb(n17854), .dout(n17858));
  jnot g17559(.din(n17259), .dout(n17859));
  jnot g17560(.din(n17261), .dout(n17860));
  jand g17561(.dina(asqrt[6] ), .dinb(n17255), .dout(n17861));
  jand g17562(.dina(n17861), .dinb(n17860), .dout(n17862));
  jor  g17563(.dina(n17862), .dinb(n17859), .dout(n17863));
  jnot g17564(.din(n17262), .dout(n17864));
  jand g17565(.dina(n17861), .dinb(n17864), .dout(n17865));
  jnot g17566(.din(n17865), .dout(n17866));
  jand g17567(.dina(n17866), .dinb(n17863), .dout(n17867));
  jand g17568(.dina(n17867), .dinb(n17858), .dout(n17868));
  jor  g17569(.dina(n17868), .dinb(n17856), .dout(n17869));
  jand g17570(.dina(n17869), .dinb(asqrt[21] ), .dout(n17870));
  jxor g17571(.dina(n17263), .dinb(n10696), .dout(n17871));
  jand g17572(.dina(n17871), .dinb(asqrt[6] ), .dout(n17872));
  jxor g17573(.dina(n17872), .dinb(n17273), .dout(n17873));
  jnot g17574(.din(n17873), .dout(n17874));
  jor  g17575(.dina(n17869), .dinb(asqrt[21] ), .dout(n17875));
  jand g17576(.dina(n17875), .dinb(n17874), .dout(n17876));
  jor  g17577(.dina(n17876), .dinb(n17870), .dout(n17877));
  jand g17578(.dina(n17877), .dinb(asqrt[22] ), .dout(n17878));
  jnot g17579(.din(n17278), .dout(n17879));
  jand g17580(.dina(n17879), .dinb(n17276), .dout(n17880));
  jand g17581(.dina(n17880), .dinb(asqrt[6] ), .dout(n17881));
  jxor g17582(.dina(n17881), .dinb(n17286), .dout(n17882));
  jnot g17583(.din(n17882), .dout(n17883));
  jor  g17584(.dina(n17870), .dinb(asqrt[22] ), .dout(n17884));
  jor  g17585(.dina(n17884), .dinb(n17876), .dout(n17885));
  jand g17586(.dina(n17885), .dinb(n17883), .dout(n17886));
  jor  g17587(.dina(n17886), .dinb(n17878), .dout(n17887));
  jand g17588(.dina(n17887), .dinb(asqrt[23] ), .dout(n17888));
  jor  g17589(.dina(n17887), .dinb(asqrt[23] ), .dout(n17889));
  jnot g17590(.din(n17292), .dout(n17890));
  jnot g17591(.din(n17293), .dout(n17891));
  jand g17592(.dina(asqrt[6] ), .dinb(n17289), .dout(n17892));
  jand g17593(.dina(n17892), .dinb(n17891), .dout(n17893));
  jor  g17594(.dina(n17893), .dinb(n17890), .dout(n17894));
  jnot g17595(.din(n17294), .dout(n17895));
  jand g17596(.dina(n17892), .dinb(n17895), .dout(n17896));
  jnot g17597(.din(n17896), .dout(n17897));
  jand g17598(.dina(n17897), .dinb(n17894), .dout(n17898));
  jand g17599(.dina(n17898), .dinb(n17889), .dout(n17899));
  jor  g17600(.dina(n17899), .dinb(n17888), .dout(n17900));
  jand g17601(.dina(n17900), .dinb(asqrt[24] ), .dout(n17901));
  jor  g17602(.dina(n17888), .dinb(asqrt[24] ), .dout(n17902));
  jor  g17603(.dina(n17902), .dinb(n17899), .dout(n17903));
  jnot g17604(.din(n17300), .dout(n17904));
  jnot g17605(.din(n17302), .dout(n17905));
  jand g17606(.dina(asqrt[6] ), .dinb(n17296), .dout(n17906));
  jand g17607(.dina(n17906), .dinb(n17905), .dout(n17907));
  jor  g17608(.dina(n17907), .dinb(n17904), .dout(n17908));
  jnot g17609(.din(n17303), .dout(n17909));
  jand g17610(.dina(n17906), .dinb(n17909), .dout(n17910));
  jnot g17611(.din(n17910), .dout(n17911));
  jand g17612(.dina(n17911), .dinb(n17908), .dout(n17912));
  jand g17613(.dina(n17912), .dinb(n17903), .dout(n17913));
  jor  g17614(.dina(n17913), .dinb(n17901), .dout(n17914));
  jand g17615(.dina(n17914), .dinb(asqrt[25] ), .dout(n17915));
  jxor g17616(.dina(n17304), .dinb(n8893), .dout(n17916));
  jand g17617(.dina(n17916), .dinb(asqrt[6] ), .dout(n17917));
  jxor g17618(.dina(n17917), .dinb(n17314), .dout(n17918));
  jnot g17619(.din(n17918), .dout(n17919));
  jor  g17620(.dina(n17914), .dinb(asqrt[25] ), .dout(n17920));
  jand g17621(.dina(n17920), .dinb(n17919), .dout(n17921));
  jor  g17622(.dina(n17921), .dinb(n17915), .dout(n17922));
  jand g17623(.dina(n17922), .dinb(asqrt[26] ), .dout(n17923));
  jnot g17624(.din(n17319), .dout(n17924));
  jand g17625(.dina(n17924), .dinb(n17317), .dout(n17925));
  jand g17626(.dina(n17925), .dinb(asqrt[6] ), .dout(n17926));
  jxor g17627(.dina(n17926), .dinb(n17327), .dout(n17927));
  jnot g17628(.din(n17927), .dout(n17928));
  jor  g17629(.dina(n17915), .dinb(asqrt[26] ), .dout(n17929));
  jor  g17630(.dina(n17929), .dinb(n17921), .dout(n17930));
  jand g17631(.dina(n17930), .dinb(n17928), .dout(n17931));
  jor  g17632(.dina(n17931), .dinb(n17923), .dout(n17932));
  jand g17633(.dina(n17932), .dinb(asqrt[27] ), .dout(n17933));
  jor  g17634(.dina(n17932), .dinb(asqrt[27] ), .dout(n17934));
  jnot g17635(.din(n17333), .dout(n17935));
  jnot g17636(.din(n17334), .dout(n17936));
  jand g17637(.dina(asqrt[6] ), .dinb(n17330), .dout(n17937));
  jand g17638(.dina(n17937), .dinb(n17936), .dout(n17938));
  jor  g17639(.dina(n17938), .dinb(n17935), .dout(n17939));
  jnot g17640(.din(n17335), .dout(n17940));
  jand g17641(.dina(n17937), .dinb(n17940), .dout(n17941));
  jnot g17642(.din(n17941), .dout(n17942));
  jand g17643(.dina(n17942), .dinb(n17939), .dout(n17943));
  jand g17644(.dina(n17943), .dinb(n17934), .dout(n17944));
  jor  g17645(.dina(n17944), .dinb(n17933), .dout(n17945));
  jand g17646(.dina(n17945), .dinb(asqrt[28] ), .dout(n17946));
  jor  g17647(.dina(n17933), .dinb(asqrt[28] ), .dout(n17947));
  jor  g17648(.dina(n17947), .dinb(n17944), .dout(n17948));
  jnot g17649(.din(n17341), .dout(n17949));
  jnot g17650(.din(n17343), .dout(n17950));
  jand g17651(.dina(asqrt[6] ), .dinb(n17337), .dout(n17951));
  jand g17652(.dina(n17951), .dinb(n17950), .dout(n17952));
  jor  g17653(.dina(n17952), .dinb(n17949), .dout(n17953));
  jnot g17654(.din(n17344), .dout(n17954));
  jand g17655(.dina(n17951), .dinb(n17954), .dout(n17955));
  jnot g17656(.din(n17955), .dout(n17956));
  jand g17657(.dina(n17956), .dinb(n17953), .dout(n17957));
  jand g17658(.dina(n17957), .dinb(n17948), .dout(n17958));
  jor  g17659(.dina(n17958), .dinb(n17946), .dout(n17959));
  jand g17660(.dina(n17959), .dinb(asqrt[29] ), .dout(n17960));
  jxor g17661(.dina(n17345), .dinb(n7260), .dout(n17961));
  jand g17662(.dina(n17961), .dinb(asqrt[6] ), .dout(n17962));
  jxor g17663(.dina(n17962), .dinb(n17355), .dout(n17963));
  jnot g17664(.din(n17963), .dout(n17964));
  jor  g17665(.dina(n17959), .dinb(asqrt[29] ), .dout(n17965));
  jand g17666(.dina(n17965), .dinb(n17964), .dout(n17966));
  jor  g17667(.dina(n17966), .dinb(n17960), .dout(n17967));
  jand g17668(.dina(n17967), .dinb(asqrt[30] ), .dout(n17968));
  jnot g17669(.din(n17360), .dout(n17969));
  jand g17670(.dina(n17969), .dinb(n17358), .dout(n17970));
  jand g17671(.dina(n17970), .dinb(asqrt[6] ), .dout(n17971));
  jxor g17672(.dina(n17971), .dinb(n17368), .dout(n17972));
  jnot g17673(.din(n17972), .dout(n17973));
  jor  g17674(.dina(n17960), .dinb(asqrt[30] ), .dout(n17974));
  jor  g17675(.dina(n17974), .dinb(n17966), .dout(n17975));
  jand g17676(.dina(n17975), .dinb(n17973), .dout(n17976));
  jor  g17677(.dina(n17976), .dinb(n17968), .dout(n17977));
  jand g17678(.dina(n17977), .dinb(asqrt[31] ), .dout(n17978));
  jor  g17679(.dina(n17977), .dinb(asqrt[31] ), .dout(n17979));
  jnot g17680(.din(n17374), .dout(n17980));
  jnot g17681(.din(n17375), .dout(n17981));
  jand g17682(.dina(asqrt[6] ), .dinb(n17371), .dout(n17982));
  jand g17683(.dina(n17982), .dinb(n17981), .dout(n17983));
  jor  g17684(.dina(n17983), .dinb(n17980), .dout(n17984));
  jnot g17685(.din(n17376), .dout(n17985));
  jand g17686(.dina(n17982), .dinb(n17985), .dout(n17986));
  jnot g17687(.din(n17986), .dout(n17987));
  jand g17688(.dina(n17987), .dinb(n17984), .dout(n17988));
  jand g17689(.dina(n17988), .dinb(n17979), .dout(n17989));
  jor  g17690(.dina(n17989), .dinb(n17978), .dout(n17990));
  jand g17691(.dina(n17990), .dinb(asqrt[32] ), .dout(n17991));
  jor  g17692(.dina(n17978), .dinb(asqrt[32] ), .dout(n17992));
  jor  g17693(.dina(n17992), .dinb(n17989), .dout(n17993));
  jnot g17694(.din(n17382), .dout(n17994));
  jnot g17695(.din(n17384), .dout(n17995));
  jand g17696(.dina(asqrt[6] ), .dinb(n17378), .dout(n17996));
  jand g17697(.dina(n17996), .dinb(n17995), .dout(n17997));
  jor  g17698(.dina(n17997), .dinb(n17994), .dout(n17998));
  jnot g17699(.din(n17385), .dout(n17999));
  jand g17700(.dina(n17996), .dinb(n17999), .dout(n18000));
  jnot g17701(.din(n18000), .dout(n18001));
  jand g17702(.dina(n18001), .dinb(n17998), .dout(n18002));
  jand g17703(.dina(n18002), .dinb(n17993), .dout(n18003));
  jor  g17704(.dina(n18003), .dinb(n17991), .dout(n18004));
  jand g17705(.dina(n18004), .dinb(asqrt[33] ), .dout(n18005));
  jxor g17706(.dina(n17386), .dinb(n5788), .dout(n18006));
  jand g17707(.dina(n18006), .dinb(asqrt[6] ), .dout(n18007));
  jxor g17708(.dina(n18007), .dinb(n17396), .dout(n18008));
  jnot g17709(.din(n18008), .dout(n18009));
  jor  g17710(.dina(n18004), .dinb(asqrt[33] ), .dout(n18010));
  jand g17711(.dina(n18010), .dinb(n18009), .dout(n18011));
  jor  g17712(.dina(n18011), .dinb(n18005), .dout(n18012));
  jand g17713(.dina(n18012), .dinb(asqrt[34] ), .dout(n18013));
  jnot g17714(.din(n17401), .dout(n18014));
  jand g17715(.dina(n18014), .dinb(n17399), .dout(n18015));
  jand g17716(.dina(n18015), .dinb(asqrt[6] ), .dout(n18016));
  jxor g17717(.dina(n18016), .dinb(n17409), .dout(n18017));
  jnot g17718(.din(n18017), .dout(n18018));
  jor  g17719(.dina(n18005), .dinb(asqrt[34] ), .dout(n18019));
  jor  g17720(.dina(n18019), .dinb(n18011), .dout(n18020));
  jand g17721(.dina(n18020), .dinb(n18018), .dout(n18021));
  jor  g17722(.dina(n18021), .dinb(n18013), .dout(n18022));
  jand g17723(.dina(n18022), .dinb(asqrt[35] ), .dout(n18023));
  jor  g17724(.dina(n18022), .dinb(asqrt[35] ), .dout(n18024));
  jnot g17725(.din(n17415), .dout(n18025));
  jnot g17726(.din(n17416), .dout(n18026));
  jand g17727(.dina(asqrt[6] ), .dinb(n17412), .dout(n18027));
  jand g17728(.dina(n18027), .dinb(n18026), .dout(n18028));
  jor  g17729(.dina(n18028), .dinb(n18025), .dout(n18029));
  jnot g17730(.din(n17417), .dout(n18030));
  jand g17731(.dina(n18027), .dinb(n18030), .dout(n18031));
  jnot g17732(.din(n18031), .dout(n18032));
  jand g17733(.dina(n18032), .dinb(n18029), .dout(n18033));
  jand g17734(.dina(n18033), .dinb(n18024), .dout(n18034));
  jor  g17735(.dina(n18034), .dinb(n18023), .dout(n18035));
  jand g17736(.dina(n18035), .dinb(asqrt[36] ), .dout(n18036));
  jor  g17737(.dina(n18023), .dinb(asqrt[36] ), .dout(n18037));
  jor  g17738(.dina(n18037), .dinb(n18034), .dout(n18038));
  jnot g17739(.din(n17423), .dout(n18039));
  jnot g17740(.din(n17425), .dout(n18040));
  jand g17741(.dina(asqrt[6] ), .dinb(n17419), .dout(n18041));
  jand g17742(.dina(n18041), .dinb(n18040), .dout(n18042));
  jor  g17743(.dina(n18042), .dinb(n18039), .dout(n18043));
  jnot g17744(.din(n17426), .dout(n18044));
  jand g17745(.dina(n18041), .dinb(n18044), .dout(n18045));
  jnot g17746(.din(n18045), .dout(n18046));
  jand g17747(.dina(n18046), .dinb(n18043), .dout(n18047));
  jand g17748(.dina(n18047), .dinb(n18038), .dout(n18048));
  jor  g17749(.dina(n18048), .dinb(n18036), .dout(n18049));
  jand g17750(.dina(n18049), .dinb(asqrt[37] ), .dout(n18050));
  jxor g17751(.dina(n17427), .dinb(n4494), .dout(n18051));
  jand g17752(.dina(n18051), .dinb(asqrt[6] ), .dout(n18052));
  jxor g17753(.dina(n18052), .dinb(n17437), .dout(n18053));
  jnot g17754(.din(n18053), .dout(n18054));
  jor  g17755(.dina(n18049), .dinb(asqrt[37] ), .dout(n18055));
  jand g17756(.dina(n18055), .dinb(n18054), .dout(n18056));
  jor  g17757(.dina(n18056), .dinb(n18050), .dout(n18057));
  jand g17758(.dina(n18057), .dinb(asqrt[38] ), .dout(n18058));
  jnot g17759(.din(n17442), .dout(n18059));
  jand g17760(.dina(n18059), .dinb(n17440), .dout(n18060));
  jand g17761(.dina(n18060), .dinb(asqrt[6] ), .dout(n18061));
  jxor g17762(.dina(n18061), .dinb(n17450), .dout(n18062));
  jnot g17763(.din(n18062), .dout(n18063));
  jor  g17764(.dina(n18050), .dinb(asqrt[38] ), .dout(n18064));
  jor  g17765(.dina(n18064), .dinb(n18056), .dout(n18065));
  jand g17766(.dina(n18065), .dinb(n18063), .dout(n18066));
  jor  g17767(.dina(n18066), .dinb(n18058), .dout(n18067));
  jand g17768(.dina(n18067), .dinb(asqrt[39] ), .dout(n18068));
  jor  g17769(.dina(n18067), .dinb(asqrt[39] ), .dout(n18069));
  jnot g17770(.din(n17456), .dout(n18070));
  jnot g17771(.din(n17457), .dout(n18071));
  jand g17772(.dina(asqrt[6] ), .dinb(n17453), .dout(n18072));
  jand g17773(.dina(n18072), .dinb(n18071), .dout(n18073));
  jor  g17774(.dina(n18073), .dinb(n18070), .dout(n18074));
  jnot g17775(.din(n17458), .dout(n18075));
  jand g17776(.dina(n18072), .dinb(n18075), .dout(n18076));
  jnot g17777(.din(n18076), .dout(n18077));
  jand g17778(.dina(n18077), .dinb(n18074), .dout(n18078));
  jand g17779(.dina(n18078), .dinb(n18069), .dout(n18079));
  jor  g17780(.dina(n18079), .dinb(n18068), .dout(n18080));
  jand g17781(.dina(n18080), .dinb(asqrt[40] ), .dout(n18081));
  jor  g17782(.dina(n18068), .dinb(asqrt[40] ), .dout(n18082));
  jor  g17783(.dina(n18082), .dinb(n18079), .dout(n18083));
  jnot g17784(.din(n17464), .dout(n18084));
  jnot g17785(.din(n17466), .dout(n18085));
  jand g17786(.dina(asqrt[6] ), .dinb(n17460), .dout(n18086));
  jand g17787(.dina(n18086), .dinb(n18085), .dout(n18087));
  jor  g17788(.dina(n18087), .dinb(n18084), .dout(n18088));
  jnot g17789(.din(n17467), .dout(n18089));
  jand g17790(.dina(n18086), .dinb(n18089), .dout(n18090));
  jnot g17791(.din(n18090), .dout(n18091));
  jand g17792(.dina(n18091), .dinb(n18088), .dout(n18092));
  jand g17793(.dina(n18092), .dinb(n18083), .dout(n18093));
  jor  g17794(.dina(n18093), .dinb(n18081), .dout(n18094));
  jand g17795(.dina(n18094), .dinb(asqrt[41] ), .dout(n18095));
  jxor g17796(.dina(n17468), .dinb(n3371), .dout(n18096));
  jand g17797(.dina(n18096), .dinb(asqrt[6] ), .dout(n18097));
  jxor g17798(.dina(n18097), .dinb(n17478), .dout(n18098));
  jnot g17799(.din(n18098), .dout(n18099));
  jor  g17800(.dina(n18094), .dinb(asqrt[41] ), .dout(n18100));
  jand g17801(.dina(n18100), .dinb(n18099), .dout(n18101));
  jor  g17802(.dina(n18101), .dinb(n18095), .dout(n18102));
  jand g17803(.dina(n18102), .dinb(asqrt[42] ), .dout(n18103));
  jnot g17804(.din(n17483), .dout(n18104));
  jand g17805(.dina(n18104), .dinb(n17481), .dout(n18105));
  jand g17806(.dina(n18105), .dinb(asqrt[6] ), .dout(n18106));
  jxor g17807(.dina(n18106), .dinb(n17491), .dout(n18107));
  jnot g17808(.din(n18107), .dout(n18108));
  jor  g17809(.dina(n18095), .dinb(asqrt[42] ), .dout(n18109));
  jor  g17810(.dina(n18109), .dinb(n18101), .dout(n18110));
  jand g17811(.dina(n18110), .dinb(n18108), .dout(n18111));
  jor  g17812(.dina(n18111), .dinb(n18103), .dout(n18112));
  jand g17813(.dina(n18112), .dinb(asqrt[43] ), .dout(n18113));
  jor  g17814(.dina(n18112), .dinb(asqrt[43] ), .dout(n18114));
  jnot g17815(.din(n17497), .dout(n18115));
  jnot g17816(.din(n17498), .dout(n18116));
  jand g17817(.dina(asqrt[6] ), .dinb(n17494), .dout(n18117));
  jand g17818(.dina(n18117), .dinb(n18116), .dout(n18118));
  jor  g17819(.dina(n18118), .dinb(n18115), .dout(n18119));
  jnot g17820(.din(n17499), .dout(n18120));
  jand g17821(.dina(n18117), .dinb(n18120), .dout(n18121));
  jnot g17822(.din(n18121), .dout(n18122));
  jand g17823(.dina(n18122), .dinb(n18119), .dout(n18123));
  jand g17824(.dina(n18123), .dinb(n18114), .dout(n18124));
  jor  g17825(.dina(n18124), .dinb(n18113), .dout(n18125));
  jand g17826(.dina(n18125), .dinb(asqrt[44] ), .dout(n18126));
  jor  g17827(.dina(n18113), .dinb(asqrt[44] ), .dout(n18127));
  jor  g17828(.dina(n18127), .dinb(n18124), .dout(n18128));
  jnot g17829(.din(n17505), .dout(n18129));
  jnot g17830(.din(n17507), .dout(n18130));
  jand g17831(.dina(asqrt[6] ), .dinb(n17501), .dout(n18131));
  jand g17832(.dina(n18131), .dinb(n18130), .dout(n18132));
  jor  g17833(.dina(n18132), .dinb(n18129), .dout(n18133));
  jnot g17834(.din(n17508), .dout(n18134));
  jand g17835(.dina(n18131), .dinb(n18134), .dout(n18135));
  jnot g17836(.din(n18135), .dout(n18136));
  jand g17837(.dina(n18136), .dinb(n18133), .dout(n18137));
  jand g17838(.dina(n18137), .dinb(n18128), .dout(n18138));
  jor  g17839(.dina(n18138), .dinb(n18126), .dout(n18139));
  jand g17840(.dina(n18139), .dinb(asqrt[45] ), .dout(n18140));
  jxor g17841(.dina(n17509), .dinb(n2420), .dout(n18141));
  jand g17842(.dina(n18141), .dinb(asqrt[6] ), .dout(n18142));
  jxor g17843(.dina(n18142), .dinb(n17519), .dout(n18143));
  jnot g17844(.din(n18143), .dout(n18144));
  jor  g17845(.dina(n18139), .dinb(asqrt[45] ), .dout(n18145));
  jand g17846(.dina(n18145), .dinb(n18144), .dout(n18146));
  jor  g17847(.dina(n18146), .dinb(n18140), .dout(n18147));
  jand g17848(.dina(n18147), .dinb(asqrt[46] ), .dout(n18148));
  jnot g17849(.din(n17524), .dout(n18149));
  jand g17850(.dina(n18149), .dinb(n17522), .dout(n18150));
  jand g17851(.dina(n18150), .dinb(asqrt[6] ), .dout(n18151));
  jxor g17852(.dina(n18151), .dinb(n17532), .dout(n18152));
  jnot g17853(.din(n18152), .dout(n18153));
  jor  g17854(.dina(n18140), .dinb(asqrt[46] ), .dout(n18154));
  jor  g17855(.dina(n18154), .dinb(n18146), .dout(n18155));
  jand g17856(.dina(n18155), .dinb(n18153), .dout(n18156));
  jor  g17857(.dina(n18156), .dinb(n18148), .dout(n18157));
  jand g17858(.dina(n18157), .dinb(asqrt[47] ), .dout(n18158));
  jor  g17859(.dina(n18157), .dinb(asqrt[47] ), .dout(n18159));
  jnot g17860(.din(n17538), .dout(n18160));
  jnot g17861(.din(n17539), .dout(n18161));
  jand g17862(.dina(asqrt[6] ), .dinb(n17535), .dout(n18162));
  jand g17863(.dina(n18162), .dinb(n18161), .dout(n18163));
  jor  g17864(.dina(n18163), .dinb(n18160), .dout(n18164));
  jnot g17865(.din(n17540), .dout(n18165));
  jand g17866(.dina(n18162), .dinb(n18165), .dout(n18166));
  jnot g17867(.din(n18166), .dout(n18167));
  jand g17868(.dina(n18167), .dinb(n18164), .dout(n18168));
  jand g17869(.dina(n18168), .dinb(n18159), .dout(n18169));
  jor  g17870(.dina(n18169), .dinb(n18158), .dout(n18170));
  jand g17871(.dina(n18170), .dinb(asqrt[48] ), .dout(n18171));
  jor  g17872(.dina(n18158), .dinb(asqrt[48] ), .dout(n18172));
  jor  g17873(.dina(n18172), .dinb(n18169), .dout(n18173));
  jnot g17874(.din(n17546), .dout(n18174));
  jnot g17875(.din(n17548), .dout(n18175));
  jand g17876(.dina(asqrt[6] ), .dinb(n17542), .dout(n18176));
  jand g17877(.dina(n18176), .dinb(n18175), .dout(n18177));
  jor  g17878(.dina(n18177), .dinb(n18174), .dout(n18178));
  jnot g17879(.din(n17549), .dout(n18179));
  jand g17880(.dina(n18176), .dinb(n18179), .dout(n18180));
  jnot g17881(.din(n18180), .dout(n18181));
  jand g17882(.dina(n18181), .dinb(n18178), .dout(n18182));
  jand g17883(.dina(n18182), .dinb(n18173), .dout(n18183));
  jor  g17884(.dina(n18183), .dinb(n18171), .dout(n18184));
  jand g17885(.dina(n18184), .dinb(asqrt[49] ), .dout(n18185));
  jxor g17886(.dina(n17550), .dinb(n1641), .dout(n18186));
  jand g17887(.dina(n18186), .dinb(asqrt[6] ), .dout(n18187));
  jxor g17888(.dina(n18187), .dinb(n17560), .dout(n18188));
  jnot g17889(.din(n18188), .dout(n18189));
  jor  g17890(.dina(n18184), .dinb(asqrt[49] ), .dout(n18190));
  jand g17891(.dina(n18190), .dinb(n18189), .dout(n18191));
  jor  g17892(.dina(n18191), .dinb(n18185), .dout(n18192));
  jand g17893(.dina(n18192), .dinb(asqrt[50] ), .dout(n18193));
  jnot g17894(.din(n17565), .dout(n18194));
  jand g17895(.dina(n18194), .dinb(n17563), .dout(n18195));
  jand g17896(.dina(n18195), .dinb(asqrt[6] ), .dout(n18196));
  jxor g17897(.dina(n18196), .dinb(n17573), .dout(n18197));
  jnot g17898(.din(n18197), .dout(n18198));
  jor  g17899(.dina(n18185), .dinb(asqrt[50] ), .dout(n18199));
  jor  g17900(.dina(n18199), .dinb(n18191), .dout(n18200));
  jand g17901(.dina(n18200), .dinb(n18198), .dout(n18201));
  jor  g17902(.dina(n18201), .dinb(n18193), .dout(n18202));
  jand g17903(.dina(n18202), .dinb(asqrt[51] ), .dout(n18203));
  jor  g17904(.dina(n18202), .dinb(asqrt[51] ), .dout(n18204));
  jnot g17905(.din(n17579), .dout(n18205));
  jnot g17906(.din(n17580), .dout(n18206));
  jand g17907(.dina(asqrt[6] ), .dinb(n17576), .dout(n18207));
  jand g17908(.dina(n18207), .dinb(n18206), .dout(n18208));
  jor  g17909(.dina(n18208), .dinb(n18205), .dout(n18209));
  jnot g17910(.din(n17581), .dout(n18210));
  jand g17911(.dina(n18207), .dinb(n18210), .dout(n18211));
  jnot g17912(.din(n18211), .dout(n18212));
  jand g17913(.dina(n18212), .dinb(n18209), .dout(n18213));
  jand g17914(.dina(n18213), .dinb(n18204), .dout(n18214));
  jor  g17915(.dina(n18214), .dinb(n18203), .dout(n18215));
  jand g17916(.dina(n18215), .dinb(asqrt[52] ), .dout(n18216));
  jor  g17917(.dina(n18203), .dinb(asqrt[52] ), .dout(n18217));
  jor  g17918(.dina(n18217), .dinb(n18214), .dout(n18218));
  jnot g17919(.din(n17587), .dout(n18219));
  jnot g17920(.din(n17589), .dout(n18220));
  jand g17921(.dina(asqrt[6] ), .dinb(n17583), .dout(n18221));
  jand g17922(.dina(n18221), .dinb(n18220), .dout(n18222));
  jor  g17923(.dina(n18222), .dinb(n18219), .dout(n18223));
  jnot g17924(.din(n17590), .dout(n18224));
  jand g17925(.dina(n18221), .dinb(n18224), .dout(n18225));
  jnot g17926(.din(n18225), .dout(n18226));
  jand g17927(.dina(n18226), .dinb(n18223), .dout(n18227));
  jand g17928(.dina(n18227), .dinb(n18218), .dout(n18228));
  jor  g17929(.dina(n18228), .dinb(n18216), .dout(n18229));
  jand g17930(.dina(n18229), .dinb(asqrt[53] ), .dout(n18230));
  jxor g17931(.dina(n17591), .dinb(n1034), .dout(n18231));
  jand g17932(.dina(n18231), .dinb(asqrt[6] ), .dout(n18232));
  jxor g17933(.dina(n18232), .dinb(n17601), .dout(n18233));
  jnot g17934(.din(n18233), .dout(n18234));
  jor  g17935(.dina(n18229), .dinb(asqrt[53] ), .dout(n18235));
  jand g17936(.dina(n18235), .dinb(n18234), .dout(n18236));
  jor  g17937(.dina(n18236), .dinb(n18230), .dout(n18237));
  jand g17938(.dina(n18237), .dinb(asqrt[54] ), .dout(n18238));
  jnot g17939(.din(n17606), .dout(n18239));
  jand g17940(.dina(n18239), .dinb(n17604), .dout(n18240));
  jand g17941(.dina(n18240), .dinb(asqrt[6] ), .dout(n18241));
  jxor g17942(.dina(n18241), .dinb(n17614), .dout(n18242));
  jnot g17943(.din(n18242), .dout(n18243));
  jor  g17944(.dina(n18230), .dinb(asqrt[54] ), .dout(n18244));
  jor  g17945(.dina(n18244), .dinb(n18236), .dout(n18245));
  jand g17946(.dina(n18245), .dinb(n18243), .dout(n18246));
  jor  g17947(.dina(n18246), .dinb(n18238), .dout(n18247));
  jand g17948(.dina(n18247), .dinb(asqrt[55] ), .dout(n18248));
  jor  g17949(.dina(n18247), .dinb(asqrt[55] ), .dout(n18249));
  jnot g17950(.din(n17620), .dout(n18250));
  jnot g17951(.din(n17621), .dout(n18251));
  jand g17952(.dina(asqrt[6] ), .dinb(n17617), .dout(n18252));
  jand g17953(.dina(n18252), .dinb(n18251), .dout(n18253));
  jor  g17954(.dina(n18253), .dinb(n18250), .dout(n18254));
  jnot g17955(.din(n17622), .dout(n18255));
  jand g17956(.dina(n18252), .dinb(n18255), .dout(n18256));
  jnot g17957(.din(n18256), .dout(n18257));
  jand g17958(.dina(n18257), .dinb(n18254), .dout(n18258));
  jand g17959(.dina(n18258), .dinb(n18249), .dout(n18259));
  jor  g17960(.dina(n18259), .dinb(n18248), .dout(n18260));
  jand g17961(.dina(n18260), .dinb(asqrt[56] ), .dout(n18261));
  jnot g17962(.din(n17626), .dout(n18262));
  jand g17963(.dina(n18262), .dinb(n17624), .dout(n18263));
  jand g17964(.dina(n18263), .dinb(asqrt[6] ), .dout(n18264));
  jxor g17965(.dina(n18264), .dinb(n17634), .dout(n18265));
  jnot g17966(.din(n18265), .dout(n18266));
  jor  g17967(.dina(n18248), .dinb(asqrt[56] ), .dout(n18267));
  jor  g17968(.dina(n18267), .dinb(n18259), .dout(n18268));
  jand g17969(.dina(n18268), .dinb(n18266), .dout(n18269));
  jor  g17970(.dina(n18269), .dinb(n18261), .dout(n18270));
  jand g17971(.dina(n18270), .dinb(asqrt[57] ), .dout(n18271));
  jnot g17972(.din(n17720), .dout(n18272));
  jor  g17973(.dina(n18270), .dinb(asqrt[57] ), .dout(n18273));
  jand g17974(.dina(n18273), .dinb(n18272), .dout(n18274));
  jor  g17975(.dina(n18274), .dinb(n18271), .dout(n18275));
  jand g17976(.dina(n18275), .dinb(asqrt[58] ), .dout(n18276));
  jor  g17977(.dina(n18271), .dinb(asqrt[58] ), .dout(n18277));
  jor  g17978(.dina(n18277), .dinb(n18274), .dout(n18278));
  jnot g17979(.din(n17645), .dout(n18279));
  jnot g17980(.din(n17647), .dout(n18280));
  jand g17981(.dina(asqrt[6] ), .dinb(n17641), .dout(n18281));
  jand g17982(.dina(n18281), .dinb(n18280), .dout(n18282));
  jor  g17983(.dina(n18282), .dinb(n18279), .dout(n18283));
  jnot g17984(.din(n17648), .dout(n18284));
  jand g17985(.dina(n18281), .dinb(n18284), .dout(n18285));
  jnot g17986(.din(n18285), .dout(n18286));
  jand g17987(.dina(n18286), .dinb(n18283), .dout(n18287));
  jand g17988(.dina(n18287), .dinb(n18278), .dout(n18288));
  jor  g17989(.dina(n18288), .dinb(n18276), .dout(n18289));
  jand g17990(.dina(n18289), .dinb(asqrt[59] ), .dout(n18290));
  jor  g17991(.dina(n18289), .dinb(asqrt[59] ), .dout(n18291));
  jnot g17992(.din(n17653), .dout(n18292));
  jnot g17993(.din(n17654), .dout(n18293));
  jand g17994(.dina(asqrt[6] ), .dinb(n17650), .dout(n18294));
  jand g17995(.dina(n18294), .dinb(n18293), .dout(n18295));
  jor  g17996(.dina(n18295), .dinb(n18292), .dout(n18296));
  jnot g17997(.din(n17655), .dout(n18297));
  jand g17998(.dina(n18294), .dinb(n18297), .dout(n18298));
  jnot g17999(.din(n18298), .dout(n18299));
  jand g18000(.dina(n18299), .dinb(n18296), .dout(n18300));
  jand g18001(.dina(n18300), .dinb(n18291), .dout(n18301));
  jor  g18002(.dina(n18301), .dinb(n18290), .dout(n18302));
  jand g18003(.dina(n18302), .dinb(asqrt[60] ), .dout(n18303));
  jor  g18004(.dina(n18290), .dinb(asqrt[60] ), .dout(n18304));
  jor  g18005(.dina(n18304), .dinb(n18301), .dout(n18305));
  jnot g18006(.din(n17661), .dout(n18306));
  jnot g18007(.din(n17663), .dout(n18307));
  jand g18008(.dina(asqrt[6] ), .dinb(n17657), .dout(n18308));
  jand g18009(.dina(n18308), .dinb(n18307), .dout(n18309));
  jor  g18010(.dina(n18309), .dinb(n18306), .dout(n18310));
  jnot g18011(.din(n17664), .dout(n18311));
  jand g18012(.dina(n18308), .dinb(n18311), .dout(n18312));
  jnot g18013(.din(n18312), .dout(n18313));
  jand g18014(.dina(n18313), .dinb(n18310), .dout(n18314));
  jand g18015(.dina(n18314), .dinb(n18305), .dout(n18315));
  jor  g18016(.dina(n18315), .dinb(n18303), .dout(n18316));
  jand g18017(.dina(n18316), .dinb(asqrt[61] ), .dout(n18317));
  jxor g18018(.dina(n17665), .dinb(n290), .dout(n18318));
  jand g18019(.dina(n18318), .dinb(asqrt[6] ), .dout(n18319));
  jxor g18020(.dina(n18319), .dinb(n17675), .dout(n18320));
  jnot g18021(.din(n18320), .dout(n18321));
  jor  g18022(.dina(n18316), .dinb(asqrt[61] ), .dout(n18322));
  jand g18023(.dina(n18322), .dinb(n18321), .dout(n18323));
  jor  g18024(.dina(n18323), .dinb(n18317), .dout(n18324));
  jand g18025(.dina(n18324), .dinb(asqrt[62] ), .dout(n18325));
  jnot g18026(.din(n17680), .dout(n18326));
  jand g18027(.dina(n18326), .dinb(n17678), .dout(n18327));
  jand g18028(.dina(n18327), .dinb(asqrt[6] ), .dout(n18328));
  jxor g18029(.dina(n18328), .dinb(n17688), .dout(n18329));
  jnot g18030(.din(n18329), .dout(n18330));
  jor  g18031(.dina(n18317), .dinb(asqrt[62] ), .dout(n18331));
  jor  g18032(.dina(n18331), .dinb(n18323), .dout(n18332));
  jand g18033(.dina(n18332), .dinb(n18330), .dout(n18333));
  jor  g18034(.dina(n18333), .dinb(n18325), .dout(n18334));
  jxor g18035(.dina(n17690), .dinb(n199), .dout(n18335));
  jand g18036(.dina(n18335), .dinb(asqrt[6] ), .dout(n18336));
  jxor g18037(.dina(n18336), .dinb(n17695), .dout(n18337));
  jnot g18038(.din(n17697), .dout(n18338));
  jnot g18039(.din(n17701), .dout(n18339));
  jand g18040(.dina(asqrt[6] ), .dinb(n18339), .dout(n18340));
  jand g18041(.dina(n18340), .dinb(n18338), .dout(n18341));
  jor  g18042(.dina(n18341), .dinb(n17708), .dout(n18342));
  jor  g18043(.dina(n18342), .dinb(n18337), .dout(n18343));
  jnot g18044(.din(n18343), .dout(n18344));
  jand g18045(.dina(n18344), .dinb(n18334), .dout(n18345));
  jor  g18046(.dina(n18345), .dinb(asqrt[63] ), .dout(n18346));
  jnot g18047(.din(n18337), .dout(n18347));
  jor  g18048(.dina(n18347), .dinb(n18334), .dout(n18348));
  jor  g18049(.dina(n18340), .dinb(n18338), .dout(n18349));
  jand g18050(.dina(n18339), .dinb(n18338), .dout(n18350));
  jor  g18051(.dina(n18350), .dinb(n194), .dout(n18351));
  jnot g18052(.din(n18351), .dout(n18352));
  jand g18053(.dina(n18352), .dinb(n18349), .dout(n18353));
  jnot g18054(.din(n18353), .dout(n18354));
  jand g18055(.dina(n18354), .dinb(n18348), .dout(n18355));
  jand g18056(.dina(n18355), .dinb(n18346), .dout(n18356));
  jxor g18057(.dina(n18270), .dinb(n430), .dout(n18357));
  jor  g18058(.dina(n18357), .dinb(n18356), .dout(n18358));
  jxor g18059(.dina(n18358), .dinb(n17720), .dout(n18359));
  jnot g18060(.din(asqrt[6] ), .dout(n18360));
  jor  g18061(.dina(n18356), .dinb(n17722), .dout(n18361));
  jnot g18062(.din(a[8] ), .dout(n18362));
  jnot g18063(.din(a[9] ), .dout(n18363));
  jand g18064(.dina(n17722), .dinb(n18363), .dout(n18364));
  jand g18065(.dina(n18364), .dinb(n18362), .dout(n18365));
  jnot g18066(.din(n18365), .dout(n18366));
  jand g18067(.dina(n18366), .dinb(n18361), .dout(n18367));
  jor  g18068(.dina(n18367), .dinb(n18360), .dout(n18368));
  jor  g18069(.dina(n18356), .dinb(a[10] ), .dout(n18369));
  jxor g18070(.dina(n18369), .dinb(n17723), .dout(n18370));
  jand g18071(.dina(n18367), .dinb(n18360), .dout(n18371));
  jor  g18072(.dina(n18371), .dinb(n18370), .dout(n18372));
  jand g18073(.dina(n18372), .dinb(n18368), .dout(n18373));
  jor  g18074(.dina(n18373), .dinb(n17140), .dout(n18374));
  jand g18075(.dina(n18368), .dinb(n17140), .dout(n18375));
  jand g18076(.dina(n18375), .dinb(n18372), .dout(n18376));
  jor  g18077(.dina(n18369), .dinb(a[11] ), .dout(n18377));
  jnot g18078(.din(n18356), .dout(asqrt[5] ));
  jor  g18079(.dina(asqrt[5] ), .dinb(n18360), .dout(n18379));
  jand g18080(.dina(n18379), .dinb(n18377), .dout(n18380));
  jxor g18081(.dina(n18380), .dinb(n17145), .dout(n18381));
  jor  g18082(.dina(n18381), .dinb(n18376), .dout(n18382));
  jand g18083(.dina(n18382), .dinb(n18374), .dout(n18383));
  jor  g18084(.dina(n18383), .dinb(n17135), .dout(n18384));
  jand g18085(.dina(n18383), .dinb(n17135), .dout(n18385));
  jxor g18086(.dina(n17726), .dinb(n17140), .dout(n18386));
  jor  g18087(.dina(n18386), .dinb(n18356), .dout(n18387));
  jxor g18088(.dina(n18387), .dinb(n17729), .dout(n18388));
  jor  g18089(.dina(n18388), .dinb(n18385), .dout(n18389));
  jand g18090(.dina(n18389), .dinb(n18384), .dout(n18390));
  jor  g18091(.dina(n18390), .dinb(n15955), .dout(n18391));
  jnot g18092(.din(n17735), .dout(n18392));
  jor  g18093(.dina(n18392), .dinb(n17733), .dout(n18393));
  jor  g18094(.dina(n18393), .dinb(n18356), .dout(n18394));
  jxor g18095(.dina(n18394), .dinb(n17744), .dout(n18395));
  jand g18096(.dina(n18384), .dinb(n15955), .dout(n18396));
  jand g18097(.dina(n18396), .dinb(n18389), .dout(n18397));
  jor  g18098(.dina(n18397), .dinb(n18395), .dout(n18398));
  jand g18099(.dina(n18398), .dinb(n18391), .dout(n18399));
  jor  g18100(.dina(n18399), .dinb(n15950), .dout(n18400));
  jand g18101(.dina(n18399), .dinb(n15950), .dout(n18401));
  jxor g18102(.dina(n17746), .dinb(n15955), .dout(n18402));
  jor  g18103(.dina(n18402), .dinb(n18356), .dout(n18403));
  jxor g18104(.dina(n18403), .dinb(n17751), .dout(n18404));
  jnot g18105(.din(n18404), .dout(n18405));
  jor  g18106(.dina(n18405), .dinb(n18401), .dout(n18406));
  jand g18107(.dina(n18406), .dinb(n18400), .dout(n18407));
  jor  g18108(.dina(n18407), .dinb(n14821), .dout(n18408));
  jand g18109(.dina(n18400), .dinb(n14821), .dout(n18409));
  jand g18110(.dina(n18409), .dinb(n18406), .dout(n18410));
  jnot g18111(.din(n17755), .dout(n18411));
  jand g18112(.dina(asqrt[5] ), .dinb(n18411), .dout(n18412));
  jand g18113(.dina(n18412), .dinb(n17762), .dout(n18413));
  jor  g18114(.dina(n18413), .dinb(n17760), .dout(n18414));
  jand g18115(.dina(n18412), .dinb(n17763), .dout(n18415));
  jnot g18116(.din(n18415), .dout(n18416));
  jand g18117(.dina(n18416), .dinb(n18414), .dout(n18417));
  jnot g18118(.din(n18417), .dout(n18418));
  jor  g18119(.dina(n18418), .dinb(n18410), .dout(n18419));
  jand g18120(.dina(n18419), .dinb(n18408), .dout(n18420));
  jor  g18121(.dina(n18420), .dinb(n14816), .dout(n18421));
  jand g18122(.dina(n18420), .dinb(n14816), .dout(n18422));
  jnot g18123(.din(n17770), .dout(n18423));
  jxor g18124(.dina(n17764), .dinb(n14821), .dout(n18424));
  jor  g18125(.dina(n18424), .dinb(n18356), .dout(n18425));
  jxor g18126(.dina(n18425), .dinb(n18423), .dout(n18426));
  jnot g18127(.din(n18426), .dout(n18427));
  jor  g18128(.dina(n18427), .dinb(n18422), .dout(n18428));
  jand g18129(.dina(n18428), .dinb(n18421), .dout(n18429));
  jor  g18130(.dina(n18429), .dinb(n13723), .dout(n18430));
  jnot g18131(.din(n17775), .dout(n18431));
  jor  g18132(.dina(n18431), .dinb(n17773), .dout(n18432));
  jor  g18133(.dina(n18432), .dinb(n18356), .dout(n18433));
  jxor g18134(.dina(n18433), .dinb(n17784), .dout(n18434));
  jand g18135(.dina(n18421), .dinb(n13723), .dout(n18435));
  jand g18136(.dina(n18435), .dinb(n18428), .dout(n18436));
  jor  g18137(.dina(n18436), .dinb(n18434), .dout(n18437));
  jand g18138(.dina(n18437), .dinb(n18430), .dout(n18438));
  jor  g18139(.dina(n18438), .dinb(n13718), .dout(n18439));
  jand g18140(.dina(n18438), .dinb(n13718), .dout(n18440));
  jnot g18141(.din(n17791), .dout(n18441));
  jxor g18142(.dina(n17786), .dinb(n13723), .dout(n18442));
  jor  g18143(.dina(n18442), .dinb(n18356), .dout(n18443));
  jxor g18144(.dina(n18443), .dinb(n18441), .dout(n18444));
  jnot g18145(.din(n18444), .dout(n18445));
  jor  g18146(.dina(n18445), .dinb(n18440), .dout(n18446));
  jand g18147(.dina(n18446), .dinb(n18439), .dout(n18447));
  jor  g18148(.dina(n18447), .dinb(n12675), .dout(n18448));
  jand g18149(.dina(n18439), .dinb(n12675), .dout(n18449));
  jand g18150(.dina(n18449), .dinb(n18446), .dout(n18450));
  jnot g18151(.din(n17794), .dout(n18451));
  jand g18152(.dina(asqrt[5] ), .dinb(n18451), .dout(n18452));
  jand g18153(.dina(n18452), .dinb(n17801), .dout(n18453));
  jor  g18154(.dina(n18453), .dinb(n17799), .dout(n18454));
  jand g18155(.dina(n18452), .dinb(n17802), .dout(n18455));
  jnot g18156(.din(n18455), .dout(n18456));
  jand g18157(.dina(n18456), .dinb(n18454), .dout(n18457));
  jnot g18158(.din(n18457), .dout(n18458));
  jor  g18159(.dina(n18458), .dinb(n18450), .dout(n18459));
  jand g18160(.dina(n18459), .dinb(n18448), .dout(n18460));
  jor  g18161(.dina(n18460), .dinb(n12670), .dout(n18461));
  jxor g18162(.dina(n17803), .dinb(n12675), .dout(n18462));
  jor  g18163(.dina(n18462), .dinb(n18356), .dout(n18463));
  jxor g18164(.dina(n18463), .dinb(n17808), .dout(n18464));
  jand g18165(.dina(n18460), .dinb(n12670), .dout(n18465));
  jor  g18166(.dina(n18465), .dinb(n18464), .dout(n18466));
  jand g18167(.dina(n18466), .dinb(n18461), .dout(n18467));
  jor  g18168(.dina(n18467), .dinb(n11662), .dout(n18468));
  jnot g18169(.din(n17813), .dout(n18469));
  jor  g18170(.dina(n18469), .dinb(n17811), .dout(n18470));
  jor  g18171(.dina(n18470), .dinb(n18356), .dout(n18471));
  jxor g18172(.dina(n18471), .dinb(n17822), .dout(n18472));
  jand g18173(.dina(n18461), .dinb(n11662), .dout(n18473));
  jand g18174(.dina(n18473), .dinb(n18466), .dout(n18474));
  jor  g18175(.dina(n18474), .dinb(n18472), .dout(n18475));
  jand g18176(.dina(n18475), .dinb(n18468), .dout(n18476));
  jor  g18177(.dina(n18476), .dinb(n11657), .dout(n18477));
  jand g18178(.dina(n18476), .dinb(n11657), .dout(n18478));
  jnot g18179(.din(n17825), .dout(n18479));
  jand g18180(.dina(asqrt[5] ), .dinb(n18479), .dout(n18480));
  jand g18181(.dina(n18480), .dinb(n17830), .dout(n18481));
  jor  g18182(.dina(n18481), .dinb(n17829), .dout(n18482));
  jand g18183(.dina(n18480), .dinb(n17831), .dout(n18483));
  jnot g18184(.din(n18483), .dout(n18484));
  jand g18185(.dina(n18484), .dinb(n18482), .dout(n18485));
  jnot g18186(.din(n18485), .dout(n18486));
  jor  g18187(.dina(n18486), .dinb(n18478), .dout(n18487));
  jand g18188(.dina(n18487), .dinb(n18477), .dout(n18488));
  jor  g18189(.dina(n18488), .dinb(n10701), .dout(n18489));
  jand g18190(.dina(n18477), .dinb(n10701), .dout(n18490));
  jand g18191(.dina(n18490), .dinb(n18487), .dout(n18491));
  jnot g18192(.din(n17833), .dout(n18492));
  jand g18193(.dina(asqrt[5] ), .dinb(n18492), .dout(n18493));
  jand g18194(.dina(n18493), .dinb(n17840), .dout(n18494));
  jor  g18195(.dina(n18494), .dinb(n17838), .dout(n18495));
  jand g18196(.dina(n18493), .dinb(n17841), .dout(n18496));
  jnot g18197(.din(n18496), .dout(n18497));
  jand g18198(.dina(n18497), .dinb(n18495), .dout(n18498));
  jnot g18199(.din(n18498), .dout(n18499));
  jor  g18200(.dina(n18499), .dinb(n18491), .dout(n18500));
  jand g18201(.dina(n18500), .dinb(n18489), .dout(n18501));
  jor  g18202(.dina(n18501), .dinb(n10696), .dout(n18502));
  jxor g18203(.dina(n17842), .dinb(n10701), .dout(n18503));
  jor  g18204(.dina(n18503), .dinb(n18356), .dout(n18504));
  jxor g18205(.dina(n18504), .dinb(n17853), .dout(n18505));
  jand g18206(.dina(n18501), .dinb(n10696), .dout(n18506));
  jor  g18207(.dina(n18506), .dinb(n18505), .dout(n18507));
  jand g18208(.dina(n18507), .dinb(n18502), .dout(n18508));
  jor  g18209(.dina(n18508), .dinb(n9774), .dout(n18509));
  jnot g18210(.din(n17858), .dout(n18510));
  jor  g18211(.dina(n18510), .dinb(n17856), .dout(n18511));
  jor  g18212(.dina(n18511), .dinb(n18356), .dout(n18512));
  jxor g18213(.dina(n18512), .dinb(n17867), .dout(n18513));
  jand g18214(.dina(n18502), .dinb(n9774), .dout(n18514));
  jand g18215(.dina(n18514), .dinb(n18507), .dout(n18515));
  jor  g18216(.dina(n18515), .dinb(n18513), .dout(n18516));
  jand g18217(.dina(n18516), .dinb(n18509), .dout(n18517));
  jor  g18218(.dina(n18517), .dinb(n9769), .dout(n18518));
  jand g18219(.dina(n18517), .dinb(n9769), .dout(n18519));
  jnot g18220(.din(n17870), .dout(n18520));
  jand g18221(.dina(asqrt[5] ), .dinb(n18520), .dout(n18521));
  jand g18222(.dina(n18521), .dinb(n17875), .dout(n18522));
  jor  g18223(.dina(n18522), .dinb(n17874), .dout(n18523));
  jand g18224(.dina(n18521), .dinb(n17876), .dout(n18524));
  jnot g18225(.din(n18524), .dout(n18525));
  jand g18226(.dina(n18525), .dinb(n18523), .dout(n18526));
  jnot g18227(.din(n18526), .dout(n18527));
  jor  g18228(.dina(n18527), .dinb(n18519), .dout(n18528));
  jand g18229(.dina(n18528), .dinb(n18518), .dout(n18529));
  jor  g18230(.dina(n18529), .dinb(n8898), .dout(n18530));
  jand g18231(.dina(n18518), .dinb(n8898), .dout(n18531));
  jand g18232(.dina(n18531), .dinb(n18528), .dout(n18532));
  jnot g18233(.din(n17878), .dout(n18533));
  jand g18234(.dina(asqrt[5] ), .dinb(n18533), .dout(n18534));
  jand g18235(.dina(n18534), .dinb(n17885), .dout(n18535));
  jor  g18236(.dina(n18535), .dinb(n17883), .dout(n18536));
  jand g18237(.dina(n18534), .dinb(n17886), .dout(n18537));
  jnot g18238(.din(n18537), .dout(n18538));
  jand g18239(.dina(n18538), .dinb(n18536), .dout(n18539));
  jnot g18240(.din(n18539), .dout(n18540));
  jor  g18241(.dina(n18540), .dinb(n18532), .dout(n18541));
  jand g18242(.dina(n18541), .dinb(n18530), .dout(n18542));
  jor  g18243(.dina(n18542), .dinb(n8893), .dout(n18543));
  jxor g18244(.dina(n17887), .dinb(n8898), .dout(n18544));
  jor  g18245(.dina(n18544), .dinb(n18356), .dout(n18545));
  jxor g18246(.dina(n18545), .dinb(n17898), .dout(n18546));
  jand g18247(.dina(n18542), .dinb(n8893), .dout(n18547));
  jor  g18248(.dina(n18547), .dinb(n18546), .dout(n18548));
  jand g18249(.dina(n18548), .dinb(n18543), .dout(n18549));
  jor  g18250(.dina(n18549), .dinb(n8058), .dout(n18550));
  jnot g18251(.din(n17903), .dout(n18551));
  jor  g18252(.dina(n18551), .dinb(n17901), .dout(n18552));
  jor  g18253(.dina(n18552), .dinb(n18356), .dout(n18553));
  jxor g18254(.dina(n18553), .dinb(n17912), .dout(n18554));
  jand g18255(.dina(n18543), .dinb(n8058), .dout(n18555));
  jand g18256(.dina(n18555), .dinb(n18548), .dout(n18556));
  jor  g18257(.dina(n18556), .dinb(n18554), .dout(n18557));
  jand g18258(.dina(n18557), .dinb(n18550), .dout(n18558));
  jor  g18259(.dina(n18558), .dinb(n8053), .dout(n18559));
  jand g18260(.dina(n18558), .dinb(n8053), .dout(n18560));
  jnot g18261(.din(n17915), .dout(n18561));
  jand g18262(.dina(asqrt[5] ), .dinb(n18561), .dout(n18562));
  jand g18263(.dina(n18562), .dinb(n17920), .dout(n18563));
  jor  g18264(.dina(n18563), .dinb(n17919), .dout(n18564));
  jand g18265(.dina(n18562), .dinb(n17921), .dout(n18565));
  jnot g18266(.din(n18565), .dout(n18566));
  jand g18267(.dina(n18566), .dinb(n18564), .dout(n18567));
  jnot g18268(.din(n18567), .dout(n18568));
  jor  g18269(.dina(n18568), .dinb(n18560), .dout(n18569));
  jand g18270(.dina(n18569), .dinb(n18559), .dout(n18570));
  jor  g18271(.dina(n18570), .dinb(n7265), .dout(n18571));
  jand g18272(.dina(n18559), .dinb(n7265), .dout(n18572));
  jand g18273(.dina(n18572), .dinb(n18569), .dout(n18573));
  jnot g18274(.din(n17923), .dout(n18574));
  jand g18275(.dina(asqrt[5] ), .dinb(n18574), .dout(n18575));
  jand g18276(.dina(n18575), .dinb(n17930), .dout(n18576));
  jor  g18277(.dina(n18576), .dinb(n17928), .dout(n18577));
  jand g18278(.dina(n18575), .dinb(n17931), .dout(n18578));
  jnot g18279(.din(n18578), .dout(n18579));
  jand g18280(.dina(n18579), .dinb(n18577), .dout(n18580));
  jnot g18281(.din(n18580), .dout(n18581));
  jor  g18282(.dina(n18581), .dinb(n18573), .dout(n18582));
  jand g18283(.dina(n18582), .dinb(n18571), .dout(n18583));
  jor  g18284(.dina(n18583), .dinb(n7260), .dout(n18584));
  jxor g18285(.dina(n17932), .dinb(n7265), .dout(n18585));
  jor  g18286(.dina(n18585), .dinb(n18356), .dout(n18586));
  jxor g18287(.dina(n18586), .dinb(n17943), .dout(n18587));
  jand g18288(.dina(n18583), .dinb(n7260), .dout(n18588));
  jor  g18289(.dina(n18588), .dinb(n18587), .dout(n18589));
  jand g18290(.dina(n18589), .dinb(n18584), .dout(n18590));
  jor  g18291(.dina(n18590), .dinb(n6505), .dout(n18591));
  jnot g18292(.din(n17948), .dout(n18592));
  jor  g18293(.dina(n18592), .dinb(n17946), .dout(n18593));
  jor  g18294(.dina(n18593), .dinb(n18356), .dout(n18594));
  jxor g18295(.dina(n18594), .dinb(n17957), .dout(n18595));
  jand g18296(.dina(n18584), .dinb(n6505), .dout(n18596));
  jand g18297(.dina(n18596), .dinb(n18589), .dout(n18597));
  jor  g18298(.dina(n18597), .dinb(n18595), .dout(n18598));
  jand g18299(.dina(n18598), .dinb(n18591), .dout(n18599));
  jor  g18300(.dina(n18599), .dinb(n6500), .dout(n18600));
  jand g18301(.dina(n18599), .dinb(n6500), .dout(n18601));
  jnot g18302(.din(n17960), .dout(n18602));
  jand g18303(.dina(asqrt[5] ), .dinb(n18602), .dout(n18603));
  jand g18304(.dina(n18603), .dinb(n17965), .dout(n18604));
  jor  g18305(.dina(n18604), .dinb(n17964), .dout(n18605));
  jand g18306(.dina(n18603), .dinb(n17966), .dout(n18606));
  jnot g18307(.din(n18606), .dout(n18607));
  jand g18308(.dina(n18607), .dinb(n18605), .dout(n18608));
  jnot g18309(.din(n18608), .dout(n18609));
  jor  g18310(.dina(n18609), .dinb(n18601), .dout(n18610));
  jand g18311(.dina(n18610), .dinb(n18600), .dout(n18611));
  jor  g18312(.dina(n18611), .dinb(n5793), .dout(n18612));
  jand g18313(.dina(n18600), .dinb(n5793), .dout(n18613));
  jand g18314(.dina(n18613), .dinb(n18610), .dout(n18614));
  jnot g18315(.din(n17968), .dout(n18615));
  jand g18316(.dina(asqrt[5] ), .dinb(n18615), .dout(n18616));
  jand g18317(.dina(n18616), .dinb(n17975), .dout(n18617));
  jor  g18318(.dina(n18617), .dinb(n17973), .dout(n18618));
  jand g18319(.dina(n18616), .dinb(n17976), .dout(n18619));
  jnot g18320(.din(n18619), .dout(n18620));
  jand g18321(.dina(n18620), .dinb(n18618), .dout(n18621));
  jnot g18322(.din(n18621), .dout(n18622));
  jor  g18323(.dina(n18622), .dinb(n18614), .dout(n18623));
  jand g18324(.dina(n18623), .dinb(n18612), .dout(n18624));
  jor  g18325(.dina(n18624), .dinb(n5788), .dout(n18625));
  jxor g18326(.dina(n17977), .dinb(n5793), .dout(n18626));
  jor  g18327(.dina(n18626), .dinb(n18356), .dout(n18627));
  jxor g18328(.dina(n18627), .dinb(n17988), .dout(n18628));
  jand g18329(.dina(n18624), .dinb(n5788), .dout(n18629));
  jor  g18330(.dina(n18629), .dinb(n18628), .dout(n18630));
  jand g18331(.dina(n18630), .dinb(n18625), .dout(n18631));
  jor  g18332(.dina(n18631), .dinb(n5121), .dout(n18632));
  jnot g18333(.din(n17993), .dout(n18633));
  jor  g18334(.dina(n18633), .dinb(n17991), .dout(n18634));
  jor  g18335(.dina(n18634), .dinb(n18356), .dout(n18635));
  jxor g18336(.dina(n18635), .dinb(n18002), .dout(n18636));
  jand g18337(.dina(n18625), .dinb(n5121), .dout(n18637));
  jand g18338(.dina(n18637), .dinb(n18630), .dout(n18638));
  jor  g18339(.dina(n18638), .dinb(n18636), .dout(n18639));
  jand g18340(.dina(n18639), .dinb(n18632), .dout(n18640));
  jor  g18341(.dina(n18640), .dinb(n5116), .dout(n18641));
  jand g18342(.dina(n18640), .dinb(n5116), .dout(n18642));
  jnot g18343(.din(n18005), .dout(n18643));
  jand g18344(.dina(asqrt[5] ), .dinb(n18643), .dout(n18644));
  jand g18345(.dina(n18644), .dinb(n18010), .dout(n18645));
  jor  g18346(.dina(n18645), .dinb(n18009), .dout(n18646));
  jand g18347(.dina(n18644), .dinb(n18011), .dout(n18647));
  jnot g18348(.din(n18647), .dout(n18648));
  jand g18349(.dina(n18648), .dinb(n18646), .dout(n18649));
  jnot g18350(.din(n18649), .dout(n18650));
  jor  g18351(.dina(n18650), .dinb(n18642), .dout(n18651));
  jand g18352(.dina(n18651), .dinb(n18641), .dout(n18652));
  jor  g18353(.dina(n18652), .dinb(n4499), .dout(n18653));
  jand g18354(.dina(n18641), .dinb(n4499), .dout(n18654));
  jand g18355(.dina(n18654), .dinb(n18651), .dout(n18655));
  jnot g18356(.din(n18013), .dout(n18656));
  jand g18357(.dina(asqrt[5] ), .dinb(n18656), .dout(n18657));
  jand g18358(.dina(n18657), .dinb(n18020), .dout(n18658));
  jor  g18359(.dina(n18658), .dinb(n18018), .dout(n18659));
  jand g18360(.dina(n18657), .dinb(n18021), .dout(n18660));
  jnot g18361(.din(n18660), .dout(n18661));
  jand g18362(.dina(n18661), .dinb(n18659), .dout(n18662));
  jnot g18363(.din(n18662), .dout(n18663));
  jor  g18364(.dina(n18663), .dinb(n18655), .dout(n18664));
  jand g18365(.dina(n18664), .dinb(n18653), .dout(n18665));
  jor  g18366(.dina(n18665), .dinb(n4494), .dout(n18666));
  jxor g18367(.dina(n18022), .dinb(n4499), .dout(n18667));
  jor  g18368(.dina(n18667), .dinb(n18356), .dout(n18668));
  jxor g18369(.dina(n18668), .dinb(n18033), .dout(n18669));
  jand g18370(.dina(n18665), .dinb(n4494), .dout(n18670));
  jor  g18371(.dina(n18670), .dinb(n18669), .dout(n18671));
  jand g18372(.dina(n18671), .dinb(n18666), .dout(n18672));
  jor  g18373(.dina(n18672), .dinb(n3912), .dout(n18673));
  jnot g18374(.din(n18038), .dout(n18674));
  jor  g18375(.dina(n18674), .dinb(n18036), .dout(n18675));
  jor  g18376(.dina(n18675), .dinb(n18356), .dout(n18676));
  jxor g18377(.dina(n18676), .dinb(n18047), .dout(n18677));
  jand g18378(.dina(n18666), .dinb(n3912), .dout(n18678));
  jand g18379(.dina(n18678), .dinb(n18671), .dout(n18679));
  jor  g18380(.dina(n18679), .dinb(n18677), .dout(n18680));
  jand g18381(.dina(n18680), .dinb(n18673), .dout(n18681));
  jor  g18382(.dina(n18681), .dinb(n3907), .dout(n18682));
  jand g18383(.dina(n18681), .dinb(n3907), .dout(n18683));
  jnot g18384(.din(n18050), .dout(n18684));
  jand g18385(.dina(asqrt[5] ), .dinb(n18684), .dout(n18685));
  jand g18386(.dina(n18685), .dinb(n18055), .dout(n18686));
  jor  g18387(.dina(n18686), .dinb(n18054), .dout(n18687));
  jand g18388(.dina(n18685), .dinb(n18056), .dout(n18688));
  jnot g18389(.din(n18688), .dout(n18689));
  jand g18390(.dina(n18689), .dinb(n18687), .dout(n18690));
  jnot g18391(.din(n18690), .dout(n18691));
  jor  g18392(.dina(n18691), .dinb(n18683), .dout(n18692));
  jand g18393(.dina(n18692), .dinb(n18682), .dout(n18693));
  jor  g18394(.dina(n18693), .dinb(n3376), .dout(n18694));
  jand g18395(.dina(n18682), .dinb(n3376), .dout(n18695));
  jand g18396(.dina(n18695), .dinb(n18692), .dout(n18696));
  jnot g18397(.din(n18058), .dout(n18697));
  jand g18398(.dina(asqrt[5] ), .dinb(n18697), .dout(n18698));
  jand g18399(.dina(n18698), .dinb(n18065), .dout(n18699));
  jor  g18400(.dina(n18699), .dinb(n18063), .dout(n18700));
  jand g18401(.dina(n18698), .dinb(n18066), .dout(n18701));
  jnot g18402(.din(n18701), .dout(n18702));
  jand g18403(.dina(n18702), .dinb(n18700), .dout(n18703));
  jnot g18404(.din(n18703), .dout(n18704));
  jor  g18405(.dina(n18704), .dinb(n18696), .dout(n18705));
  jand g18406(.dina(n18705), .dinb(n18694), .dout(n18706));
  jor  g18407(.dina(n18706), .dinb(n3371), .dout(n18707));
  jxor g18408(.dina(n18067), .dinb(n3376), .dout(n18708));
  jor  g18409(.dina(n18708), .dinb(n18356), .dout(n18709));
  jxor g18410(.dina(n18709), .dinb(n18078), .dout(n18710));
  jand g18411(.dina(n18706), .dinb(n3371), .dout(n18711));
  jor  g18412(.dina(n18711), .dinb(n18710), .dout(n18712));
  jand g18413(.dina(n18712), .dinb(n18707), .dout(n18713));
  jor  g18414(.dina(n18713), .dinb(n2875), .dout(n18714));
  jnot g18415(.din(n18083), .dout(n18715));
  jor  g18416(.dina(n18715), .dinb(n18081), .dout(n18716));
  jor  g18417(.dina(n18716), .dinb(n18356), .dout(n18717));
  jxor g18418(.dina(n18717), .dinb(n18092), .dout(n18718));
  jand g18419(.dina(n18707), .dinb(n2875), .dout(n18719));
  jand g18420(.dina(n18719), .dinb(n18712), .dout(n18720));
  jor  g18421(.dina(n18720), .dinb(n18718), .dout(n18721));
  jand g18422(.dina(n18721), .dinb(n18714), .dout(n18722));
  jor  g18423(.dina(n18722), .dinb(n2870), .dout(n18723));
  jand g18424(.dina(n18722), .dinb(n2870), .dout(n18724));
  jnot g18425(.din(n18095), .dout(n18725));
  jand g18426(.dina(asqrt[5] ), .dinb(n18725), .dout(n18726));
  jand g18427(.dina(n18726), .dinb(n18100), .dout(n18727));
  jor  g18428(.dina(n18727), .dinb(n18099), .dout(n18728));
  jand g18429(.dina(n18726), .dinb(n18101), .dout(n18729));
  jnot g18430(.din(n18729), .dout(n18730));
  jand g18431(.dina(n18730), .dinb(n18728), .dout(n18731));
  jnot g18432(.din(n18731), .dout(n18732));
  jor  g18433(.dina(n18732), .dinb(n18724), .dout(n18733));
  jand g18434(.dina(n18733), .dinb(n18723), .dout(n18734));
  jor  g18435(.dina(n18734), .dinb(n2425), .dout(n18735));
  jand g18436(.dina(n18723), .dinb(n2425), .dout(n18736));
  jand g18437(.dina(n18736), .dinb(n18733), .dout(n18737));
  jnot g18438(.din(n18103), .dout(n18738));
  jand g18439(.dina(asqrt[5] ), .dinb(n18738), .dout(n18739));
  jand g18440(.dina(n18739), .dinb(n18110), .dout(n18740));
  jor  g18441(.dina(n18740), .dinb(n18108), .dout(n18741));
  jand g18442(.dina(n18739), .dinb(n18111), .dout(n18742));
  jnot g18443(.din(n18742), .dout(n18743));
  jand g18444(.dina(n18743), .dinb(n18741), .dout(n18744));
  jnot g18445(.din(n18744), .dout(n18745));
  jor  g18446(.dina(n18745), .dinb(n18737), .dout(n18746));
  jand g18447(.dina(n18746), .dinb(n18735), .dout(n18747));
  jor  g18448(.dina(n18747), .dinb(n2420), .dout(n18748));
  jxor g18449(.dina(n18112), .dinb(n2425), .dout(n18749));
  jor  g18450(.dina(n18749), .dinb(n18356), .dout(n18750));
  jxor g18451(.dina(n18750), .dinb(n18123), .dout(n18751));
  jand g18452(.dina(n18747), .dinb(n2420), .dout(n18752));
  jor  g18453(.dina(n18752), .dinb(n18751), .dout(n18753));
  jand g18454(.dina(n18753), .dinb(n18748), .dout(n18754));
  jor  g18455(.dina(n18754), .dinb(n2010), .dout(n18755));
  jnot g18456(.din(n18128), .dout(n18756));
  jor  g18457(.dina(n18756), .dinb(n18126), .dout(n18757));
  jor  g18458(.dina(n18757), .dinb(n18356), .dout(n18758));
  jxor g18459(.dina(n18758), .dinb(n18137), .dout(n18759));
  jand g18460(.dina(n18748), .dinb(n2010), .dout(n18760));
  jand g18461(.dina(n18760), .dinb(n18753), .dout(n18761));
  jor  g18462(.dina(n18761), .dinb(n18759), .dout(n18762));
  jand g18463(.dina(n18762), .dinb(n18755), .dout(n18763));
  jor  g18464(.dina(n18763), .dinb(n2005), .dout(n18764));
  jand g18465(.dina(n18763), .dinb(n2005), .dout(n18765));
  jnot g18466(.din(n18140), .dout(n18766));
  jand g18467(.dina(asqrt[5] ), .dinb(n18766), .dout(n18767));
  jand g18468(.dina(n18767), .dinb(n18145), .dout(n18768));
  jor  g18469(.dina(n18768), .dinb(n18144), .dout(n18769));
  jand g18470(.dina(n18767), .dinb(n18146), .dout(n18770));
  jnot g18471(.din(n18770), .dout(n18771));
  jand g18472(.dina(n18771), .dinb(n18769), .dout(n18772));
  jnot g18473(.din(n18772), .dout(n18773));
  jor  g18474(.dina(n18773), .dinb(n18765), .dout(n18774));
  jand g18475(.dina(n18774), .dinb(n18764), .dout(n18775));
  jor  g18476(.dina(n18775), .dinb(n1646), .dout(n18776));
  jand g18477(.dina(n18764), .dinb(n1646), .dout(n18777));
  jand g18478(.dina(n18777), .dinb(n18774), .dout(n18778));
  jnot g18479(.din(n18148), .dout(n18779));
  jand g18480(.dina(asqrt[5] ), .dinb(n18779), .dout(n18780));
  jand g18481(.dina(n18780), .dinb(n18155), .dout(n18781));
  jor  g18482(.dina(n18781), .dinb(n18153), .dout(n18782));
  jand g18483(.dina(n18780), .dinb(n18156), .dout(n18783));
  jnot g18484(.din(n18783), .dout(n18784));
  jand g18485(.dina(n18784), .dinb(n18782), .dout(n18785));
  jnot g18486(.din(n18785), .dout(n18786));
  jor  g18487(.dina(n18786), .dinb(n18778), .dout(n18787));
  jand g18488(.dina(n18787), .dinb(n18776), .dout(n18788));
  jor  g18489(.dina(n18788), .dinb(n1641), .dout(n18789));
  jxor g18490(.dina(n18157), .dinb(n1646), .dout(n18790));
  jor  g18491(.dina(n18790), .dinb(n18356), .dout(n18791));
  jxor g18492(.dina(n18791), .dinb(n18168), .dout(n18792));
  jand g18493(.dina(n18788), .dinb(n1641), .dout(n18793));
  jor  g18494(.dina(n18793), .dinb(n18792), .dout(n18794));
  jand g18495(.dina(n18794), .dinb(n18789), .dout(n18795));
  jor  g18496(.dina(n18795), .dinb(n1317), .dout(n18796));
  jnot g18497(.din(n18173), .dout(n18797));
  jor  g18498(.dina(n18797), .dinb(n18171), .dout(n18798));
  jor  g18499(.dina(n18798), .dinb(n18356), .dout(n18799));
  jxor g18500(.dina(n18799), .dinb(n18182), .dout(n18800));
  jand g18501(.dina(n18789), .dinb(n1317), .dout(n18801));
  jand g18502(.dina(n18801), .dinb(n18794), .dout(n18802));
  jor  g18503(.dina(n18802), .dinb(n18800), .dout(n18803));
  jand g18504(.dina(n18803), .dinb(n18796), .dout(n18804));
  jor  g18505(.dina(n18804), .dinb(n1312), .dout(n18805));
  jand g18506(.dina(n18804), .dinb(n1312), .dout(n18806));
  jnot g18507(.din(n18185), .dout(n18807));
  jand g18508(.dina(asqrt[5] ), .dinb(n18807), .dout(n18808));
  jand g18509(.dina(n18808), .dinb(n18190), .dout(n18809));
  jor  g18510(.dina(n18809), .dinb(n18189), .dout(n18810));
  jand g18511(.dina(n18808), .dinb(n18191), .dout(n18811));
  jnot g18512(.din(n18811), .dout(n18812));
  jand g18513(.dina(n18812), .dinb(n18810), .dout(n18813));
  jnot g18514(.din(n18813), .dout(n18814));
  jor  g18515(.dina(n18814), .dinb(n18806), .dout(n18815));
  jand g18516(.dina(n18815), .dinb(n18805), .dout(n18816));
  jor  g18517(.dina(n18816), .dinb(n1039), .dout(n18817));
  jand g18518(.dina(n18805), .dinb(n1039), .dout(n18818));
  jand g18519(.dina(n18818), .dinb(n18815), .dout(n18819));
  jnot g18520(.din(n18193), .dout(n18820));
  jand g18521(.dina(asqrt[5] ), .dinb(n18820), .dout(n18821));
  jand g18522(.dina(n18821), .dinb(n18200), .dout(n18822));
  jor  g18523(.dina(n18822), .dinb(n18198), .dout(n18823));
  jand g18524(.dina(n18821), .dinb(n18201), .dout(n18824));
  jnot g18525(.din(n18824), .dout(n18825));
  jand g18526(.dina(n18825), .dinb(n18823), .dout(n18826));
  jnot g18527(.din(n18826), .dout(n18827));
  jor  g18528(.dina(n18827), .dinb(n18819), .dout(n18828));
  jand g18529(.dina(n18828), .dinb(n18817), .dout(n18829));
  jor  g18530(.dina(n18829), .dinb(n1034), .dout(n18830));
  jxor g18531(.dina(n18202), .dinb(n1039), .dout(n18831));
  jor  g18532(.dina(n18831), .dinb(n18356), .dout(n18832));
  jxor g18533(.dina(n18832), .dinb(n18213), .dout(n18833));
  jand g18534(.dina(n18829), .dinb(n1034), .dout(n18834));
  jor  g18535(.dina(n18834), .dinb(n18833), .dout(n18835));
  jand g18536(.dina(n18835), .dinb(n18830), .dout(n18836));
  jor  g18537(.dina(n18836), .dinb(n796), .dout(n18837));
  jnot g18538(.din(n18218), .dout(n18838));
  jor  g18539(.dina(n18838), .dinb(n18216), .dout(n18839));
  jor  g18540(.dina(n18839), .dinb(n18356), .dout(n18840));
  jxor g18541(.dina(n18840), .dinb(n18227), .dout(n18841));
  jand g18542(.dina(n18830), .dinb(n796), .dout(n18842));
  jand g18543(.dina(n18842), .dinb(n18835), .dout(n18843));
  jor  g18544(.dina(n18843), .dinb(n18841), .dout(n18844));
  jand g18545(.dina(n18844), .dinb(n18837), .dout(n18845));
  jor  g18546(.dina(n18845), .dinb(n791), .dout(n18846));
  jand g18547(.dina(n18845), .dinb(n791), .dout(n18847));
  jnot g18548(.din(n18230), .dout(n18848));
  jand g18549(.dina(asqrt[5] ), .dinb(n18848), .dout(n18849));
  jand g18550(.dina(n18849), .dinb(n18235), .dout(n18850));
  jor  g18551(.dina(n18850), .dinb(n18234), .dout(n18851));
  jand g18552(.dina(n18849), .dinb(n18236), .dout(n18852));
  jnot g18553(.din(n18852), .dout(n18853));
  jand g18554(.dina(n18853), .dinb(n18851), .dout(n18854));
  jnot g18555(.din(n18854), .dout(n18855));
  jor  g18556(.dina(n18855), .dinb(n18847), .dout(n18856));
  jand g18557(.dina(n18856), .dinb(n18846), .dout(n18857));
  jor  g18558(.dina(n18857), .dinb(n595), .dout(n18858));
  jand g18559(.dina(n18846), .dinb(n595), .dout(n18859));
  jand g18560(.dina(n18859), .dinb(n18856), .dout(n18860));
  jnot g18561(.din(n18238), .dout(n18861));
  jand g18562(.dina(asqrt[5] ), .dinb(n18861), .dout(n18862));
  jand g18563(.dina(n18862), .dinb(n18245), .dout(n18863));
  jor  g18564(.dina(n18863), .dinb(n18243), .dout(n18864));
  jand g18565(.dina(n18862), .dinb(n18246), .dout(n18865));
  jnot g18566(.din(n18865), .dout(n18866));
  jand g18567(.dina(n18866), .dinb(n18864), .dout(n18867));
  jnot g18568(.din(n18867), .dout(n18868));
  jor  g18569(.dina(n18868), .dinb(n18860), .dout(n18869));
  jand g18570(.dina(n18869), .dinb(n18858), .dout(n18870));
  jor  g18571(.dina(n18870), .dinb(n590), .dout(n18871));
  jxor g18572(.dina(n18247), .dinb(n595), .dout(n18872));
  jor  g18573(.dina(n18872), .dinb(n18356), .dout(n18873));
  jxor g18574(.dina(n18873), .dinb(n18258), .dout(n18874));
  jand g18575(.dina(n18870), .dinb(n590), .dout(n18875));
  jor  g18576(.dina(n18875), .dinb(n18874), .dout(n18876));
  jand g18577(.dina(n18876), .dinb(n18871), .dout(n18877));
  jor  g18578(.dina(n18877), .dinb(n430), .dout(n18878));
  jand g18579(.dina(n18871), .dinb(n430), .dout(n18879));
  jand g18580(.dina(n18879), .dinb(n18876), .dout(n18880));
  jnot g18581(.din(n18261), .dout(n18881));
  jand g18582(.dina(asqrt[5] ), .dinb(n18881), .dout(n18882));
  jand g18583(.dina(n18882), .dinb(n18268), .dout(n18883));
  jor  g18584(.dina(n18883), .dinb(n18266), .dout(n18884));
  jand g18585(.dina(n18882), .dinb(n18269), .dout(n18885));
  jnot g18586(.din(n18885), .dout(n18886));
  jand g18587(.dina(n18886), .dinb(n18884), .dout(n18887));
  jnot g18588(.din(n18887), .dout(n18888));
  jor  g18589(.dina(n18888), .dinb(n18880), .dout(n18889));
  jand g18590(.dina(n18889), .dinb(n18878), .dout(n18890));
  jor  g18591(.dina(n18890), .dinb(n425), .dout(n18891));
  jnot g18592(.din(n18359), .dout(n18892));
  jand g18593(.dina(n18890), .dinb(n425), .dout(n18893));
  jor  g18594(.dina(n18893), .dinb(n18892), .dout(n18894));
  jand g18595(.dina(n18894), .dinb(n18891), .dout(n18895));
  jor  g18596(.dina(n18895), .dinb(n305), .dout(n18896));
  jnot g18597(.din(n18278), .dout(n18897));
  jor  g18598(.dina(n18897), .dinb(n18276), .dout(n18898));
  jor  g18599(.dina(n18898), .dinb(n18356), .dout(n18899));
  jxor g18600(.dina(n18899), .dinb(n18287), .dout(n18900));
  jand g18601(.dina(n18891), .dinb(n305), .dout(n18901));
  jand g18602(.dina(n18901), .dinb(n18894), .dout(n18902));
  jor  g18603(.dina(n18902), .dinb(n18900), .dout(n18903));
  jand g18604(.dina(n18903), .dinb(n18896), .dout(n18904));
  jor  g18605(.dina(n18904), .dinb(n290), .dout(n18905));
  jxor g18606(.dina(n18289), .dinb(n305), .dout(n18906));
  jor  g18607(.dina(n18906), .dinb(n18356), .dout(n18907));
  jxor g18608(.dina(n18907), .dinb(n18300), .dout(n18908));
  jand g18609(.dina(n18904), .dinb(n290), .dout(n18909));
  jor  g18610(.dina(n18909), .dinb(n18908), .dout(n18910));
  jand g18611(.dina(n18910), .dinb(n18905), .dout(n18911));
  jor  g18612(.dina(n18911), .dinb(n223), .dout(n18912));
  jnot g18613(.din(n18305), .dout(n18913));
  jor  g18614(.dina(n18913), .dinb(n18303), .dout(n18914));
  jor  g18615(.dina(n18914), .dinb(n18356), .dout(n18915));
  jxor g18616(.dina(n18915), .dinb(n18314), .dout(n18916));
  jand g18617(.dina(n18905), .dinb(n223), .dout(n18917));
  jand g18618(.dina(n18917), .dinb(n18910), .dout(n18918));
  jor  g18619(.dina(n18918), .dinb(n18916), .dout(n18919));
  jand g18620(.dina(n18919), .dinb(n18912), .dout(n18920));
  jor  g18621(.dina(n18920), .dinb(n199), .dout(n18921));
  jand g18622(.dina(n18920), .dinb(n199), .dout(n18922));
  jnot g18623(.din(n18317), .dout(n18923));
  jand g18624(.dina(asqrt[5] ), .dinb(n18923), .dout(n18924));
  jand g18625(.dina(n18924), .dinb(n18322), .dout(n18925));
  jor  g18626(.dina(n18925), .dinb(n18321), .dout(n18926));
  jand g18627(.dina(n18924), .dinb(n18323), .dout(n18927));
  jnot g18628(.din(n18927), .dout(n18928));
  jand g18629(.dina(n18928), .dinb(n18926), .dout(n18929));
  jnot g18630(.din(n18929), .dout(n18930));
  jor  g18631(.dina(n18930), .dinb(n18922), .dout(n18931));
  jand g18632(.dina(n18931), .dinb(n18921), .dout(n18932));
  jnot g18633(.din(n18325), .dout(n18933));
  jand g18634(.dina(asqrt[5] ), .dinb(n18933), .dout(n18934));
  jand g18635(.dina(n18934), .dinb(n18332), .dout(n18935));
  jor  g18636(.dina(n18935), .dinb(n18330), .dout(n18936));
  jand g18637(.dina(n18934), .dinb(n18333), .dout(n18937));
  jnot g18638(.din(n18937), .dout(n18938));
  jand g18639(.dina(n18938), .dinb(n18936), .dout(n18939));
  jnot g18640(.din(n18939), .dout(n18940));
  jnot g18641(.din(n18348), .dout(n18941));
  jand g18642(.dina(asqrt[5] ), .dinb(n18347), .dout(n18942));
  jand g18643(.dina(n18942), .dinb(n18334), .dout(n18943));
  jor  g18644(.dina(n18943), .dinb(n18941), .dout(n18944));
  jor  g18645(.dina(n18944), .dinb(n18940), .dout(n18945));
  jor  g18646(.dina(n18945), .dinb(n18932), .dout(n18946));
  jand g18647(.dina(n18946), .dinb(n194), .dout(n18947));
  jand g18648(.dina(n18940), .dinb(n18932), .dout(n18948));
  jor  g18649(.dina(n18942), .dinb(n18334), .dout(n18949));
  jand g18650(.dina(n18347), .dinb(n18334), .dout(n18950));
  jor  g18651(.dina(n18950), .dinb(n194), .dout(n18951));
  jnot g18652(.din(n18951), .dout(n18952));
  jand g18653(.dina(n18952), .dinb(n18949), .dout(n18953));
  jor  g18654(.dina(n18953), .dinb(n18948), .dout(n18954));
  jor  g18655(.dina(n18954), .dinb(n18947), .dout(asqrt[4] ));
  jxor g18656(.dina(n18890), .dinb(n425), .dout(n18956));
  jand g18657(.dina(n18956), .dinb(asqrt[4] ), .dout(n18957));
  jxor g18658(.dina(n18957), .dinb(n18359), .dout(n18958));
  jnot g18659(.din(n18958), .dout(n18959));
  jand g18660(.dina(asqrt[4] ), .dinb(a[8] ), .dout(n18960));
  jnot g18661(.din(a[6] ), .dout(n18961));
  jnot g18662(.din(a[7] ), .dout(n18962));
  jand g18663(.dina(n18362), .dinb(n18962), .dout(n18963));
  jand g18664(.dina(n18963), .dinb(n18961), .dout(n18964));
  jor  g18665(.dina(n18964), .dinb(n18960), .dout(n18965));
  jand g18666(.dina(n18965), .dinb(asqrt[5] ), .dout(n18966));
  jand g18667(.dina(asqrt[4] ), .dinb(n18362), .dout(n18967));
  jxor g18668(.dina(n18967), .dinb(n18363), .dout(n18968));
  jor  g18669(.dina(n18965), .dinb(asqrt[5] ), .dout(n18969));
  jand g18670(.dina(n18969), .dinb(n18968), .dout(n18970));
  jor  g18671(.dina(n18970), .dinb(n18966), .dout(n18971));
  jand g18672(.dina(n18971), .dinb(asqrt[6] ), .dout(n18972));
  jor  g18673(.dina(n18966), .dinb(asqrt[6] ), .dout(n18973));
  jor  g18674(.dina(n18973), .dinb(n18970), .dout(n18974));
  jand g18675(.dina(n18967), .dinb(n18363), .dout(n18975));
  jnot g18676(.din(asqrt[4] ), .dout(n18976));
  jand g18677(.dina(n18976), .dinb(asqrt[5] ), .dout(n18977));
  jor  g18678(.dina(n18977), .dinb(n18975), .dout(n18978));
  jxor g18679(.dina(n18978), .dinb(n17722), .dout(n18979));
  jand g18680(.dina(n18979), .dinb(n18974), .dout(n18980));
  jor  g18681(.dina(n18980), .dinb(n18972), .dout(n18981));
  jand g18682(.dina(n18981), .dinb(asqrt[7] ), .dout(n18982));
  jor  g18683(.dina(n18981), .dinb(asqrt[7] ), .dout(n18983));
  jxor g18684(.dina(n18367), .dinb(n18360), .dout(n18984));
  jand g18685(.dina(n18984), .dinb(asqrt[4] ), .dout(n18985));
  jxor g18686(.dina(n18985), .dinb(n18370), .dout(n18986));
  jnot g18687(.din(n18986), .dout(n18987));
  jand g18688(.dina(n18987), .dinb(n18983), .dout(n18988));
  jor  g18689(.dina(n18988), .dinb(n18982), .dout(n18989));
  jand g18690(.dina(n18989), .dinb(asqrt[8] ), .dout(n18990));
  jnot g18691(.din(n18376), .dout(n18991));
  jand g18692(.dina(n18991), .dinb(n18374), .dout(n18992));
  jand g18693(.dina(n18992), .dinb(asqrt[4] ), .dout(n18993));
  jxor g18694(.dina(n18993), .dinb(n18381), .dout(n18994));
  jnot g18695(.din(n18994), .dout(n18995));
  jor  g18696(.dina(n18982), .dinb(asqrt[8] ), .dout(n18996));
  jor  g18697(.dina(n18996), .dinb(n18988), .dout(n18997));
  jand g18698(.dina(n18997), .dinb(n18995), .dout(n18998));
  jor  g18699(.dina(n18998), .dinb(n18990), .dout(n18999));
  jand g18700(.dina(n18999), .dinb(asqrt[9] ), .dout(n19000));
  jor  g18701(.dina(n18999), .dinb(asqrt[9] ), .dout(n19001));
  jnot g18702(.din(n18388), .dout(n19002));
  jxor g18703(.dina(n18383), .dinb(n17135), .dout(n19003));
  jand g18704(.dina(n19003), .dinb(asqrt[4] ), .dout(n19004));
  jxor g18705(.dina(n19004), .dinb(n19002), .dout(n19005));
  jand g18706(.dina(n19005), .dinb(n19001), .dout(n19006));
  jor  g18707(.dina(n19006), .dinb(n19000), .dout(n19007));
  jand g18708(.dina(n19007), .dinb(asqrt[10] ), .dout(n19008));
  jor  g18709(.dina(n19000), .dinb(asqrt[10] ), .dout(n19009));
  jor  g18710(.dina(n19009), .dinb(n19006), .dout(n19010));
  jnot g18711(.din(n18395), .dout(n19011));
  jnot g18712(.din(n18397), .dout(n19012));
  jand g18713(.dina(asqrt[4] ), .dinb(n18391), .dout(n19013));
  jand g18714(.dina(n19013), .dinb(n19012), .dout(n19014));
  jor  g18715(.dina(n19014), .dinb(n19011), .dout(n19015));
  jnot g18716(.din(n18398), .dout(n19016));
  jand g18717(.dina(n19013), .dinb(n19016), .dout(n19017));
  jnot g18718(.din(n19017), .dout(n19018));
  jand g18719(.dina(n19018), .dinb(n19015), .dout(n19019));
  jand g18720(.dina(n19019), .dinb(n19010), .dout(n19020));
  jor  g18721(.dina(n19020), .dinb(n19008), .dout(n19021));
  jand g18722(.dina(n19021), .dinb(asqrt[11] ), .dout(n19022));
  jor  g18723(.dina(n19021), .dinb(asqrt[11] ), .dout(n19023));
  jxor g18724(.dina(n18399), .dinb(n15950), .dout(n19024));
  jand g18725(.dina(n19024), .dinb(asqrt[4] ), .dout(n19025));
  jxor g18726(.dina(n19025), .dinb(n18404), .dout(n19026));
  jand g18727(.dina(n19026), .dinb(n19023), .dout(n19027));
  jor  g18728(.dina(n19027), .dinb(n19022), .dout(n19028));
  jand g18729(.dina(n19028), .dinb(asqrt[12] ), .dout(n19029));
  jnot g18730(.din(n18410), .dout(n19030));
  jand g18731(.dina(n19030), .dinb(n18408), .dout(n19031));
  jand g18732(.dina(n19031), .dinb(asqrt[4] ), .dout(n19032));
  jxor g18733(.dina(n19032), .dinb(n18418), .dout(n19033));
  jnot g18734(.din(n19033), .dout(n19034));
  jor  g18735(.dina(n19022), .dinb(asqrt[12] ), .dout(n19035));
  jor  g18736(.dina(n19035), .dinb(n19027), .dout(n19036));
  jand g18737(.dina(n19036), .dinb(n19034), .dout(n19037));
  jor  g18738(.dina(n19037), .dinb(n19029), .dout(n19038));
  jand g18739(.dina(n19038), .dinb(asqrt[13] ), .dout(n19039));
  jor  g18740(.dina(n19038), .dinb(asqrt[13] ), .dout(n19040));
  jxor g18741(.dina(n18420), .dinb(n14816), .dout(n19041));
  jand g18742(.dina(n19041), .dinb(asqrt[4] ), .dout(n19042));
  jxor g18743(.dina(n19042), .dinb(n18426), .dout(n19043));
  jand g18744(.dina(n19043), .dinb(n19040), .dout(n19044));
  jor  g18745(.dina(n19044), .dinb(n19039), .dout(n19045));
  jand g18746(.dina(n19045), .dinb(asqrt[14] ), .dout(n19046));
  jor  g18747(.dina(n19039), .dinb(asqrt[14] ), .dout(n19047));
  jor  g18748(.dina(n19047), .dinb(n19044), .dout(n19048));
  jnot g18749(.din(n18434), .dout(n19049));
  jnot g18750(.din(n18436), .dout(n19050));
  jand g18751(.dina(asqrt[4] ), .dinb(n18430), .dout(n19051));
  jand g18752(.dina(n19051), .dinb(n19050), .dout(n19052));
  jor  g18753(.dina(n19052), .dinb(n19049), .dout(n19053));
  jnot g18754(.din(n18437), .dout(n19054));
  jand g18755(.dina(n19051), .dinb(n19054), .dout(n19055));
  jnot g18756(.din(n19055), .dout(n19056));
  jand g18757(.dina(n19056), .dinb(n19053), .dout(n19057));
  jand g18758(.dina(n19057), .dinb(n19048), .dout(n19058));
  jor  g18759(.dina(n19058), .dinb(n19046), .dout(n19059));
  jand g18760(.dina(n19059), .dinb(asqrt[15] ), .dout(n19060));
  jxor g18761(.dina(n18438), .dinb(n13718), .dout(n19061));
  jand g18762(.dina(n19061), .dinb(asqrt[4] ), .dout(n19062));
  jxor g18763(.dina(n19062), .dinb(n18445), .dout(n19063));
  jnot g18764(.din(n19063), .dout(n19064));
  jor  g18765(.dina(n19059), .dinb(asqrt[15] ), .dout(n19065));
  jand g18766(.dina(n19065), .dinb(n19064), .dout(n19066));
  jor  g18767(.dina(n19066), .dinb(n19060), .dout(n19067));
  jand g18768(.dina(n19067), .dinb(asqrt[16] ), .dout(n19068));
  jnot g18769(.din(n18450), .dout(n19069));
  jand g18770(.dina(n19069), .dinb(n18448), .dout(n19070));
  jand g18771(.dina(n19070), .dinb(asqrt[4] ), .dout(n19071));
  jxor g18772(.dina(n19071), .dinb(n18458), .dout(n19072));
  jnot g18773(.din(n19072), .dout(n19073));
  jor  g18774(.dina(n19060), .dinb(asqrt[16] ), .dout(n19074));
  jor  g18775(.dina(n19074), .dinb(n19066), .dout(n19075));
  jand g18776(.dina(n19075), .dinb(n19073), .dout(n19076));
  jor  g18777(.dina(n19076), .dinb(n19068), .dout(n19077));
  jand g18778(.dina(n19077), .dinb(asqrt[17] ), .dout(n19078));
  jor  g18779(.dina(n19077), .dinb(asqrt[17] ), .dout(n19079));
  jnot g18780(.din(n18464), .dout(n19080));
  jnot g18781(.din(n18465), .dout(n19081));
  jand g18782(.dina(asqrt[4] ), .dinb(n18461), .dout(n19082));
  jand g18783(.dina(n19082), .dinb(n19081), .dout(n19083));
  jor  g18784(.dina(n19083), .dinb(n19080), .dout(n19084));
  jnot g18785(.din(n18466), .dout(n19085));
  jand g18786(.dina(n19082), .dinb(n19085), .dout(n19086));
  jnot g18787(.din(n19086), .dout(n19087));
  jand g18788(.dina(n19087), .dinb(n19084), .dout(n19088));
  jand g18789(.dina(n19088), .dinb(n19079), .dout(n19089));
  jor  g18790(.dina(n19089), .dinb(n19078), .dout(n19090));
  jand g18791(.dina(n19090), .dinb(asqrt[18] ), .dout(n19091));
  jor  g18792(.dina(n19078), .dinb(asqrt[18] ), .dout(n19092));
  jor  g18793(.dina(n19092), .dinb(n19089), .dout(n19093));
  jnot g18794(.din(n18472), .dout(n19094));
  jnot g18795(.din(n18474), .dout(n19095));
  jand g18796(.dina(asqrt[4] ), .dinb(n18468), .dout(n19096));
  jand g18797(.dina(n19096), .dinb(n19095), .dout(n19097));
  jor  g18798(.dina(n19097), .dinb(n19094), .dout(n19098));
  jnot g18799(.din(n18475), .dout(n19099));
  jand g18800(.dina(n19096), .dinb(n19099), .dout(n19100));
  jnot g18801(.din(n19100), .dout(n19101));
  jand g18802(.dina(n19101), .dinb(n19098), .dout(n19102));
  jand g18803(.dina(n19102), .dinb(n19093), .dout(n19103));
  jor  g18804(.dina(n19103), .dinb(n19091), .dout(n19104));
  jand g18805(.dina(n19104), .dinb(asqrt[19] ), .dout(n19105));
  jxor g18806(.dina(n18476), .dinb(n11657), .dout(n19106));
  jand g18807(.dina(n19106), .dinb(asqrt[4] ), .dout(n19107));
  jxor g18808(.dina(n19107), .dinb(n18486), .dout(n19108));
  jnot g18809(.din(n19108), .dout(n19109));
  jor  g18810(.dina(n19104), .dinb(asqrt[19] ), .dout(n19110));
  jand g18811(.dina(n19110), .dinb(n19109), .dout(n19111));
  jor  g18812(.dina(n19111), .dinb(n19105), .dout(n19112));
  jand g18813(.dina(n19112), .dinb(asqrt[20] ), .dout(n19113));
  jnot g18814(.din(n18491), .dout(n19114));
  jand g18815(.dina(n19114), .dinb(n18489), .dout(n19115));
  jand g18816(.dina(n19115), .dinb(asqrt[4] ), .dout(n19116));
  jxor g18817(.dina(n19116), .dinb(n18499), .dout(n19117));
  jnot g18818(.din(n19117), .dout(n19118));
  jor  g18819(.dina(n19105), .dinb(asqrt[20] ), .dout(n19119));
  jor  g18820(.dina(n19119), .dinb(n19111), .dout(n19120));
  jand g18821(.dina(n19120), .dinb(n19118), .dout(n19121));
  jor  g18822(.dina(n19121), .dinb(n19113), .dout(n19122));
  jand g18823(.dina(n19122), .dinb(asqrt[21] ), .dout(n19123));
  jor  g18824(.dina(n19122), .dinb(asqrt[21] ), .dout(n19124));
  jnot g18825(.din(n18505), .dout(n19125));
  jnot g18826(.din(n18506), .dout(n19126));
  jand g18827(.dina(asqrt[4] ), .dinb(n18502), .dout(n19127));
  jand g18828(.dina(n19127), .dinb(n19126), .dout(n19128));
  jor  g18829(.dina(n19128), .dinb(n19125), .dout(n19129));
  jnot g18830(.din(n18507), .dout(n19130));
  jand g18831(.dina(n19127), .dinb(n19130), .dout(n19131));
  jnot g18832(.din(n19131), .dout(n19132));
  jand g18833(.dina(n19132), .dinb(n19129), .dout(n19133));
  jand g18834(.dina(n19133), .dinb(n19124), .dout(n19134));
  jor  g18835(.dina(n19134), .dinb(n19123), .dout(n19135));
  jand g18836(.dina(n19135), .dinb(asqrt[22] ), .dout(n19136));
  jor  g18837(.dina(n19123), .dinb(asqrt[22] ), .dout(n19137));
  jor  g18838(.dina(n19137), .dinb(n19134), .dout(n19138));
  jnot g18839(.din(n18513), .dout(n19139));
  jnot g18840(.din(n18515), .dout(n19140));
  jand g18841(.dina(asqrt[4] ), .dinb(n18509), .dout(n19141));
  jand g18842(.dina(n19141), .dinb(n19140), .dout(n19142));
  jor  g18843(.dina(n19142), .dinb(n19139), .dout(n19143));
  jnot g18844(.din(n18516), .dout(n19144));
  jand g18845(.dina(n19141), .dinb(n19144), .dout(n19145));
  jnot g18846(.din(n19145), .dout(n19146));
  jand g18847(.dina(n19146), .dinb(n19143), .dout(n19147));
  jand g18848(.dina(n19147), .dinb(n19138), .dout(n19148));
  jor  g18849(.dina(n19148), .dinb(n19136), .dout(n19149));
  jand g18850(.dina(n19149), .dinb(asqrt[23] ), .dout(n19150));
  jxor g18851(.dina(n18517), .dinb(n9769), .dout(n19151));
  jand g18852(.dina(n19151), .dinb(asqrt[4] ), .dout(n19152));
  jxor g18853(.dina(n19152), .dinb(n18527), .dout(n19153));
  jnot g18854(.din(n19153), .dout(n19154));
  jor  g18855(.dina(n19149), .dinb(asqrt[23] ), .dout(n19155));
  jand g18856(.dina(n19155), .dinb(n19154), .dout(n19156));
  jor  g18857(.dina(n19156), .dinb(n19150), .dout(n19157));
  jand g18858(.dina(n19157), .dinb(asqrt[24] ), .dout(n19158));
  jnot g18859(.din(n18532), .dout(n19159));
  jand g18860(.dina(n19159), .dinb(n18530), .dout(n19160));
  jand g18861(.dina(n19160), .dinb(asqrt[4] ), .dout(n19161));
  jxor g18862(.dina(n19161), .dinb(n18540), .dout(n19162));
  jnot g18863(.din(n19162), .dout(n19163));
  jor  g18864(.dina(n19150), .dinb(asqrt[24] ), .dout(n19164));
  jor  g18865(.dina(n19164), .dinb(n19156), .dout(n19165));
  jand g18866(.dina(n19165), .dinb(n19163), .dout(n19166));
  jor  g18867(.dina(n19166), .dinb(n19158), .dout(n19167));
  jand g18868(.dina(n19167), .dinb(asqrt[25] ), .dout(n19168));
  jor  g18869(.dina(n19167), .dinb(asqrt[25] ), .dout(n19169));
  jnot g18870(.din(n18546), .dout(n19170));
  jnot g18871(.din(n18547), .dout(n19171));
  jand g18872(.dina(asqrt[4] ), .dinb(n18543), .dout(n19172));
  jand g18873(.dina(n19172), .dinb(n19171), .dout(n19173));
  jor  g18874(.dina(n19173), .dinb(n19170), .dout(n19174));
  jnot g18875(.din(n18548), .dout(n19175));
  jand g18876(.dina(n19172), .dinb(n19175), .dout(n19176));
  jnot g18877(.din(n19176), .dout(n19177));
  jand g18878(.dina(n19177), .dinb(n19174), .dout(n19178));
  jand g18879(.dina(n19178), .dinb(n19169), .dout(n19179));
  jor  g18880(.dina(n19179), .dinb(n19168), .dout(n19180));
  jand g18881(.dina(n19180), .dinb(asqrt[26] ), .dout(n19181));
  jor  g18882(.dina(n19168), .dinb(asqrt[26] ), .dout(n19182));
  jor  g18883(.dina(n19182), .dinb(n19179), .dout(n19183));
  jnot g18884(.din(n18554), .dout(n19184));
  jnot g18885(.din(n18556), .dout(n19185));
  jand g18886(.dina(asqrt[4] ), .dinb(n18550), .dout(n19186));
  jand g18887(.dina(n19186), .dinb(n19185), .dout(n19187));
  jor  g18888(.dina(n19187), .dinb(n19184), .dout(n19188));
  jnot g18889(.din(n18557), .dout(n19189));
  jand g18890(.dina(n19186), .dinb(n19189), .dout(n19190));
  jnot g18891(.din(n19190), .dout(n19191));
  jand g18892(.dina(n19191), .dinb(n19188), .dout(n19192));
  jand g18893(.dina(n19192), .dinb(n19183), .dout(n19193));
  jor  g18894(.dina(n19193), .dinb(n19181), .dout(n19194));
  jand g18895(.dina(n19194), .dinb(asqrt[27] ), .dout(n19195));
  jxor g18896(.dina(n18558), .dinb(n8053), .dout(n19196));
  jand g18897(.dina(n19196), .dinb(asqrt[4] ), .dout(n19197));
  jxor g18898(.dina(n19197), .dinb(n18568), .dout(n19198));
  jnot g18899(.din(n19198), .dout(n19199));
  jor  g18900(.dina(n19194), .dinb(asqrt[27] ), .dout(n19200));
  jand g18901(.dina(n19200), .dinb(n19199), .dout(n19201));
  jor  g18902(.dina(n19201), .dinb(n19195), .dout(n19202));
  jand g18903(.dina(n19202), .dinb(asqrt[28] ), .dout(n19203));
  jnot g18904(.din(n18573), .dout(n19204));
  jand g18905(.dina(n19204), .dinb(n18571), .dout(n19205));
  jand g18906(.dina(n19205), .dinb(asqrt[4] ), .dout(n19206));
  jxor g18907(.dina(n19206), .dinb(n18581), .dout(n19207));
  jnot g18908(.din(n19207), .dout(n19208));
  jor  g18909(.dina(n19195), .dinb(asqrt[28] ), .dout(n19209));
  jor  g18910(.dina(n19209), .dinb(n19201), .dout(n19210));
  jand g18911(.dina(n19210), .dinb(n19208), .dout(n19211));
  jor  g18912(.dina(n19211), .dinb(n19203), .dout(n19212));
  jand g18913(.dina(n19212), .dinb(asqrt[29] ), .dout(n19213));
  jor  g18914(.dina(n19212), .dinb(asqrt[29] ), .dout(n19214));
  jnot g18915(.din(n18587), .dout(n19215));
  jnot g18916(.din(n18588), .dout(n19216));
  jand g18917(.dina(asqrt[4] ), .dinb(n18584), .dout(n19217));
  jand g18918(.dina(n19217), .dinb(n19216), .dout(n19218));
  jor  g18919(.dina(n19218), .dinb(n19215), .dout(n19219));
  jnot g18920(.din(n18589), .dout(n19220));
  jand g18921(.dina(n19217), .dinb(n19220), .dout(n19221));
  jnot g18922(.din(n19221), .dout(n19222));
  jand g18923(.dina(n19222), .dinb(n19219), .dout(n19223));
  jand g18924(.dina(n19223), .dinb(n19214), .dout(n19224));
  jor  g18925(.dina(n19224), .dinb(n19213), .dout(n19225));
  jand g18926(.dina(n19225), .dinb(asqrt[30] ), .dout(n19226));
  jor  g18927(.dina(n19213), .dinb(asqrt[30] ), .dout(n19227));
  jor  g18928(.dina(n19227), .dinb(n19224), .dout(n19228));
  jnot g18929(.din(n18595), .dout(n19229));
  jnot g18930(.din(n18597), .dout(n19230));
  jand g18931(.dina(asqrt[4] ), .dinb(n18591), .dout(n19231));
  jand g18932(.dina(n19231), .dinb(n19230), .dout(n19232));
  jor  g18933(.dina(n19232), .dinb(n19229), .dout(n19233));
  jnot g18934(.din(n18598), .dout(n19234));
  jand g18935(.dina(n19231), .dinb(n19234), .dout(n19235));
  jnot g18936(.din(n19235), .dout(n19236));
  jand g18937(.dina(n19236), .dinb(n19233), .dout(n19237));
  jand g18938(.dina(n19237), .dinb(n19228), .dout(n19238));
  jor  g18939(.dina(n19238), .dinb(n19226), .dout(n19239));
  jand g18940(.dina(n19239), .dinb(asqrt[31] ), .dout(n19240));
  jxor g18941(.dina(n18599), .dinb(n6500), .dout(n19241));
  jand g18942(.dina(n19241), .dinb(asqrt[4] ), .dout(n19242));
  jxor g18943(.dina(n19242), .dinb(n18609), .dout(n19243));
  jnot g18944(.din(n19243), .dout(n19244));
  jor  g18945(.dina(n19239), .dinb(asqrt[31] ), .dout(n19245));
  jand g18946(.dina(n19245), .dinb(n19244), .dout(n19246));
  jor  g18947(.dina(n19246), .dinb(n19240), .dout(n19247));
  jand g18948(.dina(n19247), .dinb(asqrt[32] ), .dout(n19248));
  jnot g18949(.din(n18614), .dout(n19249));
  jand g18950(.dina(n19249), .dinb(n18612), .dout(n19250));
  jand g18951(.dina(n19250), .dinb(asqrt[4] ), .dout(n19251));
  jxor g18952(.dina(n19251), .dinb(n18622), .dout(n19252));
  jnot g18953(.din(n19252), .dout(n19253));
  jor  g18954(.dina(n19240), .dinb(asqrt[32] ), .dout(n19254));
  jor  g18955(.dina(n19254), .dinb(n19246), .dout(n19255));
  jand g18956(.dina(n19255), .dinb(n19253), .dout(n19256));
  jor  g18957(.dina(n19256), .dinb(n19248), .dout(n19257));
  jand g18958(.dina(n19257), .dinb(asqrt[33] ), .dout(n19258));
  jor  g18959(.dina(n19257), .dinb(asqrt[33] ), .dout(n19259));
  jnot g18960(.din(n18628), .dout(n19260));
  jnot g18961(.din(n18629), .dout(n19261));
  jand g18962(.dina(asqrt[4] ), .dinb(n18625), .dout(n19262));
  jand g18963(.dina(n19262), .dinb(n19261), .dout(n19263));
  jor  g18964(.dina(n19263), .dinb(n19260), .dout(n19264));
  jnot g18965(.din(n18630), .dout(n19265));
  jand g18966(.dina(n19262), .dinb(n19265), .dout(n19266));
  jnot g18967(.din(n19266), .dout(n19267));
  jand g18968(.dina(n19267), .dinb(n19264), .dout(n19268));
  jand g18969(.dina(n19268), .dinb(n19259), .dout(n19269));
  jor  g18970(.dina(n19269), .dinb(n19258), .dout(n19270));
  jand g18971(.dina(n19270), .dinb(asqrt[34] ), .dout(n19271));
  jor  g18972(.dina(n19258), .dinb(asqrt[34] ), .dout(n19272));
  jor  g18973(.dina(n19272), .dinb(n19269), .dout(n19273));
  jnot g18974(.din(n18636), .dout(n19274));
  jnot g18975(.din(n18638), .dout(n19275));
  jand g18976(.dina(asqrt[4] ), .dinb(n18632), .dout(n19276));
  jand g18977(.dina(n19276), .dinb(n19275), .dout(n19277));
  jor  g18978(.dina(n19277), .dinb(n19274), .dout(n19278));
  jnot g18979(.din(n18639), .dout(n19279));
  jand g18980(.dina(n19276), .dinb(n19279), .dout(n19280));
  jnot g18981(.din(n19280), .dout(n19281));
  jand g18982(.dina(n19281), .dinb(n19278), .dout(n19282));
  jand g18983(.dina(n19282), .dinb(n19273), .dout(n19283));
  jor  g18984(.dina(n19283), .dinb(n19271), .dout(n19284));
  jand g18985(.dina(n19284), .dinb(asqrt[35] ), .dout(n19285));
  jxor g18986(.dina(n18640), .dinb(n5116), .dout(n19286));
  jand g18987(.dina(n19286), .dinb(asqrt[4] ), .dout(n19287));
  jxor g18988(.dina(n19287), .dinb(n18650), .dout(n19288));
  jnot g18989(.din(n19288), .dout(n19289));
  jor  g18990(.dina(n19284), .dinb(asqrt[35] ), .dout(n19290));
  jand g18991(.dina(n19290), .dinb(n19289), .dout(n19291));
  jor  g18992(.dina(n19291), .dinb(n19285), .dout(n19292));
  jand g18993(.dina(n19292), .dinb(asqrt[36] ), .dout(n19293));
  jnot g18994(.din(n18655), .dout(n19294));
  jand g18995(.dina(n19294), .dinb(n18653), .dout(n19295));
  jand g18996(.dina(n19295), .dinb(asqrt[4] ), .dout(n19296));
  jxor g18997(.dina(n19296), .dinb(n18663), .dout(n19297));
  jnot g18998(.din(n19297), .dout(n19298));
  jor  g18999(.dina(n19285), .dinb(asqrt[36] ), .dout(n19299));
  jor  g19000(.dina(n19299), .dinb(n19291), .dout(n19300));
  jand g19001(.dina(n19300), .dinb(n19298), .dout(n19301));
  jor  g19002(.dina(n19301), .dinb(n19293), .dout(n19302));
  jand g19003(.dina(n19302), .dinb(asqrt[37] ), .dout(n19303));
  jor  g19004(.dina(n19302), .dinb(asqrt[37] ), .dout(n19304));
  jnot g19005(.din(n18669), .dout(n19305));
  jnot g19006(.din(n18670), .dout(n19306));
  jand g19007(.dina(asqrt[4] ), .dinb(n18666), .dout(n19307));
  jand g19008(.dina(n19307), .dinb(n19306), .dout(n19308));
  jor  g19009(.dina(n19308), .dinb(n19305), .dout(n19309));
  jnot g19010(.din(n18671), .dout(n19310));
  jand g19011(.dina(n19307), .dinb(n19310), .dout(n19311));
  jnot g19012(.din(n19311), .dout(n19312));
  jand g19013(.dina(n19312), .dinb(n19309), .dout(n19313));
  jand g19014(.dina(n19313), .dinb(n19304), .dout(n19314));
  jor  g19015(.dina(n19314), .dinb(n19303), .dout(n19315));
  jand g19016(.dina(n19315), .dinb(asqrt[38] ), .dout(n19316));
  jor  g19017(.dina(n19303), .dinb(asqrt[38] ), .dout(n19317));
  jor  g19018(.dina(n19317), .dinb(n19314), .dout(n19318));
  jnot g19019(.din(n18677), .dout(n19319));
  jnot g19020(.din(n18679), .dout(n19320));
  jand g19021(.dina(asqrt[4] ), .dinb(n18673), .dout(n19321));
  jand g19022(.dina(n19321), .dinb(n19320), .dout(n19322));
  jor  g19023(.dina(n19322), .dinb(n19319), .dout(n19323));
  jnot g19024(.din(n18680), .dout(n19324));
  jand g19025(.dina(n19321), .dinb(n19324), .dout(n19325));
  jnot g19026(.din(n19325), .dout(n19326));
  jand g19027(.dina(n19326), .dinb(n19323), .dout(n19327));
  jand g19028(.dina(n19327), .dinb(n19318), .dout(n19328));
  jor  g19029(.dina(n19328), .dinb(n19316), .dout(n19329));
  jand g19030(.dina(n19329), .dinb(asqrt[39] ), .dout(n19330));
  jxor g19031(.dina(n18681), .dinb(n3907), .dout(n19331));
  jand g19032(.dina(n19331), .dinb(asqrt[4] ), .dout(n19332));
  jxor g19033(.dina(n19332), .dinb(n18691), .dout(n19333));
  jnot g19034(.din(n19333), .dout(n19334));
  jor  g19035(.dina(n19329), .dinb(asqrt[39] ), .dout(n19335));
  jand g19036(.dina(n19335), .dinb(n19334), .dout(n19336));
  jor  g19037(.dina(n19336), .dinb(n19330), .dout(n19337));
  jand g19038(.dina(n19337), .dinb(asqrt[40] ), .dout(n19338));
  jnot g19039(.din(n18696), .dout(n19339));
  jand g19040(.dina(n19339), .dinb(n18694), .dout(n19340));
  jand g19041(.dina(n19340), .dinb(asqrt[4] ), .dout(n19341));
  jxor g19042(.dina(n19341), .dinb(n18704), .dout(n19342));
  jnot g19043(.din(n19342), .dout(n19343));
  jor  g19044(.dina(n19330), .dinb(asqrt[40] ), .dout(n19344));
  jor  g19045(.dina(n19344), .dinb(n19336), .dout(n19345));
  jand g19046(.dina(n19345), .dinb(n19343), .dout(n19346));
  jor  g19047(.dina(n19346), .dinb(n19338), .dout(n19347));
  jand g19048(.dina(n19347), .dinb(asqrt[41] ), .dout(n19348));
  jor  g19049(.dina(n19347), .dinb(asqrt[41] ), .dout(n19349));
  jnot g19050(.din(n18710), .dout(n19350));
  jnot g19051(.din(n18711), .dout(n19351));
  jand g19052(.dina(asqrt[4] ), .dinb(n18707), .dout(n19352));
  jand g19053(.dina(n19352), .dinb(n19351), .dout(n19353));
  jor  g19054(.dina(n19353), .dinb(n19350), .dout(n19354));
  jnot g19055(.din(n18712), .dout(n19355));
  jand g19056(.dina(n19352), .dinb(n19355), .dout(n19356));
  jnot g19057(.din(n19356), .dout(n19357));
  jand g19058(.dina(n19357), .dinb(n19354), .dout(n19358));
  jand g19059(.dina(n19358), .dinb(n19349), .dout(n19359));
  jor  g19060(.dina(n19359), .dinb(n19348), .dout(n19360));
  jand g19061(.dina(n19360), .dinb(asqrt[42] ), .dout(n19361));
  jor  g19062(.dina(n19348), .dinb(asqrt[42] ), .dout(n19362));
  jor  g19063(.dina(n19362), .dinb(n19359), .dout(n19363));
  jnot g19064(.din(n18718), .dout(n19364));
  jnot g19065(.din(n18720), .dout(n19365));
  jand g19066(.dina(asqrt[4] ), .dinb(n18714), .dout(n19366));
  jand g19067(.dina(n19366), .dinb(n19365), .dout(n19367));
  jor  g19068(.dina(n19367), .dinb(n19364), .dout(n19368));
  jnot g19069(.din(n18721), .dout(n19369));
  jand g19070(.dina(n19366), .dinb(n19369), .dout(n19370));
  jnot g19071(.din(n19370), .dout(n19371));
  jand g19072(.dina(n19371), .dinb(n19368), .dout(n19372));
  jand g19073(.dina(n19372), .dinb(n19363), .dout(n19373));
  jor  g19074(.dina(n19373), .dinb(n19361), .dout(n19374));
  jand g19075(.dina(n19374), .dinb(asqrt[43] ), .dout(n19375));
  jxor g19076(.dina(n18722), .dinb(n2870), .dout(n19376));
  jand g19077(.dina(n19376), .dinb(asqrt[4] ), .dout(n19377));
  jxor g19078(.dina(n19377), .dinb(n18732), .dout(n19378));
  jnot g19079(.din(n19378), .dout(n19379));
  jor  g19080(.dina(n19374), .dinb(asqrt[43] ), .dout(n19380));
  jand g19081(.dina(n19380), .dinb(n19379), .dout(n19381));
  jor  g19082(.dina(n19381), .dinb(n19375), .dout(n19382));
  jand g19083(.dina(n19382), .dinb(asqrt[44] ), .dout(n19383));
  jnot g19084(.din(n18737), .dout(n19384));
  jand g19085(.dina(n19384), .dinb(n18735), .dout(n19385));
  jand g19086(.dina(n19385), .dinb(asqrt[4] ), .dout(n19386));
  jxor g19087(.dina(n19386), .dinb(n18745), .dout(n19387));
  jnot g19088(.din(n19387), .dout(n19388));
  jor  g19089(.dina(n19375), .dinb(asqrt[44] ), .dout(n19389));
  jor  g19090(.dina(n19389), .dinb(n19381), .dout(n19390));
  jand g19091(.dina(n19390), .dinb(n19388), .dout(n19391));
  jor  g19092(.dina(n19391), .dinb(n19383), .dout(n19392));
  jand g19093(.dina(n19392), .dinb(asqrt[45] ), .dout(n19393));
  jor  g19094(.dina(n19392), .dinb(asqrt[45] ), .dout(n19394));
  jnot g19095(.din(n18751), .dout(n19395));
  jnot g19096(.din(n18752), .dout(n19396));
  jand g19097(.dina(asqrt[4] ), .dinb(n18748), .dout(n19397));
  jand g19098(.dina(n19397), .dinb(n19396), .dout(n19398));
  jor  g19099(.dina(n19398), .dinb(n19395), .dout(n19399));
  jnot g19100(.din(n18753), .dout(n19400));
  jand g19101(.dina(n19397), .dinb(n19400), .dout(n19401));
  jnot g19102(.din(n19401), .dout(n19402));
  jand g19103(.dina(n19402), .dinb(n19399), .dout(n19403));
  jand g19104(.dina(n19403), .dinb(n19394), .dout(n19404));
  jor  g19105(.dina(n19404), .dinb(n19393), .dout(n19405));
  jand g19106(.dina(n19405), .dinb(asqrt[46] ), .dout(n19406));
  jor  g19107(.dina(n19393), .dinb(asqrt[46] ), .dout(n19407));
  jor  g19108(.dina(n19407), .dinb(n19404), .dout(n19408));
  jnot g19109(.din(n18759), .dout(n19409));
  jnot g19110(.din(n18761), .dout(n19410));
  jand g19111(.dina(asqrt[4] ), .dinb(n18755), .dout(n19411));
  jand g19112(.dina(n19411), .dinb(n19410), .dout(n19412));
  jor  g19113(.dina(n19412), .dinb(n19409), .dout(n19413));
  jnot g19114(.din(n18762), .dout(n19414));
  jand g19115(.dina(n19411), .dinb(n19414), .dout(n19415));
  jnot g19116(.din(n19415), .dout(n19416));
  jand g19117(.dina(n19416), .dinb(n19413), .dout(n19417));
  jand g19118(.dina(n19417), .dinb(n19408), .dout(n19418));
  jor  g19119(.dina(n19418), .dinb(n19406), .dout(n19419));
  jand g19120(.dina(n19419), .dinb(asqrt[47] ), .dout(n19420));
  jxor g19121(.dina(n18763), .dinb(n2005), .dout(n19421));
  jand g19122(.dina(n19421), .dinb(asqrt[4] ), .dout(n19422));
  jxor g19123(.dina(n19422), .dinb(n18773), .dout(n19423));
  jnot g19124(.din(n19423), .dout(n19424));
  jor  g19125(.dina(n19419), .dinb(asqrt[47] ), .dout(n19425));
  jand g19126(.dina(n19425), .dinb(n19424), .dout(n19426));
  jor  g19127(.dina(n19426), .dinb(n19420), .dout(n19427));
  jand g19128(.dina(n19427), .dinb(asqrt[48] ), .dout(n19428));
  jnot g19129(.din(n18778), .dout(n19429));
  jand g19130(.dina(n19429), .dinb(n18776), .dout(n19430));
  jand g19131(.dina(n19430), .dinb(asqrt[4] ), .dout(n19431));
  jxor g19132(.dina(n19431), .dinb(n18786), .dout(n19432));
  jnot g19133(.din(n19432), .dout(n19433));
  jor  g19134(.dina(n19420), .dinb(asqrt[48] ), .dout(n19434));
  jor  g19135(.dina(n19434), .dinb(n19426), .dout(n19435));
  jand g19136(.dina(n19435), .dinb(n19433), .dout(n19436));
  jor  g19137(.dina(n19436), .dinb(n19428), .dout(n19437));
  jand g19138(.dina(n19437), .dinb(asqrt[49] ), .dout(n19438));
  jor  g19139(.dina(n19437), .dinb(asqrt[49] ), .dout(n19439));
  jnot g19140(.din(n18792), .dout(n19440));
  jnot g19141(.din(n18793), .dout(n19441));
  jand g19142(.dina(asqrt[4] ), .dinb(n18789), .dout(n19442));
  jand g19143(.dina(n19442), .dinb(n19441), .dout(n19443));
  jor  g19144(.dina(n19443), .dinb(n19440), .dout(n19444));
  jnot g19145(.din(n18794), .dout(n19445));
  jand g19146(.dina(n19442), .dinb(n19445), .dout(n19446));
  jnot g19147(.din(n19446), .dout(n19447));
  jand g19148(.dina(n19447), .dinb(n19444), .dout(n19448));
  jand g19149(.dina(n19448), .dinb(n19439), .dout(n19449));
  jor  g19150(.dina(n19449), .dinb(n19438), .dout(n19450));
  jand g19151(.dina(n19450), .dinb(asqrt[50] ), .dout(n19451));
  jor  g19152(.dina(n19438), .dinb(asqrt[50] ), .dout(n19452));
  jor  g19153(.dina(n19452), .dinb(n19449), .dout(n19453));
  jnot g19154(.din(n18800), .dout(n19454));
  jnot g19155(.din(n18802), .dout(n19455));
  jand g19156(.dina(asqrt[4] ), .dinb(n18796), .dout(n19456));
  jand g19157(.dina(n19456), .dinb(n19455), .dout(n19457));
  jor  g19158(.dina(n19457), .dinb(n19454), .dout(n19458));
  jnot g19159(.din(n18803), .dout(n19459));
  jand g19160(.dina(n19456), .dinb(n19459), .dout(n19460));
  jnot g19161(.din(n19460), .dout(n19461));
  jand g19162(.dina(n19461), .dinb(n19458), .dout(n19462));
  jand g19163(.dina(n19462), .dinb(n19453), .dout(n19463));
  jor  g19164(.dina(n19463), .dinb(n19451), .dout(n19464));
  jand g19165(.dina(n19464), .dinb(asqrt[51] ), .dout(n19465));
  jxor g19166(.dina(n18804), .dinb(n1312), .dout(n19466));
  jand g19167(.dina(n19466), .dinb(asqrt[4] ), .dout(n19467));
  jxor g19168(.dina(n19467), .dinb(n18814), .dout(n19468));
  jnot g19169(.din(n19468), .dout(n19469));
  jor  g19170(.dina(n19464), .dinb(asqrt[51] ), .dout(n19470));
  jand g19171(.dina(n19470), .dinb(n19469), .dout(n19471));
  jor  g19172(.dina(n19471), .dinb(n19465), .dout(n19472));
  jand g19173(.dina(n19472), .dinb(asqrt[52] ), .dout(n19473));
  jnot g19174(.din(n18819), .dout(n19474));
  jand g19175(.dina(n19474), .dinb(n18817), .dout(n19475));
  jand g19176(.dina(n19475), .dinb(asqrt[4] ), .dout(n19476));
  jxor g19177(.dina(n19476), .dinb(n18827), .dout(n19477));
  jnot g19178(.din(n19477), .dout(n19478));
  jor  g19179(.dina(n19465), .dinb(asqrt[52] ), .dout(n19479));
  jor  g19180(.dina(n19479), .dinb(n19471), .dout(n19480));
  jand g19181(.dina(n19480), .dinb(n19478), .dout(n19481));
  jor  g19182(.dina(n19481), .dinb(n19473), .dout(n19482));
  jand g19183(.dina(n19482), .dinb(asqrt[53] ), .dout(n19483));
  jor  g19184(.dina(n19482), .dinb(asqrt[53] ), .dout(n19484));
  jnot g19185(.din(n18833), .dout(n19485));
  jnot g19186(.din(n18834), .dout(n19486));
  jand g19187(.dina(asqrt[4] ), .dinb(n18830), .dout(n19487));
  jand g19188(.dina(n19487), .dinb(n19486), .dout(n19488));
  jor  g19189(.dina(n19488), .dinb(n19485), .dout(n19489));
  jnot g19190(.din(n18835), .dout(n19490));
  jand g19191(.dina(n19487), .dinb(n19490), .dout(n19491));
  jnot g19192(.din(n19491), .dout(n19492));
  jand g19193(.dina(n19492), .dinb(n19489), .dout(n19493));
  jand g19194(.dina(n19493), .dinb(n19484), .dout(n19494));
  jor  g19195(.dina(n19494), .dinb(n19483), .dout(n19495));
  jand g19196(.dina(n19495), .dinb(asqrt[54] ), .dout(n19496));
  jor  g19197(.dina(n19483), .dinb(asqrt[54] ), .dout(n19497));
  jor  g19198(.dina(n19497), .dinb(n19494), .dout(n19498));
  jnot g19199(.din(n18841), .dout(n19499));
  jnot g19200(.din(n18843), .dout(n19500));
  jand g19201(.dina(asqrt[4] ), .dinb(n18837), .dout(n19501));
  jand g19202(.dina(n19501), .dinb(n19500), .dout(n19502));
  jor  g19203(.dina(n19502), .dinb(n19499), .dout(n19503));
  jnot g19204(.din(n18844), .dout(n19504));
  jand g19205(.dina(n19501), .dinb(n19504), .dout(n19505));
  jnot g19206(.din(n19505), .dout(n19506));
  jand g19207(.dina(n19506), .dinb(n19503), .dout(n19507));
  jand g19208(.dina(n19507), .dinb(n19498), .dout(n19508));
  jor  g19209(.dina(n19508), .dinb(n19496), .dout(n19509));
  jand g19210(.dina(n19509), .dinb(asqrt[55] ), .dout(n19510));
  jxor g19211(.dina(n18845), .dinb(n791), .dout(n19511));
  jand g19212(.dina(n19511), .dinb(asqrt[4] ), .dout(n19512));
  jxor g19213(.dina(n19512), .dinb(n18855), .dout(n19513));
  jnot g19214(.din(n19513), .dout(n19514));
  jor  g19215(.dina(n19509), .dinb(asqrt[55] ), .dout(n19515));
  jand g19216(.dina(n19515), .dinb(n19514), .dout(n19516));
  jor  g19217(.dina(n19516), .dinb(n19510), .dout(n19517));
  jand g19218(.dina(n19517), .dinb(asqrt[56] ), .dout(n19518));
  jnot g19219(.din(n18860), .dout(n19519));
  jand g19220(.dina(n19519), .dinb(n18858), .dout(n19520));
  jand g19221(.dina(n19520), .dinb(asqrt[4] ), .dout(n19521));
  jxor g19222(.dina(n19521), .dinb(n18868), .dout(n19522));
  jnot g19223(.din(n19522), .dout(n19523));
  jor  g19224(.dina(n19510), .dinb(asqrt[56] ), .dout(n19524));
  jor  g19225(.dina(n19524), .dinb(n19516), .dout(n19525));
  jand g19226(.dina(n19525), .dinb(n19523), .dout(n19526));
  jor  g19227(.dina(n19526), .dinb(n19518), .dout(n19527));
  jand g19228(.dina(n19527), .dinb(asqrt[57] ), .dout(n19528));
  jor  g19229(.dina(n19527), .dinb(asqrt[57] ), .dout(n19529));
  jnot g19230(.din(n18874), .dout(n19530));
  jnot g19231(.din(n18875), .dout(n19531));
  jand g19232(.dina(asqrt[4] ), .dinb(n18871), .dout(n19532));
  jand g19233(.dina(n19532), .dinb(n19531), .dout(n19533));
  jor  g19234(.dina(n19533), .dinb(n19530), .dout(n19534));
  jnot g19235(.din(n18876), .dout(n19535));
  jand g19236(.dina(n19532), .dinb(n19535), .dout(n19536));
  jnot g19237(.din(n19536), .dout(n19537));
  jand g19238(.dina(n19537), .dinb(n19534), .dout(n19538));
  jand g19239(.dina(n19538), .dinb(n19529), .dout(n19539));
  jor  g19240(.dina(n19539), .dinb(n19528), .dout(n19540));
  jand g19241(.dina(n19540), .dinb(asqrt[58] ), .dout(n19541));
  jnot g19242(.din(n18880), .dout(n19542));
  jand g19243(.dina(n19542), .dinb(n18878), .dout(n19543));
  jand g19244(.dina(n19543), .dinb(asqrt[4] ), .dout(n19544));
  jxor g19245(.dina(n19544), .dinb(n18888), .dout(n19545));
  jnot g19246(.din(n19545), .dout(n19546));
  jor  g19247(.dina(n19528), .dinb(asqrt[58] ), .dout(n19547));
  jor  g19248(.dina(n19547), .dinb(n19539), .dout(n19548));
  jand g19249(.dina(n19548), .dinb(n19546), .dout(n19549));
  jor  g19250(.dina(n19549), .dinb(n19541), .dout(n19550));
  jand g19251(.dina(n19550), .dinb(asqrt[59] ), .dout(n19551));
  jor  g19252(.dina(n19550), .dinb(asqrt[59] ), .dout(n19552));
  jand g19253(.dina(n19552), .dinb(n18958), .dout(n19553));
  jor  g19254(.dina(n19553), .dinb(n19551), .dout(n19554));
  jand g19255(.dina(n19554), .dinb(asqrt[60] ), .dout(n19555));
  jor  g19256(.dina(n19551), .dinb(asqrt[60] ), .dout(n19556));
  jor  g19257(.dina(n19556), .dinb(n19553), .dout(n19557));
  jnot g19258(.din(n18900), .dout(n19558));
  jnot g19259(.din(n18902), .dout(n19559));
  jand g19260(.dina(asqrt[4] ), .dinb(n18896), .dout(n19560));
  jand g19261(.dina(n19560), .dinb(n19559), .dout(n19561));
  jor  g19262(.dina(n19561), .dinb(n19558), .dout(n19562));
  jnot g19263(.din(n18903), .dout(n19563));
  jand g19264(.dina(n19560), .dinb(n19563), .dout(n19564));
  jnot g19265(.din(n19564), .dout(n19565));
  jand g19266(.dina(n19565), .dinb(n19562), .dout(n19566));
  jand g19267(.dina(n19566), .dinb(n19557), .dout(n19567));
  jor  g19268(.dina(n19567), .dinb(n19555), .dout(n19568));
  jand g19269(.dina(n19568), .dinb(asqrt[61] ), .dout(n19569));
  jor  g19270(.dina(n19568), .dinb(asqrt[61] ), .dout(n19570));
  jnot g19271(.din(n18908), .dout(n19571));
  jnot g19272(.din(n18909), .dout(n19572));
  jand g19273(.dina(asqrt[4] ), .dinb(n18905), .dout(n19573));
  jand g19274(.dina(n19573), .dinb(n19572), .dout(n19574));
  jor  g19275(.dina(n19574), .dinb(n19571), .dout(n19575));
  jnot g19276(.din(n18910), .dout(n19576));
  jand g19277(.dina(n19573), .dinb(n19576), .dout(n19577));
  jnot g19278(.din(n19577), .dout(n19578));
  jand g19279(.dina(n19578), .dinb(n19575), .dout(n19579));
  jand g19280(.dina(n19579), .dinb(n19570), .dout(n19580));
  jor  g19281(.dina(n19580), .dinb(n19569), .dout(n19581));
  jand g19282(.dina(n19581), .dinb(asqrt[62] ), .dout(n19582));
  jor  g19283(.dina(n19569), .dinb(asqrt[62] ), .dout(n19583));
  jor  g19284(.dina(n19583), .dinb(n19580), .dout(n19584));
  jnot g19285(.din(n18916), .dout(n19585));
  jnot g19286(.din(n18918), .dout(n19586));
  jand g19287(.dina(asqrt[4] ), .dinb(n18912), .dout(n19587));
  jand g19288(.dina(n19587), .dinb(n19586), .dout(n19588));
  jor  g19289(.dina(n19588), .dinb(n19585), .dout(n19589));
  jnot g19290(.din(n18919), .dout(n19590));
  jand g19291(.dina(n19587), .dinb(n19590), .dout(n19591));
  jnot g19292(.din(n19591), .dout(n19592));
  jand g19293(.dina(n19592), .dinb(n19589), .dout(n19593));
  jand g19294(.dina(n19593), .dinb(n19584), .dout(n19594));
  jor  g19295(.dina(n19594), .dinb(n19582), .dout(n19595));
  jxor g19296(.dina(n18920), .dinb(n199), .dout(n19596));
  jand g19297(.dina(n19596), .dinb(asqrt[4] ), .dout(n19597));
  jxor g19298(.dina(n19597), .dinb(n18930), .dout(n19598));
  jnot g19299(.din(n18932), .dout(n19599));
  jand g19300(.dina(asqrt[4] ), .dinb(n18939), .dout(n19600));
  jand g19301(.dina(n19600), .dinb(n19599), .dout(n19601));
  jor  g19302(.dina(n19601), .dinb(n18948), .dout(n19602));
  jor  g19303(.dina(n19602), .dinb(n19598), .dout(n19603));
  jnot g19304(.din(n19603), .dout(n19604));
  jand g19305(.dina(n19604), .dinb(n19595), .dout(n19605));
  jor  g19306(.dina(n19605), .dinb(asqrt[63] ), .dout(n19606));
  jnot g19307(.din(n19598), .dout(n19607));
  jor  g19308(.dina(n19607), .dinb(n19595), .dout(n19608));
  jor  g19309(.dina(n19600), .dinb(n19599), .dout(n19609));
  jand g19310(.dina(n18939), .dinb(n19599), .dout(n19610));
  jor  g19311(.dina(n19610), .dinb(n194), .dout(n19611));
  jnot g19312(.din(n19611), .dout(n19612));
  jand g19313(.dina(n19612), .dinb(n19609), .dout(n19613));
  jnot g19314(.din(n19613), .dout(n19614));
  jand g19315(.dina(n19614), .dinb(n19608), .dout(n19615));
  jand g19316(.dina(n19615), .dinb(n19606), .dout(n19616));
  jxor g19317(.dina(n19550), .dinb(n305), .dout(n19617));
  jor  g19318(.dina(n19617), .dinb(n19616), .dout(n19618));
  jxor g19319(.dina(n19618), .dinb(n18959), .dout(n19619));
  jnot g19320(.din(n19619), .dout(n19620));
  jor  g19321(.dina(n19616), .dinb(n18961), .dout(n19621));
  jnot g19322(.din(a[4] ), .dout(n19622));
  jnot g19323(.din(a[5] ), .dout(n19623));
  jand g19324(.dina(n18961), .dinb(n19623), .dout(n19624));
  jand g19325(.dina(n19624), .dinb(n19622), .dout(n19625));
  jnot g19326(.din(n19625), .dout(n19626));
  jand g19327(.dina(n19626), .dinb(n19621), .dout(n19627));
  jor  g19328(.dina(n19627), .dinb(n18976), .dout(n19628));
  jor  g19329(.dina(n19616), .dinb(a[6] ), .dout(n19629));
  jxor g19330(.dina(n19629), .dinb(n18962), .dout(n19630));
  jand g19331(.dina(n19627), .dinb(n18976), .dout(n19631));
  jor  g19332(.dina(n19631), .dinb(n19630), .dout(n19632));
  jand g19333(.dina(n19632), .dinb(n19628), .dout(n19633));
  jor  g19334(.dina(n19633), .dinb(n18356), .dout(n19634));
  jand g19335(.dina(n19628), .dinb(n18356), .dout(n19635));
  jand g19336(.dina(n19635), .dinb(n19632), .dout(n19636));
  jor  g19337(.dina(n19629), .dinb(a[7] ), .dout(n19637));
  jnot g19338(.din(n19616), .dout(asqrt[3] ));
  jor  g19339(.dina(asqrt[3] ), .dinb(n18976), .dout(n19639));
  jand g19340(.dina(n19639), .dinb(n19637), .dout(n19640));
  jxor g19341(.dina(n19640), .dinb(n18362), .dout(n19641));
  jor  g19342(.dina(n19641), .dinb(n19636), .dout(n19642));
  jand g19343(.dina(n19642), .dinb(n19634), .dout(n19643));
  jor  g19344(.dina(n19643), .dinb(n18360), .dout(n19644));
  jand g19345(.dina(n19643), .dinb(n18360), .dout(n19645));
  jxor g19346(.dina(n18965), .dinb(n18356), .dout(n19646));
  jor  g19347(.dina(n19646), .dinb(n19616), .dout(n19647));
  jxor g19348(.dina(n19647), .dinb(n18968), .dout(n19648));
  jor  g19349(.dina(n19648), .dinb(n19645), .dout(n19649));
  jand g19350(.dina(n19649), .dinb(n19644), .dout(n19650));
  jor  g19351(.dina(n19650), .dinb(n17140), .dout(n19651));
  jnot g19352(.din(n18974), .dout(n19652));
  jor  g19353(.dina(n19652), .dinb(n18972), .dout(n19653));
  jor  g19354(.dina(n19653), .dinb(n19616), .dout(n19654));
  jxor g19355(.dina(n19654), .dinb(n18979), .dout(n19655));
  jand g19356(.dina(n19644), .dinb(n17140), .dout(n19656));
  jand g19357(.dina(n19656), .dinb(n19649), .dout(n19657));
  jor  g19358(.dina(n19657), .dinb(n19655), .dout(n19658));
  jand g19359(.dina(n19658), .dinb(n19651), .dout(n19659));
  jor  g19360(.dina(n19659), .dinb(n17135), .dout(n19660));
  jand g19361(.dina(n19659), .dinb(n17135), .dout(n19661));
  jxor g19362(.dina(n18981), .dinb(n17140), .dout(n19662));
  jor  g19363(.dina(n19662), .dinb(n19616), .dout(n19663));
  jxor g19364(.dina(n19663), .dinb(n18986), .dout(n19664));
  jnot g19365(.din(n19664), .dout(n19665));
  jor  g19366(.dina(n19665), .dinb(n19661), .dout(n19666));
  jand g19367(.dina(n19666), .dinb(n19660), .dout(n19667));
  jor  g19368(.dina(n19667), .dinb(n15955), .dout(n19668));
  jand g19369(.dina(n19660), .dinb(n15955), .dout(n19669));
  jand g19370(.dina(n19669), .dinb(n19666), .dout(n19670));
  jnot g19371(.din(n18990), .dout(n19671));
  jand g19372(.dina(asqrt[3] ), .dinb(n19671), .dout(n19672));
  jand g19373(.dina(n19672), .dinb(n18997), .dout(n19673));
  jor  g19374(.dina(n19673), .dinb(n18995), .dout(n19674));
  jand g19375(.dina(n19672), .dinb(n18998), .dout(n19675));
  jnot g19376(.din(n19675), .dout(n19676));
  jand g19377(.dina(n19676), .dinb(n19674), .dout(n19677));
  jnot g19378(.din(n19677), .dout(n19678));
  jor  g19379(.dina(n19678), .dinb(n19670), .dout(n19679));
  jand g19380(.dina(n19679), .dinb(n19668), .dout(n19680));
  jor  g19381(.dina(n19680), .dinb(n15950), .dout(n19681));
  jand g19382(.dina(n19680), .dinb(n15950), .dout(n19682));
  jnot g19383(.din(n19005), .dout(n19683));
  jxor g19384(.dina(n18999), .dinb(n15955), .dout(n19684));
  jor  g19385(.dina(n19684), .dinb(n19616), .dout(n19685));
  jxor g19386(.dina(n19685), .dinb(n19683), .dout(n19686));
  jnot g19387(.din(n19686), .dout(n19687));
  jor  g19388(.dina(n19687), .dinb(n19682), .dout(n19688));
  jand g19389(.dina(n19688), .dinb(n19681), .dout(n19689));
  jor  g19390(.dina(n19689), .dinb(n14821), .dout(n19690));
  jnot g19391(.din(n19010), .dout(n19691));
  jor  g19392(.dina(n19691), .dinb(n19008), .dout(n19692));
  jor  g19393(.dina(n19692), .dinb(n19616), .dout(n19693));
  jxor g19394(.dina(n19693), .dinb(n19019), .dout(n19694));
  jand g19395(.dina(n19681), .dinb(n14821), .dout(n19695));
  jand g19396(.dina(n19695), .dinb(n19688), .dout(n19696));
  jor  g19397(.dina(n19696), .dinb(n19694), .dout(n19697));
  jand g19398(.dina(n19697), .dinb(n19690), .dout(n19698));
  jor  g19399(.dina(n19698), .dinb(n14816), .dout(n19699));
  jand g19400(.dina(n19698), .dinb(n14816), .dout(n19700));
  jnot g19401(.din(n19026), .dout(n19701));
  jxor g19402(.dina(n19021), .dinb(n14821), .dout(n19702));
  jor  g19403(.dina(n19702), .dinb(n19616), .dout(n19703));
  jxor g19404(.dina(n19703), .dinb(n19701), .dout(n19704));
  jnot g19405(.din(n19704), .dout(n19705));
  jor  g19406(.dina(n19705), .dinb(n19700), .dout(n19706));
  jand g19407(.dina(n19706), .dinb(n19699), .dout(n19707));
  jor  g19408(.dina(n19707), .dinb(n13723), .dout(n19708));
  jand g19409(.dina(n19699), .dinb(n13723), .dout(n19709));
  jand g19410(.dina(n19709), .dinb(n19706), .dout(n19710));
  jnot g19411(.din(n19029), .dout(n19711));
  jand g19412(.dina(asqrt[3] ), .dinb(n19711), .dout(n19712));
  jand g19413(.dina(n19712), .dinb(n19036), .dout(n19713));
  jor  g19414(.dina(n19713), .dinb(n19034), .dout(n19714));
  jand g19415(.dina(n19712), .dinb(n19037), .dout(n19715));
  jnot g19416(.din(n19715), .dout(n19716));
  jand g19417(.dina(n19716), .dinb(n19714), .dout(n19717));
  jnot g19418(.din(n19717), .dout(n19718));
  jor  g19419(.dina(n19718), .dinb(n19710), .dout(n19719));
  jand g19420(.dina(n19719), .dinb(n19708), .dout(n19720));
  jor  g19421(.dina(n19720), .dinb(n13718), .dout(n19721));
  jxor g19422(.dina(n19038), .dinb(n13723), .dout(n19722));
  jor  g19423(.dina(n19722), .dinb(n19616), .dout(n19723));
  jxor g19424(.dina(n19723), .dinb(n19043), .dout(n19724));
  jand g19425(.dina(n19720), .dinb(n13718), .dout(n19725));
  jor  g19426(.dina(n19725), .dinb(n19724), .dout(n19726));
  jand g19427(.dina(n19726), .dinb(n19721), .dout(n19727));
  jor  g19428(.dina(n19727), .dinb(n12675), .dout(n19728));
  jnot g19429(.din(n19048), .dout(n19729));
  jor  g19430(.dina(n19729), .dinb(n19046), .dout(n19730));
  jor  g19431(.dina(n19730), .dinb(n19616), .dout(n19731));
  jxor g19432(.dina(n19731), .dinb(n19057), .dout(n19732));
  jand g19433(.dina(n19721), .dinb(n12675), .dout(n19733));
  jand g19434(.dina(n19733), .dinb(n19726), .dout(n19734));
  jor  g19435(.dina(n19734), .dinb(n19732), .dout(n19735));
  jand g19436(.dina(n19735), .dinb(n19728), .dout(n19736));
  jor  g19437(.dina(n19736), .dinb(n12670), .dout(n19737));
  jand g19438(.dina(n19736), .dinb(n12670), .dout(n19738));
  jnot g19439(.din(n19060), .dout(n19739));
  jand g19440(.dina(asqrt[3] ), .dinb(n19739), .dout(n19740));
  jand g19441(.dina(n19740), .dinb(n19065), .dout(n19741));
  jor  g19442(.dina(n19741), .dinb(n19064), .dout(n19742));
  jand g19443(.dina(n19740), .dinb(n19066), .dout(n19743));
  jnot g19444(.din(n19743), .dout(n19744));
  jand g19445(.dina(n19744), .dinb(n19742), .dout(n19745));
  jnot g19446(.din(n19745), .dout(n19746));
  jor  g19447(.dina(n19746), .dinb(n19738), .dout(n19747));
  jand g19448(.dina(n19747), .dinb(n19737), .dout(n19748));
  jor  g19449(.dina(n19748), .dinb(n11662), .dout(n19749));
  jand g19450(.dina(n19737), .dinb(n11662), .dout(n19750));
  jand g19451(.dina(n19750), .dinb(n19747), .dout(n19751));
  jnot g19452(.din(n19068), .dout(n19752));
  jand g19453(.dina(asqrt[3] ), .dinb(n19752), .dout(n19753));
  jand g19454(.dina(n19753), .dinb(n19075), .dout(n19754));
  jor  g19455(.dina(n19754), .dinb(n19073), .dout(n19755));
  jand g19456(.dina(n19753), .dinb(n19076), .dout(n19756));
  jnot g19457(.din(n19756), .dout(n19757));
  jand g19458(.dina(n19757), .dinb(n19755), .dout(n19758));
  jnot g19459(.din(n19758), .dout(n19759));
  jor  g19460(.dina(n19759), .dinb(n19751), .dout(n19760));
  jand g19461(.dina(n19760), .dinb(n19749), .dout(n19761));
  jor  g19462(.dina(n19761), .dinb(n11657), .dout(n19762));
  jxor g19463(.dina(n19077), .dinb(n11662), .dout(n19763));
  jor  g19464(.dina(n19763), .dinb(n19616), .dout(n19764));
  jxor g19465(.dina(n19764), .dinb(n19088), .dout(n19765));
  jand g19466(.dina(n19761), .dinb(n11657), .dout(n19766));
  jor  g19467(.dina(n19766), .dinb(n19765), .dout(n19767));
  jand g19468(.dina(n19767), .dinb(n19762), .dout(n19768));
  jor  g19469(.dina(n19768), .dinb(n10701), .dout(n19769));
  jnot g19470(.din(n19093), .dout(n19770));
  jor  g19471(.dina(n19770), .dinb(n19091), .dout(n19771));
  jor  g19472(.dina(n19771), .dinb(n19616), .dout(n19772));
  jxor g19473(.dina(n19772), .dinb(n19102), .dout(n19773));
  jand g19474(.dina(n19762), .dinb(n10701), .dout(n19774));
  jand g19475(.dina(n19774), .dinb(n19767), .dout(n19775));
  jor  g19476(.dina(n19775), .dinb(n19773), .dout(n19776));
  jand g19477(.dina(n19776), .dinb(n19769), .dout(n19777));
  jor  g19478(.dina(n19777), .dinb(n10696), .dout(n19778));
  jand g19479(.dina(n19777), .dinb(n10696), .dout(n19779));
  jnot g19480(.din(n19105), .dout(n19780));
  jand g19481(.dina(asqrt[3] ), .dinb(n19780), .dout(n19781));
  jand g19482(.dina(n19781), .dinb(n19110), .dout(n19782));
  jor  g19483(.dina(n19782), .dinb(n19109), .dout(n19783));
  jand g19484(.dina(n19781), .dinb(n19111), .dout(n19784));
  jnot g19485(.din(n19784), .dout(n19785));
  jand g19486(.dina(n19785), .dinb(n19783), .dout(n19786));
  jnot g19487(.din(n19786), .dout(n19787));
  jor  g19488(.dina(n19787), .dinb(n19779), .dout(n19788));
  jand g19489(.dina(n19788), .dinb(n19778), .dout(n19789));
  jor  g19490(.dina(n19789), .dinb(n9774), .dout(n19790));
  jand g19491(.dina(n19778), .dinb(n9774), .dout(n19791));
  jand g19492(.dina(n19791), .dinb(n19788), .dout(n19792));
  jnot g19493(.din(n19113), .dout(n19793));
  jand g19494(.dina(asqrt[3] ), .dinb(n19793), .dout(n19794));
  jand g19495(.dina(n19794), .dinb(n19120), .dout(n19795));
  jor  g19496(.dina(n19795), .dinb(n19118), .dout(n19796));
  jand g19497(.dina(n19794), .dinb(n19121), .dout(n19797));
  jnot g19498(.din(n19797), .dout(n19798));
  jand g19499(.dina(n19798), .dinb(n19796), .dout(n19799));
  jnot g19500(.din(n19799), .dout(n19800));
  jor  g19501(.dina(n19800), .dinb(n19792), .dout(n19801));
  jand g19502(.dina(n19801), .dinb(n19790), .dout(n19802));
  jor  g19503(.dina(n19802), .dinb(n9769), .dout(n19803));
  jxor g19504(.dina(n19122), .dinb(n9774), .dout(n19804));
  jor  g19505(.dina(n19804), .dinb(n19616), .dout(n19805));
  jxor g19506(.dina(n19805), .dinb(n19133), .dout(n19806));
  jand g19507(.dina(n19802), .dinb(n9769), .dout(n19807));
  jor  g19508(.dina(n19807), .dinb(n19806), .dout(n19808));
  jand g19509(.dina(n19808), .dinb(n19803), .dout(n19809));
  jor  g19510(.dina(n19809), .dinb(n8898), .dout(n19810));
  jnot g19511(.din(n19138), .dout(n19811));
  jor  g19512(.dina(n19811), .dinb(n19136), .dout(n19812));
  jor  g19513(.dina(n19812), .dinb(n19616), .dout(n19813));
  jxor g19514(.dina(n19813), .dinb(n19147), .dout(n19814));
  jand g19515(.dina(n19803), .dinb(n8898), .dout(n19815));
  jand g19516(.dina(n19815), .dinb(n19808), .dout(n19816));
  jor  g19517(.dina(n19816), .dinb(n19814), .dout(n19817));
  jand g19518(.dina(n19817), .dinb(n19810), .dout(n19818));
  jor  g19519(.dina(n19818), .dinb(n8893), .dout(n19819));
  jand g19520(.dina(n19818), .dinb(n8893), .dout(n19820));
  jnot g19521(.din(n19150), .dout(n19821));
  jand g19522(.dina(asqrt[3] ), .dinb(n19821), .dout(n19822));
  jand g19523(.dina(n19822), .dinb(n19155), .dout(n19823));
  jor  g19524(.dina(n19823), .dinb(n19154), .dout(n19824));
  jand g19525(.dina(n19822), .dinb(n19156), .dout(n19825));
  jnot g19526(.din(n19825), .dout(n19826));
  jand g19527(.dina(n19826), .dinb(n19824), .dout(n19827));
  jnot g19528(.din(n19827), .dout(n19828));
  jor  g19529(.dina(n19828), .dinb(n19820), .dout(n19829));
  jand g19530(.dina(n19829), .dinb(n19819), .dout(n19830));
  jor  g19531(.dina(n19830), .dinb(n8058), .dout(n19831));
  jand g19532(.dina(n19819), .dinb(n8058), .dout(n19832));
  jand g19533(.dina(n19832), .dinb(n19829), .dout(n19833));
  jnot g19534(.din(n19158), .dout(n19834));
  jand g19535(.dina(asqrt[3] ), .dinb(n19834), .dout(n19835));
  jand g19536(.dina(n19835), .dinb(n19165), .dout(n19836));
  jor  g19537(.dina(n19836), .dinb(n19163), .dout(n19837));
  jand g19538(.dina(n19835), .dinb(n19166), .dout(n19838));
  jnot g19539(.din(n19838), .dout(n19839));
  jand g19540(.dina(n19839), .dinb(n19837), .dout(n19840));
  jnot g19541(.din(n19840), .dout(n19841));
  jor  g19542(.dina(n19841), .dinb(n19833), .dout(n19842));
  jand g19543(.dina(n19842), .dinb(n19831), .dout(n19843));
  jor  g19544(.dina(n19843), .dinb(n8053), .dout(n19844));
  jxor g19545(.dina(n19167), .dinb(n8058), .dout(n19845));
  jor  g19546(.dina(n19845), .dinb(n19616), .dout(n19846));
  jxor g19547(.dina(n19846), .dinb(n19178), .dout(n19847));
  jand g19548(.dina(n19843), .dinb(n8053), .dout(n19848));
  jor  g19549(.dina(n19848), .dinb(n19847), .dout(n19849));
  jand g19550(.dina(n19849), .dinb(n19844), .dout(n19850));
  jor  g19551(.dina(n19850), .dinb(n7265), .dout(n19851));
  jnot g19552(.din(n19183), .dout(n19852));
  jor  g19553(.dina(n19852), .dinb(n19181), .dout(n19853));
  jor  g19554(.dina(n19853), .dinb(n19616), .dout(n19854));
  jxor g19555(.dina(n19854), .dinb(n19192), .dout(n19855));
  jand g19556(.dina(n19844), .dinb(n7265), .dout(n19856));
  jand g19557(.dina(n19856), .dinb(n19849), .dout(n19857));
  jor  g19558(.dina(n19857), .dinb(n19855), .dout(n19858));
  jand g19559(.dina(n19858), .dinb(n19851), .dout(n19859));
  jor  g19560(.dina(n19859), .dinb(n7260), .dout(n19860));
  jand g19561(.dina(n19859), .dinb(n7260), .dout(n19861));
  jnot g19562(.din(n19195), .dout(n19862));
  jand g19563(.dina(asqrt[3] ), .dinb(n19862), .dout(n19863));
  jand g19564(.dina(n19863), .dinb(n19200), .dout(n19864));
  jor  g19565(.dina(n19864), .dinb(n19199), .dout(n19865));
  jand g19566(.dina(n19863), .dinb(n19201), .dout(n19866));
  jnot g19567(.din(n19866), .dout(n19867));
  jand g19568(.dina(n19867), .dinb(n19865), .dout(n19868));
  jnot g19569(.din(n19868), .dout(n19869));
  jor  g19570(.dina(n19869), .dinb(n19861), .dout(n19870));
  jand g19571(.dina(n19870), .dinb(n19860), .dout(n19871));
  jor  g19572(.dina(n19871), .dinb(n6505), .dout(n19872));
  jand g19573(.dina(n19860), .dinb(n6505), .dout(n19873));
  jand g19574(.dina(n19873), .dinb(n19870), .dout(n19874));
  jnot g19575(.din(n19203), .dout(n19875));
  jand g19576(.dina(asqrt[3] ), .dinb(n19875), .dout(n19876));
  jand g19577(.dina(n19876), .dinb(n19210), .dout(n19877));
  jor  g19578(.dina(n19877), .dinb(n19208), .dout(n19878));
  jand g19579(.dina(n19876), .dinb(n19211), .dout(n19879));
  jnot g19580(.din(n19879), .dout(n19880));
  jand g19581(.dina(n19880), .dinb(n19878), .dout(n19881));
  jnot g19582(.din(n19881), .dout(n19882));
  jor  g19583(.dina(n19882), .dinb(n19874), .dout(n19883));
  jand g19584(.dina(n19883), .dinb(n19872), .dout(n19884));
  jor  g19585(.dina(n19884), .dinb(n6500), .dout(n19885));
  jxor g19586(.dina(n19212), .dinb(n6505), .dout(n19886));
  jor  g19587(.dina(n19886), .dinb(n19616), .dout(n19887));
  jxor g19588(.dina(n19887), .dinb(n19223), .dout(n19888));
  jand g19589(.dina(n19884), .dinb(n6500), .dout(n19889));
  jor  g19590(.dina(n19889), .dinb(n19888), .dout(n19890));
  jand g19591(.dina(n19890), .dinb(n19885), .dout(n19891));
  jor  g19592(.dina(n19891), .dinb(n5793), .dout(n19892));
  jnot g19593(.din(n19228), .dout(n19893));
  jor  g19594(.dina(n19893), .dinb(n19226), .dout(n19894));
  jor  g19595(.dina(n19894), .dinb(n19616), .dout(n19895));
  jxor g19596(.dina(n19895), .dinb(n19237), .dout(n19896));
  jand g19597(.dina(n19885), .dinb(n5793), .dout(n19897));
  jand g19598(.dina(n19897), .dinb(n19890), .dout(n19898));
  jor  g19599(.dina(n19898), .dinb(n19896), .dout(n19899));
  jand g19600(.dina(n19899), .dinb(n19892), .dout(n19900));
  jor  g19601(.dina(n19900), .dinb(n5788), .dout(n19901));
  jand g19602(.dina(n19900), .dinb(n5788), .dout(n19902));
  jnot g19603(.din(n19240), .dout(n19903));
  jand g19604(.dina(asqrt[3] ), .dinb(n19903), .dout(n19904));
  jand g19605(.dina(n19904), .dinb(n19245), .dout(n19905));
  jor  g19606(.dina(n19905), .dinb(n19244), .dout(n19906));
  jand g19607(.dina(n19904), .dinb(n19246), .dout(n19907));
  jnot g19608(.din(n19907), .dout(n19908));
  jand g19609(.dina(n19908), .dinb(n19906), .dout(n19909));
  jnot g19610(.din(n19909), .dout(n19910));
  jor  g19611(.dina(n19910), .dinb(n19902), .dout(n19911));
  jand g19612(.dina(n19911), .dinb(n19901), .dout(n19912));
  jor  g19613(.dina(n19912), .dinb(n5121), .dout(n19913));
  jand g19614(.dina(n19901), .dinb(n5121), .dout(n19914));
  jand g19615(.dina(n19914), .dinb(n19911), .dout(n19915));
  jnot g19616(.din(n19248), .dout(n19916));
  jand g19617(.dina(asqrt[3] ), .dinb(n19916), .dout(n19917));
  jand g19618(.dina(n19917), .dinb(n19255), .dout(n19918));
  jor  g19619(.dina(n19918), .dinb(n19253), .dout(n19919));
  jand g19620(.dina(n19917), .dinb(n19256), .dout(n19920));
  jnot g19621(.din(n19920), .dout(n19921));
  jand g19622(.dina(n19921), .dinb(n19919), .dout(n19922));
  jnot g19623(.din(n19922), .dout(n19923));
  jor  g19624(.dina(n19923), .dinb(n19915), .dout(n19924));
  jand g19625(.dina(n19924), .dinb(n19913), .dout(n19925));
  jor  g19626(.dina(n19925), .dinb(n5116), .dout(n19926));
  jxor g19627(.dina(n19257), .dinb(n5121), .dout(n19927));
  jor  g19628(.dina(n19927), .dinb(n19616), .dout(n19928));
  jxor g19629(.dina(n19928), .dinb(n19268), .dout(n19929));
  jand g19630(.dina(n19925), .dinb(n5116), .dout(n19930));
  jor  g19631(.dina(n19930), .dinb(n19929), .dout(n19931));
  jand g19632(.dina(n19931), .dinb(n19926), .dout(n19932));
  jor  g19633(.dina(n19932), .dinb(n4499), .dout(n19933));
  jnot g19634(.din(n19273), .dout(n19934));
  jor  g19635(.dina(n19934), .dinb(n19271), .dout(n19935));
  jor  g19636(.dina(n19935), .dinb(n19616), .dout(n19936));
  jxor g19637(.dina(n19936), .dinb(n19282), .dout(n19937));
  jand g19638(.dina(n19926), .dinb(n4499), .dout(n19938));
  jand g19639(.dina(n19938), .dinb(n19931), .dout(n19939));
  jor  g19640(.dina(n19939), .dinb(n19937), .dout(n19940));
  jand g19641(.dina(n19940), .dinb(n19933), .dout(n19941));
  jor  g19642(.dina(n19941), .dinb(n4494), .dout(n19942));
  jand g19643(.dina(n19941), .dinb(n4494), .dout(n19943));
  jnot g19644(.din(n19285), .dout(n19944));
  jand g19645(.dina(asqrt[3] ), .dinb(n19944), .dout(n19945));
  jand g19646(.dina(n19945), .dinb(n19290), .dout(n19946));
  jor  g19647(.dina(n19946), .dinb(n19289), .dout(n19947));
  jand g19648(.dina(n19945), .dinb(n19291), .dout(n19948));
  jnot g19649(.din(n19948), .dout(n19949));
  jand g19650(.dina(n19949), .dinb(n19947), .dout(n19950));
  jnot g19651(.din(n19950), .dout(n19951));
  jor  g19652(.dina(n19951), .dinb(n19943), .dout(n19952));
  jand g19653(.dina(n19952), .dinb(n19942), .dout(n19953));
  jor  g19654(.dina(n19953), .dinb(n3912), .dout(n19954));
  jand g19655(.dina(n19942), .dinb(n3912), .dout(n19955));
  jand g19656(.dina(n19955), .dinb(n19952), .dout(n19956));
  jnot g19657(.din(n19293), .dout(n19957));
  jand g19658(.dina(asqrt[3] ), .dinb(n19957), .dout(n19958));
  jand g19659(.dina(n19958), .dinb(n19300), .dout(n19959));
  jor  g19660(.dina(n19959), .dinb(n19298), .dout(n19960));
  jand g19661(.dina(n19958), .dinb(n19301), .dout(n19961));
  jnot g19662(.din(n19961), .dout(n19962));
  jand g19663(.dina(n19962), .dinb(n19960), .dout(n19963));
  jnot g19664(.din(n19963), .dout(n19964));
  jor  g19665(.dina(n19964), .dinb(n19956), .dout(n19965));
  jand g19666(.dina(n19965), .dinb(n19954), .dout(n19966));
  jor  g19667(.dina(n19966), .dinb(n3907), .dout(n19967));
  jxor g19668(.dina(n19302), .dinb(n3912), .dout(n19968));
  jor  g19669(.dina(n19968), .dinb(n19616), .dout(n19969));
  jxor g19670(.dina(n19969), .dinb(n19313), .dout(n19970));
  jand g19671(.dina(n19966), .dinb(n3907), .dout(n19971));
  jor  g19672(.dina(n19971), .dinb(n19970), .dout(n19972));
  jand g19673(.dina(n19972), .dinb(n19967), .dout(n19973));
  jor  g19674(.dina(n19973), .dinb(n3376), .dout(n19974));
  jnot g19675(.din(n19318), .dout(n19975));
  jor  g19676(.dina(n19975), .dinb(n19316), .dout(n19976));
  jor  g19677(.dina(n19976), .dinb(n19616), .dout(n19977));
  jxor g19678(.dina(n19977), .dinb(n19327), .dout(n19978));
  jand g19679(.dina(n19967), .dinb(n3376), .dout(n19979));
  jand g19680(.dina(n19979), .dinb(n19972), .dout(n19980));
  jor  g19681(.dina(n19980), .dinb(n19978), .dout(n19981));
  jand g19682(.dina(n19981), .dinb(n19974), .dout(n19982));
  jor  g19683(.dina(n19982), .dinb(n3371), .dout(n19983));
  jand g19684(.dina(n19982), .dinb(n3371), .dout(n19984));
  jnot g19685(.din(n19330), .dout(n19985));
  jand g19686(.dina(asqrt[3] ), .dinb(n19985), .dout(n19986));
  jand g19687(.dina(n19986), .dinb(n19335), .dout(n19987));
  jor  g19688(.dina(n19987), .dinb(n19334), .dout(n19988));
  jand g19689(.dina(n19986), .dinb(n19336), .dout(n19989));
  jnot g19690(.din(n19989), .dout(n19990));
  jand g19691(.dina(n19990), .dinb(n19988), .dout(n19991));
  jnot g19692(.din(n19991), .dout(n19992));
  jor  g19693(.dina(n19992), .dinb(n19984), .dout(n19993));
  jand g19694(.dina(n19993), .dinb(n19983), .dout(n19994));
  jor  g19695(.dina(n19994), .dinb(n2875), .dout(n19995));
  jand g19696(.dina(n19983), .dinb(n2875), .dout(n19996));
  jand g19697(.dina(n19996), .dinb(n19993), .dout(n19997));
  jnot g19698(.din(n19338), .dout(n19998));
  jand g19699(.dina(asqrt[3] ), .dinb(n19998), .dout(n19999));
  jand g19700(.dina(n19999), .dinb(n19345), .dout(n20000));
  jor  g19701(.dina(n20000), .dinb(n19343), .dout(n20001));
  jand g19702(.dina(n19999), .dinb(n19346), .dout(n20002));
  jnot g19703(.din(n20002), .dout(n20003));
  jand g19704(.dina(n20003), .dinb(n20001), .dout(n20004));
  jnot g19705(.din(n20004), .dout(n20005));
  jor  g19706(.dina(n20005), .dinb(n19997), .dout(n20006));
  jand g19707(.dina(n20006), .dinb(n19995), .dout(n20007));
  jor  g19708(.dina(n20007), .dinb(n2870), .dout(n20008));
  jxor g19709(.dina(n19347), .dinb(n2875), .dout(n20009));
  jor  g19710(.dina(n20009), .dinb(n19616), .dout(n20010));
  jxor g19711(.dina(n20010), .dinb(n19358), .dout(n20011));
  jand g19712(.dina(n20007), .dinb(n2870), .dout(n20012));
  jor  g19713(.dina(n20012), .dinb(n20011), .dout(n20013));
  jand g19714(.dina(n20013), .dinb(n20008), .dout(n20014));
  jor  g19715(.dina(n20014), .dinb(n2425), .dout(n20015));
  jnot g19716(.din(n19363), .dout(n20016));
  jor  g19717(.dina(n20016), .dinb(n19361), .dout(n20017));
  jor  g19718(.dina(n20017), .dinb(n19616), .dout(n20018));
  jxor g19719(.dina(n20018), .dinb(n19372), .dout(n20019));
  jand g19720(.dina(n20008), .dinb(n2425), .dout(n20020));
  jand g19721(.dina(n20020), .dinb(n20013), .dout(n20021));
  jor  g19722(.dina(n20021), .dinb(n20019), .dout(n20022));
  jand g19723(.dina(n20022), .dinb(n20015), .dout(n20023));
  jor  g19724(.dina(n20023), .dinb(n2420), .dout(n20024));
  jand g19725(.dina(n20023), .dinb(n2420), .dout(n20025));
  jnot g19726(.din(n19375), .dout(n20026));
  jand g19727(.dina(asqrt[3] ), .dinb(n20026), .dout(n20027));
  jand g19728(.dina(n20027), .dinb(n19380), .dout(n20028));
  jor  g19729(.dina(n20028), .dinb(n19379), .dout(n20029));
  jand g19730(.dina(n20027), .dinb(n19381), .dout(n20030));
  jnot g19731(.din(n20030), .dout(n20031));
  jand g19732(.dina(n20031), .dinb(n20029), .dout(n20032));
  jnot g19733(.din(n20032), .dout(n20033));
  jor  g19734(.dina(n20033), .dinb(n20025), .dout(n20034));
  jand g19735(.dina(n20034), .dinb(n20024), .dout(n20035));
  jor  g19736(.dina(n20035), .dinb(n2010), .dout(n20036));
  jand g19737(.dina(n20024), .dinb(n2010), .dout(n20037));
  jand g19738(.dina(n20037), .dinb(n20034), .dout(n20038));
  jnot g19739(.din(n19383), .dout(n20039));
  jand g19740(.dina(asqrt[3] ), .dinb(n20039), .dout(n20040));
  jand g19741(.dina(n20040), .dinb(n19390), .dout(n20041));
  jor  g19742(.dina(n20041), .dinb(n19388), .dout(n20042));
  jand g19743(.dina(n20040), .dinb(n19391), .dout(n20043));
  jnot g19744(.din(n20043), .dout(n20044));
  jand g19745(.dina(n20044), .dinb(n20042), .dout(n20045));
  jnot g19746(.din(n20045), .dout(n20046));
  jor  g19747(.dina(n20046), .dinb(n20038), .dout(n20047));
  jand g19748(.dina(n20047), .dinb(n20036), .dout(n20048));
  jor  g19749(.dina(n20048), .dinb(n2005), .dout(n20049));
  jxor g19750(.dina(n19392), .dinb(n2010), .dout(n20050));
  jor  g19751(.dina(n20050), .dinb(n19616), .dout(n20051));
  jxor g19752(.dina(n20051), .dinb(n19403), .dout(n20052));
  jand g19753(.dina(n20048), .dinb(n2005), .dout(n20053));
  jor  g19754(.dina(n20053), .dinb(n20052), .dout(n20054));
  jand g19755(.dina(n20054), .dinb(n20049), .dout(n20055));
  jor  g19756(.dina(n20055), .dinb(n1646), .dout(n20056));
  jnot g19757(.din(n19408), .dout(n20057));
  jor  g19758(.dina(n20057), .dinb(n19406), .dout(n20058));
  jor  g19759(.dina(n20058), .dinb(n19616), .dout(n20059));
  jxor g19760(.dina(n20059), .dinb(n19417), .dout(n20060));
  jand g19761(.dina(n20049), .dinb(n1646), .dout(n20061));
  jand g19762(.dina(n20061), .dinb(n20054), .dout(n20062));
  jor  g19763(.dina(n20062), .dinb(n20060), .dout(n20063));
  jand g19764(.dina(n20063), .dinb(n20056), .dout(n20064));
  jor  g19765(.dina(n20064), .dinb(n1641), .dout(n20065));
  jand g19766(.dina(n20064), .dinb(n1641), .dout(n20066));
  jnot g19767(.din(n19420), .dout(n20067));
  jand g19768(.dina(asqrt[3] ), .dinb(n20067), .dout(n20068));
  jand g19769(.dina(n20068), .dinb(n19425), .dout(n20069));
  jor  g19770(.dina(n20069), .dinb(n19424), .dout(n20070));
  jand g19771(.dina(n20068), .dinb(n19426), .dout(n20071));
  jnot g19772(.din(n20071), .dout(n20072));
  jand g19773(.dina(n20072), .dinb(n20070), .dout(n20073));
  jnot g19774(.din(n20073), .dout(n20074));
  jor  g19775(.dina(n20074), .dinb(n20066), .dout(n20075));
  jand g19776(.dina(n20075), .dinb(n20065), .dout(n20076));
  jor  g19777(.dina(n20076), .dinb(n1317), .dout(n20077));
  jand g19778(.dina(n20065), .dinb(n1317), .dout(n20078));
  jand g19779(.dina(n20078), .dinb(n20075), .dout(n20079));
  jnot g19780(.din(n19428), .dout(n20080));
  jand g19781(.dina(asqrt[3] ), .dinb(n20080), .dout(n20081));
  jand g19782(.dina(n20081), .dinb(n19435), .dout(n20082));
  jor  g19783(.dina(n20082), .dinb(n19433), .dout(n20083));
  jand g19784(.dina(n20081), .dinb(n19436), .dout(n20084));
  jnot g19785(.din(n20084), .dout(n20085));
  jand g19786(.dina(n20085), .dinb(n20083), .dout(n20086));
  jnot g19787(.din(n20086), .dout(n20087));
  jor  g19788(.dina(n20087), .dinb(n20079), .dout(n20088));
  jand g19789(.dina(n20088), .dinb(n20077), .dout(n20089));
  jor  g19790(.dina(n20089), .dinb(n1312), .dout(n20090));
  jxor g19791(.dina(n19437), .dinb(n1317), .dout(n20091));
  jor  g19792(.dina(n20091), .dinb(n19616), .dout(n20092));
  jxor g19793(.dina(n20092), .dinb(n19448), .dout(n20093));
  jand g19794(.dina(n20089), .dinb(n1312), .dout(n20094));
  jor  g19795(.dina(n20094), .dinb(n20093), .dout(n20095));
  jand g19796(.dina(n20095), .dinb(n20090), .dout(n20096));
  jor  g19797(.dina(n20096), .dinb(n1039), .dout(n20097));
  jnot g19798(.din(n19453), .dout(n20098));
  jor  g19799(.dina(n20098), .dinb(n19451), .dout(n20099));
  jor  g19800(.dina(n20099), .dinb(n19616), .dout(n20100));
  jxor g19801(.dina(n20100), .dinb(n19462), .dout(n20101));
  jand g19802(.dina(n20090), .dinb(n1039), .dout(n20102));
  jand g19803(.dina(n20102), .dinb(n20095), .dout(n20103));
  jor  g19804(.dina(n20103), .dinb(n20101), .dout(n20104));
  jand g19805(.dina(n20104), .dinb(n20097), .dout(n20105));
  jor  g19806(.dina(n20105), .dinb(n1034), .dout(n20106));
  jand g19807(.dina(n20105), .dinb(n1034), .dout(n20107));
  jnot g19808(.din(n19465), .dout(n20108));
  jand g19809(.dina(asqrt[3] ), .dinb(n20108), .dout(n20109));
  jand g19810(.dina(n20109), .dinb(n19470), .dout(n20110));
  jor  g19811(.dina(n20110), .dinb(n19469), .dout(n20111));
  jand g19812(.dina(n20109), .dinb(n19471), .dout(n20112));
  jnot g19813(.din(n20112), .dout(n20113));
  jand g19814(.dina(n20113), .dinb(n20111), .dout(n20114));
  jnot g19815(.din(n20114), .dout(n20115));
  jor  g19816(.dina(n20115), .dinb(n20107), .dout(n20116));
  jand g19817(.dina(n20116), .dinb(n20106), .dout(n20117));
  jor  g19818(.dina(n20117), .dinb(n796), .dout(n20118));
  jand g19819(.dina(n20106), .dinb(n796), .dout(n20119));
  jand g19820(.dina(n20119), .dinb(n20116), .dout(n20120));
  jnot g19821(.din(n19473), .dout(n20121));
  jand g19822(.dina(asqrt[3] ), .dinb(n20121), .dout(n20122));
  jand g19823(.dina(n20122), .dinb(n19480), .dout(n20123));
  jor  g19824(.dina(n20123), .dinb(n19478), .dout(n20124));
  jand g19825(.dina(n20122), .dinb(n19481), .dout(n20125));
  jnot g19826(.din(n20125), .dout(n20126));
  jand g19827(.dina(n20126), .dinb(n20124), .dout(n20127));
  jnot g19828(.din(n20127), .dout(n20128));
  jor  g19829(.dina(n20128), .dinb(n20120), .dout(n20129));
  jand g19830(.dina(n20129), .dinb(n20118), .dout(n20130));
  jor  g19831(.dina(n20130), .dinb(n791), .dout(n20131));
  jxor g19832(.dina(n19482), .dinb(n796), .dout(n20132));
  jor  g19833(.dina(n20132), .dinb(n19616), .dout(n20133));
  jxor g19834(.dina(n20133), .dinb(n19493), .dout(n20134));
  jand g19835(.dina(n20130), .dinb(n791), .dout(n20135));
  jor  g19836(.dina(n20135), .dinb(n20134), .dout(n20136));
  jand g19837(.dina(n20136), .dinb(n20131), .dout(n20137));
  jor  g19838(.dina(n20137), .dinb(n595), .dout(n20138));
  jnot g19839(.din(n19498), .dout(n20139));
  jor  g19840(.dina(n20139), .dinb(n19496), .dout(n20140));
  jor  g19841(.dina(n20140), .dinb(n19616), .dout(n20141));
  jxor g19842(.dina(n20141), .dinb(n19507), .dout(n20142));
  jand g19843(.dina(n20131), .dinb(n595), .dout(n20143));
  jand g19844(.dina(n20143), .dinb(n20136), .dout(n20144));
  jor  g19845(.dina(n20144), .dinb(n20142), .dout(n20145));
  jand g19846(.dina(n20145), .dinb(n20138), .dout(n20146));
  jor  g19847(.dina(n20146), .dinb(n590), .dout(n20147));
  jand g19848(.dina(n20146), .dinb(n590), .dout(n20148));
  jnot g19849(.din(n19510), .dout(n20149));
  jand g19850(.dina(asqrt[3] ), .dinb(n20149), .dout(n20150));
  jand g19851(.dina(n20150), .dinb(n19515), .dout(n20151));
  jor  g19852(.dina(n20151), .dinb(n19514), .dout(n20152));
  jand g19853(.dina(n20150), .dinb(n19516), .dout(n20153));
  jnot g19854(.din(n20153), .dout(n20154));
  jand g19855(.dina(n20154), .dinb(n20152), .dout(n20155));
  jnot g19856(.din(n20155), .dout(n20156));
  jor  g19857(.dina(n20156), .dinb(n20148), .dout(n20157));
  jand g19858(.dina(n20157), .dinb(n20147), .dout(n20158));
  jor  g19859(.dina(n20158), .dinb(n430), .dout(n20159));
  jand g19860(.dina(n20147), .dinb(n430), .dout(n20160));
  jand g19861(.dina(n20160), .dinb(n20157), .dout(n20161));
  jnot g19862(.din(n19518), .dout(n20162));
  jand g19863(.dina(asqrt[3] ), .dinb(n20162), .dout(n20163));
  jand g19864(.dina(n20163), .dinb(n19525), .dout(n20164));
  jor  g19865(.dina(n20164), .dinb(n19523), .dout(n20165));
  jand g19866(.dina(n20163), .dinb(n19526), .dout(n20166));
  jnot g19867(.din(n20166), .dout(n20167));
  jand g19868(.dina(n20167), .dinb(n20165), .dout(n20168));
  jnot g19869(.din(n20168), .dout(n20169));
  jor  g19870(.dina(n20169), .dinb(n20161), .dout(n20170));
  jand g19871(.dina(n20170), .dinb(n20159), .dout(n20171));
  jor  g19872(.dina(n20171), .dinb(n425), .dout(n20172));
  jxor g19873(.dina(n19527), .dinb(n430), .dout(n20173));
  jor  g19874(.dina(n20173), .dinb(n19616), .dout(n20174));
  jxor g19875(.dina(n20174), .dinb(n19538), .dout(n20175));
  jand g19876(.dina(n20171), .dinb(n425), .dout(n20176));
  jor  g19877(.dina(n20176), .dinb(n20175), .dout(n20177));
  jand g19878(.dina(n20177), .dinb(n20172), .dout(n20178));
  jor  g19879(.dina(n20178), .dinb(n305), .dout(n20179));
  jand g19880(.dina(n20172), .dinb(n305), .dout(n20180));
  jand g19881(.dina(n20180), .dinb(n20177), .dout(n20181));
  jnot g19882(.din(n19541), .dout(n20182));
  jand g19883(.dina(asqrt[3] ), .dinb(n20182), .dout(n20183));
  jand g19884(.dina(n20183), .dinb(n19548), .dout(n20184));
  jor  g19885(.dina(n20184), .dinb(n19546), .dout(n20185));
  jand g19886(.dina(n20183), .dinb(n19549), .dout(n20186));
  jnot g19887(.din(n20186), .dout(n20187));
  jand g19888(.dina(n20187), .dinb(n20185), .dout(n20188));
  jnot g19889(.din(n20188), .dout(n20189));
  jor  g19890(.dina(n20189), .dinb(n20181), .dout(n20190));
  jand g19891(.dina(n20190), .dinb(n20179), .dout(n20191));
  jor  g19892(.dina(n20191), .dinb(n290), .dout(n20192));
  jand g19893(.dina(n20191), .dinb(n290), .dout(n20193));
  jor  g19894(.dina(n20193), .dinb(n19620), .dout(n20194));
  jand g19895(.dina(n20194), .dinb(n20192), .dout(n20195));
  jor  g19896(.dina(n20195), .dinb(n223), .dout(n20196));
  jnot g19897(.din(n19557), .dout(n20197));
  jor  g19898(.dina(n20197), .dinb(n19555), .dout(n20198));
  jor  g19899(.dina(n20198), .dinb(n19616), .dout(n20199));
  jxor g19900(.dina(n20199), .dinb(n19566), .dout(n20200));
  jand g19901(.dina(n20192), .dinb(n223), .dout(n20201));
  jand g19902(.dina(n20201), .dinb(n20194), .dout(n20202));
  jor  g19903(.dina(n20202), .dinb(n20200), .dout(n20203));
  jand g19904(.dina(n20203), .dinb(n20196), .dout(n20204));
  jor  g19905(.dina(n20204), .dinb(n199), .dout(n20205));
  jand g19906(.dina(n20204), .dinb(n199), .dout(n20206));
  jxor g19907(.dina(n19568), .dinb(n223), .dout(n20207));
  jor  g19908(.dina(n20207), .dinb(n19616), .dout(n20208));
  jxor g19909(.dina(n20208), .dinb(n19579), .dout(n20209));
  jor  g19910(.dina(n20209), .dinb(n20206), .dout(n20210));
  jand g19911(.dina(n20210), .dinb(n20205), .dout(n20211));
  jnot g19912(.din(n19584), .dout(n20212));
  jor  g19913(.dina(n20212), .dinb(n19582), .dout(n20213));
  jor  g19914(.dina(n20213), .dinb(n19616), .dout(n20214));
  jxor g19915(.dina(n20214), .dinb(n19593), .dout(n20215));
  jnot g19916(.din(n19608), .dout(n20216));
  jand g19917(.dina(asqrt[3] ), .dinb(n19607), .dout(n20217));
  jand g19918(.dina(n20217), .dinb(n19595), .dout(n20218));
  jor  g19919(.dina(n20218), .dinb(n20216), .dout(n20219));
  jor  g19920(.dina(n20219), .dinb(n20215), .dout(n20220));
  jor  g19921(.dina(n20220), .dinb(n20211), .dout(n20221));
  jand g19922(.dina(n20221), .dinb(n194), .dout(n20222));
  jand g19923(.dina(n20215), .dinb(n20211), .dout(n20223));
  jor  g19924(.dina(n20217), .dinb(n19595), .dout(n20224));
  jand g19925(.dina(n19607), .dinb(n19595), .dout(n20225));
  jor  g19926(.dina(n20225), .dinb(n194), .dout(n20226));
  jnot g19927(.din(n20226), .dout(n20227));
  jand g19928(.dina(n20227), .dinb(n20224), .dout(n20228));
  jor  g19929(.dina(n20228), .dinb(n20223), .dout(n20229));
  jor  g19930(.dina(n20229), .dinb(n20222), .dout(asqrt[2] ));
  jxor g19931(.dina(n20191), .dinb(n290), .dout(n20231));
  jand g19932(.dina(n20231), .dinb(asqrt[2] ), .dout(n20232));
  jxor g19933(.dina(n20232), .dinb(n19620), .dout(n20233));
  jnot g19934(.din(n20233), .dout(n20234));
  jand g19935(.dina(asqrt[2] ), .dinb(a[4] ), .dout(n20235));
  jnot g19936(.din(a[2] ), .dout(n20236));
  jnot g19937(.din(a[3] ), .dout(n20237));
  jand g19938(.dina(n19622), .dinb(n20237), .dout(n20238));
  jand g19939(.dina(n20238), .dinb(n20236), .dout(n20239));
  jor  g19940(.dina(n20239), .dinb(n20235), .dout(n20240));
  jand g19941(.dina(n20240), .dinb(asqrt[3] ), .dout(n20241));
  jand g19942(.dina(asqrt[2] ), .dinb(n19622), .dout(n20242));
  jxor g19943(.dina(n20242), .dinb(n19623), .dout(n20243));
  jor  g19944(.dina(n20240), .dinb(asqrt[3] ), .dout(n20244));
  jand g19945(.dina(n20244), .dinb(n20243), .dout(n20245));
  jor  g19946(.dina(n20245), .dinb(n20241), .dout(n20246));
  jand g19947(.dina(n20246), .dinb(asqrt[4] ), .dout(n20247));
  jor  g19948(.dina(n20241), .dinb(asqrt[4] ), .dout(n20248));
  jor  g19949(.dina(n20248), .dinb(n20245), .dout(n20249));
  jand g19950(.dina(n20242), .dinb(n19623), .dout(n20250));
  jnot g19951(.din(asqrt[2] ), .dout(n20251));
  jand g19952(.dina(n20251), .dinb(asqrt[3] ), .dout(n20252));
  jor  g19953(.dina(n20252), .dinb(n20250), .dout(n20253));
  jxor g19954(.dina(n20253), .dinb(n18961), .dout(n20254));
  jand g19955(.dina(n20254), .dinb(n20249), .dout(n20255));
  jor  g19956(.dina(n20255), .dinb(n20247), .dout(n20256));
  jand g19957(.dina(n20256), .dinb(asqrt[5] ), .dout(n20257));
  jor  g19958(.dina(n20256), .dinb(asqrt[5] ), .dout(n20258));
  jxor g19959(.dina(n19627), .dinb(n18976), .dout(n20259));
  jand g19960(.dina(n20259), .dinb(asqrt[2] ), .dout(n20260));
  jxor g19961(.dina(n20260), .dinb(n19630), .dout(n20261));
  jnot g19962(.din(n20261), .dout(n20262));
  jand g19963(.dina(n20262), .dinb(n20258), .dout(n20263));
  jor  g19964(.dina(n20263), .dinb(n20257), .dout(n20264));
  jand g19965(.dina(n20264), .dinb(asqrt[6] ), .dout(n20265));
  jnot g19966(.din(n19636), .dout(n20266));
  jand g19967(.dina(n20266), .dinb(n19634), .dout(n20267));
  jand g19968(.dina(n20267), .dinb(asqrt[2] ), .dout(n20268));
  jxor g19969(.dina(n20268), .dinb(n19641), .dout(n20269));
  jnot g19970(.din(n20269), .dout(n20270));
  jor  g19971(.dina(n20257), .dinb(asqrt[6] ), .dout(n20271));
  jor  g19972(.dina(n20271), .dinb(n20263), .dout(n20272));
  jand g19973(.dina(n20272), .dinb(n20270), .dout(n20273));
  jor  g19974(.dina(n20273), .dinb(n20265), .dout(n20274));
  jand g19975(.dina(n20274), .dinb(asqrt[7] ), .dout(n20275));
  jor  g19976(.dina(n20274), .dinb(asqrt[7] ), .dout(n20276));
  jnot g19977(.din(n19648), .dout(n20277));
  jxor g19978(.dina(n19643), .dinb(n18360), .dout(n20278));
  jand g19979(.dina(n20278), .dinb(asqrt[2] ), .dout(n20279));
  jxor g19980(.dina(n20279), .dinb(n20277), .dout(n20280));
  jand g19981(.dina(n20280), .dinb(n20276), .dout(n20281));
  jor  g19982(.dina(n20281), .dinb(n20275), .dout(n20282));
  jand g19983(.dina(n20282), .dinb(asqrt[8] ), .dout(n20283));
  jor  g19984(.dina(n20275), .dinb(asqrt[8] ), .dout(n20284));
  jor  g19985(.dina(n20284), .dinb(n20281), .dout(n20285));
  jnot g19986(.din(n19655), .dout(n20286));
  jnot g19987(.din(n19657), .dout(n20287));
  jand g19988(.dina(asqrt[2] ), .dinb(n19651), .dout(n20288));
  jand g19989(.dina(n20288), .dinb(n20287), .dout(n20289));
  jor  g19990(.dina(n20289), .dinb(n20286), .dout(n20290));
  jnot g19991(.din(n19658), .dout(n20291));
  jand g19992(.dina(n20288), .dinb(n20291), .dout(n20292));
  jnot g19993(.din(n20292), .dout(n20293));
  jand g19994(.dina(n20293), .dinb(n20290), .dout(n20294));
  jand g19995(.dina(n20294), .dinb(n20285), .dout(n20295));
  jor  g19996(.dina(n20295), .dinb(n20283), .dout(n20296));
  jand g19997(.dina(n20296), .dinb(asqrt[9] ), .dout(n20297));
  jor  g19998(.dina(n20296), .dinb(asqrt[9] ), .dout(n20298));
  jxor g19999(.dina(n19659), .dinb(n17135), .dout(n20299));
  jand g20000(.dina(n20299), .dinb(asqrt[2] ), .dout(n20300));
  jxor g20001(.dina(n20300), .dinb(n19664), .dout(n20301));
  jand g20002(.dina(n20301), .dinb(n20298), .dout(n20302));
  jor  g20003(.dina(n20302), .dinb(n20297), .dout(n20303));
  jand g20004(.dina(n20303), .dinb(asqrt[10] ), .dout(n20304));
  jnot g20005(.din(n19670), .dout(n20305));
  jand g20006(.dina(n20305), .dinb(n19668), .dout(n20306));
  jand g20007(.dina(n20306), .dinb(asqrt[2] ), .dout(n20307));
  jxor g20008(.dina(n20307), .dinb(n19678), .dout(n20308));
  jnot g20009(.din(n20308), .dout(n20309));
  jor  g20010(.dina(n20297), .dinb(asqrt[10] ), .dout(n20310));
  jor  g20011(.dina(n20310), .dinb(n20302), .dout(n20311));
  jand g20012(.dina(n20311), .dinb(n20309), .dout(n20312));
  jor  g20013(.dina(n20312), .dinb(n20304), .dout(n20313));
  jand g20014(.dina(n20313), .dinb(asqrt[11] ), .dout(n20314));
  jor  g20015(.dina(n20313), .dinb(asqrt[11] ), .dout(n20315));
  jxor g20016(.dina(n19680), .dinb(n15950), .dout(n20316));
  jand g20017(.dina(n20316), .dinb(asqrt[2] ), .dout(n20317));
  jxor g20018(.dina(n20317), .dinb(n19686), .dout(n20318));
  jand g20019(.dina(n20318), .dinb(n20315), .dout(n20319));
  jor  g20020(.dina(n20319), .dinb(n20314), .dout(n20320));
  jand g20021(.dina(n20320), .dinb(asqrt[12] ), .dout(n20321));
  jor  g20022(.dina(n20314), .dinb(asqrt[12] ), .dout(n20322));
  jor  g20023(.dina(n20322), .dinb(n20319), .dout(n20323));
  jnot g20024(.din(n19694), .dout(n20324));
  jnot g20025(.din(n19696), .dout(n20325));
  jand g20026(.dina(asqrt[2] ), .dinb(n19690), .dout(n20326));
  jand g20027(.dina(n20326), .dinb(n20325), .dout(n20327));
  jor  g20028(.dina(n20327), .dinb(n20324), .dout(n20328));
  jnot g20029(.din(n19697), .dout(n20329));
  jand g20030(.dina(n20326), .dinb(n20329), .dout(n20330));
  jnot g20031(.din(n20330), .dout(n20331));
  jand g20032(.dina(n20331), .dinb(n20328), .dout(n20332));
  jand g20033(.dina(n20332), .dinb(n20323), .dout(n20333));
  jor  g20034(.dina(n20333), .dinb(n20321), .dout(n20334));
  jand g20035(.dina(n20334), .dinb(asqrt[13] ), .dout(n20335));
  jxor g20036(.dina(n19698), .dinb(n14816), .dout(n20336));
  jand g20037(.dina(n20336), .dinb(asqrt[2] ), .dout(n20337));
  jxor g20038(.dina(n20337), .dinb(n19705), .dout(n20338));
  jnot g20039(.din(n20338), .dout(n20339));
  jor  g20040(.dina(n20334), .dinb(asqrt[13] ), .dout(n20340));
  jand g20041(.dina(n20340), .dinb(n20339), .dout(n20341));
  jor  g20042(.dina(n20341), .dinb(n20335), .dout(n20342));
  jand g20043(.dina(n20342), .dinb(asqrt[14] ), .dout(n20343));
  jnot g20044(.din(n19710), .dout(n20344));
  jand g20045(.dina(n20344), .dinb(n19708), .dout(n20345));
  jand g20046(.dina(n20345), .dinb(asqrt[2] ), .dout(n20346));
  jxor g20047(.dina(n20346), .dinb(n19718), .dout(n20347));
  jnot g20048(.din(n20347), .dout(n20348));
  jor  g20049(.dina(n20335), .dinb(asqrt[14] ), .dout(n20349));
  jor  g20050(.dina(n20349), .dinb(n20341), .dout(n20350));
  jand g20051(.dina(n20350), .dinb(n20348), .dout(n20351));
  jor  g20052(.dina(n20351), .dinb(n20343), .dout(n20352));
  jand g20053(.dina(n20352), .dinb(asqrt[15] ), .dout(n20353));
  jor  g20054(.dina(n20352), .dinb(asqrt[15] ), .dout(n20354));
  jnot g20055(.din(n19724), .dout(n20355));
  jnot g20056(.din(n19725), .dout(n20356));
  jand g20057(.dina(asqrt[2] ), .dinb(n19721), .dout(n20357));
  jand g20058(.dina(n20357), .dinb(n20356), .dout(n20358));
  jor  g20059(.dina(n20358), .dinb(n20355), .dout(n20359));
  jnot g20060(.din(n19726), .dout(n20360));
  jand g20061(.dina(n20357), .dinb(n20360), .dout(n20361));
  jnot g20062(.din(n20361), .dout(n20362));
  jand g20063(.dina(n20362), .dinb(n20359), .dout(n20363));
  jand g20064(.dina(n20363), .dinb(n20354), .dout(n20364));
  jor  g20065(.dina(n20364), .dinb(n20353), .dout(n20365));
  jand g20066(.dina(n20365), .dinb(asqrt[16] ), .dout(n20366));
  jor  g20067(.dina(n20353), .dinb(asqrt[16] ), .dout(n20367));
  jor  g20068(.dina(n20367), .dinb(n20364), .dout(n20368));
  jnot g20069(.din(n19732), .dout(n20369));
  jnot g20070(.din(n19734), .dout(n20370));
  jand g20071(.dina(asqrt[2] ), .dinb(n19728), .dout(n20371));
  jand g20072(.dina(n20371), .dinb(n20370), .dout(n20372));
  jor  g20073(.dina(n20372), .dinb(n20369), .dout(n20373));
  jnot g20074(.din(n19735), .dout(n20374));
  jand g20075(.dina(n20371), .dinb(n20374), .dout(n20375));
  jnot g20076(.din(n20375), .dout(n20376));
  jand g20077(.dina(n20376), .dinb(n20373), .dout(n20377));
  jand g20078(.dina(n20377), .dinb(n20368), .dout(n20378));
  jor  g20079(.dina(n20378), .dinb(n20366), .dout(n20379));
  jand g20080(.dina(n20379), .dinb(asqrt[17] ), .dout(n20380));
  jxor g20081(.dina(n19736), .dinb(n12670), .dout(n20381));
  jand g20082(.dina(n20381), .dinb(asqrt[2] ), .dout(n20382));
  jxor g20083(.dina(n20382), .dinb(n19746), .dout(n20383));
  jnot g20084(.din(n20383), .dout(n20384));
  jor  g20085(.dina(n20379), .dinb(asqrt[17] ), .dout(n20385));
  jand g20086(.dina(n20385), .dinb(n20384), .dout(n20386));
  jor  g20087(.dina(n20386), .dinb(n20380), .dout(n20387));
  jand g20088(.dina(n20387), .dinb(asqrt[18] ), .dout(n20388));
  jnot g20089(.din(n19751), .dout(n20389));
  jand g20090(.dina(n20389), .dinb(n19749), .dout(n20390));
  jand g20091(.dina(n20390), .dinb(asqrt[2] ), .dout(n20391));
  jxor g20092(.dina(n20391), .dinb(n19759), .dout(n20392));
  jnot g20093(.din(n20392), .dout(n20393));
  jor  g20094(.dina(n20380), .dinb(asqrt[18] ), .dout(n20394));
  jor  g20095(.dina(n20394), .dinb(n20386), .dout(n20395));
  jand g20096(.dina(n20395), .dinb(n20393), .dout(n20396));
  jor  g20097(.dina(n20396), .dinb(n20388), .dout(n20397));
  jand g20098(.dina(n20397), .dinb(asqrt[19] ), .dout(n20398));
  jor  g20099(.dina(n20397), .dinb(asqrt[19] ), .dout(n20399));
  jnot g20100(.din(n19765), .dout(n20400));
  jnot g20101(.din(n19766), .dout(n20401));
  jand g20102(.dina(asqrt[2] ), .dinb(n19762), .dout(n20402));
  jand g20103(.dina(n20402), .dinb(n20401), .dout(n20403));
  jor  g20104(.dina(n20403), .dinb(n20400), .dout(n20404));
  jnot g20105(.din(n19767), .dout(n20405));
  jand g20106(.dina(n20402), .dinb(n20405), .dout(n20406));
  jnot g20107(.din(n20406), .dout(n20407));
  jand g20108(.dina(n20407), .dinb(n20404), .dout(n20408));
  jand g20109(.dina(n20408), .dinb(n20399), .dout(n20409));
  jor  g20110(.dina(n20409), .dinb(n20398), .dout(n20410));
  jand g20111(.dina(n20410), .dinb(asqrt[20] ), .dout(n20411));
  jor  g20112(.dina(n20398), .dinb(asqrt[20] ), .dout(n20412));
  jor  g20113(.dina(n20412), .dinb(n20409), .dout(n20413));
  jnot g20114(.din(n19773), .dout(n20414));
  jnot g20115(.din(n19775), .dout(n20415));
  jand g20116(.dina(asqrt[2] ), .dinb(n19769), .dout(n20416));
  jand g20117(.dina(n20416), .dinb(n20415), .dout(n20417));
  jor  g20118(.dina(n20417), .dinb(n20414), .dout(n20418));
  jnot g20119(.din(n19776), .dout(n20419));
  jand g20120(.dina(n20416), .dinb(n20419), .dout(n20420));
  jnot g20121(.din(n20420), .dout(n20421));
  jand g20122(.dina(n20421), .dinb(n20418), .dout(n20422));
  jand g20123(.dina(n20422), .dinb(n20413), .dout(n20423));
  jor  g20124(.dina(n20423), .dinb(n20411), .dout(n20424));
  jand g20125(.dina(n20424), .dinb(asqrt[21] ), .dout(n20425));
  jxor g20126(.dina(n19777), .dinb(n10696), .dout(n20426));
  jand g20127(.dina(n20426), .dinb(asqrt[2] ), .dout(n20427));
  jxor g20128(.dina(n20427), .dinb(n19787), .dout(n20428));
  jnot g20129(.din(n20428), .dout(n20429));
  jor  g20130(.dina(n20424), .dinb(asqrt[21] ), .dout(n20430));
  jand g20131(.dina(n20430), .dinb(n20429), .dout(n20431));
  jor  g20132(.dina(n20431), .dinb(n20425), .dout(n20432));
  jand g20133(.dina(n20432), .dinb(asqrt[22] ), .dout(n20433));
  jnot g20134(.din(n19792), .dout(n20434));
  jand g20135(.dina(n20434), .dinb(n19790), .dout(n20435));
  jand g20136(.dina(n20435), .dinb(asqrt[2] ), .dout(n20436));
  jxor g20137(.dina(n20436), .dinb(n19800), .dout(n20437));
  jnot g20138(.din(n20437), .dout(n20438));
  jor  g20139(.dina(n20425), .dinb(asqrt[22] ), .dout(n20439));
  jor  g20140(.dina(n20439), .dinb(n20431), .dout(n20440));
  jand g20141(.dina(n20440), .dinb(n20438), .dout(n20441));
  jor  g20142(.dina(n20441), .dinb(n20433), .dout(n20442));
  jand g20143(.dina(n20442), .dinb(asqrt[23] ), .dout(n20443));
  jor  g20144(.dina(n20442), .dinb(asqrt[23] ), .dout(n20444));
  jnot g20145(.din(n19806), .dout(n20445));
  jnot g20146(.din(n19807), .dout(n20446));
  jand g20147(.dina(asqrt[2] ), .dinb(n19803), .dout(n20447));
  jand g20148(.dina(n20447), .dinb(n20446), .dout(n20448));
  jor  g20149(.dina(n20448), .dinb(n20445), .dout(n20449));
  jnot g20150(.din(n19808), .dout(n20450));
  jand g20151(.dina(n20447), .dinb(n20450), .dout(n20451));
  jnot g20152(.din(n20451), .dout(n20452));
  jand g20153(.dina(n20452), .dinb(n20449), .dout(n20453));
  jand g20154(.dina(n20453), .dinb(n20444), .dout(n20454));
  jor  g20155(.dina(n20454), .dinb(n20443), .dout(n20455));
  jand g20156(.dina(n20455), .dinb(asqrt[24] ), .dout(n20456));
  jor  g20157(.dina(n20443), .dinb(asqrt[24] ), .dout(n20457));
  jor  g20158(.dina(n20457), .dinb(n20454), .dout(n20458));
  jnot g20159(.din(n19814), .dout(n20459));
  jnot g20160(.din(n19816), .dout(n20460));
  jand g20161(.dina(asqrt[2] ), .dinb(n19810), .dout(n20461));
  jand g20162(.dina(n20461), .dinb(n20460), .dout(n20462));
  jor  g20163(.dina(n20462), .dinb(n20459), .dout(n20463));
  jnot g20164(.din(n19817), .dout(n20464));
  jand g20165(.dina(n20461), .dinb(n20464), .dout(n20465));
  jnot g20166(.din(n20465), .dout(n20466));
  jand g20167(.dina(n20466), .dinb(n20463), .dout(n20467));
  jand g20168(.dina(n20467), .dinb(n20458), .dout(n20468));
  jor  g20169(.dina(n20468), .dinb(n20456), .dout(n20469));
  jand g20170(.dina(n20469), .dinb(asqrt[25] ), .dout(n20470));
  jxor g20171(.dina(n19818), .dinb(n8893), .dout(n20471));
  jand g20172(.dina(n20471), .dinb(asqrt[2] ), .dout(n20472));
  jxor g20173(.dina(n20472), .dinb(n19828), .dout(n20473));
  jnot g20174(.din(n20473), .dout(n20474));
  jor  g20175(.dina(n20469), .dinb(asqrt[25] ), .dout(n20475));
  jand g20176(.dina(n20475), .dinb(n20474), .dout(n20476));
  jor  g20177(.dina(n20476), .dinb(n20470), .dout(n20477));
  jand g20178(.dina(n20477), .dinb(asqrt[26] ), .dout(n20478));
  jnot g20179(.din(n19833), .dout(n20479));
  jand g20180(.dina(n20479), .dinb(n19831), .dout(n20480));
  jand g20181(.dina(n20480), .dinb(asqrt[2] ), .dout(n20481));
  jxor g20182(.dina(n20481), .dinb(n19841), .dout(n20482));
  jnot g20183(.din(n20482), .dout(n20483));
  jor  g20184(.dina(n20470), .dinb(asqrt[26] ), .dout(n20484));
  jor  g20185(.dina(n20484), .dinb(n20476), .dout(n20485));
  jand g20186(.dina(n20485), .dinb(n20483), .dout(n20486));
  jor  g20187(.dina(n20486), .dinb(n20478), .dout(n20487));
  jand g20188(.dina(n20487), .dinb(asqrt[27] ), .dout(n20488));
  jor  g20189(.dina(n20487), .dinb(asqrt[27] ), .dout(n20489));
  jnot g20190(.din(n19847), .dout(n20490));
  jnot g20191(.din(n19848), .dout(n20491));
  jand g20192(.dina(asqrt[2] ), .dinb(n19844), .dout(n20492));
  jand g20193(.dina(n20492), .dinb(n20491), .dout(n20493));
  jor  g20194(.dina(n20493), .dinb(n20490), .dout(n20494));
  jnot g20195(.din(n19849), .dout(n20495));
  jand g20196(.dina(n20492), .dinb(n20495), .dout(n20496));
  jnot g20197(.din(n20496), .dout(n20497));
  jand g20198(.dina(n20497), .dinb(n20494), .dout(n20498));
  jand g20199(.dina(n20498), .dinb(n20489), .dout(n20499));
  jor  g20200(.dina(n20499), .dinb(n20488), .dout(n20500));
  jand g20201(.dina(n20500), .dinb(asqrt[28] ), .dout(n20501));
  jor  g20202(.dina(n20488), .dinb(asqrt[28] ), .dout(n20502));
  jor  g20203(.dina(n20502), .dinb(n20499), .dout(n20503));
  jnot g20204(.din(n19855), .dout(n20504));
  jnot g20205(.din(n19857), .dout(n20505));
  jand g20206(.dina(asqrt[2] ), .dinb(n19851), .dout(n20506));
  jand g20207(.dina(n20506), .dinb(n20505), .dout(n20507));
  jor  g20208(.dina(n20507), .dinb(n20504), .dout(n20508));
  jnot g20209(.din(n19858), .dout(n20509));
  jand g20210(.dina(n20506), .dinb(n20509), .dout(n20510));
  jnot g20211(.din(n20510), .dout(n20511));
  jand g20212(.dina(n20511), .dinb(n20508), .dout(n20512));
  jand g20213(.dina(n20512), .dinb(n20503), .dout(n20513));
  jor  g20214(.dina(n20513), .dinb(n20501), .dout(n20514));
  jand g20215(.dina(n20514), .dinb(asqrt[29] ), .dout(n20515));
  jxor g20216(.dina(n19859), .dinb(n7260), .dout(n20516));
  jand g20217(.dina(n20516), .dinb(asqrt[2] ), .dout(n20517));
  jxor g20218(.dina(n20517), .dinb(n19869), .dout(n20518));
  jnot g20219(.din(n20518), .dout(n20519));
  jor  g20220(.dina(n20514), .dinb(asqrt[29] ), .dout(n20520));
  jand g20221(.dina(n20520), .dinb(n20519), .dout(n20521));
  jor  g20222(.dina(n20521), .dinb(n20515), .dout(n20522));
  jand g20223(.dina(n20522), .dinb(asqrt[30] ), .dout(n20523));
  jnot g20224(.din(n19874), .dout(n20524));
  jand g20225(.dina(n20524), .dinb(n19872), .dout(n20525));
  jand g20226(.dina(n20525), .dinb(asqrt[2] ), .dout(n20526));
  jxor g20227(.dina(n20526), .dinb(n19882), .dout(n20527));
  jnot g20228(.din(n20527), .dout(n20528));
  jor  g20229(.dina(n20515), .dinb(asqrt[30] ), .dout(n20529));
  jor  g20230(.dina(n20529), .dinb(n20521), .dout(n20530));
  jand g20231(.dina(n20530), .dinb(n20528), .dout(n20531));
  jor  g20232(.dina(n20531), .dinb(n20523), .dout(n20532));
  jand g20233(.dina(n20532), .dinb(asqrt[31] ), .dout(n20533));
  jor  g20234(.dina(n20532), .dinb(asqrt[31] ), .dout(n20534));
  jnot g20235(.din(n19888), .dout(n20535));
  jnot g20236(.din(n19889), .dout(n20536));
  jand g20237(.dina(asqrt[2] ), .dinb(n19885), .dout(n20537));
  jand g20238(.dina(n20537), .dinb(n20536), .dout(n20538));
  jor  g20239(.dina(n20538), .dinb(n20535), .dout(n20539));
  jnot g20240(.din(n19890), .dout(n20540));
  jand g20241(.dina(n20537), .dinb(n20540), .dout(n20541));
  jnot g20242(.din(n20541), .dout(n20542));
  jand g20243(.dina(n20542), .dinb(n20539), .dout(n20543));
  jand g20244(.dina(n20543), .dinb(n20534), .dout(n20544));
  jor  g20245(.dina(n20544), .dinb(n20533), .dout(n20545));
  jand g20246(.dina(n20545), .dinb(asqrt[32] ), .dout(n20546));
  jor  g20247(.dina(n20533), .dinb(asqrt[32] ), .dout(n20547));
  jor  g20248(.dina(n20547), .dinb(n20544), .dout(n20548));
  jnot g20249(.din(n19896), .dout(n20549));
  jnot g20250(.din(n19898), .dout(n20550));
  jand g20251(.dina(asqrt[2] ), .dinb(n19892), .dout(n20551));
  jand g20252(.dina(n20551), .dinb(n20550), .dout(n20552));
  jor  g20253(.dina(n20552), .dinb(n20549), .dout(n20553));
  jnot g20254(.din(n19899), .dout(n20554));
  jand g20255(.dina(n20551), .dinb(n20554), .dout(n20555));
  jnot g20256(.din(n20555), .dout(n20556));
  jand g20257(.dina(n20556), .dinb(n20553), .dout(n20557));
  jand g20258(.dina(n20557), .dinb(n20548), .dout(n20558));
  jor  g20259(.dina(n20558), .dinb(n20546), .dout(n20559));
  jand g20260(.dina(n20559), .dinb(asqrt[33] ), .dout(n20560));
  jxor g20261(.dina(n19900), .dinb(n5788), .dout(n20561));
  jand g20262(.dina(n20561), .dinb(asqrt[2] ), .dout(n20562));
  jxor g20263(.dina(n20562), .dinb(n19910), .dout(n20563));
  jnot g20264(.din(n20563), .dout(n20564));
  jor  g20265(.dina(n20559), .dinb(asqrt[33] ), .dout(n20565));
  jand g20266(.dina(n20565), .dinb(n20564), .dout(n20566));
  jor  g20267(.dina(n20566), .dinb(n20560), .dout(n20567));
  jand g20268(.dina(n20567), .dinb(asqrt[34] ), .dout(n20568));
  jnot g20269(.din(n19915), .dout(n20569));
  jand g20270(.dina(n20569), .dinb(n19913), .dout(n20570));
  jand g20271(.dina(n20570), .dinb(asqrt[2] ), .dout(n20571));
  jxor g20272(.dina(n20571), .dinb(n19923), .dout(n20572));
  jnot g20273(.din(n20572), .dout(n20573));
  jor  g20274(.dina(n20560), .dinb(asqrt[34] ), .dout(n20574));
  jor  g20275(.dina(n20574), .dinb(n20566), .dout(n20575));
  jand g20276(.dina(n20575), .dinb(n20573), .dout(n20576));
  jor  g20277(.dina(n20576), .dinb(n20568), .dout(n20577));
  jand g20278(.dina(n20577), .dinb(asqrt[35] ), .dout(n20578));
  jor  g20279(.dina(n20577), .dinb(asqrt[35] ), .dout(n20579));
  jnot g20280(.din(n19929), .dout(n20580));
  jnot g20281(.din(n19930), .dout(n20581));
  jand g20282(.dina(asqrt[2] ), .dinb(n19926), .dout(n20582));
  jand g20283(.dina(n20582), .dinb(n20581), .dout(n20583));
  jor  g20284(.dina(n20583), .dinb(n20580), .dout(n20584));
  jnot g20285(.din(n19931), .dout(n20585));
  jand g20286(.dina(n20582), .dinb(n20585), .dout(n20586));
  jnot g20287(.din(n20586), .dout(n20587));
  jand g20288(.dina(n20587), .dinb(n20584), .dout(n20588));
  jand g20289(.dina(n20588), .dinb(n20579), .dout(n20589));
  jor  g20290(.dina(n20589), .dinb(n20578), .dout(n20590));
  jand g20291(.dina(n20590), .dinb(asqrt[36] ), .dout(n20591));
  jor  g20292(.dina(n20578), .dinb(asqrt[36] ), .dout(n20592));
  jor  g20293(.dina(n20592), .dinb(n20589), .dout(n20593));
  jnot g20294(.din(n19937), .dout(n20594));
  jnot g20295(.din(n19939), .dout(n20595));
  jand g20296(.dina(asqrt[2] ), .dinb(n19933), .dout(n20596));
  jand g20297(.dina(n20596), .dinb(n20595), .dout(n20597));
  jor  g20298(.dina(n20597), .dinb(n20594), .dout(n20598));
  jnot g20299(.din(n19940), .dout(n20599));
  jand g20300(.dina(n20596), .dinb(n20599), .dout(n20600));
  jnot g20301(.din(n20600), .dout(n20601));
  jand g20302(.dina(n20601), .dinb(n20598), .dout(n20602));
  jand g20303(.dina(n20602), .dinb(n20593), .dout(n20603));
  jor  g20304(.dina(n20603), .dinb(n20591), .dout(n20604));
  jand g20305(.dina(n20604), .dinb(asqrt[37] ), .dout(n20605));
  jxor g20306(.dina(n19941), .dinb(n4494), .dout(n20606));
  jand g20307(.dina(n20606), .dinb(asqrt[2] ), .dout(n20607));
  jxor g20308(.dina(n20607), .dinb(n19951), .dout(n20608));
  jnot g20309(.din(n20608), .dout(n20609));
  jor  g20310(.dina(n20604), .dinb(asqrt[37] ), .dout(n20610));
  jand g20311(.dina(n20610), .dinb(n20609), .dout(n20611));
  jor  g20312(.dina(n20611), .dinb(n20605), .dout(n20612));
  jand g20313(.dina(n20612), .dinb(asqrt[38] ), .dout(n20613));
  jnot g20314(.din(n19956), .dout(n20614));
  jand g20315(.dina(n20614), .dinb(n19954), .dout(n20615));
  jand g20316(.dina(n20615), .dinb(asqrt[2] ), .dout(n20616));
  jxor g20317(.dina(n20616), .dinb(n19964), .dout(n20617));
  jnot g20318(.din(n20617), .dout(n20618));
  jor  g20319(.dina(n20605), .dinb(asqrt[38] ), .dout(n20619));
  jor  g20320(.dina(n20619), .dinb(n20611), .dout(n20620));
  jand g20321(.dina(n20620), .dinb(n20618), .dout(n20621));
  jor  g20322(.dina(n20621), .dinb(n20613), .dout(n20622));
  jand g20323(.dina(n20622), .dinb(asqrt[39] ), .dout(n20623));
  jor  g20324(.dina(n20622), .dinb(asqrt[39] ), .dout(n20624));
  jnot g20325(.din(n19970), .dout(n20625));
  jnot g20326(.din(n19971), .dout(n20626));
  jand g20327(.dina(asqrt[2] ), .dinb(n19967), .dout(n20627));
  jand g20328(.dina(n20627), .dinb(n20626), .dout(n20628));
  jor  g20329(.dina(n20628), .dinb(n20625), .dout(n20629));
  jnot g20330(.din(n19972), .dout(n20630));
  jand g20331(.dina(n20627), .dinb(n20630), .dout(n20631));
  jnot g20332(.din(n20631), .dout(n20632));
  jand g20333(.dina(n20632), .dinb(n20629), .dout(n20633));
  jand g20334(.dina(n20633), .dinb(n20624), .dout(n20634));
  jor  g20335(.dina(n20634), .dinb(n20623), .dout(n20635));
  jand g20336(.dina(n20635), .dinb(asqrt[40] ), .dout(n20636));
  jor  g20337(.dina(n20623), .dinb(asqrt[40] ), .dout(n20637));
  jor  g20338(.dina(n20637), .dinb(n20634), .dout(n20638));
  jnot g20339(.din(n19978), .dout(n20639));
  jnot g20340(.din(n19980), .dout(n20640));
  jand g20341(.dina(asqrt[2] ), .dinb(n19974), .dout(n20641));
  jand g20342(.dina(n20641), .dinb(n20640), .dout(n20642));
  jor  g20343(.dina(n20642), .dinb(n20639), .dout(n20643));
  jnot g20344(.din(n19981), .dout(n20644));
  jand g20345(.dina(n20641), .dinb(n20644), .dout(n20645));
  jnot g20346(.din(n20645), .dout(n20646));
  jand g20347(.dina(n20646), .dinb(n20643), .dout(n20647));
  jand g20348(.dina(n20647), .dinb(n20638), .dout(n20648));
  jor  g20349(.dina(n20648), .dinb(n20636), .dout(n20649));
  jand g20350(.dina(n20649), .dinb(asqrt[41] ), .dout(n20650));
  jxor g20351(.dina(n19982), .dinb(n3371), .dout(n20651));
  jand g20352(.dina(n20651), .dinb(asqrt[2] ), .dout(n20652));
  jxor g20353(.dina(n20652), .dinb(n19992), .dout(n20653));
  jnot g20354(.din(n20653), .dout(n20654));
  jor  g20355(.dina(n20649), .dinb(asqrt[41] ), .dout(n20655));
  jand g20356(.dina(n20655), .dinb(n20654), .dout(n20656));
  jor  g20357(.dina(n20656), .dinb(n20650), .dout(n20657));
  jand g20358(.dina(n20657), .dinb(asqrt[42] ), .dout(n20658));
  jnot g20359(.din(n19997), .dout(n20659));
  jand g20360(.dina(n20659), .dinb(n19995), .dout(n20660));
  jand g20361(.dina(n20660), .dinb(asqrt[2] ), .dout(n20661));
  jxor g20362(.dina(n20661), .dinb(n20005), .dout(n20662));
  jnot g20363(.din(n20662), .dout(n20663));
  jor  g20364(.dina(n20650), .dinb(asqrt[42] ), .dout(n20664));
  jor  g20365(.dina(n20664), .dinb(n20656), .dout(n20665));
  jand g20366(.dina(n20665), .dinb(n20663), .dout(n20666));
  jor  g20367(.dina(n20666), .dinb(n20658), .dout(n20667));
  jand g20368(.dina(n20667), .dinb(asqrt[43] ), .dout(n20668));
  jor  g20369(.dina(n20667), .dinb(asqrt[43] ), .dout(n20669));
  jnot g20370(.din(n20011), .dout(n20670));
  jnot g20371(.din(n20012), .dout(n20671));
  jand g20372(.dina(asqrt[2] ), .dinb(n20008), .dout(n20672));
  jand g20373(.dina(n20672), .dinb(n20671), .dout(n20673));
  jor  g20374(.dina(n20673), .dinb(n20670), .dout(n20674));
  jnot g20375(.din(n20013), .dout(n20675));
  jand g20376(.dina(n20672), .dinb(n20675), .dout(n20676));
  jnot g20377(.din(n20676), .dout(n20677));
  jand g20378(.dina(n20677), .dinb(n20674), .dout(n20678));
  jand g20379(.dina(n20678), .dinb(n20669), .dout(n20679));
  jor  g20380(.dina(n20679), .dinb(n20668), .dout(n20680));
  jand g20381(.dina(n20680), .dinb(asqrt[44] ), .dout(n20681));
  jor  g20382(.dina(n20668), .dinb(asqrt[44] ), .dout(n20682));
  jor  g20383(.dina(n20682), .dinb(n20679), .dout(n20683));
  jnot g20384(.din(n20019), .dout(n20684));
  jnot g20385(.din(n20021), .dout(n20685));
  jand g20386(.dina(asqrt[2] ), .dinb(n20015), .dout(n20686));
  jand g20387(.dina(n20686), .dinb(n20685), .dout(n20687));
  jor  g20388(.dina(n20687), .dinb(n20684), .dout(n20688));
  jnot g20389(.din(n20022), .dout(n20689));
  jand g20390(.dina(n20686), .dinb(n20689), .dout(n20690));
  jnot g20391(.din(n20690), .dout(n20691));
  jand g20392(.dina(n20691), .dinb(n20688), .dout(n20692));
  jand g20393(.dina(n20692), .dinb(n20683), .dout(n20693));
  jor  g20394(.dina(n20693), .dinb(n20681), .dout(n20694));
  jand g20395(.dina(n20694), .dinb(asqrt[45] ), .dout(n20695));
  jxor g20396(.dina(n20023), .dinb(n2420), .dout(n20696));
  jand g20397(.dina(n20696), .dinb(asqrt[2] ), .dout(n20697));
  jxor g20398(.dina(n20697), .dinb(n20033), .dout(n20698));
  jnot g20399(.din(n20698), .dout(n20699));
  jor  g20400(.dina(n20694), .dinb(asqrt[45] ), .dout(n20700));
  jand g20401(.dina(n20700), .dinb(n20699), .dout(n20701));
  jor  g20402(.dina(n20701), .dinb(n20695), .dout(n20702));
  jand g20403(.dina(n20702), .dinb(asqrt[46] ), .dout(n20703));
  jnot g20404(.din(n20038), .dout(n20704));
  jand g20405(.dina(n20704), .dinb(n20036), .dout(n20705));
  jand g20406(.dina(n20705), .dinb(asqrt[2] ), .dout(n20706));
  jxor g20407(.dina(n20706), .dinb(n20046), .dout(n20707));
  jnot g20408(.din(n20707), .dout(n20708));
  jor  g20409(.dina(n20695), .dinb(asqrt[46] ), .dout(n20709));
  jor  g20410(.dina(n20709), .dinb(n20701), .dout(n20710));
  jand g20411(.dina(n20710), .dinb(n20708), .dout(n20711));
  jor  g20412(.dina(n20711), .dinb(n20703), .dout(n20712));
  jand g20413(.dina(n20712), .dinb(asqrt[47] ), .dout(n20713));
  jor  g20414(.dina(n20712), .dinb(asqrt[47] ), .dout(n20714));
  jnot g20415(.din(n20052), .dout(n20715));
  jnot g20416(.din(n20053), .dout(n20716));
  jand g20417(.dina(asqrt[2] ), .dinb(n20049), .dout(n20717));
  jand g20418(.dina(n20717), .dinb(n20716), .dout(n20718));
  jor  g20419(.dina(n20718), .dinb(n20715), .dout(n20719));
  jnot g20420(.din(n20054), .dout(n20720));
  jand g20421(.dina(n20717), .dinb(n20720), .dout(n20721));
  jnot g20422(.din(n20721), .dout(n20722));
  jand g20423(.dina(n20722), .dinb(n20719), .dout(n20723));
  jand g20424(.dina(n20723), .dinb(n20714), .dout(n20724));
  jor  g20425(.dina(n20724), .dinb(n20713), .dout(n20725));
  jand g20426(.dina(n20725), .dinb(asqrt[48] ), .dout(n20726));
  jor  g20427(.dina(n20713), .dinb(asqrt[48] ), .dout(n20727));
  jor  g20428(.dina(n20727), .dinb(n20724), .dout(n20728));
  jnot g20429(.din(n20060), .dout(n20729));
  jnot g20430(.din(n20062), .dout(n20730));
  jand g20431(.dina(asqrt[2] ), .dinb(n20056), .dout(n20731));
  jand g20432(.dina(n20731), .dinb(n20730), .dout(n20732));
  jor  g20433(.dina(n20732), .dinb(n20729), .dout(n20733));
  jnot g20434(.din(n20063), .dout(n20734));
  jand g20435(.dina(n20731), .dinb(n20734), .dout(n20735));
  jnot g20436(.din(n20735), .dout(n20736));
  jand g20437(.dina(n20736), .dinb(n20733), .dout(n20737));
  jand g20438(.dina(n20737), .dinb(n20728), .dout(n20738));
  jor  g20439(.dina(n20738), .dinb(n20726), .dout(n20739));
  jand g20440(.dina(n20739), .dinb(asqrt[49] ), .dout(n20740));
  jxor g20441(.dina(n20064), .dinb(n1641), .dout(n20741));
  jand g20442(.dina(n20741), .dinb(asqrt[2] ), .dout(n20742));
  jxor g20443(.dina(n20742), .dinb(n20074), .dout(n20743));
  jnot g20444(.din(n20743), .dout(n20744));
  jor  g20445(.dina(n20739), .dinb(asqrt[49] ), .dout(n20745));
  jand g20446(.dina(n20745), .dinb(n20744), .dout(n20746));
  jor  g20447(.dina(n20746), .dinb(n20740), .dout(n20747));
  jand g20448(.dina(n20747), .dinb(asqrt[50] ), .dout(n20748));
  jnot g20449(.din(n20079), .dout(n20749));
  jand g20450(.dina(n20749), .dinb(n20077), .dout(n20750));
  jand g20451(.dina(n20750), .dinb(asqrt[2] ), .dout(n20751));
  jxor g20452(.dina(n20751), .dinb(n20087), .dout(n20752));
  jnot g20453(.din(n20752), .dout(n20753));
  jor  g20454(.dina(n20740), .dinb(asqrt[50] ), .dout(n20754));
  jor  g20455(.dina(n20754), .dinb(n20746), .dout(n20755));
  jand g20456(.dina(n20755), .dinb(n20753), .dout(n20756));
  jor  g20457(.dina(n20756), .dinb(n20748), .dout(n20757));
  jand g20458(.dina(n20757), .dinb(asqrt[51] ), .dout(n20758));
  jor  g20459(.dina(n20757), .dinb(asqrt[51] ), .dout(n20759));
  jnot g20460(.din(n20093), .dout(n20760));
  jnot g20461(.din(n20094), .dout(n20761));
  jand g20462(.dina(asqrt[2] ), .dinb(n20090), .dout(n20762));
  jand g20463(.dina(n20762), .dinb(n20761), .dout(n20763));
  jor  g20464(.dina(n20763), .dinb(n20760), .dout(n20764));
  jnot g20465(.din(n20095), .dout(n20765));
  jand g20466(.dina(n20762), .dinb(n20765), .dout(n20766));
  jnot g20467(.din(n20766), .dout(n20767));
  jand g20468(.dina(n20767), .dinb(n20764), .dout(n20768));
  jand g20469(.dina(n20768), .dinb(n20759), .dout(n20769));
  jor  g20470(.dina(n20769), .dinb(n20758), .dout(n20770));
  jand g20471(.dina(n20770), .dinb(asqrt[52] ), .dout(n20771));
  jor  g20472(.dina(n20758), .dinb(asqrt[52] ), .dout(n20772));
  jor  g20473(.dina(n20772), .dinb(n20769), .dout(n20773));
  jnot g20474(.din(n20101), .dout(n20774));
  jnot g20475(.din(n20103), .dout(n20775));
  jand g20476(.dina(asqrt[2] ), .dinb(n20097), .dout(n20776));
  jand g20477(.dina(n20776), .dinb(n20775), .dout(n20777));
  jor  g20478(.dina(n20777), .dinb(n20774), .dout(n20778));
  jnot g20479(.din(n20104), .dout(n20779));
  jand g20480(.dina(n20776), .dinb(n20779), .dout(n20780));
  jnot g20481(.din(n20780), .dout(n20781));
  jand g20482(.dina(n20781), .dinb(n20778), .dout(n20782));
  jand g20483(.dina(n20782), .dinb(n20773), .dout(n20783));
  jor  g20484(.dina(n20783), .dinb(n20771), .dout(n20784));
  jand g20485(.dina(n20784), .dinb(asqrt[53] ), .dout(n20785));
  jxor g20486(.dina(n20105), .dinb(n1034), .dout(n20786));
  jand g20487(.dina(n20786), .dinb(asqrt[2] ), .dout(n20787));
  jxor g20488(.dina(n20787), .dinb(n20115), .dout(n20788));
  jnot g20489(.din(n20788), .dout(n20789));
  jor  g20490(.dina(n20784), .dinb(asqrt[53] ), .dout(n20790));
  jand g20491(.dina(n20790), .dinb(n20789), .dout(n20791));
  jor  g20492(.dina(n20791), .dinb(n20785), .dout(n20792));
  jand g20493(.dina(n20792), .dinb(asqrt[54] ), .dout(n20793));
  jnot g20494(.din(n20120), .dout(n20794));
  jand g20495(.dina(n20794), .dinb(n20118), .dout(n20795));
  jand g20496(.dina(n20795), .dinb(asqrt[2] ), .dout(n20796));
  jxor g20497(.dina(n20796), .dinb(n20128), .dout(n20797));
  jnot g20498(.din(n20797), .dout(n20798));
  jor  g20499(.dina(n20785), .dinb(asqrt[54] ), .dout(n20799));
  jor  g20500(.dina(n20799), .dinb(n20791), .dout(n20800));
  jand g20501(.dina(n20800), .dinb(n20798), .dout(n20801));
  jor  g20502(.dina(n20801), .dinb(n20793), .dout(n20802));
  jand g20503(.dina(n20802), .dinb(asqrt[55] ), .dout(n20803));
  jor  g20504(.dina(n20802), .dinb(asqrt[55] ), .dout(n20804));
  jnot g20505(.din(n20134), .dout(n20805));
  jnot g20506(.din(n20135), .dout(n20806));
  jand g20507(.dina(asqrt[2] ), .dinb(n20131), .dout(n20807));
  jand g20508(.dina(n20807), .dinb(n20806), .dout(n20808));
  jor  g20509(.dina(n20808), .dinb(n20805), .dout(n20809));
  jnot g20510(.din(n20136), .dout(n20810));
  jand g20511(.dina(n20807), .dinb(n20810), .dout(n20811));
  jnot g20512(.din(n20811), .dout(n20812));
  jand g20513(.dina(n20812), .dinb(n20809), .dout(n20813));
  jand g20514(.dina(n20813), .dinb(n20804), .dout(n20814));
  jor  g20515(.dina(n20814), .dinb(n20803), .dout(n20815));
  jand g20516(.dina(n20815), .dinb(asqrt[56] ), .dout(n20816));
  jor  g20517(.dina(n20803), .dinb(asqrt[56] ), .dout(n20817));
  jor  g20518(.dina(n20817), .dinb(n20814), .dout(n20818));
  jnot g20519(.din(n20142), .dout(n20819));
  jnot g20520(.din(n20144), .dout(n20820));
  jand g20521(.dina(asqrt[2] ), .dinb(n20138), .dout(n20821));
  jand g20522(.dina(n20821), .dinb(n20820), .dout(n20822));
  jor  g20523(.dina(n20822), .dinb(n20819), .dout(n20823));
  jnot g20524(.din(n20145), .dout(n20824));
  jand g20525(.dina(n20821), .dinb(n20824), .dout(n20825));
  jnot g20526(.din(n20825), .dout(n20826));
  jand g20527(.dina(n20826), .dinb(n20823), .dout(n20827));
  jand g20528(.dina(n20827), .dinb(n20818), .dout(n20828));
  jor  g20529(.dina(n20828), .dinb(n20816), .dout(n20829));
  jand g20530(.dina(n20829), .dinb(asqrt[57] ), .dout(n20830));
  jxor g20531(.dina(n20146), .dinb(n590), .dout(n20831));
  jand g20532(.dina(n20831), .dinb(asqrt[2] ), .dout(n20832));
  jxor g20533(.dina(n20832), .dinb(n20156), .dout(n20833));
  jnot g20534(.din(n20833), .dout(n20834));
  jor  g20535(.dina(n20829), .dinb(asqrt[57] ), .dout(n20835));
  jand g20536(.dina(n20835), .dinb(n20834), .dout(n20836));
  jor  g20537(.dina(n20836), .dinb(n20830), .dout(n20837));
  jand g20538(.dina(n20837), .dinb(asqrt[58] ), .dout(n20838));
  jnot g20539(.din(n20161), .dout(n20839));
  jand g20540(.dina(n20839), .dinb(n20159), .dout(n20840));
  jand g20541(.dina(n20840), .dinb(asqrt[2] ), .dout(n20841));
  jxor g20542(.dina(n20841), .dinb(n20169), .dout(n20842));
  jnot g20543(.din(n20842), .dout(n20843));
  jor  g20544(.dina(n20830), .dinb(asqrt[58] ), .dout(n20844));
  jor  g20545(.dina(n20844), .dinb(n20836), .dout(n20845));
  jand g20546(.dina(n20845), .dinb(n20843), .dout(n20846));
  jor  g20547(.dina(n20846), .dinb(n20838), .dout(n20847));
  jand g20548(.dina(n20847), .dinb(asqrt[59] ), .dout(n20848));
  jor  g20549(.dina(n20847), .dinb(asqrt[59] ), .dout(n20849));
  jnot g20550(.din(n20175), .dout(n20850));
  jnot g20551(.din(n20176), .dout(n20851));
  jand g20552(.dina(asqrt[2] ), .dinb(n20172), .dout(n20852));
  jand g20553(.dina(n20852), .dinb(n20851), .dout(n20853));
  jor  g20554(.dina(n20853), .dinb(n20850), .dout(n20854));
  jnot g20555(.din(n20177), .dout(n20855));
  jand g20556(.dina(n20852), .dinb(n20855), .dout(n20856));
  jnot g20557(.din(n20856), .dout(n20857));
  jand g20558(.dina(n20857), .dinb(n20854), .dout(n20858));
  jand g20559(.dina(n20858), .dinb(n20849), .dout(n20859));
  jor  g20560(.dina(n20859), .dinb(n20848), .dout(n20860));
  jand g20561(.dina(n20860), .dinb(asqrt[60] ), .dout(n20861));
  jnot g20562(.din(n20181), .dout(n20862));
  jand g20563(.dina(n20862), .dinb(n20179), .dout(n20863));
  jand g20564(.dina(n20863), .dinb(asqrt[2] ), .dout(n20864));
  jxor g20565(.dina(n20864), .dinb(n20189), .dout(n20865));
  jnot g20566(.din(n20865), .dout(n20866));
  jor  g20567(.dina(n20848), .dinb(asqrt[60] ), .dout(n20867));
  jor  g20568(.dina(n20867), .dinb(n20859), .dout(n20868));
  jand g20569(.dina(n20868), .dinb(n20866), .dout(n20869));
  jor  g20570(.dina(n20869), .dinb(n20861), .dout(n20870));
  jand g20571(.dina(n20870), .dinb(asqrt[61] ), .dout(n20871));
  jor  g20572(.dina(n20870), .dinb(asqrt[61] ), .dout(n20872));
  jand g20573(.dina(n20872), .dinb(n20234), .dout(n20873));
  jor  g20574(.dina(n20873), .dinb(n20871), .dout(n20874));
  jand g20575(.dina(n20874), .dinb(asqrt[62] ), .dout(n20875));
  jor  g20576(.dina(n20871), .dinb(asqrt[62] ), .dout(n20876));
  jor  g20577(.dina(n20876), .dinb(n20873), .dout(n20877));
  jnot g20578(.din(n20200), .dout(n20878));
  jnot g20579(.din(n20202), .dout(n20879));
  jand g20580(.dina(asqrt[2] ), .dinb(n20196), .dout(n20880));
  jand g20581(.dina(n20880), .dinb(n20879), .dout(n20881));
  jor  g20582(.dina(n20881), .dinb(n20878), .dout(n20882));
  jnot g20583(.din(n20203), .dout(n20883));
  jand g20584(.dina(n20880), .dinb(n20883), .dout(n20884));
  jnot g20585(.din(n20884), .dout(n20885));
  jand g20586(.dina(n20885), .dinb(n20882), .dout(n20886));
  jand g20587(.dina(n20886), .dinb(n20877), .dout(n20887));
  jor  g20588(.dina(n20887), .dinb(n20875), .dout(n20888));
  jxor g20589(.dina(n20204), .dinb(n199), .dout(n20889));
  jand g20590(.dina(n20889), .dinb(asqrt[2] ), .dout(n20890));
  jxor g20591(.dina(n20890), .dinb(n20209), .dout(n20891));
  jnot g20592(.din(n20211), .dout(n20892));
  jnot g20593(.din(n20215), .dout(n20893));
  jand g20594(.dina(asqrt[2] ), .dinb(n20893), .dout(n20894));
  jand g20595(.dina(n20894), .dinb(n20892), .dout(n20895));
  jor  g20596(.dina(n20895), .dinb(n20223), .dout(n20896));
  jor  g20597(.dina(n20896), .dinb(n20891), .dout(n20897));
  jnot g20598(.din(n20897), .dout(n20898));
  jand g20599(.dina(n20898), .dinb(n20888), .dout(n20899));
  jor  g20600(.dina(n20899), .dinb(asqrt[63] ), .dout(n20900));
  jnot g20601(.din(n20891), .dout(n20901));
  jor  g20602(.dina(n20901), .dinb(n20888), .dout(n20902));
  jor  g20603(.dina(n20894), .dinb(n20892), .dout(n20903));
  jand g20604(.dina(n20893), .dinb(n20892), .dout(n20904));
  jor  g20605(.dina(n20904), .dinb(n194), .dout(n20905));
  jnot g20606(.din(n20905), .dout(n20906));
  jand g20607(.dina(n20906), .dinb(n20903), .dout(n20907));
  jnot g20608(.din(n20907), .dout(n20908));
  jand g20609(.dina(n20908), .dinb(n20902), .dout(n20909));
  jand g20610(.dina(n20909), .dinb(n20900), .dout(n20910));
  jxor g20611(.dina(n20870), .dinb(n223), .dout(n20911));
  jor  g20612(.dina(n20911), .dinb(n20910), .dout(n20912));
  jxor g20613(.dina(n20912), .dinb(n20234), .dout(n20913));
  jor  g20614(.dina(n20913), .dinb(n199), .dout(n20914));
  jor  g20615(.dina(a[1] ), .dinb(a[0] ), .dout(n20915));
  jand g20616(.dina(n20915), .dinb(n20236), .dout(n20916));
  jand g20617(.dina(n20910), .dinb(a[2] ), .dout(n20917));
  jor  g20618(.dina(n20917), .dinb(n20916), .dout(n20918));
  jand g20619(.dina(n20918), .dinb(n20251), .dout(n20919));
  jor  g20620(.dina(n20918), .dinb(n20251), .dout(n20920));
  jor  g20621(.dina(n20910), .dinb(a[2] ), .dout(n20921));
  jxor g20622(.dina(n20921), .dinb(n20237), .dout(n20922));
  jand g20623(.dina(n20922), .dinb(n20920), .dout(n20923));
  jor  g20624(.dina(n20923), .dinb(n20919), .dout(n20924));
  jor  g20625(.dina(n20924), .dinb(n19616), .dout(n20925));
  jor  g20626(.dina(n20921), .dinb(a[3] ), .dout(n20926));
  jnot g20627(.din(n20910), .dout(asqrt[1] ));
  jor  g20628(.dina(asqrt[1] ), .dinb(n20251), .dout(n20928));
  jand g20629(.dina(n20928), .dinb(n20926), .dout(n20929));
  jxor g20630(.dina(n20929), .dinb(n19622), .dout(n20930));
  jand g20631(.dina(n20930), .dinb(n20925), .dout(n20931));
  jxor g20632(.dina(n20240), .dinb(n19616), .dout(n20932));
  jor  g20633(.dina(n20932), .dinb(n20910), .dout(n20933));
  jxor g20634(.dina(n20933), .dinb(n20243), .dout(n20934));
  jand g20635(.dina(n20934), .dinb(n18976), .dout(n20935));
  jand g20636(.dina(n20924), .dinb(n19616), .dout(n20936));
  jor  g20637(.dina(n20936), .dinb(n20935), .dout(n20937));
  jor  g20638(.dina(n20937), .dinb(n20931), .dout(n20938));
  jnot g20639(.din(n20249), .dout(n20939));
  jor  g20640(.dina(n20939), .dinb(n20247), .dout(n20940));
  jor  g20641(.dina(n20940), .dinb(n20910), .dout(n20941));
  jxor g20642(.dina(n20941), .dinb(n20254), .dout(n20942));
  jor  g20643(.dina(n20942), .dinb(n18356), .dout(n20943));
  jor  g20644(.dina(n20934), .dinb(n18976), .dout(n20944));
  jand g20645(.dina(n20944), .dinb(n20943), .dout(n20945));
  jand g20646(.dina(n20945), .dinb(n20938), .dout(n20946));
  jand g20647(.dina(n20942), .dinb(n18356), .dout(n20947));
  jxor g20648(.dina(n20256), .dinb(n18356), .dout(n20948));
  jor  g20649(.dina(n20948), .dinb(n20910), .dout(n20949));
  jxor g20650(.dina(n20949), .dinb(n20262), .dout(n20950));
  jand g20651(.dina(n20950), .dinb(n18360), .dout(n20951));
  jor  g20652(.dina(n20951), .dinb(n20947), .dout(n20952));
  jor  g20653(.dina(n20952), .dinb(n20946), .dout(n20953));
  jnot g20654(.din(n20272), .dout(n20954));
  jor  g20655(.dina(n20910), .dinb(n20265), .dout(n20955));
  jor  g20656(.dina(n20955), .dinb(n20954), .dout(n20956));
  jand g20657(.dina(n20956), .dinb(n20269), .dout(n20957));
  jnot g20658(.din(n20955), .dout(n20958));
  jand g20659(.dina(n20958), .dinb(n20273), .dout(n20959));
  jor  g20660(.dina(n20959), .dinb(n20957), .dout(n20960));
  jor  g20661(.dina(n20960), .dinb(n17140), .dout(n20961));
  jor  g20662(.dina(n20950), .dinb(n18360), .dout(n20962));
  jand g20663(.dina(n20962), .dinb(n20961), .dout(n20963));
  jand g20664(.dina(n20963), .dinb(n20953), .dout(n20964));
  jxor g20665(.dina(n20274), .dinb(n17140), .dout(n20965));
  jor  g20666(.dina(n20965), .dinb(n20910), .dout(n20966));
  jxor g20667(.dina(n20966), .dinb(n20280), .dout(n20967));
  jand g20668(.dina(n20967), .dinb(n17135), .dout(n20968));
  jand g20669(.dina(n20960), .dinb(n17140), .dout(n20969));
  jor  g20670(.dina(n20969), .dinb(n20968), .dout(n20970));
  jor  g20671(.dina(n20970), .dinb(n20964), .dout(n20971));
  jnot g20672(.din(n20285), .dout(n20972));
  jor  g20673(.dina(n20972), .dinb(n20283), .dout(n20973));
  jor  g20674(.dina(n20973), .dinb(n20910), .dout(n20974));
  jxor g20675(.dina(n20974), .dinb(n20294), .dout(n20975));
  jor  g20676(.dina(n20975), .dinb(n15955), .dout(n20976));
  jor  g20677(.dina(n20967), .dinb(n17135), .dout(n20977));
  jand g20678(.dina(n20977), .dinb(n20976), .dout(n20978));
  jand g20679(.dina(n20978), .dinb(n20971), .dout(n20979));
  jxor g20680(.dina(n20296), .dinb(n15955), .dout(n20980));
  jor  g20681(.dina(n20980), .dinb(n20910), .dout(n20981));
  jxor g20682(.dina(n20981), .dinb(n20301), .dout(n20982));
  jand g20683(.dina(n20982), .dinb(n15950), .dout(n20983));
  jand g20684(.dina(n20975), .dinb(n15955), .dout(n20984));
  jor  g20685(.dina(n20984), .dinb(n20983), .dout(n20985));
  jor  g20686(.dina(n20985), .dinb(n20979), .dout(n20986));
  jnot g20687(.din(n20311), .dout(n20987));
  jnot g20688(.din(n20304), .dout(n20988));
  jand g20689(.dina(asqrt[1] ), .dinb(n20988), .dout(n20989));
  jnot g20690(.din(n20989), .dout(n20990));
  jor  g20691(.dina(n20990), .dinb(n20987), .dout(n20991));
  jand g20692(.dina(n20991), .dinb(n20308), .dout(n20992));
  jand g20693(.dina(n20989), .dinb(n20312), .dout(n20993));
  jor  g20694(.dina(n20993), .dinb(n20992), .dout(n20994));
  jor  g20695(.dina(n20994), .dinb(n14821), .dout(n20995));
  jor  g20696(.dina(n20982), .dinb(n15950), .dout(n20996));
  jand g20697(.dina(n20996), .dinb(n20995), .dout(n20997));
  jand g20698(.dina(n20997), .dinb(n20986), .dout(n20998));
  jxor g20699(.dina(n20313), .dinb(n14821), .dout(n20999));
  jor  g20700(.dina(n20999), .dinb(n20910), .dout(n21000));
  jxor g20701(.dina(n21000), .dinb(n20318), .dout(n21001));
  jand g20702(.dina(n21001), .dinb(n14816), .dout(n21002));
  jand g20703(.dina(n20994), .dinb(n14821), .dout(n21003));
  jor  g20704(.dina(n21003), .dinb(n21002), .dout(n21004));
  jor  g20705(.dina(n21004), .dinb(n20998), .dout(n21005));
  jnot g20706(.din(n20323), .dout(n21006));
  jor  g20707(.dina(n21006), .dinb(n20321), .dout(n21007));
  jor  g20708(.dina(n21007), .dinb(n20910), .dout(n21008));
  jxor g20709(.dina(n21008), .dinb(n20332), .dout(n21009));
  jor  g20710(.dina(n21009), .dinb(n13723), .dout(n21010));
  jor  g20711(.dina(n21001), .dinb(n14816), .dout(n21011));
  jand g20712(.dina(n21011), .dinb(n21010), .dout(n21012));
  jand g20713(.dina(n21012), .dinb(n21005), .dout(n21013));
  jnot g20714(.din(n20340), .dout(n21014));
  jnot g20715(.din(n20335), .dout(n21015));
  jand g20716(.dina(asqrt[1] ), .dinb(n21015), .dout(n21016));
  jnot g20717(.din(n21016), .dout(n21017));
  jor  g20718(.dina(n21017), .dinb(n21014), .dout(n21018));
  jand g20719(.dina(n21018), .dinb(n20338), .dout(n21019));
  jand g20720(.dina(n21016), .dinb(n20341), .dout(n21020));
  jor  g20721(.dina(n21020), .dinb(n21019), .dout(n21021));
  jand g20722(.dina(n21021), .dinb(n13718), .dout(n21022));
  jand g20723(.dina(n21009), .dinb(n13723), .dout(n21023));
  jor  g20724(.dina(n21023), .dinb(n21022), .dout(n21024));
  jor  g20725(.dina(n21024), .dinb(n21013), .dout(n21025));
  jnot g20726(.din(n20350), .dout(n21026));
  jnot g20727(.din(n20343), .dout(n21027));
  jand g20728(.dina(asqrt[1] ), .dinb(n21027), .dout(n21028));
  jnot g20729(.din(n21028), .dout(n21029));
  jor  g20730(.dina(n21029), .dinb(n21026), .dout(n21030));
  jand g20731(.dina(n21030), .dinb(n20347), .dout(n21031));
  jand g20732(.dina(n21028), .dinb(n20351), .dout(n21032));
  jor  g20733(.dina(n21032), .dinb(n21031), .dout(n21033));
  jor  g20734(.dina(n21033), .dinb(n12675), .dout(n21034));
  jor  g20735(.dina(n21021), .dinb(n13718), .dout(n21035));
  jand g20736(.dina(n21035), .dinb(n21034), .dout(n21036));
  jand g20737(.dina(n21036), .dinb(n21025), .dout(n21037));
  jxor g20738(.dina(n20352), .dinb(n12675), .dout(n21038));
  jor  g20739(.dina(n21038), .dinb(n20910), .dout(n21039));
  jxor g20740(.dina(n21039), .dinb(n20363), .dout(n21040));
  jand g20741(.dina(n21040), .dinb(n12670), .dout(n21041));
  jand g20742(.dina(n21033), .dinb(n12675), .dout(n21042));
  jor  g20743(.dina(n21042), .dinb(n21041), .dout(n21043));
  jor  g20744(.dina(n21043), .dinb(n21037), .dout(n21044));
  jnot g20745(.din(n20368), .dout(n21045));
  jor  g20746(.dina(n21045), .dinb(n20366), .dout(n21046));
  jor  g20747(.dina(n21046), .dinb(n20910), .dout(n21047));
  jxor g20748(.dina(n21047), .dinb(n20377), .dout(n21048));
  jor  g20749(.dina(n21048), .dinb(n11662), .dout(n21049));
  jor  g20750(.dina(n21040), .dinb(n12670), .dout(n21050));
  jand g20751(.dina(n21050), .dinb(n21049), .dout(n21051));
  jand g20752(.dina(n21051), .dinb(n21044), .dout(n21052));
  jnot g20753(.din(n20385), .dout(n21053));
  jnot g20754(.din(n20380), .dout(n21054));
  jand g20755(.dina(asqrt[1] ), .dinb(n21054), .dout(n21055));
  jnot g20756(.din(n21055), .dout(n21056));
  jor  g20757(.dina(n21056), .dinb(n21053), .dout(n21057));
  jand g20758(.dina(n21057), .dinb(n20383), .dout(n21058));
  jand g20759(.dina(n21055), .dinb(n20386), .dout(n21059));
  jor  g20760(.dina(n21059), .dinb(n21058), .dout(n21060));
  jand g20761(.dina(n21060), .dinb(n11657), .dout(n21061));
  jand g20762(.dina(n21048), .dinb(n11662), .dout(n21062));
  jor  g20763(.dina(n21062), .dinb(n21061), .dout(n21063));
  jor  g20764(.dina(n21063), .dinb(n21052), .dout(n21064));
  jnot g20765(.din(n20395), .dout(n21065));
  jnot g20766(.din(n20388), .dout(n21066));
  jand g20767(.dina(asqrt[1] ), .dinb(n21066), .dout(n21067));
  jnot g20768(.din(n21067), .dout(n21068));
  jor  g20769(.dina(n21068), .dinb(n21065), .dout(n21069));
  jand g20770(.dina(n21069), .dinb(n20392), .dout(n21070));
  jand g20771(.dina(n21067), .dinb(n20396), .dout(n21071));
  jor  g20772(.dina(n21071), .dinb(n21070), .dout(n21072));
  jor  g20773(.dina(n21072), .dinb(n10701), .dout(n21073));
  jor  g20774(.dina(n21060), .dinb(n11657), .dout(n21074));
  jand g20775(.dina(n21074), .dinb(n21073), .dout(n21075));
  jand g20776(.dina(n21075), .dinb(n21064), .dout(n21076));
  jxor g20777(.dina(n20397), .dinb(n10701), .dout(n21077));
  jor  g20778(.dina(n21077), .dinb(n20910), .dout(n21078));
  jxor g20779(.dina(n21078), .dinb(n20408), .dout(n21079));
  jand g20780(.dina(n21079), .dinb(n10696), .dout(n21080));
  jand g20781(.dina(n21072), .dinb(n10701), .dout(n21081));
  jor  g20782(.dina(n21081), .dinb(n21080), .dout(n21082));
  jor  g20783(.dina(n21082), .dinb(n21076), .dout(n21083));
  jnot g20784(.din(n20413), .dout(n21084));
  jor  g20785(.dina(n21084), .dinb(n20411), .dout(n21085));
  jor  g20786(.dina(n21085), .dinb(n20910), .dout(n21086));
  jxor g20787(.dina(n21086), .dinb(n20422), .dout(n21087));
  jor  g20788(.dina(n21087), .dinb(n9774), .dout(n21088));
  jor  g20789(.dina(n21079), .dinb(n10696), .dout(n21089));
  jand g20790(.dina(n21089), .dinb(n21088), .dout(n21090));
  jand g20791(.dina(n21090), .dinb(n21083), .dout(n21091));
  jnot g20792(.din(n20430), .dout(n21092));
  jnot g20793(.din(n20425), .dout(n21093));
  jand g20794(.dina(asqrt[1] ), .dinb(n21093), .dout(n21094));
  jnot g20795(.din(n21094), .dout(n21095));
  jor  g20796(.dina(n21095), .dinb(n21092), .dout(n21096));
  jand g20797(.dina(n21096), .dinb(n20428), .dout(n21097));
  jand g20798(.dina(n21094), .dinb(n20431), .dout(n21098));
  jor  g20799(.dina(n21098), .dinb(n21097), .dout(n21099));
  jand g20800(.dina(n21099), .dinb(n9769), .dout(n21100));
  jand g20801(.dina(n21087), .dinb(n9774), .dout(n21101));
  jor  g20802(.dina(n21101), .dinb(n21100), .dout(n21102));
  jor  g20803(.dina(n21102), .dinb(n21091), .dout(n21103));
  jnot g20804(.din(n20440), .dout(n21104));
  jnot g20805(.din(n20433), .dout(n21105));
  jand g20806(.dina(asqrt[1] ), .dinb(n21105), .dout(n21106));
  jnot g20807(.din(n21106), .dout(n21107));
  jor  g20808(.dina(n21107), .dinb(n21104), .dout(n21108));
  jand g20809(.dina(n21108), .dinb(n20437), .dout(n21109));
  jand g20810(.dina(n21106), .dinb(n20441), .dout(n21110));
  jor  g20811(.dina(n21110), .dinb(n21109), .dout(n21111));
  jor  g20812(.dina(n21111), .dinb(n8898), .dout(n21112));
  jor  g20813(.dina(n21099), .dinb(n9769), .dout(n21113));
  jand g20814(.dina(n21113), .dinb(n21112), .dout(n21114));
  jand g20815(.dina(n21114), .dinb(n21103), .dout(n21115));
  jxor g20816(.dina(n20442), .dinb(n8898), .dout(n21116));
  jor  g20817(.dina(n21116), .dinb(n20910), .dout(n21117));
  jxor g20818(.dina(n21117), .dinb(n20453), .dout(n21118));
  jand g20819(.dina(n21118), .dinb(n8893), .dout(n21119));
  jand g20820(.dina(n21111), .dinb(n8898), .dout(n21120));
  jor  g20821(.dina(n21120), .dinb(n21119), .dout(n21121));
  jor  g20822(.dina(n21121), .dinb(n21115), .dout(n21122));
  jnot g20823(.din(n20458), .dout(n21123));
  jor  g20824(.dina(n21123), .dinb(n20456), .dout(n21124));
  jor  g20825(.dina(n21124), .dinb(n20910), .dout(n21125));
  jxor g20826(.dina(n21125), .dinb(n20467), .dout(n21126));
  jor  g20827(.dina(n21126), .dinb(n8058), .dout(n21127));
  jor  g20828(.dina(n21118), .dinb(n8893), .dout(n21128));
  jand g20829(.dina(n21128), .dinb(n21127), .dout(n21129));
  jand g20830(.dina(n21129), .dinb(n21122), .dout(n21130));
  jnot g20831(.din(n20475), .dout(n21131));
  jnot g20832(.din(n20470), .dout(n21132));
  jand g20833(.dina(asqrt[1] ), .dinb(n21132), .dout(n21133));
  jnot g20834(.din(n21133), .dout(n21134));
  jor  g20835(.dina(n21134), .dinb(n21131), .dout(n21135));
  jand g20836(.dina(n21135), .dinb(n20473), .dout(n21136));
  jand g20837(.dina(n21133), .dinb(n20476), .dout(n21137));
  jor  g20838(.dina(n21137), .dinb(n21136), .dout(n21138));
  jand g20839(.dina(n21138), .dinb(n8053), .dout(n21139));
  jand g20840(.dina(n21126), .dinb(n8058), .dout(n21140));
  jor  g20841(.dina(n21140), .dinb(n21139), .dout(n21141));
  jor  g20842(.dina(n21141), .dinb(n21130), .dout(n21142));
  jnot g20843(.din(n20485), .dout(n21143));
  jnot g20844(.din(n20478), .dout(n21144));
  jand g20845(.dina(asqrt[1] ), .dinb(n21144), .dout(n21145));
  jnot g20846(.din(n21145), .dout(n21146));
  jor  g20847(.dina(n21146), .dinb(n21143), .dout(n21147));
  jand g20848(.dina(n21147), .dinb(n20482), .dout(n21148));
  jand g20849(.dina(n21145), .dinb(n20486), .dout(n21149));
  jor  g20850(.dina(n21149), .dinb(n21148), .dout(n21150));
  jor  g20851(.dina(n21150), .dinb(n7265), .dout(n21151));
  jor  g20852(.dina(n21138), .dinb(n8053), .dout(n21152));
  jand g20853(.dina(n21152), .dinb(n21151), .dout(n21153));
  jand g20854(.dina(n21153), .dinb(n21142), .dout(n21154));
  jxor g20855(.dina(n20487), .dinb(n7265), .dout(n21155));
  jor  g20856(.dina(n21155), .dinb(n20910), .dout(n21156));
  jxor g20857(.dina(n21156), .dinb(n20498), .dout(n21157));
  jand g20858(.dina(n21157), .dinb(n7260), .dout(n21158));
  jand g20859(.dina(n21150), .dinb(n7265), .dout(n21159));
  jor  g20860(.dina(n21159), .dinb(n21158), .dout(n21160));
  jor  g20861(.dina(n21160), .dinb(n21154), .dout(n21161));
  jnot g20862(.din(n20503), .dout(n21162));
  jor  g20863(.dina(n21162), .dinb(n20501), .dout(n21163));
  jor  g20864(.dina(n21163), .dinb(n20910), .dout(n21164));
  jxor g20865(.dina(n21164), .dinb(n20512), .dout(n21165));
  jor  g20866(.dina(n21165), .dinb(n6505), .dout(n21166));
  jor  g20867(.dina(n21157), .dinb(n7260), .dout(n21167));
  jand g20868(.dina(n21167), .dinb(n21166), .dout(n21168));
  jand g20869(.dina(n21168), .dinb(n21161), .dout(n21169));
  jnot g20870(.din(n20520), .dout(n21170));
  jnot g20871(.din(n20515), .dout(n21171));
  jand g20872(.dina(asqrt[1] ), .dinb(n21171), .dout(n21172));
  jnot g20873(.din(n21172), .dout(n21173));
  jor  g20874(.dina(n21173), .dinb(n21170), .dout(n21174));
  jand g20875(.dina(n21174), .dinb(n20518), .dout(n21175));
  jand g20876(.dina(n21172), .dinb(n20521), .dout(n21176));
  jor  g20877(.dina(n21176), .dinb(n21175), .dout(n21177));
  jand g20878(.dina(n21177), .dinb(n6500), .dout(n21178));
  jand g20879(.dina(n21165), .dinb(n6505), .dout(n21179));
  jor  g20880(.dina(n21179), .dinb(n21178), .dout(n21180));
  jor  g20881(.dina(n21180), .dinb(n21169), .dout(n21181));
  jnot g20882(.din(n20530), .dout(n21182));
  jnot g20883(.din(n20523), .dout(n21183));
  jand g20884(.dina(asqrt[1] ), .dinb(n21183), .dout(n21184));
  jnot g20885(.din(n21184), .dout(n21185));
  jor  g20886(.dina(n21185), .dinb(n21182), .dout(n21186));
  jand g20887(.dina(n21186), .dinb(n20527), .dout(n21187));
  jand g20888(.dina(n21184), .dinb(n20531), .dout(n21188));
  jor  g20889(.dina(n21188), .dinb(n21187), .dout(n21189));
  jor  g20890(.dina(n21189), .dinb(n5793), .dout(n21190));
  jor  g20891(.dina(n21177), .dinb(n6500), .dout(n21191));
  jand g20892(.dina(n21191), .dinb(n21190), .dout(n21192));
  jand g20893(.dina(n21192), .dinb(n21181), .dout(n21193));
  jxor g20894(.dina(n20532), .dinb(n5793), .dout(n21194));
  jor  g20895(.dina(n21194), .dinb(n20910), .dout(n21195));
  jxor g20896(.dina(n21195), .dinb(n20543), .dout(n21196));
  jand g20897(.dina(n21196), .dinb(n5788), .dout(n21197));
  jand g20898(.dina(n21189), .dinb(n5793), .dout(n21198));
  jor  g20899(.dina(n21198), .dinb(n21197), .dout(n21199));
  jor  g20900(.dina(n21199), .dinb(n21193), .dout(n21200));
  jnot g20901(.din(n20548), .dout(n21201));
  jor  g20902(.dina(n21201), .dinb(n20546), .dout(n21202));
  jor  g20903(.dina(n21202), .dinb(n20910), .dout(n21203));
  jxor g20904(.dina(n21203), .dinb(n20557), .dout(n21204));
  jor  g20905(.dina(n21204), .dinb(n5121), .dout(n21205));
  jor  g20906(.dina(n21196), .dinb(n5788), .dout(n21206));
  jand g20907(.dina(n21206), .dinb(n21205), .dout(n21207));
  jand g20908(.dina(n21207), .dinb(n21200), .dout(n21208));
  jnot g20909(.din(n20565), .dout(n21209));
  jnot g20910(.din(n20560), .dout(n21210));
  jand g20911(.dina(asqrt[1] ), .dinb(n21210), .dout(n21211));
  jnot g20912(.din(n21211), .dout(n21212));
  jor  g20913(.dina(n21212), .dinb(n21209), .dout(n21213));
  jand g20914(.dina(n21213), .dinb(n20563), .dout(n21214));
  jand g20915(.dina(n21211), .dinb(n20566), .dout(n21215));
  jor  g20916(.dina(n21215), .dinb(n21214), .dout(n21216));
  jand g20917(.dina(n21216), .dinb(n5116), .dout(n21217));
  jand g20918(.dina(n21204), .dinb(n5121), .dout(n21218));
  jor  g20919(.dina(n21218), .dinb(n21217), .dout(n21219));
  jor  g20920(.dina(n21219), .dinb(n21208), .dout(n21220));
  jnot g20921(.din(n20575), .dout(n21221));
  jnot g20922(.din(n20568), .dout(n21222));
  jand g20923(.dina(asqrt[1] ), .dinb(n21222), .dout(n21223));
  jnot g20924(.din(n21223), .dout(n21224));
  jor  g20925(.dina(n21224), .dinb(n21221), .dout(n21225));
  jand g20926(.dina(n21225), .dinb(n20572), .dout(n21226));
  jand g20927(.dina(n21223), .dinb(n20576), .dout(n21227));
  jor  g20928(.dina(n21227), .dinb(n21226), .dout(n21228));
  jor  g20929(.dina(n21228), .dinb(n4499), .dout(n21229));
  jor  g20930(.dina(n21216), .dinb(n5116), .dout(n21230));
  jand g20931(.dina(n21230), .dinb(n21229), .dout(n21231));
  jand g20932(.dina(n21231), .dinb(n21220), .dout(n21232));
  jxor g20933(.dina(n20577), .dinb(n4499), .dout(n21233));
  jor  g20934(.dina(n21233), .dinb(n20910), .dout(n21234));
  jxor g20935(.dina(n21234), .dinb(n20588), .dout(n21235));
  jand g20936(.dina(n21235), .dinb(n4494), .dout(n21236));
  jand g20937(.dina(n21228), .dinb(n4499), .dout(n21237));
  jor  g20938(.dina(n21237), .dinb(n21236), .dout(n21238));
  jor  g20939(.dina(n21238), .dinb(n21232), .dout(n21239));
  jnot g20940(.din(n20593), .dout(n21240));
  jor  g20941(.dina(n21240), .dinb(n20591), .dout(n21241));
  jor  g20942(.dina(n21241), .dinb(n20910), .dout(n21242));
  jxor g20943(.dina(n21242), .dinb(n20602), .dout(n21243));
  jor  g20944(.dina(n21243), .dinb(n3912), .dout(n21244));
  jor  g20945(.dina(n21235), .dinb(n4494), .dout(n21245));
  jand g20946(.dina(n21245), .dinb(n21244), .dout(n21246));
  jand g20947(.dina(n21246), .dinb(n21239), .dout(n21247));
  jnot g20948(.din(n20610), .dout(n21248));
  jnot g20949(.din(n20605), .dout(n21249));
  jand g20950(.dina(asqrt[1] ), .dinb(n21249), .dout(n21250));
  jnot g20951(.din(n21250), .dout(n21251));
  jor  g20952(.dina(n21251), .dinb(n21248), .dout(n21252));
  jand g20953(.dina(n21252), .dinb(n20608), .dout(n21253));
  jand g20954(.dina(n21250), .dinb(n20611), .dout(n21254));
  jor  g20955(.dina(n21254), .dinb(n21253), .dout(n21255));
  jand g20956(.dina(n21255), .dinb(n3907), .dout(n21256));
  jand g20957(.dina(n21243), .dinb(n3912), .dout(n21257));
  jor  g20958(.dina(n21257), .dinb(n21256), .dout(n21258));
  jor  g20959(.dina(n21258), .dinb(n21247), .dout(n21259));
  jnot g20960(.din(n20620), .dout(n21260));
  jnot g20961(.din(n20613), .dout(n21261));
  jand g20962(.dina(asqrt[1] ), .dinb(n21261), .dout(n21262));
  jnot g20963(.din(n21262), .dout(n21263));
  jor  g20964(.dina(n21263), .dinb(n21260), .dout(n21264));
  jand g20965(.dina(n21264), .dinb(n20617), .dout(n21265));
  jand g20966(.dina(n21262), .dinb(n20621), .dout(n21266));
  jor  g20967(.dina(n21266), .dinb(n21265), .dout(n21267));
  jor  g20968(.dina(n21267), .dinb(n3376), .dout(n21268));
  jor  g20969(.dina(n21255), .dinb(n3907), .dout(n21269));
  jand g20970(.dina(n21269), .dinb(n21268), .dout(n21270));
  jand g20971(.dina(n21270), .dinb(n21259), .dout(n21271));
  jxor g20972(.dina(n20622), .dinb(n3376), .dout(n21272));
  jor  g20973(.dina(n21272), .dinb(n20910), .dout(n21273));
  jxor g20974(.dina(n21273), .dinb(n20633), .dout(n21274));
  jand g20975(.dina(n21274), .dinb(n3371), .dout(n21275));
  jand g20976(.dina(n21267), .dinb(n3376), .dout(n21276));
  jor  g20977(.dina(n21276), .dinb(n21275), .dout(n21277));
  jor  g20978(.dina(n21277), .dinb(n21271), .dout(n21278));
  jnot g20979(.din(n20638), .dout(n21279));
  jor  g20980(.dina(n21279), .dinb(n20636), .dout(n21280));
  jor  g20981(.dina(n21280), .dinb(n20910), .dout(n21281));
  jxor g20982(.dina(n21281), .dinb(n20647), .dout(n21282));
  jor  g20983(.dina(n21282), .dinb(n2875), .dout(n21283));
  jor  g20984(.dina(n21274), .dinb(n3371), .dout(n21284));
  jand g20985(.dina(n21284), .dinb(n21283), .dout(n21285));
  jand g20986(.dina(n21285), .dinb(n21278), .dout(n21286));
  jnot g20987(.din(n20655), .dout(n21287));
  jnot g20988(.din(n20650), .dout(n21288));
  jand g20989(.dina(asqrt[1] ), .dinb(n21288), .dout(n21289));
  jnot g20990(.din(n21289), .dout(n21290));
  jor  g20991(.dina(n21290), .dinb(n21287), .dout(n21291));
  jand g20992(.dina(n21291), .dinb(n20653), .dout(n21292));
  jand g20993(.dina(n21289), .dinb(n20656), .dout(n21293));
  jor  g20994(.dina(n21293), .dinb(n21292), .dout(n21294));
  jand g20995(.dina(n21294), .dinb(n2870), .dout(n21295));
  jand g20996(.dina(n21282), .dinb(n2875), .dout(n21296));
  jor  g20997(.dina(n21296), .dinb(n21295), .dout(n21297));
  jor  g20998(.dina(n21297), .dinb(n21286), .dout(n21298));
  jnot g20999(.din(n20665), .dout(n21299));
  jnot g21000(.din(n20658), .dout(n21300));
  jand g21001(.dina(asqrt[1] ), .dinb(n21300), .dout(n21301));
  jnot g21002(.din(n21301), .dout(n21302));
  jor  g21003(.dina(n21302), .dinb(n21299), .dout(n21303));
  jand g21004(.dina(n21303), .dinb(n20662), .dout(n21304));
  jand g21005(.dina(n21301), .dinb(n20666), .dout(n21305));
  jor  g21006(.dina(n21305), .dinb(n21304), .dout(n21306));
  jor  g21007(.dina(n21306), .dinb(n2425), .dout(n21307));
  jor  g21008(.dina(n21294), .dinb(n2870), .dout(n21308));
  jand g21009(.dina(n21308), .dinb(n21307), .dout(n21309));
  jand g21010(.dina(n21309), .dinb(n21298), .dout(n21310));
  jxor g21011(.dina(n20667), .dinb(n2425), .dout(n21311));
  jor  g21012(.dina(n21311), .dinb(n20910), .dout(n21312));
  jxor g21013(.dina(n21312), .dinb(n20678), .dout(n21313));
  jand g21014(.dina(n21313), .dinb(n2420), .dout(n21314));
  jand g21015(.dina(n21306), .dinb(n2425), .dout(n21315));
  jor  g21016(.dina(n21315), .dinb(n21314), .dout(n21316));
  jor  g21017(.dina(n21316), .dinb(n21310), .dout(n21317));
  jnot g21018(.din(n20683), .dout(n21318));
  jor  g21019(.dina(n21318), .dinb(n20681), .dout(n21319));
  jor  g21020(.dina(n21319), .dinb(n20910), .dout(n21320));
  jxor g21021(.dina(n21320), .dinb(n20692), .dout(n21321));
  jor  g21022(.dina(n21321), .dinb(n2010), .dout(n21322));
  jor  g21023(.dina(n21313), .dinb(n2420), .dout(n21323));
  jand g21024(.dina(n21323), .dinb(n21322), .dout(n21324));
  jand g21025(.dina(n21324), .dinb(n21317), .dout(n21325));
  jnot g21026(.din(n20700), .dout(n21326));
  jnot g21027(.din(n20695), .dout(n21327));
  jand g21028(.dina(asqrt[1] ), .dinb(n21327), .dout(n21328));
  jnot g21029(.din(n21328), .dout(n21329));
  jor  g21030(.dina(n21329), .dinb(n21326), .dout(n21330));
  jand g21031(.dina(n21330), .dinb(n20698), .dout(n21331));
  jand g21032(.dina(n21328), .dinb(n20701), .dout(n21332));
  jor  g21033(.dina(n21332), .dinb(n21331), .dout(n21333));
  jand g21034(.dina(n21333), .dinb(n2005), .dout(n21334));
  jand g21035(.dina(n21321), .dinb(n2010), .dout(n21335));
  jor  g21036(.dina(n21335), .dinb(n21334), .dout(n21336));
  jor  g21037(.dina(n21336), .dinb(n21325), .dout(n21337));
  jnot g21038(.din(n20710), .dout(n21338));
  jnot g21039(.din(n20703), .dout(n21339));
  jand g21040(.dina(asqrt[1] ), .dinb(n21339), .dout(n21340));
  jnot g21041(.din(n21340), .dout(n21341));
  jor  g21042(.dina(n21341), .dinb(n21338), .dout(n21342));
  jand g21043(.dina(n21342), .dinb(n20707), .dout(n21343));
  jand g21044(.dina(n21340), .dinb(n20711), .dout(n21344));
  jor  g21045(.dina(n21344), .dinb(n21343), .dout(n21345));
  jor  g21046(.dina(n21345), .dinb(n1646), .dout(n21346));
  jor  g21047(.dina(n21333), .dinb(n2005), .dout(n21347));
  jand g21048(.dina(n21347), .dinb(n21346), .dout(n21348));
  jand g21049(.dina(n21348), .dinb(n21337), .dout(n21349));
  jxor g21050(.dina(n20712), .dinb(n1646), .dout(n21350));
  jor  g21051(.dina(n21350), .dinb(n20910), .dout(n21351));
  jxor g21052(.dina(n21351), .dinb(n20723), .dout(n21352));
  jand g21053(.dina(n21352), .dinb(n1641), .dout(n21353));
  jand g21054(.dina(n21345), .dinb(n1646), .dout(n21354));
  jor  g21055(.dina(n21354), .dinb(n21353), .dout(n21355));
  jor  g21056(.dina(n21355), .dinb(n21349), .dout(n21356));
  jnot g21057(.din(n20728), .dout(n21357));
  jor  g21058(.dina(n21357), .dinb(n20726), .dout(n21358));
  jor  g21059(.dina(n21358), .dinb(n20910), .dout(n21359));
  jxor g21060(.dina(n21359), .dinb(n20737), .dout(n21360));
  jor  g21061(.dina(n21360), .dinb(n1317), .dout(n21361));
  jor  g21062(.dina(n21352), .dinb(n1641), .dout(n21362));
  jand g21063(.dina(n21362), .dinb(n21361), .dout(n21363));
  jand g21064(.dina(n21363), .dinb(n21356), .dout(n21364));
  jnot g21065(.din(n20745), .dout(n21365));
  jnot g21066(.din(n20740), .dout(n21366));
  jand g21067(.dina(asqrt[1] ), .dinb(n21366), .dout(n21367));
  jnot g21068(.din(n21367), .dout(n21368));
  jor  g21069(.dina(n21368), .dinb(n21365), .dout(n21369));
  jand g21070(.dina(n21369), .dinb(n20743), .dout(n21370));
  jand g21071(.dina(n21367), .dinb(n20746), .dout(n21371));
  jor  g21072(.dina(n21371), .dinb(n21370), .dout(n21372));
  jand g21073(.dina(n21372), .dinb(n1312), .dout(n21373));
  jand g21074(.dina(n21360), .dinb(n1317), .dout(n21374));
  jor  g21075(.dina(n21374), .dinb(n21373), .dout(n21375));
  jor  g21076(.dina(n21375), .dinb(n21364), .dout(n21376));
  jnot g21077(.din(n20755), .dout(n21377));
  jnot g21078(.din(n20748), .dout(n21378));
  jand g21079(.dina(asqrt[1] ), .dinb(n21378), .dout(n21379));
  jnot g21080(.din(n21379), .dout(n21380));
  jor  g21081(.dina(n21380), .dinb(n21377), .dout(n21381));
  jand g21082(.dina(n21381), .dinb(n20752), .dout(n21382));
  jand g21083(.dina(n21379), .dinb(n20756), .dout(n21383));
  jor  g21084(.dina(n21383), .dinb(n21382), .dout(n21384));
  jor  g21085(.dina(n21384), .dinb(n1039), .dout(n21385));
  jor  g21086(.dina(n21372), .dinb(n1312), .dout(n21386));
  jand g21087(.dina(n21386), .dinb(n21385), .dout(n21387));
  jand g21088(.dina(n21387), .dinb(n21376), .dout(n21388));
  jxor g21089(.dina(n20757), .dinb(n1039), .dout(n21389));
  jor  g21090(.dina(n21389), .dinb(n20910), .dout(n21390));
  jxor g21091(.dina(n21390), .dinb(n20768), .dout(n21391));
  jand g21092(.dina(n21391), .dinb(n1034), .dout(n21392));
  jand g21093(.dina(n21384), .dinb(n1039), .dout(n21393));
  jor  g21094(.dina(n21393), .dinb(n21392), .dout(n21394));
  jor  g21095(.dina(n21394), .dinb(n21388), .dout(n21395));
  jnot g21096(.din(n20773), .dout(n21396));
  jor  g21097(.dina(n21396), .dinb(n20771), .dout(n21397));
  jor  g21098(.dina(n21397), .dinb(n20910), .dout(n21398));
  jxor g21099(.dina(n21398), .dinb(n20782), .dout(n21399));
  jor  g21100(.dina(n21399), .dinb(n796), .dout(n21400));
  jor  g21101(.dina(n21391), .dinb(n1034), .dout(n21401));
  jand g21102(.dina(n21401), .dinb(n21400), .dout(n21402));
  jand g21103(.dina(n21402), .dinb(n21395), .dout(n21403));
  jnot g21104(.din(n20790), .dout(n21404));
  jnot g21105(.din(n20785), .dout(n21405));
  jand g21106(.dina(asqrt[1] ), .dinb(n21405), .dout(n21406));
  jnot g21107(.din(n21406), .dout(n21407));
  jor  g21108(.dina(n21407), .dinb(n21404), .dout(n21408));
  jand g21109(.dina(n21408), .dinb(n20788), .dout(n21409));
  jand g21110(.dina(n21406), .dinb(n20791), .dout(n21410));
  jor  g21111(.dina(n21410), .dinb(n21409), .dout(n21411));
  jand g21112(.dina(n21411), .dinb(n791), .dout(n21412));
  jand g21113(.dina(n21399), .dinb(n796), .dout(n21413));
  jor  g21114(.dina(n21413), .dinb(n21412), .dout(n21414));
  jor  g21115(.dina(n21414), .dinb(n21403), .dout(n21415));
  jnot g21116(.din(n20800), .dout(n21416));
  jnot g21117(.din(n20793), .dout(n21417));
  jand g21118(.dina(asqrt[1] ), .dinb(n21417), .dout(n21418));
  jnot g21119(.din(n21418), .dout(n21419));
  jor  g21120(.dina(n21419), .dinb(n21416), .dout(n21420));
  jand g21121(.dina(n21420), .dinb(n20797), .dout(n21421));
  jand g21122(.dina(n21418), .dinb(n20801), .dout(n21422));
  jor  g21123(.dina(n21422), .dinb(n21421), .dout(n21423));
  jor  g21124(.dina(n21423), .dinb(n595), .dout(n21424));
  jor  g21125(.dina(n21411), .dinb(n791), .dout(n21425));
  jand g21126(.dina(n21425), .dinb(n21424), .dout(n21426));
  jand g21127(.dina(n21426), .dinb(n21415), .dout(n21427));
  jxor g21128(.dina(n20802), .dinb(n595), .dout(n21428));
  jor  g21129(.dina(n21428), .dinb(n20910), .dout(n21429));
  jxor g21130(.dina(n21429), .dinb(n20813), .dout(n21430));
  jand g21131(.dina(n21430), .dinb(n590), .dout(n21431));
  jand g21132(.dina(n21423), .dinb(n595), .dout(n21432));
  jor  g21133(.dina(n21432), .dinb(n21431), .dout(n21433));
  jor  g21134(.dina(n21433), .dinb(n21427), .dout(n21434));
  jnot g21135(.din(n20818), .dout(n21435));
  jor  g21136(.dina(n21435), .dinb(n20816), .dout(n21436));
  jor  g21137(.dina(n21436), .dinb(n20910), .dout(n21437));
  jxor g21138(.dina(n21437), .dinb(n20827), .dout(n21438));
  jor  g21139(.dina(n21438), .dinb(n430), .dout(n21439));
  jor  g21140(.dina(n21430), .dinb(n590), .dout(n21440));
  jand g21141(.dina(n21440), .dinb(n21439), .dout(n21441));
  jand g21142(.dina(n21441), .dinb(n21434), .dout(n21442));
  jnot g21143(.din(n20835), .dout(n21443));
  jnot g21144(.din(n20830), .dout(n21444));
  jand g21145(.dina(asqrt[1] ), .dinb(n21444), .dout(n21445));
  jnot g21146(.din(n21445), .dout(n21446));
  jor  g21147(.dina(n21446), .dinb(n21443), .dout(n21447));
  jand g21148(.dina(n21447), .dinb(n20833), .dout(n21448));
  jand g21149(.dina(n21445), .dinb(n20836), .dout(n21449));
  jor  g21150(.dina(n21449), .dinb(n21448), .dout(n21450));
  jand g21151(.dina(n21450), .dinb(n425), .dout(n21451));
  jand g21152(.dina(n21438), .dinb(n430), .dout(n21452));
  jor  g21153(.dina(n21452), .dinb(n21451), .dout(n21453));
  jor  g21154(.dina(n21453), .dinb(n21442), .dout(n21454));
  jnot g21155(.din(n20845), .dout(n21455));
  jnot g21156(.din(n20838), .dout(n21456));
  jand g21157(.dina(asqrt[1] ), .dinb(n21456), .dout(n21457));
  jnot g21158(.din(n21457), .dout(n21458));
  jor  g21159(.dina(n21458), .dinb(n21455), .dout(n21459));
  jand g21160(.dina(n21459), .dinb(n20842), .dout(n21460));
  jand g21161(.dina(n21457), .dinb(n20846), .dout(n21461));
  jor  g21162(.dina(n21461), .dinb(n21460), .dout(n21462));
  jor  g21163(.dina(n21462), .dinb(n305), .dout(n21463));
  jor  g21164(.dina(n21450), .dinb(n425), .dout(n21464));
  jand g21165(.dina(n21464), .dinb(n21463), .dout(n21465));
  jand g21166(.dina(n21465), .dinb(n21454), .dout(n21466));
  jxor g21167(.dina(n20847), .dinb(n305), .dout(n21467));
  jor  g21168(.dina(n21467), .dinb(n20910), .dout(n21468));
  jxor g21169(.dina(n21468), .dinb(n20858), .dout(n21469));
  jand g21170(.dina(n21469), .dinb(n290), .dout(n21470));
  jand g21171(.dina(n21462), .dinb(n305), .dout(n21471));
  jor  g21172(.dina(n21471), .dinb(n21470), .dout(n21472));
  jor  g21173(.dina(n21472), .dinb(n21466), .dout(n21473));
  jnot g21174(.din(n20868), .dout(n21474));
  jnot g21175(.din(n20861), .dout(n21475));
  jand g21176(.dina(asqrt[1] ), .dinb(n21475), .dout(n21476));
  jnot g21177(.din(n21476), .dout(n21477));
  jor  g21178(.dina(n21477), .dinb(n21474), .dout(n21478));
  jand g21179(.dina(n21478), .dinb(n20865), .dout(n21479));
  jand g21180(.dina(n21476), .dinb(n20869), .dout(n21480));
  jor  g21181(.dina(n21480), .dinb(n21479), .dout(n21481));
  jor  g21182(.dina(n21481), .dinb(n223), .dout(n21482));
  jor  g21183(.dina(n21469), .dinb(n290), .dout(n21483));
  jand g21184(.dina(n21483), .dinb(n21482), .dout(n21484));
  jand g21185(.dina(n21484), .dinb(n21473), .dout(n21485));
  jand g21186(.dina(n20913), .dinb(n199), .dout(n21486));
  jand g21187(.dina(n21481), .dinb(n223), .dout(n21487));
  jor  g21188(.dina(n21487), .dinb(n21486), .dout(n21488));
  jor  g21189(.dina(n21488), .dinb(n21485), .dout(n21489));
  jand g21190(.dina(n21489), .dinb(n20914), .dout(n21490));
  jnot g21191(.din(n20877), .dout(n21491));
  jor  g21192(.dina(n21491), .dinb(n20875), .dout(n21492));
  jor  g21193(.dina(n21492), .dinb(n20910), .dout(n21493));
  jxor g21194(.dina(n21493), .dinb(n20886), .dout(n21494));
  jnot g21195(.din(n20902), .dout(n21495));
  jand g21196(.dina(asqrt[1] ), .dinb(n20901), .dout(n21496));
  jand g21197(.dina(n21496), .dinb(n20888), .dout(n21497));
  jor  g21198(.dina(n21497), .dinb(n21495), .dout(n21498));
  jor  g21199(.dina(n21498), .dinb(n21494), .dout(n21499));
  jor  g21200(.dina(n21499), .dinb(n21490), .dout(n21500));
  jand g21201(.dina(n21500), .dinb(n194), .dout(n21501));
  jand g21202(.dina(n21494), .dinb(n21490), .dout(n21502));
  jor  g21203(.dina(n21496), .dinb(n20888), .dout(n21503));
  jnot g21204(.din(n20888), .dout(n21504));
  jor  g21205(.dina(n20891), .dinb(n21504), .dout(n21505));
  jand g21206(.dina(n21505), .dinb(asqrt[63] ), .dout(n21506));
  jand g21207(.dina(n21506), .dinb(n21503), .dout(n21507));
  jor  g21208(.dina(n21507), .dinb(n21502), .dout(n21508));
  jor  g21209(.dina(n21508), .dinb(n21501), .dout(asqrt[0] ));
endmodule


