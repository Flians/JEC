module gf_c432(G115gat, G108gat, G102gat, G99gat, G112gat, G95gat, G92gat, G105gat, G37gat, G4gat, G69gat, G17gat, G34gat, G1gat, G79gat, G30gat, G14gat, G21gat, G53gat, G60gat, G8gat, G63gat, G11gat, G24gat, G40gat, G43gat, G82gat, G47gat, G50gat, G56gat, G66gat, G73gat, G89gat, G76gat, G27gat, G86gat, G432gat, G430gat, G421gat, G431gat, G370gat, G329gat, G223gat);
    input G115gat, G108gat, G102gat, G99gat, G112gat, G95gat, G92gat, G105gat, G37gat, G4gat, G69gat, G17gat, G34gat, G1gat, G79gat, G30gat, G14gat, G21gat, G53gat, G60gat, G8gat, G63gat, G11gat, G24gat, G40gat, G43gat, G82gat, G47gat, G50gat, G56gat, G66gat, G73gat, G89gat, G76gat, G27gat, G86gat;
    output G432gat, G430gat, G421gat, G431gat, G370gat, G329gat, G223gat;
    wire n45;
    wire n49;
    wire n52;
    wire n56;
    wire n59;
    wire n63;
    wire n66;
    wire n70;
    wire n73;
    wire n77;
    wire n81;
    wire n84;
    wire n88;
    wire n91;
    wire n95;
    wire n99;
    wire n103;
    wire n106;
    wire n110;
    wire n113;
    wire n117;
    wire n120;
    wire n124;
    wire n128;
    wire n132;
    wire n136;
    wire n140;
    wire n143;
    wire n146;
    wire n150;
    wire n153;
    wire n157;
    wire n160;
    wire n164;
    wire n168;
    wire n171;
    wire n175;
    wire n178;
    wire n182;
    wire n186;
    wire n190;
    wire n193;
    wire n197;
    wire n200;
    wire n204;
    wire n207;
    wire n211;
    wire n215;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n242;
    wire n246;
    wire n250;
    wire n254;
    wire n258;
    wire n261;
    wire n265;
    wire n269;
    wire n273;
    wire n276;
    wire n280;
    wire n284;
    wire n288;
    wire n292;
    wire n295;
    wire n299;
    wire n303;
    wire n307;
    wire n311;
    wire n315;
    wire n318;
    wire n322;
    wire n326;
    wire n330;
    wire n333;
    wire n337;
    wire n341;
    wire n345;
    wire n348;
    wire n352;
    wire n356;
    wire n360;
    wire n363;
    wire n367;
    wire n371;
    wire n375;
    wire n379;
    wire n383;
    wire n387;
    wire n391;
    wire n395;
    wire n399;
    wire n403;
    wire n407;
    wire n411;
    wire n414;
    wire n418;
    wire n421;
    wire n424;
    wire n428;
    wire n432;
    wire n436;
    wire n439;
    wire n443;
    wire n447;
    wire n451;
    wire n455;
    wire n459;
    wire n463;
    wire n467;
    wire n471;
    wire n475;
    wire n479;
    wire n483;
    wire n487;
    wire n490;
    wire n494;
    wire n498;
    wire n502;
    wire n506;
    wire n510;
    wire n513;
    wire n517;
    wire n521;
    wire n525;
    wire n529;
    wire n533;
    wire n537;
    wire n541;
    wire n545;
    wire n549;
    wire n553;
    wire n557;
    wire n561;
    wire n565;
    wire n569;
    wire n573;
    wire n577;
    wire n580;
    wire n584;
    wire n588;
    wire n592;
    wire n596;
    wire n599;
    wire n603;
    wire n607;
    wire n611;
    wire n614;
    wire n618;
    wire n622;
    wire n626;
    wire n630;
    wire n634;
    wire n637;
    wire n641;
    wire n645;
    wire n649;
    wire n652;
    wire n656;
    wire n660;
    wire n664;
    wire n668;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n687;
    wire n691;
    wire n695;
    wire n698;
    wire n702;
    wire n706;
    wire n710;
    wire n714;
    wire n717;
    wire n721;
    wire n725;
    wire n729;
    wire n733;
    wire n737;
    wire n741;
    wire n745;
    wire n749;
    wire n753;
    wire n757;
    wire n761;
    wire n765;
    wire n769;
    wire n773;
    wire n777;
    wire n781;
    wire n785;
    wire n789;
    wire n793;
    wire n797;
    wire n801;
    wire n805;
    wire n809;
    wire n813;
    wire n817;
    wire n821;
    wire n825;
    wire n829;
    wire n833;
    wire n837;
    wire n841;
    wire n845;
    wire n849;
    wire n853;
    wire n857;
    wire n861;
    wire n864;
    wire n868;
    wire n872;
    wire n876;
    wire n880;
    wire n884;
    wire n888;
    wire n891;
    wire n894;
    wire n897;
    wire n901;
    wire n905;
    wire n909;
    wire n913;
    wire n917;
    wire n921;
    wire n925;
    wire n929;
    wire n933;
    wire n937;
    wire n941;
    wire n945;
    wire n952;
    wire n956;
    wire n959;
    wire n963;
    wire n967;
    wire n971;
    wire n975;
    wire n979;
    wire n983;
    wire n987;
    wire n991;
    wire n995;
    wire n1003;
    wire n1007;
    wire n1011;
    wire n1015;
    wire n1466;
    wire n1469;
    wire n1472;
    wire n1475;
    wire n1478;
    wire n1481;
    wire n1484;
    wire n1487;
    wire n1490;
    wire n1493;
    wire n1495;
    wire n1499;
    wire n1501;
    wire n1505;
    wire n1508;
    wire n1511;
    wire n1514;
    wire n1517;
    wire n1520;
    wire n1523;
    wire n1526;
    wire n1529;
    wire n1532;
    wire n1535;
    wire n1538;
    wire n1541;
    wire n1544;
    wire n1547;
    wire n1550;
    wire n1553;
    wire n1556;
    wire n1559;
    wire n1562;
    wire n1565;
    wire n1568;
    wire n1571;
    wire n1574;
    wire n1577;
    wire n1579;
    wire n1582;
    wire n1585;
    wire n1589;
    wire n1591;
    wire n1594;
    wire n1597;
    wire n1600;
    wire n1603;
    wire n1606;
    wire n1610;
    wire n1613;
    wire n1616;
    wire n1619;
    wire n1622;
    wire n1625;
    wire n1628;
    wire n1631;
    wire n1634;
    wire n1637;
    wire n1640;
    wire n1642;
    wire n1645;
    wire n1648;
    wire n1651;
    wire n1654;
    wire n1658;
    wire n1661;
    wire n1663;
    wire n1666;
    wire n1669;
    wire n1672;
    wire n1675;
    wire n1678;
    wire n1681;
    wire n1684;
    wire n1687;
    wire n1690;
    wire n1693;
    wire n1697;
    wire n1700;
    wire n1703;
    wire n1706;
    wire n1709;
    wire n1712;
    wire n1715;
    wire n1718;
    wire n1721;
    wire n1724;
    wire n1727;
    wire n1730;
    wire n1733;
    wire n1736;
    wire n1738;
    wire n1741;
    wire n1744;
    wire n1747;
    wire n1750;
    wire n1753;
    wire n1756;
    wire n1759;
    wire n1762;
    wire n1765;
    wire n1768;
    wire n1772;
    wire n1775;
    wire n1778;
    wire n1781;
    wire n1784;
    wire n1787;
    wire n1790;
    wire n1793;
    wire n1796;
    wire n1799;
    wire n1802;
    wire n1805;
    wire n1808;
    wire n1811;
    wire n1814;
    wire n1817;
    wire n1820;
    wire n1823;
    wire n1826;
    wire n1829;
    wire n1832;
    wire n1835;
    wire n1838;
    wire n1841;
    wire n1844;
    wire n1847;
    wire n1850;
    wire n1853;
    wire n1856;
    wire n1859;
    wire n1862;
    wire n1865;
    wire n1868;
    wire n1871;
    wire n1874;
    wire n1877;
    wire n1880;
    wire n1883;
    wire n1886;
    wire n1889;
    wire n1892;
    wire n1895;
    wire n1897;
    wire n1900;
    wire n1903;
    wire n1906;
    wire n1909;
    wire n1913;
    wire n1916;
    wire n1919;
    wire n1922;
    wire n1925;
    wire n1928;
    wire n1931;
    wire n1934;
    wire n1937;
    wire n1940;
    wire n1943;
    wire n1946;
    wire n1949;
    wire n1952;
    wire n1955;
    wire n1957;
    wire n1960;
    wire n1963;
    wire n1966;
    wire n1969;
    wire n1973;
    wire n1976;
    wire n1979;
    wire n1982;
    wire n1985;
    wire n1988;
    wire n1991;
    wire n1994;
    wire n1997;
    wire n2000;
    wire n2003;
    wire n2006;
    wire n2009;
    wire n2012;
    wire n2014;
    wire n2017;
    wire n2020;
    wire n2023;
    wire n2026;
    wire n2029;
    wire n2032;
    wire n2035;
    wire n2038;
    wire n2042;
    wire n2045;
    wire n2047;
    wire n2050;
    wire n2053;
    wire n2056;
    wire n2059;
    wire n2062;
    wire n2065;
    wire n2068;
    wire n2071;
    wire n2074;
    wire n2077;
    wire n2080;
    wire n2083;
    wire n2086;
    wire n2089;
    wire n2092;
    wire n2095;
    wire n2098;
    wire n2101;
    wire n2104;
    wire n2107;
    wire n2110;
    wire n2113;
    wire n2116;
    wire n2119;
    wire n2122;
    wire n2125;
    wire n2128;
    wire n2131;
    wire n2134;
    wire n2137;
    wire n2140;
    wire n2143;
    wire n2146;
    wire n2149;
    wire n2152;
    wire n2155;
    wire n2158;
    wire n2161;
    wire n2164;
    wire n2167;
    wire n2170;
    wire n2173;
    wire n2176;
    wire n2179;
    wire n2182;
    wire n2185;
    wire n2188;
    wire n2191;
    wire n2194;
    wire n2197;
    wire n2200;
    wire n2203;
    wire n2206;
    wire n2209;
    wire n2212;
    wire n2215;
    wire n2218;
    wire n2221;
    wire n2224;
    wire n2227;
    wire n2230;
    wire n2233;
    wire n2236;
    wire n2239;
    wire n2242;
    wire n2245;
    wire n2248;
    wire n2251;
    wire n2254;
    wire n2257;
    wire n2260;
    wire n2263;
    wire n2266;
    wire n2269;
    wire n2272;
    wire n2275;
    wire n2278;
    wire n2281;
    wire n2284;
    wire n2287;
    wire n2290;
    wire n2293;
    wire n2296;
    wire n2299;
    wire n2302;
    wire n2305;
    wire n2308;
    wire n2311;
    wire n2314;
    wire n2317;
    wire n2320;
    wire n2323;
    wire n2326;
    wire n2329;
    wire n2332;
    wire n2335;
    wire n2338;
    wire n2341;
    wire n2344;
    wire n2347;
    wire n2350;
    wire n2353;
    wire n2356;
    wire n2359;
    wire n2362;
    wire n2365;
    wire n2368;
    wire n2371;
    wire n2374;
    wire n2377;
    wire n2380;
    wire n2384;
    wire n2387;
    wire n2390;
    wire n2393;
    wire n2396;
    wire n2398;
    wire n2401;
    wire n2404;
    wire n2407;
    wire n2410;
    wire n2413;
    wire n2416;
    wire n2419;
    wire n2422;
    wire n2425;
    wire n2428;
    wire n2431;
    wire n2434;
    wire n2437;
    wire n2440;
    wire n2443;
    wire n2446;
    wire n2449;
    wire n2452;
    wire n2455;
    wire n2458;
    wire n2461;
    wire n2464;
    wire n2467;
    wire n2470;
    wire n2473;
    wire n2476;
    wire n2479;
    wire n2482;
    wire n2485;
    wire n2488;
    wire n2491;
    wire n2494;
    wire n2497;
    wire n2500;
    wire n2503;
    wire n2506;
    wire n2509;
    wire n2512;
    wire n2515;
    wire n2518;
    wire n2521;
    wire n2524;
    wire n2527;
    wire n2530;
    wire n2533;
    wire n2536;
    wire n2539;
    wire n2542;
    wire n2545;
    wire n2548;
    wire n2552;
    wire n2555;
    wire n2558;
    wire n2561;
    wire n2564;
    wire n2567;
    wire n2569;
    wire n2572;
    wire n2575;
    wire n2578;
    wire n2581;
    wire n2584;
    wire n2587;
    wire n2590;
    wire n2593;
    wire n2596;
    wire n2599;
    wire n2602;
    wire n2606;
    wire n2609;
    wire n2612;
    wire n2615;
    wire n2618;
    wire n2621;
    wire n2624;
    wire n2626;
    wire n2629;
    wire n2632;
    wire n2635;
    wire n2638;
    wire n2641;
    wire n2644;
    wire n2647;
    wire n2650;
    wire n2653;
    wire n2656;
    wire n2659;
    wire n2662;
    wire n2665;
    wire n2668;
    wire n2671;
    wire n2674;
    wire n2677;
    wire n2680;
    wire n2683;
    wire n2686;
    wire n2690;
    wire n2693;
    wire n2696;
    wire n2699;
    wire n2702;
    wire n2705;
    wire n2708;
    wire n2711;
    wire n2713;
    wire n2716;
    wire n2719;
    wire n2722;
    wire n2725;
    wire n2728;
    wire n2731;
    wire n2734;
    wire n2737;
    wire n2740;
    wire n2743;
    wire n2746;
    wire n2749;
    wire n2752;
    wire n2755;
    wire n2758;
    wire n2761;
    wire n2764;
    wire n2768;
    wire n2771;
    wire n2774;
    wire n2777;
    wire n2780;
    wire n2783;
    wire n2786;
    wire n2788;
    wire n2791;
    wire n2794;
    wire n2797;
    wire n2800;
    wire n2803;
    wire n2806;
    wire n2809;
    wire n2812;
    wire n2815;
    wire n2818;
    wire n2822;
    wire n2825;
    wire n2828;
    wire n2831;
    wire n2834;
    wire n2837;
    wire n2840;
    wire n2843;
    wire n2846;
    wire n2848;
    wire n2851;
    wire n2854;
    wire n2857;
    wire n2860;
    wire n2863;
    wire n2866;
    wire n2869;
    wire n2872;
    wire n2875;
    wire n2878;
    wire n2882;
    wire n2885;
    wire n2888;
    wire n2891;
    wire n2894;
    wire n2897;
    wire n2900;
    wire n2902;
    wire n2905;
    wire n2908;
    wire n2911;
    wire n2914;
    wire n2917;
    wire n2920;
    wire n2923;
    wire n2926;
    wire n2929;
    wire n2932;
    wire n2936;
    wire n2939;
    wire n2942;
    wire n2945;
    wire n2948;
    wire n2951;
    wire n2954;
    wire n2957;
    wire n2960;
    wire n2963;
    wire n2966;
    wire n2969;
    wire n2972;
    wire n2975;
    wire n2977;
    wire n2980;
    wire n2983;
    wire n2986;
    wire n2989;
    wire n2992;
    wire n2995;
    wire n2998;
    wire n3001;
    wire n3004;
    wire n3007;
    wire n3011;
    wire n3014;
    wire n3017;
    wire n3020;
    wire n3023;
    wire n3026;
    wire n3029;
    wire n3031;
    wire n3034;
    wire n3037;
    wire n3040;
    wire n3043;
    wire n3046;
    wire n3049;
    wire n3052;
    wire n3055;
    wire n3058;
    wire n3061;
    wire n3064;
    wire n3067;
    wire n3070;
    wire n3073;
    wire n3076;
    wire n3079;
    wire n3082;
    wire n3085;
    wire n3088;
    wire n3092;
    wire n3095;
    wire n3098;
    wire n3101;
    wire n3104;
    wire n3107;
    wire n3110;
    wire n3113;
    wire n3116;
    wire n3119;
    wire n3122;
    wire n3125;
    wire n3128;
    wire n3131;
    wire n3133;
    wire n3136;
    wire n3139;
    wire n3142;
    wire n3145;
    wire n3148;
    wire n3151;
    wire n3154;
    wire n3157;
    wire n3160;
    wire n3163;
    wire n3166;
    wire n3169;
    wire n3172;
    wire n3175;
    wire n3178;
    wire n3181;
    wire n3184;
    wire n3187;
    wire n3190;
    wire n3193;
    wire n3197;
    wire n3200;
    wire n3202;
    wire n3205;
    wire n3208;
    wire n3211;
    wire n3214;
    wire n3217;
    wire n3220;
    wire n3223;
    wire n3226;
    wire n3229;
    wire n3232;
    wire n3235;
    wire n3238;
    wire n3241;
    wire n3244;
    wire n3247;
    wire n3250;
    wire n3253;
    wire n3256;
    wire n3259;
    wire n3262;
    wire n3265;
    wire n3268;
    wire n3271;
    wire n3274;
    wire n3277;
    wire n3280;
    wire n3283;
    wire n3286;
    wire n3289;
    wire n3292;
    wire n3295;
    wire n3298;
    wire n3301;
    wire n3304;
    wire n3307;
    wire n3310;
    wire n3313;
    wire n3316;
    wire n3319;
    wire n3322;
    wire n3325;
    wire n3328;
    wire n3331;
    wire n3334;
    wire n3337;
    wire n3340;
    wire n3343;
    wire n3346;
    wire n3349;
    wire n3352;
    wire n3355;
    wire n3358;
    wire n3361;
    wire n3364;
    wire n3367;
    wire n3370;
    wire n3373;
    wire n3376;
    wire n3379;
    wire n3382;
    wire n3385;
    wire n3388;
    wire n3391;
    wire n3394;
    wire n3397;
    wire n3400;
    wire n3403;
    wire n3406;
    wire n3409;
    wire n3412;
    wire n3415;
    wire n3418;
    wire n3421;
    wire n3424;
    wire n3427;
    wire n3430;
    wire n3433;
    wire n3436;
    wire n3439;
    wire n3442;
    wire n3445;
    wire n3448;
    wire n3451;
    wire n3454;
    wire n3457;
    wire n3460;
    wire n3463;
    wire n3467;
    wire n3470;
    wire n3473;
    wire n3476;
    wire n3479;
    wire n3482;
    wire n3485;
    wire n3487;
    wire n3490;
    wire n3493;
    wire n3496;
    wire n3499;
    wire n3502;
    wire n3505;
    wire n3508;
    wire n3511;
    wire n3514;
    wire n3517;
    wire n3520;
    wire n3523;
    wire n3527;
    wire n3530;
    wire n3532;
    wire n3535;
    wire n3538;
    wire n3541;
    wire n3544;
    wire n3547;
    wire n3551;
    wire n3554;
    wire n3557;
    wire n3560;
    wire n3563;
    wire n3566;
    wire n3568;
    wire n3571;
    wire n3574;
    wire n3577;
    wire n3580;
    wire n3583;
    wire n3586;
    wire n3589;
    wire n3592;
    wire n3595;
    wire n3598;
    wire n3601;
    wire n3604;
    wire n3607;
    wire n3610;
    wire n3613;
    wire n3616;
    wire n3619;
    wire n3622;
    wire n3625;
    wire n3628;
    wire n3631;
    wire n3634;
    wire n3637;
    wire n3640;
    wire n3643;
    wire n3646;
    wire n3649;
    wire n3652;
    wire n3655;
    wire n3658;
    wire n3661;
    wire n3664;
    wire n3667;
    wire n3670;
    wire n3673;
    wire n3676;
    wire n3679;
    wire n3682;
    wire n3685;
    wire n3688;
    wire n3691;
    wire n3694;
    wire n3697;
    wire n3700;
    wire n3703;
    wire n3706;
    wire n3709;
    wire n3712;
    wire n3715;
    wire n3718;
    wire n3721;
    wire n3724;
    wire n3727;
    wire n3730;
    wire n3733;
    wire n3736;
    wire n3739;
    wire n3742;
    wire n3745;
    wire n3748;
    wire n3751;
    wire n3754;
    wire n3757;
    wire n3760;
    wire n3763;
    wire n3766;
    wire n3769;
    wire n3772;
    wire n3775;
    wire n3778;
    wire n3781;
    wire n3784;
    wire n3787;
    wire n3790;
    wire n3793;
    wire n3796;
    wire n3799;
    wire n3802;
    wire n3805;
    wire n3808;
    wire n3811;
    wire n3814;
    wire n3817;
    wire n3820;
    wire n3823;
    wire n3826;
    wire n3830;
    wire n3833;
    wire n3835;
    wire n3838;
    wire n3841;
    wire n3844;
    wire n3847;
    wire n3850;
    wire n3853;
    wire n3856;
    wire n3859;
    wire n3862;
    wire n3865;
    wire n3868;
    wire n3871;
    wire n3874;
    wire n3877;
    wire n3880;
    wire n3883;
    wire n3886;
    wire n3889;
    wire n3892;
    wire n3895;
    wire n3898;
    wire n3901;
    wire n3904;
    wire n3907;
    wire n3910;
    wire n3913;
    wire n3916;
    wire n3919;
    wire n3922;
    wire n3925;
    wire n3928;
    wire n3931;
    wire n3934;
    wire n3937;
    wire n3940;
    wire n3943;
    wire n3946;
    wire n3949;
    wire n3952;
    wire n3955;
    wire n3958;
    wire n3961;
    wire n3964;
    wire n3967;
    wire n3970;
    wire n3973;
    wire n3976;
    wire n3979;
    wire n3982;
    wire n3985;
    wire n3988;
    wire n3991;
    wire n3994;
    wire n3997;
    wire n4000;
    wire n4003;
    wire n4006;
    wire n4010;
    wire n4013;
    wire n4016;
    wire n4019;
    wire n4022;
    wire n4025;
    wire n4028;
    wire n4030;
    wire n4033;
    wire n4036;
    wire n4039;
    wire n4042;
    wire n4045;
    wire n4048;
    wire n4051;
    wire n4054;
    wire n4057;
    wire n4060;
    wire n4063;
    wire n4066;
    wire n4069;
    wire n4072;
    wire n4075;
    wire n4078;
    wire n4081;
    wire n4084;
    wire n4087;
    wire n4090;
    wire n4093;
    wire n4096;
    wire n4099;
    wire n4102;
    wire n4105;
    wire n4108;
    wire n4112;
    wire n4115;
    wire n4117;
    wire n4120;
    wire n4123;
    wire n4126;
    wire n4129;
    wire n4132;
    wire n4135;
    wire n4138;
    wire n4141;
    wire n4144;
    wire n4147;
    wire n4150;
    wire n4153;
    wire n4156;
    wire n4159;
    wire n4162;
    wire n4165;
    wire n4168;
    wire n4171;
    wire n4174;
    wire n4177;
    wire n4180;
    wire n4183;
    wire n4186;
    wire n4189;
    wire n4192;
    wire n4195;
    wire n4198;
    wire n4201;
    wire n4204;
    wire n4207;
    wire n4210;
    wire n4213;
    wire n4216;
    wire n4219;
    wire n4222;
    wire n4225;
    wire n4228;
    wire n4231;
    wire n4234;
    wire n4237;
    wire n4240;
    wire n4243;
    wire n4246;
    wire n4249;
    wire n4252;
    wire n4255;
    wire n4258;
    wire n4261;
    wire n4264;
    wire n4267;
    wire n4270;
    wire n4273;
    wire n4276;
    wire n4279;
    wire n4282;
    wire n4285;
    wire n4288;
    wire n4291;
    wire n4294;
    wire n4297;
    wire n4300;
    wire n4303;
    wire n4306;
    wire n4309;
    wire n4312;
    wire n4315;
    wire n4318;
    wire n4321;
    wire n4324;
    wire n4327;
    wire n4330;
    wire n4333;
    wire n4336;
    wire n4339;
    wire n4342;
    wire n4345;
    wire n4348;
    wire n4351;
    wire n4354;
    wire n4357;
    wire n4360;
    wire n4363;
    wire n4366;
    wire n4369;
    wire n4372;
    wire n4375;
    wire n4378;
    wire n4381;
    wire n4384;
    wire n4387;
    wire n4390;
    wire n4393;
    wire n4396;
    wire n4399;
    wire n4402;
    wire n4405;
    wire n4408;
    wire n4411;
    wire n4414;
    wire n4417;
    wire n4420;
    wire n4423;
    wire n4426;
    wire n4429;
    wire n4432;
    wire n4435;
    wire n4438;
    wire n4441;
    wire n4444;
    wire n4447;
    wire n4450;
    wire n4453;
    wire n4456;
    wire n4459;
    wire n4462;
    wire n4465;
    wire n4468;
    wire n4471;
    wire n4474;
    wire n4477;
    wire n4480;
    wire n4483;
    wire n4486;
    wire n4489;
    wire n4492;
    wire n4495;
    wire n4498;
    wire n4501;
    wire n4504;
    wire n4507;
    wire n4510;
    wire n4513;
    wire n4516;
    wire n4519;
    wire n4522;
    wire n4525;
    wire n4528;
    wire n4531;
    wire n4534;
    wire n4537;
    wire n4540;
    wire n4543;
    wire n4546;
    wire n4549;
    wire n4552;
    wire n4555;
    wire n4558;
    wire n4561;
    wire n4564;
    wire n4567;
    wire n4570;
    wire n4573;
    wire n4576;
    wire n4579;
    wire n4582;
    wire n4585;
    wire n4588;
    wire n4591;
    wire n4594;
    wire n4597;
    wire n4600;
    wire n4603;
    wire n4606;
    wire n4609;
    wire n4612;
    wire n4615;
    wire n4618;
    wire n4621;
    wire n4624;
    wire n4627;
    wire n4630;
    wire n4633;
    wire n4636;
    wire n4639;
    wire n4642;
    wire n4645;
    wire n4648;
    wire n4651;
    wire n4654;
    wire n4658;
    wire n4660;
    wire n4663;
    wire n4666;
    wire n4669;
    wire n4672;
    wire n4675;
    wire n4678;
    wire n4681;
    wire n4684;
    wire n4687;
    wire n4690;
    wire n4693;
    wire n4696;
    wire n4699;
    wire n4702;
    wire n4705;
    wire n4708;
    wire n4711;
    wire n4714;
    wire n4717;
    wire n4720;
    wire n4723;
    wire n4726;
    wire n4729;
    wire n4732;
    wire n4735;
    wire n4738;
    wire n4741;
    wire n4744;
    wire n4747;
    wire n4750;
    wire n4753;
    wire n4756;
    wire n4759;
    wire n4762;
    wire n4765;
    wire n4768;
    wire n4771;
    wire n4774;
    wire n4777;
    wire n4780;
    wire n4783;
    wire n4786;
    wire n4789;
    wire n4792;
    wire n4795;
    wire n4798;
    wire n4801;
    wire n4804;
    wire n4807;
    wire n4810;
    wire n4813;
    wire n4816;
    wire n4819;
    wire n4822;
    wire n4825;
    wire n4828;
    wire n4831;
    wire n4834;
    wire n4837;
    wire n4840;
    wire n4843;
    wire n4846;
    wire n4849;
    wire n4852;
    wire n4858;
    wire n4861;
    wire n4864;
    wire n4867;
    wire n4870;
    wire n4873;
    wire n4876;
    wire n4879;
    wire n4882;
    wire n4885;
    wire n4888;
    wire n4891;
    wire n4894;
    wire n4900;
    wire n4903;
    wire n4906;
    wire n4909;
    wire n4912;
    wire n4915;
    wire n4921;
    jnot g000(.din(G102gat), .dout(n45));
    jand g001(.dinb(n45), .dina(n4723), .dout(n49));
    jnot g002(.din(G43gat), .dout(n52));
    jor g003(.dinb(n4658), .dina(n52), .dout(n56));
    jnot g004(.din(n56), .dout(n59));
    jor g005(.dinb(n4699), .dina(n59), .dout(n63));
    jnot g006(.din(G63gat), .dout(n66));
    jand g007(.dinb(n66), .dina(n4639), .dout(n70));
    jnot g008(.din(G11gat), .dout(n73));
    jand g009(.dinb(n73), .dina(n4576), .dout(n77));
    jor g010(.dinb(n70), .dina(n77), .dout(n81));
    jnot g011(.din(G24gat), .dout(n84));
    jand g012(.dinb(n84), .dina(n4513), .dout(n88));
    jnot g013(.din(G50gat), .dout(n91));
    jand g014(.dinb(n91), .dina(n4381), .dout(n95));
    jor g015(.dinb(n88), .dina(n95), .dout(n99));
    jor g016(.dinb(n81), .dina(n99), .dout(n103));
    jnot g017(.din(G1gat), .dout(n106));
    jand g018(.dinb(n106), .dina(n4282), .dout(n110));
    jnot g019(.din(G89gat), .dout(n113));
    jand g020(.dinb(n113), .dina(n4219), .dout(n117));
    jnot g021(.din(G76gat), .dout(n120));
    jand g022(.dinb(n120), .dina(n4156), .dout(n124));
    jor g023(.dinb(n117), .dina(n124), .dout(n128));
    jor g024(.dinb(n3833), .dina(n128), .dout(n132));
    jor g025(.dinb(n103), .dina(n132), .dout(n136));
    jor g026(.dinb(n3830), .dina(n136), .dout(n140));
    jnot g027(.din(G21gat), .dout(n143));
    jnot g028(.din(n49), .dout(n146));
    jand g029(.dinb(n146), .dina(n4654), .dout(n150));
    jnot g030(.din(G69gat), .dout(n153));
    jor g031(.dinb(n4792), .dina(n153), .dout(n157));
    jnot g032(.din(G17gat), .dout(n160));
    jor g033(.dinb(n4597), .dina(n160), .dout(n164));
    jand g034(.dinb(n157), .dina(n164), .dout(n168));
    jnot g035(.din(G30gat), .dout(n171));
    jor g036(.dinb(n4534), .dina(n171), .dout(n175));
    jnot g037(.din(G56gat), .dout(n178));
    jor g038(.dinb(n4471), .dina(n178), .dout(n182));
    jand g039(.dinb(n175), .dina(n182), .dout(n186));
    jand g040(.dinb(n168), .dina(n186), .dout(n190));
    jnot g041(.din(G4gat), .dout(n193));
    jor g042(.dinb(n4303), .dina(n193), .dout(n197));
    jnot g043(.din(G95gat), .dout(n200));
    jor g044(.dinb(n4240), .dina(n200), .dout(n204));
    jnot g045(.din(G82gat), .dout(n207));
    jor g046(.dinb(n4177), .dina(n207), .dout(n211));
    jand g047(.dinb(n204), .dina(n211), .dout(n215));
    jand g048(.dinb(n4115), .dina(n215), .dout(n219));
    jand g049(.dinb(n190), .dina(n219), .dout(n223));
    jand g050(.dinb(n4112), .dina(n223), .dout(n227));
    jor g051(.dinb(n3907), .dina(n227), .dout(n231));
    jand g052(.dinb(n4555), .dina(n231), .dout(n235));
    jand g053(.dinb(n3029), .dina(n235), .dout(n239));
    jnot g054(.din(G99gat), .dout(n242));
    jor g055(.dinb(n3850), .dina(n227), .dout(n246));
    jand g056(.dinb(n4198), .dina(n246), .dout(n250));
    jand g057(.dinb(n2975), .dina(n250), .dout(n254));
    jor g058(.dinb(n239), .dina(n254), .dout(n258));
    jnot g059(.din(G73gat), .dout(n261));
    jor g060(.dinb(n4759), .dina(n227), .dout(n265));
    jand g061(.dinb(n4618), .dina(n265), .dout(n269));
    jand g062(.dinb(n4028), .dina(n269), .dout(n273));
    jnot g063(.din(G34gat), .dout(n276));
    jor g064(.dinb(n3892), .dina(n227), .dout(n280));
    jand g065(.dinb(n4492), .dina(n280), .dout(n284));
    jand g066(.dinb(n2954), .dina(n284), .dout(n288));
    jor g067(.dinb(n273), .dina(n288), .dout(n292));
    jnot g068(.din(G112gat), .dout(n295));
    jor g069(.dinb(n4726), .dina(n227), .dout(n299));
    jand g070(.dinb(n4702), .dina(n299), .dout(n303));
    jand g071(.dinb(n2900), .dina(n303), .dout(n307));
    jor g072(.dinb(n292), .dina(n2846), .dout(n311));
    jor g073(.dinb(n2843), .dina(n311), .dout(n315));
    jnot g074(.din(G60gat), .dout(n318));
    jxor g075(.dinb(n3880), .dina(n227), .dout(n322));
    jand g076(.dinb(n4450), .dina(n322), .dout(n326));
    jand g077(.dinb(n3485), .dina(n326), .dout(n330));
    jnot g078(.din(G86gat), .dout(n333));
    jor g079(.dinb(n3835), .dina(n227), .dout(n337));
    jand g080(.dinb(n4135), .dina(n337), .dout(n341));
    jand g081(.dinb(n2840), .dina(n341), .dout(n345));
    jnot g082(.din(G8gat), .dout(n348));
    jor g083(.dinb(n3865), .dina(n227), .dout(n352));
    jand g084(.dinb(n4261), .dina(n352), .dout(n356));
    jand g085(.dinb(n2786), .dina(n356), .dout(n360));
    jnot g086(.din(G47gat), .dout(n363));
    jor g087(.dinb(n3922), .dina(n227), .dout(n367));
    jand g088(.dinb(n4678), .dina(n367), .dout(n371));
    jand g089(.dinb(n2711), .dina(n371), .dout(n375));
    jor g090(.dinb(n360), .dina(n375), .dout(n379));
    jor g091(.dinb(n2690), .dina(n379), .dout(n383));
    jor g092(.dinb(n3427), .dina(n383), .dout(n387));
    jor g093(.dinb(n315), .dina(n387), .dout(n391));
    jand g094(.dinb(n4222), .dina(n140), .dout(n395));
    jor g095(.dinb(n4180), .dina(n395), .dout(n399));
    jand g096(.dinb(n3772), .dina(n391), .dout(n403));
    jor g097(.dinb(n3730), .dina(n403), .dout(n407));
    jor g098(.dinb(n3031), .dina(n407), .dout(n411));
    jnot g099(.din(n411), .dout(n414));
    jand g100(.dinb(n3226), .dina(n391), .dout(n418));
    jnot g101(.din(n418), .dout(n421));
    jnot g102(.din(G53gat), .dout(n424));
    jand g103(.dinb(n2624), .dina(n371), .dout(n428));
    jand g104(.dinb(n421), .dina(n2567), .dout(n432));
    jor g105(.dinb(n414), .dina(n2548), .dout(n436));
    jnot g106(.din(G40gat), .dout(n439));
    jand g107(.dinb(n4579), .dina(n140), .dout(n443));
    jor g108(.dinb(n4537), .dina(n443), .dout(n447));
    jor g109(.dinb(n3970), .dina(n447), .dout(n451));
    jor g110(.dinb(n3748), .dina(n399), .dout(n455));
    jand g111(.dinb(n451), .dina(n455), .dout(n459));
    jand g112(.dinb(n4774), .dina(n140), .dout(n463));
    jor g113(.dinb(n4600), .dina(n463), .dout(n467));
    jor g114(.dinb(n4069), .dina(n467), .dout(n471));
    jand g115(.dinb(n4516), .dina(n140), .dout(n475));
    jor g116(.dinb(n4474), .dina(n475), .dout(n479));
    jor g117(.dinb(n3688), .dina(n479), .dout(n483));
    jand g118(.dinb(n471), .dina(n483), .dout(n487));
    jnot g119(.din(G108gat), .dout(n490));
    jand g120(.dinb(n4741), .dina(n140), .dout(n494));
    jor g121(.dinb(n3566), .dina(n494), .dout(n498));
    jor g122(.dinb(n3607), .dina(n498), .dout(n502));
    jand g123(.dinb(n487), .dina(n3530), .dout(n506));
    jand g124(.dinb(n3527), .dina(n506), .dout(n510));
    jnot g125(.din(n330), .dout(n513));
    jand g126(.dinb(n4159), .dina(n140), .dout(n517));
    jor g127(.dinb(n4117), .dina(n517), .dout(n521));
    jor g128(.dinb(n3403), .dina(n521), .dout(n525));
    jand g129(.dinb(n4285), .dina(n140), .dout(n529));
    jor g130(.dinb(n4243), .dina(n529), .dout(n533));
    jor g131(.dinb(n3322), .dina(n533), .dout(n537));
    jand g132(.dinb(n4642), .dina(n140), .dout(n541));
    jor g133(.dinb(n4660), .dina(n541), .dout(n545));
    jor g134(.dinb(n3202), .dina(n545), .dout(n549));
    jand g135(.dinb(n537), .dina(n549), .dout(n553));
    jand g136(.dinb(n3200), .dina(n553), .dout(n557));
    jand g137(.dinb(n3197), .dina(n557), .dout(n561));
    jand g138(.dinb(n510), .dina(n561), .dout(n565));
    jor g139(.dinb(n2920), .dina(n565), .dout(n569));
    jand g140(.dinb(n2902), .dina(n569), .dout(n573));
    jand g141(.dinb(n2012), .dina(n573), .dout(n577));
    jnot g142(.din(G66gat), .dout(n580));
    jor g143(.dinb(n3451), .dina(n565), .dout(n584));
    jand g144(.dinb(n3433), .dina(n584), .dout(n588));
    jand g145(.dinb(n1952), .dina(n588), .dout(n592));
    jor g146(.dinb(n577), .dina(n592), .dout(n596));
    jnot g147(.din(G14gat), .dout(n599));
    jor g148(.dinb(n2752), .dina(n565), .dout(n603));
    jand g149(.dinb(n2734), .dina(n603), .dout(n607));
    jand g150(.dinb(n1895), .dina(n607), .dout(n611));
    jnot g151(.din(G92gat), .dout(n614));
    jor g152(.dinb(n2806), .dina(n565), .dout(n618));
    jand g153(.dinb(n2788), .dina(n618), .dout(n622));
    jand g154(.dinb(n1853), .dina(n622), .dout(n626));
    jor g155(.dinb(n611), .dina(n626), .dout(n630));
    jor g156(.dinb(n596), .dina(n630), .dout(n634));
    jnot g157(.din(G79gat), .dout(n637));
    jor g158(.dinb(n3994), .dina(n565), .dout(n641));
    jand g159(.dinb(n4093), .dina(n641), .dout(n645));
    jand g160(.dinb(n3131), .dina(n645), .dout(n649));
    jnot g161(.din(G115gat), .dout(n652));
    jor g162(.dinb(n2866), .dina(n565), .dout(n656));
    jand g163(.dinb(n2848), .dina(n656), .dout(n660));
    jand g164(.dinb(n1811), .dina(n660), .dout(n664));
    jor g165(.dinb(n649), .dina(n664), .dout(n668));
    jnot g166(.din(G27gat), .dout(n671));
    jor g167(.dinb(n2995), .dina(n565), .dout(n675));
    jand g168(.dinb(n2977), .dina(n675), .dout(n679));
    jand g169(.dinb(n1736), .dina(n679), .dout(n683));
    jor g170(.dinb(n668), .dina(n1661), .dout(n687));
    jor g171(.dinb(n634), .dina(n687), .dout(n691));
    jor g172(.dinb(n1658), .dina(n691), .dout(n695));
    jnot g173(.din(n432), .dout(n698));
    jand g174(.dinb(n2686), .dina(n698), .dout(n702));
    jand g175(.dinb(n3649), .dina(n391), .dout(n706));
    jor g176(.dinb(n3631), .dina(n706), .dout(n710));
    jor g177(.dinb(n2503), .dina(n710), .dout(n714));
    jnot g178(.din(n326), .dout(n717));
    jand g179(.dinb(n3487), .dina(n391), .dout(n721));
    jor g180(.dinb(n2396), .dina(n721), .dout(n725));
    jor g181(.dinb(n2458), .dina(n725), .dout(n729));
    jand g182(.dinb(n714), .dina(n729), .dout(n733));
    jand g183(.dinb(n3283), .dina(n391), .dout(n737));
    jor g184(.dinb(n3265), .dina(n737), .dout(n741));
    jor g185(.dinb(n2338), .dina(n741), .dout(n745));
    jand g186(.dinb(n3364), .dina(n391), .dout(n749));
    jor g187(.dinb(n3346), .dina(n749), .dout(n753));
    jor g188(.dinb(n2215), .dina(n753), .dout(n757));
    jand g189(.dinb(n745), .dina(n757), .dout(n761));
    jand g190(.dinb(n733), .dina(n761), .dout(n765));
    jand g191(.dinb(n4030), .dina(n391), .dout(n769));
    jor g192(.dinb(n3712), .dina(n769), .dout(n773));
    jor g193(.dinb(n3133), .dina(n773), .dout(n777));
    jand g194(.dinb(n3568), .dina(n391), .dout(n781));
    jor g195(.dinb(n3532), .dina(n781), .dout(n785));
    jor g196(.dinb(n2092), .dina(n785), .dout(n789));
    jand g197(.dinb(n777), .dina(n789), .dout(n793));
    jand g198(.dinb(n3931), .dina(n391), .dout(n797));
    jor g199(.dinb(n3811), .dina(n797), .dout(n801));
    jor g200(.dinb(n2047), .dina(n801), .dout(n805));
    jand g201(.dinb(n793), .dina(n2045), .dout(n809));
    jand g202(.dinb(n765), .dina(n809), .dout(n813));
    jand g203(.dinb(n2042), .dina(n813), .dout(n817));
    jor g204(.dinb(n1681), .dina(n817), .dout(n821));
    jand g205(.dinb(n1663), .dina(n821), .dout(n825));
    jor g206(.dinb(n1957), .dina(n817), .dout(n829));
    jand g207(.dinb(n2014), .dina(n829), .dout(n833));
    jor g208(.dinb(n825), .dina(n833), .dout(n837));
    jor g209(.dinb(n2569), .dina(n817), .dout(n841));
    jand g210(.dinb(n2713), .dina(n421), .dout(n845));
    jand g211(.dinb(n841), .dina(n1642), .dout(n849));
    jor g212(.dinb(n1897), .dina(n817), .dout(n853));
    jand g213(.dinb(n4306), .dina(n140), .dout(n857));
    jor g214(.dinb(n1628), .dina(n721), .dout(n861));
    jnot g215(.din(n861), .dout(n864));
    jand g216(.dinb(n853), .dina(n1490), .dout(n868));
    jand g217(.dinb(n4384), .dina(n868), .dout(n872));
    jor g218(.dinb(n1577), .dina(n872), .dout(n876));
    jor g219(.dinb(n1499), .dina(n876), .dout(n880));
    jand g220(.dinb(n2155), .dina(n695), .dout(n884));
    jor g221(.dinb(n2137), .dina(n884), .dout(n888));
    jnot g222(.din(n888), .dout(n891));
    jnot g223(.din(n407), .dout(n894));
    jnot g224(.din(G105gat), .dout(n897));
    jor g225(.dinb(n1574), .dina(n817), .dout(n901));
    jand g226(.dinb(n1517), .dina(n901), .dout(n905));
    jor g227(.dinb(n3076), .dina(n817), .dout(n909));
    jand g228(.dinb(n3178), .dina(n909), .dout(n913));
    jor g229(.dinb(n1756), .dina(n817), .dout(n917));
    jand g230(.dinb(n1738), .dina(n917), .dout(n921));
    jor g231(.dinb(n913), .dina(n921), .dout(n925));
    jor g232(.dinb(n1501), .dina(n925), .dout(n929));
    jor g233(.dinb(n1493), .dina(n929), .dout(n933));
    jor g234(.dinb(n880), .dina(n933), .dout(n937));
    jand g235(.dinb(n2278), .dina(n695), .dout(n941));
    jor g236(.dinb(n2260), .dina(n941), .dout(n945));
    jand g237(.dinb(n937), .dina(n1475), .dout(G421gat));
    jnot g238(.din(n833), .dout(n952));
    jand g239(.dinb(n2626), .dina(n695), .dout(n956));
    jnot g240(.din(n845), .dout(n959));
    jor g241(.dinb(n956), .dina(n1640), .dout(n963));
    jand g242(.dinb(n2398), .dina(n695), .dout(n967));
    jor g243(.dinb(n967), .dina(n1591), .dout(n971));
    jor g244(.dinb(n4318), .dina(n971), .dout(n975));
    jand g245(.dinb(n1589), .dina(n975), .dout(n979));
    jand g246(.dinb(n1955), .dina(n979), .dout(n983));
    jand g247(.dinb(n2032), .dina(n983), .dout(n987));
    jand g248(.dinb(n979), .dina(n1493), .dout(n991));
    jor g249(.dinb(n1495), .dina(n991), .dout(n995));
    jor g250(.dinb(n987), .dina(n995), .dout(G431gat));
    jand g251(.dinb(n888), .dina(n905), .dout(n1003));
    jor g252(.dinb(n1577), .dina(n1003), .dout(n1007));
    jand g253(.dinb(n1955), .dina(n1007), .dout(n1011));
    jor g254(.dinb(n1579), .dina(n1011), .dout(n1015));
    jor g255(.dinb(n987), .dina(n1015), .dout(G432gat));
    jdff dff_A_2cvsLWe78_0(.din(n4921), .dout(G430gat));
    jdff dff_A_azFe6ujw4_1(.din(n880), .dout(n4921));
    jdff dff_A_z3jNHQMA0_0(.din(n4915), .dout(G370gat));
    jdff dff_A_iswhRiWp5_0(.din(n4912), .dout(n4915));
    jdff dff_A_KTsi93jF9_0(.din(n4909), .dout(n4912));
    jdff dff_A_u0dyAunK0_0(.din(n4906), .dout(n4909));
    jdff dff_A_aDqauZ9T3_0(.din(n4903), .dout(n4906));
    jdff dff_A_a9rIOCa60_0(.din(n4900), .dout(n4903));
    jdff dff_A_yBeS5tNQ7_2(.din(n695), .dout(n4900));
    jdff dff_A_p8mRBsUd9_0(.din(n4894), .dout(G329gat));
    jdff dff_A_UuQOzaaV8_0(.din(n4891), .dout(n4894));
    jdff dff_A_9FNc9TVV7_0(.din(n4888), .dout(n4891));
    jdff dff_A_qXojXBgN6_0(.din(n4885), .dout(n4888));
    jdff dff_A_43gH8nQM2_0(.din(n4882), .dout(n4885));
    jdff dff_A_lrl24h1E3_0(.din(n4879), .dout(n4882));
    jdff dff_A_yhzrV6pF0_0(.din(n4876), .dout(n4879));
    jdff dff_A_NrCqfr6e4_0(.din(n4873), .dout(n4876));
    jdff dff_A_CSDyzqPJ5_0(.din(n4870), .dout(n4873));
    jdff dff_A_p08ej82O1_0(.din(n4867), .dout(n4870));
    jdff dff_A_046ZAo3f0_0(.din(n4864), .dout(n4867));
    jdff dff_A_QGRhmXyi2_0(.din(n4861), .dout(n4864));
    jdff dff_A_g5CDUu0d0_0(.din(n4858), .dout(n4861));
    jdff dff_A_n8EDLT5F7_1(.din(n391), .dout(n4858));
    jdff dff_A_7QgaQTST6_0(.din(n4852), .dout(G223gat));
    jdff dff_A_8gq10dYw0_0(.din(n4849), .dout(n4852));
    jdff dff_A_N81KYzpx5_0(.din(n4846), .dout(n4849));
    jdff dff_A_fU2MW94j0_0(.din(n4843), .dout(n4846));
    jdff dff_A_bl0NvcbN2_0(.din(n4840), .dout(n4843));
    jdff dff_A_5ANkbwFV0_0(.din(n4837), .dout(n4840));
    jdff dff_A_F6lggsDY0_0(.din(n4834), .dout(n4837));
    jdff dff_A_HrY8qfug8_0(.din(n4831), .dout(n4834));
    jdff dff_A_KSXBSmRr2_0(.din(n4828), .dout(n4831));
    jdff dff_A_mIpwl0R25_0(.din(n4825), .dout(n4828));
    jdff dff_A_uHCETZMJ0_0(.din(n4822), .dout(n4825));
    jdff dff_A_jEd241Z64_0(.din(n4819), .dout(n4822));
    jdff dff_A_cxMmrtHl2_0(.din(n4816), .dout(n4819));
    jdff dff_A_fo5d3vHc4_0(.din(n4813), .dout(n4816));
    jdff dff_A_iBZzaS8T9_0(.din(n4810), .dout(n4813));
    jdff dff_A_nxGMixCD4_0(.din(n4807), .dout(n4810));
    jdff dff_A_yAs7j40J5_0(.din(n4804), .dout(n4807));
    jdff dff_A_6RXb5wTr2_0(.din(n4801), .dout(n4804));
    jdff dff_A_W85J9Emz9_0(.din(n4798), .dout(n4801));
    jdff dff_A_FgI7NOuD4_0(.din(n4795), .dout(n4798));
    jdff dff_A_SEMGl6Zg8_1(.din(n140), .dout(n4795));
    jdff dff_A_zdoTkP3m3_1(.din(G63gat), .dout(n4792));
    jdff dff_A_usOypx327_0(.din(G63gat), .dout(n4789));
    jdff dff_A_ObiHwby38_0(.din(n4789), .dout(n4786));
    jdff dff_A_7z1ywyqd3_0(.din(n4786), .dout(n4783));
    jdff dff_A_bgSF60ae4_0(.din(n4783), .dout(n4780));
    jdff dff_A_ojfR0qZ85_0(.din(n4780), .dout(n4777));
    jdff dff_A_81gjaSbA7_0(.din(n4777), .dout(n4774));
    jdff dff_A_zUzEfCVk4_0(.din(n66), .dout(n4771));
    jdff dff_A_9vXIbKq39_0(.din(n4771), .dout(n4768));
    jdff dff_A_mWIZI3vw2_0(.din(n4768), .dout(n4765));
    jdff dff_A_cnpsrrmk0_0(.din(n4765), .dout(n4762));
    jdff dff_A_WfdLipTW7_0(.din(n4762), .dout(n4759));
    jdff dff_A_70y3XZk07_0(.din(G102gat), .dout(n4756));
    jdff dff_A_JaxLAtvC3_0(.din(n4756), .dout(n4753));
    jdff dff_A_pz45IahK8_0(.din(n4753), .dout(n4750));
    jdff dff_A_o6ixDT2s2_0(.din(n4750), .dout(n4747));
    jdff dff_A_45DDNgtQ3_0(.din(n4747), .dout(n4744));
    jdff dff_A_N65usaMv8_0(.din(n4744), .dout(n4741));
    jdff dff_A_YwwioSY85_0(.din(n45), .dout(n4738));
    jdff dff_A_TNcbctzq1_0(.din(n4738), .dout(n4735));
    jdff dff_A_UfIjYvQB1_0(.din(n4735), .dout(n4732));
    jdff dff_A_2znjptDJ4_0(.din(n4732), .dout(n4729));
    jdff dff_A_xAe2rTE61_0(.din(n4729), .dout(n4726));
    jdff dff_A_4i46PGmI0_2(.din(G108gat), .dout(n4723));
    jdff dff_A_W3svUPV46_1(.din(G108gat), .dout(n4720));
    jdff dff_A_IAtl95gj8_1(.din(n4720), .dout(n4717));
    jdff dff_A_SH013tnM8_1(.din(n4717), .dout(n4714));
    jdff dff_A_gvY4XCXn2_1(.din(n4714), .dout(n4711));
    jdff dff_A_MbjdOFz08_1(.din(n4711), .dout(n4708));
    jdff dff_A_iWOI8SEZ1_1(.din(n4708), .dout(n4705));
    jdff dff_A_NucbvHI39_1(.din(n4705), .dout(n4702));
    jdff dff_A_ebpXr9Hh7_1(.din(n49), .dout(n4699));
    jdff dff_A_MieW2VVm4_0(.din(G43gat), .dout(n4696));
    jdff dff_A_wbdwtidA6_0(.din(n4696), .dout(n4693));
    jdff dff_A_qgQcvee10_0(.din(n4693), .dout(n4690));
    jdff dff_A_PXIAEZS05_0(.din(n4690), .dout(n4687));
    jdff dff_A_gyc3Z5Gb4_0(.din(n4687), .dout(n4684));
    jdff dff_A_GRRshK6s2_0(.din(n4684), .dout(n4681));
    jdff dff_A_XNVAdMtj9_0(.din(n4681), .dout(n4678));
    jdff dff_A_q6JCB2dB3_0(.din(n52), .dout(n4675));
    jdff dff_A_sOhfZZak9_0(.din(n4675), .dout(n4672));
    jdff dff_A_Q0N3R1ey1_0(.din(n4672), .dout(n4669));
    jdff dff_A_FDkYign09_0(.din(n4669), .dout(n4666));
    jdff dff_A_OQjvPBdC0_0(.din(n4666), .dout(n4663));
    jdff dff_A_Gv5iyWLq3_0(.din(n4663), .dout(n4660));
    jdff dff_B_Ml2pD0BU8_1(.din(G37gat), .dout(n4658));
    jdff dff_A_ywAkzHm66_1(.din(n56), .dout(n4654));
    jdff dff_A_B7Epgujb4_0(.din(n56), .dout(n4651));
    jdff dff_A_ZQ72B3iZ6_0(.din(n4651), .dout(n4648));
    jdff dff_A_vP4Y4k477_0(.din(n4648), .dout(n4645));
    jdff dff_A_EMEt9F877_0(.din(n4645), .dout(n4642));
    jdff dff_A_CDaLzzUH4_2(.din(G69gat), .dout(n4639));
    jdff dff_A_7wRvwOcp8_0(.din(G69gat), .dout(n4636));
    jdff dff_A_UnP2Bxod0_0(.din(n4636), .dout(n4633));
    jdff dff_A_Jtk8u1bt3_0(.din(n4633), .dout(n4630));
    jdff dff_A_hKHameyp3_0(.din(n4630), .dout(n4627));
    jdff dff_A_A8Ooo5bE8_0(.din(n4627), .dout(n4624));
    jdff dff_A_kAOLIRaY0_0(.din(n4624), .dout(n4621));
    jdff dff_A_pOArUeeG7_0(.din(n4621), .dout(n4618));
    jdff dff_A_DfSg4lqe1_0(.din(n153), .dout(n4615));
    jdff dff_A_BvclH8Jb5_0(.din(n4615), .dout(n4612));
    jdff dff_A_tH7PkBp22_0(.din(n4612), .dout(n4609));
    jdff dff_A_cSSoVR0x0_0(.din(n4609), .dout(n4606));
    jdff dff_A_5Q2BFT2c6_0(.din(n4606), .dout(n4603));
    jdff dff_A_iICP0BMf4_0(.din(n4603), .dout(n4600));
    jdff dff_A_asY2EJUK6_1(.din(G11gat), .dout(n4597));
    jdff dff_A_X0lqFf1U5_0(.din(G11gat), .dout(n4594));
    jdff dff_A_e7Fk9voQ8_0(.din(n4594), .dout(n4591));
    jdff dff_A_gyI1bUZ51_0(.din(n4591), .dout(n4588));
    jdff dff_A_2N3DnU7i7_0(.din(n4588), .dout(n4585));
    jdff dff_A_DC01FJdH6_0(.din(n4585), .dout(n4582));
    jdff dff_A_oZF4Mh1o2_0(.din(n4582), .dout(n4579));
    jdff dff_A_2GQp74W96_2(.din(G17gat), .dout(n4576));
    jdff dff_A_KATBrZG45_0(.din(G17gat), .dout(n4573));
    jdff dff_A_i1HZzGEE2_0(.din(n4573), .dout(n4570));
    jdff dff_A_VUb1qwie9_0(.din(n4570), .dout(n4567));
    jdff dff_A_VqdGLU0k9_0(.din(n4567), .dout(n4564));
    jdff dff_A_Y53OLZNa4_0(.din(n4564), .dout(n4561));
    jdff dff_A_5hpQmw7i6_0(.din(n4561), .dout(n4558));
    jdff dff_A_1r8vJFC17_0(.din(n4558), .dout(n4555));
    jdff dff_A_jCXMQBrh3_0(.din(n160), .dout(n4552));
    jdff dff_A_HE4889sh5_0(.din(n4552), .dout(n4549));
    jdff dff_A_tN7AdNdI6_0(.din(n4549), .dout(n4546));
    jdff dff_A_52ov8LUL3_0(.din(n4546), .dout(n4543));
    jdff dff_A_CCVTszga5_0(.din(n4543), .dout(n4540));
    jdff dff_A_LaLU8o9Q5_0(.din(n4540), .dout(n4537));
    jdff dff_A_AuOKD7660_1(.din(G24gat), .dout(n4534));
    jdff dff_A_w7lt1dcp9_0(.din(G24gat), .dout(n4531));
    jdff dff_B_vwebLdyM5_0(.din(n945), .dout(n1466));
    jdff dff_B_oLBFTUv28_0(.din(n1466), .dout(n1469));
    jdff dff_B_SoG1fvF07_0(.din(n1469), .dout(n1472));
    jdff dff_B_79cmHCEP3_0(.din(n1472), .dout(n1475));
    jdff dff_B_wCIJXmYt4_0(.din(n864), .dout(n1478));
    jdff dff_B_qxQuhH704_0(.din(n1478), .dout(n1481));
    jdff dff_B_gUf4KBF24_0(.din(n1481), .dout(n1484));
    jdff dff_B_3oNaz6UP6_0(.din(n1484), .dout(n1487));
    jdff dff_B_8uzFWmwk8_0(.din(n1487), .dout(n1490));
    jdff dff_B_r4O0bDM98_2(.din(n891), .dout(n1493));
    jdff dff_A_ePfqqCRY9_0(.din(n1499), .dout(n1495));
    jdff dff_B_RfiQmJcF3_2(.din(n837), .dout(n1499));
    jdff dff_A_V53s9Bud7_1(.din(n905), .dout(n1501));
    jdff dff_B_43yBtcuU3_1(.din(n894), .dout(n1505));
    jdff dff_B_KVHQTPUU2_1(.din(n1505), .dout(n1508));
    jdff dff_B_tOvj13OK4_1(.din(n1508), .dout(n1511));
    jdff dff_B_qrDAUZOZ2_1(.din(n1511), .dout(n1514));
    jdff dff_B_FgqCtSzS2_1(.din(n1514), .dout(n1517));
    jdff dff_B_KOSLGNRT6_1(.din(n897), .dout(n1520));
    jdff dff_B_LmmiM9Xv9_1(.din(n1520), .dout(n1523));
    jdff dff_B_LfGHjFt56_1(.din(n1523), .dout(n1526));
    jdff dff_B_CPy1CaQU2_1(.din(n1526), .dout(n1529));
    jdff dff_B_25uQAo1M0_1(.din(n1529), .dout(n1532));
    jdff dff_B_hSBrOcX19_1(.din(n1532), .dout(n1535));
    jdff dff_B_E0fz8Fo44_1(.din(n1535), .dout(n1538));
    jdff dff_B_cMRFAcil9_1(.din(n1538), .dout(n1541));
    jdff dff_B_WnVUmdgl8_1(.din(n1541), .dout(n1544));
    jdff dff_B_wwQQdLiQ3_1(.din(n1544), .dout(n1547));
    jdff dff_B_yN1SrVII7_1(.din(n1547), .dout(n1550));
    jdff dff_B_O01IHSQm2_1(.din(n1550), .dout(n1553));
    jdff dff_B_szApWXCv5_1(.din(n1553), .dout(n1556));
    jdff dff_B_pOZNkinj4_1(.din(n1556), .dout(n1559));
    jdff dff_B_zQrb1Bal0_1(.din(n1559), .dout(n1562));
    jdff dff_B_ODz5wPXy6_1(.din(n1562), .dout(n1565));
    jdff dff_B_4KOH86ug3_1(.din(n1565), .dout(n1568));
    jdff dff_B_CN6R47Uy5_1(.din(n1568), .dout(n1571));
    jdff dff_B_HKO3SEqS9_1(.din(n1571), .dout(n1574));
    jdff dff_B_uui4NYYm0_2(.din(n849), .dout(n1577));
    jdff dff_A_XDeI3lnr5_0(.din(n1582), .dout(n1579));
    jdff dff_A_e9DjkIqI4_0(.din(n1585), .dout(n1582));
    jdff dff_A_svtpdesh5_0(.din(n825), .dout(n1585));
    jdff dff_B_eJEne66E0_1(.din(n963), .dout(n1589));
    jdff dff_A_GZGs2fVn7_0(.din(n1594), .dout(n1591));
    jdff dff_A_6UT3alEb7_0(.din(n1597), .dout(n1594));
    jdff dff_A_ssRhug4y7_0(.din(n1600), .dout(n1597));
    jdff dff_A_2GaXWSBg2_0(.din(n1603), .dout(n1600));
    jdff dff_A_cVOe3GPp0_0(.din(n1606), .dout(n1603));
    jdff dff_A_cQsYk8by8_0(.din(n861), .dout(n1606));
    jdff dff_B_d4byrfUW0_1(.din(n857), .dout(n1610));
    jdff dff_B_38Cgd16t7_1(.din(n1610), .dout(n1613));
    jdff dff_B_JDh6NcOG2_1(.din(n1613), .dout(n1616));
    jdff dff_B_PCjPAHOB3_1(.din(n1616), .dout(n1619));
    jdff dff_B_PLk0RNOm6_1(.din(n1619), .dout(n1622));
    jdff dff_B_6Urc5rC95_1(.din(n1622), .dout(n1625));
    jdff dff_B_3iyEOD4r6_1(.din(n1625), .dout(n1628));
    jdff dff_B_E92dO7Rk5_0(.din(n959), .dout(n1631));
    jdff dff_B_iO0msDPq8_0(.din(n1631), .dout(n1634));
    jdff dff_B_vuu4jUCe9_0(.din(n1634), .dout(n1637));
    jdff dff_B_iwDUkmAt4_0(.din(n1637), .dout(n1640));
    jdff dff_A_bwA1ag0Z4_1(.din(n1645), .dout(n1642));
    jdff dff_A_KlHbBqMD0_1(.din(n1648), .dout(n1645));
    jdff dff_A_OITiqYk01_1(.din(n1651), .dout(n1648));
    jdff dff_A_75VzJehO6_1(.din(n1654), .dout(n1651));
    jdff dff_A_e9JMKHNp3_1(.din(n845), .dout(n1654));
    jdff dff_B_K8XvReoO8_1(.din(n436), .dout(n1658));
    jdff dff_B_esJ086AR6_0(.din(n683), .dout(n1661));
    jdff dff_A_IOZJOknJ8_0(.din(n1666), .dout(n1663));
    jdff dff_A_8aKTlphy4_0(.din(n1669), .dout(n1666));
    jdff dff_A_3fXteCz35_0(.din(n1672), .dout(n1669));
    jdff dff_A_DR3j0Nzw8_0(.din(n1675), .dout(n1672));
    jdff dff_A_ZNZawBni9_0(.din(n1678), .dout(n1675));
    jdff dff_A_MtDsypUi6_0(.din(n679), .dout(n1678));
    jdff dff_A_ISmlcl4W5_0(.din(n1684), .dout(n1681));
    jdff dff_A_QEWSt3uY8_0(.din(n1687), .dout(n1684));
    jdff dff_A_emJaql312_0(.din(n1690), .dout(n1687));
    jdff dff_A_tpC5tqD67_0(.din(n1693), .dout(n1690));
    jdff dff_A_qGfc80q32_0(.din(n1736), .dout(n1693));
    jdff dff_B_7WqDrcLp1_2(.din(n671), .dout(n1697));
    jdff dff_B_9ID2y5OB1_2(.din(n1697), .dout(n1700));
    jdff dff_B_yfSETw2Y7_2(.din(n1700), .dout(n1703));
    jdff dff_B_z9yi05R28_2(.din(n1703), .dout(n1706));
    jdff dff_B_fFJEMfJy2_2(.din(n1706), .dout(n1709));
    jdff dff_B_Ri7WhaH01_2(.din(n1709), .dout(n1712));
    jdff dff_B_RGAJpQ5v8_2(.din(n1712), .dout(n1715));
    jdff dff_B_PJRQGn585_2(.din(n1715), .dout(n1718));
    jdff dff_B_88KCtT4B9_2(.din(n1718), .dout(n1721));
    jdff dff_B_KXRq1A8e9_2(.din(n1721), .dout(n1724));
    jdff dff_B_w7y06zHV5_2(.din(n1724), .dout(n1727));
    jdff dff_B_BsuvV6W49_2(.din(n1727), .dout(n1730));
    jdff dff_B_ks6N9hNk0_2(.din(n1730), .dout(n1733));
    jdff dff_B_bgzYbinz7_2(.din(n1733), .dout(n1736));
    jdff dff_A_olLEk2cE6_0(.din(n1741), .dout(n1738));
    jdff dff_A_UbvmZKng4_0(.din(n1744), .dout(n1741));
    jdff dff_A_VRvNWvrO0_0(.din(n1747), .dout(n1744));
    jdff dff_A_4fTmYll73_0(.din(n1750), .dout(n1747));
    jdff dff_A_OWTt24nJ5_0(.din(n1753), .dout(n1750));
    jdff dff_A_dbQqSDnz1_0(.din(n660), .dout(n1753));
    jdff dff_A_RhOqGTS71_0(.din(n1759), .dout(n1756));
    jdff dff_A_Q5X4imaJ6_0(.din(n1762), .dout(n1759));
    jdff dff_A_kavg2DEy0_0(.din(n1765), .dout(n1762));
    jdff dff_A_0searHjC4_0(.din(n1768), .dout(n1765));
    jdff dff_A_seRwWBH32_0(.din(n1811), .dout(n1768));
    jdff dff_B_ZgxHQ6Hk4_2(.din(n652), .dout(n1772));
    jdff dff_B_bzAcanZg5_2(.din(n1772), .dout(n1775));
    jdff dff_B_PA8Pnz9I4_2(.din(n1775), .dout(n1778));
    jdff dff_B_OGPoxPg14_2(.din(n1778), .dout(n1781));
    jdff dff_B_t73EmK7g8_2(.din(n1781), .dout(n1784));
    jdff dff_B_eg2rpMol3_2(.din(n1784), .dout(n1787));
    jdff dff_B_RYjBlcNS3_2(.din(n1787), .dout(n1790));
    jdff dff_B_0GnCNoDc7_2(.din(n1790), .dout(n1793));
    jdff dff_B_xvkXV2VS7_2(.din(n1793), .dout(n1796));
    jdff dff_B_nFb1iLfC0_2(.din(n1796), .dout(n1799));
    jdff dff_B_JKd3r0gC1_2(.din(n1799), .dout(n1802));
    jdff dff_B_17S53n1d3_2(.din(n1802), .dout(n1805));
    jdff dff_B_IwNFJkjs7_2(.din(n1805), .dout(n1808));
    jdff dff_B_JHCPCgkZ6_2(.din(n1808), .dout(n1811));
    jdff dff_B_GDaQqjpP7_1(.din(n614), .dout(n1814));
    jdff dff_B_f2VOUnh55_1(.din(n1814), .dout(n1817));
    jdff dff_B_LUQePqha0_1(.din(n1817), .dout(n1820));
    jdff dff_B_SAF5a7wU9_1(.din(n1820), .dout(n1823));
    jdff dff_B_yKHAQ7bZ8_1(.din(n1823), .dout(n1826));
    jdff dff_B_X07PlIy63_1(.din(n1826), .dout(n1829));
    jdff dff_B_m65lksJo0_1(.din(n1829), .dout(n1832));
    jdff dff_B_0erNJKzh6_1(.din(n1832), .dout(n1835));
    jdff dff_B_iZMOoaEc6_1(.din(n1835), .dout(n1838));
    jdff dff_B_R9RicJHW6_1(.din(n1838), .dout(n1841));
    jdff dff_B_aDb6Ttog1_1(.din(n1841), .dout(n1844));
    jdff dff_B_m0F1ncWq9_1(.din(n1844), .dout(n1847));
    jdff dff_B_bw5EIPSK4_1(.din(n1847), .dout(n1850));
    jdff dff_B_XRoBwbH59_1(.din(n1850), .dout(n1853));
    jdff dff_B_bwo9Ndcl8_1(.din(n599), .dout(n1856));
    jdff dff_B_O2ProZuN1_1(.din(n1856), .dout(n1859));
    jdff dff_B_tDQLSqeZ0_1(.din(n1859), .dout(n1862));
    jdff dff_B_rnxsM0XU5_1(.din(n1862), .dout(n1865));
    jdff dff_B_hikrsU7Z5_1(.din(n1865), .dout(n1868));
    jdff dff_B_8IOPiCWU6_1(.din(n1868), .dout(n1871));
    jdff dff_B_4MbmWuke4_1(.din(n1871), .dout(n1874));
    jdff dff_B_KTg1yAft1_1(.din(n1874), .dout(n1877));
    jdff dff_B_XEkyDelF6_1(.din(n1877), .dout(n1880));
    jdff dff_B_9z3QR0bs6_1(.din(n1880), .dout(n1883));
    jdff dff_B_AftZ3Wo78_1(.din(n1883), .dout(n1886));
    jdff dff_B_7nSYDCnB8_1(.din(n1886), .dout(n1889));
    jdff dff_B_GotyeNsY1_1(.din(n1889), .dout(n1892));
    jdff dff_B_PlDjCZY22_1(.din(n1892), .dout(n1895));
    jdff dff_A_PiFD3WSk3_0(.din(n1900), .dout(n1897));
    jdff dff_A_OMLjdNpq0_0(.din(n1903), .dout(n1900));
    jdff dff_A_eBwg2Bxj9_0(.din(n1906), .dout(n1903));
    jdff dff_A_TLy8opGb5_0(.din(n1909), .dout(n1906));
    jdff dff_A_zvdmaR5U2_0(.din(n1952), .dout(n1909));
    jdff dff_B_QQbq5IlY3_2(.din(n580), .dout(n1913));
    jdff dff_B_OZd97weI4_2(.din(n1913), .dout(n1916));
    jdff dff_B_P5IQ1JFW2_2(.din(n1916), .dout(n1919));
    jdff dff_B_iunqsuTI3_2(.din(n1919), .dout(n1922));
    jdff dff_B_gtk4BpM27_2(.din(n1922), .dout(n1925));
    jdff dff_B_AOsJNhcZ1_2(.din(n1925), .dout(n1928));
    jdff dff_B_pzAcnuhG5_2(.din(n1928), .dout(n1931));
    jdff dff_B_Dbx0aZZD7_2(.din(n1931), .dout(n1934));
    jdff dff_B_MnC1J1qK4_2(.din(n1934), .dout(n1937));
    jdff dff_B_dcRO4kWi7_2(.din(n1937), .dout(n1940));
    jdff dff_B_cjtuyWXx7_2(.din(n1940), .dout(n1943));
    jdff dff_B_iyYNJnsV9_2(.din(n1943), .dout(n1946));
    jdff dff_B_1JorpXEE6_2(.din(n1946), .dout(n1949));
    jdff dff_B_y54Z7sHy7_2(.din(n1949), .dout(n1952));
    jdff dff_B_oiWBOB7h9_2(.din(n952), .dout(n1955));
    jdff dff_A_DgN3MSVq3_0(.din(n1960), .dout(n1957));
    jdff dff_A_82TKdms76_0(.din(n1963), .dout(n1960));
    jdff dff_A_3SzNbMJf1_0(.din(n1966), .dout(n1963));
    jdff dff_A_jeePaV4h6_0(.din(n1969), .dout(n1966));
    jdff dff_A_xnsN78VT8_0(.din(n2012), .dout(n1969));
    jdff dff_B_GIyhLYus5_2(.din(n439), .dout(n1973));
    jdff dff_B_PwQ2kG6V7_2(.din(n1973), .dout(n1976));
    jdff dff_B_ZbC8dhtR8_2(.din(n1976), .dout(n1979));
    jdff dff_B_2SXjRmGM2_2(.din(n1979), .dout(n1982));
    jdff dff_B_LvX2UqvK5_2(.din(n1982), .dout(n1985));
    jdff dff_B_BKDMNEAh6_2(.din(n1985), .dout(n1988));
    jdff dff_B_O2oHx9JX0_2(.din(n1988), .dout(n1991));
    jdff dff_B_3IVECn2B0_2(.din(n1991), .dout(n1994));
    jdff dff_B_B5gS4YMs9_2(.din(n1994), .dout(n1997));
    jdff dff_B_Laq60N2c5_2(.din(n1997), .dout(n2000));
    jdff dff_B_TO6m9H4P8_2(.din(n2000), .dout(n2003));
    jdff dff_B_R8eM2w5n0_2(.din(n2003), .dout(n2006));
    jdff dff_B_cEebf5uW0_2(.din(n2006), .dout(n2009));
    jdff dff_B_jl8Wcy995_2(.din(n2009), .dout(n2012));
    jdff dff_A_RM1anhUw6_0(.din(n2017), .dout(n2014));
    jdff dff_A_sKthbOZ28_0(.din(n2020), .dout(n2017));
    jdff dff_A_ZcZgjok87_0(.din(n2023), .dout(n2020));
    jdff dff_A_D2pY2psu8_0(.din(n2026), .dout(n2023));
    jdff dff_A_fMuf9xEt9_0(.din(n2029), .dout(n2026));
    jdff dff_A_8Dmcj8nY2_0(.din(n573), .dout(n2029));
    jdff dff_A_UtKslg8F9_0(.din(n2035), .dout(n2032));
    jdff dff_A_1hTnlo0v1_0(.din(n2038), .dout(n2035));
    jdff dff_A_frZW8Ixb0_0(.din(n913), .dout(n2038));
    jdff dff_B_ZhxoKhHD8_1(.din(n702), .dout(n2042));
    jdff dff_B_zJt6HAym3_0(.din(n805), .dout(n2045));
    jdff dff_A_WPTe1u9q5_0(.din(n2050), .dout(n2047));
    jdff dff_A_GSNYGnTk2_0(.din(n2053), .dout(n2050));
    jdff dff_A_kqEjlvSJ1_0(.din(n2056), .dout(n2053));
    jdff dff_A_VCL4iba75_0(.din(n2059), .dout(n2056));
    jdff dff_A_1w8blDM99_0(.din(n2062), .dout(n2059));
    jdff dff_A_qWk2rJrB6_0(.din(n2065), .dout(n2062));
    jdff dff_A_DzX34acp6_0(.din(n2068), .dout(n2065));
    jdff dff_A_aCCqTrBc7_0(.din(n2071), .dout(n2068));
    jdff dff_A_SWPagyCX3_0(.din(n2074), .dout(n2071));
    jdff dff_A_QTPwGdp08_0(.din(n2077), .dout(n2074));
    jdff dff_A_Rq4e2tBh2_0(.din(n2080), .dout(n2077));
    jdff dff_A_NxpvU0VK7_0(.din(n2083), .dout(n2080));
    jdff dff_A_wgEUhDkE2_0(.din(n2086), .dout(n2083));
    jdff dff_A_arkkcmbz7_0(.din(n2089), .dout(n2086));
    jdff dff_A_mAgQsyME8_0(.din(G27gat), .dout(n2089));
    jdff dff_A_kNAQRqxn5_0(.din(n2095), .dout(n2092));
    jdff dff_A_vY8QnSd14_0(.din(n2098), .dout(n2095));
    jdff dff_A_zzuNB8Ds1_0(.din(n2101), .dout(n2098));
    jdff dff_A_FAluccEs6_0(.din(n2104), .dout(n2101));
    jdff dff_A_1gshwirA9_0(.din(n2107), .dout(n2104));
    jdff dff_A_dxkrPtun8_0(.din(n2110), .dout(n2107));
    jdff dff_A_u6BXhCcu8_0(.din(n2113), .dout(n2110));
    jdff dff_A_bsEdBsHB3_0(.din(n2116), .dout(n2113));
    jdff dff_A_UOSQooNn3_0(.din(n2119), .dout(n2116));
    jdff dff_A_1B5QYVXI4_0(.din(n2122), .dout(n2119));
    jdff dff_A_XJLVieiL0_0(.din(n2125), .dout(n2122));
    jdff dff_A_jFB0XQEE4_0(.din(n2128), .dout(n2125));
    jdff dff_A_UP0ZRpiA9_0(.din(n2131), .dout(n2128));
    jdff dff_A_iuNc7Xhb9_0(.din(n2134), .dout(n2131));
    jdff dff_A_HRDrLIPA2_0(.din(G115gat), .dout(n2134));
    jdff dff_A_yzk0Ipx60_0(.din(n2140), .dout(n2137));
    jdff dff_A_RAmVZyC48_0(.din(n2143), .dout(n2140));
    jdff dff_A_n93NZ9wV0_0(.din(n2146), .dout(n2143));
    jdff dff_A_ITq3EleO6_0(.din(n2149), .dout(n2146));
    jdff dff_A_mCrN3Lj91_0(.din(n2152), .dout(n2149));
    jdff dff_A_4hKeouNQ8_0(.din(n753), .dout(n2152));
    jdff dff_A_CQcrHCBb6_0(.din(n2158), .dout(n2155));
    jdff dff_A_C1l3zL6B5_0(.din(n2161), .dout(n2158));
    jdff dff_A_YD7hr8tY0_0(.din(n2164), .dout(n2161));
    jdff dff_A_i0KCF6q20_0(.din(n2167), .dout(n2164));
    jdff dff_A_4dtMxGzU6_0(.din(n2170), .dout(n2167));
    jdff dff_A_z1qq2N689_0(.din(n2173), .dout(n2170));
    jdff dff_A_cDTPGoMq9_0(.din(n2176), .dout(n2173));
    jdff dff_A_ieM7F0Qu8_0(.din(n2179), .dout(n2176));
    jdff dff_A_z9Dm9cNI4_0(.din(n2182), .dout(n2179));
    jdff dff_A_bNf7nTdS6_0(.din(n2185), .dout(n2182));
    jdff dff_A_67IY7bF71_0(.din(n2188), .dout(n2185));
    jdff dff_A_KCe3CFxT9_0(.din(n2191), .dout(n2188));
    jdff dff_A_V9xet9mD8_0(.din(n2194), .dout(n2191));
    jdff dff_A_Ce1tMWSv9_0(.din(n2197), .dout(n2194));
    jdff dff_A_lorB278v7_0(.din(n2200), .dout(n2197));
    jdff dff_A_8sSn4NmT8_0(.din(n2203), .dout(n2200));
    jdff dff_A_TPK5Ey768_0(.din(n2206), .dout(n2203));
    jdff dff_A_1LZv9Un12_0(.din(n2209), .dout(n2206));
    jdff dff_A_loKggvBq6_0(.din(n2212), .dout(n2209));
    jdff dff_A_FEf1B7nZ7_0(.din(G92gat), .dout(n2212));
    jdff dff_A_2uLs2c3S9_1(.din(n2218), .dout(n2215));
    jdff dff_A_AhuKunsi1_1(.din(n2221), .dout(n2218));
    jdff dff_A_pcFbUBcz9_1(.din(n2224), .dout(n2221));
    jdff dff_A_s3eF31HN8_1(.din(n2227), .dout(n2224));
    jdff dff_A_MsmPoJDb8_1(.din(n2230), .dout(n2227));
    jdff dff_A_Xfxgwyf14_1(.din(n2233), .dout(n2230));
    jdff dff_A_FFB9MV8l1_1(.din(n2236), .dout(n2233));
    jdff dff_A_LVJrnfm42_1(.din(n2239), .dout(n2236));
    jdff dff_A_14DWDvVg9_1(.din(n2242), .dout(n2239));
    jdff dff_A_3upgWeKT5_1(.din(n2245), .dout(n2242));
    jdff dff_A_kTp2LQFU5_1(.din(n2248), .dout(n2245));
    jdff dff_A_b2buw0UU4_1(.din(n2251), .dout(n2248));
    jdff dff_A_OGEALcHA6_1(.din(n2254), .dout(n2251));
    jdff dff_A_MxjzSkw00_1(.din(n2257), .dout(n2254));
    jdff dff_A_PWYb19Y21_1(.din(G92gat), .dout(n2257));
    jdff dff_A_f59jYA8P5_0(.din(n2263), .dout(n2260));
    jdff dff_A_pRmMQpeE8_0(.din(n2266), .dout(n2263));
    jdff dff_A_QIn5Lzi67_0(.din(n2269), .dout(n2266));
    jdff dff_A_AjrOsry46_0(.din(n2272), .dout(n2269));
    jdff dff_A_Qx88tkmG9_0(.din(n2275), .dout(n2272));
    jdff dff_A_l6vhJiZM3_0(.din(n741), .dout(n2275));
    jdff dff_A_isqtWgis2_0(.din(n2281), .dout(n2278));
    jdff dff_A_ITwmwsQp0_0(.din(n2284), .dout(n2281));
    jdff dff_A_wBFge4ko1_0(.din(n2287), .dout(n2284));
    jdff dff_A_ZxDfTi8f3_0(.din(n2290), .dout(n2287));
    jdff dff_A_wwlGmWnf0_0(.din(n2293), .dout(n2290));
    jdff dff_A_yTO17ioo5_0(.din(n2296), .dout(n2293));
    jdff dff_A_Cw8fn0Qz3_0(.din(n2299), .dout(n2296));
    jdff dff_A_Dgi3RNPu2_0(.din(n2302), .dout(n2299));
    jdff dff_A_tOFYThyM9_0(.din(n2305), .dout(n2302));
    jdff dff_A_AUmjnKpy6_0(.din(n2308), .dout(n2305));
    jdff dff_A_kz696BsN3_0(.din(n2311), .dout(n2308));
    jdff dff_A_PsC3Z56w8_0(.din(n2314), .dout(n2311));
    jdff dff_A_32rDj0y51_0(.din(n2317), .dout(n2314));
    jdff dff_A_awSD8oBC8_0(.din(n2320), .dout(n2317));
    jdff dff_A_bMTPEd8B3_0(.din(n2323), .dout(n2320));
    jdff dff_A_KgaLiSJk5_0(.din(n2326), .dout(n2323));
    jdff dff_A_SifZUAWh9_0(.din(n2329), .dout(n2326));
    jdff dff_A_WB3qmmwu6_0(.din(n2332), .dout(n2329));
    jdff dff_A_1mWI1GVB8_0(.din(n2335), .dout(n2332));
    jdff dff_A_X7CJlDZg1_0(.din(G14gat), .dout(n2335));
    jdff dff_A_HjH7T54d8_1(.din(n2341), .dout(n2338));
    jdff dff_A_Jjd5WVeh4_1(.din(n2344), .dout(n2341));
    jdff dff_A_vzidcSnN8_1(.din(n2347), .dout(n2344));
    jdff dff_A_0BDYz8ZI6_1(.din(n2350), .dout(n2347));
    jdff dff_A_dSPJwEna1_1(.din(n2353), .dout(n2350));
    jdff dff_A_wA5Uq0Mn6_1(.din(n2356), .dout(n2353));
    jdff dff_A_CmdJG8Ph9_1(.din(n2359), .dout(n2356));
    jdff dff_A_CzKBE1lf3_1(.din(n2362), .dout(n2359));
    jdff dff_A_J9fnEt7q1_1(.din(n2365), .dout(n2362));
    jdff dff_A_s4X9JNUG4_1(.din(n2368), .dout(n2365));
    jdff dff_A_6TGauh890_1(.din(n2371), .dout(n2368));
    jdff dff_A_4bV3bnYD5_1(.din(n2374), .dout(n2371));
    jdff dff_A_eSG4JE0Y4_1(.din(n2377), .dout(n2374));
    jdff dff_A_cyGpAo5m7_1(.din(n2380), .dout(n2377));
    jdff dff_A_zfRanZFb5_1(.din(G14gat), .dout(n2380));
    jdff dff_B_Vv1U1Xsw1_1(.din(n717), .dout(n2384));
    jdff dff_B_8QAkKt3M0_1(.din(n2384), .dout(n2387));
    jdff dff_B_355MOtrO4_1(.din(n2387), .dout(n2390));
    jdff dff_B_it2znLd43_1(.din(n2390), .dout(n2393));
    jdff dff_B_NyDAsDHa5_1(.din(n2393), .dout(n2396));
    jdff dff_A_ly6rZopT4_0(.din(n2401), .dout(n2398));
    jdff dff_A_gyXE4MHt9_0(.din(n2404), .dout(n2401));
    jdff dff_A_iWtpklWD3_0(.din(n2407), .dout(n2404));
    jdff dff_A_ukOAbM1O3_0(.din(n2410), .dout(n2407));
    jdff dff_A_KHlim5GW8_0(.din(n2413), .dout(n2410));
    jdff dff_A_o4Gn8Rp16_0(.din(n2416), .dout(n2413));
    jdff dff_A_htKJlJg06_0(.din(n2419), .dout(n2416));
    jdff dff_A_iyv5sVN33_0(.din(n2422), .dout(n2419));
    jdff dff_A_jUuZdhSc6_0(.din(n2425), .dout(n2422));
    jdff dff_A_qUxF57Qh6_0(.din(n2428), .dout(n2425));
    jdff dff_A_Q9c17TY98_0(.din(n2431), .dout(n2428));
    jdff dff_A_xKPOWsTF8_0(.din(n2434), .dout(n2431));
    jdff dff_A_C3dt0v0v1_0(.din(n2437), .dout(n2434));
    jdff dff_A_FZnNBvdh3_0(.din(n2440), .dout(n2437));
    jdff dff_A_xWYS2Qnl3_0(.din(n2443), .dout(n2440));
    jdff dff_A_WUcUq3Y59_0(.din(n2446), .dout(n2443));
    jdff dff_A_8TKz3JAl9_0(.din(n2449), .dout(n2446));
    jdff dff_A_hMc6BZEG9_0(.din(n2452), .dout(n2449));
    jdff dff_A_Qp1Rk47H9_0(.din(n2455), .dout(n2452));
    jdff dff_A_pw1kHjUz2_0(.din(G66gat), .dout(n2455));
    jdff dff_A_6mPWo1Ja7_1(.din(n2461), .dout(n2458));
    jdff dff_A_b0eEEZzx3_1(.din(n2464), .dout(n2461));
    jdff dff_A_RChVbdHd9_1(.din(n2467), .dout(n2464));
    jdff dff_A_Ug4oAg0y9_1(.din(n2470), .dout(n2467));
    jdff dff_A_CpzthAVL9_1(.din(n2473), .dout(n2470));
    jdff dff_A_r3ILZe7g6_1(.din(n2476), .dout(n2473));
    jdff dff_A_jco5sZSn2_1(.din(n2479), .dout(n2476));
    jdff dff_A_tBcWuE1L0_1(.din(n2482), .dout(n2479));
    jdff dff_A_f9fvTdNm4_1(.din(n2485), .dout(n2482));
    jdff dff_A_RzDsK4NF5_1(.din(n2488), .dout(n2485));
    jdff dff_A_ymJMnyH77_1(.din(n2491), .dout(n2488));
    jdff dff_A_8JAKO9mK3_1(.din(n2494), .dout(n2491));
    jdff dff_A_JpuSwqI38_1(.din(n2497), .dout(n2494));
    jdff dff_A_TlcIV72U0_1(.din(n2500), .dout(n2497));
    jdff dff_A_EGfukxDR9_1(.din(G66gat), .dout(n2500));
    jdff dff_A_IYKTXbQ26_0(.din(n2506), .dout(n2503));
    jdff dff_A_3MUahvAy4_0(.din(n2509), .dout(n2506));
    jdff dff_A_YYeBLsx88_0(.din(n2512), .dout(n2509));
    jdff dff_A_VYWMwE812_0(.din(n2515), .dout(n2512));
    jdff dff_A_CmjLWyko3_0(.din(n2518), .dout(n2515));
    jdff dff_A_9zRzmdzM7_0(.din(n2521), .dout(n2518));
    jdff dff_A_SyYmKoxZ3_0(.din(n2524), .dout(n2521));
    jdff dff_A_cU0uybh90_0(.din(n2527), .dout(n2524));
    jdff dff_A_FClwhfiw9_0(.din(n2530), .dout(n2527));
    jdff dff_A_gUxxbEq39_0(.din(n2533), .dout(n2530));
    jdff dff_A_Ee5Gfiu55_0(.din(n2536), .dout(n2533));
    jdff dff_A_MFKm1KjX7_0(.din(n2539), .dout(n2536));
    jdff dff_A_1MGRnFlX9_0(.din(n2542), .dout(n2539));
    jdff dff_A_rBTwsf5d4_0(.din(n2545), .dout(n2542));
    jdff dff_A_KwV5G41l5_0(.din(G40gat), .dout(n2545));
    jdff dff_A_XQDfzSS13_1(.din(n432), .dout(n2548));
    jdff dff_B_fpzEPT5I7_0(.din(n428), .dout(n2552));
    jdff dff_B_m25x534I1_0(.din(n2552), .dout(n2555));
    jdff dff_B_7DzAXQHl2_0(.din(n2555), .dout(n2558));
    jdff dff_B_LUBtFMM42_0(.din(n2558), .dout(n2561));
    jdff dff_B_JCNH5Y7g8_0(.din(n2561), .dout(n2564));
    jdff dff_B_VFPT1eVQ5_0(.din(n2564), .dout(n2567));
    jdff dff_A_cAgb6sJp5_0(.din(n2572), .dout(n2569));
    jdff dff_A_UwRY90fB9_0(.din(n2575), .dout(n2572));
    jdff dff_A_oy9L780f9_0(.din(n2578), .dout(n2575));
    jdff dff_A_YZGk8nx20_0(.din(n2581), .dout(n2578));
    jdff dff_A_XGUntYs56_0(.din(n2584), .dout(n2581));
    jdff dff_A_83uB0iM15_0(.din(n2587), .dout(n2584));
    jdff dff_A_HlQglHUY2_0(.din(n2590), .dout(n2587));
    jdff dff_A_bF9J1icF2_0(.din(n2593), .dout(n2590));
    jdff dff_A_vDrPrNMf5_0(.din(n2596), .dout(n2593));
    jdff dff_A_zbeykTCV7_0(.din(n2599), .dout(n2596));
    jdff dff_A_AsDAUV2P7_0(.din(n2602), .dout(n2599));
    jdff dff_A_MDnOkpYB1_0(.din(n2624), .dout(n2602));
    jdff dff_B_A5e2h8VR1_2(.din(n424), .dout(n2606));
    jdff dff_B_YI0AwNSz6_2(.din(n2606), .dout(n2609));
    jdff dff_B_2X8y0zbI3_2(.din(n2609), .dout(n2612));
    jdff dff_B_3tLIWoyx4_2(.din(n2612), .dout(n2615));
    jdff dff_B_ygig0ASU9_2(.din(n2615), .dout(n2618));
    jdff dff_B_VUJKNZ2w6_2(.din(n2618), .dout(n2621));
    jdff dff_B_1M8i8mw79_2(.din(n2621), .dout(n2624));
    jdff dff_A_TehYMzBl8_0(.din(n2629), .dout(n2626));
    jdff dff_A_Fn7Iv4Cx7_0(.din(n2632), .dout(n2629));
    jdff dff_A_HE2idggS8_0(.din(n2635), .dout(n2632));
    jdff dff_A_yrQ2Xsar7_0(.din(n2638), .dout(n2635));
    jdff dff_A_2vSLHRkS3_0(.din(n2641), .dout(n2638));
    jdff dff_A_2iqLDpq24_0(.din(n2644), .dout(n2641));
    jdff dff_A_OsNwv2H67_0(.din(n2647), .dout(n2644));
    jdff dff_A_KBGWrlXH4_0(.din(n2650), .dout(n2647));
    jdff dff_A_2c9lvAsF9_0(.din(n2653), .dout(n2650));
    jdff dff_A_4C9omT440_0(.din(n2656), .dout(n2653));
    jdff dff_A_9n1BOoKH9_0(.din(n2659), .dout(n2656));
    jdff dff_A_HDcVbxuz4_0(.din(n2662), .dout(n2659));
    jdff dff_A_3z2JhcZs3_0(.din(n2665), .dout(n2662));
    jdff dff_A_FMq6roSG4_0(.din(n2668), .dout(n2665));
    jdff dff_A_7U1ypy1a6_0(.din(n2671), .dout(n2668));
    jdff dff_A_WpQyq9FU3_0(.din(n2674), .dout(n2671));
    jdff dff_A_0X4VuQBb3_0(.din(n2677), .dout(n2674));
    jdff dff_A_4KdI0J6J9_0(.din(n2680), .dout(n2677));
    jdff dff_A_NXAvvox10_0(.din(n2683), .dout(n2680));
    jdff dff_A_rA6U099P1_0(.din(G53gat), .dout(n2683));
    jdff dff_A_iZIDpyIr3_0(.din(n411), .dout(n2686));
    jdff dff_B_NqK5r0uJ8_1(.din(n345), .dout(n2690));
    jdff dff_B_KqJio3Rg4_1(.din(n363), .dout(n2693));
    jdff dff_B_pYwWI0Mm8_1(.din(n2693), .dout(n2696));
    jdff dff_B_ka8Zgljp4_1(.din(n2696), .dout(n2699));
    jdff dff_B_Fyq44NgT7_1(.din(n2699), .dout(n2702));
    jdff dff_B_ZdKfvdf30_1(.din(n2702), .dout(n2705));
    jdff dff_B_447HS49Y5_1(.din(n2705), .dout(n2708));
    jdff dff_B_vJDXMRpC0_1(.din(n2708), .dout(n2711));
    jdff dff_A_ukWOq8tP3_0(.din(n2716), .dout(n2713));
    jdff dff_A_YYqfWhRq9_0(.din(n2719), .dout(n2716));
    jdff dff_A_CXIqUqbt1_0(.din(n2722), .dout(n2719));
    jdff dff_A_Rmm5znAV3_0(.din(n2725), .dout(n2722));
    jdff dff_A_iLzFQlOm1_0(.din(n2728), .dout(n2725));
    jdff dff_A_o9WJ33q89_0(.din(n2731), .dout(n2728));
    jdff dff_A_fnI5mclx4_0(.din(n371), .dout(n2731));
    jdff dff_A_DcKErPU78_0(.din(n2737), .dout(n2734));
    jdff dff_A_oBfutAC63_0(.din(n2740), .dout(n2737));
    jdff dff_A_BVrgXk641_0(.din(n2743), .dout(n2740));
    jdff dff_A_GtwakSja0_0(.din(n2746), .dout(n2743));
    jdff dff_A_8y8N3Guq4_0(.din(n2749), .dout(n2746));
    jdff dff_A_j1MTcUuX6_0(.din(n356), .dout(n2749));
    jdff dff_A_BTCMwIhv4_0(.din(n2755), .dout(n2752));
    jdff dff_A_0vTTxGiD2_0(.din(n2758), .dout(n2755));
    jdff dff_A_YR1Vi4Ty3_0(.din(n2761), .dout(n2758));
    jdff dff_A_uIcAZ2sq8_0(.din(n2764), .dout(n2761));
    jdff dff_A_sOSeQPg69_0(.din(n2786), .dout(n2764));
    jdff dff_B_ppkxjZnz4_2(.din(n348), .dout(n2768));
    jdff dff_B_MvqA1pyZ4_2(.din(n2768), .dout(n2771));
    jdff dff_B_nYPoKPki5_2(.din(n2771), .dout(n2774));
    jdff dff_B_Z878v3sO5_2(.din(n2774), .dout(n2777));
    jdff dff_B_bzuIyA295_2(.din(n2777), .dout(n2780));
    jdff dff_B_NgIky2cZ8_2(.din(n2780), .dout(n2783));
    jdff dff_B_jlkyKIwC3_2(.din(n2783), .dout(n2786));
    jdff dff_A_t0fwS1Fi4_0(.din(n2791), .dout(n2788));
    jdff dff_A_eBAMU7Fu8_0(.din(n2794), .dout(n2791));
    jdff dff_A_qiARuj7l3_0(.din(n2797), .dout(n2794));
    jdff dff_A_Fx7tNW6C3_0(.din(n2800), .dout(n2797));
    jdff dff_A_KQeLt5oc7_0(.din(n2803), .dout(n2800));
    jdff dff_A_yXhG2H8g8_0(.din(n341), .dout(n2803));
    jdff dff_A_PNEJJfWC8_0(.din(n2809), .dout(n2806));
    jdff dff_A_iXm02h9u9_0(.din(n2812), .dout(n2809));
    jdff dff_A_ZJXP5Yfj7_0(.din(n2815), .dout(n2812));
    jdff dff_A_UGzvVhbG3_0(.din(n2818), .dout(n2815));
    jdff dff_A_TNwq3u6B6_0(.din(n2840), .dout(n2818));
    jdff dff_B_IOWr197e6_2(.din(n333), .dout(n2822));
    jdff dff_B_OkO0mU4i5_2(.din(n2822), .dout(n2825));
    jdff dff_B_JbGIOMH40_2(.din(n2825), .dout(n2828));
    jdff dff_B_L9v1PK3V0_2(.din(n2828), .dout(n2831));
    jdff dff_B_uW5GfRcs4_2(.din(n2831), .dout(n2834));
    jdff dff_B_s9Nl5gDw7_2(.din(n2834), .dout(n2837));
    jdff dff_B_aWMZslLJ7_2(.din(n2837), .dout(n2840));
    jdff dff_B_tFxJeg604_1(.din(n258), .dout(n2843));
    jdff dff_B_kNpHvdbT1_0(.din(n307), .dout(n2846));
    jdff dff_A_wK59n6K32_0(.din(n2851), .dout(n2848));
    jdff dff_A_Fot6INnu1_0(.din(n2854), .dout(n2851));
    jdff dff_A_m4w3asQE4_0(.din(n2857), .dout(n2854));
    jdff dff_A_ep4zO53T7_0(.din(n2860), .dout(n2857));
    jdff dff_A_jNCJ47D70_0(.din(n2863), .dout(n2860));
    jdff dff_A_jvJV2ZFZ2_0(.din(n303), .dout(n2863));
    jdff dff_A_q0VOqsmD5_0(.din(n2869), .dout(n2866));
    jdff dff_A_oYvf3OG94_0(.din(n2872), .dout(n2869));
    jdff dff_A_qPPMUy726_0(.din(n2875), .dout(n2872));
    jdff dff_A_7Lu1vTHu9_0(.din(n2878), .dout(n2875));
    jdff dff_A_mLXAvt4n0_0(.din(n2900), .dout(n2878));
    jdff dff_B_b4dbHZai5_2(.din(n295), .dout(n2882));
    jdff dff_B_eurmNImh1_2(.din(n2882), .dout(n2885));
    jdff dff_B_Yp7sK7kU0_2(.din(n2885), .dout(n2888));
    jdff dff_B_FEn4Q8Yo7_2(.din(n2888), .dout(n2891));
    jdff dff_B_TVEWEfFY6_2(.din(n2891), .dout(n2894));
    jdff dff_B_MJmaSI9H1_2(.din(n2894), .dout(n2897));
    jdff dff_B_kRvHPEm09_2(.din(n2897), .dout(n2900));
    jdff dff_A_iJzAqBOW0_0(.din(n2905), .dout(n2902));
    jdff dff_A_UBAr06oW3_0(.din(n2908), .dout(n2905));
    jdff dff_A_zLWEIj8B8_0(.din(n2911), .dout(n2908));
    jdff dff_A_19qyuNKG3_0(.din(n2914), .dout(n2911));
    jdff dff_A_eMNfuXmO1_0(.din(n2917), .dout(n2914));
    jdff dff_A_XMNTUH095_0(.din(n284), .dout(n2917));
    jdff dff_A_hB2DIHX84_0(.din(n2923), .dout(n2920));
    jdff dff_A_tUk0OBpo4_0(.din(n2926), .dout(n2923));
    jdff dff_A_QdaKPHcP5_0(.din(n2929), .dout(n2926));
    jdff dff_A_Wkzy1KtS0_0(.din(n2932), .dout(n2929));
    jdff dff_A_V88cwFC23_0(.din(n2954), .dout(n2932));
    jdff dff_B_dA3SBpJ68_2(.din(n276), .dout(n2936));
    jdff dff_B_G1ZeSt958_2(.din(n2936), .dout(n2939));
    jdff dff_B_3aBa0O241_2(.din(n2939), .dout(n2942));
    jdff dff_B_Wus2GaKB4_2(.din(n2942), .dout(n2945));
    jdff dff_B_5oAjXXeq8_2(.din(n2945), .dout(n2948));
    jdff dff_B_U9Vb01T34_2(.din(n2948), .dout(n2951));
    jdff dff_B_93DoIoKW3_2(.din(n2951), .dout(n2954));
    jdff dff_B_4Hy0jiv52_1(.din(n242), .dout(n2957));
    jdff dff_B_ecmWlFWi7_1(.din(n2957), .dout(n2960));
    jdff dff_B_hhc665Rx5_1(.din(n2960), .dout(n2963));
    jdff dff_B_AnQhNxo99_1(.din(n2963), .dout(n2966));
    jdff dff_B_DQXU00sF7_1(.din(n2966), .dout(n2969));
    jdff dff_B_djL2IWfi4_1(.din(n2969), .dout(n2972));
    jdff dff_B_awY5TtCk8_1(.din(n2972), .dout(n2975));
    jdff dff_A_0gGFO1si5_0(.din(n2980), .dout(n2977));
    jdff dff_A_w5VXco6n2_0(.din(n2983), .dout(n2980));
    jdff dff_A_O5BubKlF6_0(.din(n2986), .dout(n2983));
    jdff dff_A_uvZBCxhN2_0(.din(n2989), .dout(n2986));
    jdff dff_A_IbJJYA8K7_0(.din(n2992), .dout(n2989));
    jdff dff_A_cRMZYc3B1_0(.din(n235), .dout(n2992));
    jdff dff_A_dAdDwizU1_0(.din(n2998), .dout(n2995));
    jdff dff_A_cIgXDEL30_0(.din(n3001), .dout(n2998));
    jdff dff_A_1e8abMSn7_0(.din(n3004), .dout(n3001));
    jdff dff_A_yCXfxgGn8_0(.din(n3007), .dout(n3004));
    jdff dff_A_dM4HeqPw5_0(.din(n3029), .dout(n3007));
    jdff dff_B_7S11WjdZ4_2(.din(n143), .dout(n3011));
    jdff dff_B_CXrh2OYW4_2(.din(n3011), .dout(n3014));
    jdff dff_B_6Cbbxs066_2(.din(n3014), .dout(n3017));
    jdff dff_B_nZFvdqNt7_2(.din(n3017), .dout(n3020));
    jdff dff_B_ubgIpsNP6_2(.din(n3020), .dout(n3023));
    jdff dff_B_WMzIhlvR0_2(.din(n3023), .dout(n3026));
    jdff dff_B_du5n4KHy9_2(.din(n3026), .dout(n3029));
    jdff dff_A_HsvVj9Sr9_1(.din(n3034), .dout(n3031));
    jdff dff_A_GfVaUSdR8_1(.din(n3037), .dout(n3034));
    jdff dff_A_TazNC8XV7_1(.din(n3040), .dout(n3037));
    jdff dff_A_QCoJQIcB1_1(.din(n3043), .dout(n3040));
    jdff dff_A_efO9Ivv29_1(.din(n3046), .dout(n3043));
    jdff dff_A_TLOHSE780_1(.din(n3049), .dout(n3046));
    jdff dff_A_gevF5jCx6_1(.din(n3052), .dout(n3049));
    jdff dff_A_W2xbkyoo0_1(.din(n3055), .dout(n3052));
    jdff dff_A_kPjP12Jp9_1(.din(n3058), .dout(n3055));
    jdff dff_A_DrfipQrw9_1(.din(n3061), .dout(n3058));
    jdff dff_A_KAZwzF9R4_1(.din(n3064), .dout(n3061));
    jdff dff_A_qrbowgNY3_1(.din(n3067), .dout(n3064));
    jdff dff_A_RC5qWVzk6_1(.din(n3070), .dout(n3067));
    jdff dff_A_SbUyfcqN9_1(.din(n3073), .dout(n3070));
    jdff dff_A_UzWk0GRm9_1(.din(G105gat), .dout(n3073));
    jdff dff_A_rN8koomI5_0(.din(n3079), .dout(n3076));
    jdff dff_A_PzEU658U9_0(.din(n3082), .dout(n3079));
    jdff dff_A_mOfbwand3_0(.din(n3085), .dout(n3082));
    jdff dff_A_AkUplPZz5_0(.din(n3088), .dout(n3085));
    jdff dff_A_UkbINEYs0_0(.din(n3131), .dout(n3088));
    jdff dff_B_i0JwDmKu3_2(.din(n637), .dout(n3092));
    jdff dff_B_nkkH4yCR3_2(.din(n3092), .dout(n3095));
    jdff dff_B_4zpay2Qy5_2(.din(n3095), .dout(n3098));
    jdff dff_B_1gHkALnk9_2(.din(n3098), .dout(n3101));
    jdff dff_B_cqrnNfOR2_2(.din(n3101), .dout(n3104));
    jdff dff_B_P2897u1Q3_2(.din(n3104), .dout(n3107));
    jdff dff_B_IaRzRIba6_2(.din(n3107), .dout(n3110));
    jdff dff_B_Q13EOOKL1_2(.din(n3110), .dout(n3113));
    jdff dff_B_1GMVD8i19_2(.din(n3113), .dout(n3116));
    jdff dff_B_J8W4Nmss9_2(.din(n3116), .dout(n3119));
    jdff dff_B_hbK7XanY0_2(.din(n3119), .dout(n3122));
    jdff dff_B_180tNT1g1_2(.din(n3122), .dout(n3125));
    jdff dff_B_KfyEUUMm8_2(.din(n3125), .dout(n3128));
    jdff dff_B_jWf3GUkZ9_2(.din(n3128), .dout(n3131));
    jdff dff_A_QD8Sn8xn6_0(.din(n3136), .dout(n3133));
    jdff dff_A_hnXEFaRo3_0(.din(n3139), .dout(n3136));
    jdff dff_A_ubLSppHX7_0(.din(n3142), .dout(n3139));
    jdff dff_A_fChuHLr85_0(.din(n3145), .dout(n3142));
    jdff dff_A_p5a7Vwgh8_0(.din(n3148), .dout(n3145));
    jdff dff_A_gj7DxBKd2_0(.din(n3151), .dout(n3148));
    jdff dff_A_xuEWtplg7_0(.din(n3154), .dout(n3151));
    jdff dff_A_gHCh00wX9_0(.din(n3157), .dout(n3154));
    jdff dff_A_56IQBdFD6_0(.din(n3160), .dout(n3157));
    jdff dff_A_Ntc4VIEX7_0(.din(n3163), .dout(n3160));
    jdff dff_A_UCyxuw599_0(.din(n3166), .dout(n3163));
    jdff dff_A_sPIJUNzg2_0(.din(n3169), .dout(n3166));
    jdff dff_A_fwbZKcqG5_0(.din(n3172), .dout(n3169));
    jdff dff_A_5Rzh4lej4_0(.din(n3175), .dout(n3172));
    jdff dff_A_PkvW4NuJ6_0(.din(G79gat), .dout(n3175));
    jdff dff_A_IQsc8pdn6_0(.din(n3181), .dout(n3178));
    jdff dff_A_qx6bSRxL0_0(.din(n3184), .dout(n3181));
    jdff dff_A_1ZnpfZau8_0(.din(n3187), .dout(n3184));
    jdff dff_A_eYlnGbmT1_0(.din(n3190), .dout(n3187));
    jdff dff_A_YZFvLYFV8_0(.din(n3193), .dout(n3190));
    jdff dff_A_4ovGi05V3_0(.din(n645), .dout(n3193));
    jdff dff_B_NQ6qWZcn7_1(.din(n513), .dout(n3197));
    jdff dff_B_MGjLvvx48_1(.din(n525), .dout(n3200));
    jdff dff_A_azkryNac6_0(.din(n3205), .dout(n3202));
    jdff dff_A_NU4en6Er5_0(.din(n3208), .dout(n3205));
    jdff dff_A_4Obfc4wf3_0(.din(n3211), .dout(n3208));
    jdff dff_A_TwTZHlF69_0(.din(n3214), .dout(n3211));
    jdff dff_A_jyiK3bZm1_0(.din(n3217), .dout(n3214));
    jdff dff_A_hGZTRHHC4_0(.din(n3220), .dout(n3217));
    jdff dff_A_CphBLeP64_0(.din(n3223), .dout(n3220));
    jdff dff_A_6LwEWqdP7_0(.din(G47gat), .dout(n3223));
    jdff dff_A_d3psj1Pa9_1(.din(n3229), .dout(n3226));
    jdff dff_A_jn0pbfpr1_1(.din(n3232), .dout(n3229));
    jdff dff_A_G66HetqF0_1(.din(n3235), .dout(n3232));
    jdff dff_A_2DcnsPvc6_1(.din(n3238), .dout(n3235));
    jdff dff_A_LL1Dh6kU8_1(.din(n3241), .dout(n3238));
    jdff dff_A_my1kK3pL0_1(.din(n3244), .dout(n3241));
    jdff dff_A_ofCS9CID6_1(.din(n3247), .dout(n3244));
    jdff dff_A_T6pXnsGV7_1(.din(n3250), .dout(n3247));
    jdff dff_A_AH4PL5i43_1(.din(n3253), .dout(n3250));
    jdff dff_A_i4JLvFh20_1(.din(n3256), .dout(n3253));
    jdff dff_A_m22eKOdL3_1(.din(n3259), .dout(n3256));
    jdff dff_A_ETi4jrU66_1(.din(n3262), .dout(n3259));
    jdff dff_A_JLloTRJ83_1(.din(G47gat), .dout(n3262));
    jdff dff_A_gnRA4fNu1_0(.din(n3268), .dout(n3265));
    jdff dff_A_7cwWfYfj1_0(.din(n3271), .dout(n3268));
    jdff dff_A_tF4grip08_0(.din(n3274), .dout(n3271));
    jdff dff_A_yEMOP4rc7_0(.din(n3277), .dout(n3274));
    jdff dff_A_7o0mONMx5_0(.din(n3280), .dout(n3277));
    jdff dff_A_Z6xDi7py5_0(.din(n533), .dout(n3280));
    jdff dff_A_keSjFFSW4_0(.din(n3286), .dout(n3283));
    jdff dff_A_FmMZyJLw4_0(.din(n3289), .dout(n3286));
    jdff dff_A_GQSUqkXk1_0(.din(n3292), .dout(n3289));
    jdff dff_A_0GQ949Hm5_0(.din(n3295), .dout(n3292));
    jdff dff_A_5LXmG0EF7_0(.din(n3298), .dout(n3295));
    jdff dff_A_OkcAVjAQ3_0(.din(n3301), .dout(n3298));
    jdff dff_A_7ZIDyrBl4_0(.din(n3304), .dout(n3301));
    jdff dff_A_tJnszgV80_0(.din(n3307), .dout(n3304));
    jdff dff_A_5K6pCmpL2_0(.din(n3310), .dout(n3307));
    jdff dff_A_e9MGPYqX1_0(.din(n3313), .dout(n3310));
    jdff dff_A_MP349w4b3_0(.din(n3316), .dout(n3313));
    jdff dff_A_F67Yb6UX5_0(.din(n3319), .dout(n3316));
    jdff dff_A_Le75QP4r4_0(.din(G8gat), .dout(n3319));
    jdff dff_A_d0c6zVx68_1(.din(n3325), .dout(n3322));
    jdff dff_A_7n9lGIWn3_1(.din(n3328), .dout(n3325));
    jdff dff_A_fBde5rFb6_1(.din(n3331), .dout(n3328));
    jdff dff_A_I8xSQwyx5_1(.din(n3334), .dout(n3331));
    jdff dff_A_sDy1bD010_1(.din(n3337), .dout(n3334));
    jdff dff_A_8JQYqsyZ2_1(.din(n3340), .dout(n3337));
    jdff dff_A_zm39boY64_1(.din(n3343), .dout(n3340));
    jdff dff_A_tttNuUrm6_1(.din(G8gat), .dout(n3343));
    jdff dff_A_Bn1RDwuN2_0(.din(n3349), .dout(n3346));
    jdff dff_A_0hA8ov3Z6_0(.din(n3352), .dout(n3349));
    jdff dff_A_4UeZc7LN8_0(.din(n3355), .dout(n3352));
    jdff dff_A_1XKNu4IG7_0(.din(n3358), .dout(n3355));
    jdff dff_A_KphDdd8P5_0(.din(n3361), .dout(n3358));
    jdff dff_A_HOZpH2xk1_0(.din(n521), .dout(n3361));
    jdff dff_A_wj4A0kFJ0_0(.din(n3367), .dout(n3364));
    jdff dff_A_lTb9FXNb9_0(.din(n3370), .dout(n3367));
    jdff dff_A_yzggL9pr8_0(.din(n3373), .dout(n3370));
    jdff dff_A_zhixABwN9_0(.din(n3376), .dout(n3373));
    jdff dff_A_8r4FoLHq8_0(.din(n3379), .dout(n3376));
    jdff dff_A_HTtol3Ui3_0(.din(n3382), .dout(n3379));
    jdff dff_A_Fw3USXt87_0(.din(n3385), .dout(n3382));
    jdff dff_A_oYqhOt2F2_0(.din(n3388), .dout(n3385));
    jdff dff_A_H7KaN3Pn9_0(.din(n3391), .dout(n3388));
    jdff dff_A_G3oHU4zl8_0(.din(n3394), .dout(n3391));
    jdff dff_A_xGqxvpuB2_0(.din(n3397), .dout(n3394));
    jdff dff_A_YPeFjJbQ3_0(.din(n3400), .dout(n3397));
    jdff dff_A_8NTOvryK9_0(.din(G86gat), .dout(n3400));
    jdff dff_A_Wj9TiAki9_1(.din(n3406), .dout(n3403));
    jdff dff_A_IxTDQcvy2_1(.din(n3409), .dout(n3406));
    jdff dff_A_0R3kRCOl1_1(.din(n3412), .dout(n3409));
    jdff dff_A_h5QL0kCJ5_1(.din(n3415), .dout(n3412));
    jdff dff_A_LYIfWeTe0_1(.din(n3418), .dout(n3415));
    jdff dff_A_ox9oGVPL0_1(.din(n3421), .dout(n3418));
    jdff dff_A_n0dbXPoS4_1(.din(n3424), .dout(n3421));
    jdff dff_A_4RTxeQTv8_1(.din(G86gat), .dout(n3424));
    jdff dff_A_CMuI8L6j7_1(.din(n3430), .dout(n3427));
    jdff dff_A_G9lrbznW0_1(.din(n330), .dout(n3430));
    jdff dff_A_KeFNm4pW6_1(.din(n3436), .dout(n3433));
    jdff dff_A_kC62ZcDW3_1(.din(n3439), .dout(n3436));
    jdff dff_A_jcY5vvGb8_1(.din(n3442), .dout(n3439));
    jdff dff_A_wRopOt5L7_1(.din(n3445), .dout(n3442));
    jdff dff_A_22tN93cK1_1(.din(n3448), .dout(n3445));
    jdff dff_A_us47lpq66_1(.din(n326), .dout(n3448));
    jdff dff_A_AC2CS2hU4_0(.din(n3454), .dout(n3451));
    jdff dff_A_shvZ5KCl4_0(.din(n3457), .dout(n3454));
    jdff dff_A_yPTK2SJA6_0(.din(n3460), .dout(n3457));
    jdff dff_A_BUk5ewy63_0(.din(n3463), .dout(n3460));
    jdff dff_A_i5tkwe6P9_0(.din(n3485), .dout(n3463));
    jdff dff_B_iEHWkATf7_2(.din(n318), .dout(n3467));
    jdff dff_B_eWavxSBs5_2(.din(n3467), .dout(n3470));
    jdff dff_B_GVnRsVxf0_2(.din(n3470), .dout(n3473));
    jdff dff_B_flLocZ0f0_2(.din(n3473), .dout(n3476));
    jdff dff_B_8H0gQXti6_2(.din(n3476), .dout(n3479));
    jdff dff_B_4MgC1ltu4_2(.din(n3479), .dout(n3482));
    jdff dff_B_A00qhiij1_2(.din(n3482), .dout(n3485));
    jdff dff_A_lolXuHU57_0(.din(n3490), .dout(n3487));
    jdff dff_A_druw62o49_0(.din(n3493), .dout(n3490));
    jdff dff_A_EWhHvAiG8_0(.din(n3496), .dout(n3493));
    jdff dff_A_Vjp4mi7i3_0(.din(n3499), .dout(n3496));
    jdff dff_A_uHBZwbJl4_0(.din(n3502), .dout(n3499));
    jdff dff_A_7h7Fu2Q37_0(.din(n3505), .dout(n3502));
    jdff dff_A_aBwOw3bx5_0(.din(n3508), .dout(n3505));
    jdff dff_A_L8UYUXoS7_0(.din(n3511), .dout(n3508));
    jdff dff_A_wOe423ER8_0(.din(n3514), .dout(n3511));
    jdff dff_A_VvECfKTc5_0(.din(n3517), .dout(n3514));
    jdff dff_A_Ca2DWTUk9_0(.din(n3520), .dout(n3517));
    jdff dff_A_WYBF2niX3_0(.din(n3523), .dout(n3520));
    jdff dff_A_Eb5WXesu6_0(.din(G60gat), .dout(n3523));
    jdff dff_B_NkP5lfii7_1(.din(n459), .dout(n3527));
    jdff dff_B_rpyFMvjf6_0(.din(n502), .dout(n3530));
    jdff dff_A_AV111u4x0_0(.din(n3535), .dout(n3532));
    jdff dff_A_wo8KVVH63_0(.din(n3538), .dout(n3535));
    jdff dff_A_ccHW2PQS0_0(.din(n3541), .dout(n3538));
    jdff dff_A_Xhx1JmBs3_0(.din(n3544), .dout(n3541));
    jdff dff_A_XsWQRDXO9_0(.din(n3547), .dout(n3544));
    jdff dff_A_4GiB9DAe3_0(.din(n498), .dout(n3547));
    jdff dff_B_ceKxluQL1_1(.din(n490), .dout(n3551));
    jdff dff_B_ixQvM5mF6_1(.din(n3551), .dout(n3554));
    jdff dff_B_rwvNWt2F9_1(.din(n3554), .dout(n3557));
    jdff dff_B_DThuhYie8_1(.din(n3557), .dout(n3560));
    jdff dff_B_rOFVomLb6_1(.din(n3560), .dout(n3563));
    jdff dff_B_KXeC1Orn6_1(.din(n3563), .dout(n3566));
    jdff dff_A_k3fKdYD15_0(.din(n3571), .dout(n3568));
    jdff dff_A_whBlaFGt4_0(.din(n3574), .dout(n3571));
    jdff dff_A_CuHV83vG7_0(.din(n3577), .dout(n3574));
    jdff dff_A_HSg7n5MY5_0(.din(n3580), .dout(n3577));
    jdff dff_A_cIuwW6t58_0(.din(n3583), .dout(n3580));
    jdff dff_A_D1ma7eyi6_0(.din(n3586), .dout(n3583));
    jdff dff_A_EdJiK31x6_0(.din(n3589), .dout(n3586));
    jdff dff_A_r3BlC9AS4_0(.din(n3592), .dout(n3589));
    jdff dff_A_Dsjj1ZWE9_0(.din(n3595), .dout(n3592));
    jdff dff_A_yUVK0bzL0_0(.din(n3598), .dout(n3595));
    jdff dff_A_bUhEWbP29_0(.din(n3601), .dout(n3598));
    jdff dff_A_07xr8NJQ7_0(.din(n3604), .dout(n3601));
    jdff dff_A_IGg9SyEP8_0(.din(G112gat), .dout(n3604));
    jdff dff_A_A4cTJAJG0_1(.din(n3610), .dout(n3607));
    jdff dff_A_VelxpJ7w3_1(.din(n3613), .dout(n3610));
    jdff dff_A_pbbzKgfQ3_1(.din(n3616), .dout(n3613));
    jdff dff_A_CrRJtig80_1(.din(n3619), .dout(n3616));
    jdff dff_A_16ISkeaI6_1(.din(n3622), .dout(n3619));
    jdff dff_A_9HJ1m68B0_1(.din(n3625), .dout(n3622));
    jdff dff_A_MRcXXCTX4_1(.din(n3628), .dout(n3625));
    jdff dff_A_Go6c1lDV5_1(.din(G112gat), .dout(n3628));
    jdff dff_A_8zIyKzcm6_0(.din(n3634), .dout(n3631));
    jdff dff_A_BXapyMDz5_0(.din(n3637), .dout(n3634));
    jdff dff_A_FBcAiRaI0_0(.din(n3640), .dout(n3637));
    jdff dff_A_jyNHHBvE5_0(.din(n3643), .dout(n3640));
    jdff dff_A_t01SNbxc5_0(.din(n3646), .dout(n3643));
    jdff dff_A_LLFs3lMj2_0(.din(n479), .dout(n3646));
    jdff dff_A_O0hk1lCZ9_0(.din(n3652), .dout(n3649));
    jdff dff_A_iy7XwnFi0_0(.din(n3655), .dout(n3652));
    jdff dff_A_9ClCkjFc1_0(.din(n3658), .dout(n3655));
    jdff dff_A_nDCd2ZVJ3_0(.din(n3661), .dout(n3658));
    jdff dff_A_PV5SEcjm8_0(.din(n3664), .dout(n3661));
    jdff dff_A_TfER06w00_0(.din(n3667), .dout(n3664));
    jdff dff_A_azgze0TS8_0(.din(n3670), .dout(n3667));
    jdff dff_A_4T1XvxtM9_0(.din(n3673), .dout(n3670));
    jdff dff_A_syqbI9W44_0(.din(n3676), .dout(n3673));
    jdff dff_A_NlPQNhwO8_0(.din(n3679), .dout(n3676));
    jdff dff_A_Cd7ZuZQ00_0(.din(n3682), .dout(n3679));
    jdff dff_A_ZMqb7ndf1_0(.din(n3685), .dout(n3682));
    jdff dff_A_qZdLlFXE3_0(.din(G34gat), .dout(n3685));
    jdff dff_A_6QRAG9CT9_1(.din(n3691), .dout(n3688));
    jdff dff_A_AcLiwcxi2_1(.din(n3694), .dout(n3691));
    jdff dff_A_qcwqUm645_1(.din(n3697), .dout(n3694));
    jdff dff_A_dYv6qkAD3_1(.din(n3700), .dout(n3697));
    jdff dff_A_dVLWKPsM2_1(.din(n3703), .dout(n3700));
    jdff dff_A_aGjZh8xo6_1(.din(n3706), .dout(n3703));
    jdff dff_A_uxhi2cct6_1(.din(n3709), .dout(n3706));
    jdff dff_A_z7fBMfWI3_1(.din(G34gat), .dout(n3709));
    jdff dff_A_2oNqJcOO7_0(.din(n3715), .dout(n3712));
    jdff dff_A_HRjeNp6v5_0(.din(n3718), .dout(n3715));
    jdff dff_A_aQ800rtG2_0(.din(n3721), .dout(n3718));
    jdff dff_A_2zq3WU0W6_0(.din(n3724), .dout(n3721));
    jdff dff_A_uV1tepnh5_0(.din(n3727), .dout(n3724));
    jdff dff_A_sKncualL7_0(.din(n467), .dout(n3727));
    jdff dff_A_5RRJF1ak2_1(.din(n3733), .dout(n3730));
    jdff dff_A_L1yUcqb50_1(.din(n3736), .dout(n3733));
    jdff dff_A_dkLUS4L14_1(.din(n3739), .dout(n3736));
    jdff dff_A_2m4pnNzZ3_1(.din(n3742), .dout(n3739));
    jdff dff_A_euCG29MY4_1(.din(n3745), .dout(n3742));
    jdff dff_A_GzJpBzPy9_1(.din(n399), .dout(n3745));
    jdff dff_A_TQUWBhtX2_0(.din(n3751), .dout(n3748));
    jdff dff_A_vJIq0LWk4_0(.din(n3754), .dout(n3751));
    jdff dff_A_NYzJIYwp2_0(.din(n3757), .dout(n3754));
    jdff dff_A_duF1Fab66_0(.din(n3760), .dout(n3757));
    jdff dff_A_HqieGEOn9_0(.din(n3763), .dout(n3760));
    jdff dff_A_STDLK6Qv8_0(.din(n3766), .dout(n3763));
    jdff dff_A_nZgFW8Dk0_0(.din(n3769), .dout(n3766));
    jdff dff_A_EV2WFCl09_0(.din(G99gat), .dout(n3769));
    jdff dff_A_MvLqRxip3_1(.din(n3775), .dout(n3772));
    jdff dff_A_wLWdPZcw9_1(.din(n3778), .dout(n3775));
    jdff dff_A_bLQHGVVf3_1(.din(n3781), .dout(n3778));
    jdff dff_A_VFNv39zM4_1(.din(n3784), .dout(n3781));
    jdff dff_A_bvzu4eKc1_1(.din(n3787), .dout(n3784));
    jdff dff_A_O7QdYVcU6_1(.din(n3790), .dout(n3787));
    jdff dff_A_NazXc7KQ6_1(.din(n3793), .dout(n3790));
    jdff dff_A_7yy3x1e71_1(.din(n3796), .dout(n3793));
    jdff dff_A_xPBJ9FAM0_1(.din(n3799), .dout(n3796));
    jdff dff_A_fQLewJoZ8_1(.din(n3802), .dout(n3799));
    jdff dff_A_9vng2tpv8_1(.din(n3805), .dout(n3802));
    jdff dff_A_chPBt41z6_1(.din(n3808), .dout(n3805));
    jdff dff_A_xwKVzm7V8_1(.din(G99gat), .dout(n3808));
    jdff dff_A_BRBQYKct3_0(.din(n3814), .dout(n3811));
    jdff dff_A_7nwawlw80_0(.din(n3817), .dout(n3814));
    jdff dff_A_IOns0ZG35_0(.din(n3820), .dout(n3817));
    jdff dff_A_0UIFhdOv2_0(.din(n3823), .dout(n3820));
    jdff dff_A_DZmf4tuv4_0(.din(n3826), .dout(n3823));
    jdff dff_A_YjxOWqGe8_0(.din(n447), .dout(n3826));
    jdff dff_B_YwTz4Rdk3_1(.din(n63), .dout(n3830));
    jdff dff_B_13jNcIH78_1(.din(n110), .dout(n3833));
    jdff dff_A_JInPuuqa8_0(.din(n3838), .dout(n3835));
    jdff dff_A_G1Aw1gSS7_0(.din(n3841), .dout(n3838));
    jdff dff_A_aNspGlsp1_0(.din(n3844), .dout(n3841));
    jdff dff_A_GDQYNaQN9_0(.din(n3847), .dout(n3844));
    jdff dff_A_kSn583jH5_0(.din(n120), .dout(n3847));
    jdff dff_A_TBubJOYM9_0(.din(n3853), .dout(n3850));
    jdff dff_A_8WMfvOJY9_0(.din(n3856), .dout(n3853));
    jdff dff_A_B6ddvVpF3_0(.din(n3859), .dout(n3856));
    jdff dff_A_IaUakkkr1_0(.din(n3862), .dout(n3859));
    jdff dff_A_fk6MrzLy9_0(.din(n113), .dout(n3862));
    jdff dff_A_UMoQmOdK2_0(.din(n3868), .dout(n3865));
    jdff dff_A_qqnjVmhM7_0(.din(n3871), .dout(n3868));
    jdff dff_A_hrgFTxrx9_0(.din(n3874), .dout(n3871));
    jdff dff_A_7AlZQU0f4_0(.din(n3877), .dout(n3874));
    jdff dff_A_9mFFV7fQ3_0(.din(n106), .dout(n3877));
    jdff dff_A_XFRjWb0e7_0(.din(n3883), .dout(n3880));
    jdff dff_A_AB5AJAx93_0(.din(n3886), .dout(n3883));
    jdff dff_A_7sx2afBE9_0(.din(n3889), .dout(n3886));
    jdff dff_A_rlN0UfkF4_0(.din(n95), .dout(n3889));
    jdff dff_A_ZeyIuTAQ0_0(.din(n3895), .dout(n3892));
    jdff dff_A_XfAAkZ0G4_0(.din(n3898), .dout(n3895));
    jdff dff_A_s1kCKJxT9_0(.din(n3901), .dout(n3898));
    jdff dff_A_JwZoJf724_0(.din(n3904), .dout(n3901));
    jdff dff_A_2sB8qnBj9_0(.din(n84), .dout(n3904));
    jdff dff_A_dmo9lwF68_0(.din(n3910), .dout(n3907));
    jdff dff_A_cN0njtaj5_0(.din(n3913), .dout(n3910));
    jdff dff_A_uwlUsmnk9_0(.din(n3916), .dout(n3913));
    jdff dff_A_CNqPklHs0_0(.din(n3919), .dout(n3916));
    jdff dff_A_EODEH6fW7_0(.din(n73), .dout(n3919));
    jdff dff_A_GjiScDiW3_0(.din(n3925), .dout(n3922));
    jdff dff_A_R73CpPBc0_0(.din(n3928), .dout(n3925));
    jdff dff_A_nhp2kmJQ0_0(.din(n59), .dout(n3928));
    jdff dff_A_X3q7bKiM4_0(.din(n3934), .dout(n3931));
    jdff dff_A_RNTOFx799_0(.din(n3937), .dout(n3934));
    jdff dff_A_SN7SJ5w29_0(.din(n3940), .dout(n3937));
    jdff dff_A_Y8ekKrsm4_0(.din(n3943), .dout(n3940));
    jdff dff_A_IqGY3AHw1_0(.din(n3946), .dout(n3943));
    jdff dff_A_bSHxnqms8_0(.din(n3949), .dout(n3946));
    jdff dff_A_anc3jKno6_0(.din(n3952), .dout(n3949));
    jdff dff_A_AOrQJtKy9_0(.din(n3955), .dout(n3952));
    jdff dff_A_YHIgEvW72_0(.din(n3958), .dout(n3955));
    jdff dff_A_M8ITuz5Y3_0(.din(n3961), .dout(n3958));
    jdff dff_A_hXIi3Tfy1_0(.din(n3964), .dout(n3961));
    jdff dff_A_ReeXbjtY2_0(.din(n3967), .dout(n3964));
    jdff dff_A_9ygUFtzK9_0(.din(G21gat), .dout(n3967));
    jdff dff_A_cGZvoynY1_1(.din(n3973), .dout(n3970));
    jdff dff_A_TPD2k8Xz9_1(.din(n3976), .dout(n3973));
    jdff dff_A_TqNdzYTj2_1(.din(n3979), .dout(n3976));
    jdff dff_A_ETYGaLcs1_1(.din(n3982), .dout(n3979));
    jdff dff_A_kkX8SL0T2_1(.din(n3985), .dout(n3982));
    jdff dff_A_1J93v6sV9_1(.din(n3988), .dout(n3985));
    jdff dff_A_uMKEEnY32_1(.din(n3991), .dout(n3988));
    jdff dff_A_2UsyUsik1_1(.din(G21gat), .dout(n3991));
    jdff dff_A_XHwaf2sQ1_0(.din(n3997), .dout(n3994));
    jdff dff_A_9NlhitPg0_0(.din(n4000), .dout(n3997));
    jdff dff_A_omjH5Oei0_0(.din(n4003), .dout(n4000));
    jdff dff_A_nhH959ff2_0(.din(n4006), .dout(n4003));
    jdff dff_A_xQEWaPFd4_0(.din(n4028), .dout(n4006));
    jdff dff_B_ixIUlemi6_2(.din(n261), .dout(n4010));
    jdff dff_B_oN58kuea0_2(.din(n4010), .dout(n4013));
    jdff dff_B_Q9b2boXO0_2(.din(n4013), .dout(n4016));
    jdff dff_B_vHmKgquF2_2(.din(n4016), .dout(n4019));
    jdff dff_B_t6OXCiwM1_2(.din(n4019), .dout(n4022));
    jdff dff_B_yn1gTL1Z5_2(.din(n4022), .dout(n4025));
    jdff dff_B_IF04gzgP6_2(.din(n4025), .dout(n4028));
    jdff dff_A_bU10WHIn3_0(.din(n4033), .dout(n4030));
    jdff dff_A_hvrbYllE2_0(.din(n4036), .dout(n4033));
    jdff dff_A_TxrgJKPe2_0(.din(n4039), .dout(n4036));
    jdff dff_A_3UCTd4K72_0(.din(n4042), .dout(n4039));
    jdff dff_A_QMSVHAYt5_0(.din(n4045), .dout(n4042));
    jdff dff_A_hyeI8XLQ6_0(.din(n4048), .dout(n4045));
    jdff dff_A_Cz0JYlKT3_0(.din(n4051), .dout(n4048));
    jdff dff_A_h8TvgjHo5_0(.din(n4054), .dout(n4051));
    jdff dff_A_GwkEOQSb7_0(.din(n4057), .dout(n4054));
    jdff dff_A_HivPc0ry6_0(.din(n4060), .dout(n4057));
    jdff dff_A_NSJpxvh96_0(.din(n4063), .dout(n4060));
    jdff dff_A_PjSU1GIe5_0(.din(n4066), .dout(n4063));
    jdff dff_A_YZreO8RO2_0(.din(G73gat), .dout(n4066));
    jdff dff_A_HUmFkQhw3_1(.din(n4072), .dout(n4069));
    jdff dff_A_EKVT5ugf1_1(.din(n4075), .dout(n4072));
    jdff dff_A_AZ5gkIHl5_1(.din(n4078), .dout(n4075));
    jdff dff_A_mj4enfqA6_1(.din(n4081), .dout(n4078));
    jdff dff_A_b3uE29Xi6_1(.din(n4084), .dout(n4081));
    jdff dff_A_SfkfkjLP5_1(.din(n4087), .dout(n4084));
    jdff dff_A_ilKvU5Xf7_1(.din(n4090), .dout(n4087));
    jdff dff_A_EE1vAm416_1(.din(G73gat), .dout(n4090));
    jdff dff_A_U9Sinh8X8_0(.din(n4096), .dout(n4093));
    jdff dff_A_1CKWLqAN1_0(.din(n4099), .dout(n4096));
    jdff dff_A_1jdCjZXD7_0(.din(n4102), .dout(n4099));
    jdff dff_A_ScTkoQ8O2_0(.din(n4105), .dout(n4102));
    jdff dff_A_4sJ3XD5G4_0(.din(n4108), .dout(n4105));
    jdff dff_A_zUsGRMpU8_0(.din(n269), .dout(n4108));
    jdff dff_B_iVWKt9F30_1(.din(n150), .dout(n4112));
    jdff dff_B_7OeTX8tP1_1(.din(n197), .dout(n4115));
    jdff dff_A_cLYJzDLR9_0(.din(n4120), .dout(n4117));
    jdff dff_A_9d8Zy8bX8_0(.din(n4123), .dout(n4120));
    jdff dff_A_I8zY70O09_0(.din(n4126), .dout(n4123));
    jdff dff_A_nKaof8P33_0(.din(n4129), .dout(n4126));
    jdff dff_A_AsYHRkx51_0(.din(n4132), .dout(n4129));
    jdff dff_A_kwJpDK9d3_0(.din(n207), .dout(n4132));
    jdff dff_A_pJCoHLR02_0(.din(n4138), .dout(n4135));
    jdff dff_A_SeAMmSL87_0(.din(n4141), .dout(n4138));
    jdff dff_A_qakHzVMB1_0(.din(n4144), .dout(n4141));
    jdff dff_A_NZCBwXPu8_0(.din(n4147), .dout(n4144));
    jdff dff_A_8Ff8nEbI3_0(.din(n4150), .dout(n4147));
    jdff dff_A_6gIMxOOk2_0(.din(n4153), .dout(n4150));
    jdff dff_A_NE6oXFhM3_0(.din(G82gat), .dout(n4153));
    jdff dff_A_jCLSgv0p3_2(.din(G82gat), .dout(n4156));
    jdff dff_A_pRmSFdzO9_0(.din(n4162), .dout(n4159));
    jdff dff_A_tW2aJNWD6_0(.din(n4165), .dout(n4162));
    jdff dff_A_eTIT3P1E9_0(.din(n4168), .dout(n4165));
    jdff dff_A_lbMIEfNe9_0(.din(n4171), .dout(n4168));
    jdff dff_A_iOnzaU6I2_0(.din(n4174), .dout(n4171));
    jdff dff_A_9dUrKNKd3_0(.din(G76gat), .dout(n4174));
    jdff dff_A_0ivgQ7UW7_1(.din(G76gat), .dout(n4177));
    jdff dff_A_sQG3aNIQ2_0(.din(n4183), .dout(n4180));
    jdff dff_A_NSLkkRcy3_0(.din(n4186), .dout(n4183));
    jdff dff_A_NZvhiyj07_0(.din(n4189), .dout(n4186));
    jdff dff_A_TtnypJFA6_0(.din(n4192), .dout(n4189));
    jdff dff_A_JuVeqah71_0(.din(n4195), .dout(n4192));
    jdff dff_A_VfX4Xf9w3_0(.din(n200), .dout(n4195));
    jdff dff_A_9RG3yveU9_0(.din(n4201), .dout(n4198));
    jdff dff_A_27ER9Jzv1_0(.din(n4204), .dout(n4201));
    jdff dff_A_tSk2aKxK9_0(.din(n4207), .dout(n4204));
    jdff dff_A_R0n8zemA2_0(.din(n4210), .dout(n4207));
    jdff dff_A_wyeJougk1_0(.din(n4213), .dout(n4210));
    jdff dff_A_rq5gl4iL9_0(.din(n4216), .dout(n4213));
    jdff dff_A_1s5F0kqf1_0(.din(G95gat), .dout(n4216));
    jdff dff_A_m3tq5pOZ7_2(.din(G95gat), .dout(n4219));
    jdff dff_A_bc99Wd5Z3_0(.din(n4225), .dout(n4222));
    jdff dff_A_vtgvAEaQ7_0(.din(n4228), .dout(n4225));
    jdff dff_A_jei1LsGN8_0(.din(n4231), .dout(n4228));
    jdff dff_A_sOO6HaqA6_0(.din(n4234), .dout(n4231));
    jdff dff_A_d2JnQgsp2_0(.din(n4237), .dout(n4234));
    jdff dff_A_lKn6yJlJ6_0(.din(G89gat), .dout(n4237));
    jdff dff_A_TRRJesDS2_1(.din(G89gat), .dout(n4240));
    jdff dff_A_xVmFd9Dm5_0(.din(n4246), .dout(n4243));
    jdff dff_A_uMGYBVYl1_0(.din(n4249), .dout(n4246));
    jdff dff_A_EiSnpKIJ6_0(.din(n4252), .dout(n4249));
    jdff dff_A_T7qDgt7E6_0(.din(n4255), .dout(n4252));
    jdff dff_A_dOTcBzwc9_0(.din(n4258), .dout(n4255));
    jdff dff_A_gGNBgYqU5_0(.din(n193), .dout(n4258));
    jdff dff_A_pcgnEsJ98_0(.din(n4264), .dout(n4261));
    jdff dff_A_GmnGWvfI8_0(.din(n4267), .dout(n4264));
    jdff dff_A_VHqVsIXk3_0(.din(n4270), .dout(n4267));
    jdff dff_A_2D6P5aMx2_0(.din(n4273), .dout(n4270));
    jdff dff_A_WiWzKvF72_0(.din(n4276), .dout(n4273));
    jdff dff_A_S1nC82Tx3_0(.din(n4279), .dout(n4276));
    jdff dff_A_u2Wkcub51_0(.din(G4gat), .dout(n4279));
    jdff dff_A_CPVaA3YE2_2(.din(G4gat), .dout(n4282));
    jdff dff_A_hl3QBdk34_0(.din(n4288), .dout(n4285));
    jdff dff_A_M4NHu0WP6_0(.din(n4291), .dout(n4288));
    jdff dff_A_2GBha37m9_0(.din(n4294), .dout(n4291));
    jdff dff_A_dTgi6XPn2_0(.din(n4297), .dout(n4294));
    jdff dff_A_7fGXVDn78_0(.din(n4300), .dout(n4297));
    jdff dff_A_9feHHqEP9_0(.din(G1gat), .dout(n4300));
    jdff dff_A_ZUmlp4ih2_1(.din(G1gat), .dout(n4303));
    jdff dff_A_893RPwEf4_0(.din(n4309), .dout(n4306));
    jdff dff_A_luoqwI3p0_0(.din(n4312), .dout(n4309));
    jdff dff_A_dZEkaBhF4_0(.din(n4315), .dout(n4312));
    jdff dff_A_QWq5YH7x7_0(.din(n182), .dout(n4315));
    jdff dff_A_s3FmS4px5_0(.din(n4321), .dout(n4318));
    jdff dff_A_2z1I5Puz3_0(.din(n4324), .dout(n4321));
    jdff dff_A_ULD4DwGY1_0(.din(n4327), .dout(n4324));
    jdff dff_A_VeGUxuiq8_0(.din(n4330), .dout(n4327));
    jdff dff_A_ZKU1lP1t1_0(.din(n4333), .dout(n4330));
    jdff dff_A_NMfp3Yml3_0(.din(n4336), .dout(n4333));
    jdff dff_A_5iMHirOA5_0(.din(n4339), .dout(n4336));
    jdff dff_A_2jtw5R4j9_0(.din(n4342), .dout(n4339));
    jdff dff_A_EcgTezgs3_0(.din(n4345), .dout(n4342));
    jdff dff_A_wfQ7uCxp3_0(.din(n4348), .dout(n4345));
    jdff dff_A_GiJdxXtb8_0(.din(n4351), .dout(n4348));
    jdff dff_A_bgcdtyLP4_0(.din(n4354), .dout(n4351));
    jdff dff_A_0bQ4fxyL7_0(.din(n4357), .dout(n4354));
    jdff dff_A_eSJpdP357_0(.din(n4360), .dout(n4357));
    jdff dff_A_C69Ak8SM2_0(.din(n4363), .dout(n4360));
    jdff dff_A_m4p2c9nk5_0(.din(n4366), .dout(n4363));
    jdff dff_A_A1f7VNc53_0(.din(n4369), .dout(n4366));
    jdff dff_A_xY1SuJ7Y7_0(.din(n4372), .dout(n4369));
    jdff dff_A_INVL3gxL2_0(.din(n4375), .dout(n4372));
    jdff dff_A_mziMIdWz5_0(.din(n4378), .dout(n4375));
    jdff dff_A_KULj1DkY4_0(.din(n178), .dout(n4378));
    jdff dff_A_dZOlZMLW4_1(.din(G56gat), .dout(n4381));
    jdff dff_A_LVGuxcLB1_1(.din(n4387), .dout(n4384));
    jdff dff_A_wmTR8ict7_1(.din(n4390), .dout(n4387));
    jdff dff_A_yFShnhJM9_1(.din(n4393), .dout(n4390));
    jdff dff_A_ZMA7FEMY9_1(.din(n4396), .dout(n4393));
    jdff dff_A_qhPKt9yi6_1(.din(n4399), .dout(n4396));
    jdff dff_A_ySmVm7jB4_1(.din(n4402), .dout(n4399));
    jdff dff_A_oiBtZd8U0_1(.din(n4405), .dout(n4402));
    jdff dff_A_FBpKnxet5_1(.din(n4408), .dout(n4405));
    jdff dff_A_fYIfsCf14_1(.din(n4411), .dout(n4408));
    jdff dff_A_xozF5Ach0_1(.din(n4414), .dout(n4411));
    jdff dff_A_pdTn0NBz5_1(.din(n4417), .dout(n4414));
    jdff dff_A_UrBp0ROh1_1(.din(n4420), .dout(n4417));
    jdff dff_A_SbqqBJrZ8_1(.din(n4423), .dout(n4420));
    jdff dff_A_PcM4HkA08_1(.din(n4426), .dout(n4423));
    jdff dff_A_Ht3awnJL8_1(.din(n4429), .dout(n4426));
    jdff dff_A_2ixDfRJv6_1(.din(n4432), .dout(n4429));
    jdff dff_A_j3CELniN6_1(.din(n4435), .dout(n4432));
    jdff dff_A_p3oH2QIB6_1(.din(n4438), .dout(n4435));
    jdff dff_A_c91kfoCy9_1(.din(n4441), .dout(n4438));
    jdff dff_A_x2trJ02B9_1(.din(n4444), .dout(n4441));
    jdff dff_A_KLpJZTcl2_1(.din(n4447), .dout(n4444));
    jdff dff_A_t52nroUK4_1(.din(G56gat), .dout(n4447));
    jdff dff_A_68hQuQow0_2(.din(n4453), .dout(n4450));
    jdff dff_A_UAyRo1Zw5_2(.din(n4456), .dout(n4453));
    jdff dff_A_cZX06fTd3_2(.din(n4459), .dout(n4456));
    jdff dff_A_rhNdrFvP2_2(.din(n4462), .dout(n4459));
    jdff dff_A_84alNLuP1_2(.din(n4465), .dout(n4462));
    jdff dff_A_3RBbZaOv7_2(.din(n4468), .dout(n4465));
    jdff dff_A_HM7Xt9M00_2(.din(G56gat), .dout(n4468));
    jdff dff_A_sns6gJAF5_0(.din(G50gat), .dout(n4471));
    jdff dff_A_ygNnZWiE9_0(.din(n4477), .dout(n4474));
    jdff dff_A_UYxhPOTK9_0(.din(n4480), .dout(n4477));
    jdff dff_A_OstBHuum1_0(.din(n4483), .dout(n4480));
    jdff dff_A_LXonWnii7_0(.din(n4486), .dout(n4483));
    jdff dff_A_ReADckMX0_0(.din(n4489), .dout(n4486));
    jdff dff_A_4tjV6s9y4_0(.din(n171), .dout(n4489));
    jdff dff_A_44Q1Hx1w5_0(.din(n4495), .dout(n4492));
    jdff dff_A_ErKFxt4K2_0(.din(n4498), .dout(n4495));
    jdff dff_A_l0mWy9y61_0(.din(n4501), .dout(n4498));
    jdff dff_A_QmPZJawy2_0(.din(n4504), .dout(n4501));
    jdff dff_A_mVgvovWA6_0(.din(n4507), .dout(n4504));
    jdff dff_A_s7Pv9KOO4_0(.din(n4510), .dout(n4507));
    jdff dff_A_TclB1t9Z4_0(.din(G30gat), .dout(n4510));
    jdff dff_A_GkEWWy088_2(.din(G30gat), .dout(n4513));
    jdff dff_A_VhMnQ70e8_0(.din(n4519), .dout(n4516));
    jdff dff_A_RbLgk9ah9_0(.din(n4522), .dout(n4519));
    jdff dff_A_NcyuVqO52_0(.din(n4525), .dout(n4522));
    jdff dff_A_FKAcYUAm7_0(.din(n4528), .dout(n4525));
    jdff dff_A_cLWxCmsI0_0(.din(n4531), .dout(n4528));
endmodule

