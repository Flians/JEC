// Benchmark "c7552" written by ABC on Wed May 27 22:06:16 2020

module gf_c7552 ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496,
    G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253,
    G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743,
    G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432,
    G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire n317, n318, n319, n320, n321, n322, n324, n325, n326, n327, n328,
    n329, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342,
    n343, n345, n347, n348, n349, n352, n353, n354, n355, n356, n357, n358,
    n359, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1078, n1079, n1080,
    n1082, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1102, n1103,
    n1105, n1106, n1107, n1108, n1109, n1110, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1347, n1348, n1349, n1351, n1352, n1353,
    n1354, n1356, n1357, n1359, n1360, n1361, n1363, n1364, n1365, n1366,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1377, n1378, n1379,
    n1380, n1381, n1384, n1385, n1387, n1388, n1389, n1390, n1394, n1395,
    n1396, n1399, n1400, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1413, n1414, n1416, n1417, n1419, n1421, n1423,
    n1424, n1426, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632;
  jnot g0000(.din(G15), .dout(G279));
  jor  g0001(.dina(G57), .dinb(G5), .dout(G402));
  jnot g0002(.din(G184), .dout(n317));
  jnot g0003(.din(G228), .dout(n318));
  jor  g0004(.dina(n318), .dinb(n317), .dout(n319));
  jnot g0005(.din(G150), .dout(n320));
  jnot g0006(.din(G240), .dout(n321));
  jor  g0007(.dina(n321), .dinb(n320), .dout(n322));
  jor  g0008(.dina(n322), .dinb(n319), .dout(G404));
  jnot g0009(.din(G210), .dout(n324));
  jnot g0010(.din(G218), .dout(n325));
  jor  g0011(.dina(n325), .dinb(n324), .dout(n326));
  jnot g0012(.din(G152), .dout(n327));
  jnot g0013(.din(G230), .dout(n328));
  jor  g0014(.dina(n328), .dinb(n327), .dout(n329));
  jor  g0015(.dina(n329), .dinb(n326), .dout(G406));
  jnot g0016(.din(G183), .dout(n331));
  jnot g0017(.din(G185), .dout(n332));
  jor  g0018(.dina(n332), .dinb(n331), .dout(n333));
  jnot g0019(.din(G182), .dout(n334));
  jnot g0020(.din(G186), .dout(n335));
  jor  g0021(.dina(n335), .dinb(n334), .dout(n336));
  jor  g0022(.dina(n336), .dinb(n333), .dout(G408));
  jnot g0023(.din(G172), .dout(n338));
  jnot g0024(.din(G188), .dout(n339));
  jor  g0025(.dina(n339), .dinb(n338), .dout(n340));
  jnot g0026(.din(G162), .dout(n341));
  jnot g0027(.din(G199), .dout(n342));
  jor  g0028(.dina(n342), .dinb(n341), .dout(n343));
  jor  g0029(.dina(n343), .dinb(n340), .dout(G410));
  jnot g0030(.din(G1197), .dout(n345));
  jor  g0031(.dina(n345), .dinb(G5), .dout(G284));
  jnot g0032(.din(G134), .dout(n347));
  jnot g0033(.din(G133), .dout(n348));
  jor  g0034(.dina(n348), .dinb(G5), .dout(n349));
  jor  g0035(.dina(n349), .dinb(n347), .dout(G292));
  jand g0036(.dina(G163), .dinb(G1), .dout(G278));
  jnot g0037(.din(G41), .dout(n352));
  jor  g0038(.dina(n352), .dinb(G18), .dout(n353));
  jor  g0039(.dina(n353), .dinb(G3701), .dout(n354));
  jnot g0040(.din(G18), .dout(n355));
  jand g0041(.dina(G3701), .dinb(n355), .dout(n356));
  jand g0042(.dina(n356), .dinb(n353), .dout(n357));
  jnot g0043(.din(n357), .dout(n358));
  jand g0044(.dina(n358), .dinb(n354), .dout(n359));
  jxor g0045(.dina(n359), .dinb(G4526), .dout(G373));
  jnot g0046(.din(G38), .dout(n361));
  jand g0047(.dina(G4528), .dinb(G1492), .dout(n362));
  jxor g0048(.dina(n362), .dinb(n361), .dout(n363));
  jand g0049(.dina(G4528), .dinb(G1496), .dout(n364));
  jor  g0050(.dina(n364), .dinb(n361), .dout(n365));
  jnot g0051(.din(G1496), .dout(n366));
  jnot g0052(.din(G4528), .dout(n367));
  jor  g0053(.dina(n367), .dinb(G38), .dout(n368));
  jor  g0054(.dina(n368), .dinb(n366), .dout(n369));
  jand g0055(.dina(n369), .dinb(n365), .dout(n370));
  jnot g0056(.din(G1486), .dout(n371));
  jand g0057(.dina(G12), .dinb(G9), .dout(n372));
  jnot g0058(.din(n372), .dout(n373));
  jor  g0059(.dina(G213), .dinb(n355), .dout(n374));
  jand g0060(.dina(n374), .dinb(n373), .dout(n375));
  jand g0061(.dina(n375), .dinb(n371), .dout(n376));
  jxor g0062(.dina(n375), .dinb(n371), .dout(n377));
  jor  g0063(.dina(G214), .dinb(n355), .dout(n378));
  jand g0064(.dina(n378), .dinb(n373), .dout(n379));
  jnot g0065(.din(n379), .dout(n380));
  jand g0066(.dina(n380), .dinb(G1480), .dout(n381));
  jnot g0067(.din(n381), .dout(n382));
  jnot g0068(.din(G1480), .dout(n383));
  jand g0069(.dina(n379), .dinb(n383), .dout(n384));
  jnot g0070(.din(G106), .dout(n385));
  jor  g0071(.dina(G215), .dinb(n355), .dout(n386));
  jand g0072(.dina(n386), .dinb(n373), .dout(n387));
  jxor g0073(.dina(n387), .dinb(n385), .dout(n388));
  jnot g0074(.din(G1462), .dout(n389));
  jor  g0075(.dina(G209), .dinb(n355), .dout(n390));
  jand g0076(.dina(n390), .dinb(n373), .dout(n391));
  jand g0077(.dina(n391), .dinb(n389), .dout(n392));
  jnot g0078(.din(G1469), .dout(n393));
  jor  g0079(.dina(G216), .dinb(n355), .dout(n394));
  jand g0080(.dina(n394), .dinb(n373), .dout(n395));
  jxor g0081(.dina(n395), .dinb(n393), .dout(n396));
  jand g0082(.dina(n396), .dinb(n392), .dout(n397));
  jand g0083(.dina(n397), .dinb(n388), .dout(n398));
  jnot g0084(.din(n398), .dout(n399));
  jand g0085(.dina(n387), .dinb(n385), .dout(n400));
  jnot g0086(.din(n400), .dout(n401));
  jnot g0087(.din(n387), .dout(n402));
  jand g0088(.dina(n402), .dinb(G106), .dout(n403));
  jand g0089(.dina(n395), .dinb(n393), .dout(n404));
  jnot g0090(.din(n404), .dout(n405));
  jor  g0091(.dina(n405), .dinb(n403), .dout(n406));
  jand g0092(.dina(n406), .dinb(n401), .dout(n407));
  jand g0093(.dina(n407), .dinb(n399), .dout(n408));
  jnot g0094(.din(n408), .dout(n409));
  jor  g0095(.dina(n409), .dinb(n384), .dout(n410));
  jand g0096(.dina(n410), .dinb(n382), .dout(n411));
  jand g0097(.dina(n411), .dinb(n377), .dout(n412));
  jor  g0098(.dina(n412), .dinb(n376), .dout(n413));
  jxor g0099(.dina(n391), .dinb(n389), .dout(n414));
  jand g0100(.dina(n414), .dinb(n396), .dout(n415));
  jxor g0101(.dina(n379), .dinb(n383), .dout(n416));
  jand g0102(.dina(n416), .dinb(n388), .dout(n417));
  jand g0103(.dina(n417), .dinb(n415), .dout(n418));
  jand g0104(.dina(n418), .dinb(n377), .dout(n419));
  jor  g0105(.dina(n419), .dinb(n413), .dout(n420));
  jnot g0106(.din(G2256), .dout(n421));
  jor  g0107(.dina(G153), .dinb(n355), .dout(n422));
  jand g0108(.dina(n422), .dinb(n373), .dout(n423));
  jand g0109(.dina(n423), .dinb(n421), .dout(n424));
  jxor g0110(.dina(n423), .dinb(n421), .dout(n425));
  jnot g0111(.din(G2253), .dout(n426));
  jor  g0112(.dina(G154), .dinb(n355), .dout(n427));
  jand g0113(.dina(n427), .dinb(n373), .dout(n428));
  jxor g0114(.dina(n428), .dinb(n426), .dout(n429));
  jnot g0115(.din(G2247), .dout(n430));
  jor  g0116(.dina(G155), .dinb(n355), .dout(n431));
  jand g0117(.dina(n431), .dinb(n373), .dout(n432));
  jxor g0118(.dina(n432), .dinb(n430), .dout(n433));
  jnot g0119(.din(G2239), .dout(n434));
  jor  g0120(.dina(G156), .dinb(n355), .dout(n435));
  jand g0121(.dina(n435), .dinb(n373), .dout(n436));
  jxor g0122(.dina(n436), .dinb(n434), .dout(n437));
  jand g0123(.dina(n437), .dinb(n433), .dout(n438));
  jand g0124(.dina(n438), .dinb(n429), .dout(n439));
  jnot g0125(.din(n428), .dout(n440));
  jand g0126(.dina(n440), .dinb(G2253), .dout(n441));
  jnot g0127(.din(n441), .dout(n442));
  jand g0128(.dina(n428), .dinb(n426), .dout(n443));
  jand g0129(.dina(n432), .dinb(n430), .dout(n444));
  jand g0130(.dina(n436), .dinb(n434), .dout(n445));
  jand g0131(.dina(n445), .dinb(n433), .dout(n446));
  jor  g0132(.dina(n446), .dinb(n444), .dout(n447));
  jor  g0133(.dina(n447), .dinb(n443), .dout(n448));
  jand g0134(.dina(n448), .dinb(n442), .dout(n449));
  jor  g0135(.dina(n449), .dinb(n439), .dout(n450));
  jnot g0136(.din(G2236), .dout(n451));
  jor  g0137(.dina(G157), .dinb(n355), .dout(n452));
  jand g0138(.dina(n452), .dinb(n373), .dout(n453));
  jand g0139(.dina(n453), .dinb(n451), .dout(n454));
  jor  g0140(.dina(n453), .dinb(n451), .dout(n455));
  jnot g0141(.din(G2230), .dout(n456));
  jand g0142(.dina(G135), .dinb(n355), .dout(n457));
  jand g0143(.dina(G158), .dinb(G18), .dout(n458));
  jor  g0144(.dina(n458), .dinb(n457), .dout(n459));
  jand g0145(.dina(n459), .dinb(n456), .dout(n460));
  jand g0146(.dina(n460), .dinb(n455), .dout(n461));
  jor  g0147(.dina(n461), .dinb(n454), .dout(n462));
  jxor g0148(.dina(n453), .dinb(n451), .dout(n463));
  jxor g0149(.dina(n459), .dinb(n456), .dout(n464));
  jand g0150(.dina(n464), .dinb(n463), .dout(n465));
  jnot g0151(.din(G2224), .dout(n466));
  jand g0152(.dina(G144), .dinb(n355), .dout(n467));
  jand g0153(.dina(G159), .dinb(G18), .dout(n468));
  jor  g0154(.dina(n468), .dinb(n467), .dout(n469));
  jxor g0155(.dina(n469), .dinb(n466), .dout(n470));
  jnot g0156(.din(G2218), .dout(n471));
  jand g0157(.dina(G138), .dinb(n355), .dout(n472));
  jand g0158(.dina(G160), .dinb(G18), .dout(n473));
  jor  g0159(.dina(n473), .dinb(n472), .dout(n474));
  jxor g0160(.dina(n474), .dinb(n471), .dout(n475));
  jnot g0161(.din(G2211), .dout(n476));
  jand g0162(.dina(G147), .dinb(n355), .dout(n477));
  jand g0163(.dina(G151), .dinb(G18), .dout(n478));
  jor  g0164(.dina(n478), .dinb(n477), .dout(n479));
  jxor g0165(.dina(n479), .dinb(n476), .dout(n480));
  jand g0166(.dina(n480), .dinb(n475), .dout(n481));
  jand g0167(.dina(n481), .dinb(n470), .dout(n482));
  jnot g0168(.din(n469), .dout(n483));
  jand g0169(.dina(n483), .dinb(G2224), .dout(n484));
  jnot g0170(.din(n474), .dout(n485));
  jand g0171(.dina(n485), .dinb(G2218), .dout(n486));
  jand g0172(.dina(n479), .dinb(n476), .dout(n487));
  jnot g0173(.din(n487), .dout(n488));
  jor  g0174(.dina(n488), .dinb(n486), .dout(n489));
  jand g0175(.dina(n469), .dinb(n466), .dout(n490));
  jand g0176(.dina(n474), .dinb(n471), .dout(n491));
  jor  g0177(.dina(n491), .dinb(n490), .dout(n492));
  jnot g0178(.din(n492), .dout(n493));
  jand g0179(.dina(n493), .dinb(n489), .dout(n494));
  jor  g0180(.dina(n494), .dinb(n484), .dout(n495));
  jnot g0181(.din(n495), .dout(n496));
  jor  g0182(.dina(n496), .dinb(n482), .dout(n497));
  jand g0183(.dina(n497), .dinb(n465), .dout(n498));
  jor  g0184(.dina(n498), .dinb(n462), .dout(n499));
  jand g0185(.dina(n496), .dinb(n465), .dout(n500));
  jnot g0186(.din(G4437), .dout(n501));
  jand g0187(.dina(G219), .dinb(G18), .dout(n502));
  jand g0188(.dina(G66), .dinb(n355), .dout(n503));
  jor  g0189(.dina(n503), .dinb(n502), .dout(n504));
  jand g0190(.dina(n504), .dinb(n501), .dout(n505));
  jnot g0191(.din(n504), .dout(n506));
  jand g0192(.dina(n506), .dinb(G4437), .dout(n507));
  jnot g0193(.din(n507), .dout(n508));
  jnot g0194(.din(G4432), .dout(n509));
  jand g0195(.dina(G220), .dinb(G18), .dout(n510));
  jand g0196(.dina(G50), .dinb(n355), .dout(n511));
  jor  g0197(.dina(n511), .dinb(n510), .dout(n512));
  jxor g0198(.dina(n512), .dinb(n509), .dout(n513));
  jnot g0199(.din(G4420), .dout(n514));
  jand g0200(.dina(G222), .dinb(G18), .dout(n515));
  jand g0201(.dina(G35), .dinb(n355), .dout(n516));
  jor  g0202(.dina(n516), .dinb(n515), .dout(n517));
  jand g0203(.dina(n517), .dinb(n514), .dout(n518));
  jnot g0204(.din(n518), .dout(n519));
  jnot g0205(.din(G4427), .dout(n520));
  jand g0206(.dina(G221), .dinb(G18), .dout(n521));
  jand g0207(.dina(G32), .dinb(n355), .dout(n522));
  jor  g0208(.dina(n522), .dinb(n521), .dout(n523));
  jxor g0209(.dina(n523), .dinb(n520), .dout(n524));
  jnot g0210(.din(n517), .dout(n525));
  jand g0211(.dina(n525), .dinb(G4420), .dout(n526));
  jnot g0212(.din(n526), .dout(n527));
  jnot g0213(.din(G4415), .dout(n528));
  jand g0214(.dina(G223), .dinb(G18), .dout(n529));
  jand g0215(.dina(G47), .dinb(n355), .dout(n530));
  jor  g0216(.dina(n530), .dinb(n529), .dout(n531));
  jand g0217(.dina(n531), .dinb(n528), .dout(n532));
  jnot g0218(.din(n531), .dout(n533));
  jand g0219(.dina(n533), .dinb(G4415), .dout(n534));
  jnot g0220(.din(n534), .dout(n535));
  jnot g0221(.din(G4410), .dout(n536));
  jand g0222(.dina(G224), .dinb(G18), .dout(n537));
  jand g0223(.dina(G121), .dinb(n355), .dout(n538));
  jor  g0224(.dina(n538), .dinb(n537), .dout(n539));
  jand g0225(.dina(n539), .dinb(n536), .dout(n540));
  jnot g0226(.din(n539), .dout(n541));
  jand g0227(.dina(n541), .dinb(G4410), .dout(n542));
  jnot g0228(.din(n542), .dout(n543));
  jnot g0229(.din(G4405), .dout(n544));
  jand g0230(.dina(G225), .dinb(G18), .dout(n545));
  jand g0231(.dina(G94), .dinb(n355), .dout(n546));
  jor  g0232(.dina(n546), .dinb(n545), .dout(n547));
  jand g0233(.dina(n547), .dinb(n544), .dout(n548));
  jnot g0234(.din(n547), .dout(n549));
  jand g0235(.dina(n549), .dinb(G4405), .dout(n550));
  jnot g0236(.din(n550), .dout(n551));
  jnot g0237(.din(G4400), .dout(n552));
  jand g0238(.dina(G226), .dinb(G18), .dout(n553));
  jand g0239(.dina(G97), .dinb(n355), .dout(n554));
  jor  g0240(.dina(n554), .dinb(n553), .dout(n555));
  jand g0241(.dina(n555), .dinb(n552), .dout(n556));
  jnot g0242(.din(n555), .dout(n557));
  jand g0243(.dina(n557), .dinb(G4400), .dout(n558));
  jnot g0244(.din(n558), .dout(n559));
  jnot g0245(.din(G4394), .dout(n560));
  jand g0246(.dina(G217), .dinb(G18), .dout(n561));
  jand g0247(.dina(G118), .dinb(n355), .dout(n562));
  jor  g0248(.dina(n562), .dinb(n561), .dout(n563));
  jand g0249(.dina(n563), .dinb(n560), .dout(n564));
  jand g0250(.dina(n564), .dinb(n559), .dout(n565));
  jor  g0251(.dina(n565), .dinb(n556), .dout(n566));
  jand g0252(.dina(n566), .dinb(n551), .dout(n567));
  jor  g0253(.dina(n567), .dinb(n548), .dout(n568));
  jand g0254(.dina(n568), .dinb(n543), .dout(n569));
  jor  g0255(.dina(n569), .dinb(n540), .dout(n570));
  jand g0256(.dina(n570), .dinb(n535), .dout(n571));
  jor  g0257(.dina(n571), .dinb(n532), .dout(n572));
  jxor g0258(.dina(n531), .dinb(n528), .dout(n573));
  jxor g0259(.dina(n555), .dinb(n552), .dout(n574));
  jxor g0260(.dina(n563), .dinb(n560), .dout(n575));
  jand g0261(.dina(n575), .dinb(n574), .dout(n576));
  jxor g0262(.dina(n539), .dinb(n536), .dout(n577));
  jxor g0263(.dina(n547), .dinb(n544), .dout(n578));
  jand g0264(.dina(n578), .dinb(n577), .dout(n579));
  jand g0265(.dina(n579), .dinb(n576), .dout(n580));
  jand g0266(.dina(n580), .dinb(n573), .dout(n581));
  jnot g0267(.din(G3749), .dout(n582));
  jand g0268(.dina(G231), .dinb(G18), .dout(n583));
  jand g0269(.dina(G100), .dinb(n355), .dout(n584));
  jor  g0270(.dina(n584), .dinb(n583), .dout(n585));
  jand g0271(.dina(n585), .dinb(n582), .dout(n586));
  jnot g0272(.din(n585), .dout(n587));
  jand g0273(.dina(n587), .dinb(G3749), .dout(n588));
  jnot g0274(.din(n588), .dout(n589));
  jnot g0275(.din(G3743), .dout(n590));
  jand g0276(.dina(G232), .dinb(G18), .dout(n591));
  jand g0277(.dina(G124), .dinb(n355), .dout(n592));
  jor  g0278(.dina(n592), .dinb(n591), .dout(n593));
  jxor g0279(.dina(n593), .dinb(n590), .dout(n594));
  jnot g0280(.din(G3737), .dout(n595));
  jand g0281(.dina(G233), .dinb(G18), .dout(n596));
  jand g0282(.dina(G127), .dinb(n355), .dout(n597));
  jor  g0283(.dina(n597), .dinb(n596), .dout(n598));
  jxor g0284(.dina(n598), .dinb(n595), .dout(n599));
  jnot g0285(.din(G3729), .dout(n600));
  jand g0286(.dina(G234), .dinb(G18), .dout(n601));
  jand g0287(.dina(G130), .dinb(n355), .dout(n602));
  jor  g0288(.dina(n602), .dinb(n601), .dout(n603));
  jxor g0289(.dina(n603), .dinb(n600), .dout(n604));
  jand g0290(.dina(n604), .dinb(n599), .dout(n605));
  jand g0291(.dina(n605), .dinb(n594), .dout(n606));
  jnot g0292(.din(n606), .dout(n607));
  jnot g0293(.din(n593), .dout(n608));
  jand g0294(.dina(n608), .dinb(G3743), .dout(n609));
  jand g0295(.dina(n593), .dinb(n590), .dout(n610));
  jnot g0296(.din(n610), .dout(n611));
  jand g0297(.dina(n598), .dinb(n595), .dout(n612));
  jand g0298(.dina(n603), .dinb(n600), .dout(n613));
  jand g0299(.dina(n613), .dinb(n599), .dout(n614));
  jor  g0300(.dina(n614), .dinb(n612), .dout(n615));
  jnot g0301(.din(n615), .dout(n616));
  jand g0302(.dina(n616), .dinb(n611), .dout(n617));
  jor  g0303(.dina(n617), .dinb(n609), .dout(n618));
  jand g0304(.dina(n618), .dinb(n607), .dout(n619));
  jnot g0305(.din(n619), .dout(n620));
  jnot g0306(.din(n618), .dout(n621));
  jnot g0307(.din(G3723), .dout(n622));
  jand g0308(.dina(G235), .dinb(G18), .dout(n623));
  jand g0309(.dina(G103), .dinb(n355), .dout(n624));
  jor  g0310(.dina(n624), .dinb(n623), .dout(n625));
  jxor g0311(.dina(n625), .dinb(n622), .dout(n626));
  jnot g0312(.din(G3717), .dout(n627));
  jand g0313(.dina(G236), .dinb(G18), .dout(n628));
  jand g0314(.dina(G23), .dinb(n355), .dout(n629));
  jor  g0315(.dina(n629), .dinb(n628), .dout(n630));
  jxor g0316(.dina(n630), .dinb(n627), .dout(n631));
  jnot g0317(.din(G3711), .dout(n632));
  jand g0318(.dina(G237), .dinb(G18), .dout(n633));
  jand g0319(.dina(G26), .dinb(n355), .dout(n634));
  jor  g0320(.dina(n634), .dinb(n633), .dout(n635));
  jxor g0321(.dina(n635), .dinb(n632), .dout(n636));
  jnot g0322(.din(G238), .dout(n637));
  jor  g0323(.dina(n637), .dinb(n355), .dout(n638));
  jnot g0324(.din(G29), .dout(n639));
  jor  g0325(.dina(n639), .dinb(G18), .dout(n640));
  jand g0326(.dina(n640), .dinb(n638), .dout(n641));
  jxor g0327(.dina(n641), .dinb(G3705), .dout(n642));
  jand g0328(.dina(n642), .dinb(n359), .dout(n643));
  jand g0329(.dina(n643), .dinb(n636), .dout(n644));
  jand g0330(.dina(n644), .dinb(n631), .dout(n645));
  jand g0331(.dina(n645), .dinb(n626), .dout(n646));
  jand g0332(.dina(n625), .dinb(n622), .dout(n647));
  jnot g0333(.din(n625), .dout(n648));
  jand g0334(.dina(n648), .dinb(G3723), .dout(n649));
  jnot g0335(.din(n649), .dout(n650));
  jnot g0336(.din(n630), .dout(n651));
  jand g0337(.dina(n651), .dinb(G3717), .dout(n652));
  jnot g0338(.din(n652), .dout(n653));
  jand g0339(.dina(n630), .dinb(n627), .dout(n654));
  jand g0340(.dina(n635), .dinb(n632), .dout(n655));
  jor  g0341(.dina(n635), .dinb(n632), .dout(n656));
  jnot g0342(.din(G3705), .dout(n657));
  jand g0343(.dina(G238), .dinb(G18), .dout(n658));
  jand g0344(.dina(G29), .dinb(n355), .dout(n659));
  jor  g0345(.dina(n659), .dinb(n658), .dout(n660));
  jor  g0346(.dina(n660), .dinb(n657), .dout(n661));
  jnot g0347(.din(G3701), .dout(n662));
  jand g0348(.dina(G41), .dinb(n355), .dout(n663));
  jand g0349(.dina(n663), .dinb(n662), .dout(n664));
  jand g0350(.dina(n660), .dinb(n657), .dout(n665));
  jor  g0351(.dina(n665), .dinb(n664), .dout(n666));
  jand g0352(.dina(n666), .dinb(n661), .dout(n667));
  jand g0353(.dina(n667), .dinb(n656), .dout(n668));
  jor  g0354(.dina(n668), .dinb(n655), .dout(n669));
  jor  g0355(.dina(n669), .dinb(n654), .dout(n670));
  jand g0356(.dina(n670), .dinb(n653), .dout(n671));
  jand g0357(.dina(n671), .dinb(n650), .dout(n672));
  jor  g0358(.dina(n672), .dinb(n647), .dout(n673));
  jor  g0359(.dina(n673), .dinb(n646), .dout(n674));
  jor  g0360(.dina(n673), .dinb(G4526), .dout(n675));
  jand g0361(.dina(n675), .dinb(n674), .dout(n676));
  jor  g0362(.dina(n676), .dinb(n621), .dout(n677));
  jand g0363(.dina(n677), .dinb(n620), .dout(n678));
  jand g0364(.dina(n678), .dinb(n589), .dout(n679));
  jor  g0365(.dina(n679), .dinb(n586), .dout(n680));
  jand g0366(.dina(n680), .dinb(n581), .dout(n681));
  jor  g0367(.dina(n681), .dinb(n572), .dout(n682));
  jand g0368(.dina(n682), .dinb(n527), .dout(n683));
  jand g0369(.dina(n683), .dinb(n524), .dout(n684));
  jand g0370(.dina(n684), .dinb(n519), .dout(n685));
  jand g0371(.dina(n685), .dinb(n513), .dout(n686));
  jand g0372(.dina(n512), .dinb(n509), .dout(n687));
  jnot g0373(.din(n687), .dout(n688));
  jnot g0374(.din(n512), .dout(n689));
  jand g0375(.dina(n689), .dinb(G4432), .dout(n690));
  jand g0376(.dina(n523), .dinb(n520), .dout(n691));
  jand g0377(.dina(n524), .dinb(n518), .dout(n692));
  jor  g0378(.dina(n692), .dinb(n691), .dout(n693));
  jnot g0379(.din(n693), .dout(n694));
  jor  g0380(.dina(n694), .dinb(n690), .dout(n695));
  jand g0381(.dina(n695), .dinb(n688), .dout(n696));
  jnot g0382(.din(n696), .dout(n697));
  jor  g0383(.dina(n697), .dinb(n686), .dout(n698));
  jand g0384(.dina(n698), .dinb(n508), .dout(n699));
  jor  g0385(.dina(n699), .dinb(n505), .dout(n700));
  jor  g0386(.dina(n700), .dinb(n462), .dout(n701));
  jor  g0387(.dina(n701), .dinb(n500), .dout(n702));
  jand g0388(.dina(n702), .dinb(n499), .dout(n703));
  jor  g0389(.dina(n703), .dinb(n449), .dout(n704));
  jand g0390(.dina(n704), .dinb(n450), .dout(n705));
  jand g0391(.dina(n705), .dinb(n425), .dout(n706));
  jor  g0392(.dina(n706), .dinb(n424), .dout(n707));
  jor  g0393(.dina(n707), .dinb(n413), .dout(n708));
  jand g0394(.dina(n708), .dinb(n420), .dout(n709));
  jand g0395(.dina(n709), .dinb(n370), .dout(n710));
  jand g0396(.dina(n710), .dinb(n363), .dout(n711));
  jnot g0397(.din(n362), .dout(n712));
  jand g0398(.dina(n712), .dinb(G38), .dout(n713));
  jand g0399(.dina(n366), .dinb(G38), .dout(n714));
  jor  g0400(.dina(n714), .dinb(n713), .dout(n715));
  jor  g0401(.dina(n715), .dinb(n711), .dout(G246));
  jand g0402(.dina(G2204), .dinb(G1455), .dout(n717));
  jor  g0403(.dina(n717), .dinb(n368), .dout(n718));
  jor  g0404(.dina(G166), .dinb(n355), .dout(n719));
  jand g0405(.dina(n719), .dinb(n373), .dout(n720));
  jor  g0406(.dina(n371), .dinb(n355), .dout(n721));
  jor  g0407(.dina(G88), .dinb(G18), .dout(n722));
  jand g0408(.dina(n722), .dinb(n721), .dout(n723));
  jxor g0409(.dina(n723), .dinb(n720), .dout(n724));
  jor  g0410(.dina(G167), .dinb(n355), .dout(n725));
  jand g0411(.dina(n725), .dinb(n373), .dout(n726));
  jor  g0412(.dina(n383), .dinb(n355), .dout(n727));
  jor  g0413(.dina(G112), .dinb(G18), .dout(n728));
  jand g0414(.dina(n728), .dinb(n727), .dout(n729));
  jor  g0415(.dina(n729), .dinb(n726), .dout(n730));
  jand g0416(.dina(n729), .dinb(n726), .dout(n731));
  jor  g0417(.dina(n389), .dinb(n355), .dout(n732));
  jor  g0418(.dina(G113), .dinb(G18), .dout(n733));
  jand g0419(.dina(n733), .dinb(n732), .dout(n734));
  jand g0420(.dina(n734), .dinb(n373), .dout(n735));
  jor  g0421(.dina(G168), .dinb(n355), .dout(n736));
  jand g0422(.dina(n736), .dinb(n373), .dout(n737));
  jand g0423(.dina(G106), .dinb(G18), .dout(n738));
  jnot g0424(.din(n738), .dout(n739));
  jor  g0425(.dina(G87), .dinb(G18), .dout(n740));
  jand g0426(.dina(n740), .dinb(n739), .dout(n741));
  jxor g0427(.dina(n741), .dinb(n737), .dout(n742));
  jor  g0428(.dina(G169), .dinb(n355), .dout(n743));
  jand g0429(.dina(n743), .dinb(n373), .dout(n744));
  jor  g0430(.dina(n393), .dinb(n355), .dout(n745));
  jor  g0431(.dina(G111), .dinb(G18), .dout(n746));
  jand g0432(.dina(n746), .dinb(n745), .dout(n747));
  jxor g0433(.dina(n747), .dinb(n744), .dout(n748));
  jand g0434(.dina(n748), .dinb(n742), .dout(n749));
  jand g0435(.dina(n749), .dinb(n735), .dout(n750));
  jor  g0436(.dina(n750), .dinb(n731), .dout(n751));
  jand g0437(.dina(n751), .dinb(n730), .dout(n752));
  jand g0438(.dina(n752), .dinb(n724), .dout(n753));
  jor  g0439(.dina(G173), .dinb(n355), .dout(n754));
  jand g0440(.dina(n754), .dinb(n373), .dout(n755));
  jor  g0441(.dina(n421), .dinb(n355), .dout(n756));
  jor  g0442(.dina(G110), .dinb(G18), .dout(n757));
  jand g0443(.dina(n757), .dinb(n756), .dout(n758));
  jxor g0444(.dina(n758), .dinb(n755), .dout(n759));
  jor  g0445(.dina(G174), .dinb(n355), .dout(n760));
  jand g0446(.dina(n760), .dinb(n373), .dout(n761));
  jor  g0447(.dina(n426), .dinb(n355), .dout(n762));
  jor  g0448(.dina(G109), .dinb(G18), .dout(n763));
  jand g0449(.dina(n763), .dinb(n762), .dout(n764));
  jxor g0450(.dina(n764), .dinb(n761), .dout(n765));
  jand g0451(.dina(n765), .dinb(n759), .dout(n766));
  jor  g0452(.dina(G175), .dinb(n355), .dout(n767));
  jand g0453(.dina(n767), .dinb(n373), .dout(n768));
  jand g0454(.dina(G2247), .dinb(G18), .dout(n769));
  jnot g0455(.din(n769), .dout(n770));
  jor  g0456(.dina(G86), .dinb(G18), .dout(n771));
  jand g0457(.dina(n771), .dinb(n770), .dout(n772));
  jand g0458(.dina(n772), .dinb(n768), .dout(n773));
  jor  g0459(.dina(n772), .dinb(n768), .dout(n774));
  jor  g0460(.dina(G176), .dinb(n355), .dout(n775));
  jand g0461(.dina(n775), .dinb(n373), .dout(n776));
  jand g0462(.dina(G2239), .dinb(G18), .dout(n777));
  jnot g0463(.din(n777), .dout(n778));
  jor  g0464(.dina(G63), .dinb(G18), .dout(n779));
  jand g0465(.dina(n779), .dinb(n778), .dout(n780));
  jand g0466(.dina(n780), .dinb(n776), .dout(n781));
  jand g0467(.dina(n781), .dinb(n774), .dout(n782));
  jor  g0468(.dina(n782), .dinb(n773), .dout(n783));
  jand g0469(.dina(n783), .dinb(n766), .dout(n784));
  jand g0470(.dina(n758), .dinb(n755), .dout(n785));
  jor  g0471(.dina(n758), .dinb(n755), .dout(n786));
  jand g0472(.dina(n764), .dinb(n761), .dout(n787));
  jand g0473(.dina(n787), .dinb(n786), .dout(n788));
  jor  g0474(.dina(n788), .dinb(n785), .dout(n789));
  jor  g0475(.dina(n789), .dinb(n784), .dout(n790));
  jnot g0476(.din(n773), .dout(n791));
  jnot g0477(.din(n781), .dout(n792));
  jand g0478(.dina(n792), .dinb(n791), .dout(n793));
  jand g0479(.dina(n793), .dinb(n766), .dout(n794));
  jor  g0480(.dina(G177), .dinb(n355), .dout(n795));
  jand g0481(.dina(n795), .dinb(n373), .dout(n796));
  jand g0482(.dina(G2236), .dinb(G18), .dout(n797));
  jnot g0483(.din(n797), .dout(n798));
  jor  g0484(.dina(G64), .dinb(G18), .dout(n799));
  jand g0485(.dina(n799), .dinb(n798), .dout(n800));
  jxor g0486(.dina(n800), .dinb(n796), .dout(n801));
  jand g0487(.dina(G178), .dinb(G18), .dout(n802));
  jor  g0488(.dina(n802), .dinb(n457), .dout(n803));
  jor  g0489(.dina(n456), .dinb(n355), .dout(n804));
  jor  g0490(.dina(G85), .dinb(G18), .dout(n805));
  jand g0491(.dina(n805), .dinb(n804), .dout(n806));
  jxor g0492(.dina(n806), .dinb(n803), .dout(n807));
  jand g0493(.dina(n807), .dinb(n801), .dout(n808));
  jand g0494(.dina(G179), .dinb(G18), .dout(n809));
  jor  g0495(.dina(n809), .dinb(n467), .dout(n810));
  jand g0496(.dina(G2224), .dinb(G18), .dout(n811));
  jnot g0497(.din(n811), .dout(n812));
  jor  g0498(.dina(G84), .dinb(G18), .dout(n813));
  jand g0499(.dina(n813), .dinb(n812), .dout(n814));
  jxor g0500(.dina(n814), .dinb(n810), .dout(n815));
  jand g0501(.dina(G180), .dinb(G18), .dout(n816));
  jor  g0502(.dina(n816), .dinb(n472), .dout(n817));
  jor  g0503(.dina(n471), .dinb(n355), .dout(n818));
  jor  g0504(.dina(G83), .dinb(G18), .dout(n819));
  jand g0505(.dina(n819), .dinb(n818), .dout(n820));
  jxor g0506(.dina(n820), .dinb(n817), .dout(n821));
  jand g0507(.dina(n821), .dinb(n815), .dout(n822));
  jand g0508(.dina(G171), .dinb(G18), .dout(n823));
  jor  g0509(.dina(n823), .dinb(n477), .dout(n824));
  jor  g0510(.dina(n476), .dinb(n355), .dout(n825));
  jor  g0511(.dina(G65), .dinb(G18), .dout(n826));
  jand g0512(.dina(n826), .dinb(n825), .dout(n827));
  jand g0513(.dina(n827), .dinb(n824), .dout(n828));
  jand g0514(.dina(n828), .dinb(n822), .dout(n829));
  jand g0515(.dina(n814), .dinb(n810), .dout(n830));
  jor  g0516(.dina(n814), .dinb(n810), .dout(n831));
  jand g0517(.dina(n820), .dinb(n817), .dout(n832));
  jand g0518(.dina(n832), .dinb(n831), .dout(n833));
  jor  g0519(.dina(n833), .dinb(n830), .dout(n834));
  jor  g0520(.dina(n834), .dinb(n829), .dout(n835));
  jand g0521(.dina(n835), .dinb(n808), .dout(n836));
  jand g0522(.dina(n800), .dinb(n796), .dout(n837));
  jor  g0523(.dina(n800), .dinb(n796), .dout(n838));
  jand g0524(.dina(n806), .dinb(n803), .dout(n839));
  jand g0525(.dina(n839), .dinb(n838), .dout(n840));
  jor  g0526(.dina(n840), .dinb(n837), .dout(n841));
  jor  g0527(.dina(n841), .dinb(n836), .dout(n842));
  jand g0528(.dina(n822), .dinb(n808), .dout(n843));
  jand g0529(.dina(G189), .dinb(G18), .dout(n844));
  jor  g0530(.dina(n844), .dinb(n503), .dout(n845));
  jor  g0531(.dina(n501), .dinb(n355), .dout(n846));
  jor  g0532(.dina(G62), .dinb(G18), .dout(n847));
  jand g0533(.dina(n847), .dinb(n846), .dout(n848));
  jxor g0534(.dina(n848), .dinb(n845), .dout(n849));
  jand g0535(.dina(G190), .dinb(G18), .dout(n850));
  jor  g0536(.dina(n850), .dinb(n511), .dout(n851));
  jor  g0537(.dina(n509), .dinb(n355), .dout(n852));
  jor  g0538(.dina(G61), .dinb(G18), .dout(n853));
  jand g0539(.dina(n853), .dinb(n852), .dout(n854));
  jxor g0540(.dina(n854), .dinb(n851), .dout(n855));
  jand g0541(.dina(n855), .dinb(n849), .dout(n856));
  jand g0542(.dina(G191), .dinb(G18), .dout(n857));
  jor  g0543(.dina(n857), .dinb(n522), .dout(n858));
  jand g0544(.dina(G4427), .dinb(G18), .dout(n859));
  jnot g0545(.din(n859), .dout(n860));
  jor  g0546(.dina(G60), .dinb(G18), .dout(n861));
  jand g0547(.dina(n861), .dinb(n860), .dout(n862));
  jand g0548(.dina(n862), .dinb(n858), .dout(n863));
  jor  g0549(.dina(n862), .dinb(n858), .dout(n864));
  jand g0550(.dina(G192), .dinb(G18), .dout(n865));
  jor  g0551(.dina(n865), .dinb(n516), .dout(n866));
  jand g0552(.dina(G4420), .dinb(G18), .dout(n867));
  jnot g0553(.din(n867), .dout(n868));
  jor  g0554(.dina(G79), .dinb(G18), .dout(n869));
  jand g0555(.dina(n869), .dinb(n868), .dout(n870));
  jand g0556(.dina(n870), .dinb(n866), .dout(n871));
  jand g0557(.dina(n871), .dinb(n864), .dout(n872));
  jor  g0558(.dina(n872), .dinb(n863), .dout(n873));
  jand g0559(.dina(n873), .dinb(n856), .dout(n874));
  jand g0560(.dina(n848), .dinb(n845), .dout(n875));
  jor  g0561(.dina(n848), .dinb(n845), .dout(n876));
  jand g0562(.dina(n854), .dinb(n851), .dout(n877));
  jand g0563(.dina(n877), .dinb(n876), .dout(n878));
  jor  g0564(.dina(n878), .dinb(n875), .dout(n879));
  jor  g0565(.dina(n879), .dinb(n874), .dout(n880));
  jor  g0566(.dina(n870), .dinb(n866), .dout(n881));
  jand g0567(.dina(n881), .dinb(n864), .dout(n882));
  jand g0568(.dina(n882), .dinb(n856), .dout(n883));
  jand g0569(.dina(G205), .dinb(G18), .dout(n884));
  jor  g0570(.dina(n884), .dinb(n629), .dout(n885));
  jor  g0571(.dina(n627), .dinb(n355), .dout(n886));
  jor  g0572(.dina(G75), .dinb(G18), .dout(n887));
  jand g0573(.dina(n887), .dinb(n886), .dout(n888));
  jor  g0574(.dina(n888), .dinb(n885), .dout(n889));
  jand g0575(.dina(G206), .dinb(G18), .dout(n890));
  jor  g0576(.dina(n890), .dinb(n634), .dout(n891));
  jor  g0577(.dina(n632), .dinb(n355), .dout(n892));
  jor  g0578(.dina(G76), .dinb(G18), .dout(n893));
  jand g0579(.dina(n893), .dinb(n892), .dout(n894));
  jand g0580(.dina(n894), .dinb(n891), .dout(n895));
  jor  g0581(.dina(G89), .dinb(G70), .dout(n896));
  jand g0582(.dina(n896), .dinb(n663), .dout(n897));
  jor  g0583(.dina(n897), .dinb(n895), .dout(n898));
  jand g0584(.dina(G207), .dinb(G18), .dout(n899));
  jor  g0585(.dina(n899), .dinb(n659), .dout(n900));
  jor  g0586(.dina(n657), .dinb(n355), .dout(n901));
  jor  g0587(.dina(G74), .dinb(G18), .dout(n902));
  jand g0588(.dina(n902), .dinb(n901), .dout(n903));
  jand g0589(.dina(n903), .dinb(n900), .dout(n904));
  jor  g0590(.dina(G70), .dinb(G18), .dout(n905));
  jand g0591(.dina(n905), .dinb(G89), .dout(n906));
  jor  g0592(.dina(n906), .dinb(n904), .dout(n907));
  jor  g0593(.dina(n907), .dinb(n898), .dout(n908));
  jor  g0594(.dina(n903), .dinb(n900), .dout(n909));
  jor  g0595(.dina(n894), .dinb(n891), .dout(n910));
  jand g0596(.dina(n910), .dinb(n909), .dout(n911));
  jor  g0597(.dina(n911), .dinb(n895), .dout(n912));
  jand g0598(.dina(n912), .dinb(n908), .dout(n913));
  jand g0599(.dina(n913), .dinb(n889), .dout(n914));
  jand g0600(.dina(G204), .dinb(G18), .dout(n915));
  jor  g0601(.dina(n915), .dinb(n624), .dout(n916));
  jor  g0602(.dina(n622), .dinb(n355), .dout(n917));
  jor  g0603(.dina(G73), .dinb(G18), .dout(n918));
  jand g0604(.dina(n918), .dinb(n917), .dout(n919));
  jand g0605(.dina(n919), .dinb(n916), .dout(n920));
  jand g0606(.dina(n888), .dinb(n885), .dout(n921));
  jor  g0607(.dina(n921), .dinb(n920), .dout(n922));
  jor  g0608(.dina(n922), .dinb(n914), .dout(n923));
  jor  g0609(.dina(n919), .dinb(n916), .dout(n924));
  jand g0610(.dina(G203), .dinb(G18), .dout(n925));
  jor  g0611(.dina(n925), .dinb(n602), .dout(n926));
  jand g0612(.dina(G3729), .dinb(G18), .dout(n927));
  jnot g0613(.din(n927), .dout(n928));
  jor  g0614(.dina(G53), .dinb(G18), .dout(n929));
  jand g0615(.dina(n929), .dinb(n928), .dout(n930));
  jor  g0616(.dina(n930), .dinb(n926), .dout(n931));
  jand g0617(.dina(n931), .dinb(n924), .dout(n932));
  jand g0618(.dina(n932), .dinb(n923), .dout(n933));
  jand g0619(.dina(G202), .dinb(G18), .dout(n934));
  jor  g0620(.dina(n934), .dinb(n597), .dout(n935));
  jor  g0621(.dina(n595), .dinb(n355), .dout(n936));
  jor  g0622(.dina(G54), .dinb(G18), .dout(n937));
  jand g0623(.dina(n937), .dinb(n936), .dout(n938));
  jand g0624(.dina(n938), .dinb(n935), .dout(n939));
  jand g0625(.dina(n930), .dinb(n926), .dout(n940));
  jor  g0626(.dina(n940), .dinb(n939), .dout(n941));
  jor  g0627(.dina(n941), .dinb(n933), .dout(n942));
  jand g0628(.dina(G201), .dinb(G18), .dout(n943));
  jor  g0629(.dina(n943), .dinb(n592), .dout(n944));
  jor  g0630(.dina(n590), .dinb(n355), .dout(n945));
  jor  g0631(.dina(G55), .dinb(G18), .dout(n946));
  jand g0632(.dina(n946), .dinb(n945), .dout(n947));
  jxor g0633(.dina(n947), .dinb(n944), .dout(n948));
  jand g0634(.dina(G200), .dinb(G18), .dout(n949));
  jor  g0635(.dina(n949), .dinb(n584), .dout(n950));
  jor  g0636(.dina(n582), .dinb(n355), .dout(n951));
  jor  g0637(.dina(G56), .dinb(G18), .dout(n952));
  jand g0638(.dina(n952), .dinb(n951), .dout(n953));
  jxor g0639(.dina(n953), .dinb(n950), .dout(n954));
  jand g0640(.dina(n954), .dinb(n948), .dout(n955));
  jor  g0641(.dina(n938), .dinb(n935), .dout(n956));
  jand g0642(.dina(n956), .dinb(n955), .dout(n957));
  jand g0643(.dina(n957), .dinb(n942), .dout(n958));
  jand g0644(.dina(n953), .dinb(n950), .dout(n959));
  jand g0645(.dina(n947), .dinb(n944), .dout(n960));
  jor  g0646(.dina(n953), .dinb(n950), .dout(n961));
  jand g0647(.dina(n961), .dinb(n960), .dout(n962));
  jor  g0648(.dina(n962), .dinb(n959), .dout(n963));
  jor  g0649(.dina(n963), .dinb(n958), .dout(n964));
  jand g0650(.dina(G187), .dinb(G18), .dout(n965));
  jor  g0651(.dina(n965), .dinb(n562), .dout(n966));
  jand g0652(.dina(G4394), .dinb(G18), .dout(n967));
  jnot g0653(.din(n967), .dout(n968));
  jor  g0654(.dina(G77), .dinb(G18), .dout(n969));
  jand g0655(.dina(n969), .dinb(n968), .dout(n970));
  jor  g0656(.dina(n970), .dinb(n966), .dout(n971));
  jand g0657(.dina(G193), .dinb(G18), .dout(n972));
  jor  g0658(.dina(n972), .dinb(n530), .dout(n973));
  jand g0659(.dina(G4415), .dinb(G18), .dout(n974));
  jnot g0660(.din(n974), .dout(n975));
  jor  g0661(.dina(G80), .dinb(G18), .dout(n976));
  jand g0662(.dina(n976), .dinb(n975), .dout(n977));
  jxor g0663(.dina(n977), .dinb(n973), .dout(n978));
  jand g0664(.dina(G194), .dinb(G18), .dout(n979));
  jor  g0665(.dina(n979), .dinb(n538), .dout(n980));
  jor  g0666(.dina(n536), .dinb(n355), .dout(n981));
  jor  g0667(.dina(G81), .dinb(G18), .dout(n982));
  jand g0668(.dina(n982), .dinb(n981), .dout(n983));
  jxor g0669(.dina(n983), .dinb(n980), .dout(n984));
  jand g0670(.dina(n984), .dinb(n978), .dout(n985));
  jand g0671(.dina(G196), .dinb(G18), .dout(n986));
  jor  g0672(.dina(n986), .dinb(n554), .dout(n987));
  jand g0673(.dina(G4400), .dinb(G18), .dout(n988));
  jnot g0674(.din(n988), .dout(n989));
  jor  g0675(.dina(G78), .dinb(G18), .dout(n990));
  jand g0676(.dina(n990), .dinb(n989), .dout(n991));
  jand g0677(.dina(n991), .dinb(n987), .dout(n992));
  jnot g0678(.din(n992), .dout(n993));
  jand g0679(.dina(G195), .dinb(G18), .dout(n994));
  jor  g0680(.dina(n994), .dinb(n546), .dout(n995));
  jand g0681(.dina(G4405), .dinb(G18), .dout(n996));
  jnot g0682(.din(n996), .dout(n997));
  jor  g0683(.dina(G59), .dinb(G18), .dout(n998));
  jand g0684(.dina(n998), .dinb(n997), .dout(n999));
  jor  g0685(.dina(n999), .dinb(n995), .dout(n1000));
  jand g0686(.dina(n1000), .dinb(n993), .dout(n1001));
  jor  g0687(.dina(n991), .dinb(n987), .dout(n1002));
  jand g0688(.dina(n999), .dinb(n995), .dout(n1003));
  jnot g0689(.din(n1003), .dout(n1004));
  jand g0690(.dina(n1004), .dinb(n1002), .dout(n1005));
  jand g0691(.dina(n1005), .dinb(n1001), .dout(n1006));
  jand g0692(.dina(n1006), .dinb(n985), .dout(n1007));
  jand g0693(.dina(n970), .dinb(n966), .dout(n1008));
  jnot g0694(.din(n1008), .dout(n1009));
  jand g0695(.dina(n1009), .dinb(n1007), .dout(n1010));
  jand g0696(.dina(n1010), .dinb(n971), .dout(n1011));
  jand g0697(.dina(n1011), .dinb(n964), .dout(n1012));
  jand g0698(.dina(n977), .dinb(n973), .dout(n1013));
  jor  g0699(.dina(n977), .dinb(n973), .dout(n1014));
  jand g0700(.dina(n983), .dinb(n980), .dout(n1015));
  jand g0701(.dina(n1015), .dinb(n1014), .dout(n1016));
  jor  g0702(.dina(n1016), .dinb(n1013), .dout(n1017));
  jand g0703(.dina(n1008), .dinb(n1007), .dout(n1018));
  jand g0704(.dina(n1000), .dinb(n992), .dout(n1019));
  jor  g0705(.dina(n1019), .dinb(n1003), .dout(n1020));
  jand g0706(.dina(n1020), .dinb(n985), .dout(n1021));
  jor  g0707(.dina(n1021), .dinb(n1018), .dout(n1022));
  jor  g0708(.dina(n1022), .dinb(n1017), .dout(n1023));
  jor  g0709(.dina(n1023), .dinb(n1012), .dout(n1024));
  jnot g0710(.din(n863), .dout(n1025));
  jnot g0711(.din(n871), .dout(n1026));
  jand g0712(.dina(n1026), .dinb(n1025), .dout(n1027));
  jand g0713(.dina(n1027), .dinb(n1024), .dout(n1028));
  jand g0714(.dina(n1028), .dinb(n883), .dout(n1029));
  jor  g0715(.dina(n1029), .dinb(n880), .dout(G252));
  jxor g0716(.dina(n827), .dinb(n824), .dout(n1031));
  jand g0717(.dina(n1031), .dinb(G252), .dout(n1032));
  jand g0718(.dina(n1032), .dinb(n843), .dout(n1033));
  jor  g0719(.dina(n1033), .dinb(n842), .dout(n1034));
  jor  g0720(.dina(n780), .dinb(n776), .dout(n1035));
  jand g0721(.dina(n1035), .dinb(n774), .dout(n1036));
  jand g0722(.dina(n1036), .dinb(n1034), .dout(n1037));
  jand g0723(.dina(n1037), .dinb(n794), .dout(n1038));
  jor  g0724(.dina(n1038), .dinb(n790), .dout(n1039));
  jxor g0725(.dina(n734), .dinb(n373), .dout(n1040));
  jxor g0726(.dina(n729), .dinb(n726), .dout(n1041));
  jand g0727(.dina(n1041), .dinb(n724), .dout(n1042));
  jand g0728(.dina(n1042), .dinb(n749), .dout(n1043));
  jand g0729(.dina(n1043), .dinb(n1040), .dout(n1044));
  jand g0730(.dina(n1044), .dinb(n1039), .dout(n1045));
  jor  g0731(.dina(G2204), .dinb(G1455), .dout(n1046));
  jor  g0732(.dina(n1046), .dinb(n367), .dout(n1047));
  jand g0733(.dina(n1047), .dinb(G38), .dout(n1048));
  jand g0734(.dina(n723), .dinb(n720), .dout(n1049));
  jand g0735(.dina(n741), .dinb(n737), .dout(n1050));
  jor  g0736(.dina(n741), .dinb(n737), .dout(n1051));
  jand g0737(.dina(n747), .dinb(n744), .dout(n1052));
  jand g0738(.dina(n1052), .dinb(n1051), .dout(n1053));
  jor  g0739(.dina(n1053), .dinb(n1050), .dout(n1054));
  jand g0740(.dina(n1054), .dinb(n1042), .dout(n1055));
  jor  g0741(.dina(n1055), .dinb(n1049), .dout(n1056));
  jor  g0742(.dina(n1056), .dinb(n1048), .dout(n1057));
  jor  g0743(.dina(n1057), .dinb(n1045), .dout(n1058));
  jor  g0744(.dina(n1058), .dinb(n753), .dout(n1059));
  jand g0745(.dina(n1059), .dinb(n718), .dout(G258));
  jnot g0746(.din(n644), .dout(n1061));
  jnot g0747(.din(n655), .dout(n1062));
  jnot g0748(.din(n656), .dout(n1063));
  jand g0749(.dina(n641), .dinb(G3705), .dout(n1064));
  jor  g0750(.dina(n641), .dinb(G3705), .dout(n1065));
  jand g0751(.dina(n1065), .dinb(n354), .dout(n1066));
  jor  g0752(.dina(n1066), .dinb(n1064), .dout(n1067));
  jor  g0753(.dina(n1067), .dinb(n1063), .dout(n1068));
  jand g0754(.dina(n1068), .dinb(n1062), .dout(n1069));
  jand g0755(.dina(n1069), .dinb(n1061), .dout(n1070));
  jnot g0756(.din(n1070), .dout(n1071));
  jor  g0757(.dina(n669), .dinb(G4526), .dout(n1072));
  jand g0758(.dina(n1072), .dinb(n1071), .dout(n1073));
  jor  g0759(.dina(n1073), .dinb(n654), .dout(n1074));
  jand g0760(.dina(n1074), .dinb(n653), .dout(n1075));
  jxor g0761(.dina(n1075), .dinb(n626), .dout(G388));
  jxor g0762(.dina(n1073), .dinb(n631), .dout(G391));
  jand g0763(.dina(n359), .dinb(G4526), .dout(n1078));
  jor  g0764(.dina(n666), .dinb(n1078), .dout(n1079));
  jand g0765(.dina(n1079), .dinb(n661), .dout(n1080));
  jxor g0766(.dina(n1080), .dinb(n636), .dout(G394));
  jor  g0767(.dina(n1078), .dinb(n664), .dout(n1082));
  jxor g0768(.dina(n1082), .dinb(n642), .dout(G397));
  jxor g0769(.dina(n585), .dinb(n582), .dout(n1084));
  jor  g0770(.dina(n1084), .dinb(n678), .dout(n1085));
  jnot g0771(.din(n646), .dout(n1086));
  jnot g0772(.din(n647), .dout(n1087));
  jnot g0773(.din(n654), .dout(n1088));
  jand g0774(.dina(n1069), .dinb(n1088), .dout(n1089));
  jor  g0775(.dina(n1089), .dinb(n652), .dout(n1090));
  jor  g0776(.dina(n1090), .dinb(n649), .dout(n1091));
  jand g0777(.dina(n1091), .dinb(n1087), .dout(n1092));
  jand g0778(.dina(n1092), .dinb(n1086), .dout(n1093));
  jnot g0779(.din(G4526), .dout(n1094));
  jand g0780(.dina(n1092), .dinb(n1094), .dout(n1095));
  jor  g0781(.dina(n1095), .dinb(n1093), .dout(n1096));
  jand g0782(.dina(n1096), .dinb(n618), .dout(n1097));
  jor  g0783(.dina(n1097), .dinb(n619), .dout(n1098));
  jor  g0784(.dina(n1098), .dinb(n588), .dout(n1099));
  jor  g0785(.dina(n1099), .dinb(n586), .dout(n1100));
  jand g0786(.dina(n1100), .dinb(n1085), .dout(G376));
  jand g0787(.dina(n676), .dinb(n605), .dout(n1102));
  jor  g0788(.dina(n1102), .dinb(n615), .dout(n1103));
  jxor g0789(.dina(n1103), .dinb(n594), .dout(G379));
  jnot g0790(.din(n599), .dout(n1105));
  jnot g0791(.din(n613), .dout(n1106));
  jnot g0792(.din(n603), .dout(n1107));
  jand g0793(.dina(n1107), .dinb(G3729), .dout(n1108));
  jor  g0794(.dina(n1096), .dinb(n1108), .dout(n1109));
  jand g0795(.dina(n1109), .dinb(n1106), .dout(n1110));
  jxor g0796(.dina(n1110), .dinb(n1105), .dout(G382));
  jxor g0797(.dina(n676), .dinb(n604), .dout(G385));
  jnot g0798(.din(n436), .dout(n1113));
  jor  g0799(.dina(n1113), .dinb(n431), .dout(n1114));
  jnot g0800(.din(n432), .dout(n1115));
  jor  g0801(.dina(n435), .dinb(n1115), .dout(n1116));
  jand g0802(.dina(n1116), .dinb(n1114), .dout(n1117));
  jnot g0803(.din(n459), .dout(n1118));
  jxor g0804(.dina(n1118), .dinb(n453), .dout(n1119));
  jxor g0805(.dina(n1119), .dinb(n1117), .dout(n1120));
  jxor g0806(.dina(n485), .dinb(n469), .dout(n1121));
  jor  g0807(.dina(n440), .dinb(n422), .dout(n1122));
  jnot g0808(.din(n423), .dout(n1123));
  jor  g0809(.dina(n427), .dinb(n1123), .dout(n1124));
  jand g0810(.dina(n1124), .dinb(n1122), .dout(n1125));
  jnot g0811(.din(G141), .dout(n1126));
  jor  g0812(.dina(n1126), .dinb(G18), .dout(n1127));
  jnot g0813(.din(G161), .dout(n1128));
  jor  g0814(.dina(n1128), .dinb(n355), .dout(n1129));
  jand g0815(.dina(n1129), .dinb(n1127), .dout(n1130));
  jxor g0816(.dina(n1130), .dinb(n479), .dout(n1131));
  jxor g0817(.dina(n1131), .dinb(n1125), .dout(n1132));
  jxor g0818(.dina(n1132), .dinb(n1121), .dout(n1133));
  jxor g0819(.dina(n1133), .dinb(n1120), .dout(n1134));
  jxor g0820(.dina(n603), .dinb(n598), .dout(n1135));
  jand g0821(.dina(G239), .dinb(G18), .dout(n1136));
  jand g0822(.dina(G44), .dinb(n355), .dout(n1137));
  jor  g0823(.dina(n1137), .dinb(n1136), .dout(n1138));
  jxor g0824(.dina(n1138), .dinb(n651), .dout(n1139));
  jxor g0825(.dina(n1139), .dinb(n1135), .dout(n1140));
  jand g0826(.dina(G229), .dinb(G18), .dout(n1141));
  jor  g0827(.dina(n1141), .dinb(n663), .dout(n1142));
  jxor g0828(.dina(n1142), .dinb(n660), .dout(n1143));
  jxor g0829(.dina(n635), .dinb(n625), .dout(n1144));
  jxor g0830(.dina(n1144), .dinb(n1143), .dout(n1145));
  jxor g0831(.dina(n593), .dinb(n585), .dout(n1146));
  jxor g0832(.dina(n1146), .dinb(n1145), .dout(n1147));
  jxor g0833(.dina(n1147), .dinb(n1140), .dout(n1148));
  jor  g0834(.dina(n1148), .dinb(n1134), .dout(n1149));
  jor  g0835(.dina(n372), .dinb(n355), .dout(n1150));
  jxor g0836(.dina(G212), .dinb(G211), .dout(n1151));
  jxor g0837(.dina(n1151), .dinb(G209), .dout(n1152));
  jor  g0838(.dina(n1152), .dinb(n1150), .dout(n1153));
  jnot g0839(.din(n386), .dout(n1154));
  jand g0840(.dina(n395), .dinb(n1154), .dout(n1155));
  jnot g0841(.din(n394), .dout(n1156));
  jand g0842(.dina(n1156), .dinb(n387), .dout(n1157));
  jor  g0843(.dina(n1157), .dinb(n1155), .dout(n1158));
  jor  g0844(.dina(n380), .dinb(n374), .dout(n1159));
  jnot g0845(.din(n375), .dout(n1160));
  jor  g0846(.dina(n378), .dinb(n1160), .dout(n1161));
  jand g0847(.dina(n1161), .dinb(n1159), .dout(n1162));
  jxor g0848(.dina(n1162), .dinb(n1158), .dout(n1163));
  jxor g0849(.dina(n1163), .dinb(n1153), .dout(n1164));
  jxor g0850(.dina(n689), .dinb(n504), .dout(n1165));
  jxor g0851(.dina(n523), .dinb(n517), .dout(n1166));
  jxor g0852(.dina(n1166), .dinb(n1165), .dout(n1167));
  jxor g0853(.dina(n555), .dinb(n539), .dout(n1168));
  jxor g0854(.dina(n547), .dinb(n531), .dout(n1169));
  jxor g0855(.dina(n1169), .dinb(n1168), .dout(n1170));
  jand g0856(.dina(G227), .dinb(G18), .dout(n1171));
  jand g0857(.dina(G115), .dinb(n355), .dout(n1172));
  jor  g0858(.dina(n1172), .dinb(n1171), .dout(n1173));
  jxor g0859(.dina(n1173), .dinb(n563), .dout(n1174));
  jxor g0860(.dina(n1174), .dinb(n1170), .dout(n1175));
  jxor g0861(.dina(n1175), .dinb(n1167), .dout(n1176));
  jor  g0862(.dina(n1176), .dinb(n1164), .dout(n1177));
  jor  g0863(.dina(n1177), .dinb(n1149), .dout(G412));
  jnot g0864(.din(n772), .dout(n1179));
  jxor g0865(.dina(n780), .dinb(n1179), .dout(n1180));
  jnot g0866(.din(G2208), .dout(n1181));
  jor  g0867(.dina(n1181), .dinb(n355), .dout(n1182));
  jor  g0868(.dina(G82), .dinb(G18), .dout(n1183));
  jand g0869(.dina(n1183), .dinb(n1182), .dout(n1184));
  jxor g0870(.dina(n1184), .dinb(n827), .dout(n1185));
  jxor g0871(.dina(n1185), .dinb(n1180), .dout(n1186));
  jxor g0872(.dina(n806), .dinb(n800), .dout(n1187));
  jxor g0873(.dina(n820), .dinb(n814), .dout(n1188));
  jxor g0874(.dina(n1188), .dinb(n1187), .dout(n1189));
  jxor g0875(.dina(n764), .dinb(n758), .dout(n1190));
  jxor g0876(.dina(n1190), .dinb(n1189), .dout(n1191));
  jxor g0877(.dina(n1191), .dinb(n1186), .dout(n1192));
  jxor g0878(.dina(n953), .dinb(n947), .dout(n1193));
  jxor g0879(.dina(n903), .dinb(n894), .dout(n1194));
  jxor g0880(.dina(n1194), .dinb(n1193), .dout(n1195));
  jnot g0881(.din(G3698), .dout(n1196));
  jor  g0882(.dina(n1196), .dinb(n355), .dout(n1197));
  jor  g0883(.dina(G69), .dinb(G18), .dout(n1198));
  jand g0884(.dina(n1198), .dinb(n1197), .dout(n1199));
  jxor g0885(.dina(n1199), .dinb(n888), .dout(n1200));
  jor  g0886(.dina(n662), .dinb(n355), .dout(n1201));
  jand g0887(.dina(n1201), .dinb(n905), .dout(n1202));
  jxor g0888(.dina(n1202), .dinb(n919), .dout(n1203));
  jxor g0889(.dina(n1203), .dinb(n1200), .dout(n1204));
  jnot g0890(.din(n930), .dout(n1205));
  jxor g0891(.dina(n938), .dinb(n1205), .dout(n1206));
  jxor g0892(.dina(n1206), .dinb(n1204), .dout(n1207));
  jxor g0893(.dina(n1207), .dinb(n1195), .dout(n1208));
  jor  g0894(.dina(n1208), .dinb(n1192), .dout(n1209));
  jxor g0895(.dina(n854), .dinb(n848), .dout(n1210));
  jxor g0896(.dina(n870), .dinb(n862), .dout(n1211));
  jxor g0897(.dina(n1211), .dinb(n1210), .dout(n1212));
  jxor g0898(.dina(n983), .dinb(n977), .dout(n1213));
  jand g0899(.dina(G4393), .dinb(G18), .dout(n1214));
  jnot g0900(.din(G58), .dout(n1215));
  jand g0901(.dina(n1215), .dinb(n355), .dout(n1216));
  jor  g0902(.dina(n1216), .dinb(n1214), .dout(n1217));
  jxor g0903(.dina(n1217), .dinb(n970), .dout(n1218));
  jxor g0904(.dina(n999), .dinb(n991), .dout(n1219));
  jxor g0905(.dina(n1219), .dinb(n1218), .dout(n1220));
  jxor g0906(.dina(n1220), .dinb(n1213), .dout(n1221));
  jxor g0907(.dina(n1221), .dinb(n1212), .dout(n1222));
  jxor g0908(.dina(n366), .dinb(G1492), .dout(n1223));
  jor  g0909(.dina(n1223), .dinb(n355), .dout(n1224));
  jnot g0910(.din(G1455), .dout(n1225));
  jxor g0911(.dina(G2204), .dinb(n1225), .dout(n1226));
  jor  g0912(.dina(n1226), .dinb(G18), .dout(n1227));
  jand g0913(.dina(n1227), .dinb(n1224), .dout(n1228));
  jxor g0914(.dina(n729), .dinb(n723), .dout(n1229));
  jxor g0915(.dina(n747), .dinb(n741), .dout(n1230));
  jxor g0916(.dina(n1230), .dinb(n1229), .dout(n1231));
  jnot g0917(.din(G1459), .dout(n1232));
  jor  g0918(.dina(n1232), .dinb(n355), .dout(n1233));
  jor  g0919(.dina(G114), .dinb(G18), .dout(n1234));
  jand g0920(.dina(n1234), .dinb(n1233), .dout(n1235));
  jxor g0921(.dina(n1235), .dinb(n734), .dout(n1236));
  jxor g0922(.dina(n1236), .dinb(n1231), .dout(n1237));
  jxor g0923(.dina(n1237), .dinb(n1228), .dout(n1238));
  jor  g0924(.dina(n1238), .dinb(n1222), .dout(n1239));
  jor  g0925(.dina(n1239), .dinb(n1209), .dout(G414));
  jnot g0926(.din(n935), .dout(n1241));
  jxor g0927(.dina(n1241), .dinb(n926), .dout(n1242));
  jxor g0928(.dina(n950), .dinb(n944), .dout(n1243));
  jxor g0929(.dina(n1243), .dinb(n1242), .dout(n1244));
  jand g0930(.dina(G208), .dinb(G18), .dout(n1245));
  jor  g0931(.dina(n1245), .dinb(n1137), .dout(n1246));
  jand g0932(.dina(G198), .dinb(G18), .dout(n1247));
  jor  g0933(.dina(n1247), .dinb(n663), .dout(n1248));
  jxor g0934(.dina(n1248), .dinb(n1246), .dout(n1249));
  jxor g0935(.dina(n916), .dinb(n885), .dout(n1250));
  jxor g0936(.dina(n1250), .dinb(n1249), .dout(n1251));
  jxor g0937(.dina(n900), .dinb(n891), .dout(n1252));
  jxor g0938(.dina(n1252), .dinb(n1251), .dout(n1253));
  jxor g0939(.dina(n1253), .dinb(n1244), .dout(n1254));
  jxor g0940(.dina(n866), .dinb(n858), .dout(n1255));
  jxor g0941(.dina(n995), .dinb(n987), .dout(n1256));
  jxor g0942(.dina(n1256), .dinb(n1255), .dout(n1257));
  jxor g0943(.dina(n980), .dinb(n973), .dout(n1258));
  jand g0944(.dina(G197), .dinb(G18), .dout(n1259));
  jor  g0945(.dina(n1259), .dinb(n1172), .dout(n1260));
  jxor g0946(.dina(n1260), .dinb(n966), .dout(n1261));
  jxor g0947(.dina(n1261), .dinb(n1258), .dout(n1262));
  jnot g0948(.din(n851), .dout(n1263));
  jxor g0949(.dina(n1263), .dinb(n845), .dout(n1264));
  jxor g0950(.dina(n1264), .dinb(n1262), .dout(n1265));
  jxor g0951(.dina(n1265), .dinb(n1257), .dout(n1266));
  jor  g0952(.dina(n1266), .dinb(n1254), .dout(n1267));
  jxor g0953(.dina(G165), .dinb(G164), .dout(n1268));
  jxor g0954(.dina(n1268), .dinb(G170), .dout(n1269));
  jor  g0955(.dina(n1269), .dinb(n1150), .dout(n1270));
  jnot g0956(.din(n736), .dout(n1271));
  jand g0957(.dina(n744), .dinb(n1271), .dout(n1272));
  jnot g0958(.din(n743), .dout(n1273));
  jand g0959(.dina(n1273), .dinb(n737), .dout(n1274));
  jor  g0960(.dina(n1274), .dinb(n1272), .dout(n1275));
  jnot g0961(.din(n726), .dout(n1276));
  jor  g0962(.dina(n1276), .dinb(n719), .dout(n1277));
  jnot g0963(.din(n720), .dout(n1278));
  jor  g0964(.dina(n725), .dinb(n1278), .dout(n1279));
  jand g0965(.dina(n1279), .dinb(n1277), .dout(n1280));
  jxor g0966(.dina(n1280), .dinb(n1275), .dout(n1281));
  jxor g0967(.dina(n1281), .dinb(n1270), .dout(n1282));
  jor  g0968(.dina(n1282), .dinb(n1267), .dout(n1283));
  jnot g0969(.din(G181), .dout(n1284));
  jor  g0970(.dina(n1284), .dinb(n355), .dout(n1285));
  jand g0971(.dina(n1285), .dinb(n1127), .dout(n1286));
  jxor g0972(.dina(n1286), .dinb(n824), .dout(n1287));
  jxor g0973(.dina(n803), .dinb(n796), .dout(n1288));
  jxor g0974(.dina(n1288), .dinb(n1287), .dout(n1289));
  jnot g0975(.din(n767), .dout(n1290));
  jand g0976(.dina(n776), .dinb(n1290), .dout(n1291));
  jnot g0977(.din(n775), .dout(n1292));
  jand g0978(.dina(n1292), .dinb(n768), .dout(n1293));
  jor  g0979(.dina(n1293), .dinb(n1291), .dout(n1294));
  jnot g0980(.din(n754), .dout(n1295));
  jand g0981(.dina(n761), .dinb(n1295), .dout(n1296));
  jnot g0982(.din(n760), .dout(n1297));
  jand g0983(.dina(n1297), .dinb(n755), .dout(n1298));
  jor  g0984(.dina(n1298), .dinb(n1296), .dout(n1299));
  jxor g0985(.dina(n1299), .dinb(n1294), .dout(n1300));
  jxor g0986(.dina(n817), .dinb(n810), .dout(n1301));
  jxor g0987(.dina(n1301), .dinb(n1300), .dout(n1302));
  jxor g0988(.dina(n1302), .dinb(n1289), .dout(n1303));
  jor  g0989(.dina(n1303), .dinb(n1283), .dout(G416));
  jnot g0990(.din(n480), .dout(n1305));
  jnot g0991(.din(n505), .dout(n1306));
  jnot g0992(.din(n513), .dout(n1307));
  jnot g0993(.din(n524), .dout(n1308));
  jnot g0994(.din(n572), .dout(n1309));
  jnot g0995(.din(n581), .dout(n1310));
  jnot g0996(.din(n586), .dout(n1311));
  jand g0997(.dina(n1099), .dinb(n1311), .dout(n1312));
  jor  g0998(.dina(n1312), .dinb(n1310), .dout(n1313));
  jand g0999(.dina(n1313), .dinb(n1309), .dout(n1314));
  jor  g1000(.dina(n1314), .dinb(n526), .dout(n1315));
  jor  g1001(.dina(n1315), .dinb(n1308), .dout(n1316));
  jor  g1002(.dina(n1316), .dinb(n518), .dout(n1317));
  jor  g1003(.dina(n1317), .dinb(n1307), .dout(n1318));
  jand g1004(.dina(n696), .dinb(n1318), .dout(n1319));
  jor  g1005(.dina(n1319), .dinb(n507), .dout(n1320));
  jand g1006(.dina(n1320), .dinb(n1306), .dout(n1321));
  jxor g1007(.dina(n1321), .dinb(n1305), .dout(G295));
  jnot g1008(.din(n414), .dout(n1323));
  jnot g1009(.din(n424), .dout(n1324));
  jnot g1010(.din(n425), .dout(n1325));
  jnot g1011(.din(n450), .dout(n1326));
  jnot g1012(.din(n449), .dout(n1327));
  jnot g1013(.din(n499), .dout(n1328));
  jnot g1014(.din(n500), .dout(n1329));
  jnot g1015(.din(n462), .dout(n1330));
  jand g1016(.dina(n1321), .dinb(n1330), .dout(n1331));
  jand g1017(.dina(n1331), .dinb(n1329), .dout(n1332));
  jor  g1018(.dina(n1332), .dinb(n1328), .dout(n1333));
  jand g1019(.dina(n1333), .dinb(n1327), .dout(n1334));
  jor  g1020(.dina(n1334), .dinb(n1326), .dout(n1335));
  jor  g1021(.dina(n1335), .dinb(n1325), .dout(n1336));
  jand g1022(.dina(n1336), .dinb(n1324), .dout(n1337));
  jxor g1023(.dina(n1337), .dinb(n1323), .dout(G324));
  jand g1024(.dina(n1118), .dinb(G2230), .dout(n1339));
  jnot g1025(.din(n1339), .dout(n1340));
  jand g1026(.dina(n1321), .dinb(n495), .dout(n1341));
  jnot g1027(.din(n1341), .dout(n1342));
  jand g1028(.dina(n1342), .dinb(n497), .dout(n1343));
  jand g1029(.dina(n1343), .dinb(n1340), .dout(n1344));
  jor  g1030(.dina(n1344), .dinb(n460), .dout(n1345));
  jxor g1031(.dina(n1345), .dinb(n463), .dout(G310));
  jor  g1032(.dina(n1343), .dinb(n464), .dout(n1347));
  jnot g1033(.din(n1344), .dout(n1348));
  jor  g1034(.dina(n1348), .dinb(n460), .dout(n1349));
  jand g1035(.dina(n1349), .dinb(n1347), .dout(G313));
  jnot g1036(.din(n489), .dout(n1351));
  jor  g1037(.dina(n1351), .dinb(n491), .dout(n1352));
  jand g1038(.dina(n700), .dinb(n481), .dout(n1353));
  jor  g1039(.dina(n1353), .dinb(n1352), .dout(n1354));
  jxor g1040(.dina(n1354), .dinb(n470), .dout(G316));
  jand g1041(.dina(n700), .dinb(n480), .dout(n1356));
  jor  g1042(.dina(n1356), .dinb(n487), .dout(n1357));
  jxor g1043(.dina(n1357), .dinb(n475), .dout(G319));
  jor  g1044(.dina(n418), .dinb(n411), .dout(n1359));
  jor  g1045(.dina(n707), .dinb(n411), .dout(n1360));
  jand g1046(.dina(n1360), .dinb(n1359), .dout(n1361));
  jxor g1047(.dina(n1361), .dinb(n377), .dout(G327));
  jand g1048(.dina(n415), .dinb(n388), .dout(n1363));
  jor  g1049(.dina(n1363), .dinb(n409), .dout(n1364));
  jor  g1050(.dina(n707), .dinb(n409), .dout(n1365));
  jand g1051(.dina(n1365), .dinb(n1364), .dout(n1366));
  jxor g1052(.dina(n1366), .dinb(n416), .dout(G330));
  jnot g1053(.din(n388), .dout(n1368));
  jnot g1054(.din(n396), .dout(n1369));
  jnot g1055(.din(n392), .dout(n1370));
  jor  g1056(.dina(n1337), .dinb(n1323), .dout(n1371));
  jand g1057(.dina(n1371), .dinb(n1370), .dout(n1372));
  jor  g1058(.dina(n1372), .dinb(n1369), .dout(n1373));
  jand g1059(.dina(n1373), .dinb(n405), .dout(n1374));
  jxor g1060(.dina(n1374), .dinb(n1368), .dout(G333));
  jxor g1061(.dina(n1372), .dinb(n1369), .dout(G336));
  jor  g1062(.dina(G416), .dinb(G414), .dout(n1377));
  jor  g1063(.dina(G408), .dinb(G404), .dout(n1378));
  jor  g1064(.dina(G410), .dinb(G406), .dout(n1379));
  jor  g1065(.dina(n1379), .dinb(G412), .dout(n1380));
  jor  g1066(.dina(n1380), .dinb(n1378), .dout(n1381));
  jor  g1067(.dina(n1381), .dinb(n1377), .dout(G418));
  jxor g1068(.dina(n705), .dinb(n425), .dout(G298));
  jand g1069(.dina(n703), .dinb(n438), .dout(n1384));
  jor  g1070(.dina(n1384), .dinb(n447), .dout(n1385));
  jxor g1071(.dina(n1385), .dinb(n429), .dout(G301));
  jand g1072(.dina(n1113), .dinb(G2239), .dout(n1387));
  jnot g1073(.din(n1387), .dout(n1388));
  jor  g1074(.dina(n703), .dinb(n445), .dout(n1389));
  jand g1075(.dina(n1389), .dinb(n1388), .dout(n1390));
  jxor g1076(.dina(n1390), .dinb(n433), .dout(G304));
  jxor g1077(.dina(n703), .dinb(n437), .dout(G307));
  jxor g1078(.dina(n680), .dinb(n575), .dout(G344));
  jor  g1079(.dina(n712), .dinb(G38), .dout(n1394));
  jor  g1080(.dina(n713), .dinb(n709), .dout(n1395));
  jand g1081(.dina(n1395), .dinb(n1394), .dout(n1396));
  jxor g1082(.dina(n1396), .dinb(n370), .dout(G422));
  jxor g1083(.dina(n709), .dinb(n363), .dout(G419));
  jand g1084(.dina(n680), .dinb(n580), .dout(n1399));
  jor  g1085(.dina(n1399), .dinb(n570), .dout(n1400));
  jxor g1086(.dina(n1400), .dinb(n573), .dout(G359));
  jnot g1087(.din(n577), .dout(n1402));
  jnot g1088(.din(n548), .dout(n1403));
  jnot g1089(.din(n566), .dout(n1404));
  jnot g1090(.din(n576), .dout(n1405));
  jand g1091(.dina(n1405), .dinb(n1404), .dout(n1406));
  jor  g1092(.dina(n1406), .dinb(n550), .dout(n1407));
  jand g1093(.dina(n1407), .dinb(n1403), .dout(n1408));
  jnot g1094(.din(n568), .dout(n1409));
  jand g1095(.dina(n1312), .dinb(n1409), .dout(n1410));
  jor  g1096(.dina(n1410), .dinb(n1408), .dout(n1411));
  jxor g1097(.dina(n1411), .dinb(n1402), .dout(G362));
  jand g1098(.dina(n680), .dinb(n576), .dout(n1413));
  jor  g1099(.dina(n1413), .dinb(n566), .dout(n1414));
  jxor g1100(.dina(n1414), .dinb(n578), .dout(G365));
  jand g1101(.dina(n680), .dinb(n575), .dout(n1416));
  jor  g1102(.dina(n1416), .dinb(n564), .dout(n1417));
  jxor g1103(.dina(n1417), .dinb(n574), .dout(G368));
  jxor g1104(.dina(n504), .dinb(n501), .dout(n1419));
  jxor g1105(.dina(n1419), .dinb(n698), .dout(G347));
  jand g1106(.dina(n694), .dinb(n1317), .dout(n1421));
  jxor g1107(.dina(n1421), .dinb(n1307), .dout(G350));
  jxor g1108(.dina(n524), .dinb(n518), .dout(n1423));
  jor  g1109(.dina(n1423), .dinb(n683), .dout(n1424));
  jand g1110(.dina(n1424), .dinb(n1316), .dout(G353));
  jxor g1111(.dina(n517), .dinb(n514), .dout(n1426));
  jxor g1112(.dina(n1426), .dinb(n682), .dout(G356));
  jxor g1113(.dina(n429), .dinb(n425), .dout(n1431));
  jor  g1114(.dina(n1388), .dinb(n444), .dout(n1432));
  jnot g1115(.din(n447), .dout(n1433));
  jor  g1116(.dina(n1433), .dinb(n1387), .dout(n1434));
  jand g1117(.dina(n1434), .dinb(n1432), .dout(n1435));
  jxor g1118(.dina(n1435), .dinb(n1431), .dout(n1436));
  jxor g1119(.dina(n449), .dinb(n433), .dout(n1437));
  jxor g1120(.dina(n1437), .dinb(n1436), .dout(n1438));
  jand g1121(.dina(n1438), .dinb(n1333), .dout(n1439));
  jxor g1122(.dina(n445), .dinb(n433), .dout(n1440));
  jnot g1123(.din(n1440), .dout(n1441));
  jand g1124(.dina(n1441), .dinb(n1433), .dout(n1442));
  jor  g1125(.dina(n437), .dinb(n444), .dout(n1443));
  jand g1126(.dina(n1443), .dinb(n1440), .dout(n1444));
  jor  g1127(.dina(n1444), .dinb(n1442), .dout(n1445));
  jxor g1128(.dina(n1431), .dinb(n450), .dout(n1446));
  jxor g1129(.dina(n1446), .dinb(n1445), .dout(n1447));
  jand g1130(.dina(n1447), .dinb(n703), .dout(n1448));
  jor  g1131(.dina(n1448), .dinb(n1439), .dout(n1449));
  jand g1132(.dina(n497), .dinb(n1340), .dout(n1450));
  jor  g1133(.dina(n1450), .dinb(n460), .dout(n1451));
  jxor g1134(.dina(n480), .dinb(n475), .dout(n1452));
  jand g1135(.dina(n1452), .dinb(n495), .dout(n1453));
  jnot g1136(.din(n1452), .dout(n1454));
  jand g1137(.dina(n1454), .dinb(n497), .dout(n1455));
  jor  g1138(.dina(n1455), .dinb(n1453), .dout(n1456));
  jnot g1139(.din(n479), .dout(n1457));
  jand g1140(.dina(n1457), .dinb(G2211), .dout(n1458));
  jnot g1141(.din(n1458), .dout(n1459));
  jor  g1142(.dina(n1459), .dinb(n491), .dout(n1460));
  jor  g1143(.dina(n1458), .dinb(n486), .dout(n1461));
  jand g1144(.dina(n1461), .dinb(n1460), .dout(n1462));
  jxor g1145(.dina(n1462), .dinb(n463), .dout(n1463));
  jxor g1146(.dina(n1463), .dinb(n1456), .dout(n1464));
  jxor g1147(.dina(n1464), .dinb(n1451), .dout(n1465));
  jand g1148(.dina(n1465), .dinb(n700), .dout(n1466));
  jand g1149(.dina(n496), .dinb(n1340), .dout(n1467));
  jor  g1150(.dina(n1467), .dinb(n460), .dout(n1468));
  jor  g1151(.dina(n487), .dinb(n491), .dout(n1469));
  jand g1152(.dina(n1469), .dinb(n489), .dout(n1470));
  jxor g1153(.dina(n1470), .dinb(n463), .dout(n1471));
  jxor g1154(.dina(n1471), .dinb(n495), .dout(n1472));
  jxor g1155(.dina(n1472), .dinb(n1452), .dout(n1473));
  jxor g1156(.dina(n1473), .dinb(n1468), .dout(n1474));
  jand g1157(.dina(n1474), .dinb(n1321), .dout(n1475));
  jor  g1158(.dina(n1475), .dinb(n1466), .dout(n1476));
  jxor g1159(.dina(n470), .dinb(n464), .dout(n1477));
  jxor g1160(.dina(n1477), .dinb(n1476), .dout(n1478));
  jxor g1161(.dina(n1478), .dinb(n1449), .dout(G321));
  jxor g1162(.dina(n416), .dinb(n388), .dout(n1480));
  jxor g1163(.dina(n411), .dinb(n377), .dout(n1481));
  jand g1164(.dina(n407), .dinb(n1370), .dout(n1482));
  jand g1165(.dina(n409), .dinb(n392), .dout(n1483));
  jor  g1166(.dina(n1483), .dinb(n1482), .dout(n1484));
  jnot g1167(.din(n397), .dout(n1485));
  jand g1168(.dina(n1485), .dinb(n405), .dout(n1486));
  jxor g1169(.dina(n414), .dinb(n396), .dout(n1487));
  jxor g1170(.dina(n1487), .dinb(n1486), .dout(n1488));
  jxor g1171(.dina(n1488), .dinb(n1484), .dout(n1489));
  jxor g1172(.dina(n1489), .dinb(n1481), .dout(n1490));
  jor  g1173(.dina(n1490), .dinb(n707), .dout(n1491));
  jor  g1174(.dina(n391), .dinb(n389), .dout(n1492));
  jor  g1175(.dina(n395), .dinb(n393), .dout(n1493));
  jand g1176(.dina(n1493), .dinb(n1492), .dout(n1494));
  jnot g1177(.din(n1492), .dout(n1495));
  jand g1178(.dina(n1486), .dinb(n1495), .dout(n1496));
  jor  g1179(.dina(n1496), .dinb(n1494), .dout(n1497));
  jxor g1180(.dina(n396), .dinb(n377), .dout(n1498));
  jxor g1181(.dina(n1498), .dinb(n1364), .dout(n1499));
  jxor g1182(.dina(n1499), .dinb(n1497), .dout(n1500));
  jxor g1183(.dina(n1500), .dinb(n414), .dout(n1501));
  jxor g1184(.dina(n1501), .dinb(n1359), .dout(n1502));
  jor  g1185(.dina(n1502), .dinb(n1337), .dout(n1503));
  jand g1186(.dina(n1503), .dinb(n1491), .dout(n1504));
  jxor g1187(.dina(n1504), .dinb(n1480), .dout(n1505));
  jand g1188(.dina(n362), .dinb(G38), .dout(n1506));
  jnot g1189(.din(n364), .dout(n1507));
  jor  g1190(.dina(n1507), .dinb(n1506), .dout(n1508));
  jnot g1191(.din(n1506), .dout(n1509));
  jor  g1192(.dina(n1509), .dinb(G1496), .dout(n1510));
  jand g1193(.dina(n1510), .dinb(n1508), .dout(n1511));
  jand g1194(.dina(n1511), .dinb(n413), .dout(n1512));
  jnot g1195(.din(n413), .dout(n1513));
  jand g1196(.dina(n712), .dinb(n361), .dout(n1514));
  jor  g1197(.dina(n364), .dinb(n1514), .dout(n1515));
  jor  g1198(.dina(n369), .dinb(G1492), .dout(n1516));
  jand g1199(.dina(n1516), .dinb(n1515), .dout(n1517));
  jand g1200(.dina(n1517), .dinb(n1513), .dout(n1518));
  jor  g1201(.dina(n1518), .dinb(n1512), .dout(n1519));
  jor  g1202(.dina(n1519), .dinb(n707), .dout(n1520));
  jnot g1203(.din(n419), .dout(n1521));
  jand g1204(.dina(n1518), .dinb(n1521), .dout(n1522));
  jand g1205(.dina(n1511), .dinb(n420), .dout(n1523));
  jor  g1206(.dina(n1523), .dinb(n1522), .dout(n1524));
  jor  g1207(.dina(n1524), .dinb(n1337), .dout(n1525));
  jand g1208(.dina(n1525), .dinb(n1520), .dout(n1526));
  jxor g1209(.dina(n1526), .dinb(n1505), .dout(G338));
  jor  g1210(.dina(n693), .dinb(n687), .dout(n1528));
  jand g1211(.dina(n1528), .dinb(n695), .dout(n1529));
  jor  g1212(.dina(n1529), .dinb(n513), .dout(n1530));
  jxor g1213(.dina(n1419), .dinb(n1308), .dout(n1531));
  jxor g1214(.dina(n1531), .dinb(n526), .dout(n1532));
  jxor g1215(.dina(n1532), .dinb(n1530), .dout(n1533));
  jand g1216(.dina(n1533), .dinb(n1309), .dout(n1534));
  jand g1217(.dina(n1534), .dinb(n1310), .dout(n1535));
  jand g1218(.dina(n1426), .dinb(n524), .dout(n1536));
  jnot g1219(.din(n1536), .dout(n1537));
  jor  g1220(.dina(n1537), .dinb(n690), .dout(n1538));
  jor  g1221(.dina(n1536), .dinb(n1529), .dout(n1539));
  jand g1222(.dina(n1539), .dinb(n1538), .dout(n1540));
  jxor g1223(.dina(n518), .dinb(n513), .dout(n1541));
  jxor g1224(.dina(n1541), .dinb(n1531), .dout(n1542));
  jxor g1225(.dina(n1542), .dinb(n1540), .dout(n1543));
  jor  g1226(.dina(n581), .dinb(n572), .dout(n1544));
  jand g1227(.dina(n1544), .dinb(n1543), .dout(n1545));
  jor  g1228(.dina(n1545), .dinb(n1535), .dout(n1546));
  jand g1229(.dina(n1546), .dinb(n680), .dout(n1547));
  jand g1230(.dina(n1543), .dinb(n572), .dout(n1548));
  jor  g1231(.dina(n1548), .dinb(n1534), .dout(n1549));
  jand g1232(.dina(n1549), .dinb(n1312), .dout(n1550));
  jor  g1233(.dina(n1550), .dinb(n1547), .dout(n1551));
  jxor g1234(.dina(n578), .dinb(n1402), .dout(n1552));
  jnot g1235(.din(n563), .dout(n1553));
  jand g1236(.dina(n1553), .dinb(G4394), .dout(n1554));
  jnot g1237(.din(n1554), .dout(n1555));
  jand g1238(.dina(n1555), .dinb(n558), .dout(n1556));
  jand g1239(.dina(n1554), .dinb(n556), .dout(n1557));
  jor  g1240(.dina(n1557), .dinb(n1556), .dout(n1558));
  jxor g1241(.dina(n1558), .dinb(n573), .dout(n1559));
  jxor g1242(.dina(n1559), .dinb(n1408), .dout(n1560));
  jnot g1243(.din(n570), .dout(n1561));
  jxor g1244(.dina(n575), .dinb(n574), .dout(n1562));
  jnot g1245(.din(n1562), .dout(n1563));
  jor  g1246(.dina(n1563), .dinb(n1561), .dout(n1564));
  jor  g1247(.dina(n1562), .dinb(n570), .dout(n1565));
  jor  g1248(.dina(n1565), .dinb(n580), .dout(n1566));
  jand g1249(.dina(n1566), .dinb(n1564), .dout(n1567));
  jxor g1250(.dina(n1567), .dinb(n1560), .dout(n1568));
  jor  g1251(.dina(n1568), .dinb(n1312), .dout(n1569));
  jxor g1252(.dina(n1562), .dinb(n570), .dout(n1570));
  jnot g1253(.din(n565), .dout(n1571));
  jor  g1254(.dina(n564), .dinb(n556), .dout(n1572));
  jand g1255(.dina(n1572), .dinb(n1571), .dout(n1573));
  jxor g1256(.dina(n1573), .dinb(n573), .dout(n1574));
  jxor g1257(.dina(n1574), .dinb(n568), .dout(n1575));
  jxor g1258(.dina(n1575), .dinb(n1570), .dout(n1576));
  jor  g1259(.dina(n1576), .dinb(n680), .dout(n1577));
  jand g1260(.dina(n1577), .dinb(n1569), .dout(n1578));
  jxor g1261(.dina(n1578), .dinb(n1552), .dout(n1579));
  jxor g1262(.dina(n1579), .dinb(n1551), .dout(G370));
  jxor g1263(.dina(n1084), .dinb(n1108), .dout(n1581));
  jxor g1264(.dina(n1581), .dinb(n1105), .dout(n1582));
  jand g1265(.dina(n616), .dinb(n609), .dout(n1583));
  jand g1266(.dina(n615), .dinb(n610), .dout(n1584));
  jor  g1267(.dina(n1584), .dinb(n1583), .dout(n1585));
  jxor g1268(.dina(n1585), .dinb(n1582), .dout(n1586));
  jand g1269(.dina(n1586), .dinb(n1092), .dout(n1587));
  jand g1270(.dina(n1587), .dinb(n1086), .dout(n1588));
  jnot g1271(.din(n598), .dout(n1589));
  jand g1272(.dina(n1589), .dinb(G3737), .dout(n1590));
  jand g1273(.dina(n1106), .dinb(n1590), .dout(n1591));
  jand g1274(.dina(n613), .dinb(n612), .dout(n1592));
  jor  g1275(.dina(n1592), .dinb(n1591), .dout(n1593));
  jor  g1276(.dina(n1593), .dinb(n605), .dout(n1594));
  jxor g1277(.dina(n1084), .dinb(n594), .dout(n1595));
  jxor g1278(.dina(n1595), .dinb(n1594), .dout(n1596));
  jxor g1279(.dina(n1596), .dinb(n619), .dout(n1597));
  jand g1280(.dina(n1597), .dinb(n674), .dout(n1598));
  jor  g1281(.dina(n1598), .dinb(n1094), .dout(n1599));
  jor  g1282(.dina(n1599), .dinb(n1588), .dout(n1600));
  jand g1283(.dina(n1597), .dinb(n673), .dout(n1601));
  jor  g1284(.dina(n1601), .dinb(n1587), .dout(n1602));
  jor  g1285(.dina(n1602), .dinb(G4526), .dout(n1603));
  jand g1286(.dina(n1603), .dinb(n1600), .dout(n1604));
  jxor g1287(.dina(n642), .dinb(n359), .dout(n1605));
  jxor g1288(.dina(n1605), .dinb(n1067), .dout(n1606));
  jxor g1289(.dina(n1606), .dinb(n1069), .dout(n1607));
  jnot g1290(.din(n1607), .dout(n1608));
  jxor g1291(.dina(n626), .dinb(n354), .dout(n1609));
  jxor g1292(.dina(n1609), .dinb(n671), .dout(n1610));
  jor  g1293(.dina(n1610), .dinb(n1608), .dout(n1611));
  jnot g1294(.din(n1610), .dout(n1612));
  jor  g1295(.dina(n1612), .dinb(n1607), .dout(n1613));
  jand g1296(.dina(n1613), .dinb(n1094), .dout(n1614));
  jand g1297(.dina(n1614), .dinb(n1611), .dout(n1615));
  jand g1298(.dina(n1067), .dinb(n357), .dout(n1616));
  jand g1299(.dina(n661), .dinb(n358), .dout(n1617));
  jor  g1300(.dina(n1617), .dinb(n1616), .dout(n1618));
  jxor g1301(.dina(n1618), .dinb(n626), .dout(n1619));
  jxor g1302(.dina(n1619), .dinb(n1070), .dout(n1620));
  jnot g1303(.din(n1620), .dout(n1621));
  jnot g1304(.din(n645), .dout(n1622));
  jand g1305(.dina(n1090), .dinb(n1622), .dout(n1623));
  jxor g1306(.dina(n1623), .dinb(n1605), .dout(n1624));
  jnot g1307(.din(n1624), .dout(n1625));
  jor  g1308(.dina(n1625), .dinb(n1621), .dout(n1626));
  jor  g1309(.dina(n1624), .dinb(n1620), .dout(n1627));
  jand g1310(.dina(n1627), .dinb(G4526), .dout(n1628));
  jand g1311(.dina(n1628), .dinb(n1626), .dout(n1629));
  jor  g1312(.dina(n1629), .dinb(n1615), .dout(n1630));
  jxor g1313(.dina(n636), .dinb(n631), .dout(n1631));
  jxor g1314(.dina(n1631), .dinb(n1630), .dout(n1632));
  jxor g1315(.dina(n1632), .dinb(n1604), .dout(G399));
  jdff  g1316(.din(G1), .dout(G2));
  jdff  g1317(.din(G1), .dout(G3));
  jdff  g1318(.din(G1459), .dout(G450));
  jdff  g1319(.din(G1469), .dout(G448));
  jdff  g1320(.din(G1480), .dout(G444));
  jdff  g1321(.din(G1486), .dout(G442));
  jdff  g1322(.din(G1492), .dout(G440));
  jdff  g1323(.din(G1496), .dout(G438));
  jdff  g1324(.din(G2208), .dout(G496));
  jdff  g1325(.din(G2218), .dout(G494));
  jdff  g1326(.din(G2224), .dout(G492));
  jdff  g1327(.din(G2230), .dout(G490));
  jdff  g1328(.din(G2236), .dout(G488));
  jdff  g1329(.din(G2239), .dout(G486));
  jdff  g1330(.din(G2247), .dout(G484));
  jdff  g1331(.din(G2253), .dout(G482));
  jdff  g1332(.din(G2256), .dout(G480));
  jdff  g1333(.din(G3698), .dout(G560));
  jdff  g1334(.din(G3701), .dout(G542));
  jdff  g1335(.din(G3705), .dout(G558));
  jdff  g1336(.din(G3711), .dout(G556));
  jdff  g1337(.din(G3717), .dout(G554));
  jdff  g1338(.din(G3723), .dout(G552));
  jdff  g1339(.din(G3729), .dout(G550));
  jdff  g1340(.din(G3737), .dout(G548));
  jdff  g1341(.din(G3743), .dout(G546));
  jdff  g1342(.din(G3749), .dout(G544));
  jdff  g1343(.din(G4393), .dout(G540));
  jdff  g1344(.din(G4400), .dout(G538));
  jdff  g1345(.din(G4405), .dout(G536));
  jdff  g1346(.din(G4410), .dout(G534));
  jdff  g1347(.din(G4415), .dout(G532));
  jdff  g1348(.din(G4420), .dout(G530));
  jdff  g1349(.din(G4427), .dout(G528));
  jdff  g1350(.din(G4432), .dout(G526));
  jdff  g1351(.din(G4437), .dout(G524));
  jdff  g1352(.din(G1462), .dout(G436));
  jdff  g1353(.din(G2211), .dout(G478));
  jdff  g1354(.din(G4394), .dout(G522));
  jdff  g1355(.din(G1), .dout(G432));
  jdff  g1356(.din(G106), .dout(G446));
  jnot g1357(.din(G15), .dout(G286));
  jor  g1358(.dina(n345), .dinb(G5), .dout(G289));
  jnot g1359(.din(G15), .dout(G341));
  jor  g1360(.dina(n349), .dinb(n347), .dout(G281));
  jdff  g1361(.din(G1), .dout(G453));
  jand g1362(.dina(n1059), .dinb(n718), .dout(G264));
  jor  g1363(.dina(n715), .dinb(n711), .dout(G270));
  jand g1364(.dina(n1059), .dinb(n718), .dout(G249));
  jor  g1365(.dina(n715), .dinb(n711), .dout(G276));
  jor  g1366(.dina(n715), .dinb(n711), .dout(G273));
  jxor g1367(.dina(n1396), .dinb(n370), .dout(G469));
  jxor g1368(.dina(n709), .dinb(n363), .dout(G471));
endmodule


