module gf_c3540(G1698, G330, G326, G343, G317, G311, G303, G294, G2897, G274, G250, G244, G238, G232, G322, G226, G223, G270, G200, G257, G77, G20, G125, G116, G283, G143, G45, G190, G68, G1, G58, G132, G33, G150, G87, G128, G97, G107, G124, G329, G264, G222, G50, G137, G159, G41, G169, G13, G179, G213, G409, G407, G381, G375, G378, G393, G353, G361, G390, G396, G351, G372, G384, G405, G358, G355, G369, G399, G364, G367, G402, G387);
    input G1698, G330, G326, G343, G317, G311, G303, G294, G2897, G274, G250, G244, G238, G232, G322, G226, G223, G270, G200, G257, G77, G20, G125, G116, G283, G143, G45, G190, G68, G1, G58, G132, G33, G150, G87, G128, G97, G107, G124, G329, G264, G222, G50, G137, G159, G41, G169, G13, G179, G213;
    output G409, G407, G381, G375, G378, G393, G353, G361, G390, G396, G351, G372, G384, G405, G358, G355, G369, G399, G364, G367, G402, G387;
    wire n74;
    wire n77;
    wire n80;
    wire n83;
    wire n87;
    wire n91;
    wire n95;
    wire n98;
    wire n101;
    wire n104;
    wire n108;
    wire n112;
    wire n115;
    wire n118;
    wire n121;
    wire n125;
    wire n129;
    wire n132;
    wire n136;
    wire n140;
    wire n144;
    wire n148;
    wire n151;
    wire n155;
    wire n158;
    wire n162;
    wire n166;
    wire n169;
    wire n173;
    wire n177;
    wire n181;
    wire n184;
    wire n188;
    wire n191;
    wire n194;
    wire n198;
    wire n202;
    wire n206;
    wire n210;
    wire n214;
    wire n217;
    wire n221;
    wire n225;
    wire n229;
    wire n233;
    wire n236;
    wire n240;
    wire n243;
    wire n247;
    wire n251;
    wire n255;
    wire n259;
    wire n263;
    wire n267;
    wire n271;
    wire n274;
    wire n278;
    wire n282;
    wire n286;
    wire n290;
    wire n294;
    wire n298;
    wire n302;
    wire n306;
    wire n310;
    wire n314;
    wire n318;
    wire n322;
    wire n326;
    wire n330;
    wire n333;
    wire n337;
    wire n341;
    wire n345;
    wire n349;
    wire n353;
    wire n356;
    wire n360;
    wire n364;
    wire n367;
    wire n371;
    wire n374;
    wire n378;
    wire n382;
    wire n386;
    wire n390;
    wire n394;
    wire n398;
    wire n402;
    wire n406;
    wire n409;
    wire n412;
    wire n416;
    wire n420;
    wire n423;
    wire n427;
    wire n431;
    wire n435;
    wire n439;
    wire n442;
    wire n446;
    wire n450;
    wire n454;
    wire n458;
    wire n461;
    wire n465;
    wire n469;
    wire n473;
    wire n477;
    wire n481;
    wire n484;
    wire n488;
    wire n492;
    wire n496;
    wire n500;
    wire n504;
    wire n507;
    wire n510;
    wire n514;
    wire n518;
    wire n522;
    wire n526;
    wire n529;
    wire n533;
    wire n537;
    wire n541;
    wire n545;
    wire n548;
    wire n552;
    wire n556;
    wire n560;
    wire n564;
    wire n567;
    wire n571;
    wire n575;
    wire n579;
    wire n582;
    wire n586;
    wire n590;
    wire n594;
    wire n598;
    wire n602;
    wire n606;
    wire n610;
    wire n614;
    wire n618;
    wire n622;
    wire n626;
    wire n630;
    wire n634;
    wire n638;
    wire n642;
    wire n646;
    wire n649;
    wire n652;
    wire n655;
    wire n659;
    wire n663;
    wire n666;
    wire n670;
    wire n674;
    wire n678;
    wire n682;
    wire n686;
    wire n690;
    wire n694;
    wire n698;
    wire n702;
    wire n706;
    wire n710;
    wire n714;
    wire n718;
    wire n721;
    wire n724;
    wire n728;
    wire n732;
    wire n736;
    wire n740;
    wire n744;
    wire n748;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n779;
    wire n783;
    wire n786;
    wire n790;
    wire n793;
    wire n797;
    wire n801;
    wire n805;
    wire n809;
    wire n813;
    wire n817;
    wire n820;
    wire n824;
    wire n828;
    wire n831;
    wire n835;
    wire n839;
    wire n842;
    wire n846;
    wire n850;
    wire n854;
    wire n858;
    wire n862;
    wire n866;
    wire n870;
    wire n873;
    wire n876;
    wire n880;
    wire n884;
    wire n888;
    wire n892;
    wire n896;
    wire n900;
    wire n904;
    wire n908;
    wire n912;
    wire n916;
    wire n920;
    wire n924;
    wire n928;
    wire n931;
    wire n935;
    wire n939;
    wire n942;
    wire n946;
    wire n950;
    wire n954;
    wire n958;
    wire n962;
    wire n966;
    wire n970;
    wire n974;
    wire n977;
    wire n981;
    wire n985;
    wire n988;
    wire n992;
    wire n996;
    wire n1000;
    wire n1004;
    wire n1008;
    wire n1012;
    wire n1016;
    wire n1020;
    wire n1024;
    wire n1028;
    wire n1032;
    wire n1036;
    wire n1040;
    wire n1044;
    wire n1048;
    wire n1052;
    wire n1056;
    wire n1060;
    wire n1064;
    wire n1068;
    wire n1071;
    wire n1074;
    wire n1078;
    wire n1082;
    wire n1086;
    wire n1090;
    wire n1094;
    wire n1097;
    wire n1101;
    wire n1105;
    wire n1109;
    wire n1113;
    wire n1117;
    wire n1121;
    wire n1125;
    wire n1129;
    wire n1133;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1147;
    wire n1151;
    wire n1154;
    wire n1158;
    wire n1162;
    wire n1166;
    wire n1170;
    wire n1174;
    wire n1177;
    wire n1181;
    wire n1185;
    wire n1189;
    wire n1193;
    wire n1196;
    wire n1200;
    wire n1204;
    wire n1208;
    wire n1212;
    wire n1216;
    wire n1220;
    wire n1224;
    wire n1227;
    wire n1231;
    wire n1234;
    wire n1238;
    wire n1242;
    wire n1246;
    wire n1250;
    wire n1254;
    wire n1257;
    wire n1261;
    wire n1265;
    wire n1269;
    wire n1272;
    wire n1276;
    wire n1279;
    wire n1283;
    wire n1287;
    wire n1291;
    wire n1295;
    wire n1298;
    wire n1302;
    wire n1306;
    wire n1310;
    wire n1314;
    wire n1318;
    wire n1322;
    wire n1326;
    wire n1330;
    wire n1334;
    wire n1337;
    wire n1341;
    wire n1345;
    wire n1349;
    wire n1353;
    wire n1357;
    wire n1361;
    wire n1365;
    wire n1369;
    wire n1373;
    wire n1377;
    wire n1381;
    wire n1385;
    wire n1389;
    wire n1393;
    wire n1397;
    wire n1401;
    wire n1405;
    wire n1409;
    wire n1413;
    wire n1416;
    wire n1420;
    wire n1424;
    wire n1428;
    wire n1431;
    wire n1435;
    wire n1438;
    wire n1441;
    wire n1444;
    wire n1448;
    wire n1452;
    wire n1456;
    wire n1460;
    wire n1464;
    wire n1468;
    wire n1472;
    wire n1476;
    wire n1480;
    wire n1483;
    wire n1487;
    wire n1491;
    wire n1495;
    wire n1498;
    wire n1502;
    wire n1506;
    wire n1510;
    wire n1513;
    wire n1516;
    wire n1520;
    wire n1523;
    wire n1527;
    wire n1531;
    wire n1535;
    wire n1538;
    wire n1542;
    wire n1546;
    wire n1550;
    wire n1554;
    wire n1558;
    wire n1562;
    wire n1566;
    wire n1570;
    wire n1573;
    wire n1576;
    wire n1580;
    wire n1584;
    wire n1588;
    wire n1592;
    wire n1596;
    wire n1600;
    wire n1604;
    wire n1608;
    wire n1612;
    wire n1616;
    wire n1620;
    wire n1624;
    wire n1628;
    wire n1632;
    wire n1635;
    wire n1639;
    wire n1642;
    wire n1645;
    wire n1649;
    wire n1653;
    wire n1657;
    wire n1661;
    wire n1664;
    wire n1668;
    wire n1672;
    wire n1676;
    wire n1679;
    wire n1683;
    wire n1686;
    wire n1690;
    wire n1694;
    wire n1698;
    wire n1702;
    wire n1706;
    wire n1710;
    wire n1714;
    wire n1717;
    wire n1721;
    wire n1724;
    wire n1728;
    wire n1732;
    wire n1736;
    wire n1740;
    wire n1744;
    wire n1748;
    wire n1752;
    wire n1755;
    wire n1759;
    wire n1762;
    wire n1766;
    wire n1770;
    wire n1774;
    wire n1777;
    wire n1781;
    wire n1785;
    wire n1789;
    wire n1793;
    wire n1796;
    wire n1800;
    wire n1804;
    wire n1808;
    wire n1811;
    wire n1815;
    wire n1819;
    wire n1823;
    wire n1827;
    wire n1830;
    wire n1834;
    wire n1838;
    wire n1842;
    wire n1846;
    wire n1850;
    wire n1854;
    wire n1858;
    wire n1862;
    wire n1866;
    wire n1870;
    wire n1874;
    wire n1878;
    wire n1882;
    wire n1886;
    wire n1890;
    wire n1894;
    wire n1897;
    wire n1900;
    wire n1904;
    wire n1907;
    wire n1910;
    wire n1913;
    wire n1917;
    wire n1921;
    wire n1925;
    wire n1929;
    wire n1933;
    wire n1936;
    wire n1940;
    wire n1944;
    wire n1948;
    wire n1952;
    wire n1956;
    wire n1959;
    wire n1962;
    wire n1965;
    wire n1969;
    wire n1973;
    wire n1977;
    wire n1981;
    wire n1985;
    wire n1989;
    wire n1993;
    wire n1997;
    wire n2001;
    wire n2005;
    wire n2009;
    wire n2013;
    wire n2017;
    wire n2020;
    wire n2024;
    wire n2028;
    wire n2031;
    wire n2035;
    wire n2039;
    wire n2043;
    wire n2047;
    wire n2051;
    wire n2055;
    wire n2059;
    wire n2063;
    wire n2067;
    wire n2071;
    wire n2074;
    wire n2078;
    wire n2082;
    wire n2085;
    wire n2089;
    wire n2092;
    wire n2096;
    wire n2100;
    wire n2104;
    wire n2108;
    wire n2112;
    wire n2116;
    wire n2120;
    wire n2124;
    wire n2127;
    wire n2131;
    wire n2134;
    wire n2138;
    wire n2142;
    wire n2146;
    wire n2150;
    wire n2153;
    wire n2157;
    wire n2161;
    wire n2164;
    wire n2168;
    wire n2171;
    wire n2175;
    wire n2178;
    wire n2182;
    wire n2186;
    wire n2190;
    wire n2193;
    wire n2197;
    wire n2201;
    wire n2205;
    wire n2208;
    wire n2212;
    wire n2216;
    wire n2220;
    wire n2224;
    wire n2228;
    wire n2232;
    wire n2236;
    wire n2240;
    wire n2243;
    wire n2247;
    wire n2251;
    wire n2255;
    wire n2259;
    wire n2263;
    wire n2267;
    wire n2271;
    wire n2275;
    wire n2279;
    wire n2283;
    wire n2287;
    wire n2291;
    wire n2295;
    wire n2298;
    wire n2302;
    wire n2305;
    wire n2309;
    wire n2313;
    wire n2317;
    wire n2321;
    wire n2325;
    wire n2329;
    wire n2333;
    wire n2337;
    wire n2341;
    wire n2345;
    wire n2349;
    wire n2353;
    wire n2357;
    wire n2361;
    wire n2365;
    wire n2369;
    wire n2373;
    wire n2377;
    wire n2381;
    wire n2384;
    wire n2388;
    wire n2392;
    wire n2396;
    wire n2400;
    wire n2403;
    wire n2407;
    wire n2411;
    wire n2414;
    wire n2418;
    wire n2421;
    wire n2425;
    wire n2429;
    wire n2433;
    wire n2437;
    wire n2441;
    wire n2445;
    wire n2448;
    wire n2452;
    wire n2456;
    wire n2460;
    wire n2464;
    wire n2468;
    wire n2472;
    wire n2475;
    wire n2479;
    wire n2482;
    wire n2486;
    wire n2490;
    wire n2494;
    wire n2498;
    wire n2502;
    wire n2506;
    wire n2510;
    wire n2514;
    wire n2518;
    wire n2522;
    wire n2526;
    wire n2530;
    wire n2534;
    wire n2538;
    wire n2542;
    wire n2546;
    wire n2550;
    wire n2554;
    wire n2558;
    wire n2562;
    wire n2566;
    wire n2570;
    wire n2574;
    wire n2578;
    wire n2582;
    wire n2586;
    wire n2590;
    wire n2594;
    wire n2598;
    wire n2602;
    wire n2606;
    wire n2610;
    wire n2614;
    wire n2617;
    wire n2621;
    wire n2625;
    wire n2628;
    wire n2632;
    wire n2636;
    wire n2640;
    wire n2643;
    wire n2647;
    wire n2651;
    wire n2655;
    wire n2658;
    wire n2662;
    wire n2666;
    wire n2670;
    wire n2674;
    wire n2678;
    wire n2682;
    wire n2686;
    wire n2690;
    wire n2693;
    wire n2696;
    wire n2700;
    wire n2703;
    wire n2707;
    wire n2711;
    wire n2715;
    wire n2718;
    wire n2722;
    wire n2725;
    wire n2729;
    wire n2733;
    wire n2736;
    wire n2740;
    wire n2744;
    wire n2748;
    wire n2752;
    wire n2756;
    wire n2760;
    wire n2764;
    wire n2768;
    wire n2772;
    wire n2776;
    wire n2780;
    wire n2784;
    wire n2788;
    wire n2792;
    wire n2796;
    wire n2800;
    wire n2804;
    wire n2808;
    wire n2812;
    wire n2816;
    wire n2820;
    wire n2824;
    wire n2828;
    wire n2832;
    wire n2836;
    wire n2840;
    wire n2844;
    wire n2847;
    wire n2851;
    wire n2854;
    wire n2858;
    wire n2862;
    wire n2866;
    wire n2870;
    wire n2874;
    wire n2878;
    wire n2882;
    wire n2886;
    wire n2890;
    wire n2894;
    wire n2898;
    wire n2902;
    wire n2906;
    wire n2910;
    wire n2914;
    wire n2918;
    wire n2922;
    wire n2926;
    wire n2930;
    wire n2934;
    wire n2938;
    wire n2942;
    wire n2946;
    wire n2950;
    wire n2954;
    wire n2958;
    wire n2962;
    wire n2966;
    wire n2970;
    wire n2974;
    wire n2978;
    wire n2982;
    wire n2986;
    wire n2990;
    wire n2994;
    wire n2998;
    wire n3002;
    wire n3006;
    wire n3010;
    wire n3014;
    wire n3017;
    wire n3021;
    wire n3025;
    wire n3028;
    wire n3032;
    wire n3036;
    wire n3040;
    wire n3044;
    wire n3048;
    wire n3052;
    wire n3056;
    wire n3060;
    wire n3064;
    wire n3068;
    wire n3071;
    wire n3075;
    wire n3079;
    wire n3083;
    wire n3086;
    wire n3090;
    wire n3094;
    wire n3098;
    wire n3102;
    wire n3106;
    wire n3110;
    wire n3114;
    wire n3118;
    wire n3121;
    wire n3125;
    wire n3129;
    wire n3133;
    wire n3137;
    wire n3141;
    wire n3145;
    wire n3149;
    wire n3153;
    wire n3157;
    wire n3161;
    wire n3165;
    wire n3169;
    wire n3172;
    wire n3176;
    wire n3179;
    wire n3183;
    wire n3186;
    wire n3190;
    wire n3194;
    wire n3198;
    wire n3202;
    wire n3206;
    wire n3210;
    wire n3213;
    wire n3217;
    wire n3221;
    wire n3224;
    wire n3228;
    wire n3232;
    wire n3236;
    wire n3240;
    wire n3244;
    wire n3248;
    wire n3252;
    wire n3256;
    wire n3260;
    wire n3264;
    wire n3268;
    wire n3272;
    wire n3276;
    wire n3280;
    wire n3284;
    wire n3288;
    wire n3292;
    wire n3296;
    wire n3300;
    wire n3303;
    wire n3306;
    wire n3310;
    wire n3313;
    wire n3317;
    wire n3321;
    wire n3325;
    wire n3329;
    wire n3332;
    wire n3336;
    wire n3340;
    wire n3344;
    wire n3348;
    wire n3352;
    wire n3356;
    wire n3360;
    wire n3364;
    wire n3368;
    wire n3372;
    wire n3375;
    wire n3379;
    wire n3382;
    wire n3385;
    wire n3388;
    wire n3392;
    wire n3396;
    wire n3400;
    wire n3404;
    wire n3407;
    wire n3411;
    wire n3415;
    wire n3419;
    wire n3423;
    wire n3427;
    wire n3431;
    wire n3435;
    wire n3439;
    wire n3443;
    wire n3447;
    wire n3451;
    wire n3455;
    wire n3459;
    wire n3463;
    wire n3467;
    wire n3471;
    wire n3475;
    wire n3479;
    wire n3483;
    wire n3487;
    wire n3491;
    wire n3495;
    wire n3499;
    wire n3503;
    wire n3507;
    wire n3511;
    wire n3515;
    wire n3519;
    wire n3523;
    wire n3527;
    wire n3531;
    wire n3535;
    wire n3539;
    wire n3543;
    wire n3547;
    wire n3551;
    wire n3555;
    wire n3559;
    wire n3563;
    wire n3566;
    wire n3570;
    wire n3574;
    wire n3577;
    wire n3581;
    wire n3584;
    wire n3588;
    wire n3592;
    wire n3596;
    wire n3600;
    wire n3604;
    wire n3608;
    wire n3612;
    wire n3616;
    wire n3620;
    wire n3624;
    wire n3628;
    wire n3632;
    wire n3636;
    wire n3640;
    wire n3644;
    wire n3648;
    wire n3652;
    wire n3656;
    wire n3660;
    wire n3664;
    wire n3668;
    wire n3672;
    wire n3676;
    wire n3680;
    wire n3684;
    wire n3688;
    wire n3692;
    wire n3696;
    wire n3700;
    wire n3704;
    wire n3708;
    wire n3712;
    wire n3715;
    wire n3719;
    wire n3723;
    wire n3727;
    wire n3730;
    wire n3734;
    wire n3738;
    wire n3741;
    wire n3745;
    wire n3748;
    wire n3752;
    wire n3756;
    wire n3760;
    wire n3764;
    wire n3768;
    wire n3772;
    wire n3776;
    wire n3780;
    wire n3784;
    wire n3788;
    wire n3792;
    wire n3796;
    wire n3800;
    wire n3804;
    wire n3807;
    wire n3810;
    wire n3814;
    wire n3818;
    wire n3822;
    wire n3826;
    wire n3830;
    wire n3833;
    wire n3837;
    wire n3841;
    wire n3845;
    wire n3849;
    wire n3853;
    wire n3857;
    wire n3861;
    wire n3865;
    wire n3869;
    wire n3873;
    wire n3877;
    wire n3881;
    wire n3885;
    wire n3888;
    wire n3892;
    wire n3896;
    wire n3900;
    wire n3904;
    wire n3908;
    wire n3912;
    wire n3916;
    wire n3920;
    wire n3924;
    wire n3928;
    wire n3932;
    wire n3936;
    wire n3940;
    wire n3944;
    wire n3948;
    wire n3952;
    wire n3956;
    wire n3960;
    wire n3964;
    wire n3968;
    wire n3972;
    wire n3975;
    wire n3979;
    wire n3982;
    wire n3986;
    wire n3990;
    wire n3994;
    wire n3998;
    wire n4002;
    wire n4006;
    wire n4010;
    wire n4014;
    wire n4017;
    wire n4021;
    wire n4025;
    wire n4028;
    wire n4032;
    wire n4036;
    wire n4040;
    wire n4044;
    wire n4047;
    wire n4051;
    wire n4055;
    wire n4059;
    wire n4062;
    wire n4066;
    wire n4069;
    wire n4073;
    wire n4076;
    wire n4080;
    wire n4084;
    wire n4088;
    wire n4092;
    wire n4096;
    wire n4100;
    wire n4104;
    wire n4108;
    wire n4112;
    wire n4116;
    wire n4120;
    wire n4124;
    wire n4128;
    wire n4132;
    wire n4136;
    wire n4140;
    wire n4144;
    wire n4148;
    wire n4152;
    wire n4156;
    wire n4160;
    wire n4164;
    wire n4168;
    wire n4172;
    wire n4176;
    wire n4180;
    wire n4184;
    wire n4188;
    wire n4192;
    wire n4196;
    wire n4200;
    wire n4204;
    wire n4207;
    wire n4211;
    wire n4215;
    wire n4219;
    wire n4222;
    wire n4226;
    wire n4229;
    wire n4233;
    wire n4237;
    wire n4241;
    wire n4244;
    wire n4248;
    wire n4252;
    wire n4256;
    wire n4259;
    wire n4263;
    wire n4267;
    wire n4271;
    wire n4275;
    wire n4278;
    wire n4281;
    wire n4285;
    wire n4288;
    wire n4292;
    wire n4300;
    wire n4304;
    wire n4308;
    wire n4312;
    wire n4316;
    wire n4320;
    wire n4324;
    wire n4327;
    wire n4331;
    wire n4335;
    wire n4339;
    wire n4343;
    wire n4351;
    wire n6381;
    wire n6384;
    wire n6387;
    wire n6390;
    wire n6393;
    wire n6396;
    wire n6399;
    wire n6402;
    wire n6405;
    wire n6408;
    wire n6411;
    wire n6414;
    wire n6417;
    wire n6420;
    wire n6423;
    wire n6426;
    wire n6429;
    wire n6432;
    wire n6435;
    wire n6438;
    wire n6441;
    wire n6444;
    wire n6447;
    wire n6450;
    wire n6453;
    wire n6456;
    wire n6459;
    wire n6462;
    wire n6465;
    wire n6468;
    wire n6471;
    wire n6474;
    wire n6477;
    wire n6480;
    wire n6483;
    wire n6486;
    wire n6489;
    wire n6492;
    wire n6495;
    wire n6498;
    wire n6501;
    wire n6504;
    wire n6507;
    wire n6510;
    wire n6513;
    wire n6516;
    wire n6519;
    wire n6522;
    wire n6525;
    wire n6528;
    wire n6531;
    wire n6534;
    wire n6537;
    wire n6540;
    wire n6543;
    wire n6546;
    wire n6548;
    wire n6551;
    wire n6554;
    wire n6558;
    wire n6561;
    wire n6564;
    wire n6567;
    wire n6570;
    wire n6573;
    wire n6576;
    wire n6579;
    wire n6582;
    wire n6585;
    wire n6588;
    wire n6591;
    wire n6594;
    wire n6597;
    wire n6600;
    wire n6603;
    wire n6606;
    wire n6609;
    wire n6612;
    wire n6615;
    wire n6617;
    wire n6621;
    wire n6624;
    wire n6627;
    wire n6630;
    wire n6633;
    wire n6636;
    wire n6639;
    wire n6642;
    wire n6645;
    wire n6648;
    wire n6651;
    wire n6654;
    wire n6657;
    wire n6660;
    wire n6663;
    wire n6666;
    wire n6669;
    wire n6672;
    wire n6675;
    wire n6678;
    wire n6681;
    wire n6684;
    wire n6687;
    wire n6690;
    wire n6693;
    wire n6696;
    wire n6699;
    wire n6702;
    wire n6705;
    wire n6708;
    wire n6711;
    wire n6714;
    wire n6716;
    wire n6720;
    wire n6723;
    wire n6726;
    wire n6729;
    wire n6732;
    wire n6735;
    wire n6738;
    wire n6741;
    wire n6744;
    wire n6747;
    wire n6750;
    wire n6753;
    wire n6756;
    wire n6759;
    wire n6762;
    wire n6765;
    wire n6768;
    wire n6771;
    wire n6774;
    wire n6777;
    wire n6780;
    wire n6783;
    wire n6786;
    wire n6789;
    wire n6792;
    wire n6795;
    wire n6798;
    wire n6801;
    wire n6804;
    wire n6807;
    wire n6810;
    wire n6813;
    wire n6816;
    wire n6819;
    wire n6822;
    wire n6825;
    wire n6828;
    wire n6831;
    wire n6834;
    wire n6837;
    wire n6840;
    wire n6843;
    wire n6846;
    wire n6849;
    wire n6852;
    wire n6855;
    wire n6858;
    wire n6861;
    wire n6864;
    wire n6867;
    wire n6870;
    wire n6873;
    wire n6875;
    wire n6878;
    wire n6881;
    wire n6884;
    wire n6887;
    wire n6890;
    wire n6893;
    wire n6896;
    wire n6899;
    wire n6902;
    wire n6905;
    wire n6908;
    wire n6911;
    wire n6914;
    wire n6917;
    wire n6920;
    wire n6923;
    wire n6926;
    wire n6929;
    wire n6932;
    wire n6935;
    wire n6938;
    wire n6941;
    wire n6944;
    wire n6947;
    wire n6950;
    wire n6953;
    wire n6956;
    wire n6959;
    wire n6962;
    wire n6965;
    wire n6968;
    wire n6971;
    wire n6974;
    wire n6977;
    wire n6980;
    wire n6983;
    wire n6986;
    wire n6989;
    wire n6992;
    wire n6995;
    wire n6998;
    wire n7001;
    wire n7004;
    wire n7007;
    wire n7010;
    wire n7013;
    wire n7016;
    wire n7019;
    wire n7022;
    wire n7025;
    wire n7028;
    wire n7032;
    wire n7035;
    wire n7038;
    wire n7041;
    wire n7044;
    wire n7047;
    wire n7050;
    wire n7053;
    wire n7056;
    wire n7059;
    wire n7062;
    wire n7065;
    wire n7068;
    wire n7071;
    wire n7074;
    wire n7077;
    wire n7080;
    wire n7083;
    wire n7086;
    wire n7089;
    wire n7092;
    wire n7095;
    wire n7098;
    wire n7101;
    wire n7104;
    wire n7107;
    wire n7110;
    wire n7113;
    wire n7116;
    wire n7119;
    wire n7122;
    wire n7125;
    wire n7128;
    wire n7131;
    wire n7134;
    wire n7137;
    wire n7140;
    wire n7143;
    wire n7146;
    wire n7149;
    wire n7151;
    wire n7154;
    wire n7157;
    wire n7160;
    wire n7163;
    wire n7166;
    wire n7169;
    wire n7172;
    wire n7176;
    wire n7179;
    wire n7182;
    wire n7185;
    wire n7188;
    wire n7191;
    wire n7194;
    wire n7197;
    wire n7200;
    wire n7203;
    wire n7205;
    wire n7208;
    wire n7211;
    wire n7215;
    wire n7218;
    wire n7221;
    wire n7224;
    wire n7227;
    wire n7230;
    wire n7233;
    wire n7236;
    wire n7239;
    wire n7242;
    wire n7245;
    wire n7248;
    wire n7251;
    wire n7254;
    wire n7257;
    wire n7260;
    wire n7262;
    wire n7265;
    wire n7269;
    wire n7272;
    wire n7274;
    wire n7277;
    wire n7280;
    wire n7283;
    wire n7286;
    wire n7289;
    wire n7292;
    wire n7295;
    wire n7299;
    wire n7302;
    wire n7304;
    wire n7308;
    wire n7311;
    wire n7314;
    wire n7317;
    wire n7320;
    wire n7323;
    wire n7326;
    wire n7329;
    wire n7332;
    wire n7335;
    wire n7338;
    wire n7341;
    wire n7344;
    wire n7347;
    wire n7350;
    wire n7353;
    wire n7356;
    wire n7359;
    wire n7362;
    wire n7364;
    wire n7368;
    wire n7371;
    wire n7374;
    wire n7376;
    wire n7379;
    wire n7382;
    wire n7385;
    wire n7388;
    wire n7391;
    wire n7394;
    wire n7397;
    wire n7400;
    wire n7403;
    wire n7406;
    wire n7409;
    wire n7412;
    wire n7415;
    wire n7419;
    wire n7422;
    wire n7425;
    wire n7428;
    wire n7431;
    wire n7434;
    wire n7437;
    wire n7440;
    wire n7443;
    wire n7446;
    wire n7449;
    wire n7451;
    wire n7454;
    wire n7457;
    wire n7460;
    wire n7463;
    wire n7466;
    wire n7470;
    wire n7473;
    wire n7476;
    wire n7479;
    wire n7482;
    wire n7485;
    wire n7487;
    wire n7491;
    wire n7493;
    wire n7496;
    wire n7499;
    wire n7502;
    wire n7505;
    wire n7508;
    wire n7511;
    wire n7514;
    wire n7517;
    wire n7520;
    wire n7524;
    wire n7527;
    wire n7530;
    wire n7533;
    wire n7536;
    wire n7539;
    wire n7542;
    wire n7545;
    wire n7547;
    wire n7550;
    wire n7554;
    wire n7556;
    wire n7559;
    wire n7562;
    wire n7565;
    wire n7568;
    wire n7571;
    wire n7575;
    wire n7577;
    wire n7580;
    wire n7584;
    wire n7587;
    wire n7589;
    wire n7592;
    wire n7595;
    wire n7598;
    wire n7602;
    wire n7604;
    wire n7607;
    wire n7610;
    wire n7613;
    wire n7616;
    wire n7619;
    wire n7622;
    wire n7625;
    wire n7629;
    wire n7632;
    wire n7635;
    wire n7638;
    wire n7641;
    wire n7644;
    wire n7647;
    wire n7650;
    wire n7653;
    wire n7656;
    wire n7659;
    wire n7662;
    wire n7665;
    wire n7668;
    wire n7671;
    wire n7674;
    wire n7677;
    wire n7680;
    wire n7683;
    wire n7686;
    wire n7689;
    wire n7692;
    wire n7694;
    wire n7698;
    wire n7701;
    wire n7704;
    wire n7706;
    wire n7709;
    wire n7712;
    wire n7715;
    wire n7718;
    wire n7722;
    wire n7725;
    wire n7727;
    wire n7730;
    wire n7733;
    wire n7737;
    wire n7740;
    wire n7742;
    wire n7745;
    wire n7748;
    wire n7751;
    wire n7754;
    wire n7758;
    wire n7761;
    wire n7764;
    wire n7767;
    wire n7769;
    wire n7772;
    wire n7775;
    wire n7779;
    wire n7782;
    wire n7785;
    wire n7788;
    wire n7790;
    wire n7793;
    wire n7796;
    wire n7799;
    wire n7802;
    wire n7805;
    wire n7808;
    wire n7812;
    wire n7814;
    wire n7818;
    wire n7821;
    wire n7824;
    wire n7826;
    wire n7829;
    wire n7832;
    wire n7835;
    wire n7838;
    wire n7841;
    wire n7844;
    wire n7847;
    wire n7850;
    wire n7854;
    wire n7857;
    wire n7860;
    wire n7863;
    wire n7865;
    wire n7868;
    wire n7871;
    wire n7875;
    wire n7878;
    wire n7881;
    wire n7884;
    wire n7887;
    wire n7890;
    wire n7893;
    wire n7896;
    wire n7899;
    wire n7901;
    wire n7904;
    wire n7907;
    wire n7910;
    wire n7913;
    wire n7916;
    wire n7919;
    wire n7922;
    wire n7925;
    wire n7928;
    wire n7931;
    wire n7934;
    wire n7937;
    wire n7940;
    wire n7943;
    wire n7946;
    wire n7949;
    wire n7952;
    wire n7955;
    wire n7958;
    wire n7961;
    wire n7964;
    wire n7968;
    wire n7971;
    wire n7974;
    wire n7977;
    wire n7980;
    wire n7982;
    wire n7985;
    wire n7988;
    wire n7991;
    wire n7995;
    wire n7998;
    wire n8000;
    wire n8004;
    wire n8007;
    wire n8010;
    wire n8013;
    wire n8016;
    wire n8019;
    wire n8021;
    wire n8024;
    wire n8027;
    wire n8030;
    wire n8033;
    wire n8036;
    wire n8039;
    wire n8042;
    wire n8045;
    wire n8048;
    wire n8052;
    wire n8055;
    wire n8058;
    wire n8061;
    wire n8064;
    wire n8066;
    wire n8069;
    wire n8072;
    wire n8075;
    wire n8078;
    wire n8081;
    wire n8084;
    wire n8087;
    wire n8090;
    wire n8094;
    wire n8097;
    wire n8099;
    wire n8102;
    wire n8105;
    wire n8109;
    wire n8112;
    wire n8115;
    wire n8117;
    wire n8120;
    wire n8124;
    wire n8127;
    wire n8130;
    wire n8132;
    wire n8135;
    wire n8138;
    wire n8141;
    wire n8144;
    wire n8147;
    wire n8150;
    wire n8153;
    wire n8156;
    wire n8159;
    wire n8163;
    wire n8166;
    wire n8169;
    wire n8172;
    wire n8175;
    wire n8178;
    wire n8181;
    wire n8184;
    wire n8187;
    wire n8190;
    wire n8193;
    wire n8196;
    wire n8199;
    wire n8202;
    wire n8205;
    wire n8208;
    wire n8211;
    wire n8213;
    wire n8217;
    wire n8219;
    wire n8223;
    wire n8226;
    wire n8229;
    wire n8232;
    wire n8235;
    wire n8238;
    wire n8240;
    wire n8243;
    wire n8246;
    wire n8249;
    wire n8252;
    wire n8255;
    wire n8258;
    wire n8261;
    wire n8264;
    wire n8267;
    wire n8271;
    wire n8274;
    wire n8277;
    wire n8279;
    wire n8283;
    wire n8286;
    wire n8289;
    wire n8292;
    wire n8295;
    wire n8298;
    wire n8301;
    wire n8304;
    wire n8307;
    wire n8310;
    wire n8313;
    wire n8316;
    wire n8318;
    wire n8321;
    wire n8324;
    wire n8327;
    wire n8331;
    wire n8334;
    wire n8337;
    wire n8340;
    wire n8343;
    wire n8346;
    wire n8348;
    wire n8351;
    wire n8354;
    wire n8357;
    wire n8360;
    wire n8364;
    wire n8367;
    wire n8369;
    wire n8372;
    wire n8375;
    wire n8378;
    wire n8382;
    wire n8385;
    wire n8388;
    wire n8390;
    wire n8393;
    wire n8397;
    wire n8400;
    wire n8403;
    wire n8406;
    wire n8409;
    wire n8412;
    wire n8415;
    wire n8418;
    wire n8421;
    wire n8423;
    wire n8427;
    wire n8429;
    wire n8432;
    wire n8435;
    wire n8438;
    wire n8441;
    wire n8444;
    wire n8447;
    wire n8451;
    wire n8454;
    wire n8457;
    wire n8460;
    wire n8462;
    wire n8466;
    wire n8469;
    wire n8472;
    wire n8475;
    wire n8478;
    wire n8481;
    wire n8484;
    wire n8487;
    wire n8489;
    wire n8493;
    wire n8495;
    wire n8498;
    wire n8501;
    wire n8504;
    wire n8507;
    wire n8510;
    wire n8513;
    wire n8516;
    wire n8519;
    wire n8522;
    wire n8525;
    wire n8528;
    wire n8531;
    wire n8535;
    wire n8538;
    wire n8541;
    wire n8543;
    wire n8547;
    wire n8549;
    wire n8552;
    wire n8555;
    wire n8558;
    wire n8561;
    wire n8564;
    wire n8567;
    wire n8570;
    wire n8573;
    wire n8576;
    wire n8579;
    wire n8582;
    wire n8585;
    wire n8588;
    wire n8591;
    wire n8594;
    wire n8597;
    wire n8600;
    wire n8603;
    wire n8606;
    wire n8609;
    wire n8613;
    wire n8616;
    wire n8618;
    wire n8621;
    wire n8624;
    wire n8627;
    wire n8630;
    wire n8633;
    wire n8636;
    wire n8639;
    wire n8642;
    wire n8646;
    wire n8649;
    wire n8652;
    wire n8655;
    wire n8658;
    wire n8661;
    wire n8664;
    wire n8667;
    wire n8670;
    wire n8673;
    wire n8676;
    wire n8679;
    wire n8682;
    wire n8684;
    wire n8687;
    wire n8690;
    wire n8693;
    wire n8696;
    wire n8699;
    wire n8702;
    wire n8705;
    wire n8708;
    wire n8711;
    wire n8715;
    wire n8718;
    wire n8720;
    wire n8724;
    wire n8726;
    wire n8729;
    wire n8732;
    wire n8735;
    wire n8738;
    wire n8741;
    wire n8744;
    wire n8747;
    wire n8750;
    wire n8753;
    wire n8756;
    wire n8759;
    wire n8762;
    wire n8765;
    wire n8768;
    wire n8771;
    wire n8774;
    wire n8777;
    wire n8781;
    wire n8784;
    wire n8787;
    wire n8790;
    wire n8793;
    wire n8796;
    wire n8799;
    wire n8801;
    wire n8804;
    wire n8807;
    wire n8810;
    wire n8813;
    wire n8816;
    wire n8819;
    wire n8823;
    wire n8826;
    wire n8828;
    wire n8832;
    wire n8835;
    wire n8838;
    wire n8841;
    wire n8844;
    wire n8846;
    wire n8849;
    wire n8852;
    wire n8856;
    wire n8859;
    wire n8861;
    wire n8864;
    wire n8867;
    wire n8870;
    wire n8873;
    wire n8876;
    wire n8879;
    wire n8882;
    wire n8885;
    wire n8888;
    wire n8891;
    wire n8895;
    wire n8898;
    wire n8900;
    wire n8903;
    wire n8906;
    wire n8909;
    wire n8912;
    wire n8915;
    wire n8918;
    wire n8921;
    wire n8924;
    wire n8927;
    wire n8930;
    wire n8933;
    wire n8936;
    wire n8939;
    wire n8942;
    wire n8945;
    wire n8948;
    wire n8951;
    wire n8954;
    wire n8957;
    wire n8960;
    wire n8963;
    wire n8966;
    wire n8969;
    wire n8972;
    wire n8975;
    wire n8978;
    wire n8981;
    wire n8984;
    wire n8987;
    wire n8990;
    wire n8993;
    wire n8996;
    wire n8999;
    wire n9002;
    wire n9005;
    wire n9008;
    wire n9011;
    wire n9014;
    wire n9018;
    wire n9020;
    wire n9023;
    wire n9026;
    wire n9029;
    wire n9032;
    wire n9035;
    wire n9038;
    wire n9042;
    wire n9045;
    wire n9047;
    wire n9050;
    wire n9053;
    wire n9056;
    wire n9059;
    wire n9062;
    wire n9066;
    wire n9069;
    wire n9072;
    wire n9074;
    wire n9077;
    wire n9081;
    wire n9084;
    wire n9086;
    wire n9089;
    wire n9092;
    wire n9095;
    wire n9098;
    wire n9101;
    wire n9104;
    wire n9107;
    wire n9111;
    wire n9113;
    wire n9116;
    wire n9120;
    wire n9122;
    wire n9125;
    wire n9128;
    wire n9131;
    wire n9134;
    wire n9137;
    wire n9140;
    wire n9143;
    wire n9146;
    wire n9149;
    wire n9152;
    wire n9155;
    wire n9158;
    wire n9161;
    wire n9164;
    wire n9167;
    wire n9170;
    wire n9173;
    wire n9176;
    wire n9179;
    wire n9182;
    wire n9185;
    wire n9188;
    wire n9191;
    wire n9194;
    wire n9197;
    wire n9200;
    wire n9203;
    wire n9206;
    wire n9209;
    wire n9212;
    wire n9215;
    wire n9219;
    wire n9222;
    wire n9224;
    wire n9227;
    wire n9230;
    wire n9233;
    wire n9236;
    wire n9239;
    wire n9242;
    wire n9245;
    wire n9248;
    wire n9251;
    wire n9254;
    wire n9257;
    wire n9260;
    wire n9263;
    wire n9266;
    wire n9269;
    wire n9272;
    wire n9275;
    wire n9278;
    wire n9281;
    wire n9284;
    wire n9287;
    wire n9290;
    wire n9293;
    wire n9296;
    wire n9299;
    wire n9302;
    wire n9305;
    wire n9308;
    wire n9311;
    wire n9314;
    wire n9317;
    wire n9320;
    wire n9323;
    wire n9326;
    wire n9329;
    wire n9332;
    wire n9335;
    wire n9338;
    wire n9341;
    wire n9344;
    wire n9347;
    wire n9350;
    wire n9353;
    wire n9356;
    wire n9359;
    wire n9363;
    wire n9365;
    wire n9369;
    wire n9372;
    wire n9375;
    wire n9377;
    wire n9380;
    wire n9383;
    wire n9386;
    wire n9389;
    wire n9392;
    wire n9396;
    wire n9399;
    wire n9402;
    wire n9405;
    wire n9408;
    wire n9410;
    wire n9413;
    wire n9416;
    wire n9419;
    wire n9422;
    wire n9425;
    wire n9428;
    wire n9431;
    wire n9434;
    wire n9437;
    wire n9440;
    wire n9443;
    wire n9446;
    wire n9449;
    wire n9452;
    wire n9455;
    wire n9459;
    wire n9461;
    wire n9465;
    wire n9468;
    wire n9470;
    wire n9473;
    wire n9477;
    wire n9480;
    wire n9482;
    wire n9485;
    wire n9489;
    wire n9491;
    wire n9494;
    wire n9497;
    wire n9500;
    wire n9503;
    wire n9506;
    wire n9509;
    wire n9512;
    wire n9515;
    wire n9518;
    wire n9521;
    wire n9524;
    wire n9527;
    wire n9530;
    wire n9533;
    wire n9536;
    wire n9539;
    wire n9542;
    wire n9545;
    wire n9548;
    wire n9551;
    wire n9555;
    wire n9558;
    wire n9561;
    wire n9564;
    wire n9567;
    wire n9570;
    wire n9572;
    wire n9575;
    wire n9579;
    wire n9582;
    wire n9585;
    wire n9588;
    wire n9591;
    wire n9594;
    wire n9597;
    wire n9600;
    wire n9603;
    wire n9606;
    wire n9608;
    wire n9611;
    wire n9614;
    wire n9617;
    wire n9620;
    wire n9623;
    wire n9626;
    wire n9629;
    wire n9632;
    wire n9635;
    wire n9638;
    wire n9641;
    wire n9644;
    wire n9647;
    wire n9650;
    wire n9653;
    wire n9656;
    wire n9659;
    wire n9662;
    wire n9665;
    wire n9668;
    wire n9671;
    wire n9674;
    wire n9677;
    wire n9680;
    wire n9683;
    wire n9686;
    wire n9689;
    wire n9692;
    wire n9695;
    wire n9698;
    wire n9701;
    wire n9704;
    wire n9707;
    wire n9710;
    wire n9713;
    wire n9716;
    wire n9719;
    wire n9722;
    wire n9725;
    wire n9728;
    wire n9731;
    wire n9735;
    wire n9738;
    wire n9741;
    wire n9744;
    wire n9746;
    wire n9749;
    wire n9752;
    wire n9755;
    wire n9758;
    wire n9761;
    wire n9764;
    wire n9767;
    wire n9770;
    wire n9773;
    wire n9776;
    wire n9779;
    wire n9782;
    wire n9785;
    wire n9788;
    wire n9791;
    wire n9794;
    wire n9797;
    wire n9800;
    wire n9803;
    wire n9806;
    wire n9809;
    wire n9812;
    wire n9815;
    wire n9818;
    wire n9821;
    wire n9824;
    wire n9827;
    wire n9830;
    wire n9833;
    wire n9836;
    wire n9839;
    wire n9842;
    wire n9845;
    wire n9848;
    wire n9851;
    wire n9854;
    wire n9857;
    wire n9860;
    wire n9863;
    wire n9866;
    wire n9869;
    wire n9872;
    wire n9875;
    wire n9878;
    wire n9881;
    wire n9884;
    wire n9887;
    wire n9890;
    wire n9893;
    wire n9896;
    wire n9899;
    wire n9902;
    wire n9905;
    wire n9908;
    wire n9911;
    wire n9914;
    wire n9917;
    wire n9920;
    wire n9923;
    wire n9926;
    wire n9929;
    wire n9932;
    wire n9935;
    wire n9938;
    wire n9941;
    wire n9944;
    wire n9947;
    wire n9950;
    wire n9953;
    wire n9956;
    wire n9959;
    wire n9962;
    wire n9965;
    wire n9968;
    wire n9971;
    wire n9974;
    wire n9977;
    wire n9980;
    wire n9983;
    wire n9986;
    wire n9989;
    wire n9992;
    wire n9995;
    wire n9999;
    wire n10002;
    wire n10005;
    wire n10008;
    wire n10011;
    wire n10014;
    wire n10017;
    wire n10019;
    wire n10023;
    wire n10026;
    wire n10029;
    wire n10031;
    wire n10035;
    wire n10038;
    wire n10041;
    wire n10044;
    wire n10047;
    wire n10050;
    wire n10053;
    wire n10056;
    wire n10059;
    wire n10061;
    wire n10065;
    wire n10068;
    wire n10071;
    wire n10074;
    wire n10076;
    wire n10079;
    wire n10082;
    wire n10085;
    wire n10088;
    wire n10091;
    wire n10094;
    wire n10097;
    wire n10100;
    wire n10103;
    wire n10106;
    wire n10110;
    wire n10113;
    wire n10116;
    wire n10119;
    wire n10122;
    wire n10125;
    wire n10127;
    wire n10130;
    wire n10133;
    wire n10136;
    wire n10139;
    wire n10142;
    wire n10145;
    wire n10148;
    wire n10151;
    wire n10154;
    wire n10157;
    wire n10160;
    wire n10163;
    wire n10166;
    wire n10169;
    wire n10172;
    wire n10175;
    wire n10178;
    wire n10181;
    wire n10184;
    wire n10187;
    wire n10190;
    wire n10193;
    wire n10196;
    wire n10199;
    wire n10202;
    wire n10205;
    wire n10208;
    wire n10211;
    wire n10214;
    wire n10218;
    wire n10221;
    wire n10223;
    wire n10226;
    wire n10229;
    wire n10232;
    wire n10235;
    wire n10238;
    wire n10241;
    wire n10244;
    wire n10247;
    wire n10250;
    wire n10253;
    wire n10256;
    wire n10259;
    wire n10262;
    wire n10265;
    wire n10268;
    wire n10271;
    wire n10274;
    wire n10277;
    wire n10280;
    wire n10283;
    wire n10286;
    wire n10289;
    wire n10292;
    wire n10295;
    wire n10298;
    wire n10301;
    wire n10304;
    wire n10307;
    wire n10310;
    wire n10313;
    wire n10316;
    wire n10319;
    wire n10322;
    wire n10325;
    wire n10328;
    wire n10331;
    wire n10334;
    wire n10337;
    wire n10340;
    wire n10343;
    wire n10346;
    wire n10349;
    wire n10352;
    wire n10355;
    wire n10358;
    wire n10361;
    wire n10364;
    wire n10367;
    wire n10370;
    wire n10373;
    wire n10376;
    wire n10379;
    wire n10382;
    wire n10385;
    wire n10388;
    wire n10392;
    wire n10394;
    wire n10397;
    wire n10400;
    wire n10403;
    wire n10406;
    wire n10409;
    wire n10412;
    wire n10415;
    wire n10418;
    wire n10421;
    wire n10424;
    wire n10427;
    wire n10430;
    wire n10433;
    wire n10436;
    wire n10439;
    wire n10442;
    wire n10445;
    wire n10448;
    wire n10451;
    wire n10454;
    wire n10457;
    wire n10460;
    wire n10463;
    wire n10466;
    wire n10469;
    wire n10472;
    wire n10475;
    wire n10478;
    wire n10481;
    wire n10484;
    wire n10487;
    wire n10490;
    wire n10493;
    wire n10496;
    wire n10499;
    wire n10502;
    wire n10505;
    wire n10508;
    wire n10511;
    wire n10514;
    wire n10517;
    wire n10520;
    wire n10523;
    wire n10526;
    wire n10529;
    wire n10532;
    wire n10535;
    wire n10538;
    wire n10541;
    wire n10544;
    wire n10547;
    wire n10550;
    wire n10553;
    wire n10556;
    wire n10559;
    wire n10562;
    wire n10565;
    wire n10568;
    wire n10571;
    wire n10574;
    wire n10577;
    wire n10580;
    wire n10583;
    wire n10586;
    wire n10589;
    wire n10592;
    wire n10595;
    wire n10598;
    wire n10601;
    wire n10604;
    wire n10607;
    wire n10610;
    wire n10613;
    wire n10616;
    wire n10619;
    wire n10622;
    wire n10625;
    wire n10628;
    wire n10631;
    wire n10634;
    wire n10637;
    wire n10640;
    wire n10643;
    wire n10646;
    wire n10649;
    wire n10652;
    wire n10655;
    wire n10658;
    wire n10661;
    wire n10664;
    wire n10667;
    wire n10670;
    wire n10673;
    wire n10676;
    wire n10679;
    wire n10682;
    wire n10685;
    wire n10688;
    wire n10691;
    wire n10694;
    wire n10697;
    wire n10700;
    wire n10703;
    wire n10706;
    wire n10709;
    wire n10712;
    wire n10715;
    wire n10718;
    wire n10721;
    wire n10724;
    wire n10727;
    wire n10731;
    wire n10734;
    wire n10737;
    wire n10740;
    wire n10743;
    wire n10746;
    wire n10749;
    wire n10752;
    wire n10755;
    wire n10758;
    wire n10761;
    wire n10764;
    wire n10766;
    wire n10769;
    wire n10772;
    wire n10775;
    wire n10778;
    wire n10781;
    wire n10784;
    wire n10787;
    wire n10790;
    wire n10793;
    wire n10796;
    wire n10799;
    wire n10802;
    wire n10805;
    wire n10808;
    wire n10811;
    wire n10814;
    wire n10817;
    wire n10820;
    wire n10823;
    wire n10826;
    wire n10829;
    wire n10832;
    wire n10835;
    wire n10838;
    wire n10841;
    wire n10844;
    wire n10847;
    wire n10850;
    wire n10853;
    wire n10856;
    wire n10859;
    wire n10862;
    wire n10865;
    wire n10868;
    wire n10871;
    wire n10874;
    wire n10877;
    wire n10880;
    wire n10883;
    wire n10886;
    wire n10889;
    wire n10892;
    wire n10895;
    wire n10899;
    wire n10902;
    wire n10904;
    wire n10907;
    wire n10910;
    wire n10913;
    wire n10916;
    wire n10919;
    wire n10922;
    wire n10925;
    wire n10928;
    wire n10931;
    wire n10934;
    wire n10937;
    wire n10940;
    wire n10943;
    wire n10946;
    wire n10949;
    wire n10952;
    wire n10955;
    wire n10958;
    wire n10961;
    wire n10964;
    wire n10967;
    wire n10970;
    wire n10973;
    wire n10976;
    wire n10979;
    wire n10982;
    wire n10986;
    wire n10989;
    wire n10991;
    wire n10994;
    wire n10997;
    wire n11000;
    wire n11003;
    wire n11006;
    wire n11009;
    wire n11012;
    wire n11015;
    wire n11018;
    wire n11021;
    wire n11024;
    wire n11027;
    wire n11030;
    wire n11033;
    wire n11036;
    wire n11039;
    wire n11042;
    wire n11045;
    wire n11048;
    wire n11051;
    wire n11054;
    wire n11057;
    wire n11060;
    wire n11063;
    wire n11066;
    wire n11069;
    wire n11072;
    wire n11075;
    wire n11078;
    wire n11081;
    wire n11084;
    wire n11087;
    wire n11090;
    wire n11093;
    wire n11096;
    wire n11099;
    wire n11102;
    wire n11105;
    wire n11108;
    wire n11112;
    wire n11114;
    wire n11117;
    wire n11120;
    wire n11123;
    wire n11127;
    wire n11130;
    wire n11133;
    wire n11135;
    wire n11138;
    wire n11141;
    wire n11144;
    wire n11147;
    wire n11150;
    wire n11153;
    wire n11156;
    wire n11159;
    wire n11162;
    wire n11165;
    wire n11168;
    wire n11171;
    wire n11174;
    wire n11177;
    wire n11180;
    wire n11183;
    wire n11186;
    wire n11189;
    wire n11192;
    wire n11195;
    wire n11198;
    wire n11201;
    wire n11204;
    wire n11207;
    wire n11210;
    wire n11213;
    wire n11216;
    wire n11219;
    wire n11222;
    wire n11225;
    wire n11228;
    wire n11231;
    wire n11234;
    wire n11237;
    wire n11240;
    wire n11243;
    wire n11246;
    wire n11249;
    wire n11253;
    wire n11255;
    wire n11258;
    wire n11261;
    wire n11264;
    wire n11267;
    wire n11270;
    wire n11273;
    wire n11276;
    wire n11279;
    wire n11282;
    wire n11285;
    wire n11288;
    wire n11291;
    wire n11294;
    wire n11297;
    wire n11300;
    wire n11303;
    wire n11306;
    wire n11309;
    wire n11312;
    wire n11315;
    wire n11318;
    wire n11321;
    wire n11324;
    wire n11327;
    wire n11330;
    wire n11333;
    wire n11336;
    wire n11339;
    wire n11342;
    wire n11345;
    wire n11348;
    wire n11351;
    wire n11354;
    wire n11357;
    wire n11360;
    wire n11363;
    wire n11366;
    wire n11369;
    wire n11372;
    wire n11375;
    wire n11378;
    wire n11381;
    wire n11384;
    wire n11387;
    wire n11391;
    wire n11394;
    wire n11396;
    wire n11399;
    wire n11402;
    wire n11405;
    wire n11408;
    wire n11411;
    wire n11414;
    wire n11418;
    wire n11421;
    wire n11424;
    wire n11426;
    wire n11429;
    wire n11432;
    wire n11435;
    wire n11438;
    wire n11441;
    wire n11444;
    wire n11447;
    wire n11450;
    wire n11453;
    wire n11456;
    wire n11459;
    wire n11462;
    wire n11465;
    wire n11468;
    wire n11471;
    wire n11474;
    wire n11477;
    wire n11480;
    wire n11483;
    wire n11486;
    wire n11489;
    wire n11492;
    wire n11495;
    wire n11498;
    wire n11501;
    wire n11504;
    wire n11507;
    wire n11510;
    wire n11513;
    wire n11516;
    wire n11519;
    wire n11522;
    wire n11525;
    wire n11528;
    wire n11531;
    wire n11534;
    wire n11537;
    wire n11540;
    wire n11544;
    wire n11547;
    wire n11549;
    wire n11552;
    wire n11555;
    wire n11558;
    wire n11561;
    wire n11564;
    wire n11567;
    wire n11570;
    wire n11573;
    wire n11576;
    wire n11579;
    wire n11582;
    wire n11585;
    wire n11588;
    wire n11591;
    wire n11594;
    wire n11597;
    wire n11600;
    wire n11603;
    wire n11606;
    wire n11609;
    wire n11612;
    wire n11615;
    wire n11618;
    wire n11621;
    wire n11624;
    wire n11627;
    wire n11630;
    wire n11633;
    wire n11636;
    wire n11640;
    wire n11643;
    wire n11646;
    wire n11649;
    wire n11652;
    wire n11655;
    wire n11658;
    wire n11661;
    wire n11664;
    wire n11667;
    wire n11670;
    wire n11673;
    wire n11676;
    wire n11678;
    wire n11681;
    wire n11684;
    wire n11687;
    wire n11690;
    wire n11693;
    wire n11696;
    wire n11699;
    wire n11702;
    wire n11705;
    wire n11708;
    wire n11711;
    wire n11714;
    wire n11717;
    wire n11720;
    wire n11723;
    wire n11726;
    wire n11729;
    wire n11732;
    wire n11735;
    wire n11738;
    wire n11741;
    wire n11744;
    wire n11747;
    wire n11750;
    wire n11753;
    wire n11756;
    wire n11759;
    wire n11762;
    wire n11765;
    wire n11768;
    wire n11771;
    wire n11774;
    wire n11777;
    wire n11780;
    wire n11783;
    wire n11786;
    wire n11789;
    wire n11792;
    wire n11795;
    wire n11798;
    wire n11801;
    wire n11804;
    wire n11807;
    wire n11810;
    wire n11813;
    wire n11816;
    wire n11819;
    wire n11822;
    wire n11825;
    wire n11828;
    wire n11831;
    wire n11834;
    wire n11837;
    wire n11840;
    wire n11843;
    wire n11846;
    wire n11849;
    wire n11852;
    wire n11855;
    wire n11858;
    wire n11861;
    wire n11864;
    wire n11867;
    wire n11870;
    wire n11873;
    wire n11876;
    wire n11879;
    wire n11882;
    wire n11885;
    wire n11888;
    wire n11891;
    wire n11894;
    wire n11897;
    wire n11900;
    wire n11903;
    wire n11906;
    wire n11909;
    wire n11912;
    wire n11915;
    wire n11918;
    wire n11921;
    wire n11924;
    wire n11927;
    wire n11930;
    wire n11933;
    wire n11936;
    wire n11939;
    wire n11942;
    wire n11945;
    wire n11948;
    wire n11951;
    wire n11954;
    wire n11957;
    wire n11960;
    wire n11964;
    wire n11966;
    wire n11969;
    wire n11972;
    wire n11975;
    wire n11978;
    wire n11981;
    wire n11984;
    wire n11987;
    wire n11990;
    wire n11993;
    wire n11996;
    wire n11999;
    wire n12002;
    wire n12005;
    wire n12008;
    wire n12011;
    wire n12014;
    wire n12017;
    wire n12020;
    wire n12023;
    wire n12026;
    wire n12029;
    wire n12032;
    wire n12035;
    wire n12038;
    wire n12041;
    wire n12044;
    wire n12047;
    wire n12050;
    wire n12053;
    wire n12056;
    wire n12059;
    wire n12062;
    wire n12065;
    wire n12068;
    wire n12071;
    wire n12074;
    wire n12077;
    wire n12080;
    wire n12083;
    wire n12086;
    wire n12089;
    wire n12092;
    wire n12095;
    wire n12098;
    wire n12101;
    wire n12104;
    wire n12107;
    wire n12110;
    wire n12113;
    wire n12116;
    wire n12119;
    wire n12122;
    wire n12125;
    wire n12128;
    wire n12131;
    wire n12134;
    wire n12137;
    wire n12140;
    wire n12143;
    wire n12146;
    wire n12149;
    wire n12152;
    wire n12155;
    wire n12158;
    wire n12161;
    wire n12164;
    wire n12167;
    wire n12170;
    wire n12173;
    wire n12176;
    wire n12179;
    wire n12182;
    wire n12185;
    wire n12188;
    wire n12191;
    wire n12194;
    wire n12197;
    wire n12200;
    wire n12203;
    wire n12206;
    wire n12209;
    wire n12212;
    wire n12215;
    wire n12218;
    wire n12221;
    wire n12224;
    wire n12227;
    wire n12230;
    wire n12233;
    wire n12236;
    wire n12239;
    wire n12242;
    wire n12245;
    wire n12248;
    wire n12251;
    wire n12254;
    wire n12257;
    wire n12260;
    wire n12263;
    wire n12266;
    wire n12269;
    wire n12272;
    wire n12275;
    wire n12278;
    wire n12284;
    wire n12287;
    wire n12290;
    wire n12293;
    wire n12296;
    wire n12299;
    wire n12302;
    wire n12305;
    wire n12308;
    wire n12311;
    wire n12314;
    wire n12317;
    wire n12320;
    wire n12323;
    wire n12326;
    wire n12329;
    wire n12332;
    wire n12335;
    wire n12338;
    wire n12341;
    wire n12344;
    wire n12347;
    wire n12350;
    wire n12353;
    wire n12356;
    wire n12359;
    wire n12362;
    wire n12368;
    wire n12371;
    wire n12374;
    wire n12377;
    wire n12380;
    wire n12383;
    wire n12386;
    wire n12389;
    wire n12392;
    wire n12395;
    wire n12398;
    wire n12401;
    wire n12404;
    wire n12407;
    wire n12410;
    wire n12413;
    wire n12416;
    wire n12419;
    wire n12422;
    wire n12425;
    wire n12428;
    wire n12431;
    wire n12437;
    wire n12440;
    wire n12443;
    wire n12446;
    wire n12449;
    wire n12452;
    wire n12455;
    wire n12458;
    wire n12461;
    wire n12464;
    wire n12467;
    wire n12470;
    wire n12473;
    wire n12476;
    wire n12479;
    wire n12482;
    wire n12485;
    wire n12488;
    wire n12491;
    wire n12494;
    wire n12497;
    wire n12500;
    wire n12503;
    wire n12506;
    wire n12509;
    wire n12515;
    wire n12518;
    wire n12521;
    wire n12524;
    wire n12527;
    wire n12530;
    wire n12533;
    wire n12536;
    wire n12539;
    wire n12542;
    wire n12545;
    wire n12548;
    wire n12551;
    wire n12554;
    wire n12557;
    wire n12560;
    wire n12563;
    wire n12566;
    wire n12569;
    wire n12572;
    wire n12575;
    wire n12578;
    wire n12581;
    wire n12584;
    wire n12587;
    wire n12590;
    wire n12596;
    wire n12599;
    wire n12602;
    wire n12605;
    wire n12608;
    wire n12611;
    wire n12614;
    wire n12617;
    wire n12620;
    wire n12623;
    wire n12626;
    wire n12629;
    wire n12632;
    wire n12638;
    wire n12641;
    wire n12644;
    wire n12647;
    wire n12650;
    wire n12653;
    wire n12656;
    wire n12659;
    wire n12662;
    wire n12665;
    wire n12668;
    wire n12674;
    wire n12677;
    wire n12680;
    wire n12683;
    wire n12686;
    wire n12689;
    wire n12692;
    wire n12695;
    wire n12698;
    wire n12701;
    wire n12704;
    wire n12707;
    wire n12710;
    wire n12716;
    wire n12719;
    wire n12722;
    wire n12725;
    wire n12728;
    wire n12731;
    wire n12734;
    wire n12737;
    wire n12743;
    wire n12746;
    wire n12749;
    wire n12752;
    wire n12755;
    wire n12758;
    wire n12761;
    wire n12764;
    wire n12767;
    wire n12770;
    wire n12773;
    wire n12776;
    wire n12782;
    wire n12785;
    wire n12788;
    wire n12791;
    wire n12794;
    wire n12797;
    wire n12800;
    wire n12806;
    wire n12809;
    wire n12812;
    wire n12815;
    wire n12818;
    wire n12821;
    wire n12827;
    wire n12830;
    wire n12833;
    wire n12836;
    wire n12839;
    wire n12845;
    wire n12848;
    wire n12851;
    wire n12854;
    wire n12857;
    wire n12860;
    wire n12866;
    wire n12869;
    wire n12872;
    wire n12875;
    wire n12878;
    wire n12884;
    wire n12887;
    wire n12890;
    wire n12896;
    wire n12899;
    wire n12902;
    wire n12908;
    wire n12911;
    wire n12914;
    wire n12923;
    jnot g0000(.din(G77), .dout(n74));
    jnot g0001(.din(G50), .dout(n77));
    jnot g0002(.din(G58), .dout(n80));
    jnot g0003(.din(G68), .dout(n83));
    jand g0004(.dinb(n80), .dina(n83), .dout(n87));
    jand g0005(.dinb(n7565), .dina(n87), .dout(n91));
    jand g0006(.dinb(n9122), .dina(n91), .dout(n95));
    jnot g0007(.din(G87), .dout(n98));
    jnot g0008(.din(G97), .dout(n101));
    jnot g0009(.din(G107), .dout(n104));
    jand g0010(.dinb(n101), .dina(n104), .dout(n108));
    jor g0011(.dinb(n9722), .dina(n108), .dout(n112));
    jnot g0012(.din(G250), .dout(n115));
    jnot g0013(.din(G257), .dout(n118));
    jnot g0014(.din(G264), .dout(n121));
    jand g0015(.dinb(n118), .dina(n121), .dout(n125));
    jor g0016(.dinb(n9506), .dina(n125), .dout(n129));
    jnot g0017(.din(G13), .dout(n132));
    jand g0018(.dinb(n12131), .dina(n132), .dout(n136));
    jand g0019(.dinb(n12152), .dina(n136), .dout(n140));
    jand g0020(.dinb(n129), .dina(n140), .dout(n144));
    jor g0021(.dinb(n101), .dina(n118), .dout(n148));
    jnot g0022(.din(G244), .dout(n151));
    jor g0023(.dinb(n74), .dina(n151), .dout(n155));
    jnot g0024(.din(G238), .dout(n158));
    jor g0025(.dinb(n83), .dina(n158), .dout(n162));
    jand g0026(.dinb(n155), .dina(n162), .dout(n166));
    jnot g0027(.din(G226), .dout(n169));
    jor g0028(.dinb(n77), .dina(n169), .dout(n173));
    jand g0029(.dinb(n166), .dina(n6402), .dout(n177));
    jand g0030(.dinb(n6399), .dina(n177), .dout(n181));
    jnot g0031(.din(G232), .dout(n184));
    jor g0032(.dinb(n80), .dina(n184), .dout(n188));
    jnot g0033(.din(G116), .dout(n191));
    jnot g0034(.din(G270), .dout(n194));
    jor g0035(.dinb(n191), .dina(n194), .dout(n198));
    jand g0036(.dinb(n188), .dina(n198), .dout(n202));
    jor g0037(.dinb(n104), .dina(n121), .dout(n206));
    jand g0038(.dinb(n202), .dina(n6393), .dout(n210));
    jand g0039(.dinb(G1), .dina(G20), .dout(n214));
    jnot g0040(.din(n214), .dout(n217));
    jor g0041(.dinb(n98), .dina(n115), .dout(n221));
    jand g0042(.dinb(n217), .dina(n221), .dout(n225));
    jand g0043(.dinb(n210), .dina(n6390), .dout(n229));
    jand g0044(.dinb(n181), .dina(n229), .dout(n233));
    jnot g0045(.din(n87), .dout(n236));
    jand g0046(.dinb(n9842), .dina(n236), .dout(n240));
    jnot g0047(.din(n240), .dout(n243));
    jand g0048(.dinb(n12128), .dina(n214), .dout(n247));
    jand g0049(.dinb(n243), .dina(n6548), .dout(n251));
    jor g0050(.dinb(n233), .dina(n251), .dout(n255));
    jor g0051(.dinb(n6387), .dina(n255), .dout(n259));
    jxor g0052(.dinb(n121), .dina(n11123), .dout(n263));
    jxor g0053(.dinb(G250), .dina(G257), .dout(n267));
    jxor g0054(.dinb(n263), .dina(n8547), .dout(n271));
    jnot g0055(.din(n271), .dout(n274));
    jxor g0056(.dinb(n158), .dina(n9191), .dout(n278));
    jxor g0057(.dinb(G226), .dina(G232), .dout(n282));
    jxor g0058(.dinb(n278), .dina(n8724), .dout(n286));
    jxor g0059(.dinb(n274), .dina(n8720), .dout(n290));
    jxor g0060(.dinb(G50), .dina(G58), .dout(n294));
    jxor g0061(.dinb(G68), .dina(G77), .dout(n298));
    jxor g0062(.dinb(n294), .dina(n298), .dout(n302));
    jxor g0063(.dinb(n104), .dina(n11603), .dout(n306));
    jxor g0064(.dinb(G87), .dina(G97), .dout(n310));
    jxor g0065(.dinb(n306), .dina(n8283), .dout(n314));
    jxor g0066(.dinb(n9809), .dina(n314), .dout(n318));
    jand g0067(.dinb(G1), .dina(G13), .dout(n322));
    jand g0068(.dinb(n11558), .dina(n214), .dout(n326));
    jor g0069(.dinb(n11573), .dina(n326), .dout(n330));
    jnot g0070(.din(G1), .dout(n333));
    jand g0071(.dinb(n333), .dina(n11582), .dout(n337));
    jand g0072(.dinb(n12146), .dina(n337), .dout(n341));
    jor g0073(.dinb(n330), .dina(n341), .dout(n345));
    jand g0074(.dinb(n333), .dina(n11555), .dout(n349));
    jor g0075(.dinb(n345), .dina(n11547), .dout(n353));
    jnot g0076(.din(n353), .dout(n356));
    jand g0077(.dinb(n11585), .dina(n356), .dout(n360));
    jand g0078(.dinb(G20), .dina(G116), .dout(n364));
    jnot g0079(.din(G20), .dout(n367));
    jand g0080(.dinb(G33), .dina(G283), .dout(n371));
    jnot g0081(.din(G33), .dout(n374));
    jand g0082(.dinb(n374), .dina(n11426), .dout(n378));
    jor g0083(.dinb(n11483), .dina(n378), .dout(n382));
    jand g0084(.dinb(n11528), .dina(n382), .dout(n386));
    jor g0085(.dinb(n11424), .dina(n386), .dout(n390));
    jand g0086(.dinb(n11549), .dina(n390), .dout(n394));
    jand g0087(.dinb(n11396), .dina(n341), .dout(n398));
    jor g0088(.dinb(n394), .dina(n11394), .dout(n402));
    jor g0089(.dinb(n360), .dina(n402), .dout(n406));
    jnot g0090(.din(n406), .dout(n409));
    jnot g0091(.din(G41), .dout(n412));
    jand g0092(.dinb(n333), .dina(n11276), .dout(n416));
    jand g0093(.dinb(n11333), .dina(n416), .dout(n420));
    jnot g0094(.din(n322), .dout(n423));
    jand g0095(.dinb(G33), .dina(G41), .dout(n427));
    jor g0096(.dinb(n423), .dina(n11255), .dout(n431));
    jand g0097(.dinb(n11264), .dina(n431), .dout(n435));
    jand g0098(.dinb(n11273), .dina(n435), .dout(n439));
    jnot g0099(.din(n427), .dout(n442));
    jand g0100(.dinb(n11570), .dina(n442), .dout(n446));
    jand g0101(.dinb(n374), .dina(n11195), .dout(n450));
    jand g0102(.dinb(n11207), .dina(n450), .dout(n454));
    jand g0103(.dinb(G33), .dina(G303), .dout(n458));
    jnot g0104(.din(G1698), .dout(n461));
    jand g0105(.dinb(n374), .dina(n461), .dout(n465));
    jand g0106(.dinb(n11135), .dina(n465), .dout(n469));
    jor g0107(.dinb(n11133), .dina(n469), .dout(n473));
    jor g0108(.dinb(n11127), .dina(n473), .dout(n477));
    jand g0109(.dinb(n11219), .dina(n477), .dout(n481));
    jnot g0110(.din(n420), .dout(n484));
    jand g0111(.dinb(n11114), .dina(n431), .dout(n488));
    jand g0112(.dinb(n484), .dina(n488), .dout(n492));
    jor g0113(.dinb(n481), .dina(n11112), .dout(n496));
    jor g0114(.dinb(n11249), .dina(n496), .dout(n500));
    jand g0115(.dinb(n11336), .dina(n500), .dout(n504));
    jnot g0116(.din(n504), .dout(n507));
    jnot g0117(.din(G179), .dout(n510));
    jor g0118(.dinb(n10997), .dina(n500), .dout(n514));
    jand g0119(.dinb(n507), .dina(n10991), .dout(n518));
    jor g0120(.dinb(n10989), .dina(n518), .dout(n522));
    jand g0121(.dinb(n10955), .dina(n500), .dout(n526));
    jnot g0122(.din(n500), .dout(n529));
    jand g0123(.dinb(n10907), .dina(n529), .dout(n533));
    jor g0124(.dinb(n11384), .dina(n533), .dout(n537));
    jor g0125(.dinb(n10902), .dina(n537), .dout(n541));
    jand g0126(.dinb(n522), .dina(n541), .dout(n545));
    jnot g0127(.din(G169), .dout(n548));
    jand g0128(.dinb(n11198), .dina(n431), .dout(n552));
    jand g0129(.dinb(n484), .dina(n552), .dout(n556));
    jand g0130(.dinb(n11150), .dina(n450), .dout(n560));
    jand g0131(.dinb(G33), .dina(G294), .dout(n564));
    jnot g0132(.din(n564), .dout(n567));
    jor g0133(.dinb(G33), .dina(G1698), .dout(n571));
    jor g0134(.dinb(n115), .dina(n571), .dout(n575));
    jand g0135(.dinb(n567), .dina(n575), .dout(n579));
    jnot g0136(.din(n579), .dout(n582));
    jor g0137(.dinb(n9521), .dina(n582), .dout(n586));
    jand g0138(.dinb(n11213), .dina(n586), .dout(n590));
    jor g0139(.dinb(n11253), .dina(n590), .dout(n594));
    jor g0140(.dinb(n9524), .dina(n594), .dout(n598));
    jand g0141(.dinb(n9551), .dina(n598), .dout(n602));
    jand g0142(.dinb(n9656), .dina(n356), .dout(n606));
    jor g0143(.dinb(n11576), .dina(n326), .dout(n610));
    jand g0144(.dinb(n11984), .dina(n104), .dout(n614));
    jand g0145(.dinb(n610), .dina(n9489), .dout(n618));
    jand g0146(.dinb(G33), .dina(G116), .dout(n622));
    jand g0147(.dinb(n374), .dina(n9731), .dout(n626));
    jor g0148(.dinb(n9482), .dina(n626), .dout(n630));
    jand g0149(.dinb(n330), .dina(n630), .dout(n634));
    jand g0150(.dinb(n11522), .dina(n634), .dout(n638));
    jor g0151(.dinb(n9480), .dina(n638), .dout(n642));
    jor g0152(.dinb(n606), .dina(n9477), .dout(n646));
    jnot g0153(.din(n646), .dout(n649));
    jnot g0154(.din(n556), .dout(n652));
    jnot g0155(.din(G274), .dout(n655));
    jor g0156(.dinb(n9468), .dina(n446), .dout(n659));
    jor g0157(.dinb(n484), .dina(n659), .dout(n663));
    jnot g0158(.din(n560), .dout(n666));
    jand g0159(.dinb(n666), .dina(n9503), .dout(n670));
    jor g0160(.dinb(n9536), .dina(n670), .dout(n674));
    jand g0161(.dinb(n9461), .dina(n674), .dout(n678));
    jand g0162(.dinb(n9459), .dina(n678), .dout(n682));
    jand g0163(.dinb(n10994), .dina(n682), .dout(n686));
    jor g0164(.dinb(n649), .dina(n686), .dout(n690));
    jor g0165(.dinb(n9494), .dina(n690), .dout(n694));
    jand g0166(.dinb(n10904), .dina(n682), .dout(n698));
    jand g0167(.dinb(n10955), .dina(n598), .dout(n702));
    jor g0168(.dinb(n9470), .dina(n702), .dout(n706));
    jor g0169(.dinb(n9440), .dina(n706), .dout(n710));
    jand g0170(.dinb(n694), .dina(n710), .dout(n714));
    jand g0171(.dinb(n9326), .dina(n450), .dout(n718));
    jnot g0172(.din(n718), .dout(n721));
    jnot g0173(.din(n622), .dout(n724));
    jor g0174(.dinb(n158), .dina(n571), .dout(n728));
    jand g0175(.dinb(n724), .dina(n728), .dout(n732));
    jand g0176(.dinb(n721), .dina(n9299), .dout(n736));
    jand g0177(.dinb(n11243), .dina(n736), .dout(n740));
    jor g0178(.dinb(n9512), .dina(n416), .dout(n744));
    jand g0179(.dinb(n11258), .dina(n416), .dout(n748));
    jnot g0180(.din(n748), .dout(n751));
    jand g0181(.dinb(n9296), .dina(n751), .dout(n755));
    jand g0182(.dinb(n9530), .dina(n755), .dout(n759));
    jor g0183(.dinb(n740), .dina(n759), .dout(n763));
    jand g0184(.dinb(n11018), .dina(n763), .dout(n767));
    jor g0185(.dinb(n9710), .dina(n353), .dout(n771));
    jand g0186(.dinb(n98), .dina(n101), .dout(n775));
    jand g0187(.dinb(n9491), .dina(n775), .dout(n779));
    jand g0188(.dinb(n9281), .dina(n779), .dout(n783));
    jnot g0189(.din(n330), .dout(n786));
    jand g0190(.dinb(G33), .dina(G97), .dout(n790));
    jnot g0191(.din(n790), .dout(n793));
    jor g0192(.dinb(n9272), .dina(n83), .dout(n797));
    jand g0193(.dinb(n11525), .dina(n797), .dout(n801));
    jand g0194(.dinb(n9222), .dina(n801), .dout(n805));
    jor g0195(.dinb(n786), .dina(n805), .dout(n809));
    jor g0196(.dinb(n9275), .dina(n809), .dout(n813));
    jand g0197(.dinb(n9725), .dina(n341), .dout(n817));
    jnot g0198(.din(n817), .dout(n820));
    jand g0199(.dinb(n813), .dina(n9219), .dout(n824));
    jand g0200(.dinb(n9287), .dina(n824), .dout(n828));
    jnot g0201(.din(n732), .dout(n831));
    jor g0202(.dinb(n9317), .dina(n831), .dout(n835));
    jor g0203(.dinb(n9245), .dina(n835), .dout(n839));
    jnot g0204(.din(n744), .dout(n842));
    jor g0205(.dinb(n842), .dina(n9293), .dout(n846));
    jor g0206(.dinb(n11243), .dina(n846), .dout(n850));
    jand g0207(.dinb(n839), .dina(n850), .dout(n854));
    jand g0208(.dinb(n9570), .dina(n854), .dout(n858));
    jor g0209(.dinb(n828), .dina(n858), .dout(n862));
    jor g0210(.dinb(n9290), .dina(n862), .dout(n866));
    jand g0211(.dinb(n10325), .dina(n854), .dout(n870));
    jnot g0212(.din(n771), .dout(n873));
    jnot g0213(.din(n783), .dout(n876));
    jand g0214(.dinb(n374), .dina(n9827), .dout(n880));
    jor g0215(.dinb(n9278), .dina(n880), .dout(n884));
    jor g0216(.dinb(n9263), .dina(n884), .dout(n888));
    jand g0217(.dinb(n9485), .dina(n888), .dout(n892));
    jand g0218(.dinb(n876), .dina(n892), .dout(n896));
    jor g0219(.dinb(n896), .dina(n9251), .dout(n900));
    jor g0220(.dinb(n873), .dina(n900), .dout(n904));
    jand g0221(.dinb(n10913), .dina(n763), .dout(n908));
    jor g0222(.dinb(n904), .dina(n908), .dout(n912));
    jor g0223(.dinb(n9239), .dina(n912), .dout(n916));
    jand g0224(.dinb(n866), .dina(n916), .dout(n920));
    jand g0225(.dinb(n11141), .dina(n431), .dout(n924));
    jand g0226(.dinb(n484), .dina(n924), .dout(n928));
    jnot g0227(.din(n928), .dout(n931));
    jor g0228(.dinb(n9269), .dina(n461), .dout(n935));
    jor g0229(.dinb(n9509), .dina(n935), .dout(n939));
    jnot g0230(.din(n371), .dout(n942));
    jor g0231(.dinb(n151), .dina(n571), .dout(n946));
    jand g0232(.dinb(n942), .dina(n946), .dout(n950));
    jand g0233(.dinb(n939), .dina(n950), .dout(n954));
    jor g0234(.dinb(n9242), .dina(n954), .dout(n958));
    jand g0235(.dinb(n663), .dina(n958), .dout(n962));
    jand g0236(.dinb(n931), .dina(n962), .dout(n966));
    jand g0237(.dinb(n10934), .dina(n966), .dout(n970));
    jor g0238(.dinb(n9698), .dina(n353), .dout(n974));
    jnot g0239(.din(n974), .dout(n977));
    jxor g0240(.dinb(G97), .dina(G107), .dout(n981));
    jand g0241(.dinb(n12158), .dina(n981), .dout(n985));
    jnot g0242(.din(n985), .dout(n988));
    jand g0243(.dinb(G33), .dina(G107), .dout(n992));
    jand g0244(.dinb(n374), .dina(n9812), .dout(n996));
    jor g0245(.dinb(n9086), .dina(n996), .dout(n1000));
    jor g0246(.dinb(n9152), .dina(n1000), .dout(n1004));
    jand g0247(.dinb(n9092), .dina(n1004), .dout(n1008));
    jand g0248(.dinb(n9084), .dina(n1008), .dout(n1012));
    jand g0249(.dinb(n9692), .dina(n341), .dout(n1016));
    jor g0250(.dinb(n1012), .dina(n9113), .dout(n1020));
    jor g0251(.dinb(n977), .dina(n1020), .dout(n1024));
    jand g0252(.dinb(n9515), .dina(n450), .dout(n1028));
    jand g0253(.dinb(n9320), .dina(n465), .dout(n1032));
    jor g0254(.dinb(n11477), .dina(n1032), .dout(n1036));
    jor g0255(.dinb(n9072), .dina(n1036), .dout(n1040));
    jand g0256(.dinb(n11243), .dina(n1040), .dout(n1044));
    jor g0257(.dinb(n11253), .dina(n1044), .dout(n1048));
    jor g0258(.dinb(n9194), .dina(n1048), .dout(n1052));
    jand g0259(.dinb(n10301), .dina(n1052), .dout(n1056));
    jor g0260(.dinb(n9077), .dina(n1056), .dout(n1060));
    jor g0261(.dinb(n9176), .dina(n1060), .dout(n1064));
    jor g0262(.dinb(n11363), .dina(n966), .dout(n1068));
    jnot g0263(.din(n1068), .dout(n1071));
    jnot g0264(.din(n992), .dout(n1074));
    jor g0265(.dinb(n9158), .dina(n74), .dout(n1078));
    jand g0266(.dinb(n11525), .dina(n1078), .dout(n1082));
    jand g0267(.dinb(n9120), .dina(n1082), .dout(n1086));
    jor g0268(.dinb(n786), .dina(n1086), .dout(n1090));
    jor g0269(.dinb(n9161), .dina(n1090), .dout(n1094));
    jnot g0270(.din(n1016), .dout(n1097));
    jand g0271(.dinb(n1094), .dina(n9111), .dout(n1101));
    jand g0272(.dinb(n9173), .dina(n1101), .dout(n1105));
    jand g0273(.dinb(n11000), .dina(n966), .dout(n1109));
    jor g0274(.dinb(n1105), .dina(n1109), .dout(n1113));
    jor g0275(.dinb(n1071), .dina(n1113), .dout(n1117));
    jand g0276(.dinb(n1064), .dina(n9053), .dout(n1121));
    jand g0277(.dinb(n7863), .dina(n1121), .dout(n1125));
    jand g0278(.dinb(n9437), .dina(n1125), .dout(n1129));
    jand g0279(.dinb(n10895), .dina(n1129), .dout(n1133));
    jnot g0280(.din(G45), .dout(n1136));
    jand g0281(.dinb(n412), .dina(n1136), .dout(n1140));
    jor g0282(.dinb(n11990), .dina(n1140), .dout(n1144));
    jnot g0283(.din(n1144), .dout(n1147));
    jand g0284(.dinb(n435), .dina(n1147), .dout(n1151));
    jnot g0285(.din(n1151), .dout(n1154));
    jand g0286(.dinb(n9311), .dina(n450), .dout(n1158));
    jand g0287(.dinb(n8726), .dina(n465), .dout(n1162));
    jor g0288(.dinb(n9146), .dina(n1162), .dout(n1166));
    jor g0289(.dinb(n8130), .dina(n1166), .dout(n1170));
    jand g0290(.dinb(n11237), .dina(n1170), .dout(n1174));
    jnot g0291(.din(n1174), .dout(n1177));
    jor g0292(.dinb(n9182), .dina(n1147), .dout(n1181));
    jor g0293(.dinb(n11237), .dina(n1181), .dout(n1185));
    jand g0294(.dinb(n1177), .dina(n8127), .dout(n1189));
    jand g0295(.dinb(n8132), .dina(n1189), .dout(n1193));
    jnot g0296(.din(n1193), .dout(n1196));
    jand g0297(.dinb(n9542), .dina(n1196), .dout(n1200));
    jand g0298(.dinb(G33), .dina(G87), .dout(n1204));
    jand g0299(.dinb(n374), .dina(n9839), .dout(n1208));
    jor g0300(.dinb(n8124), .dina(n1208), .dout(n1212));
    jand g0301(.dinb(n9224), .dina(n1212), .dout(n1216));
    jand g0302(.dinb(n9089), .dina(n1216), .dout(n1220));
    jand g0303(.dinb(n367), .dina(n322), .dout(n1224));
    jnot g0304(.din(n1224), .dout(n1227));
    jand g0305(.dinb(n333), .dina(n12161), .dout(n1231));
    jnot g0306(.din(n1231), .dout(n1234));
    jand g0307(.dinb(n10355), .dina(n1234), .dout(n1238));
    jand g0308(.dinb(n8115), .dina(n1238), .dout(n1242));
    jand g0309(.dinb(n9140), .dina(n341), .dout(n1246));
    jor g0310(.dinb(n1242), .dina(n8112), .dout(n1250));
    jor g0311(.dinb(n8109), .dina(n1250), .dout(n1254));
    jnot g0312(.din(n1254), .dout(n1257));
    jand g0313(.dinb(n9056), .dina(n1193), .dout(n1261));
    jor g0314(.dinb(n8097), .dina(n1261), .dout(n1265));
    jor g0315(.dinb(n1200), .dina(n1265), .dout(n1269));
    jnot g0316(.din(G200), .dout(n1272));
    jor g0317(.dinb(n8090), .dina(n1193), .dout(n1276));
    jnot g0318(.din(n1276), .dout(n1279));
    jand g0319(.dinb(n9206), .dina(n1193), .dout(n1283));
    jor g0320(.dinb(n8099), .dina(n1283), .dout(n1287));
    jor g0321(.dinb(n1279), .dina(n1287), .dout(n1291));
    jand g0322(.dinb(n1269), .dina(n1291), .dout(n1295));
    jnot g0323(.din(n1295), .dout(n1298));
    jand g0324(.dinb(n9302), .dina(n431), .dout(n1302));
    jand g0325(.dinb(n8147), .dina(n1302), .dout(n1306));
    jand g0326(.dinb(n8741), .dina(n450), .dout(n1310));
    jand g0327(.dinb(n8747), .dina(n465), .dout(n1314));
    jor g0328(.dinb(n9257), .dina(n1314), .dout(n1318));
    jor g0329(.dinb(n7824), .dina(n1318), .dout(n1322));
    jand g0330(.dinb(n11237), .dina(n1322), .dout(n1326));
    jor g0331(.dinb(n8138), .dina(n1326), .dout(n1330));
    jor g0332(.dinb(n7821), .dina(n1330), .dout(n1334));
    jnot g0333(.din(n1334), .dout(n1337));
    jor g0334(.dinb(n9104), .dina(n1337), .dout(n1341));
    jand g0335(.dinb(G33), .dina(G77), .dout(n1345));
    jand g0336(.dinb(n374), .dina(n10154), .dout(n1349));
    jor g0337(.dinb(n7814), .dina(n1349), .dout(n1353));
    jand g0338(.dinb(n330), .dina(n1353), .dout(n1357));
    jand g0339(.dinb(n9989), .dina(n1357), .dout(n1361));
    jand g0340(.dinb(n12161), .dina(n83), .dout(n1365));
    jand g0341(.dinb(n610), .dina(n7812), .dout(n1369));
    jand g0342(.dinb(n786), .dina(n8117), .dout(n1373));
    jand g0343(.dinb(n7796), .dina(n1373), .dout(n1377));
    jor g0344(.dinb(n7788), .dina(n1377), .dout(n1381));
    jor g0345(.dinb(n7782), .dina(n1381), .dout(n1385));
    jor g0346(.dinb(n11060), .dina(n1334), .dout(n1389));
    jand g0347(.dinb(n7775), .dina(n1389), .dout(n1393));
    jand g0348(.dinb(n1341), .dina(n1393), .dout(n1397));
    jand g0349(.dinb(n9200), .dina(n1337), .dout(n1401));
    jand g0350(.dinb(n10424), .dina(n1334), .dout(n1405));
    jor g0351(.dinb(n7772), .dina(n1405), .dout(n1409));
    jor g0352(.dinb(n1401), .dina(n1409), .dout(n1413));
    jnot g0353(.din(n1413), .dout(n1416));
    jor g0354(.dinb(n7769), .dina(n1416), .dout(n1420));
    jand g0355(.dinb(n8759), .dina(n431), .dout(n1424));
    jand g0356(.dinb(n8153), .dina(n1424), .dout(n1428));
    jnot g0357(.din(n1428), .dout(n1431));
    jand g0358(.dinb(n7587), .dina(n450), .dout(n1435));
    jnot g0359(.din(n1435), .dout(n1438));
    jnot g0360(.din(n1345), .dout(n1441));
    jnot g0361(.din(G222), .dout(n1444));
    jor g0362(.dinb(n1444), .dina(n571), .dout(n1448));
    jand g0363(.dinb(n1441), .dina(n1448), .dout(n1452));
    jand g0364(.dinb(n1438), .dina(n7577), .dout(n1456));
    jor g0365(.dinb(n7826), .dina(n1456), .dout(n1460));
    jand g0366(.dinb(n1154), .dina(n1460), .dout(n1464));
    jand g0367(.dinb(n7575), .dina(n1464), .dout(n1468));
    jor g0368(.dinb(n9101), .dina(n1468), .dout(n1472));
    jand g0369(.dinb(n367), .dina(n10388), .dout(n1476));
    jand g0370(.dinb(n10199), .dina(n1476), .dout(n1480));
    jnot g0371(.din(n1480), .dout(n1483));
    jor g0372(.dinb(n7568), .dina(n91), .dout(n1487));
    jand g0373(.dinb(n367), .dina(n374), .dout(n1491));
    jand g0374(.dinb(n8859), .dina(n1491), .dout(n1495));
    jnot g0375(.din(n1495), .dout(n1498));
    jand g0376(.dinb(n1487), .dina(n1498), .dout(n1502));
    jand g0377(.dinb(n7554), .dina(n1502), .dout(n1506));
    jor g0378(.dinb(n9233), .dina(n1506), .dout(n1510));
    jnot g0379(.din(n1510), .dout(n1513));
    jnot g0380(.din(n341), .dout(n1516));
    jand g0381(.dinb(n7556), .dina(n1516), .dout(n1520));
    jnot g0382(.din(n1520), .dout(n1523));
    jor g0383(.dinb(n8690), .dina(n1373), .dout(n1527));
    jand g0384(.dinb(n1523), .dina(n1527), .dout(n1531));
    jor g0385(.dinb(n1513), .dina(n7547), .dout(n1535));
    jnot g0386(.din(n1452), .dout(n1538));
    jor g0387(.dinb(n7580), .dina(n1538), .dout(n1542));
    jand g0388(.dinb(n11231), .dina(n1542), .dout(n1546));
    jor g0389(.dinb(n8144), .dina(n1546), .dout(n1550));
    jor g0390(.dinb(n7589), .dina(n1550), .dout(n1554));
    jor g0391(.dinb(n11036), .dina(n1554), .dout(n1558));
    jand g0392(.dinb(n1535), .dina(n1558), .dout(n1562));
    jand g0393(.dinb(n7491), .dina(n1562), .dout(n1566));
    jand g0394(.dinb(n10484), .dina(n1468), .dout(n1570));
    jnot g0395(.din(n1570), .dout(n1573));
    jnot g0396(.din(n1531), .dout(n1576));
    jand g0397(.dinb(n7550), .dina(n1576), .dout(n1580));
    jor g0398(.dinb(n10280), .dina(n1468), .dout(n1584));
    jand g0399(.dinb(n1580), .dina(n1584), .dout(n1588));
    jand g0400(.dinb(n1573), .dina(n1588), .dout(n1592));
    jor g0401(.dinb(n1566), .dina(n1592), .dout(n1596));
    jand g0402(.dinb(n8732), .dina(n431), .dout(n1600));
    jand g0403(.dinb(n8150), .dina(n1600), .dout(n1604));
    jand g0404(.dinb(n8753), .dina(n450), .dout(n1608));
    jand g0405(.dinb(n7587), .dina(n465), .dout(n1612));
    jor g0406(.dinb(n8120), .dina(n1612), .dout(n1616));
    jor g0407(.dinb(n7545), .dina(n1616), .dout(n1620));
    jand g0408(.dinb(n11225), .dina(n1620), .dout(n1624));
    jor g0409(.dinb(n8141), .dina(n1624), .dout(n1628));
    jor g0410(.dinb(n7542), .dina(n1628), .dout(n1632));
    jnot g0411(.din(n1632), .dout(n1635));
    jor g0412(.dinb(n9965), .dina(n1635), .dout(n1639));
    jnot g0413(.din(G159), .dout(n1642));
    jnot g0414(.din(n1491), .dout(n1645));
    jor g0415(.dinb(n7536), .dina(n1645), .dout(n1649));
    jxor g0416(.dinb(G58), .dina(G68), .dout(n1653));
    jor g0417(.dinb(n367), .dina(n1653), .dout(n1657));
    jand g0418(.dinb(n7790), .dina(n1476), .dout(n1661));
    jnot g0419(.din(n1661), .dout(n1664));
    jand g0420(.dinb(n7530), .dina(n1664), .dout(n1668));
    jand g0421(.dinb(n7524), .dina(n1668), .dout(n1672));
    jor g0422(.dinb(n9227), .dina(n1672), .dout(n1676));
    jnot g0423(.din(n1676), .dout(n1679));
    jand g0424(.dinb(n7511), .dina(n1516), .dout(n1683));
    jnot g0425(.din(n1683), .dout(n1686));
    jor g0426(.dinb(n7499), .dina(n1373), .dout(n1690));
    jand g0427(.dinb(n1686), .dina(n1690), .dout(n1694));
    jor g0428(.dinb(n1679), .dina(n7496), .dout(n1698));
    jor g0429(.dinb(n11084), .dina(n1632), .dout(n1702));
    jand g0430(.dinb(n1698), .dina(n1702), .dout(n1706));
    jand g0431(.dinb(n1639), .dina(n1706), .dout(n1710));
    jor g0432(.dinb(n9335), .dina(n1635), .dout(n1714));
    jnot g0433(.din(n1694), .dout(n1717));
    jand g0434(.dinb(n7520), .dina(n1717), .dout(n1721));
    jnot g0435(.din(G190), .dout(n1724));
    jor g0436(.dinb(n9215), .dina(n1632), .dout(n1728));
    jand g0437(.dinb(n1721), .dina(n1728), .dout(n1732));
    jand g0438(.dinb(n1714), .dina(n1732), .dout(n1736));
    jor g0439(.dinb(n1710), .dina(n1736), .dout(n1740));
    jor g0440(.dinb(n1596), .dina(n1740), .dout(n1744));
    jor g0441(.dinb(n1420), .dina(n1744), .dout(n1748));
    jor g0442(.dinb(n1298), .dina(n1748), .dout(n1752));
    jnot g0443(.din(n1752), .dout(n1755));
    jand g0444(.dinb(n7604), .dina(n1755), .dout(n1759));
    jnot g0445(.din(n602), .dout(n1762));
    jor g0446(.dinb(n11084), .dina(n598), .dout(n1766));
    jand g0447(.dinb(n9473), .dina(n1766), .dout(n1770));
    jand g0448(.dinb(n1762), .dina(n1770), .dout(n1774));
    jnot g0449(.din(n698), .dout(n1777));
    jor g0450(.dinb(n9332), .dina(n682), .dout(n1781));
    jand g0451(.dinb(n649), .dina(n1781), .dout(n1785));
    jand g0452(.dinb(n1777), .dina(n1785), .dout(n1789));
    jor g0453(.dinb(n1774), .dina(n1789), .dout(n1793));
    jnot g0454(.din(n767), .dout(n1796));
    jor g0455(.dinb(n9947), .dina(n763), .dout(n1800));
    jand g0456(.dinb(n904), .dina(n1800), .dout(n1804));
    jand g0457(.dinb(n1796), .dina(n1804), .dout(n1808));
    jnot g0458(.din(n870), .dout(n1811));
    jor g0459(.dinb(n10457), .dina(n854), .dout(n1815));
    jand g0460(.dinb(n828), .dina(n1815), .dout(n1819));
    jand g0461(.dinb(n1811), .dina(n1819), .dout(n1823));
    jor g0462(.dinb(n1808), .dina(n1823), .dout(n1827));
    jnot g0463(.din(n970), .dout(n1830));
    jor g0464(.dinb(n10262), .dina(n966), .dout(n1834));
    jand g0465(.dinb(n1105), .dina(n1834), .dout(n1838));
    jand g0466(.dinb(n1830), .dina(n1838), .dout(n1842));
    jor g0467(.dinb(n11084), .dina(n1052), .dout(n1846));
    jand g0468(.dinb(n9074), .dina(n1846), .dout(n1850));
    jand g0469(.dinb(n9095), .dina(n1850), .dout(n1854));
    jor g0470(.dinb(n9069), .dina(n1854), .dout(n1858));
    jor g0471(.dinb(n9212), .dina(n1858), .dout(n1862));
    jor g0472(.dinb(n9066), .dina(n1862), .dout(n1866));
    jor g0473(.dinb(n10979), .dina(n1866), .dout(n1870));
    jor g0474(.dinb(n9443), .dina(n1862), .dout(n1874));
    jor g0475(.dinb(n1823), .dina(n1117), .dout(n1878));
    jand g0476(.dinb(n9062), .dina(n1878), .dout(n1882));
    jand g0477(.dinb(n1874), .dina(n9047), .dout(n1886));
    jand g0478(.dinb(n1870), .dina(n1886), .dout(n1890));
    jor g0479(.dinb(n7451), .dina(n1890), .dout(n1894));
    jnot g0480(.din(n1894), .dout(n1897));
    jnot g0481(.din(n1592), .dout(n1900));
    jand g0482(.dinb(n1900), .dina(n7493), .dout(n1904));
    jnot g0483(.din(n1904), .dout(n1907));
    jnot g0484(.din(n1566), .dout(n1910));
    jnot g0485(.din(n1397), .dout(n1913));
    jor g0486(.dinb(n1269), .dina(n1416), .dout(n1917));
    jand g0487(.dinb(n7485), .dina(n1917), .dout(n1921));
    jor g0488(.dinb(n7487), .dina(n1921), .dout(n1925));
    jand g0489(.dinb(n7482), .dina(n1925), .dout(n1929));
    jand g0490(.dinb(n7473), .dina(n1929), .dout(n1933));
    jnot g0491(.din(n1933), .dout(n1936));
    jor g0492(.dinb(n1897), .dina(n1936), .dout(n1940));
    jand g0493(.dinb(n10877), .dina(n337), .dout(n1944));
    jand g0494(.dinb(n11978), .dina(n1944), .dout(n1948));
    jand g0495(.dinb(n10883), .dina(n1948), .dout(n1952));
    jor g0496(.dinb(n694), .dina(n9410), .dout(n1956));
    jnot g0497(.din(n1956), .dout(n1959));
    jnot g0498(.din(n522), .dout(n1962));
    jnot g0499(.din(n1952), .dout(n1965));
    jand g0500(.dinb(n1962), .dina(n9383), .dout(n1969));
    jand g0501(.dinb(n9431), .dina(n1969), .dout(n1973));
    jor g0502(.dinb(n8348), .dina(n1973), .dout(n1977));
    jand g0503(.dinb(n406), .dina(n10790), .dout(n1981));
    jxor g0504(.dinb(n545), .dina(n10764), .dout(n1985));
    jand g0505(.dinb(n11636), .dina(n1985), .dout(n1989));
    jand g0506(.dinb(n646), .dina(n10790), .dout(n1993));
    jxor g0507(.dinb(n714), .dina(n9375), .dout(n1997));
    jand g0508(.dinb(n1989), .dina(n8390), .dout(n2001));
    jor g0509(.dinb(n1977), .dina(n2001), .dout(n2005));
    jand g0510(.dinb(n12197), .dina(n140), .dout(n2009));
    jand g0511(.dinb(n240), .dina(n2009), .dout(n2013));
    jor g0512(.dinb(n1890), .dina(n10766), .dout(n2017));
    jnot g0513(.din(n545), .dout(n2020));
    jor g0514(.dinb(n2020), .dina(n1866), .dout(n2024));
    jand g0515(.dinb(n2024), .dina(n9377), .dout(n2028));
    jnot g0516(.din(n514), .dout(n2031));
    jand g0517(.dinb(n763), .dina(n966), .dout(n2035));
    jand g0518(.dinb(n2031), .dina(n9045), .dout(n2039));
    jand g0519(.dinb(n9449), .dina(n2039), .dout(n2043));
    jand g0520(.dinb(n11000), .dina(n854), .dout(n2047));
    jand g0521(.dinb(n1052), .dina(n2047), .dout(n2051));
    jand g0522(.dinb(n11108), .dina(n2051), .dout(n2055));
    jand g0523(.dinb(n9497), .dina(n2055), .dout(n2059));
    jor g0524(.dinb(n9408), .dina(n2059), .dout(n2063));
    jor g0525(.dinb(n2043), .dina(n2063), .dout(n2067));
    jand g0526(.dinb(n11676), .dina(n2067), .dout(n2071));
    jnot g0527(.din(n2071), .dout(n2074));
    jor g0528(.dinb(n2028), .dina(n9018), .dout(n2078));
    jand g0529(.dinb(n2017), .dina(n2078), .dout(n2082));
    jnot g0530(.din(n2082), .dout(n2085));
    jand g0531(.dinb(n11279), .dina(n2085), .dout(n2089));
    jnot g0532(.din(n2009), .dout(n2092));
    jand g0533(.dinb(n11411), .dina(n779), .dout(n2096));
    jand g0534(.dinb(n12134), .dina(n2096), .dout(n2100));
    jand g0535(.dinb(n2092), .dina(n2100), .dout(n2104));
    jor g0536(.dinb(n2089), .dina(n6492), .dout(n2108));
    jor g0537(.dinb(n6450), .dina(n2108), .dout(n2112));
    jand g0538(.dinb(G13), .dina(G45), .dout(n2116));
    jand g0539(.dinb(n367), .dina(n2116), .dout(n2120));
    jor g0540(.dinb(n11987), .dina(n2120), .dout(n2124));
    jnot g0541(.din(n2124), .dout(n2127));
    jand g0542(.dinb(n2092), .dina(n11964), .dout(n2131));
    jnot g0543(.din(n2131), .dout(n2134));
    jxor g0544(.dinb(n11633), .dina(n1985), .dout(n2138));
    jand g0545(.dinb(n10752), .dina(n2138), .dout(n2142));
    jand g0546(.dinb(n132), .dina(n374), .dout(n2146));
    jand g0547(.dinb(n11975), .dina(n2146), .dout(n2150));
    jnot g0548(.din(n2150), .dout(n2153));
    jor g0549(.dinb(n1985), .dina(n10550), .dout(n2157));
    jand g0550(.dinb(n10508), .dina(n1724), .dout(n2161));
    jnot g0551(.din(n2161), .dout(n2164));
    jand g0552(.dinb(G20), .dina(G200), .dout(n2168));
    jnot g0553(.din(n2168), .dout(n2171));
    jand g0554(.dinb(G20), .dina(G179), .dout(n2175));
    jnot g0555(.din(n2175), .dout(n2178));
    jand g0556(.dinb(n2171), .dina(n2178), .dout(n2182));
    jand g0557(.dinb(n2164), .dina(n2182), .dout(n2186));
    jand g0558(.dinb(n10511), .dina(n2186), .dout(n2190));
    jnot g0559(.din(n2190), .dout(n2193));
    jand g0560(.dinb(n510), .dina(n2168), .dout(n2197));
    jand g0561(.dinb(n10478), .dina(n2197), .dout(n2201));
    jand g0562(.dinb(n10403), .dina(n2201), .dout(n2205));
    jnot g0563(.din(n2205), .dout(n2208));
    jand g0564(.dinb(n2193), .dina(n10392), .dout(n2212));
    jand g0565(.dinb(n1272), .dina(n2175), .dout(n2216));
    jand g0566(.dinb(n10454), .dina(n2216), .dout(n2220));
    jand g0567(.dinb(n10346), .dina(n2220), .dout(n2224));
    jand g0568(.dinb(n10448), .dina(n2182), .dout(n2228));
    jand g0569(.dinb(n10232), .dina(n2228), .dout(n2232));
    jor g0570(.dinb(n10221), .dina(n2232), .dout(n2236));
    jor g0571(.dinb(n10370), .dina(n2236), .dout(n2240));
    jnot g0572(.din(n2240), .dout(n2243));
    jand g0573(.dinb(n10218), .dina(n2243), .dout(n2247));
    jand g0574(.dinb(n10928), .dina(n2216), .dout(n2251));
    jand g0575(.dinb(n10190), .dina(n2251), .dout(n2255));
    jand g0576(.dinb(n10451), .dina(n2197), .dout(n2259));
    jand g0577(.dinb(n10172), .dina(n2259), .dout(n2263));
    jand g0578(.dinb(n10421), .dina(n2175), .dout(n2267));
    jand g0579(.dinb(n10928), .dina(n2267), .dout(n2271));
    jand g0580(.dinb(n10148), .dina(n2271), .dout(n2275));
    jand g0581(.dinb(n10475), .dina(n2267), .dout(n2279));
    jand g0582(.dinb(n10133), .dina(n2279), .dout(n2283));
    jor g0583(.dinb(n2275), .dina(n2283), .dout(n2287));
    jor g0584(.dinb(n10169), .dina(n2287), .dout(n2291));
    jor g0585(.dinb(n10125), .dina(n2291), .dout(n2295));
    jnot g0586(.din(n2295), .dout(n2298));
    jand g0587(.dinb(n2247), .dina(n10119), .dout(n2302));
    jnot g0588(.din(n2302), .dout(n2305));
    jand g0589(.dinb(n10116), .dina(n2251), .dout(n2309));
    jand g0590(.dinb(n11165), .dina(n2201), .dout(n2313));
    jand g0591(.dinb(n10076), .dina(n2186), .dout(n2317));
    jor g0592(.dinb(n10074), .dina(n2317), .dout(n2321));
    jand g0593(.dinb(n10071), .dina(n2271), .dout(n2325));
    jor g0594(.dinb(n2321), .dina(n10059), .dout(n2329));
    jand g0595(.dinb(n10053), .dina(n2228), .dout(n2333));
    jor g0596(.dinb(n10712), .dina(n2333), .dout(n2337));
    jand g0597(.dinb(n10041), .dina(n2220), .dout(n2341));
    jand g0598(.dinb(n10029), .dina(n2279), .dout(n2345));
    jor g0599(.dinb(n2341), .dina(n2345), .dout(n2349));
    jand g0600(.dinb(n11495), .dina(n2259), .dout(n2353));
    jor g0601(.dinb(n2349), .dina(n10017), .dout(n2357));
    jor g0602(.dinb(n2337), .dina(n2357), .dout(n2361));
    jor g0603(.dinb(n2329), .dina(n2361), .dout(n2365));
    jor g0604(.dinb(n10014), .dina(n2365), .dout(n2369));
    jand g0605(.dinb(n2305), .dina(n10002), .dout(n2373));
    jand g0606(.dinb(n11360), .dina(n322), .dout(n2377));
    jor g0607(.dinb(n1224), .dina(n2377), .dout(n2381));
    jnot g0608(.din(n2381), .dout(n2384));
    jor g0609(.dinb(n2373), .dina(n9887), .dout(n2388));
    jand g0610(.dinb(n2153), .dina(n2384), .dout(n2392));
    jor g0611(.dinb(n9851), .dina(n302), .dout(n2396));
    jand g0612(.dinb(n11561), .dina(n140), .dout(n2400));
    jnot g0613(.din(n2400), .dout(n2403));
    jand g0614(.dinb(n9866), .dina(n240), .dout(n2407));
    jor g0615(.dinb(n2403), .dina(n2407), .dout(n2411));
    jnot g0616(.din(n2411), .dout(n2414));
    jand g0617(.dinb(n9744), .dina(n2414), .dout(n2418));
    jnot g0618(.din(n140), .dout(n2421));
    jand g0619(.dinb(n11402), .dina(n2421), .dout(n2425));
    jand g0620(.dinb(n10724), .dina(n140), .dout(n2429));
    jand g0621(.dinb(n9644), .dina(n2429), .dout(n2433));
    jor g0622(.dinb(n2425), .dina(n2433), .dout(n2437));
    jor g0623(.dinb(n2418), .dina(n9606), .dout(n2441));
    jand g0624(.dinb(n9875), .dina(n2441), .dout(n2445));
    jnot g0625(.din(n2445), .dout(n2448));
    jand g0626(.dinb(n2388), .dina(n9600), .dout(n2452));
    jand g0627(.dinb(n2157), .dina(n9594), .dout(n2456));
    jand g0628(.dinb(n11678), .dina(n2456), .dout(n2460));
    jor g0629(.dinb(n9591), .dina(n2460), .dout(n2464));
    jand g0630(.dinb(n1254), .dina(n10838), .dout(n2468));
    jxor g0631(.dinb(n1295), .dina(n8064), .dout(n2472));
    jnot g0632(.din(n2472), .dout(n2475));
    jand g0633(.dinb(n10637), .dina(n2475), .dout(n2479));
    jnot g0634(.din(n2479), .dout(n2482));
    jand g0635(.dinb(n8021), .dina(n2279), .dout(n2486));
    jand g0636(.dinb(n8472), .dina(n2271), .dout(n2490));
    jand g0637(.dinb(n10142), .dina(n2201), .dout(n2494));
    jor g0638(.dinb(n2490), .dina(n2494), .dout(n2498));
    jand g0639(.dinb(n8457), .dina(n2251), .dout(n2502));
    jor g0640(.dinb(n2498), .dina(n8019), .dout(n2506));
    jor g0641(.dinb(n8016), .dina(n2506), .dout(n2510));
    jand g0642(.dinb(n10223), .dina(n2220), .dout(n2514));
    jand g0643(.dinb(n8000), .dina(n2228), .dout(n2518));
    jor g0644(.dinb(n7998), .dina(n2518), .dout(n2522));
    jand g0645(.dinb(n8438), .dina(n2186), .dout(n2526));
    jand g0646(.dinb(n10127), .dina(n2259), .dout(n2530));
    jor g0647(.dinb(n2526), .dina(n7995), .dout(n2534));
    jor g0648(.dinb(n9788), .dina(n2534), .dout(n2538));
    jor g0649(.dinb(n7980), .dina(n2538), .dout(n2542));
    jor g0650(.dinb(n7977), .dina(n2542), .dout(n2546));
    jand g0651(.dinb(n11486), .dina(n2279), .dout(n2550));
    jand g0652(.dinb(n10031), .dina(n2228), .dout(n2554));
    jor g0653(.dinb(n7974), .dina(n2554), .dout(n2558));
    jand g0654(.dinb(n10181), .dina(n2201), .dout(n2562));
    jor g0655(.dinb(n2190), .dina(n7971), .dout(n2566));
    jor g0656(.dinb(n2558), .dina(n2566), .dout(n2570));
    jand g0657(.dinb(n10097), .dina(n2251), .dout(n2574));
    jand g0658(.dinb(n11534), .dina(n2220), .dout(n2578));
    jor g0659(.dinb(n2574), .dina(n2578), .dout(n2582));
    jand g0660(.dinb(n11156), .dina(n2271), .dout(n2586));
    jand g0661(.dinb(n10394), .dina(n2259), .dout(n2590));
    jor g0662(.dinb(n2586), .dina(n2590), .dout(n2594));
    jor g0663(.dinb(n2582), .dina(n2594), .dout(n2598));
    jor g0664(.dinb(n2570), .dina(n7968), .dout(n2602));
    jor g0665(.dinb(n9629), .dina(n2602), .dout(n2606));
    jand g0666(.dinb(n2546), .dina(n2606), .dout(n2610));
    jor g0667(.dinb(n8516), .dina(n2610), .dout(n2614));
    jnot g0668(.din(n2146), .dout(n2617));
    jand g0669(.dinb(n7899), .dina(n2384), .dout(n2621));
    jand g0670(.dinb(n9128), .dina(n2621), .dout(n2625));
    jnot g0671(.din(n2625), .dout(n2628));
    jand g0672(.dinb(n2614), .dina(n7896), .dout(n2632));
    jand g0673(.dinb(n8585), .dina(n2632), .dout(n2636));
    jand g0674(.dinb(n2482), .dina(n7884), .dout(n2640));
    jnot g0675(.din(n2640), .dout(n2643));
    jor g0676(.dinb(n7865), .dina(n2017), .dout(n2647));
    jand g0677(.dinb(n9428), .dina(n1129), .dout(n2651));
    jand g0678(.dinb(n9341), .dina(n1125), .dout(n2655));
    jnot g0679(.din(n1882), .dout(n2658));
    jor g0680(.dinb(n2655), .dina(n7860), .dout(n2662));
    jor g0681(.dinb(n2651), .dina(n2662), .dout(n2666));
    jand g0682(.dinb(n2666), .dina(n9026), .dout(n2670));
    jor g0683(.dinb(n2670), .dina(n8030), .dout(n2674));
    jand g0684(.dinb(n2647), .dina(n2674), .dout(n2678));
    jxor g0685(.dinb(n9011), .dina(n2678), .dout(n2682));
    jor g0686(.dinb(n8549), .dina(n2682), .dout(n2686));
    jand g0687(.dinb(n7857), .dina(n2686), .dout(n2690));
    jnot g0688(.din(n2690), .dout(n2693));
    jnot g0689(.din(n136), .dout(n2696));
    jand g0690(.dinb(n2696), .dina(n6617), .dout(n2700));
    jnot g0691(.din(n1948), .dout(n2703));
    jand g0692(.dinb(n1710), .dina(n7230), .dout(n2707));
    jand g0693(.dinb(n1698), .dina(n10859), .dout(n2711));
    jxor g0694(.dinb(n1740), .dina(n7422), .dout(n2715));
    jnot g0695(.din(n2715), .dout(n2718));
    jor g0696(.dinb(n1921), .dina(n8069), .dout(n2722));
    jnot g0697(.din(n2722), .dout(n2725));
    jand g0698(.dinb(n1385), .dina(n8066), .dout(n2729));
    jxor g0699(.dinb(n1420), .dina(n7767), .dout(n2733));
    jnot g0700(.din(n2733), .dout(n2736));
    jand g0701(.dinb(n8048), .dina(n2736), .dout(n2740));
    jand g0702(.dinb(n2670), .dina(n7274), .dout(n2744));
    jor g0703(.dinb(n7272), .dina(n2744), .dout(n2748));
    jand g0704(.dinb(n7205), .dina(n2748), .dout(n2752));
    jor g0705(.dinb(n7203), .dina(n2752), .dout(n2756));
    jand g0706(.dinb(n7302), .dina(n2740), .dout(n2760));
    jxor g0707(.dinb(n7460), .dina(n2760), .dout(n2764));
    jor g0708(.dinb(n9008), .dina(n2764), .dout(n2768));
    jor g0709(.dinb(n1894), .dina(n8618), .dout(n2772));
    jand g0710(.dinb(n7466), .dina(n2772), .dout(n2776));
    jxor g0711(.dinb(n2768), .dina(n2776), .dout(n2780));
    jxor g0712(.dinb(n2756), .dina(n6615), .dout(n2784));
    jand g0713(.dinb(n6612), .dina(n2784), .dout(n2788));
    jor g0714(.dinb(n80), .dina(n83), .dout(n2792));
    jand g0715(.dinb(n10364), .dina(n2792), .dout(n2796));
    jor g0716(.dinb(n8684), .dina(n2796), .dout(n2800));
    jand g0717(.dinb(G50), .dina(G58), .dout(n2804));
    jor g0718(.dinb(n10139), .dina(n2804), .dout(n2808));
    jand g0719(.dinb(n136), .dina(n2808), .dout(n2812));
    jand g0720(.dinb(n2800), .dina(n6558), .dout(n2816));
    jand g0721(.dinb(n247), .dina(n9170), .dout(n2820));
    jand g0722(.dinb(n11624), .dina(n2820), .dout(n2824));
    jor g0723(.dinb(n2816), .dina(n6546), .dout(n2828));
    jor g0724(.dinb(n2788), .dina(n6543), .dout(n2832));
    jand g0725(.dinb(n904), .dina(n10829), .dout(n2836));
    jxor g0726(.dinb(n1827), .dina(n8616), .dout(n2840));
    jand g0727(.dinb(n10610), .dina(n2840), .dout(n2844));
    jnot g0728(.din(n2844), .dout(n2847));
    jand g0729(.dinb(n8543), .dina(n2400), .dout(n2851));
    jnot g0730(.din(n2392), .dout(n2854));
    jand g0731(.dinb(n8891), .dina(n2421), .dout(n2858));
    jor g0732(.dinb(n2854), .dina(n8541), .dout(n2862));
    jor g0733(.dinb(n8538), .dina(n2862), .dout(n2866));
    jand g0734(.dinb(n11708), .dina(n2866), .dout(n2870));
    jand g0735(.dinb(n11174), .dina(n2251), .dout(n2874));
    jand g0736(.dinb(n11513), .dina(n2220), .dout(n2878));
    jor g0737(.dinb(n2874), .dina(n2878), .dout(n2882));
    jand g0738(.dinb(n10041), .dina(n2271), .dout(n2886));
    jand g0739(.dinb(n11624), .dina(n2201), .dout(n2890));
    jor g0740(.dinb(n2886), .dina(n2890), .dout(n2894));
    jand g0741(.dinb(n10097), .dina(n2279), .dout(n2898));
    jand g0742(.dinb(n10019), .dina(n2228), .dout(n2902));
    jor g0743(.dinb(n8493), .dina(n2902), .dout(n2906));
    jand g0744(.dinb(n8489), .dina(n2186), .dout(n2910));
    jand g0745(.dinb(n11447), .dina(n2259), .dout(n2914));
    jor g0746(.dinb(n2910), .dina(n8921), .dout(n2918));
    jor g0747(.dinb(n2906), .dina(n2918), .dout(n2922));
    jor g0748(.dinb(n8487), .dina(n2922), .dout(n2926));
    jor g0749(.dinb(n8481), .dina(n2926), .dout(n2930));
    jand g0750(.dinb(n9770), .dina(n2930), .dout(n2934));
    jand g0751(.dinb(n8870), .dina(n2220), .dout(n2938));
    jand g0752(.dinb(n8462), .dina(n2228), .dout(n2942));
    jor g0753(.dinb(n8460), .dina(n2942), .dout(n2946));
    jand g0754(.dinb(n8457), .dina(n2271), .dout(n2950));
    jand g0755(.dinb(n10253), .dina(n2279), .dout(n2954));
    jor g0756(.dinb(n2950), .dina(n2954), .dout(n2958));
    jand g0757(.dinb(n8429), .dina(n2201), .dout(n2962));
    jand g0758(.dinb(n8909), .dina(n2186), .dout(n2966));
    jor g0759(.dinb(n8427), .dina(n2966), .dout(n2970));
    jand g0760(.dinb(n8852), .dina(n2251), .dout(n2974));
    jand g0761(.dinb(n8885), .dina(n2259), .dout(n2978));
    jor g0762(.dinb(n2974), .dina(n2978), .dout(n2982));
    jor g0763(.dinb(n2970), .dina(n8421), .dout(n2986));
    jor g0764(.dinb(n8418), .dina(n2986), .dout(n2990));
    jor g0765(.dinb(n8412), .dina(n2990), .dout(n2994));
    jand g0766(.dinb(n9611), .dina(n2994), .dout(n2998));
    jor g0767(.dinb(n2934), .dina(n2998), .dout(n3002));
    jor g0768(.dinb(n8495), .dina(n3002), .dout(n3006));
    jand g0769(.dinb(n8406), .dina(n3006), .dout(n3010));
    jand g0770(.dinb(n2847), .dina(n8397), .dout(n3014));
    jnot g0771(.din(n3014), .dout(n3017));
    jand g0772(.dinb(n1024), .dina(n10829), .dout(n3021));
    jxor g0773(.dinb(n1858), .dina(n8388), .dout(n3025));
    jnot g0774(.din(n3025), .dout(n3028));
    jand g0775(.dinb(n2001), .dina(n8367), .dout(n3032));
    jand g0776(.dinb(n1854), .dina(n9408), .dout(n3036));
    jand g0777(.dinb(n8354), .dina(n1997), .dout(n3040));
    jand g0778(.dinb(n1969), .dina(n3040), .dout(n3044));
    jand g0779(.dinb(n8357), .dina(n1959), .dout(n3048));
    jor g0780(.dinb(n3044), .dina(n8346), .dout(n3052));
    jor g0781(.dinb(n8343), .dina(n3052), .dout(n3056));
    jxor g0782(.dinb(n8597), .dina(n3056), .dout(n3060));
    jxor g0783(.dinb(n8331), .dina(n3060), .dout(n3064));
    jor g0784(.dinb(n11825), .dina(n3064), .dout(n3068));
    jnot g0785(.din(n1973), .dout(n3071));
    jor g0786(.dinb(n1969), .dina(n9365), .dout(n3075));
    jand g0787(.dinb(n3071), .dina(n9363), .dout(n3079));
    jxor g0788(.dinb(n9572), .dina(n3079), .dout(n3083));
    jnot g0789(.din(n3083), .dout(n3086));
    jxor g0790(.dinb(n1977), .dina(n2001), .dout(n3090));
    jxor g0791(.dinb(n8369), .dina(n3090), .dout(n3094));
    jor g0792(.dinb(n3086), .dina(n8327), .dout(n3098));
    jand g0793(.dinb(n9002), .dina(n3098), .dout(n3102));
    jor g0794(.dinb(n11996), .dina(n3064), .dout(n3106));
    jor g0795(.dinb(n3102), .dina(n8316), .dout(n3110));
    jand g0796(.dinb(n8313), .dina(n3110), .dout(n3114));
    jand g0797(.dinb(n8307), .dina(n3114), .dout(n3118));
    jnot g0798(.din(n3118), .dout(n3121));
    jor g0799(.dinb(n12038), .dina(n2085), .dout(n3125));
    jand g0800(.dinb(n9359), .dina(n3125), .dout(n3129));
    jand g0801(.dinb(n2082), .dina(n3083), .dout(n3133));
    jand g0802(.dinb(n11783), .dina(n3133), .dout(n3137));
    jor g0803(.dinb(n8975), .dina(n3137), .dout(n3141));
    jor g0804(.dinb(n3129), .dina(n3141), .dout(n3145));
    jor g0805(.dinb(n1997), .dina(n10523), .dout(n3149));
    jand g0806(.dinb(n8942), .dina(n2279), .dout(n3153));
    jand g0807(.dinb(n8900), .dina(n2220), .dout(n3157));
    jor g0808(.dinb(n2914), .dina(n3157), .dout(n3161));
    jor g0809(.dinb(n9803), .dina(n3161), .dout(n3165));
    jor g0810(.dinb(n8898), .dina(n3165), .dout(n3169));
    jnot g0811(.din(n3169), .dout(n3172));
    jand g0812(.dinb(n8888), .dina(n2186), .dout(n3176));
    jnot g0813(.din(n3176), .dout(n3179));
    jand g0814(.dinb(n8882), .dina(n2201), .dout(n3183));
    jnot g0815(.din(n3183), .dout(n3186));
    jand g0816(.dinb(n3179), .dina(n8879), .dout(n3190));
    jand g0817(.dinb(n8861), .dina(n2251), .dout(n3194));
    jand g0818(.dinb(n8846), .dina(n2228), .dout(n3198));
    jor g0819(.dinb(n8844), .dina(n3198), .dout(n3202));
    jand g0820(.dinb(n10253), .dina(n2271), .dout(n3206));
    jor g0821(.dinb(n3202), .dina(n8841), .dout(n3210));
    jnot g0822(.din(n3210), .dout(n3213));
    jand g0823(.dinb(n8835), .dina(n3213), .dout(n3217));
    jand g0824(.dinb(n8832), .dina(n3217), .dout(n3221));
    jnot g0825(.din(n3221), .dout(n3224));
    jand g0826(.dinb(n10041), .dina(n2279), .dout(n3228));
    jand g0827(.dinb(n10097), .dina(n2201), .dout(n3232));
    jand g0828(.dinb(n8828), .dina(n2186), .dout(n3236));
    jor g0829(.dinb(n8826), .dina(n3236), .dout(n3240));
    jand g0830(.dinb(n10116), .dina(n2271), .dout(n3244));
    jand g0831(.dinb(n10061), .dina(n2228), .dout(n3248));
    jor g0832(.dinb(n8823), .dina(n3248), .dout(n3252));
    jor g0833(.dinb(n3240), .dina(n3252), .dout(n3256));
    jand g0834(.dinb(n11174), .dina(n2220), .dout(n3260));
    jand g0835(.dinb(n11624), .dina(n2259), .dout(n3264));
    jor g0836(.dinb(n3260), .dina(n3264), .dout(n3268));
    jand g0837(.dinb(n10029), .dina(n2251), .dout(n3272));
    jor g0838(.dinb(n3268), .dina(n8799), .dout(n3276));
    jor g0839(.dinb(n8816), .dina(n3276), .dout(n3280));
    jor g0840(.dinb(n3256), .dina(n3280), .dout(n3284));
    jor g0841(.dinb(n8796), .dina(n3284), .dout(n3288));
    jand g0842(.dinb(n3224), .dina(n8784), .dout(n3292));
    jor g0843(.dinb(n8954), .dina(n3292), .dout(n3296));
    jand g0844(.dinb(n9647), .dina(n2421), .dout(n3300));
    jnot g0845(.din(n3300), .dout(n3303));
    jnot g0846(.din(n2096), .dout(n3306));
    jand g0847(.dinb(n3306), .dina(n9608), .dout(n3310));
    jnot g0848(.din(n3310), .dout(n3313));
    jand g0849(.dinb(n11966), .dina(n286), .dout(n3317));
    jor g0850(.dinb(n2403), .dina(n8718), .dout(n3321));
    jand g0851(.dinb(n3313), .dina(n8715), .dout(n3325));
    jand g0852(.dinb(G68), .dina(G77), .dout(n3329));
    jnot g0853(.din(n3329), .dout(n3332));
    jand g0854(.dinb(n77), .dina(n10214), .dout(n3336));
    jand g0855(.dinb(n3332), .dina(n3336), .dout(n3340));
    jand g0856(.dinb(n2096), .dina(n8682), .dout(n3344));
    jand g0857(.dinb(n9854), .dina(n3344), .dout(n3348));
    jor g0858(.dinb(n3325), .dina(n8679), .dout(n3352));
    jand g0859(.dinb(n8673), .dina(n3352), .dout(n3356));
    jor g0860(.dinb(n8768), .dina(n3356), .dout(n3360));
    jand g0861(.dinb(n3296), .dina(n8664), .dout(n3364));
    jand g0862(.dinb(n3149), .dina(n3364), .dout(n3368));
    jand g0863(.dinb(n8963), .dina(n3368), .dout(n3372));
    jnot g0864(.din(n3372), .dout(n3375));
    jand g0865(.dinb(n3145), .dina(n8658), .dout(n3379));
    jnot g0866(.din(n3379), .dout(n3382));
    jnot g0867(.din(n3094), .dout(n3385));
    jnot g0868(.din(n3133), .dout(n3388));
    jor g0869(.dinb(n8286), .dina(n3388), .dout(n3392));
    jor g0870(.dinb(n9353), .dina(n3392), .dout(n3396));
    jor g0871(.dinb(n8318), .dina(n3141), .dout(n3400));
    jand g0872(.dinb(n10580), .dina(n3025), .dout(n3404));
    jnot g0873(.din(n3404), .dout(n3407));
    jand g0874(.dinb(n8924), .dina(n2421), .dout(n3411));
    jand g0875(.dinb(n8279), .dina(n2400), .dout(n3415));
    jor g0876(.dinb(n2854), .dina(n8277), .dout(n3419));
    jor g0877(.dinb(n8274), .dina(n3419), .dout(n3423));
    jand g0878(.dinb(n8261), .dina(n2279), .dout(n3427));
    jand g0879(.dinb(n8936), .dina(n2220), .dout(n3431));
    jor g0880(.dinb(n3427), .dina(n3431), .dout(n3435));
    jand g0881(.dinb(n10253), .dina(n2251), .dout(n3439));
    jand g0882(.dinb(n9830), .dina(n2201), .dout(n3443));
    jor g0883(.dinb(n3439), .dina(n3443), .dout(n3447));
    jand g0884(.dinb(n8852), .dina(n2271), .dout(n3451));
    jor g0885(.dinb(n2590), .dina(n3451), .dout(n3455));
    jand g0886(.dinb(n8249), .dina(n2228), .dout(n3459));
    jand g0887(.dinb(n9815), .dina(n2186), .dout(n3463));
    jor g0888(.dinb(n3459), .dina(n3463), .dout(n3467));
    jor g0889(.dinb(n8238), .dina(n3467), .dout(n3471));
    jor g0890(.dinb(n8235), .dina(n3471), .dout(n3475));
    jor g0891(.dinb(n8229), .dina(n3475), .dout(n3479));
    jand g0892(.dinb(n8801), .dina(n3479), .dout(n3483));
    jand g0893(.dinb(n10088), .dina(n2220), .dout(n3487));
    jand g0894(.dinb(n10106), .dina(n2228), .dout(n3491));
    jor g0895(.dinb(n8217), .dina(n3491), .dout(n3495));
    jand g0896(.dinb(n10041), .dina(n2251), .dout(n3499));
    jand g0897(.dinb(n10029), .dina(n2271), .dout(n3503));
    jor g0898(.dinb(n3499), .dina(n3503), .dout(n3507));
    jand g0899(.dinb(n11174), .dina(n2279), .dout(n3511));
    jor g0900(.dinb(n2263), .dina(n3511), .dout(n3515));
    jor g0901(.dinb(n3507), .dina(n3515), .dout(n3519));
    jand g0902(.dinb(n11513), .dina(n2201), .dout(n3523));
    jand g0903(.dinb(n8213), .dina(n2186), .dout(n3527));
    jor g0904(.dinb(n8211), .dina(n3527), .dout(n3531));
    jor g0905(.dinb(n3519), .dina(n3531), .dout(n3535));
    jor g0906(.dinb(n8208), .dina(n3535), .dout(n3539));
    jand g0907(.dinb(n8927), .dina(n3539), .dout(n3543));
    jor g0908(.dinb(n9932), .dina(n3543), .dout(n3547));
    jor g0909(.dinb(n3483), .dina(n3547), .dout(n3551));
    jand g0910(.dinb(n11768), .dina(n3551), .dout(n3555));
    jand g0911(.dinb(n8205), .dina(n3555), .dout(n3559));
    jand g0912(.dinb(n3407), .dina(n8193), .dout(n3563));
    jnot g0913(.din(n3563), .dout(n3566));
    jand g0914(.dinb(n3400), .dina(n8187), .dout(n3570));
    jand g0915(.dinb(n8172), .dina(n3570), .dout(n3574));
    jnot g0916(.din(n3574), .dout(n3577));
    jand g0917(.dinb(n7934), .dina(n2715), .dout(n3581));
    jnot g0918(.din(n3581), .dout(n3584));
    jand g0919(.dinb(n7704), .dina(n2271), .dout(n3588));
    jand g0920(.dinb(n7364), .dina(n2228), .dout(n3592));
    jor g0921(.dinb(n7362), .dina(n3592), .dout(n3596));
    jand g0922(.dinb(n8252), .dina(n2259), .dout(n3600));
    jand g0923(.dinb(n8472), .dina(n2279), .dout(n3604));
    jor g0924(.dinb(n3600), .dina(n3604), .dout(n3608));
    jor g0925(.dinb(n9803), .dina(n3608), .dout(n3612));
    jor g0926(.dinb(n3596), .dina(n3612), .dout(n3616));
    jand g0927(.dinb(n8457), .dina(n2220), .dout(n3620));
    jand g0928(.dinb(n8849), .dina(n2201), .dout(n3624));
    jand g0929(.dinb(n7733), .dina(n2186), .dout(n3628));
    jand g0930(.dinb(n8010), .dina(n2251), .dout(n3632));
    jor g0931(.dinb(n3628), .dina(n7359), .dout(n3636));
    jor g0932(.dinb(n7356), .dina(n3636), .dout(n3640));
    jor g0933(.dinb(n7350), .dina(n3640), .dout(n3644));
    jor g0934(.dinb(n7341), .dina(n3644), .dout(n3648));
    jand g0935(.dinb(n11504), .dina(n2271), .dout(n3652));
    jand g0936(.dinb(n11447), .dina(n2220), .dout(n3656));
    jor g0937(.dinb(n11468), .dina(n3656), .dout(n3660));
    jor g0938(.dinb(n7338), .dina(n3660), .dout(n3664));
    jand g0939(.dinb(n11615), .dina(n2251), .dout(n3668));
    jand g0940(.dinb(n8219), .dina(n2228), .dout(n3672));
    jor g0941(.dinb(n7335), .dina(n3672), .dout(n3676));
    jand g0942(.dinb(n10181), .dina(n2279), .dout(n3680));
    jor g0943(.dinb(n2205), .dina(n3680), .dout(n3684));
    jor g0944(.dinb(n3676), .dina(n7332), .dout(n3688));
    jor g0945(.dinb(n7329), .dina(n3688), .dout(n3692));
    jor g0946(.dinb(n8240), .dina(n3692), .dout(n3696));
    jor g0947(.dinb(n7982), .dina(n3696), .dout(n3700));
    jand g0948(.dinb(n7326), .dina(n3700), .dout(n3704));
    jor g0949(.dinb(n8948), .dina(n3704), .dout(n3708));
    jand g0950(.dinb(n9758), .dina(n2621), .dout(n3712));
    jnot g0951(.din(n3712), .dout(n3715));
    jand g0952(.dinb(n3708), .dina(n7323), .dout(n3719));
    jand g0953(.dinb(n11747), .dina(n3719), .dout(n3723));
    jand g0954(.dinb(n3584), .dina(n7308), .dout(n3727));
    jnot g0955(.din(n3727), .dout(n3730));
    jor g0956(.dinb(n7454), .dina(n2078), .dout(n3734));
    jand g0957(.dinb(n2776), .dina(n7449), .dout(n3738));
    jnot g0958(.din(n1269), .dout(n3741));
    jand g0959(.dinb(n3741), .dina(n9389), .dout(n3745));
    jnot g0960(.din(n3745), .dout(n3748));
    jand g0961(.dinb(n2647), .dina(n7635), .dout(n3752));
    jor g0962(.dinb(n1133), .dina(n10799), .dout(n3756));
    jand g0963(.dinb(n3756), .dina(n9020), .dout(n3760));
    jand g0964(.dinb(n3760), .dina(n8039), .dout(n3764));
    jxor g0965(.dinb(n7616), .dina(n3764), .dout(n3768));
    jxor g0966(.dinb(n3752), .dina(n3768), .dout(n3772));
    jand g0967(.dinb(n3738), .dina(n3772), .dout(n3776));
    jor g0968(.dinb(n9347), .dina(n3776), .dout(n3780));
    jand g0969(.dinb(n11912), .dina(n3780), .dout(n3784));
    jor g0970(.dinb(n2078), .dina(n8024), .dout(n3788));
    jor g0971(.dinb(n7745), .dina(n3788), .dout(n3792));
    jxor g0972(.dinb(n7289), .dina(n2748), .dout(n3796));
    jxor g0973(.dinb(n7304), .dina(n3796), .dout(n3800));
    jor g0974(.dinb(n3784), .dina(n7262), .dout(n3804));
    jnot g0975(.din(n3776), .dout(n3807));
    jnot g0976(.din(n3792), .dout(n3810));
    jxor g0977(.dinb(n3810), .dina(n3796), .dout(n3814));
    jor g0978(.dinb(n12080), .dina(n3814), .dout(n3818));
    jor g0979(.dinb(n3807), .dina(n3818), .dout(n3822));
    jand g0980(.dinb(n3804), .dina(n7260), .dout(n3826));
    jand g0981(.dinb(n7257), .dina(n3826), .dout(n3830));
    jnot g0982(.din(n3830), .dout(n3833));
    jxor g0983(.dinb(n7607), .dina(n3764), .dout(n3837));
    jxor g0984(.dinb(n3752), .dina(n3837), .dout(n3841));
    jor g0985(.dinb(n7602), .dina(n3800), .dout(n3845));
    jand g0986(.dinb(n11867), .dina(n3738), .dout(n3849));
    jand g0987(.dinb(n3845), .dina(n7233), .dout(n3853));
    jand g0988(.dinb(n7277), .dina(n3810), .dout(n3857));
    jand g0989(.dinb(n1535), .dina(n10844), .dout(n3861));
    jxor g0990(.dinb(n1596), .dina(n7179), .dout(n3865));
    jxor g0991(.dinb(n2756), .dina(n7151), .dout(n3869));
    jxor g0992(.dinb(n7149), .dina(n3869), .dout(n3873));
    jor g0993(.dinb(n3853), .dina(n3873), .dout(n3877));
    jor g0994(.dinb(n7385), .dina(n3877), .dout(n3881));
    jand g0995(.dinb(n7901), .dina(n3865), .dout(n3885));
    jnot g0996(.din(n3885), .dout(n3888));
    jand g0997(.dinb(G41), .dina(G50), .dout(n3892));
    jor g0998(.dinb(n2384), .dina(n7146), .dout(n3896));
    jand g0999(.dinb(n8472), .dina(n2220), .dout(n3900));
    jand g1000(.dinb(n8457), .dina(n2201), .dout(n3904));
    jand g1001(.dinb(n7374), .dina(n2271), .dout(n3908));
    jor g1002(.dinb(n3904), .dina(n3908), .dout(n3912));
    jor g1003(.dinb(n7137), .dina(n3912), .dout(n3916));
    jand g1004(.dinb(n7134), .dina(n2228), .dout(n3920));
    jand g1005(.dinb(n7730), .dina(n2186), .dout(n3924));
    jand g1006(.dinb(n7704), .dina(n2251), .dout(n3928));
    jor g1007(.dinb(n3924), .dina(n7122), .dout(n3932));
    jor g1008(.dinb(n7119), .dina(n3932), .dout(n3936));
    jand g1009(.dinb(n10244), .dina(n2259), .dout(n3940));
    jand g1010(.dinb(n8010), .dina(n2279), .dout(n3944));
    jor g1011(.dinb(n3940), .dina(n3944), .dout(n3948));
    jor g1012(.dinb(n9797), .dina(n3948), .dout(n3952));
    jor g1013(.dinb(n3936), .dina(n7116), .dout(n3956));
    jor g1014(.dinb(n7113), .dina(n3956), .dout(n3960));
    jand g1015(.dinb(n11438), .dina(n2279), .dout(n3964));
    jand g1016(.dinb(n9683), .dina(n2251), .dout(n3968));
    jor g1017(.dinb(n3964), .dina(n3968), .dout(n3972));
    jnot g1018(.din(n3972), .dout(n3975));
    jand g1019(.dinb(n10205), .dina(n2259), .dout(n3979));
    jnot g1020(.din(n3979), .dout(n3982));
    jand g1021(.dinb(n3186), .dina(n3982), .dout(n3986));
    jand g1022(.dinb(n3975), .dina(n3986), .dout(n3990));
    jand g1023(.dinb(n7742), .dina(n2228), .dout(n3994));
    jor g1024(.dinb(n2966), .dina(n3994), .dout(n3998));
    jand g1025(.dinb(n11615), .dina(n2271), .dout(n4002));
    jand g1026(.dinb(n10412), .dina(n2220), .dout(n4006));
    jor g1027(.dinb(n4002), .dina(n4006), .dout(n4010));
    jor g1028(.dinb(n3998), .dina(n7107), .dout(n4014));
    jnot g1029(.din(n4014), .dout(n4017));
    jand g1030(.dinb(n7104), .dina(n4017), .dout(n4021));
    jand g1031(.dinb(n7709), .dina(n4021), .dout(n4025));
    jnot g1032(.din(n4025), .dout(n4028));
    jand g1033(.dinb(n7101), .dina(n4028), .dout(n4032));
    jand g1034(.dinb(n12164), .dina(n4032), .dout(n4036));
    jor g1035(.dinb(n7095), .dina(n4036), .dout(n4040));
    jand g1036(.dinb(n8702), .dina(n2621), .dout(n4044));
    jnot g1037(.din(n4044), .dout(n4047));
    jand g1038(.dinb(n4040), .dina(n7071), .dout(n4051));
    jand g1039(.dinb(n3888), .dina(n4051), .dout(n4055));
    jand g1040(.dinb(n7376), .dina(n4055), .dout(n4059));
    jnot g1041(.din(n4059), .dout(n4062));
    jand g1042(.dinb(n3881), .dina(n7050), .dout(n4066));
    jnot g1043(.din(n4066), .dout(n4069));
    jand g1044(.dinb(n10676), .dina(n2733), .dout(n4073));
    jnot g1045(.din(n4073), .dout(n4076));
    jand g1046(.dinb(n11504), .dina(n2251), .dout(n4080));
    jand g1047(.dinb(n11429), .dina(n2201), .dout(n4084));
    jand g1048(.dinb(n11606), .dina(n2279), .dout(n4088));
    jor g1049(.dinb(n4084), .dina(n4088), .dout(n4092));
    jand g1050(.dinb(n11183), .dina(n2228), .dout(n4096));
    jor g1051(.dinb(n4092), .dina(n4096), .dout(n4100));
    jor g1052(.dinb(n7740), .dina(n4100), .dout(n4104));
    jor g1053(.dinb(n8423), .dina(n3176), .dout(n4108));
    jand g1054(.dinb(n10088), .dina(n2271), .dout(n4112));
    jand g1055(.dinb(n9674), .dina(n2220), .dout(n4116));
    jor g1056(.dinb(n4112), .dina(n4116), .dout(n4120));
    jor g1057(.dinb(n11456), .dina(n4120), .dout(n4124));
    jor g1058(.dinb(n4108), .dina(n4124), .dout(n4128));
    jor g1059(.dinb(n4104), .dina(n4128), .dout(n4132));
    jand g1060(.dinb(n8472), .dina(n2251), .dout(n4136));
    jand g1061(.dinb(n10244), .dina(n2201), .dout(n4140));
    jand g1062(.dinb(n8849), .dina(n2220), .dout(n4144));
    jor g1063(.dinb(n4140), .dina(n4144), .dout(n4148));
    jand g1064(.dinb(n8010), .dina(n2271), .dout(n4152));
    jand g1065(.dinb(n10157), .dina(n2186), .dout(n4156));
    jor g1066(.dinb(n7727), .dina(n4156), .dout(n4160));
    jor g1067(.dinb(n7725), .dina(n4160), .dout(n4164));
    jand g1068(.dinb(n8457), .dina(n2279), .dout(n4168));
    jand g1069(.dinb(n7694), .dina(n2228), .dout(n4172));
    jor g1070(.dinb(n7692), .dina(n4172), .dout(n4176));
    jor g1071(.dinb(n7706), .dina(n4176), .dout(n4180));
    jor g1072(.dinb(n4164), .dina(n4180), .dout(n4184));
    jor g1073(.dinb(n7689), .dina(n4184), .dout(n4188));
    jor g1074(.dinb(n7680), .dina(n4188), .dout(n4192));
    jand g1075(.dinb(n7665), .dina(n4192), .dout(n4196));
    jor g1076(.dinb(n9911), .dina(n4196), .dout(n4200));
    jand g1077(.dinb(n9746), .dina(n2621), .dout(n4204));
    jnot g1078(.din(n4204), .dout(n4207));
    jand g1079(.dinb(n4200), .dina(n7659), .dout(n4211));
    jand g1080(.dinb(n4076), .dina(n7644), .dout(n4215));
    jand g1081(.dinb(n11714), .dina(n4215), .dout(n4219));
    jnot g1082(.din(n4219), .dout(n4222));
    jor g1083(.dinb(n7595), .dina(n3784), .dout(n4226));
    jnot g1084(.din(n3738), .dout(n4229));
    jor g1085(.dinb(n7446), .dina(n3780), .dout(n4233));
    jand g1086(.dinb(n4226), .dina(n7443), .dout(n4237));
    jand g1087(.dinb(n7440), .dina(n4237), .dout(n4241));
    jnot g1088(.din(n4241), .dout(n4244));
    jand g1089(.dinb(n3830), .dina(n4066), .dout(n4248));
    jand g1090(.dinb(n7841), .dina(n4241), .dout(n4252));
    jand g1091(.dinb(n3118), .dina(n3574), .dout(n4256));
    jnot g1092(.din(n2464), .dout(n4259));
    jand g1093(.dinb(n9588), .dina(n3379), .dout(n4263));
    jand g1094(.dinb(n4256), .dina(n6714), .dout(n4267));
    jand g1095(.dinb(n4252), .dina(n6711), .dout(n4271));
    jand g1096(.dinb(n6716), .dina(n4271), .dout(n4275));
    jnot g1097(.din(n4275), .dout(n4278));
    jnot g1098(.din(G343), .dout(n4281));
    jand g1099(.dinb(n6953), .dina(n4248), .dout(n4285));
    jnot g1100(.din(G213), .dout(n4288));
    jor g1101(.dinb(n6708), .dina(n4275), .dout(n4292));
    jor g1102(.dinb(n6624), .dina(n4292), .dout(G409));
    jxor g1103(.dinb(n9588), .dina(n3379), .dout(n4300));
    jxor g1104(.dinb(n3118), .dina(n3574), .dout(n4304));
    jxor g1105(.dinb(n8169), .dina(n4304), .dout(n4308));
    jand g1106(.dinb(n10874), .dina(n4281), .dout(n4312));
    jxor g1107(.dinb(n7832), .dina(n4241), .dout(n4316));
    jxor g1108(.dinb(n6873), .dina(n4316), .dout(n4320));
    jand g1109(.dinb(n6875), .dina(n4320), .dout(n4324));
    jnot g1110(.din(n4312), .dout(n4327));
    jxor g1111(.dinb(n3830), .dina(n4066), .dout(n4331));
    jxor g1112(.dinb(n4316), .dina(n4331), .dout(n4335));
    jand g1113(.dinb(n6792), .dina(n4335), .dout(n4339));
    jor g1114(.dinb(n4324), .dina(n4339), .dout(n4343));
    jxor g1115(.dinb(n8156), .dina(n4343), .dout(G405));
    jxor g1116(.dinb(n8166), .dina(n4335), .dout(n4351));
    jdff dff_A_c0IRpd548_0(.din(n12923), .dout(G402));
    jdff dff_A_nMRnQXEZ3_2(.din(n4351), .dout(n12923));
    jdff dff_A_U9Dhhxdh2_1(.din(n4278), .dout(G407));
    jdff dff_A_Pr5W43mi1_0(.din(n12914), .dout(G381));
    jdff dff_A_ntiPQ6aK5_0(.din(n12911), .dout(n12914));
    jdff dff_A_GLrwuIti6_0(.din(n12908), .dout(n12911));
    jdff dff_A_ZFDj4KzA8_1(.din(n4244), .dout(n12908));
    jdff dff_A_OFjJ8rbw8_0(.din(n12902), .dout(G375));
    jdff dff_A_ZtU3tyDA1_0(.din(n12899), .dout(n12902));
    jdff dff_A_0f7I85Sz6_0(.din(n12896), .dout(n12899));
    jdff dff_A_1rpzyvbw3_1(.din(n4069), .dout(n12896));
    jdff dff_A_Tyi4ypDL0_0(.din(n12890), .dout(G378));
    jdff dff_A_zrE6ZEQR2_0(.din(n12887), .dout(n12890));
    jdff dff_A_eOvyUM789_0(.din(n12884), .dout(n12887));
    jdff dff_A_lKt9RnS31_1(.din(n3833), .dout(n12884));
    jdff dff_A_C38MetWn2_0(.din(n12878), .dout(G390));
    jdff dff_A_DlL4fp6E6_0(.din(n12875), .dout(n12878));
    jdff dff_A_wsfjiJc34_0(.din(n12872), .dout(n12875));
    jdff dff_A_K8cjy4tB5_0(.din(n12869), .dout(n12872));
    jdff dff_A_70oyHGSA9_0(.din(n12866), .dout(n12869));
    jdff dff_A_4z7A7QZb0_1(.din(n3577), .dout(n12866));
    jdff dff_A_Jq6zQMHU6_0(.din(n12860), .dout(G393));
    jdff dff_A_21LJ38qi8_0(.din(n12857), .dout(n12860));
    jdff dff_A_P1VdzwAK9_0(.din(n12854), .dout(n12857));
    jdff dff_A_cdgl24GK6_0(.din(n12851), .dout(n12854));
    jdff dff_A_bEHImB6t9_0(.din(n12848), .dout(n12851));
    jdff dff_A_P9xmPpsY4_0(.din(n12845), .dout(n12848));
    jdff dff_A_AxGVX6TL1_1(.din(n3382), .dout(n12845));
    jdff dff_A_ebIqPRx40_0(.din(n12839), .dout(G387));
    jdff dff_A_2VS1HYFM1_0(.din(n12836), .dout(n12839));
    jdff dff_A_BPJNqi4P9_0(.din(n12833), .dout(n12836));
    jdff dff_A_XsprfBTq5_0(.din(n12830), .dout(n12833));
    jdff dff_A_Bt9wVzTt8_0(.din(n12827), .dout(n12830));
    jdff dff_A_9T1uPaDL7_1(.din(n3121), .dout(n12827));
    jdff dff_A_L68NbBTi7_0(.din(n12821), .dout(G367));
    jdff dff_A_hKoYBXx60_0(.din(n12818), .dout(n12821));
    jdff dff_A_Egy2GMK16_0(.din(n12815), .dout(n12818));
    jdff dff_A_KKwkaz148_0(.din(n12812), .dout(n12815));
    jdff dff_A_Za09WhNt1_0(.din(n12809), .dout(n12812));
    jdff dff_A_xIPw46ed7_0(.din(n12806), .dout(n12809));
    jdff dff_A_s1BWpEPJ7_2(.din(n2832), .dout(n12806));
    jdff dff_A_iP8xR4Dp5_0(.din(n12800), .dout(G384));
    jdff dff_A_Qw83aOJF4_0(.din(n12797), .dout(n12800));
    jdff dff_A_zwwGGmF66_0(.din(n12794), .dout(n12797));
    jdff dff_A_kxVVvueZ2_0(.din(n12791), .dout(n12794));
    jdff dff_A_Hs7YH4XS1_0(.din(n12788), .dout(n12791));
    jdff dff_A_OsULOYGU0_0(.din(n12785), .dout(n12788));
    jdff dff_A_s3gw2Kpf0_0(.din(n12782), .dout(n12785));
    jdff dff_A_w0ospIK34_1(.din(n2693), .dout(n12782));
    jdff dff_A_pYpDbVvt6_0(.din(n12776), .dout(G396));
    jdff dff_A_TJTCX4ic6_0(.din(n12773), .dout(n12776));
    jdff dff_A_RWQgGR7b9_0(.din(n12770), .dout(n12773));
    jdff dff_A_B1rZOdhm8_0(.din(n12767), .dout(n12770));
    jdff dff_A_C3fHhtX00_0(.din(n12764), .dout(n12767));
    jdff dff_A_xToQ7eE15_0(.din(n12761), .dout(n12764));
    jdff dff_A_2mzac4AP3_0(.din(n12758), .dout(n12761));
    jdff dff_A_fjYciVHo3_0(.din(n12755), .dout(n12758));
    jdff dff_A_zaFEr2Qo4_0(.din(n12752), .dout(n12755));
    jdff dff_A_1XaNwXtd4_0(.din(n12749), .dout(n12752));
    jdff dff_A_gpCErC2J7_0(.din(n12746), .dout(n12749));
    jdff dff_A_OFpUOMpJ2_0(.din(n12743), .dout(n12746));
    jdff dff_A_0XfjDTOX8_1(.din(n2464), .dout(n12743));
    jdff dff_A_qFi8lNVn2_0(.din(n12737), .dout(G364));
    jdff dff_A_aDbrixL86_0(.din(n12734), .dout(n12737));
    jdff dff_A_izzAIYDC1_0(.din(n12731), .dout(n12734));
    jdff dff_A_s9buAJxf5_0(.din(n12728), .dout(n12731));
    jdff dff_A_KRnIQjkJ0_0(.din(n12725), .dout(n12728));
    jdff dff_A_GDYQeMP93_0(.din(n12722), .dout(n12725));
    jdff dff_A_GkwRoEH73_0(.din(n12719), .dout(n12722));
    jdff dff_A_Mib1ZxWW6_0(.din(n12716), .dout(n12719));
    jdff dff_A_PHITdRC31_2(.din(n2112), .dout(n12716));
    jdff dff_A_Q2ojPoe65_0(.din(n12710), .dout(G399));
    jdff dff_A_cDq0uFlu5_0(.din(n12707), .dout(n12710));
    jdff dff_A_e250Ta4u5_0(.din(n12704), .dout(n12707));
    jdff dff_A_s7KFIQBH1_0(.din(n12701), .dout(n12704));
    jdff dff_A_EdHWmoz13_0(.din(n12698), .dout(n12701));
    jdff dff_A_hok2NpAF2_0(.din(n12695), .dout(n12698));
    jdff dff_A_6yVs5rtw8_0(.din(n12692), .dout(n12695));
    jdff dff_A_m3L8a7Bg5_0(.din(n12689), .dout(n12692));
    jdff dff_A_ZVNovf346_0(.din(n12686), .dout(n12689));
    jdff dff_A_lgoO7Orz8_0(.din(n12683), .dout(n12686));
    jdff dff_A_ZLF4pp3d5_0(.din(n12680), .dout(n12683));
    jdff dff_A_BN5PaiSn9_0(.din(n12677), .dout(n12680));
    jdff dff_A_KjTc5jEp4_0(.din(n12674), .dout(n12677));
    jdff dff_A_UHzT0RaE1_2(.din(n2005), .dout(n12674));
    jdff dff_A_4m1UV7fw5_0(.din(n12668), .dout(G369));
    jdff dff_A_o8MDBcjX5_0(.din(n12665), .dout(n12668));
    jdff dff_A_FFSEMvOO7_0(.din(n12662), .dout(n12665));
    jdff dff_A_a4QoQGjb7_0(.din(n12659), .dout(n12662));
    jdff dff_A_oEKfbMSB8_0(.din(n12656), .dout(n12659));
    jdff dff_A_5GmK2co63_0(.din(n12653), .dout(n12656));
    jdff dff_A_85QK85lL7_0(.din(n12650), .dout(n12653));
    jdff dff_A_fknHQfj16_0(.din(n12647), .dout(n12650));
    jdff dff_A_7Zfn1xMY5_0(.din(n12644), .dout(n12647));
    jdff dff_A_c0es5wGK8_0(.din(n12641), .dout(n12644));
    jdff dff_A_OyvXMKs59_0(.din(n12638), .dout(n12641));
    jdff dff_A_qRdAfI1F8_2(.din(n1940), .dout(n12638));
    jdff dff_A_S4Ge7OwR4_0(.din(n12632), .dout(G372));
    jdff dff_A_iCJ2GGev6_0(.din(n12629), .dout(n12632));
    jdff dff_A_C4EbJt2q8_0(.din(n12626), .dout(n12629));
    jdff dff_A_4gVZ4j902_0(.din(n12623), .dout(n12626));
    jdff dff_A_urGzhT8P2_0(.din(n12620), .dout(n12623));
    jdff dff_A_XzLmBfRQ1_0(.din(n12617), .dout(n12620));
    jdff dff_A_VmKEePlN2_0(.din(n12614), .dout(n12617));
    jdff dff_A_lFczkg4K6_0(.din(n12611), .dout(n12614));
    jdff dff_A_85CUouSP3_0(.din(n12608), .dout(n12611));
    jdff dff_A_d6sMEsnZ6_0(.din(n12605), .dout(n12608));
    jdff dff_A_FAjOD6Oi6_0(.din(n12602), .dout(n12605));
    jdff dff_A_gjrpNmAA2_0(.din(n12599), .dout(n12602));
    jdff dff_A_EoICxVBu2_0(.din(n12596), .dout(n12599));
    jdff dff_A_JAByGg7B5_2(.din(n1759), .dout(n12596));
    jdff dff_A_HJpBciPx2_0(.din(n12590), .dout(G351));
    jdff dff_A_HbUE7IYu9_0(.din(n12587), .dout(n12590));
    jdff dff_A_cmSYvPGX9_0(.din(n12584), .dout(n12587));
    jdff dff_A_meWnGMiq9_0(.din(n12581), .dout(n12584));
    jdff dff_A_Cq8yWShR4_0(.din(n12578), .dout(n12581));
    jdff dff_A_qP85N9KR9_0(.din(n12575), .dout(n12578));
    jdff dff_A_9FAkzqTC5_0(.din(n12572), .dout(n12575));
    jdff dff_A_946hA4991_0(.din(n12569), .dout(n12572));
    jdff dff_A_MoOazLC59_0(.din(n12566), .dout(n12569));
    jdff dff_A_HdJhXA425_0(.din(n12563), .dout(n12566));
    jdff dff_A_QmxGzTpy0_0(.din(n12560), .dout(n12563));
    jdff dff_A_AJaRT1qj2_0(.din(n12557), .dout(n12560));
    jdff dff_A_j1ky04Bg4_0(.din(n12554), .dout(n12557));
    jdff dff_A_Ojk52XmW4_0(.din(n12551), .dout(n12554));
    jdff dff_A_YmqN1DgV8_0(.din(n12548), .dout(n12551));
    jdff dff_A_1csAG2rb0_0(.din(n12545), .dout(n12548));
    jdff dff_A_ueyEnQai1_0(.din(n12542), .dout(n12545));
    jdff dff_A_xGH5Ivs95_0(.din(n12539), .dout(n12542));
    jdff dff_A_kMvDyWg85_0(.din(n12536), .dout(n12539));
    jdff dff_A_O5cozlGr7_0(.din(n12533), .dout(n12536));
    jdff dff_A_8mzykBEF3_0(.din(n12530), .dout(n12533));
    jdff dff_A_qjN0MhyM1_0(.din(n12527), .dout(n12530));
    jdff dff_A_k5TFpQE33_0(.din(n12524), .dout(n12527));
    jdff dff_A_tJd3NBRk9_0(.din(n12521), .dout(n12524));
    jdff dff_A_sMhKaenh0_0(.din(n12518), .dout(n12521));
    jdff dff_A_2lCTvU9h2_0(.din(n12515), .dout(n12518));
    jdff dff_A_jxO7Gb1E1_2(.din(n318), .dout(n12515));
    jdff dff_A_q1pa0OsA6_0(.din(n12509), .dout(G358));
    jdff dff_A_qiXxe7Fc9_0(.din(n12506), .dout(n12509));
    jdff dff_A_QrDGQSQd8_0(.din(n12503), .dout(n12506));
    jdff dff_A_qRv3Kthb3_0(.din(n12500), .dout(n12503));
    jdff dff_A_K9ynOQIK4_0(.din(n12497), .dout(n12500));
    jdff dff_A_Y3Md220M2_0(.din(n12494), .dout(n12497));
    jdff dff_A_mvxanOFS4_0(.din(n12491), .dout(n12494));
    jdff dff_A_RToiNRdE6_0(.din(n12488), .dout(n12491));
    jdff dff_A_UFIMXzq03_0(.din(n12485), .dout(n12488));
    jdff dff_A_8RHrabNL8_0(.din(n12482), .dout(n12485));
    jdff dff_A_VyaPxz1f2_0(.din(n12479), .dout(n12482));
    jdff dff_A_uzyAGsou2_0(.din(n12476), .dout(n12479));
    jdff dff_A_AGd7AVLH3_0(.din(n12473), .dout(n12476));
    jdff dff_A_fhGLWfSZ6_0(.din(n12470), .dout(n12473));
    jdff dff_A_vqd355fq0_0(.din(n12467), .dout(n12470));
    jdff dff_A_UAe7Fu759_0(.din(n12464), .dout(n12467));
    jdff dff_A_Nihax5y29_0(.din(n12461), .dout(n12464));
    jdff dff_A_qUW0RoQM1_0(.din(n12458), .dout(n12461));
    jdff dff_A_dHku9i8q2_0(.din(n12455), .dout(n12458));
    jdff dff_A_6xS7V23c1_0(.din(n12452), .dout(n12455));
    jdff dff_A_mRQio0LQ0_0(.din(n12449), .dout(n12452));
    jdff dff_A_cK1OG4ZC5_0(.din(n12446), .dout(n12449));
    jdff dff_A_viKuLYhm9_0(.din(n12443), .dout(n12446));
    jdff dff_A_SxW2B5cl0_0(.din(n12440), .dout(n12443));
    jdff dff_A_CFNiCZF28_0(.din(n12437), .dout(n12440));
    jdff dff_A_LguSs9EC9_2(.din(n290), .dout(n12437));
    jdff dff_A_1F2vq7cY6_0(.din(n12431), .dout(G361));
    jdff dff_A_S8FkLZxb3_0(.din(n12428), .dout(n12431));
    jdff dff_A_MiEXD3jG9_0(.din(n12425), .dout(n12428));
    jdff dff_A_ADLAh3eJ8_0(.din(n12422), .dout(n12425));
    jdff dff_A_SJifkAxx4_0(.din(n12419), .dout(n12422));
    jdff dff_A_eylU7JFY2_0(.din(n12416), .dout(n12419));
    jdff dff_A_MLO4bTuK9_0(.din(n12413), .dout(n12416));
    jdff dff_A_5iZI7iGb1_0(.din(n12410), .dout(n12413));
    jdff dff_A_mVa35RVi0_0(.din(n12407), .dout(n12410));
    jdff dff_A_TWoDI0xq5_0(.din(n12404), .dout(n12407));
    jdff dff_A_wNyduM9r0_0(.din(n12401), .dout(n12404));
    jdff dff_A_5KRr7hOJ1_0(.din(n12398), .dout(n12401));
    jdff dff_A_fXDVISIz7_0(.din(n12395), .dout(n12398));
    jdff dff_A_WMmrDgGo0_0(.din(n12392), .dout(n12395));
    jdff dff_A_xeiXKon84_0(.din(n12389), .dout(n12392));
    jdff dff_A_zWpc0EmV8_0(.din(n12386), .dout(n12389));
    jdff dff_A_8qzrIc9S6_0(.din(n12383), .dout(n12386));
    jdff dff_A_OKX3pUMK6_0(.din(n12380), .dout(n12383));
    jdff dff_A_k3cg0RrP9_0(.din(n12377), .dout(n12380));
    jdff dff_A_2tAQ40B94_0(.din(n12374), .dout(n12377));
    jdff dff_A_eOMG95CX1_0(.din(n12371), .dout(n12374));
    jdff dff_A_2JWF9wm07_0(.din(n12368), .dout(n12371));
    jdff dff_A_dcDQDPxH8_2(.din(n259), .dout(n12368));
    jdff dff_A_MhNMV9bW1_0(.din(n12362), .dout(G355));
    jdff dff_A_09oKH6DA8_0(.din(n12359), .dout(n12362));
    jdff dff_A_mE5NcZom7_0(.din(n12356), .dout(n12359));
    jdff dff_A_8mTF0rtj6_0(.din(n12353), .dout(n12356));
    jdff dff_A_WhhtPLAe0_0(.din(n12350), .dout(n12353));
    jdff dff_A_p1L3MV9H0_0(.din(n12347), .dout(n12350));
    jdff dff_A_rmUqLk1b0_0(.din(n12344), .dout(n12347));
    jdff dff_A_7zuE67D02_0(.din(n12341), .dout(n12344));
    jdff dff_A_mknWWI8a5_0(.din(n12338), .dout(n12341));
    jdff dff_A_N0on1wpE3_0(.din(n12335), .dout(n12338));
    jdff dff_A_1GVJ6AsH9_0(.din(n12332), .dout(n12335));
    jdff dff_A_O3bEJz710_0(.din(n12329), .dout(n12332));
    jdff dff_A_VQDCUjM34_0(.din(n12326), .dout(n12329));
    jdff dff_A_CqozIHur5_0(.din(n12323), .dout(n12326));
    jdff dff_A_ZTSJahtc0_0(.din(n12320), .dout(n12323));
    jdff dff_A_T1Ru8qFm5_0(.din(n12317), .dout(n12320));
    jdff dff_A_nRxvoZy43_0(.din(n12314), .dout(n12317));
    jdff dff_A_fxx806kt2_0(.din(n12311), .dout(n12314));
    jdff dff_A_C5vjGe879_0(.din(n12308), .dout(n12311));
    jdff dff_A_1bFkcBog0_0(.din(n12305), .dout(n12308));
    jdff dff_A_P98P93Vo1_0(.din(n12302), .dout(n12305));
    jdff dff_A_BM61Geu76_0(.din(n12299), .dout(n12302));
    jdff dff_A_4Z0zJ60r3_0(.din(n12296), .dout(n12299));
    jdff dff_A_3ouQPzKh8_0(.din(n12293), .dout(n12296));
    jdff dff_A_zSHMdOlg5_0(.din(n12290), .dout(n12293));
    jdff dff_A_oBlulQxO4_0(.din(n12287), .dout(n12290));
    jdff dff_A_6FpreaDL9_0(.din(n12284), .dout(n12287));
    jdff dff_A_heHbqSsj6_1(.din(n112), .dout(n12284));
    jdff dff_A_kWSj6xz52_0(.din(n12278), .dout(G353));
    jdff dff_A_E6yqJQNg3_0(.din(n12275), .dout(n12278));
    jdff dff_A_3NHEjUHK0_0(.din(n12272), .dout(n12275));
    jdff dff_A_xiulzJwB2_0(.din(n12269), .dout(n12272));
    jdff dff_A_IRyFOeZM1_0(.din(n12266), .dout(n12269));
    jdff dff_A_jOVPISwb2_0(.din(n12263), .dout(n12266));
    jdff dff_A_QyRcSd7n2_0(.din(n12260), .dout(n12263));
    jdff dff_A_Q01RmBgn9_0(.din(n12257), .dout(n12260));
    jdff dff_A_eOJ13Mva0_0(.din(n12254), .dout(n12257));
    jdff dff_A_USFsF0Q75_0(.din(n12251), .dout(n12254));
    jdff dff_A_bC1ONhvq0_0(.din(n12248), .dout(n12251));
    jdff dff_A_jn2ogL1S9_0(.din(n12245), .dout(n12248));
    jdff dff_A_MFrcOJQK7_0(.din(n12242), .dout(n12245));
    jdff dff_A_Vpq56JlK0_0(.din(n12239), .dout(n12242));
    jdff dff_A_ugjitDbz9_0(.din(n12236), .dout(n12239));
    jdff dff_A_ICHD9OEJ4_0(.din(n12233), .dout(n12236));
    jdff dff_A_il6Dvlg90_0(.din(n12230), .dout(n12233));
    jdff dff_A_EuImGtAL1_0(.din(n12227), .dout(n12230));
    jdff dff_A_bzLOMo5p2_0(.din(n12224), .dout(n12227));
    jdff dff_A_AVbjljYj0_0(.din(n12221), .dout(n12224));
    jdff dff_A_tz7QtjWd6_0(.din(n12218), .dout(n12221));
    jdff dff_A_SOvO5oUh8_0(.din(n12215), .dout(n12218));
    jdff dff_A_c8gsiFJd5_0(.din(n12212), .dout(n12215));
    jdff dff_A_S5KM9Trm0_0(.din(n12209), .dout(n12212));
    jdff dff_A_6BjZhAeX9_0(.din(n12206), .dout(n12209));
    jdff dff_A_8wK8UJoV2_0(.din(n12203), .dout(n12206));
    jdff dff_A_Ai93AJFG8_2(.din(n95), .dout(n12203));
    jdff dff_A_jIXxqQBl5_2(.din(n412), .dout(n12200));
    jdff dff_A_nTFcBRwC5_2(.din(n12200), .dout(n12197));
    jdff dff_A_Ug09h26b1_1(.din(n412), .dout(n12194));
    jdff dff_A_RBGcIbgw2_1(.din(n12194), .dout(n12191));
    jdff dff_A_cY9hvLqp3_1(.din(n12191), .dout(n12188));
    jdff dff_A_DGZgzgEp6_1(.din(n12188), .dout(n12185));
    jdff dff_A_T1y13SqN0_1(.din(n12185), .dout(n12182));
    jdff dff_A_4vkk07dQ3_1(.din(n12182), .dout(n12179));
    jdff dff_A_jkhOXIw50_1(.din(n12179), .dout(n12176));
    jdff dff_A_xir4isHr5_1(.din(n12176), .dout(n12173));
    jdff dff_A_skFdznOb0_1(.din(n12173), .dout(n12170));
    jdff dff_A_qD6GtDDf0_1(.din(n12170), .dout(n12167));
    jdff dff_A_kTSf2yCF4_1(.din(n12167), .dout(n12164));
    jdff dff_A_4X5ktXLG6_2(.din(G20), .dout(n12161));
    jdff dff_A_umfdCvHV8_0(.din(G20), .dout(n12158));
    jdff dff_A_WDaLdjET0_2(.din(G20), .dout(n12155));
    jdff dff_A_K1JJceJN9_2(.din(n12155), .dout(n12152));
    jdff dff_A_4naE8Tex9_0(.din(G20), .dout(n12149));
    jdff dff_A_8ZETPY5M4_0(.din(n12149), .dout(n12146));
    jdff dff_A_Z3J2hJSb1_2(.din(G1), .dout(n12143));
    jdff dff_A_rq0kkRTd8_2(.din(n12143), .dout(n12140));
    jdff dff_A_5tQGUpOt2_2(.din(n12140), .dout(n12137));
    jdff dff_A_NOPU9yVk7_2(.din(n12137), .dout(n12134));
    jdff dff_A_aAR6pYCz9_1(.din(G1), .dout(n12131));
    jdff dff_A_e3s8cSwM6_0(.din(G13), .dout(n12128));
    jdff dff_A_guTVlD6N5_2(.din(n2092), .dout(n12125));
    jdff dff_A_wDowTD480_2(.din(n12125), .dout(n12122));
    jdff dff_A_4RapG7jq9_2(.din(n12122), .dout(n12119));
    jdff dff_A_XeLfyT332_2(.din(n12119), .dout(n12116));
    jdff dff_A_ezUndS1G2_2(.din(n12116), .dout(n12113));
    jdff dff_A_dyi1Gi8L2_2(.din(n12113), .dout(n12110));
    jdff dff_A_dUxOj9k29_2(.din(n12110), .dout(n12107));
    jdff dff_A_obwNyN3M3_2(.din(n12107), .dout(n12104));
    jdff dff_A_G9GbJgRh8_2(.din(n12104), .dout(n12101));
    jdff dff_A_isP7eMnG7_2(.din(n12101), .dout(n12098));
    jdff dff_A_N1HLg4Qb8_2(.din(n12098), .dout(n12095));
    jdff dff_A_hTCvXI2g6_2(.din(n12095), .dout(n12092));
    jdff dff_A_j50Xlt662_2(.din(n12092), .dout(n12089));
    jdff dff_A_NQJiFtDC4_2(.din(n12089), .dout(n12086));
    jdff dff_A_2noCDfoW2_2(.din(n12086), .dout(n12083));
    jdff dff_A_3cnhfRbG6_2(.din(n12083), .dout(n12080));
    jdff dff_A_0NHp2NW70_0(.din(n2092), .dout(n12077));
    jdff dff_A_PUd3i7Rp2_0(.din(n12077), .dout(n12074));
    jdff dff_A_61jEzgoa0_0(.din(n12074), .dout(n12071));
    jdff dff_A_1aQXot4l1_0(.din(n12071), .dout(n12068));
    jdff dff_A_WDZpszBJ8_0(.din(n12068), .dout(n12065));
    jdff dff_A_96EuYVYl3_0(.din(n12065), .dout(n12062));
    jdff dff_A_Tszw1cSD1_0(.din(n12062), .dout(n12059));
    jdff dff_A_taupPDeH9_0(.din(n12059), .dout(n12056));
    jdff dff_A_Abwx3fK25_0(.din(n12056), .dout(n12053));
    jdff dff_A_RHuUdByJ7_0(.din(n12053), .dout(n12050));
    jdff dff_A_wQHYfsYp4_0(.din(n12050), .dout(n12047));
    jdff dff_A_p3nTqZD10_0(.din(n12047), .dout(n12044));
    jdff dff_A_wmUZLzCh4_0(.din(n12044), .dout(n12041));
    jdff dff_A_2J4xUV9f5_0(.din(n12041), .dout(n12038));
    jdff dff_A_InXusHiD4_0(.din(n2092), .dout(n12035));
    jdff dff_A_HDp4Rv4b7_0(.din(n12035), .dout(n12032));
    jdff dff_A_79mn2xNf3_0(.din(n12032), .dout(n12029));
    jdff dff_A_1qPTpA1q6_0(.din(n12029), .dout(n12026));
    jdff dff_A_AX1G0bb44_0(.din(n12026), .dout(n12023));
    jdff dff_A_wEp1EegM7_0(.din(n12023), .dout(n12020));
    jdff dff_A_YTEdMcQC8_0(.din(n12020), .dout(n12017));
    jdff dff_A_ywYiSN8k3_0(.din(n12017), .dout(n12014));
    jdff dff_A_cWYLC7ju0_0(.din(n12014), .dout(n12011));
    jdff dff_A_iVRRV7Sw1_0(.din(n12011), .dout(n12008));
    jdff dff_A_F7ERN3hQ1_0(.din(n12008), .dout(n12005));
    jdff dff_A_aI1RUtP61_0(.din(n12005), .dout(n12002));
    jdff dff_A_H35nGzRP5_0(.din(n12002), .dout(n11999));
    jdff dff_A_qSKEbZh49_0(.din(n11999), .dout(n11996));
    jdff dff_A_N5jP9i6U3_0(.din(G1), .dout(n11993));
    jdff dff_A_yAMMVBFC6_0(.din(n11993), .dout(n11990));
    jdff dff_A_VsLbwrtO3_2(.din(n333), .dout(n11987));
    jdff dff_A_S8Ex2UsS9_0(.din(G20), .dout(n11984));
    jdff dff_A_0bioxm1z1_2(.din(n367), .dout(n11981));
    jdff dff_A_XHe6xMWF4_2(.din(n11981), .dout(n11978));
    jdff dff_A_6jCIhLww4_0(.din(n367), .dout(n11975));
    jdff dff_A_aZAttY8G0_1(.din(G45), .dout(n11972));
    jdff dff_A_JMvy7szU2_1(.din(n11972), .dout(n11969));
    jdff dff_A_egaZa6cr5_1(.din(n11969), .dout(n11966));
    jdff dff_B_ZKL3QDgj6_3(.din(n2127), .dout(n11964));
    jdff dff_A_qEGBsBzK4_2(.din(n11964), .dout(n11960));
    jdff dff_A_Rj63iQgT8_2(.din(n11960), .dout(n11957));
    jdff dff_A_JXIXWcGo8_2(.din(n11957), .dout(n11954));
    jdff dff_A_4G8okOjd0_2(.din(n11954), .dout(n11951));
    jdff dff_A_AJeI4UoQ8_2(.din(n11951), .dout(n11948));
    jdff dff_A_VrYoCOTw7_2(.din(n11948), .dout(n11945));
    jdff dff_A_M8HdTe4Q8_2(.din(n11945), .dout(n11942));
    jdff dff_A_IHTSHDyC1_2(.din(n11942), .dout(n11939));
    jdff dff_A_GsdaWvN54_2(.din(n11939), .dout(n11936));
    jdff dff_A_4DpscUuV9_2(.din(n11936), .dout(n11933));
    jdff dff_A_0CweugFC8_2(.din(n11933), .dout(n11930));
    jdff dff_A_fOGu7ZWA5_2(.din(n11930), .dout(n11927));
    jdff dff_A_496hTPo42_2(.din(n11927), .dout(n11924));
    jdff dff_A_0wVrAMwP3_2(.din(n11924), .dout(n11921));
    jdff dff_A_d4rvyG4T9_2(.din(n11921), .dout(n11918));
    jdff dff_A_wA86aAFS4_2(.din(n11918), .dout(n11915));
    jdff dff_A_kFe3LRGZ8_2(.din(n11915), .dout(n11912));
    jdff dff_A_e63nU98t4_1(.din(n11964), .dout(n11909));
    jdff dff_A_KoqiKnEX4_1(.din(n11909), .dout(n11906));
    jdff dff_A_2x6djRsS9_1(.din(n11906), .dout(n11903));
    jdff dff_A_5C1hva4C5_1(.din(n11903), .dout(n11900));
    jdff dff_A_v9xiFeg96_1(.din(n11900), .dout(n11897));
    jdff dff_A_CtcEoa8n2_1(.din(n11897), .dout(n11894));
    jdff dff_A_x1s2U30T8_1(.din(n11894), .dout(n11891));
    jdff dff_A_nqPUHYk00_1(.din(n11891), .dout(n11888));
    jdff dff_A_vfWf3gR25_1(.din(n11888), .dout(n11885));
    jdff dff_A_DQGtUc2l6_1(.din(n11885), .dout(n11882));
    jdff dff_A_tkGJ9t5y6_1(.din(n11882), .dout(n11879));
    jdff dff_A_V4OFxZ083_1(.din(n11879), .dout(n11876));
    jdff dff_A_WbCy81H91_1(.din(n11876), .dout(n11873));
    jdff dff_A_VIhe6DUA7_1(.din(n11873), .dout(n11870));
    jdff dff_A_wuQD9Hzj0_1(.din(n11870), .dout(n11867));
    jdff dff_A_zKqqXszk4_1(.din(n11964), .dout(n11864));
    jdff dff_A_9VP9IOha1_1(.din(n11864), .dout(n11861));
    jdff dff_A_QF5aFoH61_1(.din(n11861), .dout(n11858));
    jdff dff_A_iVqHq4Hr1_1(.din(n11858), .dout(n11855));
    jdff dff_A_VaePAUu87_1(.din(n11855), .dout(n11852));
    jdff dff_A_GY1MIUoT5_1(.din(n11852), .dout(n11849));
    jdff dff_A_9Coo9IHi9_1(.din(n11849), .dout(n11846));
    jdff dff_A_eUW2J06r9_1(.din(n11846), .dout(n11843));
    jdff dff_A_r1h7pgr00_1(.din(n11843), .dout(n11840));
    jdff dff_A_DlW4a4Wk7_1(.din(n11840), .dout(n11837));
    jdff dff_A_x3oAx41T3_1(.din(n11837), .dout(n11834));
    jdff dff_A_C23dacP67_1(.din(n11834), .dout(n11831));
    jdff dff_A_tFYi5S421_1(.din(n11831), .dout(n11828));
    jdff dff_A_aSvgI4nP6_1(.din(n11828), .dout(n11825));
    jdff dff_A_WPwKHGLe3_0(.din(n11964), .dout(n11822));
    jdff dff_A_5zyMBQ4e6_0(.din(n11822), .dout(n11819));
    jdff dff_A_6cth4LiG5_0(.din(n11819), .dout(n11816));
    jdff dff_A_MyorrT4o6_0(.din(n11816), .dout(n11813));
    jdff dff_A_TpMP28h14_0(.din(n11813), .dout(n11810));
    jdff dff_A_OkecXknK2_0(.din(n11810), .dout(n11807));
    jdff dff_A_n64U0nQk4_0(.din(n11807), .dout(n11804));
    jdff dff_A_NnUSno4B3_0(.din(n11804), .dout(n11801));
    jdff dff_A_8AQttcRs1_0(.din(n11801), .dout(n11798));
    jdff dff_A_s2AiT7Rh9_0(.din(n11798), .dout(n11795));
    jdff dff_A_AelXYhZ19_0(.din(n11795), .dout(n11792));
    jdff dff_A_sfT8hdn89_0(.din(n11792), .dout(n11789));
    jdff dff_A_eOOd4Wzs3_0(.din(n11789), .dout(n11786));
    jdff dff_A_9O5Nxu9W0_0(.din(n11786), .dout(n11783));
    jdff dff_A_pMifdcYw3_2(.din(n2131), .dout(n11780));
    jdff dff_A_fOMhSwhw7_2(.din(n11780), .dout(n11777));
    jdff dff_A_FcQcbM5U6_2(.din(n11777), .dout(n11774));
    jdff dff_A_qshZv7hQ7_2(.din(n11774), .dout(n11771));
    jdff dff_A_fp8UZbm02_2(.din(n11771), .dout(n11768));
    jdff dff_A_TQSST8xv0_1(.din(n2131), .dout(n11765));
    jdff dff_A_8v5wyk799_1(.din(n11765), .dout(n11762));
    jdff dff_A_X7aHFhnq1_1(.din(n11762), .dout(n11759));
    jdff dff_A_dRxpiVZy0_1(.din(n11759), .dout(n11756));
    jdff dff_A_L1rxmO587_1(.din(n11756), .dout(n11753));
    jdff dff_A_1ETxCsuV3_1(.din(n11753), .dout(n11750));
    jdff dff_A_LJbc8UgO7_1(.din(n11750), .dout(n11747));
    jdff dff_A_OF6GhCY34_2(.din(n2131), .dout(n11744));
    jdff dff_A_2eUFjgy66_2(.din(n11744), .dout(n11741));
    jdff dff_A_gidrEGX38_2(.din(n11741), .dout(n11738));
    jdff dff_A_sucSOSwM4_2(.din(n11738), .dout(n11735));
    jdff dff_A_lWijELjg8_2(.din(n11735), .dout(n11732));
    jdff dff_A_NgFE8Z6K9_2(.din(n11732), .dout(n11729));
    jdff dff_A_ZWk61n8A7_2(.din(n11729), .dout(n11726));
    jdff dff_A_fOXKGzIH2_2(.din(n11726), .dout(n11723));
    jdff dff_A_8c6wB8ym4_2(.din(n11723), .dout(n11720));
    jdff dff_A_NtHf2mZN3_2(.din(n11720), .dout(n11717));
    jdff dff_A_riJUsCaV4_2(.din(n11717), .dout(n11714));
    jdff dff_A_ax2aeJKe0_0(.din(n2131), .dout(n11711));
    jdff dff_A_pe4VyM901_0(.din(n11711), .dout(n11708));
    jdff dff_A_uHCxWV2a9_0(.din(n2131), .dout(n11705));
    jdff dff_A_Rnhv3WZw1_0(.din(n11705), .dout(n11702));
    jdff dff_A_nMsuSsbP8_0(.din(n11702), .dout(n11699));
    jdff dff_A_yc5yqWwW4_0(.din(n11699), .dout(n11696));
    jdff dff_A_PednxCB11_0(.din(n11696), .dout(n11693));
    jdff dff_A_tYyIqU8I4_0(.din(n11693), .dout(n11690));
    jdff dff_A_tOSKmY9K7_0(.din(n11690), .dout(n11687));
    jdff dff_A_VPZDvZ3B7_0(.din(n11687), .dout(n11684));
    jdff dff_A_QGN3FYtA1_0(.din(n11684), .dout(n11681));
    jdff dff_A_EIouoLnc5_0(.din(n11681), .dout(n11678));
    jdff dff_B_LllyakdK2_3(.din(n11673), .dout(n11676));
    jdff dff_B_XISZZfl35_3(.din(n11670), .dout(n11673));
    jdff dff_B_D5Bx6L4k1_3(.din(n11667), .dout(n11670));
    jdff dff_B_9VXUoVH00_3(.din(n11664), .dout(n11667));
    jdff dff_B_3lrWq1ZZ2_3(.din(n11661), .dout(n11664));
    jdff dff_B_MahJQJth5_3(.din(n11658), .dout(n11661));
    jdff dff_B_qbxsD1Wv8_3(.din(n11655), .dout(n11658));
    jdff dff_B_5gC5FILO3_3(.din(n11652), .dout(n11655));
    jdff dff_B_90HfVKk17_3(.din(n11649), .dout(n11652));
    jdff dff_B_rHPmGMoo8_3(.din(n11646), .dout(n11649));
    jdff dff_B_6bk3x7n79_3(.din(n11643), .dout(n11646));
    jdff dff_B_ni0jTr7x7_3(.din(n11640), .dout(n11643));
    jdff dff_B_KJmYe58O5_3(.din(G330), .dout(n11640));
    jdff dff_A_2LB4S6lL1_2(.din(n11676), .dout(n11636));
    jdff dff_A_92WyQHFf7_0(.din(n11676), .dout(n11633));
    jdff dff_A_7SiU0GIE8_2(.din(G116), .dout(n11630));
    jdff dff_A_OWUQhYUJ5_2(.din(n11630), .dout(n11627));
    jdff dff_A_v6Tm0TTV7_2(.din(n11627), .dout(n11624));
    jdff dff_A_6Jnib6tG3_1(.din(G116), .dout(n11621));
    jdff dff_A_wYohYmHl8_1(.din(n11621), .dout(n11618));
    jdff dff_A_1mvVggJS4_1(.din(n11618), .dout(n11615));
    jdff dff_A_7FnPaeON8_2(.din(G116), .dout(n11612));
    jdff dff_A_FPq6sE740_2(.din(n11612), .dout(n11609));
    jdff dff_A_AhkhnfD37_2(.din(n11609), .dout(n11606));
    jdff dff_A_VKaiihHm3_1(.din(G116), .dout(n11603));
    jdff dff_A_cIXMQj1C0_0(.din(G116), .dout(n11600));
    jdff dff_A_Y9rTJxB16_0(.din(n11600), .dout(n11597));
    jdff dff_A_ksJxD0uI3_0(.din(n11597), .dout(n11594));
    jdff dff_A_t1IPvC8r1_0(.din(n11594), .dout(n11591));
    jdff dff_A_fBrIb4Yj7_0(.din(n11591), .dout(n11588));
    jdff dff_A_XtbjMlao6_0(.din(n11588), .dout(n11585));
    jdff dff_A_DU8SRIU89_1(.din(G13), .dout(n11582));
    jdff dff_A_a2pL4i4R6_0(.din(G13), .dout(n11579));
    jdff dff_A_TYwDA2GO3_0(.din(n11579), .dout(n11576));
    jdff dff_A_Xf56kWhH1_2(.din(n322), .dout(n11573));
    jdff dff_A_4m3fVzqZ7_0(.din(n322), .dout(n11570));
    jdff dff_A_Fe2KaN991_0(.din(G33), .dout(n11567));
    jdff dff_A_7hmPxE388_0(.din(n11567), .dout(n11564));
    jdff dff_A_JUyi6zAp5_0(.din(n11564), .dout(n11561));
    jdff dff_A_6UMkh2iw9_2(.din(G33), .dout(n11558));
    jdff dff_A_4G19A59n2_1(.din(G33), .dout(n11555));
    jdff dff_A_H7EoIeNt4_0(.din(n330), .dout(n11552));
    jdff dff_A_1QcmdyLC6_0(.din(n11552), .dout(n11549));
    jdff dff_B_TWpw5Lkn9_0(.din(n11544), .dout(n11547));
    jdff dff_B_myevPPDS9_0(.din(n349), .dout(n11544));
    jdff dff_A_aCfmhJLD5_0(.din(G116), .dout(n11540));
    jdff dff_A_rrN7MSkv5_0(.din(n11540), .dout(n11537));
    jdff dff_A_rB8oE75a0_0(.din(n11537), .dout(n11534));
    jdff dff_A_J6xfLXCV2_2(.din(n367), .dout(n11531));
    jdff dff_A_rMTa615l0_2(.din(n11531), .dout(n11528));
    jdff dff_A_QoYS69xf0_1(.din(n367), .dout(n11525));
    jdff dff_A_lypYdccR6_0(.din(n11528), .dout(n11522));
    jdff dff_A_IrXp32UJ4_1(.din(G283), .dout(n11519));
    jdff dff_A_W7JmUWlk9_1(.din(n11519), .dout(n11516));
    jdff dff_A_raukKi4E5_1(.din(n11516), .dout(n11513));
    jdff dff_A_G7tY3cCa7_0(.din(G283), .dout(n11510));
    jdff dff_A_DXX6RVdY6_0(.din(n11510), .dout(n11507));
    jdff dff_A_NqqpT5bS4_0(.din(n11507), .dout(n11504));
    jdff dff_A_OcKfnYpe3_1(.din(G283), .dout(n11501));
    jdff dff_A_0daeuNOR1_1(.din(n11501), .dout(n11498));
    jdff dff_A_VPcXu3Td2_1(.din(n11498), .dout(n11495));
    jdff dff_A_UMyuYaC41_0(.din(G283), .dout(n11492));
    jdff dff_A_DcWhLFiX8_0(.din(n11492), .dout(n11489));
    jdff dff_A_bxpFVpxw1_0(.din(n11489), .dout(n11486));
    jdff dff_A_UWfbyl1h1_2(.din(n371), .dout(n11483));
    jdff dff_A_oJeBx24G4_0(.din(n371), .dout(n11480));
    jdff dff_A_9ngiHv6q8_0(.din(n11480), .dout(n11477));
    jdff dff_A_y8uCNX1z9_2(.din(n374), .dout(n11474));
    jdff dff_A_tJ7Qxpoe3_2(.din(n11474), .dout(n11471));
    jdff dff_A_Xo8Car738_2(.din(n11471), .dout(n11468));
    jdff dff_A_dZAaiECU3_2(.din(n374), .dout(n11465));
    jdff dff_A_hPOLBwJu3_2(.din(n11465), .dout(n11462));
    jdff dff_A_wGwwfJCx9_2(.din(n11462), .dout(n11459));
    jdff dff_A_p63nj3rN5_2(.din(n11459), .dout(n11456));
    jdff dff_A_ytpqUgnf0_1(.din(G97), .dout(n11453));
    jdff dff_A_0EFK6krm0_1(.din(n11453), .dout(n11450));
    jdff dff_A_jbusTZln6_1(.din(n11450), .dout(n11447));
    jdff dff_A_6yYBYou13_2(.din(G97), .dout(n11444));
    jdff dff_A_xewqMdmD6_2(.din(n11444), .dout(n11441));
    jdff dff_A_Yg7is76d4_2(.din(n11441), .dout(n11438));
    jdff dff_A_l8TPzBcC4_1(.din(G97), .dout(n11435));
    jdff dff_A_CueYVveM3_1(.din(n11435), .dout(n11432));
    jdff dff_A_WKeEDn6S5_1(.din(n11432), .dout(n11429));
    jdff dff_A_sDaQeqU74_0(.din(G97), .dout(n11426));
    jdff dff_B_QKp3wjYK2_1(.din(n11421), .dout(n11424));
    jdff dff_B_FzHTR9pu7_1(.din(n11418), .dout(n11421));
    jdff dff_B_ZZIFyYAI8_1(.din(n364), .dout(n11418));
    jdff dff_A_p1Lv5tZs8_2(.din(n191), .dout(n11414));
    jdff dff_A_6gcDyPwH1_2(.din(n11414), .dout(n11411));
    jdff dff_A_TB5hfQ0o8_1(.din(n191), .dout(n11408));
    jdff dff_A_AzWh0D143_1(.din(n11408), .dout(n11405));
    jdff dff_A_awxo882Y8_1(.din(n11405), .dout(n11402));
    jdff dff_A_qgWVCfvQ1_0(.din(n191), .dout(n11399));
    jdff dff_A_wyilZyJB0_0(.din(n11399), .dout(n11396));
    jdff dff_B_M2hcu2Iu9_0(.din(n11391), .dout(n11394));
    jdff dff_B_izbAE8qO7_0(.din(n398), .dout(n11391));
    jdff dff_A_agZidya10_1(.din(n406), .dout(n11387));
    jdff dff_A_N0M2Dwtu1_1(.din(n11387), .dout(n11384));
    jdff dff_A_Gi5qJDve0_1(.din(G169), .dout(n11381));
    jdff dff_A_Zd6KN2l20_1(.din(n11381), .dout(n11378));
    jdff dff_A_iyrgdOn12_1(.din(n11378), .dout(n11375));
    jdff dff_A_ON8lIAsy5_1(.din(n11375), .dout(n11372));
    jdff dff_A_yt34euw66_1(.din(n11372), .dout(n11369));
    jdff dff_A_lQQRhe7H8_1(.din(n11369), .dout(n11366));
    jdff dff_A_QgG4Hyin7_1(.din(n11366), .dout(n11363));
    jdff dff_A_GBIGJCYs5_0(.din(G169), .dout(n11360));
    jdff dff_A_53LigxUI3_1(.din(G169), .dout(n11357));
    jdff dff_A_WrA9bOyU1_1(.din(n11357), .dout(n11354));
    jdff dff_A_OEB2aHrV7_1(.din(n11354), .dout(n11351));
    jdff dff_A_9MtHASw25_1(.din(n11351), .dout(n11348));
    jdff dff_A_wP7iAD9G9_1(.din(n11348), .dout(n11345));
    jdff dff_A_SFIRQzNx1_1(.din(n11345), .dout(n11342));
    jdff dff_A_BVNBrHJ22_1(.din(n11342), .dout(n11339));
    jdff dff_A_XM8BCtkG6_1(.din(n11339), .dout(n11336));
    jdff dff_A_Ehupaxh00_1(.din(n412), .dout(n11333));
    jdff dff_A_RfddQYn10_0(.din(n333), .dout(n11330));
    jdff dff_A_F2uvRqSV5_0(.din(n11330), .dout(n11327));
    jdff dff_A_LwCLSk4Q9_0(.din(n11327), .dout(n11324));
    jdff dff_A_DdA5je7k2_0(.din(n11324), .dout(n11321));
    jdff dff_A_p9d7fzAb5_0(.din(n11321), .dout(n11318));
    jdff dff_A_4moNnSnd2_0(.din(n11318), .dout(n11315));
    jdff dff_A_fqjEorEV0_0(.din(n11315), .dout(n11312));
    jdff dff_A_XdMqc9jc1_0(.din(n11312), .dout(n11309));
    jdff dff_A_ei1SxWmQ4_0(.din(n11309), .dout(n11306));
    jdff dff_A_8yMCUGnd6_0(.din(n11306), .dout(n11303));
    jdff dff_A_H7Vs399g6_0(.din(n11303), .dout(n11300));
    jdff dff_A_duVIurAX0_0(.din(n11300), .dout(n11297));
    jdff dff_A_xCWnU4zI3_0(.din(n11297), .dout(n11294));
    jdff dff_A_pLAuYhxD6_0(.din(n11294), .dout(n11291));
    jdff dff_A_gw5ysKeH9_0(.din(n11291), .dout(n11288));
    jdff dff_A_MncSweYv9_0(.din(n11288), .dout(n11285));
    jdff dff_A_NeFbVxgv6_0(.din(n11285), .dout(n11282));
    jdff dff_A_jjyOFsE86_0(.din(n11282), .dout(n11279));
    jdff dff_A_gIp1idMr6_1(.din(G45), .dout(n11276));
    jdff dff_A_kNaDVNSq3_1(.din(n420), .dout(n11273));
    jdff dff_A_GSO5PdCL6_2(.din(G274), .dout(n11270));
    jdff dff_A_03ahk3n16_2(.din(n11270), .dout(n11267));
    jdff dff_A_NSZ2h9dl9_2(.din(n11267), .dout(n11264));
    jdff dff_A_u6jQZWCN8_0(.din(G274), .dout(n11261));
    jdff dff_A_yD4Oi5hU0_0(.din(n11261), .dout(n11258));
    jdff dff_A_XTFGpIVr3_1(.din(n427), .dout(n11255));
    jdff dff_B_j1gpmBTM4_3(.din(n439), .dout(n11253));
    jdff dff_A_YJlh3oE04_2(.din(n11253), .dout(n11249));
    jdff dff_A_rPcvYyJw0_2(.din(n446), .dout(n11246));
    jdff dff_A_4NqUh69t6_2(.din(n11246), .dout(n11243));
    jdff dff_A_a7OroNKR0_1(.din(n446), .dout(n11240));
    jdff dff_B_ynZ5YnHd1_1(.din(n144), .dout(n6381));
    jdff dff_B_xrbgYCPy3_1(.din(n6381), .dout(n6384));
    jdff dff_B_Pb9h1aHH6_1(.din(n6384), .dout(n6387));
    jdff dff_B_q71j2OGx8_0(.din(n225), .dout(n6390));
    jdff dff_B_udMr7RwF5_0(.din(n206), .dout(n6393));
    jdff dff_B_9z3KwyPI0_1(.din(n148), .dout(n6396));
    jdff dff_B_hbZGDMrg3_1(.din(n6396), .dout(n6399));
    jdff dff_B_zCONiVVC8_0(.din(n173), .dout(n6402));
    jdff dff_B_WG4S1uzv0_1(.din(n2013), .dout(n6405));
    jdff dff_B_e4hfOEbK7_1(.din(n6405), .dout(n6408));
    jdff dff_B_ZbTG51FI0_1(.din(n6408), .dout(n6411));
    jdff dff_B_t6YLDsJf6_1(.din(n6411), .dout(n6414));
    jdff dff_B_JHWAjE433_1(.din(n6414), .dout(n6417));
    jdff dff_B_Ws5GYjEw0_1(.din(n6417), .dout(n6420));
    jdff dff_B_xB1RSBq43_1(.din(n6420), .dout(n6423));
    jdff dff_B_rpt2txpk2_1(.din(n6423), .dout(n6426));
    jdff dff_B_CXcfAsYh9_1(.din(n6426), .dout(n6429));
    jdff dff_B_8FKXV26O9_1(.din(n6429), .dout(n6432));
    jdff dff_B_N9BGqFE76_1(.din(n6432), .dout(n6435));
    jdff dff_B_VtB1sIV48_1(.din(n6435), .dout(n6438));
    jdff dff_B_mL75RmLX6_1(.din(n6438), .dout(n6441));
    jdff dff_B_N6Lw2OXO1_1(.din(n6441), .dout(n6444));
    jdff dff_B_S51GjHWv7_1(.din(n6444), .dout(n6447));
    jdff dff_B_prADZb7W6_1(.din(n6447), .dout(n6450));
    jdff dff_B_fHOwcBxf0_0(.din(n2104), .dout(n6453));
    jdff dff_B_Jvtvvq538_0(.din(n6453), .dout(n6456));
    jdff dff_B_3M27IcLs1_0(.din(n6456), .dout(n6459));
    jdff dff_B_I7gb4k2j7_0(.din(n6459), .dout(n6462));
    jdff dff_B_Q0OU1C3u7_0(.din(n6462), .dout(n6465));
    jdff dff_B_cFVEODNb8_0(.din(n6465), .dout(n6468));
    jdff dff_B_jOwdAJi95_0(.din(n6468), .dout(n6471));
    jdff dff_B_1m3mqAGi7_0(.din(n6471), .dout(n6474));
    jdff dff_B_jnU9okez8_0(.din(n6474), .dout(n6477));
    jdff dff_B_oyimtRpZ0_0(.din(n6477), .dout(n6480));
    jdff dff_B_EAroxufK9_0(.din(n6480), .dout(n6483));
    jdff dff_B_0OMFfL6U4_0(.din(n6483), .dout(n6486));
    jdff dff_B_kUcR5PsM8_0(.din(n6486), .dout(n6489));
    jdff dff_B_mOPif1fF3_0(.din(n6489), .dout(n6492));
    jdff dff_B_bLAKcHKe6_0(.din(n2828), .dout(n6495));
    jdff dff_B_SPiR5Gfq0_0(.din(n6495), .dout(n6498));
    jdff dff_B_40lhxiL72_0(.din(n6498), .dout(n6501));
    jdff dff_B_U7NvSjUt8_0(.din(n6501), .dout(n6504));
    jdff dff_B_c7m59G2O8_0(.din(n6504), .dout(n6507));
    jdff dff_B_lUWwwYmu7_0(.din(n6507), .dout(n6510));
    jdff dff_B_H9wIZlfo4_0(.din(n6510), .dout(n6513));
    jdff dff_B_1EC4mkL36_0(.din(n6513), .dout(n6516));
    jdff dff_B_sNMgBzfb4_0(.din(n6516), .dout(n6519));
    jdff dff_B_dYU2wWJk4_0(.din(n6519), .dout(n6522));
    jdff dff_B_KCoETwj26_0(.din(n6522), .dout(n6525));
    jdff dff_B_347UTkUS3_0(.din(n6525), .dout(n6528));
    jdff dff_B_6RgXlCOo7_0(.din(n6528), .dout(n6531));
    jdff dff_B_huhjNFeY1_0(.din(n6531), .dout(n6534));
    jdff dff_B_1TU4w3Jl0_0(.din(n6534), .dout(n6537));
    jdff dff_B_fHVw0UMH6_0(.din(n6537), .dout(n6540));
    jdff dff_B_eyzArHIQ3_0(.din(n6540), .dout(n6543));
    jdff dff_B_sq671Pcx0_0(.din(n2824), .dout(n6546));
    jdff dff_A_rwvnvfyK3_1(.din(n6551), .dout(n6548));
    jdff dff_A_Gv04fcjb4_1(.din(n6554), .dout(n6551));
    jdff dff_A_fqJ0YkIr5_1(.din(n247), .dout(n6554));
    jdff dff_B_AVjPnWhX9_0(.din(n2812), .dout(n6558));
    jdff dff_B_KpnIjPAZ5_1(.din(n2700), .dout(n6561));
    jdff dff_B_TwPIIMOM4_1(.din(n6561), .dout(n6564));
    jdff dff_B_cYnRrgGN4_1(.din(n6564), .dout(n6567));
    jdff dff_B_QsOWg22Z7_1(.din(n6567), .dout(n6570));
    jdff dff_B_9puWg91t9_1(.din(n6570), .dout(n6573));
    jdff dff_B_pdUogo6x0_1(.din(n6573), .dout(n6576));
    jdff dff_B_7P58rKmj8_1(.din(n6576), .dout(n6579));
    jdff dff_B_k6DQEmqy0_1(.din(n6579), .dout(n6582));
    jdff dff_B_KAQ6kGp86_1(.din(n6582), .dout(n6585));
    jdff dff_B_mfgfwltP7_1(.din(n6585), .dout(n6588));
    jdff dff_B_IiyhBUHa3_1(.din(n6588), .dout(n6591));
    jdff dff_B_xGeWlfHP1_1(.din(n6591), .dout(n6594));
    jdff dff_B_F7txf4wl7_1(.din(n6594), .dout(n6597));
    jdff dff_B_FMWNkpb43_1(.din(n6597), .dout(n6600));
    jdff dff_B_rDYpXZLK3_1(.din(n6600), .dout(n6603));
    jdff dff_B_F6XMW7zK9_1(.din(n6603), .dout(n6606));
    jdff dff_B_mCBbpt9J8_1(.din(n6606), .dout(n6609));
    jdff dff_B_mirvIYcZ8_1(.din(n6609), .dout(n6612));
    jdff dff_B_NNpb1PAP1_0(.din(n2780), .dout(n6615));
    jdff dff_A_VV0G5Xfi3_0(.din(n217), .dout(n6617));
    jdff dff_B_MOGcl5UV4_1(.din(n4285), .dout(n6621));
    jdff dff_B_pLHv3hyp7_1(.din(n6621), .dout(n6624));
    jdff dff_B_HfCFKUce9_1(.din(n4288), .dout(n6627));
    jdff dff_B_oUye4lm36_1(.din(n6627), .dout(n6630));
    jdff dff_B_ccCmc88O3_1(.din(n6630), .dout(n6633));
    jdff dff_B_Oyyhcu7R7_1(.din(n6633), .dout(n6636));
    jdff dff_B_3yH9xtxp0_1(.din(n6636), .dout(n6639));
    jdff dff_B_fVa69rRd2_1(.din(n6639), .dout(n6642));
    jdff dff_B_ISIuAwLU4_1(.din(n6642), .dout(n6645));
    jdff dff_B_MiPcuc7d1_1(.din(n6645), .dout(n6648));
    jdff dff_B_i56ZNTFD4_1(.din(n6648), .dout(n6651));
    jdff dff_B_Yg9QwWVa5_1(.din(n6651), .dout(n6654));
    jdff dff_B_uh65DdRn2_1(.din(n6654), .dout(n6657));
    jdff dff_B_lkpLCRPL1_1(.din(n6657), .dout(n6660));
    jdff dff_B_OHSAB6HG1_1(.din(n6660), .dout(n6663));
    jdff dff_B_j1VOoZqi5_1(.din(n6663), .dout(n6666));
    jdff dff_B_LFokzkIg5_1(.din(n6666), .dout(n6669));
    jdff dff_B_GcFzOQHz3_1(.din(n6669), .dout(n6672));
    jdff dff_B_CP8Qiqn29_1(.din(n6672), .dout(n6675));
    jdff dff_B_ZhLnKxlj9_1(.din(n6675), .dout(n6678));
    jdff dff_B_CE4hUIpS1_1(.din(n6678), .dout(n6681));
    jdff dff_B_yqcq7O9G2_1(.din(n6681), .dout(n6684));
    jdff dff_B_FoniNyag2_1(.din(n6684), .dout(n6687));
    jdff dff_B_1tFGnpYG7_1(.din(n6687), .dout(n6690));
    jdff dff_B_iQ6wkzeT9_1(.din(n6690), .dout(n6693));
    jdff dff_B_bFmJ5DuS4_1(.din(n6693), .dout(n6696));
    jdff dff_B_HkKtItOb4_1(.din(n6696), .dout(n6699));
    jdff dff_B_LvvcfnQ51_1(.din(n6699), .dout(n6702));
    jdff dff_B_9RlCuJE84_1(.din(n6702), .dout(n6705));
    jdff dff_B_jy3F7UiK7_1(.din(n6705), .dout(n6708));
    jdff dff_B_NZyNgzld3_0(.din(n4267), .dout(n6711));
    jdff dff_B_HSI4VBVl1_0(.din(n4263), .dout(n6714));
    jdff dff_A_NlX6DN6V3_1(.din(n4248), .dout(n6716));
    jdff dff_B_4Jva4wWJ7_1(.din(n4327), .dout(n6720));
    jdff dff_B_Yp126YZE0_1(.din(n6720), .dout(n6723));
    jdff dff_B_WjTJ54NR6_1(.din(n6723), .dout(n6726));
    jdff dff_B_KxS9j7Ct8_1(.din(n6726), .dout(n6729));
    jdff dff_B_ooJVhPtl4_1(.din(n6729), .dout(n6732));
    jdff dff_B_Swa2GdbL7_1(.din(n6732), .dout(n6735));
    jdff dff_B_Gp7nP9S90_1(.din(n6735), .dout(n6738));
    jdff dff_B_XY1pnQ3s1_1(.din(n6738), .dout(n6741));
    jdff dff_B_JRXFOd4X2_1(.din(n6741), .dout(n6744));
    jdff dff_B_VWEfQuec5_1(.din(n6744), .dout(n6747));
    jdff dff_B_hkHyVgjx6_1(.din(n6747), .dout(n6750));
    jdff dff_B_ElenyalL8_1(.din(n6750), .dout(n6753));
    jdff dff_B_LL1UC17n5_1(.din(n6753), .dout(n6756));
    jdff dff_B_onvbfAJl0_1(.din(n6756), .dout(n6759));
    jdff dff_B_7GqXLUBk4_1(.din(n6759), .dout(n6762));
    jdff dff_B_TJrrlA0t2_1(.din(n6762), .dout(n6765));
    jdff dff_B_QJSsaXGL6_1(.din(n6765), .dout(n6768));
    jdff dff_B_AvtvG76D6_1(.din(n6768), .dout(n6771));
    jdff dff_B_4YD8iW2l7_1(.din(n6771), .dout(n6774));
    jdff dff_B_EZATfHu78_1(.din(n6774), .dout(n6777));
    jdff dff_B_rPPpTlqc4_1(.din(n6777), .dout(n6780));
    jdff dff_B_YTkb88oz0_1(.din(n6780), .dout(n6783));
    jdff dff_B_hRMMJKQr8_1(.din(n6783), .dout(n6786));
    jdff dff_B_0ug2eyZl8_1(.din(n6786), .dout(n6789));
    jdff dff_B_ep09lUf91_1(.din(n6789), .dout(n6792));
    jdff dff_B_tCTyTYsZ1_1(.din(G2897), .dout(n6795));
    jdff dff_B_nNZ0GruW3_1(.din(n6795), .dout(n6798));
    jdff dff_B_Sb1jYBl36_1(.din(n6798), .dout(n6801));
    jdff dff_B_FoKlvykA8_1(.din(n6801), .dout(n6804));
    jdff dff_B_92NfxHvE5_1(.din(n6804), .dout(n6807));
    jdff dff_B_akcrgVn10_1(.din(n6807), .dout(n6810));
    jdff dff_B_LkkgUbfh9_1(.din(n6810), .dout(n6813));
    jdff dff_B_DdU91plB6_1(.din(n6813), .dout(n6816));
    jdff dff_B_NkrRuS4v6_1(.din(n6816), .dout(n6819));
    jdff dff_B_kGzofVkP0_1(.din(n6819), .dout(n6822));
    jdff dff_B_FkDjUroM5_1(.din(n6822), .dout(n6825));
    jdff dff_B_a5qsdpPl0_1(.din(n6825), .dout(n6828));
    jdff dff_B_geszqRin9_1(.din(n6828), .dout(n6831));
    jdff dff_B_XPPkmska3_1(.din(n6831), .dout(n6834));
    jdff dff_B_q6xrlLHy0_1(.din(n6834), .dout(n6837));
    jdff dff_B_u4YvyHno2_1(.din(n6837), .dout(n6840));
    jdff dff_B_oiUAum5a2_1(.din(n6840), .dout(n6843));
    jdff dff_B_Dj4EA9br3_1(.din(n6843), .dout(n6846));
    jdff dff_B_AVlSSToM7_1(.din(n6846), .dout(n6849));
    jdff dff_B_2wh4DxzF3_1(.din(n6849), .dout(n6852));
    jdff dff_B_kqcm35Et6_1(.din(n6852), .dout(n6855));
    jdff dff_B_9Lneeevi3_1(.din(n6855), .dout(n6858));
    jdff dff_B_SccqQPVF0_1(.din(n6858), .dout(n6861));
    jdff dff_B_DpKEq05N3_1(.din(n6861), .dout(n6864));
    jdff dff_B_CkLQh78X3_1(.din(n6864), .dout(n6867));
    jdff dff_B_UM0Lkz9K1_1(.din(n6867), .dout(n6870));
    jdff dff_B_PsF3JsDJ6_1(.din(n6870), .dout(n6873));
    jdff dff_A_ILeDfsuw7_1(.din(n6878), .dout(n6875));
    jdff dff_A_pxawqQ3a3_1(.din(n6881), .dout(n6878));
    jdff dff_A_D2wsoZKF9_1(.din(n6884), .dout(n6881));
    jdff dff_A_Inn18rz07_1(.din(n6887), .dout(n6884));
    jdff dff_A_FXi9Q7wi5_1(.din(n6890), .dout(n6887));
    jdff dff_A_AIxfc44U1_1(.din(n6893), .dout(n6890));
    jdff dff_A_iS0tUClF8_1(.din(n6896), .dout(n6893));
    jdff dff_A_OXTVixPV4_1(.din(n6899), .dout(n6896));
    jdff dff_A_kx9jF2yE1_1(.din(n6902), .dout(n6899));
    jdff dff_A_f5EBb4x37_1(.din(n6905), .dout(n6902));
    jdff dff_A_KaqR2Yu58_1(.din(n6908), .dout(n6905));
    jdff dff_A_pEQqklk58_1(.din(n6911), .dout(n6908));
    jdff dff_A_PLmr5Ubr7_1(.din(n6914), .dout(n6911));
    jdff dff_A_fApyZn363_1(.din(n6917), .dout(n6914));
    jdff dff_A_sTXFaWHj3_1(.din(n6920), .dout(n6917));
    jdff dff_A_OmsWeqas0_1(.din(n6923), .dout(n6920));
    jdff dff_A_KKksWgzY0_1(.din(n6926), .dout(n6923));
    jdff dff_A_hFSP9obF9_1(.din(n6929), .dout(n6926));
    jdff dff_A_YzSysODz5_1(.din(n6932), .dout(n6929));
    jdff dff_A_YGXs8kLG2_1(.din(n6935), .dout(n6932));
    jdff dff_A_Q9MBdEoW4_1(.din(n6938), .dout(n6935));
    jdff dff_A_oiDLfZe90_1(.din(n6941), .dout(n6938));
    jdff dff_A_FqziWXfs7_1(.din(n6944), .dout(n6941));
    jdff dff_A_ZZi18SpG5_1(.din(n6947), .dout(n6944));
    jdff dff_A_HODbHNBK8_1(.din(n6950), .dout(n6947));
    jdff dff_A_cebzNpmp2_1(.din(n4312), .dout(n6950));
    jdff dff_A_5IgX0xir6_1(.din(n6956), .dout(n6953));
    jdff dff_A_vyPi09V38_1(.din(n6959), .dout(n6956));
    jdff dff_A_9BDr473e2_1(.din(n6962), .dout(n6959));
    jdff dff_A_5ynAQ5FP8_1(.din(n6965), .dout(n6962));
    jdff dff_A_3QWOje9G8_1(.din(n6968), .dout(n6965));
    jdff dff_A_Dw1jRvsm7_1(.din(n6971), .dout(n6968));
    jdff dff_A_rYyvzy0h3_1(.din(n6974), .dout(n6971));
    jdff dff_A_CK34gOZr6_1(.din(n6977), .dout(n6974));
    jdff dff_A_JoU1LoiZ6_1(.din(n6980), .dout(n6977));
    jdff dff_A_348Mxk9U0_1(.din(n6983), .dout(n6980));
    jdff dff_A_WvnTDaGw9_1(.din(n6986), .dout(n6983));
    jdff dff_A_Y29Mh8P43_1(.din(n6989), .dout(n6986));
    jdff dff_A_34Hh8ZaC5_1(.din(n6992), .dout(n6989));
    jdff dff_A_6j09Spgg0_1(.din(n6995), .dout(n6992));
    jdff dff_A_ksMFUMwP3_1(.din(n6998), .dout(n6995));
    jdff dff_A_MagO818t6_1(.din(n7001), .dout(n6998));
    jdff dff_A_VdYA3Qjv1_1(.din(n7004), .dout(n7001));
    jdff dff_A_mRX1fxRK9_1(.din(n7007), .dout(n7004));
    jdff dff_A_Zm5e9g7P5_1(.din(n7010), .dout(n7007));
    jdff dff_A_O5r1H6216_1(.din(n7013), .dout(n7010));
    jdff dff_A_1gOiWsKn6_1(.din(n7016), .dout(n7013));
    jdff dff_A_3dzdKn6K9_1(.din(n7019), .dout(n7016));
    jdff dff_A_agWKvC6d4_1(.din(n7022), .dout(n7019));
    jdff dff_A_6kZ25O5i0_1(.din(n7025), .dout(n7022));
    jdff dff_A_pKK2AQ8o9_1(.din(n7028), .dout(n7025));
    jdff dff_A_WWo1OGan9_1(.din(n4281), .dout(n7028));
    jdff dff_B_9IOKiBPx3_0(.din(n4062), .dout(n7032));
    jdff dff_B_AmBrGIhR0_0(.din(n7032), .dout(n7035));
    jdff dff_B_M6ZwTmD70_0(.din(n7035), .dout(n7038));
    jdff dff_B_8kcLwFOF0_0(.din(n7038), .dout(n7041));
    jdff dff_B_FXcr77hx2_0(.din(n7041), .dout(n7044));
    jdff dff_B_yGoT3d7y9_0(.din(n7044), .dout(n7047));
    jdff dff_B_yX29Iaal8_0(.din(n7047), .dout(n7050));
    jdff dff_B_2PGtm2bd1_0(.din(n4047), .dout(n7053));
    jdff dff_B_b2c5cbPb0_0(.din(n7053), .dout(n7056));
    jdff dff_B_etvtQCR71_0(.din(n7056), .dout(n7059));
    jdff dff_B_xIkmAwaF3_0(.din(n7059), .dout(n7062));
    jdff dff_B_14GPHnhZ5_0(.din(n7062), .dout(n7065));
    jdff dff_B_1bzYNzPb2_0(.din(n7065), .dout(n7068));
    jdff dff_B_LpNv12ZK0_0(.din(n7068), .dout(n7071));
    jdff dff_B_2YJIO6bP1_1(.din(n3896), .dout(n7074));
    jdff dff_B_TVj34eH45_1(.din(n7074), .dout(n7077));
    jdff dff_B_a2suvZFA7_1(.din(n7077), .dout(n7080));
    jdff dff_B_vCoqdJZO5_1(.din(n7080), .dout(n7083));
    jdff dff_B_qwclzErK5_1(.din(n7083), .dout(n7086));
    jdff dff_B_fmH78Oyd7_1(.din(n7086), .dout(n7089));
    jdff dff_B_WQ2yBKPr1_1(.din(n7089), .dout(n7092));
    jdff dff_B_jY1lzMXy0_1(.din(n7092), .dout(n7095));
    jdff dff_B_AgLcT7f60_1(.din(n3960), .dout(n7098));
    jdff dff_B_UcePQ7nO9_1(.din(n7098), .dout(n7101));
    jdff dff_B_6p2TD6t02_1(.din(n3990), .dout(n7104));
    jdff dff_B_vIG23IUk8_0(.din(n4010), .dout(n7107));
    jdff dff_B_PAQIdhXW3_1(.din(n3916), .dout(n7110));
    jdff dff_B_seMa3UNg8_1(.din(n7110), .dout(n7113));
    jdff dff_B_SRmOgYXh7_0(.din(n3952), .dout(n7116));
    jdff dff_B_q2JofDlD2_1(.din(n3920), .dout(n7119));
    jdff dff_B_TdsIXP264_0(.din(n3928), .dout(n7122));
    jdff dff_B_7SvklPTh7_1(.din(G124), .dout(n7125));
    jdff dff_B_eqVYmkLb8_1(.din(n7125), .dout(n7128));
    jdff dff_B_sDZ488Y14_1(.din(n7128), .dout(n7131));
    jdff dff_B_C7SLVvkC7_1(.din(n7131), .dout(n7134));
    jdff dff_B_dfAUOGxt2_1(.din(n3900), .dout(n7137));
    jdff dff_B_Vn3lvBwj6_0(.din(n3892), .dout(n7140));
    jdff dff_B_f72n7whF8_0(.din(n7140), .dout(n7143));
    jdff dff_B_dIaU5zlH8_0(.din(n7143), .dout(n7146));
    jdff dff_B_jIOqZmB33_1(.din(n3857), .dout(n7149));
    jdff dff_A_AQjdfNJy3_1(.din(n7154), .dout(n7151));
    jdff dff_A_RYql7SpD6_1(.din(n7157), .dout(n7154));
    jdff dff_A_M7cIU7oP7_1(.din(n7160), .dout(n7157));
    jdff dff_A_g66tHovf5_1(.din(n7163), .dout(n7160));
    jdff dff_A_OD4kqRMI8_1(.din(n7166), .dout(n7163));
    jdff dff_A_gBPuj7GC2_1(.din(n7169), .dout(n7166));
    jdff dff_A_4E3ZfTzQ6_1(.din(n7172), .dout(n7169));
    jdff dff_A_NvbC047F9_1(.din(n3865), .dout(n7172));
    jdff dff_B_t3YZ9YNv1_0(.din(n3861), .dout(n7176));
    jdff dff_B_QnLRwrnw8_0(.din(n7176), .dout(n7179));
    jdff dff_B_nCJnhmBj5_1(.din(n2707), .dout(n7182));
    jdff dff_B_6uSLkFyL4_1(.din(n7182), .dout(n7185));
    jdff dff_B_vXSWPy6C5_1(.din(n7185), .dout(n7188));
    jdff dff_B_SfkCUuyu4_1(.din(n7188), .dout(n7191));
    jdff dff_B_E6LEHatv5_1(.din(n7191), .dout(n7194));
    jdff dff_B_9mUJs9TO4_1(.din(n7194), .dout(n7197));
    jdff dff_B_uCU5BhTa0_1(.din(n7197), .dout(n7200));
    jdff dff_B_4HRWX6FB9_1(.din(n7200), .dout(n7203));
    jdff dff_A_Iys6T4A83_1(.din(n7208), .dout(n7205));
    jdff dff_A_i2Gbulu39_1(.din(n7211), .dout(n7208));
    jdff dff_A_JEo4JplL4_1(.din(n7302), .dout(n7211));
    jdff dff_B_MzbukCNK4_0(.din(n2703), .dout(n7215));
    jdff dff_B_s8dXbXUQ9_0(.din(n7215), .dout(n7218));
    jdff dff_B_qQRl7ORa8_0(.din(n7218), .dout(n7221));
    jdff dff_B_6xmW4B3f8_0(.din(n7221), .dout(n7224));
    jdff dff_B_mDHgUgxZ7_0(.din(n7224), .dout(n7227));
    jdff dff_B_uxtRcIsy7_0(.din(n7227), .dout(n7230));
    jdff dff_B_XZ06BLZb3_0(.din(n3849), .dout(n7233));
    jdff dff_B_soZKWZSH9_1(.din(n3730), .dout(n7236));
    jdff dff_B_DVJbvddl0_1(.din(n7236), .dout(n7239));
    jdff dff_B_t14mZ7Wt6_1(.din(n7239), .dout(n7242));
    jdff dff_B_TKIzkszB4_1(.din(n7242), .dout(n7245));
    jdff dff_B_YmC8U9uy1_1(.din(n7245), .dout(n7248));
    jdff dff_B_NEDV5Qq39_1(.din(n7248), .dout(n7251));
    jdff dff_B_O181L9ZS5_1(.din(n7251), .dout(n7254));
    jdff dff_B_4uF57oCj4_1(.din(n7254), .dout(n7257));
    jdff dff_B_1N7T31AP7_0(.din(n3822), .dout(n7260));
    jdff dff_A_L99Ypaxn3_1(.din(n7265), .dout(n7262));
    jdff dff_A_qSzqW1xY9_1(.din(n3800), .dout(n7265));
    jdff dff_B_Go0Z7t8Q7_1(.din(n2725), .dout(n7269));
    jdff dff_B_ED5gFEA37_1(.din(n7269), .dout(n7272));
    jdff dff_A_vvtvW8iE0_1(.din(n2740), .dout(n7274));
    jdff dff_A_XTyFZhMw1_1(.din(n7280), .dout(n7277));
    jdff dff_A_PocpNMT54_1(.din(n7283), .dout(n7280));
    jdff dff_A_Mo2Sva0V8_1(.din(n7286), .dout(n7283));
    jdff dff_A_Ney4EExm3_1(.din(n7302), .dout(n7286));
    jdff dff_A_ggCuepbO8_2(.din(n7292), .dout(n7289));
    jdff dff_A_mAfW15vs4_2(.din(n7295), .dout(n7292));
    jdff dff_A_z0M12BCP9_2(.din(n7302), .dout(n7295));
    jdff dff_B_nasyWk486_3(.din(n2718), .dout(n7299));
    jdff dff_B_p5X6eS3F5_3(.din(n7299), .dout(n7302));
    jdff dff_A_pXjCxg399_1(.din(n3792), .dout(n7304));
    jdff dff_B_B2gUorcj5_0(.din(n3723), .dout(n7308));
    jdff dff_B_6UKKzey64_0(.din(n3715), .dout(n7311));
    jdff dff_B_8GJiAsB33_0(.din(n7311), .dout(n7314));
    jdff dff_B_ELkhX7KN4_0(.din(n7314), .dout(n7317));
    jdff dff_B_t3fUfV9F2_0(.din(n7317), .dout(n7320));
    jdff dff_B_QKTeOl1e3_0(.din(n7320), .dout(n7323));
    jdff dff_B_m88xIWPw1_1(.din(n3648), .dout(n7326));
    jdff dff_B_8gPGC0Fu6_1(.din(n3664), .dout(n7329));
    jdff dff_B_AaXitViX9_0(.din(n3684), .dout(n7332));
    jdff dff_B_Jp6T2fN52_1(.din(n3668), .dout(n7335));
    jdff dff_B_CLm81odN6_1(.din(n3652), .dout(n7338));
    jdff dff_B_CkUcccqP4_1(.din(n3616), .dout(n7341));
    jdff dff_B_eEs0hkWs3_1(.din(n3620), .dout(n7344));
    jdff dff_B_4qBjV5F97_1(.din(n7344), .dout(n7347));
    jdff dff_B_8UkSvFVL7_1(.din(n7347), .dout(n7350));
    jdff dff_B_0ccWCGf52_1(.din(n3624), .dout(n7353));
    jdff dff_B_mpEZYCdW1_1(.din(n7353), .dout(n7356));
    jdff dff_B_qpyT6lIT2_0(.din(n3632), .dout(n7359));
    jdff dff_B_MemRcEoA6_1(.din(n3588), .dout(n7362));
    jdff dff_A_6fwpVXDc5_1(.din(n7374), .dout(n7364));
    jdff dff_B_kYAY9cCE3_2(.din(G125), .dout(n7368));
    jdff dff_B_DvAMv9hV5_2(.din(n7368), .dout(n7371));
    jdff dff_B_osGoo7l30_2(.din(n7371), .dout(n7374));
    jdff dff_A_ctnulHmK7_0(.din(n7379), .dout(n7376));
    jdff dff_A_wsO9wAL21_0(.din(n7382), .dout(n7379));
    jdff dff_A_peMkkoOB8_0(.din(n11747), .dout(n7382));
    jdff dff_A_lBHOKvxP8_1(.din(n7388), .dout(n7385));
    jdff dff_A_lN4oWSO32_1(.din(n7391), .dout(n7388));
    jdff dff_A_zJXLAHkh2_1(.din(n7394), .dout(n7391));
    jdff dff_A_6XkRdgC42_1(.din(n7397), .dout(n7394));
    jdff dff_A_UPHyR0D85_1(.din(n7400), .dout(n7397));
    jdff dff_A_IId9JDG40_1(.din(n7403), .dout(n7400));
    jdff dff_A_8vlSL97B9_1(.din(n7406), .dout(n7403));
    jdff dff_A_TkQ626Ep1_1(.din(n7409), .dout(n7406));
    jdff dff_A_Eq3uJins8_1(.din(n7412), .dout(n7409));
    jdff dff_A_e0sy6Ty21_1(.din(n7415), .dout(n7412));
    jdff dff_A_gps9NreM1_1(.din(n11747), .dout(n7415));
    jdff dff_B_kwjGrP3X0_0(.din(n2711), .dout(n7419));
    jdff dff_B_pgpnDPot6_0(.din(n7419), .dout(n7422));
    jdff dff_B_bbDuC9hg5_1(.din(n4222), .dout(n7425));
    jdff dff_B_tofmwiV27_1(.din(n7425), .dout(n7428));
    jdff dff_B_O2CbvBPK1_1(.din(n7428), .dout(n7431));
    jdff dff_B_Q26YwzAT5_1(.din(n7431), .dout(n7434));
    jdff dff_B_zb8rwFO40_1(.din(n7434), .dout(n7437));
    jdff dff_B_aPConhyT7_1(.din(n7437), .dout(n7440));
    jdff dff_B_DuplOqxG0_0(.din(n4233), .dout(n7443));
    jdff dff_B_wko8F1q72_1(.din(n4229), .dout(n7446));
    jdff dff_B_zOWbBvLs7_0(.din(n3734), .dout(n7449));
    jdff dff_A_obDpq9Wc4_0(.din(n1752), .dout(n7451));
    jdff dff_A_KtaDcr6o2_1(.din(n7457), .dout(n7454));
    jdff dff_A_YS7cNnUb6_1(.din(n1752), .dout(n7457));
    jdff dff_A_76GUKfTK9_2(.din(n7463), .dout(n7460));
    jdff dff_A_6ypzyubQ1_2(.din(n1752), .dout(n7463));
    jdff dff_A_Vep6fdi22_0(.din(n1933), .dout(n7466));
    jdff dff_B_codiG89P1_1(.din(n1907), .dout(n7470));
    jdff dff_B_a6D3DV1K1_1(.din(n7470), .dout(n7473));
    jdff dff_B_Xsm9xh5N4_1(.din(n1910), .dout(n7476));
    jdff dff_B_3wtckWVD5_1(.din(n7476), .dout(n7479));
    jdff dff_B_K3A7R6M86_1(.din(n7479), .dout(n7482));
    jdff dff_B_GHDibozC2_1(.din(n1913), .dout(n7485));
    jdff dff_A_vSDsysS30_0(.din(n1744), .dout(n7487));
    jdff dff_B_gWM7VLxp7_1(.din(n1472), .dout(n7491));
    jdff dff_A_W5Ogq3VP7_1(.din(n1710), .dout(n7493));
    jdff dff_A_I33LFH801_1(.din(n1694), .dout(n7496));
    jdff dff_A_JrOA0bvg9_1(.din(n7502), .dout(n7499));
    jdff dff_A_jLEg05hM1_1(.din(n7505), .dout(n7502));
    jdff dff_A_0KyCEXJH5_1(.din(n7508), .dout(n7505));
    jdff dff_A_JEG8Zf214_1(.din(n80), .dout(n7508));
    jdff dff_A_196A7o9u3_2(.din(n7514), .dout(n7511));
    jdff dff_A_XwUXAtVT4_2(.din(n7517), .dout(n7514));
    jdff dff_A_jI0YuI4j5_2(.din(n80), .dout(n7517));
    jdff dff_A_uPxZXOvn9_0(.din(n1676), .dout(n7520));
    jdff dff_B_eapyrZRK4_1(.din(n1649), .dout(n7524));
    jdff dff_B_s7xqtnNw8_1(.din(n1657), .dout(n7527));
    jdff dff_B_fPSynR9i2_1(.din(n7527), .dout(n7530));
    jdff dff_B_mDqj1ljP3_1(.din(n1642), .dout(n7533));
    jdff dff_B_IOgjobww9_1(.din(n7533), .dout(n7536));
    jdff dff_B_GY5YBRnb7_1(.din(n1604), .dout(n7539));
    jdff dff_B_uAVr2jzw7_1(.din(n7539), .dout(n7542));
    jdff dff_B_G3EgqqmC4_1(.din(n1608), .dout(n7545));
    jdff dff_A_n48ZFbuf3_1(.din(n1531), .dout(n7547));
    jdff dff_A_NLrLty692_0(.din(n1510), .dout(n7550));
    jdff dff_B_OKK6X1Xx9_1(.din(n1483), .dout(n7554));
    jdff dff_A_ETyHwJZZ6_0(.din(n7559), .dout(n7556));
    jdff dff_A_5GUiSh0H6_0(.din(n7562), .dout(n7559));
    jdff dff_A_0l8nIW9H9_0(.din(n77), .dout(n7562));
    jdff dff_A_o7WcTBV71_2(.din(n77), .dout(n7565));
    jdff dff_A_kLHkaF9J4_2(.din(n7571), .dout(n7568));
    jdff dff_A_PzhApn8n0_2(.din(n367), .dout(n7571));
    jdff dff_B_HPDhHTvl3_1(.din(n1431), .dout(n7575));
    jdff dff_A_Zh3LZqwt0_1(.din(n1452), .dout(n7577));
    jdff dff_A_Cqut5Hol2_0(.din(n1435), .dout(n7580));
    jdff dff_B_QuYqfTew0_2(.din(G223), .dout(n7584));
    jdff dff_B_zdMtXarI8_2(.din(n7584), .dout(n7587));
    jdff dff_A_nzPHUKnK0_0(.din(n7592), .dout(n7589));
    jdff dff_A_UbfmXpYv9_0(.din(n1428), .dout(n7592));
    jdff dff_A_MpttRNvE6_0(.din(n7598), .dout(n7595));
    jdff dff_A_VvKWeSn83_0(.din(n7602), .dout(n7598));
    jdff dff_B_IF4NufHq0_2(.din(n3841), .dout(n7602));
    jdff dff_A_UUzuMJy37_1(.din(n1133), .dout(n7604));
    jdff dff_A_FtBHihML4_0(.din(n7610), .dout(n7607));
    jdff dff_A_D96Dk9uZ6_0(.din(n7613), .dout(n7610));
    jdff dff_A_Z55c4btw4_0(.din(n2736), .dout(n7613));
    jdff dff_A_aZSTRNcR3_0(.din(n7619), .dout(n7616));
    jdff dff_A_Fv85uBtG6_0(.din(n7622), .dout(n7619));
    jdff dff_A_M6D2HWEZ2_0(.din(n7625), .dout(n7622));
    jdff dff_A_EPTeD56R1_0(.din(n2733), .dout(n7625));
    jdff dff_B_wMi9uOsJ9_0(.din(n3748), .dout(n7629));
    jdff dff_B_4ZkfhsuZ8_0(.din(n7629), .dout(n7632));
    jdff dff_B_Uz0lf2br0_0(.din(n7632), .dout(n7635));
    jdff dff_B_CrutxyLd1_0(.din(n4211), .dout(n7638));
    jdff dff_B_kSpOWxbn2_0(.din(n7638), .dout(n7641));
    jdff dff_B_pgnI3aQB0_0(.din(n7641), .dout(n7644));
    jdff dff_B_PQ6gA8B69_0(.din(n4207), .dout(n7647));
    jdff dff_B_EGXmiC7J3_0(.din(n7647), .dout(n7650));
    jdff dff_B_kfpXk8sW5_0(.din(n7650), .dout(n7653));
    jdff dff_B_hFunX7DE5_0(.din(n7653), .dout(n7656));
    jdff dff_B_Alqur92y5_0(.din(n7656), .dout(n7659));
    jdff dff_B_mz2u4UQD9_1(.din(n4132), .dout(n7662));
    jdff dff_B_UeGz7vFO4_1(.din(n7662), .dout(n7665));
    jdff dff_B_VI8urFpX0_1(.din(n4136), .dout(n7668));
    jdff dff_B_qI34WO6Q9_1(.din(n7668), .dout(n7671));
    jdff dff_B_WtBCHLNl5_1(.din(n7671), .dout(n7674));
    jdff dff_B_I96gKeLI7_1(.din(n7674), .dout(n7677));
    jdff dff_B_OckltRcT2_1(.din(n7677), .dout(n7680));
    jdff dff_B_cBcHvVMM1_1(.din(n4148), .dout(n7683));
    jdff dff_B_c4620I9v0_1(.din(n7683), .dout(n7686));
    jdff dff_B_PXEpW0aS6_1(.din(n7686), .dout(n7689));
    jdff dff_B_KZ9JUhvf0_1(.din(n4168), .dout(n7692));
    jdff dff_A_YWRtBQ7V5_0(.din(n7704), .dout(n7694));
    jdff dff_B_W3iuT2RV1_3(.din(G128), .dout(n7698));
    jdff dff_B_8O9yucme6_3(.din(n7698), .dout(n7701));
    jdff dff_B_aXjaDQ4M0_3(.din(n7701), .dout(n7704));
    jdff dff_A_5O647Yik4_0(.din(n9797), .dout(n7706));
    jdff dff_A_2F2Oudh08_1(.din(n7712), .dout(n7709));
    jdff dff_A_XtQxDIXw9_1(.din(n7715), .dout(n7712));
    jdff dff_A_LOuZt1hJ2_1(.din(n7718), .dout(n7715));
    jdff dff_A_90HwEfKC6_1(.din(n9797), .dout(n7718));
    jdff dff_B_FptpMnwi7_1(.din(n4152), .dout(n7722));
    jdff dff_B_JeNg2Ljz2_1(.din(n7722), .dout(n7725));
    jdff dff_A_0yyXrzMH2_0(.din(n3979), .dout(n7727));
    jdff dff_A_JIa7x4XB8_1(.din(n8849), .dout(n7730));
    jdff dff_A_oAPZEv3J5_2(.din(n10244), .dout(n7733));
    jdff dff_B_YPROuvuL0_1(.din(n4080), .dout(n7737));
    jdff dff_B_JxhsXLS99_1(.din(n7737), .dout(n7740));
    jdff dff_A_bvHEwYPn0_1(.din(n11504), .dout(n7742));
    jdff dff_A_NcO9Sjbo1_2(.din(n7748), .dout(n7745));
    jdff dff_A_6eiINvJZ3_2(.din(n7751), .dout(n7748));
    jdff dff_A_mdZgBqlb2_2(.din(n7754), .dout(n7751));
    jdff dff_A_TJwIehfe4_2(.din(n2733), .dout(n7754));
    jdff dff_B_5c9wZdRa0_0(.din(n2729), .dout(n7758));
    jdff dff_B_IWopkhLh1_0(.din(n7758), .dout(n7761));
    jdff dff_B_ZNbHQtQH4_0(.din(n7761), .dout(n7764));
    jdff dff_B_hQIfFVma4_0(.din(n7764), .dout(n7767));
    jdff dff_A_FcdkyXoc5_1(.din(n1397), .dout(n7769));
    jdff dff_A_Oh91G41R4_1(.din(n1385), .dout(n7772));
    jdff dff_A_SKxkA4gY1_2(.din(n1385), .dout(n7775));
    jdff dff_B_9sgztSk90_1(.din(n1361), .dout(n7779));
    jdff dff_B_bH0fzxpY2_1(.din(n7779), .dout(n7782));
    jdff dff_B_mqMdDvCO3_1(.din(n1369), .dout(n7785));
    jdff dff_B_BhPBEMs71_1(.din(n7785), .dout(n7788));
    jdff dff_A_MchgcMM65_0(.din(n7793), .dout(n7790));
    jdff dff_A_vb2mpHcf6_0(.din(G68), .dout(n7793));
    jdff dff_A_SfnC8UI12_2(.din(n7799), .dout(n7796));
    jdff dff_A_0msoXEw23_2(.din(n7802), .dout(n7799));
    jdff dff_A_IMx4AmGF3_2(.din(n7805), .dout(n7802));
    jdff dff_A_gwvRXqe98_2(.din(n7808), .dout(n7805));
    jdff dff_A_OE7sgIuQ1_2(.din(G68), .dout(n7808));
    jdff dff_B_lrgl6soP5_0(.din(n1365), .dout(n7812));
    jdff dff_A_xc49V2yN9_1(.din(n1345), .dout(n7814));
    jdff dff_B_Vz7Z6xjQ8_1(.din(n1306), .dout(n7818));
    jdff dff_B_947c0t5M6_1(.din(n7818), .dout(n7821));
    jdff dff_B_EwVOvqLO1_1(.din(n1310), .dout(n7824));
    jdff dff_A_ZrygzSyX5_0(.din(n7829), .dout(n7826));
    jdff dff_A_9QBz8RYs5_0(.din(n431), .dout(n7829));
    jdff dff_A_e5E483ow0_0(.din(n7835), .dout(n7832));
    jdff dff_A_Q2U1rWYC3_0(.din(n7838), .dout(n7835));
    jdff dff_A_UDsUAlsV2_0(.din(n2693), .dout(n7838));
    jdff dff_A_g5xzbAJs4_0(.din(n7844), .dout(n7841));
    jdff dff_A_vgLnRoeq5_0(.din(n7847), .dout(n7844));
    jdff dff_A_UydSEI1R7_0(.din(n7850), .dout(n7847));
    jdff dff_A_akZQpuOp2_0(.din(n2690), .dout(n7850));
    jdff dff_B_rh4QLE558_1(.din(n2643), .dout(n7854));
    jdff dff_B_WE9fOSRN4_1(.din(n7854), .dout(n7857));
    jdff dff_B_UcjOiyLY9_0(.din(n2658), .dout(n7860));
    jdff dff_B_7B0RoYiB7_1(.din(n920), .dout(n7863));
    jdff dff_A_EmMFb6Ux0_0(.din(n7868), .dout(n7865));
    jdff dff_A_zDloW7fa1_0(.din(n7871), .dout(n7868));
    jdff dff_A_YTi8Dgu26_0(.din(n1298), .dout(n7871));
    jdff dff_B_hVfg89iI1_0(.din(n2636), .dout(n7875));
    jdff dff_B_yiifLGK53_0(.din(n7875), .dout(n7878));
    jdff dff_B_vhBtoQwU7_0(.din(n7878), .dout(n7881));
    jdff dff_B_iNYb9PqW3_0(.din(n7881), .dout(n7884));
    jdff dff_B_6axqDvYD6_0(.din(n2628), .dout(n7887));
    jdff dff_B_a4VQMPiO2_0(.din(n7887), .dout(n7890));
    jdff dff_B_yOlpVy2k4_0(.din(n7890), .dout(n7893));
    jdff dff_B_vaDBoLY89_0(.din(n7893), .dout(n7896));
    jdff dff_B_QeiMDT8I5_1(.din(n2617), .dout(n7899));
    jdff dff_A_czxibepF3_0(.din(n7904), .dout(n7901));
    jdff dff_A_YimUmIaL6_0(.din(n7907), .dout(n7904));
    jdff dff_A_40nzIkoe9_0(.din(n7910), .dout(n7907));
    jdff dff_A_yXd4Uuu18_0(.din(n7913), .dout(n7910));
    jdff dff_A_YXZheSm79_0(.din(n7916), .dout(n7913));
    jdff dff_A_D0lwcCld0_0(.din(n7919), .dout(n7916));
    jdff dff_A_QGPlReu91_0(.din(n7922), .dout(n7919));
    jdff dff_A_82kfVSlJ5_0(.din(n7925), .dout(n7922));
    jdff dff_A_vqqHyQld4_0(.din(n7928), .dout(n7925));
    jdff dff_A_SCvhVDYY6_0(.din(n7931), .dout(n7928));
    jdff dff_A_vp9rvH7c9_0(.din(n2146), .dout(n7931));
    jdff dff_A_xgxKAMrc7_1(.din(n7937), .dout(n7934));
    jdff dff_A_W6tDfEn78_1(.din(n7940), .dout(n7937));
    jdff dff_A_sWjbEFMw4_1(.din(n7943), .dout(n7940));
    jdff dff_A_3WDz4osr6_1(.din(n7946), .dout(n7943));
    jdff dff_A_xlixRGKu3_1(.din(n7949), .dout(n7946));
    jdff dff_A_VM8dThXw0_1(.din(n7952), .dout(n7949));
    jdff dff_A_pOrw0prw5_1(.din(n7955), .dout(n7952));
    jdff dff_A_eWucBi366_1(.din(n7958), .dout(n7955));
    jdff dff_A_u5hNhmDB3_1(.din(n7961), .dout(n7958));
    jdff dff_A_Dz7BMP8p7_1(.din(n7964), .dout(n7961));
    jdff dff_A_om1uan588_1(.din(n2146), .dout(n7964));
    jdff dff_B_OhgEfmRx3_0(.din(n2598), .dout(n7968));
    jdff dff_B_c4JQbR9H5_0(.din(n2562), .dout(n7971));
    jdff dff_B_Qgk1zIAq1_1(.din(n2550), .dout(n7974));
    jdff dff_B_oCrH7Lgx0_1(.din(n2510), .dout(n7977));
    jdff dff_B_LPi0uogA1_1(.din(n2522), .dout(n7980));
    jdff dff_A_n5GY4sdo6_0(.din(n7985), .dout(n7982));
    jdff dff_A_9ipMDwCo7_0(.din(n7988), .dout(n7985));
    jdff dff_A_1uyzNcr30_0(.din(n7991), .dout(n7988));
    jdff dff_A_tpD3wjjN6_0(.din(n7995), .dout(n7991));
    jdff dff_B_5UdxwxRG3_2(.din(n2530), .dout(n7995));
    jdff dff_B_l3j8OZvY8_1(.din(n2514), .dout(n7998));
    jdff dff_A_97lxGxD29_1(.din(n8010), .dout(n8000));
    jdff dff_B_WfF5hDW57_3(.din(G132), .dout(n8004));
    jdff dff_B_wPFcyzwI9_3(.din(n8004), .dout(n8007));
    jdff dff_B_EDPlRGQZ8_3(.din(n8007), .dout(n8010));
    jdff dff_B_yO4odglo3_1(.din(n2486), .dout(n8013));
    jdff dff_B_CsOHDHJM3_1(.din(n8013), .dout(n8016));
    jdff dff_B_0YsiHeIC6_0(.din(n2502), .dout(n8019));
    jdff dff_A_nbkZK3gz7_0(.din(n8859), .dout(n8021));
    jdff dff_A_226JHW4E9_0(.din(n8027), .dout(n8024));
    jdff dff_A_JH3Amltv7_0(.din(n2475), .dout(n8027));
    jdff dff_A_TXIsUPNy8_0(.din(n8033), .dout(n8030));
    jdff dff_A_39XrxDvY6_0(.din(n8036), .dout(n8033));
    jdff dff_A_iOdcPdRN2_0(.din(n2472), .dout(n8036));
    jdff dff_A_mjcIPlYI2_1(.din(n8042), .dout(n8039));
    jdff dff_A_W95K5KKG3_1(.din(n8045), .dout(n8042));
    jdff dff_A_ByPGuawY7_1(.din(n2472), .dout(n8045));
    jdff dff_A_qHvtVqkT7_2(.din(n2472), .dout(n8048));
    jdff dff_B_vI1890VH2_0(.din(n2468), .dout(n8052));
    jdff dff_B_gmxxOQzu0_0(.din(n8052), .dout(n8055));
    jdff dff_B_tIvO4YzW4_0(.din(n8055), .dout(n8058));
    jdff dff_B_oEGQHARh0_0(.din(n8058), .dout(n8061));
    jdff dff_B_LzxIiMpc8_0(.din(n8061), .dout(n8064));
    jdff dff_A_sdMQGsvz6_0(.din(n10838), .dout(n8066));
    jdff dff_A_ruwX4sgZ3_1(.din(n8072), .dout(n8069));
    jdff dff_A_wWlgZZ4S2_1(.din(n8075), .dout(n8072));
    jdff dff_A_RLsYC9xP9_1(.din(n8078), .dout(n8075));
    jdff dff_A_t9pnQjqb7_1(.din(n8081), .dout(n8078));
    jdff dff_A_1cZgT8FT3_1(.din(n8084), .dout(n8081));
    jdff dff_A_aYTPkeyl4_1(.din(n8087), .dout(n8084));
    jdff dff_A_dTjGelrD5_1(.din(n10838), .dout(n8087));
    jdff dff_A_LR5W7OFQ5_1(.din(n10280), .dout(n8090));
    jdff dff_B_qhibm7nF7_1(.din(n1257), .dout(n8094));
    jdff dff_B_IAH45NQo8_1(.din(n8094), .dout(n8097));
    jdff dff_A_UZ27vMAF8_1(.din(n8102), .dout(n8099));
    jdff dff_A_GdC3iBAj1_1(.din(n8105), .dout(n8102));
    jdff dff_A_PSySrwr68_1(.din(n1254), .dout(n8105));
    jdff dff_B_2DwCmg7O1_1(.din(n1220), .dout(n8109));
    jdff dff_B_2c83vRPV0_0(.din(n1246), .dout(n8112));
    jdff dff_B_aEtb0mcV1_1(.din(n1227), .dout(n8115));
    jdff dff_A_pgfK9uma1_0(.din(n1234), .dout(n8117));
    jdff dff_A_34WEawZK6_0(.din(n8124), .dout(n8120));
    jdff dff_B_gHQTSLrz0_2(.din(n1204), .dout(n8124));
    jdff dff_B_jLV0ghFw1_0(.din(n1185), .dout(n8127));
    jdff dff_B_pGicBI5G6_1(.din(n1158), .dout(n8130));
    jdff dff_A_jxVQlUsh1_1(.din(n8135), .dout(n8132));
    jdff dff_A_u0zShoW77_1(.din(n1154), .dout(n8135));
    jdff dff_A_Mi458JfJ5_0(.din(n1151), .dout(n8138));
    jdff dff_A_LB2BJLy78_1(.din(n1151), .dout(n8141));
    jdff dff_A_CwoR9y7N7_2(.din(n1151), .dout(n8144));
    jdff dff_A_uEuoVxFA7_0(.din(n1144), .dout(n8147));
    jdff dff_A_NDct26XZ8_1(.din(n1144), .dout(n8150));
    jdff dff_A_zzA9gOhC2_2(.din(n1144), .dout(n8153));
    jdff dff_A_7H2DEj1c7_1(.din(n8159), .dout(n8156));
    jdff dff_A_Lz3Y5PGp7_1(.din(n8166), .dout(n8159));
    jdff dff_B_hpwzkZhz7_2(.din(n4308), .dout(n8163));
    jdff dff_B_Dq2Xk9Zs5_2(.din(n8163), .dout(n8166));
    jdff dff_B_cRQ7BKJr4_1(.din(n4300), .dout(n8169));
    jdff dff_B_76G1R80I7_1(.din(n3396), .dout(n8172));
    jdff dff_B_MW8Bjtcc4_0(.din(n3566), .dout(n8175));
    jdff dff_B_EEa8Na864_0(.din(n8175), .dout(n8178));
    jdff dff_B_lnQ8HUb74_0(.din(n8178), .dout(n8181));
    jdff dff_B_L79gYsFG0_0(.din(n8181), .dout(n8184));
    jdff dff_B_JC0CyPB34_0(.din(n8184), .dout(n8187));
    jdff dff_B_gNQYeVZj1_0(.din(n3559), .dout(n8190));
    jdff dff_B_Og2VNfOO6_0(.din(n8190), .dout(n8193));
    jdff dff_B_Q6ihH8472_1(.din(n3423), .dout(n8196));
    jdff dff_B_p0uyDgDK6_1(.din(n8196), .dout(n8199));
    jdff dff_B_LpW2euEs6_1(.din(n8199), .dout(n8202));
    jdff dff_B_7g4tZBYO7_1(.din(n8202), .dout(n8205));
    jdff dff_B_7whsfyG25_1(.din(n3495), .dout(n8208));
    jdff dff_B_Y3pctb3y9_1(.din(n3523), .dout(n8211));
    jdff dff_A_cUW9NY2e1_2(.din(n11615), .dout(n8213));
    jdff dff_B_QGb6dHNc8_1(.din(n3487), .dout(n8217));
    jdff dff_A_p726uaCi3_1(.din(n10088), .dout(n8219));
    jdff dff_B_oesYkrT41_1(.din(n3435), .dout(n8223));
    jdff dff_B_1o1k8E266_1(.din(n8223), .dout(n8226));
    jdff dff_B_2fzj4tTD7_1(.din(n8226), .dout(n8229));
    jdff dff_B_00tOmlcV1_1(.din(n3447), .dout(n8232));
    jdff dff_B_yRAbqoPj3_1(.din(n8232), .dout(n8235));
    jdff dff_B_3538W6Se4_1(.din(n3455), .dout(n8238));
    jdff dff_A_n1qPfFTw9_0(.din(n8243), .dout(n8240));
    jdff dff_A_ceXLqub56_0(.din(n8246), .dout(n8243));
    jdff dff_A_AvSlXyCe7_0(.din(n3463), .dout(n8246));
    jdff dff_A_0FXdgbTT2_2(.din(n8457), .dout(n8249));
    jdff dff_A_Fweb03Sm6_1(.din(n8255), .dout(n8252));
    jdff dff_A_zkS5FPqg8_1(.din(n8258), .dout(n8255));
    jdff dff_A_N4Y2Mr3N2_1(.din(G50), .dout(n8258));
    jdff dff_A_0JtXnC2e8_2(.din(n8264), .dout(n8261));
    jdff dff_A_q93wIPSs7_2(.din(n8267), .dout(n8264));
    jdff dff_A_nLJPHWsy8_2(.din(G50), .dout(n8267));
    jdff dff_B_lm0hFwU34_1(.din(n3411), .dout(n8271));
    jdff dff_B_LY7bYntw8_1(.din(n8271), .dout(n8274));
    jdff dff_B_AwPZqyvy3_0(.din(n3415), .dout(n8277));
    jdff dff_A_NxLNoeNl9_0(.din(n314), .dout(n8279));
    jdff dff_B_DZJ2aS4s0_0(.din(n310), .dout(n8283));
    jdff dff_B_bmkZyDxZ1_1(.din(n3385), .dout(n8286));
    jdff dff_B_JvjjaOGR2_1(.din(n3017), .dout(n8289));
    jdff dff_B_P5QO7Brl0_1(.din(n8289), .dout(n8292));
    jdff dff_B_wnA5m0lB7_1(.din(n8292), .dout(n8295));
    jdff dff_B_vujsMn4w8_1(.din(n8295), .dout(n8298));
    jdff dff_B_pMhcoQm33_1(.din(n8298), .dout(n8301));
    jdff dff_B_u5krdrV44_1(.din(n8301), .dout(n8304));
    jdff dff_B_vSBWEpvC8_1(.din(n8304), .dout(n8307));
    jdff dff_B_DrZ5NFFL2_1(.din(n3068), .dout(n8310));
    jdff dff_B_EYZKU5ko9_1(.din(n8310), .dout(n8313));
    jdff dff_B_2qZ3BbhQ9_0(.din(n3106), .dout(n8316));
    jdff dff_A_ufV6lJRQ8_0(.din(n8321), .dout(n8318));
    jdff dff_A_oowgKUsw6_0(.din(n8324), .dout(n8321));
    jdff dff_A_lbuSIHpA8_0(.din(n3094), .dout(n8324));
    jdff dff_A_gfTtQOA63_2(.din(n3094), .dout(n8327));
    jdff dff_B_YAk8KxDc6_1(.din(n3032), .dout(n8331));
    jdff dff_B_FRUsGpKl3_1(.din(n3036), .dout(n8334));
    jdff dff_B_500HLwzz0_1(.din(n8334), .dout(n8337));
    jdff dff_B_8phYCkmE0_1(.din(n8337), .dout(n8340));
    jdff dff_B_ZAfep1yA9_1(.din(n8340), .dout(n8343));
    jdff dff_B_drb9tgyI3_0(.din(n3048), .dout(n8346));
    jdff dff_A_6SXdzCnI2_1(.din(n8351), .dout(n8348));
    jdff dff_A_WfzRtcFC0_1(.din(n1959), .dout(n8351));
    jdff dff_A_CrFou7NL0_0(.din(n1121), .dout(n8354));
    jdff dff_A_AcbZ4Tay0_0(.din(n8360), .dout(n8357));
    jdff dff_A_JS0Y1SzS9_0(.din(n1064), .dout(n8360));
    jdff dff_B_tascgUPq3_0(.din(n3028), .dout(n8364));
    jdff dff_B_olPxfAgE5_0(.din(n8364), .dout(n8367));
    jdff dff_A_zBDMi8J16_1(.din(n8372), .dout(n8369));
    jdff dff_A_41v9qUwg2_1(.din(n8375), .dout(n8372));
    jdff dff_A_jsVmobp23_1(.din(n8378), .dout(n8375));
    jdff dff_A_OG8upKwM1_1(.din(n3025), .dout(n8378));
    jdff dff_B_tDkrTTgd8_0(.din(n3021), .dout(n8382));
    jdff dff_B_XrN8ujoq0_0(.din(n8382), .dout(n8385));
    jdff dff_B_JiavlIFh1_0(.din(n8385), .dout(n8388));
    jdff dff_A_yxo8XTQb4_1(.din(n8393), .dout(n8390));
    jdff dff_A_nBTj7VM28_1(.din(n1997), .dout(n8393));
    jdff dff_B_reR9chzK7_0(.din(n3010), .dout(n8397));
    jdff dff_B_lryXG1jZ6_1(.din(n2870), .dout(n8400));
    jdff dff_B_dnmNCXeR4_1(.din(n8400), .dout(n8403));
    jdff dff_B_tbPUkQaw0_1(.din(n8403), .dout(n8406));
    jdff dff_B_3oQ96Ro83_1(.din(n2946), .dout(n8409));
    jdff dff_B_PwACYx4m9_1(.din(n8409), .dout(n8412));
    jdff dff_B_wcfSg0N25_1(.din(n2958), .dout(n8415));
    jdff dff_B_RxJFYEeT9_1(.din(n8415), .dout(n8418));
    jdff dff_B_evK5ALlS6_0(.din(n2982), .dout(n8421));
    jdff dff_A_1gSwhNQf5_0(.din(n2978), .dout(n8423));
    jdff dff_B_xumulVta2_1(.din(n2962), .dout(n8427));
    jdff dff_A_RooK4Q3D0_0(.din(n8432), .dout(n8429));
    jdff dff_A_bG2djZ6W8_0(.din(n8435), .dout(n8432));
    jdff dff_A_QDZZMnUA1_0(.din(G58), .dout(n8435));
    jdff dff_A_YJiz5Z9H3_2(.din(n8441), .dout(n8438));
    jdff dff_A_3ZEmc1Qq4_2(.din(n8444), .dout(n8441));
    jdff dff_A_GR0woiLp9_2(.din(n8447), .dout(n8444));
    jdff dff_A_ziTFnVBC9_2(.din(G58), .dout(n8447));
    jdff dff_B_OSTqnc9o9_3(.din(G143), .dout(n8451));
    jdff dff_B_yZBK22iS5_3(.din(n8451), .dout(n8454));
    jdff dff_B_2fQBAMhR4_3(.din(n8454), .dout(n8457));
    jdff dff_B_J4G9mpnt1_1(.din(n2938), .dout(n8460));
    jdff dff_A_8cGpDfv52_1(.din(n8472), .dout(n8462));
    jdff dff_B_3A6t9QDM7_3(.din(G137), .dout(n8466));
    jdff dff_B_Ux9afbeq9_3(.din(n8466), .dout(n8469));
    jdff dff_B_24faEiGY7_3(.din(n8469), .dout(n8472));
    jdff dff_B_Pa7mNo931_1(.din(n2882), .dout(n8475));
    jdff dff_B_E0lqSfHI1_1(.din(n8475), .dout(n8478));
    jdff dff_B_ITBo9cRh8_1(.din(n8478), .dout(n8481));
    jdff dff_B_tBpgZeHR6_1(.din(n2894), .dout(n8484));
    jdff dff_B_IcFqzFcb4_1(.din(n8484), .dout(n8487));
    jdff dff_A_GugwOcEI1_1(.din(n10181), .dout(n8489));
    jdff dff_B_ORF3evCs4_1(.din(n2898), .dout(n8493));
    jdff dff_A_s7wx6l3t2_0(.din(n8498), .dout(n8495));
    jdff dff_A_Hn3xa1Rf4_0(.din(n8501), .dout(n8498));
    jdff dff_A_HKxft28O8_0(.din(n8504), .dout(n8501));
    jdff dff_A_TQ8QPLsV9_0(.din(n8507), .dout(n8504));
    jdff dff_A_oyhoAt5v5_0(.din(n8510), .dout(n8507));
    jdff dff_A_XaaQSeDR1_0(.din(n8513), .dout(n8510));
    jdff dff_A_GbYdWwlj5_0(.din(n2384), .dout(n8513));
    jdff dff_A_UNfPpoSj7_2(.din(n8519), .dout(n8516));
    jdff dff_A_xDs9WJzV1_2(.din(n8522), .dout(n8519));
    jdff dff_A_JMSQkLdp9_2(.din(n8525), .dout(n8522));
    jdff dff_A_1xwARsnp4_2(.din(n8528), .dout(n8525));
    jdff dff_A_n8K1NTCA0_2(.din(n8531), .dout(n8528));
    jdff dff_A_JmyOfB7B1_2(.din(n2384), .dout(n8531));
    jdff dff_B_3EdAInlv4_1(.din(n2851), .dout(n8535));
    jdff dff_B_9kC6cd7E5_1(.din(n8535), .dout(n8538));
    jdff dff_B_jHdHPdUh9_0(.din(n2858), .dout(n8541));
    jdff dff_A_oZ09gIbv8_0(.din(n271), .dout(n8543));
    jdff dff_B_PHRg72GV4_0(.din(n267), .dout(n8547));
    jdff dff_A_f2O2TfQE2_1(.din(n8552), .dout(n8549));
    jdff dff_A_ROk1wMdd7_1(.din(n8555), .dout(n8552));
    jdff dff_A_O1iMba9j5_1(.din(n8558), .dout(n8555));
    jdff dff_A_N5L1lzpW5_1(.din(n8561), .dout(n8558));
    jdff dff_A_QjXIX3JX3_1(.din(n8564), .dout(n8561));
    jdff dff_A_q4424rMo6_1(.din(n8567), .dout(n8564));
    jdff dff_A_qQHdypN76_1(.din(n8570), .dout(n8567));
    jdff dff_A_p8ELpzs83_1(.din(n8573), .dout(n8570));
    jdff dff_A_NPPMvooM8_1(.din(n8576), .dout(n8573));
    jdff dff_A_zsDmacJB5_1(.din(n8579), .dout(n8576));
    jdff dff_A_7SMRNitG2_1(.din(n8582), .dout(n8579));
    jdff dff_A_aBqoN1gC4_1(.din(n11708), .dout(n8582));
    jdff dff_A_rhnNNtjf9_2(.din(n8588), .dout(n8585));
    jdff dff_A_TuA7yQBL6_2(.din(n8591), .dout(n8588));
    jdff dff_A_U4G2hbYB4_2(.din(n8594), .dout(n8591));
    jdff dff_A_VZajrdVB7_2(.din(n11708), .dout(n8594));
    jdff dff_A_FNF8GtI49_0(.din(n8600), .dout(n8597));
    jdff dff_A_cda3Ibtk0_0(.din(n8603), .dout(n8600));
    jdff dff_A_ZoqZzlTJ5_0(.din(n8606), .dout(n8603));
    jdff dff_A_PY053j2E3_0(.din(n8609), .dout(n8606));
    jdff dff_A_NWjxawI12_0(.din(n2840), .dout(n8609));
    jdff dff_B_aw7lozyC2_0(.din(n2836), .dout(n8613));
    jdff dff_B_n68jINf37_0(.din(n8613), .dout(n8616));
    jdff dff_A_CsKIKhNk8_2(.din(n8621), .dout(n8618));
    jdff dff_A_6ClywbqX8_2(.din(n8624), .dout(n8621));
    jdff dff_A_yv9RxOo11_2(.din(n8627), .dout(n8624));
    jdff dff_A_oCgTu8PU1_2(.din(n8630), .dout(n8627));
    jdff dff_A_om3QB3IG7_2(.din(n8633), .dout(n8630));
    jdff dff_A_kIFH2Ysa1_2(.din(n8636), .dout(n8633));
    jdff dff_A_b1lHgAcI0_2(.din(n8639), .dout(n8636));
    jdff dff_A_OKjBty4r9_2(.din(n8642), .dout(n8639));
    jdff dff_A_RsAMSWpq3_2(.din(n10829), .dout(n8642));
    jdff dff_B_mBIfwTu57_0(.din(n3375), .dout(n8646));
    jdff dff_B_HxCQNKHB7_0(.din(n8646), .dout(n8649));
    jdff dff_B_Qes4Prln1_0(.din(n8649), .dout(n8652));
    jdff dff_B_9gG2pNCA3_0(.din(n8652), .dout(n8655));
    jdff dff_B_jlxAK9nM9_0(.din(n8655), .dout(n8658));
    jdff dff_B_9cMgXHwX2_0(.din(n3360), .dout(n8661));
    jdff dff_B_t2YV5ulg4_0(.din(n8661), .dout(n8664));
    jdff dff_B_RF4hpguR9_1(.din(n3303), .dout(n8667));
    jdff dff_B_A3jLiNuo4_1(.din(n8667), .dout(n8670));
    jdff dff_B_BNt8wNsu8_1(.din(n8670), .dout(n8673));
    jdff dff_B_tyQKaLlA7_0(.din(n3348), .dout(n8676));
    jdff dff_B_KdZ70WhS7_0(.din(n8676), .dout(n8679));
    jdff dff_B_7ESZrZng0_0(.din(n3340), .dout(n8682));
    jdff dff_A_8psWY8rS6_1(.din(n8687), .dout(n8684));
    jdff dff_A_YyiYAuhi0_1(.din(n77), .dout(n8687));
    jdff dff_A_XMNBXna95_2(.din(n8693), .dout(n8690));
    jdff dff_A_6uaoxXlx0_2(.din(n8696), .dout(n8693));
    jdff dff_A_DSLseczh2_2(.din(n8699), .dout(n8696));
    jdff dff_A_FadPCto76_2(.din(n77), .dout(n8699));
    jdff dff_A_4iOF6mXk2_2(.din(n8705), .dout(n8702));
    jdff dff_A_Sd7ZNSfY2_2(.din(n8708), .dout(n8705));
    jdff dff_A_CVp4pTp89_2(.din(n8711), .dout(n8708));
    jdff dff_A_8fctjVtq2_2(.din(n77), .dout(n8711));
    jdff dff_B_6MfxNJ1F1_0(.din(n3321), .dout(n8715));
    jdff dff_B_Q4nvGl6c1_0(.din(n3317), .dout(n8718));
    jdff dff_A_K5y6vMox0_1(.din(n286), .dout(n8720));
    jdff dff_B_3f5k93LL3_0(.din(n282), .dout(n8724));
    jdff dff_A_iXiu8ig33_0(.din(n8729), .dout(n8726));
    jdff dff_A_40PAzvkt0_0(.din(G232), .dout(n8729));
    jdff dff_A_rNztm4fG1_1(.din(n8735), .dout(n8732));
    jdff dff_A_De6k9eKv4_1(.din(n8738), .dout(n8735));
    jdff dff_A_5mpRZrMx0_1(.din(G232), .dout(n8738));
    jdff dff_A_PfoVU7vB4_2(.din(n8744), .dout(n8741));
    jdff dff_A_rGcJMBIj6_2(.din(G232), .dout(n8744));
    jdff dff_A_WPNxCxhU7_0(.din(n8750), .dout(n8747));
    jdff dff_A_wBv5RdHQ9_0(.din(G226), .dout(n8750));
    jdff dff_A_OHByhVgl2_1(.din(n8756), .dout(n8753));
    jdff dff_A_8DaOgCE19_1(.din(G226), .dout(n8756));
    jdff dff_A_Sn8UzVX90_2(.din(n8762), .dout(n8759));
    jdff dff_A_AEw2G3VR6_2(.din(n8765), .dout(n8762));
    jdff dff_A_cOKP08oN6_2(.din(G226), .dout(n8765));
    jdff dff_A_e6d3Dqpr7_1(.din(n8771), .dout(n8768));
    jdff dff_A_fJHbRvmw7_1(.din(n8774), .dout(n8771));
    jdff dff_A_gH7AkekS8_1(.din(n8777), .dout(n8774));
    jdff dff_A_eiDE24Oq2_1(.din(n2854), .dout(n8777));
    jdff dff_B_LDgdsH4j0_0(.din(n3288), .dout(n8781));
    jdff dff_B_mJyPI1ZB7_0(.din(n8781), .dout(n8784));
    jdff dff_B_K0aRBr5x9_1(.din(n3228), .dout(n8787));
    jdff dff_B_TGNX02BM7_1(.din(n8787), .dout(n8790));
    jdff dff_B_XsJZ1J8F9_1(.din(n8790), .dout(n8793));
    jdff dff_B_gNEDBGez0_1(.din(n8793), .dout(n8796));
    jdff dff_B_USA1XYU61_0(.din(n3272), .dout(n8799));
    jdff dff_A_JHKb9dFG7_1(.din(n8804), .dout(n8801));
    jdff dff_A_aPMWqlyr2_1(.din(n8807), .dout(n8804));
    jdff dff_A_AszVSaBX6_1(.din(n8810), .dout(n8807));
    jdff dff_A_qFW8mvb81_1(.din(n8813), .dout(n8810));
    jdff dff_A_tsGL62uo6_1(.din(n11468), .dout(n8813));
    jdff dff_A_yoJMUpJN0_2(.din(n8819), .dout(n8816));
    jdff dff_A_x9FcaIIF3_2(.din(n11468), .dout(n8819));
    jdff dff_B_ITkbkyJf1_1(.din(n3244), .dout(n8823));
    jdff dff_B_uJOhXaQ34_1(.din(n3232), .dout(n8826));
    jdff dff_A_XgHMaMKJ0_1(.din(n11513), .dout(n8828));
    jdff dff_B_PERCOOkK4_1(.din(n3172), .dout(n8832));
    jdff dff_B_h4qqhYoZ3_1(.din(n3190), .dout(n8835));
    jdff dff_B_O3Odp1da0_0(.din(n3206), .dout(n8838));
    jdff dff_B_v9iNmF707_0(.din(n8838), .dout(n8841));
    jdff dff_B_RwoL5VWu8_1(.din(n3194), .dout(n8844));
    jdff dff_A_sDiaw4jP0_1(.din(n8852), .dout(n8846));
    jdff dff_A_xY4JYrGU6_0(.din(n8859), .dout(n8849));
    jdff dff_A_fhwY2GGF7_1(.din(n8859), .dout(n8852));
    jdff dff_B_lOVN20O51_3(.din(G150), .dout(n8856));
    jdff dff_B_rVxBzmCT4_3(.din(n8856), .dout(n8859));
    jdff dff_A_CxId2X4p1_0(.din(n8864), .dout(n8861));
    jdff dff_A_YeNUUbk43_0(.din(n8867), .dout(n8864));
    jdff dff_A_Yq1g9EbF9_0(.din(G50), .dout(n8867));
    jdff dff_A_QovUWjK44_1(.din(n8873), .dout(n8870));
    jdff dff_A_PCgw152I9_1(.din(n8876), .dout(n8873));
    jdff dff_A_W5vhrWtU2_1(.din(G50), .dout(n8876));
    jdff dff_A_xR7b1os08_1(.din(n3186), .dout(n8879));
    jdff dff_A_PcNxiZVX6_0(.din(n10364), .dout(n8882));
    jdff dff_A_IIsPcozW7_1(.din(n10364), .dout(n8885));
    jdff dff_A_O0UPS0rg6_1(.din(n10412), .dout(n8888));
    jdff dff_A_u3LkBAgE3_2(.din(n10412), .dout(n8891));
    jdff dff_B_UF5t5H872_1(.din(n3153), .dout(n8895));
    jdff dff_B_8Vywqy5C4_1(.din(n8895), .dout(n8898));
    jdff dff_A_C1qcDK9h2_1(.din(n8903), .dout(n8900));
    jdff dff_A_vSeCGvWH5_1(.din(n8906), .dout(n8903));
    jdff dff_A_xOXKEPir9_1(.din(G68), .dout(n8906));
    jdff dff_A_A5yn995E5_2(.din(n8912), .dout(n8909));
    jdff dff_A_5zADzc499_2(.din(n8915), .dout(n8912));
    jdff dff_A_8LkxneID7_2(.din(n8918), .dout(n8915));
    jdff dff_A_V27RGjLX5_2(.din(G68), .dout(n8918));
    jdff dff_A_jZ8bFWoo9_1(.din(n2914), .dout(n8921));
    jdff dff_A_YnKQKoVh5_1(.din(n11447), .dout(n8924));
    jdff dff_A_MzxxoxCA9_1(.din(n8930), .dout(n8927));
    jdff dff_A_DVdKI9wv2_1(.din(n8933), .dout(n8930));
    jdff dff_A_yuAZQRgU4_1(.din(n9803), .dout(n8933));
    jdff dff_A_ef7BMETH9_0(.din(n8939), .dout(n8936));
    jdff dff_A_tuXdhDwY1_0(.din(n10214), .dout(n8939));
    jdff dff_A_Ipm7vSBl0_2(.din(n8945), .dout(n8942));
    jdff dff_A_bAIyhmRv0_2(.din(n10214), .dout(n8945));
    jdff dff_A_JvW1s6wj8_0(.din(n8951), .dout(n8948));
    jdff dff_A_U5NGfB3C5_0(.din(n9932), .dout(n8951));
    jdff dff_A_4jPOWda36_2(.din(n8957), .dout(n8954));
    jdff dff_A_VXiDgnTl0_2(.din(n8960), .dout(n8957));
    jdff dff_A_mQ5PH6K54_2(.din(n9932), .dout(n8960));
    jdff dff_A_BZKHOI4D0_1(.din(n8966), .dout(n8963));
    jdff dff_A_w0RmUAOp6_1(.din(n8969), .dout(n8966));
    jdff dff_A_qcIAzvu09_1(.din(n8972), .dout(n8969));
    jdff dff_A_uhmDajlO9_1(.din(n11768), .dout(n8972));
    jdff dff_A_dHVanQTw5_2(.din(n8978), .dout(n8975));
    jdff dff_A_Nyew7vER2_2(.din(n8981), .dout(n8978));
    jdff dff_A_wqkhJfN54_2(.din(n8984), .dout(n8981));
    jdff dff_A_Zi7TV5ts4_2(.din(n8987), .dout(n8984));
    jdff dff_A_hwu55APx7_2(.din(n8990), .dout(n8987));
    jdff dff_A_K1yCmZ129_2(.din(n8993), .dout(n8990));
    jdff dff_A_FmQ1WqRS3_2(.din(n8996), .dout(n8993));
    jdff dff_A_nkb3mWIg6_2(.din(n8999), .dout(n8996));
    jdff dff_A_XOHknlG88_2(.din(n11768), .dout(n8999));
    jdff dff_A_Lq4xPcLF3_1(.din(n9005), .dout(n9002));
    jdff dff_A_GsUCtSeh1_1(.din(n2082), .dout(n9005));
    jdff dff_A_rV0vbByL7_0(.din(n2078), .dout(n9008));
    jdff dff_A_mUoU2YLO5_1(.din(n9014), .dout(n9011));
    jdff dff_A_wN72twRj6_1(.din(n2078), .dout(n9014));
    jdff dff_B_STIrPms96_0(.din(n2074), .dout(n9018));
    jdff dff_A_psZ4pvPn6_0(.din(n9023), .dout(n9020));
    jdff dff_A_mGCpcx5X1_0(.din(n2071), .dout(n9023));
    jdff dff_A_xy45DvJ30_1(.din(n9029), .dout(n9026));
    jdff dff_A_D6gbvKTe2_1(.din(n9032), .dout(n9029));
    jdff dff_A_dcoKiQBF6_1(.din(n9035), .dout(n9032));
    jdff dff_A_BlOSIGtz5_1(.din(n9038), .dout(n9035));
    jdff dff_A_UDYrwmQr2_1(.din(n9408), .dout(n9038));
    jdff dff_B_vcISusnL7_0(.din(n2035), .dout(n9042));
    jdff dff_B_rBoAC2sS8_0(.din(n9042), .dout(n9045));
    jdff dff_A_WW3mbcMB1_1(.din(n9050), .dout(n9047));
    jdff dff_A_fFhQYuH08_1(.din(n1882), .dout(n9050));
    jdff dff_A_I6SmfvYh6_1(.din(n1117), .dout(n9053));
    jdff dff_A_I6R4qOpr9_1(.din(n9059), .dout(n9056));
    jdff dff_A_CwkCNF3L1_1(.din(n11000), .dout(n9059));
    jdff dff_A_IvJ5Yk489_0(.din(n866), .dout(n9062));
    jdff dff_B_OrLSHVmi8_1(.din(n1793), .dout(n9066));
    jdff dff_B_azq4YLDP6_1(.din(n1842), .dout(n9069));
    jdff dff_B_acPEU2UT6_1(.din(n1028), .dout(n9072));
    jdff dff_A_8l4yuvmS0_1(.din(n1024), .dout(n9074));
    jdff dff_A_BhmWJ5Xk8_2(.din(n1024), .dout(n9077));
    jdff dff_B_L6k4xnL21_1(.din(n988), .dout(n9081));
    jdff dff_B_RxrF3lmL5_1(.din(n9081), .dout(n9084));
    jdff dff_A_CJmQAE0W4_2(.din(n12161), .dout(n9086));
    jdff dff_A_uBod4A164_1(.din(n330), .dout(n9089));
    jdff dff_A_6qfkpFnA6_2(.din(n330), .dout(n9092));
    jdff dff_A_VOUHRpC53_0(.din(n9098), .dout(n9095));
    jdff dff_A_iYvogae46_0(.din(n1068), .dout(n9098));
    jdff dff_A_gaaqrNnu9_0(.din(n11363), .dout(n9101));
    jdff dff_A_myzdZv9H0_1(.din(n9107), .dout(n9104));
    jdff dff_A_CZyKlEfI8_1(.din(n11363), .dout(n9107));
    jdff dff_B_vGb3QaKr3_0(.din(n1097), .dout(n9111));
    jdff dff_A_UH2mw9IG9_1(.din(n9116), .dout(n9113));
    jdff dff_A_v6Kexx641_1(.din(n1016), .dout(n9116));
    jdff dff_B_aDt2lZxg4_1(.din(n1074), .dout(n9120));
    jdff dff_A_lGjIW0tb1_2(.din(n9125), .dout(n9122));
    jdff dff_A_ZVkHsFxW5_2(.din(n74), .dout(n9125));
    jdff dff_A_Wn6G64x50_1(.din(n9131), .dout(n9128));
    jdff dff_A_P5CCnnsY7_1(.din(n9134), .dout(n9131));
    jdff dff_A_vIN32VZI0_1(.din(n9137), .dout(n9134));
    jdff dff_A_UjcH846S9_1(.din(n74), .dout(n9137));
    jdff dff_A_ugurzdDE3_2(.din(n9143), .dout(n9140));
    jdff dff_A_AOrGp42Y8_2(.din(n74), .dout(n9143));
    jdff dff_A_4IRxXou16_0(.din(n9149), .dout(n9146));
    jdff dff_A_4u1g0nRA4_0(.din(n992), .dout(n9149));
    jdff dff_A_c0kaHqI69_2(.din(n9155), .dout(n9152));
    jdff dff_A_sABhtlWN3_2(.din(n992), .dout(n9155));
    jdff dff_A_ugfSWE8Z0_1(.din(G33), .dout(n9158));
    jdff dff_A_S3P8vT1S3_0(.din(n9164), .dout(n9161));
    jdff dff_A_hyYF8zgZ9_0(.din(n9167), .dout(n9164));
    jdff dff_A_PoKWS1oL5_0(.din(n985), .dout(n9167));
    jdff dff_A_4f98VY5J0_0(.din(n981), .dout(n9170));
    jdff dff_A_r52exDBL5_0(.din(n974), .dout(n9173));
    jdff dff_A_UL17uMyz6_1(.din(n9179), .dout(n9176));
    jdff dff_A_lCjPuVzC0_1(.din(n970), .dout(n9179));
    jdff dff_A_zQqKriJB3_0(.din(n9185), .dout(n9182));
    jdff dff_A_KOZBvQqa7_0(.din(n9188), .dout(n9185));
    jdff dff_A_2fVsdO4y2_0(.din(n151), .dout(n9188));
    jdff dff_A_DBtIjgyf7_0(.din(G244), .dout(n9191));
    jdff dff_A_T04A5Jm83_0(.din(n9197), .dout(n9194));
    jdff dff_A_09glOBoH0_0(.din(n928), .dout(n9197));
    jdff dff_A_EW6FVQyj1_0(.din(n9203), .dout(n9200));
    jdff dff_A_pI5UWDYu8_0(.din(n10934), .dout(n9203));
    jdff dff_A_K3q8J32N3_1(.din(n9209), .dout(n9206));
    jdff dff_A_rkfMiR059_1(.din(n10934), .dout(n9209));
    jdff dff_A_Gm4CyLtF8_1(.din(n1827), .dout(n9212));
    jdff dff_A_V6jSsjcw7_1(.din(n10457), .dout(n9215));
    jdff dff_B_zLrZuBmg2_0(.din(n820), .dout(n9219));
    jdff dff_B_0yChTZMT8_1(.din(n793), .dout(n9222));
    jdff dff_A_WruRIkvC8_0(.din(n11525), .dout(n9224));
    jdff dff_A_Maqp9vwT3_1(.din(n9230), .dout(n9227));
    jdff dff_A_7UT1Tdcn2_1(.din(n786), .dout(n9230));
    jdff dff_A_IAiOz3ZI6_2(.din(n9236), .dout(n9233));
    jdff dff_A_FZAOHU4A3_2(.din(n786), .dout(n9236));
    jdff dff_A_HKxjezPj9_1(.din(n870), .dout(n9239));
    jdff dff_A_0C1uqOXc6_0(.din(n431), .dout(n9242));
    jdff dff_A_ojfbe8eC4_2(.din(n9248), .dout(n9245));
    jdff dff_A_aIBsKakw8_2(.din(n431), .dout(n9248));
    jdff dff_A_Q4Evzbr60_0(.din(n9254), .dout(n9251));
    jdff dff_A_ZNRnTKv70_0(.din(n817), .dout(n9254));
    jdff dff_A_s9hBFqu00_0(.din(n9260), .dout(n9257));
    jdff dff_A_HmUdrO5U0_0(.din(n790), .dout(n9260));
    jdff dff_A_cu6nqP592_1(.din(n9266), .dout(n9263));
    jdff dff_A_jIEF3LPd4_1(.din(n790), .dout(n9266));
    jdff dff_A_LFqTsjbc6_0(.din(G33), .dout(n9269));
    jdff dff_A_YBop4ogN4_1(.din(G33), .dout(n9272));
    jdff dff_A_d4Ac9V5o7_1(.din(n783), .dout(n9275));
    jdff dff_A_Mk9d0q7l7_1(.din(n12158), .dout(n9278));
    jdff dff_A_ptBuZUVv8_2(.din(n9284), .dout(n9281));
    jdff dff_A_bzBoME3G6_2(.din(n12158), .dout(n9284));
    jdff dff_A_Q2RwdHnB6_1(.din(n771), .dout(n9287));
    jdff dff_A_y6QJ2NYk0_1(.din(n767), .dout(n9290));
    jdff dff_A_LKGd0RP57_0(.din(n748), .dout(n9293));
    jdff dff_A_5pvZ8Iej6_1(.din(n744), .dout(n9296));
    jdff dff_A_jJRwyNRU9_1(.din(n732), .dout(n9299));
    jdff dff_A_VMpsqkN26_0(.din(n9305), .dout(n9302));
    jdff dff_A_MgaHJqQP3_0(.din(n9308), .dout(n9305));
    jdff dff_A_WGcIau8i4_0(.din(G238), .dout(n9308));
    jdff dff_A_kslexxj42_1(.din(n9314), .dout(n9311));
    jdff dff_A_vm0PmMfd2_1(.din(G238), .dout(n9314));
    jdff dff_A_lUeRqMzZ6_0(.din(n718), .dout(n9317));
    jdff dff_A_Lyne1nuA5_1(.din(n9323), .dout(n9320));
    jdff dff_A_xBgHXuCO4_1(.din(G244), .dout(n9323));
    jdff dff_A_Yh9u04z25_2(.din(n9329), .dout(n9326));
    jdff dff_A_a4qbyPcr0_2(.din(G244), .dout(n9329));
    jdff dff_A_ONNWueaN8_1(.din(n10262), .dout(n9332));
    jdff dff_A_JHn4h5fV4_2(.din(n9338), .dout(n9335));
    jdff dff_A_JoHpLu1U0_2(.din(n10262), .dout(n9338));
    jdff dff_A_xbHy7meL8_0(.din(n9344), .dout(n9341));
    jdff dff_A_SqJOrxYE3_0(.din(n1774), .dout(n9344));
    jdff dff_A_h97w8Uuz8_0(.din(n9350), .dout(n9347));
    jdff dff_A_q04uKjDl0_0(.din(n12038), .dout(n9350));
    jdff dff_A_XbByAM9Z5_1(.din(n9356), .dout(n9353));
    jdff dff_A_VK0Jemwn8_1(.din(n12038), .dout(n9356));
    jdff dff_A_lk2PBJq41_0(.din(n3086), .dout(n9359));
    jdff dff_B_Fsh1G4pF3_0(.din(n3075), .dout(n9363));
    jdff dff_A_4EkeUj953_2(.din(n1997), .dout(n9365));
    jdff dff_B_7izUGPf87_0(.din(n1993), .dout(n9369));
    jdff dff_B_7kdH1aLg2_0(.din(n9369), .dout(n9372));
    jdff dff_B_YHsPo9ub3_0(.din(n9372), .dout(n9375));
    jdff dff_A_pyvMT0dW7_0(.din(n9380), .dout(n9377));
    jdff dff_A_ubAFFJDR1_0(.din(n9383), .dout(n9380));
    jdff dff_A_eNjzWxfS2_1(.din(n9386), .dout(n9383));
    jdff dff_A_0YNUmbHB5_1(.din(n9408), .dout(n9386));
    jdff dff_A_BeM6e52w4_2(.din(n9392), .dout(n9389));
    jdff dff_A_tA6eYaIu4_2(.din(n9408), .dout(n9392));
    jdff dff_B_FCYgFZDb8_3(.din(n1965), .dout(n9396));
    jdff dff_B_Dgf2wMUK4_3(.din(n9396), .dout(n9399));
    jdff dff_B_0mSZYAmZ8_3(.din(n9399), .dout(n9402));
    jdff dff_B_leZnMZJz3_3(.din(n9402), .dout(n9405));
    jdff dff_B_fj0fuCCv9_3(.din(n9405), .dout(n9408));
    jdff dff_A_C6mqboJQ1_1(.din(n9413), .dout(n9410));
    jdff dff_A_yg7TGh7s4_1(.din(n9416), .dout(n9413));
    jdff dff_A_dMFM4oPT9_1(.din(n9419), .dout(n9416));
    jdff dff_A_0v9d9oYZ3_1(.din(n9422), .dout(n9419));
    jdff dff_A_Nbk5Aqs47_1(.din(n9425), .dout(n9422));
    jdff dff_A_fRorsgP65_1(.din(n1952), .dout(n9425));
    jdff dff_A_b8cO9g9e4_0(.din(n1962), .dout(n9428));
    jdff dff_A_Gva2bMP27_1(.din(n9434), .dout(n9431));
    jdff dff_A_MeHRTeA34_1(.din(n714), .dout(n9434));
    jdff dff_A_tCXveOjQ6_2(.din(n714), .dout(n9437));
    jdff dff_A_pbCCveUn4_1(.din(n698), .dout(n9440));
    jdff dff_A_UM007gqd4_1(.din(n9446), .dout(n9443));
    jdff dff_A_1H4g7aOH3_1(.din(n694), .dout(n9446));
    jdff dff_A_sSWuGHby9_1(.din(n9452), .dout(n9449));
    jdff dff_A_KXepKQry7_1(.din(n9455), .dout(n9452));
    jdff dff_A_Bc6Smvon8_1(.din(n682), .dout(n9455));
    jdff dff_B_H5DWbEEY9_1(.din(n652), .dout(n9459));
    jdff dff_A_ehyGtSRL7_1(.din(n663), .dout(n9461));
    jdff dff_B_l6ynPKtQ1_1(.din(n655), .dout(n9465));
    jdff dff_B_vjIuho306_1(.din(n9465), .dout(n9468));
    jdff dff_A_m0U3yfr82_0(.din(n646), .dout(n9470));
    jdff dff_A_t9qhoLV72_2(.din(n646), .dout(n9473));
    jdff dff_B_3956jpsI0_0(.din(n642), .dout(n9477));
    jdff dff_B_v4umk7t39_1(.din(n618), .dout(n9480));
    jdff dff_A_jTypQ46G6_1(.din(n622), .dout(n9482));
    jdff dff_A_y5iOTmpa2_0(.din(n330), .dout(n9485));
    jdff dff_B_b6QY8yMK0_0(.din(n614), .dout(n9489));
    jdff dff_A_wpDTwxvd2_0(.din(n104), .dout(n9491));
    jdff dff_A_hlo8UFjr6_1(.din(n602), .dout(n9494));
    jdff dff_A_E0X6eWJ73_1(.din(n9500), .dout(n9497));
    jdff dff_A_BlTCyyYc9_1(.din(n598), .dout(n9500));
    jdff dff_A_bViPQEmR9_0(.din(n579), .dout(n9503));
    jdff dff_A_JqIje15q7_2(.din(n115), .dout(n9506));
    jdff dff_A_4Z7QsvPG7_1(.din(n115), .dout(n9509));
    jdff dff_A_9Zcfe4AD1_2(.din(n115), .dout(n9512));
    jdff dff_A_XtgaX3F38_0(.din(n9518), .dout(n9515));
    jdff dff_A_UifMbqcT0_0(.din(G250), .dout(n9518));
    jdff dff_A_eQ84Agja2_1(.din(n560), .dout(n9521));
    jdff dff_A_GS59ELfG3_1(.din(n9527), .dout(n9524));
    jdff dff_A_smOwfoRH9_1(.din(n556), .dout(n9527));
    jdff dff_A_dZlq84rC4_0(.din(n9533), .dout(n9530));
    jdff dff_A_ezplO8FG1_0(.din(n431), .dout(n9533));
    jdff dff_A_9GkQ8nxk7_1(.din(n9539), .dout(n9536));
    jdff dff_A_UT5E5WLW6_1(.din(n431), .dout(n9539));
    jdff dff_A_zwpxlafl6_0(.din(n9545), .dout(n9542));
    jdff dff_A_mCUAmSWn7_0(.din(n9548), .dout(n9545));
    jdff dff_A_kq9R0Hx92_0(.din(n9570), .dout(n9548));
    jdff dff_A_d9JyWCYQ8_2(.din(n9570), .dout(n9551));
    jdff dff_B_1o0b1wRq7_3(.din(n548), .dout(n9555));
    jdff dff_B_2fIvKTzI6_3(.din(n9555), .dout(n9558));
    jdff dff_B_n66BveGg3_3(.din(n9558), .dout(n9561));
    jdff dff_B_dQmmLHRO0_3(.din(n9561), .dout(n9564));
    jdff dff_B_kMTbtHbg6_3(.din(n9564), .dout(n9567));
    jdff dff_B_ffUfftvl6_3(.din(n9567), .dout(n9570));
    jdff dff_A_2TRl5kqn1_0(.din(n9575), .dout(n9572));
    jdff dff_A_f3ju7Xvn3_0(.din(n1989), .dout(n9575));
    jdff dff_B_iXyxHpsb3_2(.din(n4259), .dout(n9579));
    jdff dff_B_mXIarFpT2_2(.din(n9579), .dout(n9582));
    jdff dff_B_CnME2FJ40_2(.din(n9582), .dout(n9585));
    jdff dff_B_W7UKalJt1_2(.din(n9585), .dout(n9588));
    jdff dff_B_7dexFQRr4_1(.din(n2142), .dout(n9591));
    jdff dff_B_3KsAx5iO0_0(.din(n2452), .dout(n9594));
    jdff dff_B_hoiOK8je7_0(.din(n2448), .dout(n9597));
    jdff dff_B_eIU6FKJH2_0(.din(n9597), .dout(n9600));
    jdff dff_B_H2ok2CHD2_0(.din(n2437), .dout(n9603));
    jdff dff_B_2uiw1TE68_0(.din(n9603), .dout(n9606));
    jdff dff_A_Icil9oyk6_0(.din(n2429), .dout(n9608));
    jdff dff_A_HV5MqwNv4_0(.din(n9614), .dout(n9611));
    jdff dff_A_wCY4BIU75_0(.din(n9617), .dout(n9614));
    jdff dff_A_FJXwIsoD3_0(.din(n9620), .dout(n9617));
    jdff dff_A_B099aipu7_0(.din(n9623), .dout(n9620));
    jdff dff_A_I9OoPHr58_0(.din(n9626), .dout(n9623));
    jdff dff_A_3RdTVT158_0(.din(n10724), .dout(n9626));
    jdff dff_A_0mHxmi5c9_1(.din(n9632), .dout(n9629));
    jdff dff_A_prntjCou7_1(.din(n9635), .dout(n9632));
    jdff dff_A_YJ7N1I1O6_1(.din(n9638), .dout(n9635));
    jdff dff_A_u93sXQNP5_1(.din(n9641), .dout(n9638));
    jdff dff_A_zIyt1ZDW7_1(.din(n10724), .dout(n9641));
    jdff dff_A_2tQIXM091_0(.din(n112), .dout(n9644));
    jdff dff_A_BXp19r1I9_2(.din(n9650), .dout(n9647));
    jdff dff_A_Gtl4BAO57_2(.din(n9653), .dout(n9650));
    jdff dff_A_NKXy33Zt9_2(.din(n104), .dout(n9653));
    jdff dff_A_FSrO6w4K0_0(.din(n9659), .dout(n9656));
    jdff dff_A_bZCkoJDo6_0(.din(n9662), .dout(n9659));
    jdff dff_A_6VTTiOdz4_0(.din(n9665), .dout(n9662));
    jdff dff_A_Y0dcH6Gw9_0(.din(n9668), .dout(n9665));
    jdff dff_A_DcO9EYeb0_0(.din(n9671), .dout(n9668));
    jdff dff_A_ieJJYPRg7_0(.din(G107), .dout(n9671));
    jdff dff_A_VBAT3ybe9_1(.din(n9677), .dout(n9674));
    jdff dff_A_2Ub4ESG99_1(.din(n9680), .dout(n9677));
    jdff dff_A_6ineyHI54_1(.din(G107), .dout(n9680));
    jdff dff_A_zThGJpvx2_2(.din(n9686), .dout(n9683));
    jdff dff_A_diHCYZvR4_2(.din(n9689), .dout(n9686));
    jdff dff_A_AfTxsI4D4_2(.din(G107), .dout(n9689));
    jdff dff_A_ZqrpNP8R5_1(.din(n9695), .dout(n9692));
    jdff dff_A_sukh36C02_1(.din(n101), .dout(n9695));
    jdff dff_A_uCHG4j7O2_2(.din(n9701), .dout(n9698));
    jdff dff_A_hrCraXZX3_2(.din(n9704), .dout(n9701));
    jdff dff_A_D9v8rz468_2(.din(n9707), .dout(n9704));
    jdff dff_A_pK4nazjv8_2(.din(n101), .dout(n9707));
    jdff dff_A_AUfBtQ1c5_0(.din(n9713), .dout(n9710));
    jdff dff_A_PPGohfHm8_0(.din(n9716), .dout(n9713));
    jdff dff_A_Ib35Ox4U7_0(.din(n9719), .dout(n9716));
    jdff dff_A_OFeyg3eT2_0(.din(n98), .dout(n9719));
    jdff dff_A_PRuOSv1q6_2(.din(n98), .dout(n9722));
    jdff dff_A_pJD95jjG5_1(.din(n9728), .dout(n9725));
    jdff dff_A_N68nDtWQ1_1(.din(n98), .dout(n9728));
    jdff dff_A_FMuI1CcA8_0(.din(G87), .dout(n9731));
    jdff dff_B_g2BUHUmX1_1(.din(n2396), .dout(n9735));
    jdff dff_B_AroFzrwl4_1(.din(n9735), .dout(n9738));
    jdff dff_B_EOO2UkWM2_1(.din(n9738), .dout(n9741));
    jdff dff_B_zs0to0HM6_1(.din(n9741), .dout(n9744));
    jdff dff_A_JrF3vsGJ7_2(.din(n9749), .dout(n9746));
    jdff dff_A_Gul787wf1_2(.din(n9752), .dout(n9749));
    jdff dff_A_N1DAoVzM8_2(.din(n9755), .dout(n9752));
    jdff dff_A_Evudwhde2_2(.din(n83), .dout(n9755));
    jdff dff_A_KpwcKUwN2_2(.din(n9761), .dout(n9758));
    jdff dff_A_gusQRcRR1_2(.din(n9764), .dout(n9761));
    jdff dff_A_Pgt8R5mk2_2(.din(n9767), .dout(n9764));
    jdff dff_A_Q82G0qZs0_2(.din(n80), .dout(n9767));
    jdff dff_A_xSsMCRBr7_0(.din(n9773), .dout(n9770));
    jdff dff_A_lW4jTWas2_0(.din(n9776), .dout(n9773));
    jdff dff_A_3elhcIgK5_0(.din(n9779), .dout(n9776));
    jdff dff_A_Qz9JojIl6_0(.din(n9782), .dout(n9779));
    jdff dff_A_FvVptbhJ6_0(.din(n9785), .dout(n9782));
    jdff dff_A_tvZyrkCr1_0(.din(n11561), .dout(n9785));
    jdff dff_A_SprqBrJ81_1(.din(n9791), .dout(n9788));
    jdff dff_A_jlWWod3j4_1(.din(n9794), .dout(n9791));
    jdff dff_A_4ED3xgM51_1(.din(n11561), .dout(n9794));
    jdff dff_A_iVZsRrpd7_0(.din(n9800), .dout(n9797));
    jdff dff_A_2SGy3vXE7_0(.din(n11561), .dout(n9800));
    jdff dff_A_UfpkqPRw4_1(.din(n9806), .dout(n9803));
    jdff dff_A_iCkZqIXJ7_1(.din(n11561), .dout(n9806));
    jdff dff_A_IfmgPiJs5_1(.din(n302), .dout(n9809));
    jdff dff_A_66Lb5xL71_0(.din(G77), .dout(n9812));
    jdff dff_A_kk3grUL39_1(.din(n9818), .dout(n9815));
    jdff dff_A_DLOvlq2Y9_1(.din(n9821), .dout(n9818));
    jdff dff_A_U3yMFeo12_1(.din(n9824), .dout(n9821));
    jdff dff_A_t101vT8I6_1(.din(G77), .dout(n9824));
    jdff dff_A_GYNZU5xm9_0(.din(G68), .dout(n9827));
    jdff dff_A_Z5goGDQd7_2(.din(n9833), .dout(n9830));
    jdff dff_A_ywlBQ1Eu4_2(.din(n9836), .dout(n9833));
    jdff dff_A_atCkOc2f6_2(.din(G68), .dout(n9836));
    jdff dff_A_4T2OBKU75_0(.din(G58), .dout(n9839));
    jdff dff_A_uevzUhaB9_1(.din(n9845), .dout(n9842));
    jdff dff_A_YHrPatvI4_1(.din(n9848), .dout(n9845));
    jdff dff_A_5FfXtKws4_1(.din(G50), .dout(n9848));
    jdff dff_A_Ur4fGXuz7_0(.din(n1136), .dout(n9851));
    jdff dff_A_tvIXBdGs1_1(.din(n9857), .dout(n9854));
    jdff dff_A_Om6iWjaW9_1(.din(n9860), .dout(n9857));
    jdff dff_A_skZTG5Uq4_1(.din(n9863), .dout(n9860));
    jdff dff_A_l5QVFNa52_1(.din(n1136), .dout(n9863));
    jdff dff_A_3kGape6e9_2(.din(n9869), .dout(n9866));
    jdff dff_A_Igq2p78F1_2(.din(n9872), .dout(n9869));
    jdff dff_A_OVOzVEbJ0_2(.din(n1136), .dout(n9872));
    jdff dff_A_HR4uFf1G5_1(.din(n9878), .dout(n9875));
    jdff dff_A_jvgRanVX8_1(.din(n9881), .dout(n9878));
    jdff dff_A_W5TRT1jw1_1(.din(n9884), .dout(n9881));
    jdff dff_A_sHAus9Hg6_1(.din(n2392), .dout(n9884));
    jdff dff_A_6lkBff8a2_1(.din(n9890), .dout(n9887));
    jdff dff_A_r3xTgCrX5_1(.din(n9893), .dout(n9890));
    jdff dff_A_cHLg8j5i1_1(.din(n9896), .dout(n9893));
    jdff dff_A_KxzTbend0_1(.din(n9899), .dout(n9896));
    jdff dff_A_L1OUvBOX5_1(.din(n9902), .dout(n9899));
    jdff dff_A_gLdsm9MT0_1(.din(n9905), .dout(n9902));
    jdff dff_A_vOdaRpIR9_1(.din(n9908), .dout(n9905));
    jdff dff_A_wVzkdJBF7_1(.din(n2384), .dout(n9908));
    jdff dff_A_WB1iM4RD7_1(.din(n9914), .dout(n9911));
    jdff dff_A_HlhaDl444_1(.din(n9917), .dout(n9914));
    jdff dff_A_bUjDrnwq9_1(.din(n9920), .dout(n9917));
    jdff dff_A_Uld5ZWv42_1(.din(n9923), .dout(n9920));
    jdff dff_A_pB17JVLV8_1(.din(n9926), .dout(n9923));
    jdff dff_A_RYyAyxtK4_1(.din(n9929), .dout(n9926));
    jdff dff_A_AieAZqdi9_1(.din(n2384), .dout(n9929));
    jdff dff_A_3UeoD8xh0_1(.din(n9935), .dout(n9932));
    jdff dff_A_mJel1wGl0_1(.din(n9938), .dout(n9935));
    jdff dff_A_iTbNsJcu3_1(.din(n9941), .dout(n9938));
    jdff dff_A_VLgwlKXU5_1(.din(n9944), .dout(n9941));
    jdff dff_A_sQCRFlbg1_1(.din(n2384), .dout(n9944));
    jdff dff_A_pilupIAD1_1(.din(n9950), .dout(n9947));
    jdff dff_A_LlXQbDvJ1_1(.din(n9953), .dout(n9950));
    jdff dff_A_3QuVspq13_1(.din(n9956), .dout(n9953));
    jdff dff_A_qabvBadO0_1(.din(n9959), .dout(n9956));
    jdff dff_A_vBIy6OKn2_1(.din(n9962), .dout(n9959));
    jdff dff_A_Zq0Bc14H4_1(.din(n11360), .dout(n9962));
    jdff dff_A_S1Gy7Grj3_2(.din(n9968), .dout(n9965));
    jdff dff_A_oXYJQoHw7_2(.din(n9971), .dout(n9968));
    jdff dff_A_PVds1BQh4_2(.din(n9974), .dout(n9971));
    jdff dff_A_VG8jbie57_2(.din(n9977), .dout(n9974));
    jdff dff_A_Eibqprn34_2(.din(n9980), .dout(n9977));
    jdff dff_A_abaKJPaS9_2(.din(n9983), .dout(n9980));
    jdff dff_A_huDPOu0W6_2(.din(n9986), .dout(n9983));
    jdff dff_A_n08iQj1A2_2(.din(n11360), .dout(n9986));
    jdff dff_A_NOo5No7a1_1(.din(n9992), .dout(n9989));
    jdff dff_A_ja4D9moc2_1(.din(n9995), .dout(n9992));
    jdff dff_A_4MwNiXOn4_1(.din(n367), .dout(n9995));
    jdff dff_B_epnIwufb4_0(.din(n2369), .dout(n9999));
    jdff dff_B_IPXw9dON6_0(.din(n9999), .dout(n10002));
    jdff dff_B_zQEgkBVr2_1(.din(n2309), .dout(n10005));
    jdff dff_B_SI3vpvEF0_1(.din(n10005), .dout(n10008));
    jdff dff_B_duIrmeBB7_1(.din(n10008), .dout(n10011));
    jdff dff_B_2WX1sdRp1_1(.din(n10011), .dout(n10014));
    jdff dff_B_PGB7mGTc7_0(.din(n2353), .dout(n10017));
    jdff dff_A_wFVyREYN6_0(.din(n10029), .dout(n10019));
    jdff dff_B_15zbGLLk8_3(.din(G317), .dout(n10023));
    jdff dff_B_PFBmPIhI2_3(.din(n10023), .dout(n10026));
    jdff dff_B_aZT4eAIR2_3(.din(n10026), .dout(n10029));
    jdff dff_A_FduAQ6k65_1(.din(n10041), .dout(n10031));
    jdff dff_B_YFWQiIGl2_3(.din(G311), .dout(n10035));
    jdff dff_B_b8tum4Cb1_3(.din(n10035), .dout(n10038));
    jdff dff_B_DleL7hkB5_3(.din(n10038), .dout(n10041));
    jdff dff_B_Qoi6h4hS8_1(.din(G329), .dout(n10044));
    jdff dff_B_MkNT7zZD7_1(.din(n10044), .dout(n10047));
    jdff dff_B_hpPNEX8y4_1(.din(n10047), .dout(n10050));
    jdff dff_B_U5SKTSDO0_1(.din(n10050), .dout(n10053));
    jdff dff_B_s0siIhop1_0(.din(n2325), .dout(n10056));
    jdff dff_B_Xa6NuVoZ9_0(.din(n10056), .dout(n10059));
    jdff dff_A_UAHBuC8a9_0(.din(n10071), .dout(n10061));
    jdff dff_B_ctEQa78R7_2(.din(G326), .dout(n10065));
    jdff dff_B_uWuWFUxP0_2(.din(n10065), .dout(n10068));
    jdff dff_B_3IYLQbVv5_2(.din(n10068), .dout(n10071));
    jdff dff_B_MdHqP3XU9_1(.din(n2313), .dout(n10074));
    jdff dff_A_RvwD4hSX8_0(.din(n10079), .dout(n10076));
    jdff dff_A_HFE3nYvt1_0(.din(n10082), .dout(n10079));
    jdff dff_A_InUxnsUw6_0(.din(n10085), .dout(n10082));
    jdff dff_A_7KXAvexG1_0(.din(G294), .dout(n10085));
    jdff dff_A_nCtp9fmY5_0(.din(n10091), .dout(n10088));
    jdff dff_A_imFC1NFv1_0(.din(n10094), .dout(n10091));
    jdff dff_A_M8PDc24u2_0(.din(G294), .dout(n10094));
    jdff dff_A_dfPF7vOD9_1(.din(n10100), .dout(n10097));
    jdff dff_A_XA49QrCj3_1(.din(n10103), .dout(n10100));
    jdff dff_A_UGB6UDPz6_1(.din(G294), .dout(n10103));
    jdff dff_A_IgwH6UHi3_0(.din(n10116), .dout(n10106));
    jdff dff_B_nT9B3m7w1_3(.din(G322), .dout(n10110));
    jdff dff_B_DuNi19WN8_3(.din(n10110), .dout(n10113));
    jdff dff_B_76RyYuVJ5_3(.din(n10113), .dout(n10116));
    jdff dff_B_XZYEa8my8_0(.din(n2298), .dout(n10119));
    jdff dff_B_ZpGwgD9l5_1(.din(n2255), .dout(n10122));
    jdff dff_B_WwaOHHlo8_1(.din(n10122), .dout(n10125));
    jdff dff_A_Rpv7GXwZ4_1(.din(n10130), .dout(n10127));
    jdff dff_A_gkhyvNus0_1(.din(n10139), .dout(n10130));
    jdff dff_A_99bYBXMd5_2(.din(n10136), .dout(n10133));
    jdff dff_A_YbKn54312_2(.din(n10139), .dout(n10136));
    jdff dff_A_hIy1Evbj3_2(.din(G68), .dout(n10139));
    jdff dff_A_Lvr95I756_0(.din(n10145), .dout(n10142));
    jdff dff_A_myzgEm6o4_0(.din(n10154), .dout(n10145));
    jdff dff_A_bPu9byLN0_1(.din(n10151), .dout(n10148));
    jdff dff_A_IatAuJ4D8_1(.din(n10154), .dout(n10151));
    jdff dff_A_uRXQAEmO4_0(.din(G50), .dout(n10154));
    jdff dff_A_TYmLuvgm0_2(.din(n10160), .dout(n10157));
    jdff dff_A_iPQOF0Vq4_2(.din(n10163), .dout(n10160));
    jdff dff_A_PLpIwZTf2_2(.din(n10166), .dout(n10163));
    jdff dff_A_TfYO4oLX8_2(.din(G50), .dout(n10166));
    jdff dff_A_BaM0tXbx0_1(.din(n2263), .dout(n10169));
    jdff dff_A_rwpDjkM27_0(.din(n10175), .dout(n10172));
    jdff dff_A_u7tOXK7N1_0(.din(n10178), .dout(n10175));
    jdff dff_A_1053Xzse9_0(.din(G107), .dout(n10178));
    jdff dff_A_PSu8SQtN0_1(.din(n10184), .dout(n10181));
    jdff dff_A_mLeTIMsk2_1(.din(n10187), .dout(n10184));
    jdff dff_A_JOflgydm7_1(.din(G107), .dout(n10187));
    jdff dff_A_lbRvUuZh2_0(.din(n10193), .dout(n10190));
    jdff dff_A_GjeJFaG75_0(.din(n10196), .dout(n10193));
    jdff dff_A_JDcLtCSU8_0(.din(G58), .dout(n10196));
    jdff dff_A_jcmTerpl0_2(.din(n10202), .dout(n10199));
    jdff dff_A_ga0eICyE4_2(.din(G58), .dout(n10202));
    jdff dff_A_S2EvNYYq9_2(.din(n10208), .dout(n10205));
    jdff dff_A_a8oYTciW2_2(.din(n10211), .dout(n10208));
    jdff dff_A_oDEU0Bbw2_2(.din(G58), .dout(n10211));
    jdff dff_A_ID44LOwM4_1(.din(G58), .dout(n10214));
    jdff dff_B_cx0kmtJb8_1(.din(n2212), .dout(n10218));
    jdff dff_B_cTi4cvda5_1(.din(n2224), .dout(n10221));
    jdff dff_A_Ud0i2WQE0_0(.din(n10226), .dout(n10223));
    jdff dff_A_LySYsfzo0_0(.din(n10229), .dout(n10226));
    jdff dff_A_uCHVmEAR2_0(.din(G159), .dout(n10229));
    jdff dff_A_RRvMJjBr1_1(.din(n10235), .dout(n10232));
    jdff dff_A_easMpTaD7_1(.din(n10238), .dout(n10235));
    jdff dff_A_wBMgzwlS3_1(.din(n10241), .dout(n10238));
    jdff dff_A_OjRpaYTH3_1(.din(G159), .dout(n10241));
    jdff dff_A_jPZB0Uh39_0(.din(n10247), .dout(n10244));
    jdff dff_A_fgpOljVt1_0(.din(n10250), .dout(n10247));
    jdff dff_A_gTmJHqmw8_0(.din(G159), .dout(n10250));
    jdff dff_A_BoUr2vNR5_1(.din(n10256), .dout(n10253));
    jdff dff_A_7aLUCqxE7_1(.din(n10259), .dout(n10256));
    jdff dff_A_02gL5xdu7_1(.din(G159), .dout(n10259));
    jdff dff_A_FNTuUT801_0(.din(n10265), .dout(n10262));
    jdff dff_A_HTBDeNDf9_0(.din(n10268), .dout(n10265));
    jdff dff_A_VJu7bfcK9_0(.din(n10271), .dout(n10268));
    jdff dff_A_rJbWsbZI0_0(.din(n10274), .dout(n10271));
    jdff dff_A_dhPSkfWg5_0(.din(n10277), .dout(n10274));
    jdff dff_A_hvqDGvPG2_0(.din(n1272), .dout(n10277));
    jdff dff_A_0DNBLfcy6_1(.din(n10283), .dout(n10280));
    jdff dff_A_roSSWwob9_1(.din(n10286), .dout(n10283));
    jdff dff_A_Gn1Ngk807_1(.din(n10289), .dout(n10286));
    jdff dff_A_wRJmGnUW9_1(.din(n10292), .dout(n10289));
    jdff dff_A_nEejx1Yk7_1(.din(n10295), .dout(n10292));
    jdff dff_A_eFTL9DI97_1(.din(n10298), .dout(n10295));
    jdff dff_A_5ZUteJJl5_1(.din(n1272), .dout(n10298));
    jdff dff_A_OVgrBv1T6_1(.din(n10304), .dout(n10301));
    jdff dff_A_CtOhJ50s6_1(.din(n10307), .dout(n10304));
    jdff dff_A_NnTjfPfF4_1(.din(n10310), .dout(n10307));
    jdff dff_A_Z8NYjraw5_1(.din(n10313), .dout(n10310));
    jdff dff_A_VaIGOAew9_1(.din(n10316), .dout(n10313));
    jdff dff_A_cNXzxi6f5_1(.din(n10319), .dout(n10316));
    jdff dff_A_9LhzQicR2_1(.din(n10322), .dout(n10319));
    jdff dff_A_JVEiqZj74_1(.din(G200), .dout(n10322));
    jdff dff_A_juqI9PiX2_2(.din(n10328), .dout(n10325));
    jdff dff_A_dv0y0SBw3_2(.din(n10331), .dout(n10328));
    jdff dff_A_uf482u1O4_2(.din(n10334), .dout(n10331));
    jdff dff_A_ZGUTahiJ3_2(.din(n10337), .dout(n10334));
    jdff dff_A_9gTQKhFJ3_2(.din(n10340), .dout(n10337));
    jdff dff_A_ddD7f9Uq0_2(.din(n10343), .dout(n10340));
    jdff dff_A_RuwTxlmp4_2(.din(G200), .dout(n10343));
    jdff dff_A_7bb0sUTJ1_0(.din(n10349), .dout(n10346));
    jdff dff_A_50Fg1vgp4_0(.din(n10352), .dout(n10349));
    jdff dff_A_RnLehcsx9_0(.din(G77), .dout(n10352));
    jdff dff_A_i9CGDgPG3_2(.din(n10358), .dout(n10355));
    jdff dff_A_MlJChBlm4_2(.din(n10361), .dout(n10358));
    jdff dff_A_6R5e6Vpw8_2(.din(G77), .dout(n10361));
    jdff dff_A_H00ab9SS9_1(.din(n10367), .dout(n10364));
    jdff dff_A_TlHlMIDS6_1(.din(G77), .dout(n10367));
    jdff dff_A_WHNRDtKO3_0(.din(n10373), .dout(n10370));
    jdff dff_A_QzjSqOyr6_0(.din(n10376), .dout(n10373));
    jdff dff_A_iZdiPAK29_0(.din(n10379), .dout(n10376));
    jdff dff_A_i9Y28Gpo5_0(.din(n10382), .dout(n10379));
    jdff dff_A_eH5pr1Dt4_0(.din(n10385), .dout(n10382));
    jdff dff_A_KAokJYo86_0(.din(G33), .dout(n10385));
    jdff dff_A_awdv05eE1_1(.din(G33), .dout(n10388));
    jdff dff_B_HSexzlMl6_0(.din(n2208), .dout(n10392));
    jdff dff_A_f6htjZ0h2_0(.din(n10397), .dout(n10394));
    jdff dff_A_ctYTbV0I7_0(.din(n10400), .dout(n10397));
    jdff dff_A_lb8DHTMQ0_0(.din(G87), .dout(n10400));
    jdff dff_A_2w6f3LV65_1(.din(n10406), .dout(n10403));
    jdff dff_A_8vQCB9x34_1(.din(n10409), .dout(n10406));
    jdff dff_A_sCFfnYDW2_1(.din(G87), .dout(n10409));
    jdff dff_A_1cN0h2PT2_0(.din(n10415), .dout(n10412));
    jdff dff_A_gV5tDO9v0_0(.din(n10418), .dout(n10415));
    jdff dff_A_tP0ttjuI6_0(.din(G87), .dout(n10418));
    jdff dff_A_WuJdh9tN4_0(.din(G200), .dout(n10421));
    jdff dff_A_2SLOiQmU2_2(.din(n10427), .dout(n10424));
    jdff dff_A_JTPDVDkf9_2(.din(n10430), .dout(n10427));
    jdff dff_A_5qPkdKiB1_2(.din(n10433), .dout(n10430));
    jdff dff_A_oMVEQn4J3_2(.din(n10436), .dout(n10433));
    jdff dff_A_naVGPcSL9_2(.din(n10439), .dout(n10436));
    jdff dff_A_jcyD8gAL9_2(.din(n10442), .dout(n10439));
    jdff dff_A_tyIazhTB1_2(.din(n10445), .dout(n10442));
    jdff dff_A_qJJ0psJq6_2(.din(G200), .dout(n10445));
    jdff dff_A_LNnhatrx2_0(.din(n2161), .dout(n10448));
    jdff dff_A_EdOHaFaB2_0(.din(n1724), .dout(n10451));
    jdff dff_A_HegGS2qX4_1(.din(n1724), .dout(n10454));
    jdff dff_A_aJvojiDY3_1(.din(n10460), .dout(n10457));
    jdff dff_A_NSxwuF543_1(.din(n10463), .dout(n10460));
    jdff dff_A_EgUzCAux4_1(.din(n10466), .dout(n10463));
    jdff dff_A_UZiJZi3v3_1(.din(n10469), .dout(n10466));
    jdff dff_A_yLXqfWQo9_1(.din(n10472), .dout(n10469));
    jdff dff_A_qdkzIen67_1(.din(n1724), .dout(n10472));
    jdff dff_A_kt9eReKY6_2(.din(n1724), .dout(n10475));
    jdff dff_A_U5zeaEBP4_0(.din(n10481), .dout(n10478));
    jdff dff_A_mj3y81XF0_0(.din(G190), .dout(n10481));
    jdff dff_A_CirbFGOI2_2(.din(n10487), .dout(n10484));
    jdff dff_A_G1XrAQAe4_2(.din(n10490), .dout(n10487));
    jdff dff_A_kwMSiL5q6_2(.din(n10493), .dout(n10490));
    jdff dff_A_VbPXRntC0_2(.din(n10496), .dout(n10493));
    jdff dff_A_QiMpmbzV4_2(.din(n10499), .dout(n10496));
    jdff dff_A_ggKQXFRs6_2(.din(n10502), .dout(n10499));
    jdff dff_A_wOdYPzuO0_2(.din(n10505), .dout(n10502));
    jdff dff_A_exnGLAXE9_2(.din(G190), .dout(n10505));
    jdff dff_A_Za5J4EeW1_2(.din(G20), .dout(n10508));
    jdff dff_A_uAnlLjrn6_0(.din(n10514), .dout(n10511));
    jdff dff_A_uhWG3V3B0_0(.din(n10517), .dout(n10514));
    jdff dff_A_bKjz2g4f0_0(.din(n10520), .dout(n10517));
    jdff dff_A_P9BlaCSh4_0(.din(G97), .dout(n10520));
    jdff dff_A_SdTEQVUl4_0(.din(n10526), .dout(n10523));
    jdff dff_A_EuxU2Int0_0(.din(n10529), .dout(n10526));
    jdff dff_A_tmBL4v1l1_0(.din(n10532), .dout(n10529));
    jdff dff_A_SZgxCPfN6_0(.din(n10535), .dout(n10532));
    jdff dff_A_2QJJym2f7_0(.din(n10538), .dout(n10535));
    jdff dff_A_AiEo29PQ1_0(.din(n10541), .dout(n10538));
    jdff dff_A_Gqltzonz4_0(.din(n10544), .dout(n10541));
    jdff dff_A_6RJezA6N7_0(.din(n10547), .dout(n10544));
    jdff dff_A_cLTLoYju5_0(.din(n2153), .dout(n10547));
    jdff dff_A_xbB1niDx1_2(.din(n10553), .dout(n10550));
    jdff dff_A_HzjUXLGv1_2(.din(n10556), .dout(n10553));
    jdff dff_A_uX9FTeu49_2(.din(n10559), .dout(n10556));
    jdff dff_A_xm2zcuXS4_2(.din(n10562), .dout(n10559));
    jdff dff_A_z9eqSGSK2_2(.din(n10565), .dout(n10562));
    jdff dff_A_6U9VqsfF3_2(.din(n10568), .dout(n10565));
    jdff dff_A_sH8FbVQ41_2(.din(n10571), .dout(n10568));
    jdff dff_A_ejUtGVit9_2(.din(n10574), .dout(n10571));
    jdff dff_A_hh3UPOJj3_2(.din(n10577), .dout(n10574));
    jdff dff_A_M3oKymkX0_2(.din(n2153), .dout(n10577));
    jdff dff_A_pAH16aaE0_0(.din(n10583), .dout(n10580));
    jdff dff_A_EhRKcNdn1_0(.din(n10586), .dout(n10583));
    jdff dff_A_kbRTm1KI5_0(.din(n10589), .dout(n10586));
    jdff dff_A_3F6v94TU0_0(.din(n10592), .dout(n10589));
    jdff dff_A_jiZw6dXz8_0(.din(n10595), .dout(n10592));
    jdff dff_A_gyGu27sC8_0(.din(n10598), .dout(n10595));
    jdff dff_A_HzuVDqZY0_0(.din(n10601), .dout(n10598));
    jdff dff_A_5ahwCGFI4_0(.din(n10604), .dout(n10601));
    jdff dff_A_pNIealtt9_0(.din(n10607), .dout(n10604));
    jdff dff_A_gUS2zuK58_0(.din(n2150), .dout(n10607));
    jdff dff_A_FigNKfxo7_1(.din(n10613), .dout(n10610));
    jdff dff_A_260bEBTC6_1(.din(n10616), .dout(n10613));
    jdff dff_A_VEn8q4z92_1(.din(n10619), .dout(n10616));
    jdff dff_A_msprWaCP2_1(.din(n10622), .dout(n10619));
    jdff dff_A_zdJ6DOrn3_1(.din(n10625), .dout(n10622));
    jdff dff_A_2mkDxWwO8_1(.din(n10628), .dout(n10625));
    jdff dff_A_XVHiTYCN8_1(.din(n10631), .dout(n10628));
    jdff dff_A_Gr4gVzGG9_1(.din(n10634), .dout(n10631));
    jdff dff_A_pRUa8Ttq1_1(.din(n2150), .dout(n10634));
    jdff dff_A_zJ3ZWgMV1_0(.din(n10640), .dout(n10637));
    jdff dff_A_4yptJBWd6_0(.din(n10643), .dout(n10640));
    jdff dff_A_yjrrCu7o5_0(.din(n10646), .dout(n10643));
    jdff dff_A_ibZVVIeY2_0(.din(n10649), .dout(n10646));
    jdff dff_A_DuypDAPN2_0(.din(n10652), .dout(n10649));
    jdff dff_A_2kPYGMWC2_0(.din(n10655), .dout(n10652));
    jdff dff_A_35poXltV8_0(.din(n10658), .dout(n10655));
    jdff dff_A_TwCJsRjF2_0(.din(n10661), .dout(n10658));
    jdff dff_A_SgxLCfYC5_0(.din(n10664), .dout(n10661));
    jdff dff_A_tFbVVaAs8_0(.din(n10667), .dout(n10664));
    jdff dff_A_oUZrYATW0_0(.din(n10670), .dout(n10667));
    jdff dff_A_QFvgbUU20_0(.din(n10673), .dout(n10670));
    jdff dff_A_8kOfjuPP0_0(.din(n2146), .dout(n10673));
    jdff dff_A_k7wsKiL36_2(.din(n10679), .dout(n10676));
    jdff dff_A_xf7JuvVR3_2(.din(n10682), .dout(n10679));
    jdff dff_A_qemMsgKK9_2(.din(n10685), .dout(n10682));
    jdff dff_A_HYhoACAY5_2(.din(n10688), .dout(n10685));
    jdff dff_A_w3mQjxe81_2(.din(n10691), .dout(n10688));
    jdff dff_A_zCGulpcr7_2(.din(n10694), .dout(n10691));
    jdff dff_A_0NDY6e3v0_2(.din(n10697), .dout(n10694));
    jdff dff_A_W0WBHR8e2_2(.din(n10700), .dout(n10697));
    jdff dff_A_K0Pad6Ns8_2(.din(n10703), .dout(n10700));
    jdff dff_A_4kzqbnWJ8_2(.din(n10706), .dout(n10703));
    jdff dff_A_yjipZPyy5_2(.din(n10709), .dout(n10706));
    jdff dff_A_V5rlJOz46_2(.din(n2146), .dout(n10709));
    jdff dff_A_I9dstlAO9_0(.din(n10715), .dout(n10712));
    jdff dff_A_JEtBTcVc0_0(.din(n10718), .dout(n10715));
    jdff dff_A_xWn1uct69_0(.din(n10721), .dout(n10718));
    jdff dff_A_uk6JKueg4_0(.din(n374), .dout(n10721));
    jdff dff_A_cj41HD791_0(.din(n10727), .dout(n10724));
    jdff dff_A_RNoxb2dK4_0(.din(n374), .dout(n10727));
    jdff dff_B_w3v2F4oM6_1(.din(n2134), .dout(n10731));
    jdff dff_B_HIhbgpsC2_1(.din(n10731), .dout(n10734));
    jdff dff_B_mV0nW1Tm9_1(.din(n10734), .dout(n10737));
    jdff dff_B_60ChBBxI3_1(.din(n10737), .dout(n10740));
    jdff dff_B_FKThuiyb9_1(.din(n10740), .dout(n10743));
    jdff dff_B_Od5Gk1gw0_1(.din(n10743), .dout(n10746));
    jdff dff_B_B3u4cSBY8_1(.din(n10746), .dout(n10749));
    jdff dff_B_q8k9MOuf7_1(.din(n10749), .dout(n10752));
    jdff dff_B_KvJ7e3XT4_0(.din(n1981), .dout(n10755));
    jdff dff_B_0Vssa9tt8_0(.din(n10755), .dout(n10758));
    jdff dff_B_7xDTL5ru8_0(.din(n10758), .dout(n10761));
    jdff dff_B_jvbrpiFg4_0(.din(n10761), .dout(n10764));
    jdff dff_A_m7ctGy0p4_0(.din(n10769), .dout(n10766));
    jdff dff_A_QGRxRHqV0_0(.din(n10772), .dout(n10769));
    jdff dff_A_NClwg5zS3_0(.din(n10775), .dout(n10772));
    jdff dff_A_28EEJ0Sn8_0(.din(n10778), .dout(n10775));
    jdff dff_A_3rZZEYLc6_0(.din(n10781), .dout(n10778));
    jdff dff_A_MEGH1NvO4_0(.din(n10784), .dout(n10781));
    jdff dff_A_uCmTs7TH7_0(.din(n10787), .dout(n10784));
    jdff dff_A_6TImLwIf6_0(.din(n10790), .dout(n10787));
    jdff dff_A_kYHBqgOM8_0(.din(n10793), .dout(n10790));
    jdff dff_A_VWP2JInt9_0(.din(n10796), .dout(n10793));
    jdff dff_A_H10i0gnZ4_0(.din(n1952), .dout(n10796));
    jdff dff_A_UdIxKefW1_2(.din(n10802), .dout(n10799));
    jdff dff_A_RFYth3pu9_2(.din(n10805), .dout(n10802));
    jdff dff_A_O7ydR7cm8_2(.din(n10808), .dout(n10805));
    jdff dff_A_OV09zMKu6_2(.din(n10811), .dout(n10808));
    jdff dff_A_0HMKhCxd2_2(.din(n10814), .dout(n10811));
    jdff dff_A_393srodo3_2(.din(n10817), .dout(n10814));
    jdff dff_A_LTo0MXWQ5_2(.din(n10820), .dout(n10817));
    jdff dff_A_BovatdL55_2(.din(n10823), .dout(n10820));
    jdff dff_A_icapLlXC4_2(.din(n10826), .dout(n10823));
    jdff dff_A_hqzJ7BUz0_2(.din(n1952), .dout(n10826));
    jdff dff_A_zyQLVVjd6_1(.din(n10832), .dout(n10829));
    jdff dff_A_Oye7c9t85_1(.din(n10835), .dout(n10832));
    jdff dff_A_AaWsLxke0_1(.din(n1952), .dout(n10835));
    jdff dff_A_cByZCHFb3_2(.din(n10841), .dout(n10838));
    jdff dff_A_MzwhkeoN1_2(.din(n1952), .dout(n10841));
    jdff dff_A_VwmtA1gA7_1(.din(n10847), .dout(n10844));
    jdff dff_A_Z2XBsqBC9_1(.din(n10850), .dout(n10847));
    jdff dff_A_AfCrQjjM0_1(.din(n10853), .dout(n10850));
    jdff dff_A_PuTXQgIf1_1(.din(n10856), .dout(n10853));
    jdff dff_A_az5jMjMD1_1(.din(n1948), .dout(n10856));
    jdff dff_A_q0CypoSz6_2(.din(n10862), .dout(n10859));
    jdff dff_A_QXZO0qHl4_2(.din(n10865), .dout(n10862));
    jdff dff_A_IHj1ibR70_2(.din(n10868), .dout(n10865));
    jdff dff_A_JJmQXtTo5_2(.din(n10871), .dout(n10868));
    jdff dff_A_00kALzpj4_2(.din(n1948), .dout(n10871));
    jdff dff_A_lJ5nagS34_0(.din(G213), .dout(n10874));
    jdff dff_A_fFX9Wa6W5_2(.din(n10880), .dout(n10877));
    jdff dff_A_raF79JIE4_2(.din(G213), .dout(n10880));
    jdff dff_A_5xFSuWWJ2_1(.din(n10886), .dout(n10883));
    jdff dff_A_VH4fbc1h7_1(.din(n10889), .dout(n10886));
    jdff dff_A_mLMEhh1X3_1(.din(n10892), .dout(n10889));
    jdff dff_A_aA2Efb6n2_1(.din(G343), .dout(n10892));
    jdff dff_A_PyGxFW0l7_2(.din(n545), .dout(n10895));
    jdff dff_B_GES3CfPU6_1(.din(n526), .dout(n10899));
    jdff dff_B_tISGEVh33_1(.din(n10899), .dout(n10902));
    jdff dff_A_3jLZoVp15_1(.din(n10913), .dout(n10904));
    jdff dff_A_ZmYTtGjP7_2(.din(n10910), .dout(n10907));
    jdff dff_A_hxtQ4qkq4_2(.din(n10913), .dout(n10910));
    jdff dff_A_eXXOSfVr4_0(.din(n10916), .dout(n10913));
    jdff dff_A_pg2YfUI82_0(.din(n10919), .dout(n10916));
    jdff dff_A_gKdiZiIb8_0(.din(n10922), .dout(n10919));
    jdff dff_A_25PEjoF99_0(.din(n10925), .dout(n10922));
    jdff dff_A_e7aAggJJ6_0(.din(n10928), .dout(n10925));
    jdff dff_A_oUdYKSkV9_0(.din(n10931), .dout(n10928));
    jdff dff_A_AOAazSbn8_0(.din(G190), .dout(n10931));
    jdff dff_A_268u0N709_2(.din(n10937), .dout(n10934));
    jdff dff_A_KUBNllBB7_2(.din(n10940), .dout(n10937));
    jdff dff_A_ZC8WDYmo0_2(.din(n10943), .dout(n10940));
    jdff dff_A_mrfJpwXB4_2(.din(n10946), .dout(n10943));
    jdff dff_A_WrRtgUhA4_2(.din(n10949), .dout(n10946));
    jdff dff_A_Xcuel7Tg7_2(.din(n10952), .dout(n10949));
    jdff dff_A_TufCRslF2_2(.din(G190), .dout(n10952));
    jdff dff_A_iPX7Z4Cu9_2(.din(n10958), .dout(n10955));
    jdff dff_A_VefTAxdH1_2(.din(n10961), .dout(n10958));
    jdff dff_A_cXO4wwz39_2(.din(n10964), .dout(n10961));
    jdff dff_A_Ldn2NI1j8_2(.din(n10967), .dout(n10964));
    jdff dff_A_ttA7cKY37_2(.din(n10970), .dout(n10967));
    jdff dff_A_jOAji8bc1_2(.din(n10973), .dout(n10970));
    jdff dff_A_8rxErzIf8_2(.din(n10976), .dout(n10973));
    jdff dff_A_7TIFVRkI6_2(.din(G200), .dout(n10976));
    jdff dff_A_NUfNMVn58_1(.din(n10982), .dout(n10979));
    jdff dff_A_oAfHk9in3_1(.din(n522), .dout(n10982));
    jdff dff_B_2RLYosgE9_1(.din(n409), .dout(n10986));
    jdff dff_B_4iA5VZ472_1(.din(n10986), .dout(n10989));
    jdff dff_A_Uw9rA5Q79_1(.din(n514), .dout(n10991));
    jdff dff_A_maUN2Flg6_1(.din(n11018), .dout(n10994));
    jdff dff_A_gb7dweU23_2(.din(n11018), .dout(n10997));
    jdff dff_A_PeA8ptfg2_0(.din(n11003), .dout(n11000));
    jdff dff_A_VNirrpwN2_0(.din(n11006), .dout(n11003));
    jdff dff_A_50kHApfg2_0(.din(n11009), .dout(n11006));
    jdff dff_A_o4b01Lh21_0(.din(n11012), .dout(n11009));
    jdff dff_A_Ji9HKJb18_0(.din(n11015), .dout(n11012));
    jdff dff_A_oKT7Ez0f7_0(.din(n510), .dout(n11015));
    jdff dff_A_xpS69ZrS3_1(.din(n11021), .dout(n11018));
    jdff dff_A_yJts9i7G6_1(.din(n11024), .dout(n11021));
    jdff dff_A_2yzE9Y8S6_1(.din(n11027), .dout(n11024));
    jdff dff_A_eM4pA4l30_1(.din(n11030), .dout(n11027));
    jdff dff_A_vn0SLuPI6_1(.din(n11033), .dout(n11030));
    jdff dff_A_FPx0BJSn6_1(.din(n510), .dout(n11033));
    jdff dff_A_UFx35RBF0_0(.din(n11039), .dout(n11036));
    jdff dff_A_uVC9z8PY3_0(.din(n11042), .dout(n11039));
    jdff dff_A_HS9Rn81n8_0(.din(n11045), .dout(n11042));
    jdff dff_A_bSnjeapd9_0(.din(n11048), .dout(n11045));
    jdff dff_A_Gbdxrt8p0_0(.din(n11051), .dout(n11048));
    jdff dff_A_jzvCaJzW7_0(.din(n11054), .dout(n11051));
    jdff dff_A_W5jceAN66_0(.din(n11057), .dout(n11054));
    jdff dff_A_adNHm5Ts5_0(.din(G179), .dout(n11057));
    jdff dff_A_VNW6KaN29_1(.din(n11063), .dout(n11060));
    jdff dff_A_Pncs4or61_1(.din(n11066), .dout(n11063));
    jdff dff_A_cQgTutSB9_1(.din(n11069), .dout(n11066));
    jdff dff_A_n8LNq6bN8_1(.din(n11072), .dout(n11069));
    jdff dff_A_JGeeLpHH8_1(.din(n11075), .dout(n11072));
    jdff dff_A_6CZSu0Gw2_1(.din(n11078), .dout(n11075));
    jdff dff_A_zdPn62Q54_1(.din(n11081), .dout(n11078));
    jdff dff_A_C1uqPPe31_1(.din(G179), .dout(n11081));
    jdff dff_A_9CGFR2918_0(.din(n11087), .dout(n11084));
    jdff dff_A_cB6r0kEd9_0(.din(n11090), .dout(n11087));
    jdff dff_A_PJ0ANXx23_0(.din(n11093), .dout(n11090));
    jdff dff_A_d28yZRUN3_0(.din(n11096), .dout(n11093));
    jdff dff_A_8qmwtbr90_0(.din(n11099), .dout(n11096));
    jdff dff_A_dJhGqiUZ6_0(.din(n11102), .dout(n11099));
    jdff dff_A_RyIK6iYs2_0(.din(n11105), .dout(n11102));
    jdff dff_A_kBLVlvFw4_0(.din(G179), .dout(n11105));
    jdff dff_A_SyzkO7SL4_1(.din(n500), .dout(n11108));
    jdff dff_B_GcnqWhjj5_0(.din(n492), .dout(n11112));
    jdff dff_A_21LTCwyy0_0(.din(n11117), .dout(n11114));
    jdff dff_A_5Os4Co0L7_0(.din(n11120), .dout(n11117));
    jdff dff_A_D30XsiAm4_0(.din(G270), .dout(n11120));
    jdff dff_A_AYEVyLfQ3_1(.din(G270), .dout(n11123));
    jdff dff_B_dI5peQw07_1(.din(n454), .dout(n11127));
    jdff dff_B_SJl0iTHM2_1(.din(n458), .dout(n11130));
    jdff dff_B_BgZDjfnJ5_1(.din(n11130), .dout(n11133));
    jdff dff_A_Yay1H0sT4_0(.din(n11138), .dout(n11135));
    jdff dff_A_XjVZ48HX4_0(.din(G257), .dout(n11138));
    jdff dff_A_8O7tS3tU4_1(.din(n11144), .dout(n11141));
    jdff dff_A_axQXsGFK3_1(.din(n11147), .dout(n11144));
    jdff dff_A_LseBYIOK8_1(.din(G257), .dout(n11147));
    jdff dff_A_DwDyRc4z4_2(.din(n11153), .dout(n11150));
    jdff dff_A_TGsmLIqQ6_2(.din(G257), .dout(n11153));
    jdff dff_A_sAjQKnIV0_0(.din(n11159), .dout(n11156));
    jdff dff_A_25Ixg5Bz5_0(.din(n11162), .dout(n11159));
    jdff dff_A_hMpawB0o6_0(.din(G303), .dout(n11162));
    jdff dff_A_J7DcwswV9_1(.din(n11168), .dout(n11165));
    jdff dff_A_VvwDY8HE4_1(.din(n11171), .dout(n11168));
    jdff dff_A_Z1eKN7YO8_1(.din(G303), .dout(n11171));
    jdff dff_A_tA4WwVps9_0(.din(n11177), .dout(n11174));
    jdff dff_A_MY4gmzcB6_0(.din(n11180), .dout(n11177));
    jdff dff_A_5em3aR5A7_0(.din(G303), .dout(n11180));
    jdff dff_A_Yu7uDWyd5_2(.din(n11186), .dout(n11183));
    jdff dff_A_jhzE4bo43_2(.din(n11189), .dout(n11186));
    jdff dff_A_K6oeFYj22_2(.din(n11192), .dout(n11189));
    jdff dff_A_qt1GiljN0_2(.din(G303), .dout(n11192));
    jdff dff_A_rzrEgui05_2(.din(G1698), .dout(n11195));
    jdff dff_A_m34ss2Ex2_0(.din(n11201), .dout(n11198));
    jdff dff_A_2kBUp0gP7_0(.din(n11204), .dout(n11201));
    jdff dff_A_B212phLv9_0(.din(G264), .dout(n11204));
    jdff dff_A_iK7dFzir4_1(.din(n11210), .dout(n11207));
    jdff dff_A_ahXSG8UL4_1(.din(G264), .dout(n11210));
    jdff dff_A_ceBD7C2p2_1(.din(n11216), .dout(n11213));
    jdff dff_A_re8iwzaB9_1(.din(n446), .dout(n11216));
    jdff dff_A_GVkq5jlA9_2(.din(n11222), .dout(n11219));
    jdff dff_A_qhl06zxv1_2(.din(n446), .dout(n11222));
    jdff dff_A_XKjLqvyA4_1(.din(n11228), .dout(n11225));
    jdff dff_A_NwQFKoZl5_1(.din(n446), .dout(n11228));
    jdff dff_A_bW7EyHf57_2(.din(n11234), .dout(n11231));
    jdff dff_A_dZmAmqcr4_2(.din(n446), .dout(n11234));
    jdff dff_A_MW926Uyt6_1(.din(n11240), .dout(n11237));
endmodule

