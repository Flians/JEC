/*
rf_max:
	jspl: 725
	jspl3: 1027
	jnot: 1034
	jand: 1780
	jor: 1381

Summary:
	jspl: 725
	jspl3: 1027
	jnot: 1034
	jand: 1780
	jor: 1381

The maximum logic level gap of any gate:
	rf_max: 106
*/

module rf_max(gclk, in0, in1, in2, in3, result, address);
	input gclk;
	input [127:0] in0;
	input [127:0] in1;
	input [127:0] in2;
	input [127:0] in3;
	output [127:0] result;
	output [1:0] address;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1903;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1921;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1976;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1994;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2006;
	wire n2007;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2011;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2049;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2067;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2102;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2122;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2140;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2195;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2204;
	wire n2205;
	wire n2206;
	wire n2207;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2213;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2230;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2237;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2247;
	wire n2248;
	wire n2249;
	wire n2250;
	wire n2251;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2264;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2268;
	wire n2269;
	wire n2270;
	wire n2271;
	wire n2272;
	wire n2273;
	wire n2274;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2281;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2298;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2315;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2332;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2341;
	wire n2342;
	wire n2343;
	wire n2344;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2349;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2366;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2383;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2400;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2414;
	wire n2415;
	wire n2416;
	wire n2417;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2421;
	wire n2422;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2426;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2431;
	wire n2432;
	wire n2433;
	wire n2434;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2448;
	wire n2449;
	wire n2450;
	wire n2451;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2465;
	wire n2466;
	wire n2467;
	wire n2468;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2482;
	wire n2483;
	wire n2484;
	wire n2485;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2499;
	wire n2500;
	wire n2501;
	wire n2502;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2516;
	wire n2517;
	wire n2518;
	wire n2519;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2533;
	wire n2534;
	wire n2535;
	wire n2536;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2550;
	wire n2551;
	wire n2552;
	wire n2553;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2562;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2567;
	wire n2568;
	wire n2569;
	wire n2570;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2584;
	wire n2585;
	wire n2586;
	wire n2587;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2601;
	wire n2602;
	wire n2603;
	wire n2604;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2618;
	wire n2619;
	wire n2620;
	wire n2621;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2631;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2635;
	wire n2636;
	wire n2637;
	wire n2638;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2652;
	wire n2653;
	wire n2654;
	wire n2655;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2669;
	wire n2670;
	wire n2671;
	wire n2672;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2686;
	wire n2687;
	wire n2688;
	wire n2689;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2703;
	wire n2704;
	wire n2705;
	wire n2706;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2718;
	wire n2719;
	wire n2720;
	wire n2721;
	wire n2722;
	wire n2723;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2731;
	wire n2732;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2737;
	wire n2738;
	wire n2739;
	wire n2740;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2745;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2754;
	wire n2755;
	wire n2756;
	wire n2757;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2771;
	wire n2772;
	wire n2773;
	wire n2774;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2788;
	wire n2789;
	wire n2790;
	wire n2791;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2805;
	wire n2806;
	wire n2807;
	wire n2808;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2822;
	wire n2823;
	wire n2824;
	wire n2825;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2832;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2839;
	wire n2840;
	wire n2841;
	wire n2842;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2856;
	wire n2857;
	wire n2858;
	wire n2859;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2871;
	wire n2872;
	wire n2873;
	wire n2874;
	wire n2875;
	wire n2876;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2890;
	wire n2891;
	wire n2892;
	wire n2893;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2907;
	wire n2908;
	wire n2909;
	wire n2910;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2924;
	wire n2925;
	wire n2926;
	wire n2927;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2941;
	wire n2942;
	wire n2943;
	wire n2944;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2958;
	wire n2959;
	wire n2960;
	wire n2961;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2975;
	wire n2976;
	wire n2977;
	wire n2978;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2992;
	wire n2993;
	wire n2994;
	wire n2995;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3009;
	wire n3010;
	wire n3011;
	wire n3012;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3026;
	wire n3027;
	wire n3028;
	wire n3029;
	wire n3030;
	wire n3031;
	wire n3032;
	wire n3033;
	wire n3034;
	wire n3035;
	wire n3036;
	wire n3037;
	wire n3038;
	wire n3039;
	wire n3040;
	wire n3041;
	wire n3042;
	wire n3043;
	wire n3044;
	wire n3045;
	wire n3046;
	wire n3047;
	wire n3048;
	wire n3049;
	wire n3050;
	wire n3051;
	wire n3052;
	wire n3053;
	wire n3054;
	wire n3055;
	wire n3056;
	wire n3057;
	wire n3058;
	wire n3059;
	wire n3060;
	wire n3061;
	wire n3062;
	wire n3063;
	wire n3064;
	wire n3065;
	wire n3066;
	wire n3067;
	wire n3068;
	wire n3069;
	wire n3070;
	wire n3071;
	wire n3072;
	wire n3073;
	wire n3074;
	wire n3075;
	wire n3076;
	wire n3077;
	wire n3078;
	wire n3079;
	wire n3080;
	wire n3081;
	wire n3082;
	wire n3083;
	wire n3084;
	wire n3085;
	wire n3086;
	wire n3087;
	wire n3088;
	wire n3089;
	wire n3090;
	wire n3091;
	wire n3092;
	wire n3093;
	wire n3094;
	wire n3095;
	wire n3096;
	wire n3097;
	wire n3098;
	wire n3099;
	wire n3100;
	wire n3101;
	wire n3102;
	wire n3103;
	wire n3104;
	wire n3105;
	wire n3106;
	wire n3107;
	wire n3108;
	wire n3109;
	wire n3110;
	wire n3111;
	wire n3112;
	wire n3113;
	wire n3114;
	wire n3115;
	wire n3116;
	wire n3117;
	wire n3118;
	wire n3119;
	wire n3120;
	wire n3121;
	wire n3122;
	wire n3123;
	wire n3124;
	wire n3125;
	wire n3126;
	wire n3127;
	wire n3128;
	wire n3129;
	wire n3130;
	wire n3131;
	wire n3132;
	wire n3133;
	wire n3134;
	wire n3135;
	wire n3136;
	wire n3137;
	wire n3138;
	wire n3139;
	wire n3140;
	wire n3141;
	wire n3142;
	wire n3143;
	wire n3144;
	wire n3145;
	wire n3146;
	wire n3147;
	wire n3148;
	wire n3149;
	wire n3150;
	wire n3151;
	wire n3152;
	wire n3153;
	wire n3154;
	wire n3155;
	wire n3156;
	wire n3157;
	wire n3158;
	wire n3159;
	wire n3160;
	wire n3161;
	wire n3162;
	wire n3163;
	wire n3164;
	wire n3165;
	wire n3166;
	wire n3167;
	wire n3168;
	wire n3169;
	wire n3170;
	wire n3171;
	wire n3172;
	wire n3173;
	wire n3174;
	wire n3175;
	wire n3176;
	wire n3177;
	wire n3178;
	wire n3179;
	wire n3180;
	wire n3181;
	wire n3182;
	wire n3183;
	wire n3184;
	wire n3185;
	wire n3186;
	wire n3187;
	wire n3188;
	wire n3189;
	wire n3190;
	wire n3191;
	wire n3192;
	wire n3193;
	wire n3194;
	wire n3195;
	wire n3196;
	wire n3197;
	wire n3198;
	wire n3199;
	wire n3200;
	wire n3201;
	wire n3202;
	wire n3203;
	wire n3204;
	wire n3205;
	wire n3206;
	wire n3207;
	wire n3208;
	wire n3209;
	wire n3210;
	wire n3211;
	wire n3212;
	wire n3213;
	wire n3214;
	wire n3215;
	wire n3216;
	wire n3217;
	wire n3218;
	wire n3219;
	wire n3220;
	wire n3221;
	wire n3222;
	wire n3223;
	wire n3224;
	wire n3225;
	wire n3226;
	wire n3227;
	wire n3228;
	wire n3229;
	wire n3230;
	wire n3231;
	wire n3232;
	wire n3233;
	wire n3234;
	wire n3235;
	wire n3236;
	wire n3237;
	wire n3238;
	wire n3239;
	wire n3240;
	wire n3241;
	wire n3242;
	wire n3243;
	wire n3244;
	wire n3245;
	wire n3246;
	wire n3247;
	wire n3248;
	wire n3249;
	wire n3250;
	wire n3251;
	wire n3252;
	wire n3253;
	wire n3254;
	wire n3255;
	wire n3256;
	wire n3257;
	wire n3258;
	wire n3259;
	wire n3260;
	wire n3261;
	wire n3262;
	wire n3263;
	wire n3264;
	wire n3265;
	wire n3266;
	wire n3267;
	wire n3268;
	wire n3269;
	wire n3270;
	wire n3271;
	wire n3272;
	wire n3273;
	wire n3274;
	wire n3275;
	wire n3276;
	wire n3277;
	wire n3278;
	wire n3279;
	wire n3280;
	wire n3281;
	wire n3282;
	wire n3283;
	wire n3284;
	wire n3285;
	wire n3286;
	wire n3287;
	wire n3288;
	wire n3289;
	wire n3290;
	wire n3291;
	wire n3292;
	wire n3293;
	wire n3294;
	wire n3295;
	wire n3296;
	wire n3297;
	wire n3298;
	wire n3299;
	wire n3300;
	wire n3301;
	wire n3302;
	wire n3303;
	wire n3304;
	wire n3305;
	wire n3306;
	wire n3307;
	wire n3308;
	wire n3309;
	wire n3310;
	wire n3311;
	wire n3312;
	wire n3313;
	wire n3314;
	wire n3315;
	wire n3316;
	wire n3317;
	wire n3318;
	wire n3319;
	wire n3320;
	wire n3321;
	wire n3322;
	wire n3323;
	wire n3324;
	wire n3325;
	wire n3326;
	wire n3327;
	wire n3328;
	wire n3329;
	wire n3330;
	wire n3331;
	wire n3332;
	wire n3333;
	wire n3334;
	wire n3335;
	wire n3336;
	wire n3337;
	wire n3338;
	wire n3339;
	wire n3340;
	wire n3341;
	wire n3342;
	wire n3343;
	wire n3344;
	wire n3345;
	wire n3346;
	wire n3347;
	wire n3348;
	wire n3349;
	wire n3350;
	wire n3351;
	wire n3352;
	wire n3353;
	wire n3354;
	wire n3355;
	wire n3356;
	wire n3357;
	wire n3358;
	wire n3359;
	wire n3360;
	wire n3361;
	wire n3362;
	wire n3363;
	wire n3364;
	wire n3365;
	wire n3366;
	wire n3367;
	wire n3368;
	wire n3369;
	wire n3370;
	wire n3371;
	wire n3372;
	wire n3373;
	wire n3374;
	wire n3375;
	wire n3376;
	wire n3377;
	wire n3378;
	wire n3379;
	wire n3380;
	wire n3381;
	wire n3382;
	wire n3383;
	wire n3384;
	wire n3385;
	wire n3386;
	wire n3387;
	wire n3388;
	wire n3389;
	wire n3390;
	wire n3391;
	wire n3392;
	wire n3393;
	wire n3394;
	wire n3395;
	wire n3396;
	wire n3397;
	wire n3398;
	wire n3399;
	wire n3400;
	wire n3401;
	wire n3402;
	wire n3403;
	wire n3404;
	wire n3405;
	wire n3406;
	wire n3407;
	wire n3408;
	wire n3409;
	wire n3410;
	wire n3411;
	wire n3412;
	wire n3413;
	wire n3414;
	wire n3415;
	wire n3416;
	wire n3417;
	wire n3418;
	wire n3419;
	wire n3420;
	wire n3421;
	wire n3422;
	wire n3423;
	wire n3424;
	wire n3425;
	wire n3426;
	wire n3427;
	wire n3428;
	wire n3429;
	wire n3430;
	wire n3431;
	wire n3432;
	wire n3433;
	wire n3434;
	wire n3435;
	wire n3436;
	wire n3437;
	wire n3438;
	wire n3439;
	wire n3440;
	wire n3441;
	wire n3442;
	wire n3443;
	wire n3444;
	wire n3445;
	wire n3446;
	wire n3447;
	wire n3448;
	wire n3449;
	wire n3450;
	wire n3451;
	wire n3452;
	wire n3453;
	wire n3454;
	wire n3455;
	wire n3456;
	wire n3457;
	wire n3458;
	wire n3459;
	wire n3460;
	wire n3461;
	wire n3462;
	wire n3463;
	wire n3464;
	wire n3465;
	wire n3466;
	wire n3467;
	wire n3468;
	wire n3469;
	wire n3470;
	wire n3471;
	wire n3472;
	wire n3473;
	wire n3474;
	wire n3475;
	wire n3476;
	wire n3477;
	wire n3478;
	wire n3479;
	wire n3480;
	wire n3481;
	wire n3482;
	wire n3483;
	wire n3484;
	wire n3485;
	wire n3486;
	wire n3487;
	wire n3488;
	wire n3489;
	wire n3490;
	wire n3491;
	wire n3492;
	wire n3493;
	wire n3494;
	wire n3495;
	wire n3496;
	wire n3497;
	wire n3498;
	wire n3499;
	wire n3500;
	wire n3501;
	wire n3502;
	wire n3503;
	wire n3504;
	wire n3505;
	wire n3506;
	wire n3507;
	wire n3508;
	wire n3509;
	wire n3510;
	wire n3511;
	wire n3512;
	wire n3513;
	wire n3514;
	wire n3515;
	wire n3516;
	wire n3517;
	wire n3518;
	wire n3519;
	wire n3520;
	wire n3521;
	wire n3522;
	wire n3523;
	wire n3524;
	wire n3525;
	wire n3526;
	wire n3527;
	wire n3528;
	wire n3529;
	wire n3530;
	wire n3531;
	wire n3532;
	wire n3533;
	wire n3534;
	wire n3535;
	wire n3536;
	wire n3537;
	wire n3538;
	wire n3539;
	wire n3540;
	wire n3541;
	wire n3542;
	wire n3543;
	wire n3544;
	wire n3545;
	wire n3546;
	wire n3547;
	wire n3548;
	wire n3549;
	wire n3550;
	wire n3551;
	wire n3552;
	wire n3553;
	wire n3554;
	wire n3555;
	wire n3556;
	wire n3557;
	wire n3558;
	wire n3559;
	wire n3560;
	wire n3561;
	wire n3562;
	wire n3563;
	wire n3564;
	wire n3565;
	wire n3566;
	wire n3567;
	wire n3568;
	wire n3569;
	wire n3570;
	wire n3571;
	wire n3572;
	wire n3573;
	wire n3574;
	wire n3575;
	wire n3576;
	wire n3577;
	wire n3578;
	wire n3579;
	wire n3580;
	wire n3581;
	wire n3582;
	wire n3583;
	wire n3584;
	wire n3585;
	wire n3586;
	wire n3587;
	wire n3588;
	wire n3589;
	wire n3590;
	wire n3591;
	wire n3592;
	wire n3593;
	wire n3594;
	wire n3595;
	wire n3596;
	wire n3597;
	wire n3598;
	wire n3599;
	wire n3600;
	wire n3601;
	wire n3602;
	wire n3603;
	wire n3604;
	wire n3605;
	wire n3606;
	wire n3607;
	wire n3608;
	wire n3609;
	wire n3610;
	wire n3611;
	wire n3612;
	wire n3613;
	wire n3614;
	wire n3615;
	wire n3616;
	wire n3617;
	wire n3618;
	wire n3619;
	wire n3620;
	wire n3621;
	wire n3622;
	wire n3623;
	wire n3624;
	wire n3625;
	wire n3626;
	wire n3627;
	wire n3628;
	wire n3629;
	wire n3630;
	wire n3631;
	wire n3632;
	wire n3633;
	wire n3634;
	wire n3635;
	wire n3636;
	wire n3637;
	wire n3638;
	wire n3639;
	wire n3640;
	wire n3641;
	wire n3642;
	wire n3643;
	wire n3644;
	wire n3645;
	wire n3646;
	wire n3647;
	wire n3648;
	wire n3649;
	wire n3650;
	wire n3651;
	wire n3652;
	wire n3653;
	wire n3654;
	wire n3655;
	wire n3656;
	wire n3657;
	wire n3658;
	wire n3659;
	wire n3660;
	wire n3661;
	wire n3662;
	wire n3663;
	wire n3664;
	wire n3665;
	wire n3666;
	wire n3667;
	wire n3668;
	wire n3669;
	wire n3670;
	wire n3671;
	wire n3672;
	wire n3673;
	wire n3674;
	wire n3675;
	wire n3676;
	wire n3677;
	wire n3678;
	wire n3679;
	wire n3680;
	wire n3681;
	wire n3682;
	wire n3683;
	wire n3684;
	wire n3685;
	wire n3686;
	wire n3687;
	wire n3688;
	wire n3689;
	wire n3690;
	wire n3691;
	wire n3692;
	wire n3693;
	wire n3694;
	wire n3695;
	wire n3696;
	wire n3697;
	wire n3698;
	wire n3699;
	wire n3700;
	wire n3701;
	wire n3702;
	wire n3703;
	wire n3704;
	wire n3705;
	wire n3706;
	wire n3707;
	wire n3708;
	wire n3709;
	wire n3710;
	wire n3711;
	wire n3712;
	wire n3713;
	wire n3714;
	wire n3715;
	wire n3716;
	wire n3717;
	wire n3718;
	wire n3719;
	wire n3720;
	wire n3721;
	wire n3722;
	wire n3723;
	wire n3724;
	wire n3725;
	wire n3726;
	wire n3727;
	wire n3728;
	wire n3729;
	wire n3730;
	wire n3731;
	wire n3732;
	wire n3733;
	wire n3734;
	wire n3735;
	wire n3736;
	wire n3737;
	wire n3738;
	wire n3739;
	wire n3740;
	wire n3741;
	wire n3742;
	wire n3743;
	wire n3744;
	wire n3745;
	wire n3746;
	wire n3747;
	wire n3748;
	wire n3749;
	wire n3750;
	wire n3751;
	wire n3752;
	wire n3753;
	wire n3754;
	wire n3755;
	wire n3756;
	wire n3757;
	wire n3758;
	wire n3759;
	wire n3760;
	wire n3761;
	wire n3762;
	wire n3763;
	wire n3764;
	wire n3765;
	wire n3766;
	wire n3767;
	wire n3768;
	wire n3769;
	wire n3770;
	wire n3771;
	wire n3772;
	wire n3773;
	wire n3774;
	wire n3775;
	wire n3776;
	wire n3777;
	wire n3778;
	wire n3779;
	wire n3780;
	wire n3781;
	wire n3782;
	wire n3783;
	wire n3784;
	wire n3785;
	wire n3786;
	wire n3787;
	wire n3788;
	wire n3789;
	wire n3790;
	wire n3791;
	wire n3792;
	wire n3793;
	wire n3794;
	wire n3795;
	wire n3796;
	wire n3797;
	wire n3798;
	wire n3799;
	wire n3800;
	wire n3801;
	wire n3802;
	wire n3803;
	wire n3804;
	wire n3805;
	wire n3806;
	wire n3807;
	wire n3808;
	wire n3809;
	wire n3810;
	wire n3811;
	wire n3812;
	wire n3813;
	wire n3814;
	wire n3815;
	wire n3816;
	wire n3817;
	wire n3818;
	wire n3819;
	wire n3820;
	wire n3821;
	wire n3822;
	wire n3823;
	wire n3824;
	wire n3825;
	wire n3826;
	wire n3827;
	wire n3828;
	wire n3829;
	wire n3830;
	wire n3831;
	wire n3832;
	wire n3833;
	wire n3834;
	wire n3835;
	wire n3836;
	wire n3837;
	wire n3838;
	wire n3839;
	wire n3840;
	wire n3841;
	wire n3842;
	wire n3843;
	wire n3844;
	wire n3845;
	wire n3846;
	wire n3847;
	wire n3848;
	wire n3849;
	wire n3850;
	wire n3851;
	wire n3852;
	wire n3853;
	wire n3854;
	wire n3855;
	wire n3856;
	wire n3857;
	wire n3858;
	wire n3859;
	wire n3860;
	wire n3861;
	wire n3862;
	wire n3863;
	wire n3864;
	wire n3865;
	wire n3866;
	wire n3867;
	wire n3868;
	wire n3869;
	wire n3870;
	wire n3871;
	wire n3872;
	wire n3873;
	wire n3874;
	wire n3875;
	wire n3876;
	wire n3877;
	wire n3878;
	wire n3879;
	wire n3880;
	wire n3881;
	wire n3882;
	wire n3883;
	wire n3884;
	wire n3885;
	wire n3886;
	wire n3887;
	wire n3888;
	wire n3889;
	wire n3890;
	wire n3891;
	wire n3892;
	wire n3893;
	wire n3894;
	wire n3895;
	wire n3896;
	wire n3897;
	wire n3898;
	wire n3899;
	wire n3900;
	wire n3901;
	wire n3902;
	wire n3903;
	wire n3904;
	wire n3905;
	wire n3906;
	wire n3907;
	wire n3908;
	wire n3909;
	wire n3910;
	wire n3911;
	wire n3912;
	wire n3913;
	wire n3914;
	wire n3915;
	wire n3916;
	wire n3917;
	wire n3918;
	wire n3919;
	wire n3920;
	wire n3921;
	wire n3922;
	wire n3923;
	wire n3924;
	wire n3925;
	wire n3926;
	wire n3927;
	wire n3928;
	wire n3929;
	wire n3930;
	wire n3931;
	wire n3932;
	wire n3933;
	wire n3934;
	wire n3935;
	wire n3936;
	wire n3937;
	wire n3938;
	wire n3939;
	wire n3940;
	wire n3941;
	wire n3942;
	wire n3943;
	wire n3944;
	wire n3945;
	wire n3946;
	wire n3947;
	wire n3948;
	wire n3949;
	wire n3950;
	wire n3951;
	wire n3952;
	wire n3953;
	wire n3954;
	wire n3955;
	wire n3956;
	wire n3957;
	wire n3958;
	wire n3959;
	wire n3960;
	wire n3961;
	wire n3962;
	wire n3963;
	wire n3964;
	wire n3965;
	wire n3966;
	wire n3967;
	wire n3968;
	wire n3969;
	wire n3970;
	wire n3971;
	wire n3972;
	wire n3973;
	wire n3974;
	wire n3975;
	wire n3976;
	wire n3977;
	wire n3978;
	wire n3979;
	wire n3980;
	wire n3981;
	wire n3982;
	wire n3983;
	wire n3984;
	wire n3985;
	wire n3986;
	wire n3987;
	wire n3988;
	wire n3989;
	wire n3990;
	wire n3991;
	wire n3992;
	wire n3993;
	wire n3994;
	wire n3995;
	wire n3996;
	wire n3997;
	wire n3998;
	wire n3999;
	wire n4000;
	wire n4001;
	wire n4002;
	wire n4003;
	wire n4004;
	wire n4005;
	wire n4006;
	wire n4007;
	wire n4008;
	wire n4009;
	wire n4010;
	wire n4011;
	wire n4012;
	wire n4013;
	wire n4014;
	wire n4015;
	wire n4016;
	wire n4017;
	wire n4018;
	wire n4019;
	wire n4020;
	wire n4021;
	wire n4022;
	wire n4023;
	wire n4024;
	wire n4025;
	wire n4026;
	wire n4027;
	wire n4028;
	wire n4029;
	wire n4030;
	wire n4031;
	wire n4032;
	wire n4033;
	wire n4034;
	wire n4035;
	wire n4036;
	wire n4037;
	wire n4038;
	wire n4039;
	wire n4040;
	wire n4041;
	wire n4042;
	wire n4043;
	wire n4044;
	wire n4045;
	wire n4046;
	wire n4047;
	wire n4048;
	wire n4049;
	wire n4050;
	wire n4051;
	wire n4052;
	wire n4053;
	wire n4054;
	wire n4055;
	wire n4056;
	wire n4057;
	wire n4058;
	wire n4059;
	wire n4060;
	wire n4061;
	wire n4062;
	wire n4063;
	wire n4064;
	wire n4065;
	wire n4066;
	wire n4067;
	wire n4068;
	wire n4069;
	wire n4070;
	wire n4071;
	wire n4072;
	wire n4073;
	wire n4074;
	wire n4075;
	wire n4076;
	wire n4077;
	wire n4078;
	wire n4079;
	wire n4080;
	wire n4081;
	wire n4082;
	wire n4083;
	wire n4084;
	wire n4085;
	wire n4086;
	wire n4087;
	wire n4088;
	wire n4089;
	wire n4090;
	wire n4091;
	wire n4092;
	wire n4093;
	wire n4094;
	wire n4095;
	wire n4096;
	wire n4097;
	wire n4098;
	wire n4099;
	wire n4100;
	wire n4101;
	wire n4102;
	wire n4103;
	wire n4104;
	wire n4105;
	wire n4106;
	wire n4107;
	wire n4108;
	wire n4109;
	wire n4110;
	wire n4111;
	wire n4112;
	wire n4113;
	wire n4114;
	wire n4115;
	wire n4116;
	wire n4117;
	wire n4118;
	wire n4119;
	wire n4120;
	wire n4121;
	wire n4122;
	wire n4123;
	wire n4124;
	wire n4125;
	wire n4126;
	wire n4127;
	wire n4128;
	wire n4129;
	wire n4130;
	wire n4131;
	wire n4132;
	wire n4133;
	wire n4134;
	wire n4135;
	wire n4136;
	wire n4137;
	wire n4138;
	wire n4139;
	wire n4140;
	wire n4141;
	wire n4142;
	wire n4143;
	wire n4144;
	wire n4145;
	wire n4146;
	wire n4147;
	wire n4148;
	wire n4149;
	wire n4150;
	wire n4151;
	wire n4152;
	wire n4153;
	wire n4154;
	wire n4155;
	wire n4156;
	wire n4157;
	wire n4158;
	wire n4159;
	wire n4160;
	wire n4161;
	wire n4162;
	wire n4163;
	wire n4164;
	wire n4165;
	wire n4166;
	wire n4167;
	wire n4168;
	wire n4169;
	wire n4170;
	wire n4171;
	wire n4172;
	wire n4173;
	wire n4174;
	wire n4175;
	wire n4176;
	wire n4177;
	wire n4178;
	wire n4179;
	wire n4180;
	wire n4181;
	wire n4182;
	wire n4183;
	wire n4184;
	wire n4185;
	wire n4186;
	wire n4187;
	wire n4188;
	wire n4189;
	wire n4190;
	wire n4191;
	wire n4192;
	wire n4193;
	wire n4194;
	wire n4195;
	wire n4196;
	wire n4197;
	wire n4198;
	wire n4199;
	wire n4200;
	wire n4201;
	wire n4202;
	wire n4203;
	wire n4204;
	wire n4205;
	wire n4206;
	wire n4207;
	wire n4208;
	wire n4209;
	wire n4210;
	wire n4211;
	wire n4212;
	wire n4213;
	wire n4214;
	wire n4215;
	wire n4216;
	wire n4217;
	wire n4218;
	wire n4219;
	wire n4220;
	wire n4221;
	wire n4222;
	wire n4223;
	wire n4224;
	wire n4225;
	wire n4226;
	wire n4227;
	wire n4228;
	wire n4229;
	wire n4230;
	wire n4231;
	wire n4232;
	wire n4233;
	wire n4234;
	wire n4235;
	wire n4236;
	wire n4237;
	wire n4238;
	wire n4239;
	wire n4240;
	wire n4241;
	wire n4242;
	wire n4243;
	wire n4244;
	wire n4245;
	wire n4246;
	wire n4247;
	wire n4248;
	wire n4249;
	wire n4250;
	wire n4251;
	wire n4252;
	wire n4253;
	wire n4254;
	wire n4255;
	wire n4256;
	wire n4257;
	wire n4258;
	wire n4259;
	wire n4260;
	wire n4261;
	wire n4262;
	wire n4263;
	wire n4264;
	wire n4265;
	wire n4266;
	wire n4267;
	wire n4268;
	wire n4269;
	wire n4271;
	wire n4272;
	wire n4273;
	wire n4274;
	wire n4275;
	wire n4276;
	wire n4277;
	wire n4278;
	wire n4279;
	wire n4280;
	wire n4281;
	wire n4282;
	wire n4283;
	wire n4284;
	wire n4285;
	wire n4286;
	wire n4287;
	wire n4288;
	wire n4289;
	wire n4290;
	wire n4291;
	wire n4292;
	wire n4293;
	wire n4294;
	wire n4295;
	wire n4296;
	wire n4297;
	wire n4298;
	wire n4299;
	wire n4300;
	wire n4301;
	wire n4302;
	wire n4303;
	wire n4304;
	wire n4305;
	wire n4306;
	wire n4307;
	wire n4308;
	wire n4309;
	wire n4310;
	wire n4311;
	wire n4312;
	wire n4313;
	wire n4314;
	wire n4315;
	wire n4316;
	wire n4317;
	wire n4318;
	wire n4319;
	wire n4320;
	wire n4321;
	wire n4322;
	wire n4323;
	wire n4324;
	wire n4325;
	wire n4326;
	wire n4327;
	wire n4328;
	wire n4329;
	wire n4330;
	wire n4331;
	wire n4332;
	wire n4333;
	wire n4334;
	wire n4335;
	wire n4336;
	wire n4337;
	wire n4338;
	wire n4339;
	wire n4340;
	wire n4341;
	wire n4342;
	wire n4343;
	wire n4344;
	wire n4345;
	wire n4346;
	wire n4347;
	wire n4348;
	wire n4349;
	wire n4350;
	wire n4351;
	wire n4352;
	wire n4353;
	wire n4354;
	wire n4355;
	wire n4356;
	wire n4357;
	wire n4358;
	wire n4359;
	wire n4360;
	wire n4361;
	wire n4362;
	wire n4363;
	wire n4364;
	wire n4365;
	wire n4366;
	wire n4367;
	wire n4368;
	wire n4369;
	wire n4370;
	wire n4371;
	wire n4372;
	wire n4373;
	wire n4374;
	wire n4375;
	wire n4376;
	wire n4377;
	wire n4378;
	wire n4379;
	wire n4380;
	wire n4381;
	wire n4382;
	wire n4383;
	wire n4384;
	wire n4385;
	wire n4386;
	wire n4387;
	wire n4388;
	wire n4389;
	wire n4390;
	wire n4391;
	wire n4392;
	wire n4393;
	wire n4394;
	wire n4395;
	wire n4396;
	wire n4397;
	wire n4398;
	wire n4399;
	wire n4400;
	wire n4401;
	wire n4402;
	wire n4403;
	wire n4404;
	wire n4405;
	wire n4406;
	wire n4407;
	wire n4408;
	wire n4409;
	wire n4410;
	wire n4411;
	wire n4412;
	wire n4413;
	wire n4414;
	wire n4415;
	wire n4416;
	wire n4417;
	wire n4418;
	wire n4419;
	wire n4420;
	wire n4421;
	wire n4422;
	wire n4423;
	wire n4424;
	wire n4425;
	wire n4426;
	wire n4427;
	wire n4428;
	wire n4429;
	wire n4430;
	wire n4431;
	wire n4432;
	wire n4433;
	wire n4434;
	wire n4435;
	wire n4436;
	wire n4437;
	wire n4438;
	wire n4439;
	wire n4440;
	wire n4441;
	wire n4442;
	wire n4443;
	wire n4444;
	wire n4445;
	wire n4446;
	wire n4447;
	wire n4448;
	wire n4449;
	wire n4450;
	wire n4451;
	wire n4452;
	wire n4453;
	wire n4455;
	wire n4456;
	wire n4458;
	wire n4459;
	wire n4461;
	wire n4462;
	wire n4464;
	wire n4465;
	wire n4467;
	wire n4468;
	wire n4470;
	wire n4471;
	wire n4473;
	wire n4474;
	wire n4476;
	wire n4477;
	wire n4479;
	wire n4480;
	wire n4482;
	wire n4483;
	wire n4485;
	wire n4486;
	wire n4488;
	wire n4489;
	wire n4491;
	wire n4492;
	wire n4494;
	wire n4495;
	wire n4497;
	wire n4498;
	wire n4500;
	wire n4501;
	wire n4503;
	wire n4504;
	wire n4506;
	wire n4507;
	wire n4509;
	wire n4510;
	wire n4512;
	wire n4513;
	wire n4515;
	wire n4516;
	wire n4518;
	wire n4519;
	wire n4521;
	wire n4522;
	wire n4524;
	wire n4525;
	wire n4527;
	wire n4528;
	wire n4530;
	wire n4531;
	wire n4533;
	wire n4534;
	wire n4536;
	wire n4537;
	wire n4539;
	wire n4540;
	wire n4542;
	wire n4543;
	wire n4545;
	wire n4546;
	wire n4548;
	wire n4549;
	wire n4551;
	wire n4552;
	wire n4554;
	wire n4555;
	wire n4557;
	wire n4558;
	wire n4560;
	wire n4561;
	wire n4563;
	wire n4564;
	wire n4566;
	wire n4567;
	wire n4569;
	wire n4570;
	wire n4572;
	wire n4573;
	wire n4575;
	wire n4576;
	wire n4578;
	wire n4579;
	wire n4581;
	wire n4582;
	wire n4584;
	wire n4585;
	wire n4587;
	wire n4588;
	wire n4590;
	wire n4591;
	wire n4593;
	wire n4594;
	wire n4596;
	wire n4597;
	wire n4599;
	wire n4600;
	wire n4602;
	wire n4603;
	wire n4605;
	wire n4606;
	wire n4608;
	wire n4609;
	wire n4611;
	wire n4612;
	wire n4614;
	wire n4615;
	wire n4617;
	wire n4618;
	wire n4620;
	wire n4621;
	wire n4623;
	wire n4624;
	wire n4626;
	wire n4627;
	wire n4629;
	wire n4630;
	wire n4632;
	wire n4633;
	wire n4635;
	wire n4636;
	wire n4638;
	wire n4639;
	wire n4641;
	wire n4642;
	wire n4644;
	wire n4645;
	wire n4647;
	wire n4648;
	wire n4650;
	wire n4651;
	wire n4653;
	wire n4654;
	wire n4656;
	wire n4657;
	wire n4659;
	wire n4660;
	wire n4662;
	wire n4663;
	wire n4665;
	wire n4666;
	wire n4668;
	wire n4669;
	wire n4671;
	wire n4672;
	wire n4674;
	wire n4675;
	wire n4677;
	wire n4678;
	wire n4680;
	wire n4681;
	wire n4683;
	wire n4684;
	wire n4686;
	wire n4687;
	wire n4689;
	wire n4690;
	wire n4692;
	wire n4693;
	wire n4695;
	wire n4696;
	wire n4698;
	wire n4699;
	wire n4701;
	wire n4702;
	wire n4704;
	wire n4705;
	wire n4707;
	wire n4708;
	wire n4710;
	wire n4711;
	wire n4713;
	wire n4714;
	wire n4716;
	wire n4717;
	wire n4719;
	wire n4720;
	wire n4722;
	wire n4723;
	wire n4725;
	wire n4726;
	wire n4728;
	wire n4729;
	wire n4731;
	wire n4732;
	wire n4734;
	wire n4735;
	wire n4737;
	wire n4738;
	wire n4740;
	wire n4741;
	wire n4743;
	wire n4744;
	wire n4746;
	wire n4747;
	wire n4749;
	wire n4750;
	wire n4752;
	wire n4753;
	wire n4755;
	wire n4756;
	wire n4758;
	wire n4759;
	wire n4761;
	wire n4762;
	wire n4764;
	wire n4765;
	wire n4767;
	wire n4768;
	wire n4770;
	wire n4771;
	wire n4773;
	wire n4774;
	wire n4776;
	wire n4777;
	wire n4779;
	wire n4780;
	wire n4782;
	wire n4783;
	wire n4785;
	wire n4786;
	wire n4788;
	wire n4789;
	wire n4791;
	wire n4792;
	wire n4794;
	wire n4795;
	wire n4797;
	wire n4798;
	wire n4800;
	wire n4801;
	wire n4803;
	wire n4804;
	wire n4806;
	wire n4807;
	wire n4809;
	wire n4810;
	wire n4812;
	wire n4813;
	wire n4815;
	wire n4816;
	wire n4818;
	wire n4819;
	wire n4821;
	wire n4822;
	wire n4824;
	wire n4825;
	wire n4827;
	wire n4828;
	wire n4830;
	wire n4831;
	wire n4834;
	wire n4835;
	wire [2:0] w_in00_0;
	wire [2:0] w_in01_0;
	wire [1:0] w_in01_1;
	wire [2:0] w_in02_0;
	wire [2:0] w_in03_0;
	wire [2:0] w_in04_0;
	wire [2:0] w_in05_0;
	wire [2:0] w_in06_0;
	wire [2:0] w_in07_0;
	wire [2:0] w_in08_0;
	wire [2:0] w_in09_0;
	wire [2:0] w_in010_0;
	wire [2:0] w_in011_0;
	wire [2:0] w_in012_0;
	wire [2:0] w_in013_0;
	wire [2:0] w_in014_0;
	wire [2:0] w_in015_0;
	wire [2:0] w_in016_0;
	wire [2:0] w_in017_0;
	wire [2:0] w_in018_0;
	wire [2:0] w_in019_0;
	wire [2:0] w_in020_0;
	wire [2:0] w_in021_0;
	wire [2:0] w_in022_0;
	wire [2:0] w_in023_0;
	wire [2:0] w_in024_0;
	wire [2:0] w_in025_0;
	wire [2:0] w_in026_0;
	wire [2:0] w_in027_0;
	wire [2:0] w_in028_0;
	wire [2:0] w_in029_0;
	wire [2:0] w_in030_0;
	wire [2:0] w_in031_0;
	wire [2:0] w_in032_0;
	wire [2:0] w_in033_0;
	wire [2:0] w_in034_0;
	wire [2:0] w_in035_0;
	wire [2:0] w_in036_0;
	wire [2:0] w_in037_0;
	wire [2:0] w_in038_0;
	wire [2:0] w_in039_0;
	wire [2:0] w_in040_0;
	wire [2:0] w_in041_0;
	wire [2:0] w_in042_0;
	wire [2:0] w_in043_0;
	wire [2:0] w_in044_0;
	wire [2:0] w_in045_0;
	wire [2:0] w_in046_0;
	wire [2:0] w_in047_0;
	wire [2:0] w_in048_0;
	wire [2:0] w_in049_0;
	wire [2:0] w_in050_0;
	wire [2:0] w_in051_0;
	wire [2:0] w_in052_0;
	wire [2:0] w_in053_0;
	wire [2:0] w_in054_0;
	wire [2:0] w_in055_0;
	wire [2:0] w_in056_0;
	wire [2:0] w_in057_0;
	wire [2:0] w_in058_0;
	wire [2:0] w_in059_0;
	wire [2:0] w_in060_0;
	wire [2:0] w_in061_0;
	wire [2:0] w_in062_0;
	wire [2:0] w_in063_0;
	wire [2:0] w_in064_0;
	wire [2:0] w_in065_0;
	wire [2:0] w_in066_0;
	wire [2:0] w_in067_0;
	wire [2:0] w_in068_0;
	wire [2:0] w_in069_0;
	wire [2:0] w_in070_0;
	wire [2:0] w_in071_0;
	wire [2:0] w_in072_0;
	wire [2:0] w_in073_0;
	wire [2:0] w_in074_0;
	wire [2:0] w_in075_0;
	wire [2:0] w_in076_0;
	wire [2:0] w_in077_0;
	wire [2:0] w_in078_0;
	wire [2:0] w_in079_0;
	wire [2:0] w_in080_0;
	wire [2:0] w_in081_0;
	wire [2:0] w_in082_0;
	wire [2:0] w_in083_0;
	wire [2:0] w_in084_0;
	wire [2:0] w_in085_0;
	wire [2:0] w_in086_0;
	wire [2:0] w_in087_0;
	wire [2:0] w_in088_0;
	wire [2:0] w_in089_0;
	wire [2:0] w_in090_0;
	wire [2:0] w_in091_0;
	wire [2:0] w_in092_0;
	wire [2:0] w_in093_0;
	wire [2:0] w_in094_0;
	wire [2:0] w_in095_0;
	wire [2:0] w_in096_0;
	wire [2:0] w_in097_0;
	wire [2:0] w_in098_0;
	wire [2:0] w_in099_0;
	wire [2:0] w_in0100_0;
	wire [2:0] w_in0101_0;
	wire [2:0] w_in0102_0;
	wire [2:0] w_in0103_0;
	wire [2:0] w_in0104_0;
	wire [2:0] w_in0105_0;
	wire [2:0] w_in0106_0;
	wire [2:0] w_in0107_0;
	wire [2:0] w_in0108_0;
	wire [2:0] w_in0109_0;
	wire [2:0] w_in0110_0;
	wire [2:0] w_in0111_0;
	wire [2:0] w_in0112_0;
	wire [2:0] w_in0113_0;
	wire [2:0] w_in0114_0;
	wire [2:0] w_in0115_0;
	wire [2:0] w_in0116_0;
	wire [2:0] w_in0117_0;
	wire [2:0] w_in0118_0;
	wire [2:0] w_in0119_0;
	wire [2:0] w_in0120_0;
	wire [2:0] w_in0121_0;
	wire [2:0] w_in0122_0;
	wire [2:0] w_in0123_0;
	wire [2:0] w_in0124_0;
	wire [2:0] w_in0125_0;
	wire [2:0] w_in0126_0;
	wire [2:0] w_in0127_0;
	wire [2:0] w_in10_0;
	wire [2:0] w_in11_0;
	wire [1:0] w_in11_1;
	wire [2:0] w_in12_0;
	wire [2:0] w_in13_0;
	wire [2:0] w_in14_0;
	wire [2:0] w_in15_0;
	wire [2:0] w_in16_0;
	wire [2:0] w_in17_0;
	wire [2:0] w_in18_0;
	wire [2:0] w_in19_0;
	wire [2:0] w_in110_0;
	wire [2:0] w_in111_0;
	wire [2:0] w_in112_0;
	wire [2:0] w_in113_0;
	wire [2:0] w_in114_0;
	wire [2:0] w_in115_0;
	wire [2:0] w_in116_0;
	wire [2:0] w_in117_0;
	wire [2:0] w_in118_0;
	wire [2:0] w_in119_0;
	wire [2:0] w_in120_0;
	wire [2:0] w_in121_0;
	wire [2:0] w_in122_0;
	wire [2:0] w_in123_0;
	wire [2:0] w_in124_0;
	wire [2:0] w_in125_0;
	wire [2:0] w_in126_0;
	wire [2:0] w_in127_0;
	wire [2:0] w_in128_0;
	wire [2:0] w_in129_0;
	wire [2:0] w_in130_0;
	wire [2:0] w_in131_0;
	wire [2:0] w_in132_0;
	wire [2:0] w_in133_0;
	wire [2:0] w_in134_0;
	wire [2:0] w_in135_0;
	wire [2:0] w_in136_0;
	wire [2:0] w_in137_0;
	wire [2:0] w_in138_0;
	wire [2:0] w_in139_0;
	wire [2:0] w_in140_0;
	wire [2:0] w_in141_0;
	wire [2:0] w_in142_0;
	wire [2:0] w_in143_0;
	wire [2:0] w_in144_0;
	wire [2:0] w_in145_0;
	wire [2:0] w_in146_0;
	wire [2:0] w_in147_0;
	wire [2:0] w_in148_0;
	wire [2:0] w_in149_0;
	wire [2:0] w_in150_0;
	wire [2:0] w_in151_0;
	wire [1:0] w_in152_0;
	wire [2:0] w_in153_0;
	wire [2:0] w_in154_0;
	wire [2:0] w_in155_0;
	wire [2:0] w_in156_0;
	wire [2:0] w_in157_0;
	wire [2:0] w_in158_0;
	wire [2:0] w_in159_0;
	wire [2:0] w_in160_0;
	wire [2:0] w_in161_0;
	wire [2:0] w_in162_0;
	wire [2:0] w_in163_0;
	wire [2:0] w_in164_0;
	wire [2:0] w_in165_0;
	wire [2:0] w_in166_0;
	wire [2:0] w_in167_0;
	wire [2:0] w_in168_0;
	wire [2:0] w_in169_0;
	wire [2:0] w_in170_0;
	wire [2:0] w_in171_0;
	wire [2:0] w_in172_0;
	wire [2:0] w_in173_0;
	wire [2:0] w_in174_0;
	wire [2:0] w_in175_0;
	wire [2:0] w_in176_0;
	wire [2:0] w_in177_0;
	wire [2:0] w_in178_0;
	wire [2:0] w_in179_0;
	wire [2:0] w_in180_0;
	wire [2:0] w_in181_0;
	wire [2:0] w_in182_0;
	wire [2:0] w_in183_0;
	wire [2:0] w_in184_0;
	wire [2:0] w_in185_0;
	wire [2:0] w_in186_0;
	wire [2:0] w_in187_0;
	wire [2:0] w_in188_0;
	wire [2:0] w_in189_0;
	wire [2:0] w_in190_0;
	wire [2:0] w_in191_0;
	wire [2:0] w_in192_0;
	wire [2:0] w_in193_0;
	wire [2:0] w_in194_0;
	wire [2:0] w_in195_0;
	wire [2:0] w_in196_0;
	wire [2:0] w_in197_0;
	wire [2:0] w_in198_0;
	wire [2:0] w_in199_0;
	wire [2:0] w_in1100_0;
	wire [2:0] w_in1101_0;
	wire [2:0] w_in1102_0;
	wire [2:0] w_in1103_0;
	wire [2:0] w_in1104_0;
	wire [2:0] w_in1105_0;
	wire [2:0] w_in1106_0;
	wire [2:0] w_in1107_0;
	wire [2:0] w_in1108_0;
	wire [2:0] w_in1109_0;
	wire [2:0] w_in1110_0;
	wire [2:0] w_in1111_0;
	wire [2:0] w_in1112_0;
	wire [2:0] w_in1113_0;
	wire [2:0] w_in1114_0;
	wire [2:0] w_in1115_0;
	wire [2:0] w_in1116_0;
	wire [2:0] w_in1117_0;
	wire [2:0] w_in1118_0;
	wire [2:0] w_in1119_0;
	wire [2:0] w_in1120_0;
	wire [2:0] w_in1121_0;
	wire [2:0] w_in1122_0;
	wire [2:0] w_in1123_0;
	wire [2:0] w_in1124_0;
	wire [2:0] w_in1125_0;
	wire [2:0] w_in1126_0;
	wire [2:0] w_in1127_0;
	wire [2:0] w_in20_0;
	wire [2:0] w_in21_0;
	wire [1:0] w_in21_1;
	wire [2:0] w_in22_0;
	wire [2:0] w_in23_0;
	wire [2:0] w_in24_0;
	wire [2:0] w_in25_0;
	wire [2:0] w_in26_0;
	wire [2:0] w_in27_0;
	wire [2:0] w_in28_0;
	wire [2:0] w_in29_0;
	wire [2:0] w_in210_0;
	wire [2:0] w_in211_0;
	wire [2:0] w_in212_0;
	wire [2:0] w_in213_0;
	wire [2:0] w_in214_0;
	wire [2:0] w_in215_0;
	wire [2:0] w_in216_0;
	wire [2:0] w_in217_0;
	wire [2:0] w_in218_0;
	wire [2:0] w_in219_0;
	wire [2:0] w_in220_0;
	wire [2:0] w_in221_0;
	wire [2:0] w_in222_0;
	wire [2:0] w_in223_0;
	wire [2:0] w_in224_0;
	wire [2:0] w_in225_0;
	wire [2:0] w_in226_0;
	wire [2:0] w_in227_0;
	wire [2:0] w_in228_0;
	wire [2:0] w_in229_0;
	wire [2:0] w_in230_0;
	wire [2:0] w_in231_0;
	wire [2:0] w_in232_0;
	wire [2:0] w_in233_0;
	wire [2:0] w_in234_0;
	wire [2:0] w_in235_0;
	wire [2:0] w_in236_0;
	wire [2:0] w_in237_0;
	wire [2:0] w_in238_0;
	wire [2:0] w_in239_0;
	wire [2:0] w_in240_0;
	wire [2:0] w_in241_0;
	wire [2:0] w_in242_0;
	wire [2:0] w_in243_0;
	wire [2:0] w_in244_0;
	wire [2:0] w_in245_0;
	wire [2:0] w_in246_0;
	wire [2:0] w_in247_0;
	wire [2:0] w_in248_0;
	wire [2:0] w_in249_0;
	wire [2:0] w_in250_0;
	wire [2:0] w_in251_0;
	wire [2:0] w_in252_0;
	wire [2:0] w_in253_0;
	wire [2:0] w_in254_0;
	wire [2:0] w_in255_0;
	wire [2:0] w_in256_0;
	wire [2:0] w_in257_0;
	wire [2:0] w_in258_0;
	wire [2:0] w_in259_0;
	wire [2:0] w_in260_0;
	wire [2:0] w_in261_0;
	wire [2:0] w_in262_0;
	wire [2:0] w_in263_0;
	wire [2:0] w_in264_0;
	wire [2:0] w_in265_0;
	wire [2:0] w_in266_0;
	wire [2:0] w_in267_0;
	wire [2:0] w_in268_0;
	wire [2:0] w_in269_0;
	wire [2:0] w_in270_0;
	wire [2:0] w_in271_0;
	wire [2:0] w_in272_0;
	wire [2:0] w_in273_0;
	wire [2:0] w_in274_0;
	wire [2:0] w_in275_0;
	wire [2:0] w_in276_0;
	wire [2:0] w_in277_0;
	wire [2:0] w_in278_0;
	wire [2:0] w_in279_0;
	wire [2:0] w_in280_0;
	wire [2:0] w_in281_0;
	wire [2:0] w_in282_0;
	wire [2:0] w_in283_0;
	wire [2:0] w_in284_0;
	wire [2:0] w_in285_0;
	wire [2:0] w_in286_0;
	wire [2:0] w_in287_0;
	wire [2:0] w_in288_0;
	wire [2:0] w_in289_0;
	wire [2:0] w_in290_0;
	wire [2:0] w_in291_0;
	wire [2:0] w_in292_0;
	wire [2:0] w_in293_0;
	wire [2:0] w_in294_0;
	wire [2:0] w_in295_0;
	wire [2:0] w_in296_0;
	wire [2:0] w_in297_0;
	wire [2:0] w_in298_0;
	wire [2:0] w_in299_0;
	wire [2:0] w_in2100_0;
	wire [2:0] w_in2101_0;
	wire [2:0] w_in2102_0;
	wire [2:0] w_in2103_0;
	wire [2:0] w_in2104_0;
	wire [2:0] w_in2105_0;
	wire [2:0] w_in2106_0;
	wire [2:0] w_in2107_0;
	wire [2:0] w_in2108_0;
	wire [2:0] w_in2109_0;
	wire [2:0] w_in2110_0;
	wire [2:0] w_in2111_0;
	wire [2:0] w_in2112_0;
	wire [2:0] w_in2113_0;
	wire [2:0] w_in2114_0;
	wire [2:0] w_in2115_0;
	wire [2:0] w_in2116_0;
	wire [2:0] w_in2117_0;
	wire [2:0] w_in2118_0;
	wire [2:0] w_in2119_0;
	wire [2:0] w_in2120_0;
	wire [2:0] w_in2121_0;
	wire [2:0] w_in2122_0;
	wire [2:0] w_in2123_0;
	wire [2:0] w_in2124_0;
	wire [2:0] w_in2125_0;
	wire [2:0] w_in2126_0;
	wire [2:0] w_in2127_0;
	wire [2:0] w_in30_0;
	wire [2:0] w_in31_0;
	wire [1:0] w_in31_1;
	wire [2:0] w_in32_0;
	wire [2:0] w_in33_0;
	wire [2:0] w_in34_0;
	wire [2:0] w_in35_0;
	wire [2:0] w_in36_0;
	wire [2:0] w_in37_0;
	wire [2:0] w_in38_0;
	wire [2:0] w_in39_0;
	wire [2:0] w_in310_0;
	wire [2:0] w_in311_0;
	wire [2:0] w_in312_0;
	wire [2:0] w_in313_0;
	wire [2:0] w_in314_0;
	wire [2:0] w_in315_0;
	wire [2:0] w_in316_0;
	wire [2:0] w_in317_0;
	wire [2:0] w_in318_0;
	wire [2:0] w_in319_0;
	wire [2:0] w_in320_0;
	wire [2:0] w_in321_0;
	wire [2:0] w_in322_0;
	wire [2:0] w_in323_0;
	wire [2:0] w_in324_0;
	wire [2:0] w_in325_0;
	wire [2:0] w_in326_0;
	wire [2:0] w_in327_0;
	wire [2:0] w_in328_0;
	wire [2:0] w_in329_0;
	wire [2:0] w_in330_0;
	wire [2:0] w_in331_0;
	wire [2:0] w_in332_0;
	wire [2:0] w_in333_0;
	wire [2:0] w_in334_0;
	wire [2:0] w_in335_0;
	wire [2:0] w_in336_0;
	wire [2:0] w_in337_0;
	wire [2:0] w_in338_0;
	wire [2:0] w_in339_0;
	wire [2:0] w_in340_0;
	wire [2:0] w_in341_0;
	wire [2:0] w_in342_0;
	wire [2:0] w_in343_0;
	wire [2:0] w_in344_0;
	wire [2:0] w_in345_0;
	wire [2:0] w_in346_0;
	wire [2:0] w_in347_0;
	wire [2:0] w_in348_0;
	wire [2:0] w_in349_0;
	wire [2:0] w_in350_0;
	wire [2:0] w_in351_0;
	wire [1:0] w_in352_0;
	wire [2:0] w_in353_0;
	wire [2:0] w_in354_0;
	wire [2:0] w_in355_0;
	wire [2:0] w_in356_0;
	wire [2:0] w_in357_0;
	wire [2:0] w_in358_0;
	wire [2:0] w_in359_0;
	wire [2:0] w_in360_0;
	wire [2:0] w_in361_0;
	wire [2:0] w_in362_0;
	wire [2:0] w_in363_0;
	wire [2:0] w_in364_0;
	wire [2:0] w_in365_0;
	wire [2:0] w_in366_0;
	wire [2:0] w_in367_0;
	wire [2:0] w_in368_0;
	wire [2:0] w_in369_0;
	wire [2:0] w_in370_0;
	wire [2:0] w_in371_0;
	wire [2:0] w_in372_0;
	wire [2:0] w_in373_0;
	wire [2:0] w_in374_0;
	wire [2:0] w_in375_0;
	wire [2:0] w_in376_0;
	wire [2:0] w_in377_0;
	wire [2:0] w_in378_0;
	wire [2:0] w_in379_0;
	wire [2:0] w_in380_0;
	wire [2:0] w_in381_0;
	wire [2:0] w_in382_0;
	wire [2:0] w_in383_0;
	wire [2:0] w_in384_0;
	wire [2:0] w_in385_0;
	wire [2:0] w_in386_0;
	wire [2:0] w_in387_0;
	wire [2:0] w_in388_0;
	wire [2:0] w_in389_0;
	wire [2:0] w_in390_0;
	wire [2:0] w_in391_0;
	wire [2:0] w_in392_0;
	wire [2:0] w_in393_0;
	wire [2:0] w_in394_0;
	wire [2:0] w_in395_0;
	wire [2:0] w_in396_0;
	wire [2:0] w_in397_0;
	wire [2:0] w_in398_0;
	wire [2:0] w_in399_0;
	wire [2:0] w_in3100_0;
	wire [2:0] w_in3101_0;
	wire [2:0] w_in3102_0;
	wire [2:0] w_in3103_0;
	wire [2:0] w_in3104_0;
	wire [2:0] w_in3105_0;
	wire [2:0] w_in3106_0;
	wire [2:0] w_in3107_0;
	wire [2:0] w_in3108_0;
	wire [2:0] w_in3109_0;
	wire [2:0] w_in3110_0;
	wire [2:0] w_in3111_0;
	wire [2:0] w_in3112_0;
	wire [2:0] w_in3113_0;
	wire [2:0] w_in3114_0;
	wire [2:0] w_in3115_0;
	wire [2:0] w_in3116_0;
	wire [2:0] w_in3117_0;
	wire [2:0] w_in3118_0;
	wire [2:0] w_in3119_0;
	wire [2:0] w_in3120_0;
	wire [2:0] w_in3121_0;
	wire [2:0] w_in3122_0;
	wire [2:0] w_in3123_0;
	wire [2:0] w_in3124_0;
	wire [2:0] w_in3125_0;
	wire [2:0] w_in3126_0;
	wire [2:0] w_in3127_0;
	wire [2:0] w_address1_0;
	wire [2:0] w_address1_1;
	wire [2:0] w_address1_2;
	wire [2:0] w_address1_3;
	wire [2:0] w_address1_4;
	wire [2:0] w_address1_5;
	wire [2:0] w_address1_6;
	wire [2:0] w_address1_7;
	wire [2:0] w_address1_8;
	wire [2:0] w_address1_9;
	wire [2:0] w_address1_10;
	wire [2:0] w_address1_11;
	wire [2:0] w_address1_12;
	wire [2:0] w_address1_13;
	wire [2:0] w_address1_14;
	wire [2:0] w_address1_15;
	wire [2:0] w_address1_16;
	wire [2:0] w_address1_17;
	wire [2:0] w_address1_18;
	wire [2:0] w_address1_19;
	wire [2:0] w_address1_20;
	wire [2:0] w_address1_21;
	wire [2:0] w_address1_22;
	wire [2:0] w_address1_23;
	wire [2:0] w_address1_24;
	wire [2:0] w_address1_25;
	wire [2:0] w_address1_26;
	wire [2:0] w_address1_27;
	wire [2:0] w_address1_28;
	wire [2:0] w_address1_29;
	wire [2:0] w_address1_30;
	wire [2:0] w_address1_31;
	wire [2:0] w_address1_32;
	wire [2:0] w_address1_33;
	wire [2:0] w_address1_34;
	wire [2:0] w_address1_35;
	wire [2:0] w_address1_36;
	wire [2:0] w_address1_37;
	wire [2:0] w_address1_38;
	wire [2:0] w_address1_39;
	wire [2:0] w_address1_40;
	wire [2:0] w_address1_41;
	wire [2:0] w_address1_42;
	wire [2:0] w_address1_43;
	wire [2:0] w_address1_44;
	wire [2:0] w_address1_45;
	wire [2:0] w_address1_46;
	wire [2:0] w_address1_47;
	wire [2:0] w_address1_48;
	wire [2:0] w_address1_49;
	wire [2:0] w_address1_50;
	wire [2:0] w_address1_51;
	wire [2:0] w_address1_52;
	wire [2:0] w_address1_53;
	wire [2:0] w_address1_54;
	wire [2:0] w_address1_55;
	wire [2:0] w_address1_56;
	wire [2:0] w_address1_57;
	wire [2:0] w_address1_58;
	wire [2:0] w_address1_59;
	wire [2:0] w_address1_60;
	wire [2:0] w_address1_61;
	wire [2:0] w_address1_62;
	wire [1:0] w_address1_63;
	wire address_fa_1;
	wire [1:0] w_n643_0;
	wire [1:0] w_n646_0;
	wire [1:0] w_n648_0;
	wire [1:0] w_n651_0;
	wire [1:0] w_n653_0;
	wire [1:0] w_n656_0;
	wire [1:0] w_n658_0;
	wire [1:0] w_n661_0;
	wire [1:0] w_n663_0;
	wire [1:0] w_n666_0;
	wire [1:0] w_n668_0;
	wire [1:0] w_n671_0;
	wire [1:0] w_n673_0;
	wire [1:0] w_n676_0;
	wire [1:0] w_n678_0;
	wire [1:0] w_n681_0;
	wire [1:0] w_n683_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n688_0;
	wire [1:0] w_n691_0;
	wire [1:0] w_n693_0;
	wire [1:0] w_n696_0;
	wire [1:0] w_n698_0;
	wire [1:0] w_n701_0;
	wire [1:0] w_n703_0;
	wire [1:0] w_n706_0;
	wire [1:0] w_n708_0;
	wire [1:0] w_n711_0;
	wire [1:0] w_n713_0;
	wire [1:0] w_n716_0;
	wire [1:0] w_n718_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n726_0;
	wire [1:0] w_n728_0;
	wire [1:0] w_n731_0;
	wire [1:0] w_n733_0;
	wire [1:0] w_n736_0;
	wire [1:0] w_n738_0;
	wire [1:0] w_n741_0;
	wire [1:0] w_n743_0;
	wire [1:0] w_n746_0;
	wire [1:0] w_n748_0;
	wire [1:0] w_n751_0;
	wire [1:0] w_n753_0;
	wire [1:0] w_n756_0;
	wire [1:0] w_n758_0;
	wire [1:0] w_n761_0;
	wire [1:0] w_n763_0;
	wire [1:0] w_n766_0;
	wire [1:0] w_n768_0;
	wire [1:0] w_n771_0;
	wire [1:0] w_n773_0;
	wire [1:0] w_n776_0;
	wire [1:0] w_n778_0;
	wire [1:0] w_n780_0;
	wire [1:0] w_n781_0;
	wire [1:0] w_n782_0;
	wire [1:0] w_n783_0;
	wire [1:0] w_n785_0;
	wire [1:0] w_n788_0;
	wire [1:0] w_n853_0;
	wire [1:0] w_n858_0;
	wire [1:0] w_n862_0;
	wire [1:0] w_n867_0;
	wire [1:0] w_n871_0;
	wire [1:0] w_n874_0;
	wire [1:0] w_n880_0;
	wire [1:0] w_n915_0;
	wire [1:0] w_n920_0;
	wire [1:0] w_n924_0;
	wire [1:0] w_n929_0;
	wire [1:0] w_n931_0;
	wire [1:0] w_n935_0;
	wire [1:0] w_n939_0;
	wire [1:0] w_n974_0;
	wire [1:0] w_n979_0;
	wire [1:0] w_n980_0;
	wire [1:0] w_n982_0;
	wire [1:0] w_n988_0;
	wire [1:0] w_n993_0;
	wire [1:0] w_n997_0;
	wire [1:0] w_n1001_0;
	wire [1:0] w_n1032_0;
	wire [1:0] w_n1037_0;
	wire [1:0] w_n1041_0;
	wire [1:0] w_n1046_0;
	wire [1:0] w_n1048_0;
	wire [1:0] w_n1052_0;
	wire [1:0] w_n1056_0;
	wire [1:0] w_n1091_0;
	wire [1:0] w_n1097_0;
	wire [1:0] w_n1099_0;
	wire [1:0] w_n1103_0;
	wire [1:0] w_n1120_0;
	wire [1:0] w_n1127_0;
	wire [1:0] w_n1131_0;
	wire [1:0] w_n1132_0;
	wire [1:0] w_n1149_0;
	wire [1:0] w_n1155_0;
	wire [1:0] w_n1157_0;
	wire [1:0] w_n1161_0;
	wire [1:0] w_n1178_0;
	wire [1:0] w_n1185_0;
	wire [1:0] w_n1189_0;
	wire [1:0] w_n1190_0;
	wire [1:0] w_n1207_0;
	wire [1:0] w_n1213_0;
	wire [1:0] w_n1215_0;
	wire [1:0] w_n1219_0;
	wire [1:0] w_n1236_0;
	wire [1:0] w_n1243_0;
	wire [1:0] w_n1247_0;
	wire [1:0] w_n1248_0;
	wire [1:0] w_n1265_0;
	wire [1:0] w_n1271_0;
	wire [1:0] w_n1273_0;
	wire [1:0] w_n1277_0;
	wire [1:0] w_n1294_0;
	wire [1:0] w_n1301_0;
	wire [1:0] w_n1305_0;
	wire [1:0] w_n1306_0;
	wire [1:0] w_n1323_0;
	wire [1:0] w_n1329_0;
	wire [1:0] w_n1331_0;
	wire [1:0] w_n1335_0;
	wire [1:0] w_n1352_0;
	wire [1:0] w_n1359_0;
	wire [1:0] w_n1363_0;
	wire [1:0] w_n1364_0;
	wire [1:0] w_n1381_0;
	wire [1:0] w_n1387_0;
	wire [1:0] w_n1389_0;
	wire [1:0] w_n1393_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1417_0;
	wire [1:0] w_n1421_0;
	wire [1:0] w_n1422_0;
	wire [1:0] w_n1439_0;
	wire [1:0] w_n1445_0;
	wire [1:0] w_n1447_0;
	wire [1:0] w_n1451_0;
	wire [1:0] w_n1468_0;
	wire [1:0] w_n1475_0;
	wire [1:0] w_n1479_0;
	wire [1:0] w_n1480_0;
	wire [1:0] w_n1497_0;
	wire [1:0] w_n1503_0;
	wire [1:0] w_n1505_0;
	wire [1:0] w_n1509_0;
	wire [1:0] w_n1526_0;
	wire [1:0] w_n1532_0;
	wire [1:0] w_n1534_0;
	wire [1:0] w_n1538_0;
	wire [1:0] w_n1555_0;
	wire [2:0] w_n1556_0;
	wire [2:0] w_n1556_1;
	wire [2:0] w_n1556_2;
	wire [2:0] w_n1556_3;
	wire [2:0] w_n1556_4;
	wire [2:0] w_n1556_5;
	wire [2:0] w_n1556_6;
	wire [2:0] w_n1556_7;
	wire [2:0] w_n1556_8;
	wire [2:0] w_n1556_9;
	wire [2:0] w_n1556_10;
	wire [2:0] w_n1556_11;
	wire [2:0] w_n1556_12;
	wire [2:0] w_n1556_13;
	wire [2:0] w_n1556_14;
	wire [2:0] w_n1556_15;
	wire [2:0] w_n1556_16;
	wire [2:0] w_n1556_17;
	wire [2:0] w_n1556_18;
	wire [2:0] w_n1556_19;
	wire [2:0] w_n1556_20;
	wire [2:0] w_n1556_21;
	wire [2:0] w_n1556_22;
	wire [2:0] w_n1556_23;
	wire [2:0] w_n1556_24;
	wire [2:0] w_n1556_25;
	wire [2:0] w_n1556_26;
	wire [2:0] w_n1556_27;
	wire [2:0] w_n1556_28;
	wire [2:0] w_n1556_29;
	wire [2:0] w_n1556_30;
	wire [2:0] w_n1556_31;
	wire [2:0] w_n1556_32;
	wire [2:0] w_n1556_33;
	wire [2:0] w_n1556_34;
	wire [2:0] w_n1556_35;
	wire [2:0] w_n1556_36;
	wire [2:0] w_n1556_37;
	wire [2:0] w_n1556_38;
	wire [2:0] w_n1556_39;
	wire [2:0] w_n1556_40;
	wire [2:0] w_n1556_41;
	wire [2:0] w_n1556_42;
	wire [2:0] w_n1556_43;
	wire [2:0] w_n1556_44;
	wire [2:0] w_n1556_45;
	wire [2:0] w_n1556_46;
	wire [2:0] w_n1556_47;
	wire [2:0] w_n1556_48;
	wire [2:0] w_n1556_49;
	wire [2:0] w_n1556_50;
	wire [2:0] w_n1556_51;
	wire [2:0] w_n1556_52;
	wire [2:0] w_n1556_53;
	wire [2:0] w_n1556_54;
	wire [2:0] w_n1556_55;
	wire [2:0] w_n1556_56;
	wire [2:0] w_n1556_57;
	wire [2:0] w_n1556_58;
	wire [2:0] w_n1556_59;
	wire [2:0] w_n1556_60;
	wire [2:0] w_n1556_61;
	wire [2:0] w_n1556_62;
	wire [2:0] w_n1556_63;
	wire [1:0] w_n1586_0;
	wire [1:0] w_n1589_0;
	wire [2:0] w_n1711_0;
	wire [2:0] w_n1711_1;
	wire [2:0] w_n1711_2;
	wire [2:0] w_n1711_3;
	wire [2:0] w_n1711_4;
	wire [2:0] w_n1711_5;
	wire [2:0] w_n1711_6;
	wire [2:0] w_n1711_7;
	wire [2:0] w_n1711_8;
	wire [2:0] w_n1711_9;
	wire [2:0] w_n1711_10;
	wire [2:0] w_n1711_11;
	wire [2:0] w_n1711_12;
	wire [2:0] w_n1711_13;
	wire [2:0] w_n1711_14;
	wire [2:0] w_n1711_15;
	wire [2:0] w_n1711_16;
	wire [2:0] w_n1711_17;
	wire [2:0] w_n1711_18;
	wire [2:0] w_n1711_19;
	wire [2:0] w_n1711_20;
	wire [2:0] w_n1711_21;
	wire [2:0] w_n1711_22;
	wire [2:0] w_n1711_23;
	wire [2:0] w_n1711_24;
	wire [2:0] w_n1711_25;
	wire [2:0] w_n1711_26;
	wire [2:0] w_n1711_27;
	wire [2:0] w_n1711_28;
	wire [2:0] w_n1711_29;
	wire [2:0] w_n1711_30;
	wire [2:0] w_n1711_31;
	wire [2:0] w_n1711_32;
	wire [2:0] w_n1711_33;
	wire [2:0] w_n1711_34;
	wire [2:0] w_n1711_35;
	wire [2:0] w_n1711_36;
	wire [2:0] w_n1711_37;
	wire [2:0] w_n1711_38;
	wire [2:0] w_n1711_39;
	wire [2:0] w_n1711_40;
	wire [2:0] w_n1711_41;
	wire [2:0] w_n1711_42;
	wire [2:0] w_n1711_43;
	wire [2:0] w_n1711_44;
	wire [2:0] w_n1711_45;
	wire [2:0] w_n1711_46;
	wire [2:0] w_n1711_47;
	wire [2:0] w_n1711_48;
	wire [2:0] w_n1711_49;
	wire [2:0] w_n1711_50;
	wire [2:0] w_n1711_51;
	wire [2:0] w_n1711_52;
	wire [2:0] w_n1711_53;
	wire [2:0] w_n1711_54;
	wire [2:0] w_n1711_55;
	wire [2:0] w_n1711_56;
	wire [2:0] w_n1711_57;
	wire [2:0] w_n1711_58;
	wire [2:0] w_n1711_59;
	wire [2:0] w_n1711_60;
	wire [2:0] w_n1711_61;
	wire [2:0] w_n1711_62;
	wire [2:0] w_n1711_63;
	wire [1:0] w_n1711_64;
	wire [1:0] w_n1713_0;
	wire [1:0] w_n1715_0;
	wire [1:0] w_n1718_0;
	wire [1:0] w_n1720_0;
	wire [1:0] w_n1723_0;
	wire [1:0] w_n1725_0;
	wire [1:0] w_n1728_0;
	wire [1:0] w_n1730_0;
	wire [1:0] w_n1733_0;
	wire [1:0] w_n1735_0;
	wire [1:0] w_n1738_0;
	wire [1:0] w_n1740_0;
	wire [1:0] w_n1743_0;
	wire [1:0] w_n1745_0;
	wire [1:0] w_n1748_0;
	wire [1:0] w_n1750_0;
	wire [1:0] w_n1753_0;
	wire [1:0] w_n1755_0;
	wire [1:0] w_n1758_0;
	wire [1:0] w_n1760_0;
	wire [1:0] w_n1763_0;
	wire [1:0] w_n1765_0;
	wire [1:0] w_n1768_0;
	wire [1:0] w_n1770_0;
	wire [1:0] w_n1773_0;
	wire [1:0] w_n1775_0;
	wire [1:0] w_n1778_0;
	wire [1:0] w_n1780_0;
	wire [1:0] w_n1783_0;
	wire [1:0] w_n1785_0;
	wire [1:0] w_n1788_0;
	wire [1:0] w_n1790_0;
	wire [1:0] w_n1793_0;
	wire [1:0] w_n1795_0;
	wire [1:0] w_n1798_0;
	wire [1:0] w_n1800_0;
	wire [1:0] w_n1803_0;
	wire [1:0] w_n1805_0;
	wire [1:0] w_n1808_0;
	wire [1:0] w_n1810_0;
	wire [1:0] w_n1813_0;
	wire [1:0] w_n1815_0;
	wire [1:0] w_n1818_0;
	wire [1:0] w_n1820_0;
	wire [1:0] w_n1823_0;
	wire [1:0] w_n1825_0;
	wire [1:0] w_n1828_0;
	wire [1:0] w_n1830_0;
	wire [1:0] w_n1833_0;
	wire [1:0] w_n1835_0;
	wire [1:0] w_n1838_0;
	wire [1:0] w_n1840_0;
	wire [1:0] w_n1843_0;
	wire [1:0] w_n1845_0;
	wire [1:0] w_n1848_0;
	wire [1:0] w_n1850_0;
	wire [1:0] w_n1852_0;
	wire [1:0] w_n1853_0;
	wire [1:0] w_n1854_0;
	wire [1:0] w_n1855_0;
	wire [2:0] w_n1857_0;
	wire [1:0] w_n1860_0;
	wire [1:0] w_n1925_0;
	wire [1:0] w_n1930_0;
	wire [1:0] w_n1934_0;
	wire [1:0] w_n1939_0;
	wire [1:0] w_n1943_0;
	wire [1:0] w_n1946_0;
	wire [1:0] w_n1952_0;
	wire [1:0] w_n1987_0;
	wire [1:0] w_n1992_0;
	wire [1:0] w_n1996_0;
	wire [1:0] w_n2001_0;
	wire [1:0] w_n2003_0;
	wire [1:0] w_n2007_0;
	wire [1:0] w_n2011_0;
	wire [1:0] w_n2046_0;
	wire [1:0] w_n2051_0;
	wire [1:0] w_n2052_0;
	wire [1:0] w_n2054_0;
	wire [1:0] w_n2060_0;
	wire [1:0] w_n2065_0;
	wire [1:0] w_n2069_0;
	wire [1:0] w_n2073_0;
	wire [1:0] w_n2104_0;
	wire [1:0] w_n2109_0;
	wire [1:0] w_n2113_0;
	wire [1:0] w_n2118_0;
	wire [1:0] w_n2120_0;
	wire [1:0] w_n2124_0;
	wire [1:0] w_n2128_0;
	wire [1:0] w_n2163_0;
	wire [1:0] w_n2169_0;
	wire [1:0] w_n2171_0;
	wire [1:0] w_n2175_0;
	wire [1:0] w_n2192_0;
	wire [1:0] w_n2199_0;
	wire [1:0] w_n2203_0;
	wire [1:0] w_n2204_0;
	wire [1:0] w_n2221_0;
	wire [1:0] w_n2227_0;
	wire [1:0] w_n2229_0;
	wire [1:0] w_n2233_0;
	wire [1:0] w_n2250_0;
	wire [1:0] w_n2257_0;
	wire [1:0] w_n2261_0;
	wire [1:0] w_n2262_0;
	wire [1:0] w_n2279_0;
	wire [1:0] w_n2285_0;
	wire [1:0] w_n2287_0;
	wire [1:0] w_n2291_0;
	wire [1:0] w_n2308_0;
	wire [1:0] w_n2315_0;
	wire [1:0] w_n2319_0;
	wire [1:0] w_n2320_0;
	wire [1:0] w_n2337_0;
	wire [1:0] w_n2343_0;
	wire [1:0] w_n2345_0;
	wire [1:0] w_n2349_0;
	wire [1:0] w_n2366_0;
	wire [1:0] w_n2373_0;
	wire [1:0] w_n2377_0;
	wire [1:0] w_n2378_0;
	wire [1:0] w_n2395_0;
	wire [1:0] w_n2401_0;
	wire [1:0] w_n2403_0;
	wire [1:0] w_n2407_0;
	wire [1:0] w_n2424_0;
	wire [1:0] w_n2431_0;
	wire [1:0] w_n2435_0;
	wire [1:0] w_n2436_0;
	wire [1:0] w_n2453_0;
	wire [1:0] w_n2459_0;
	wire [1:0] w_n2461_0;
	wire [1:0] w_n2465_0;
	wire [1:0] w_n2482_0;
	wire [1:0] w_n2489_0;
	wire [1:0] w_n2493_0;
	wire [1:0] w_n2494_0;
	wire [1:0] w_n2511_0;
	wire [1:0] w_n2517_0;
	wire [1:0] w_n2519_0;
	wire [1:0] w_n2523_0;
	wire [1:0] w_n2540_0;
	wire [1:0] w_n2547_0;
	wire [1:0] w_n2551_0;
	wire [1:0] w_n2552_0;
	wire [1:0] w_n2569_0;
	wire [1:0] w_n2575_0;
	wire [1:0] w_n2577_0;
	wire [1:0] w_n2581_0;
	wire [1:0] w_n2598_0;
	wire [1:0] w_n2604_0;
	wire [1:0] w_n2606_0;
	wire [1:0] w_n2610_0;
	wire [1:0] w_n2627_0;
	wire [2:0] w_n2628_0;
	wire [2:0] w_n2628_1;
	wire [2:0] w_n2628_2;
	wire [2:0] w_n2628_3;
	wire [2:0] w_n2628_4;
	wire [2:0] w_n2628_5;
	wire [2:0] w_n2628_6;
	wire [2:0] w_n2628_7;
	wire [2:0] w_n2628_8;
	wire [2:0] w_n2628_9;
	wire [2:0] w_n2628_10;
	wire [2:0] w_n2628_11;
	wire [2:0] w_n2628_12;
	wire [2:0] w_n2628_13;
	wire [2:0] w_n2628_14;
	wire [2:0] w_n2628_15;
	wire [2:0] w_n2628_16;
	wire [2:0] w_n2628_17;
	wire [2:0] w_n2628_18;
	wire [2:0] w_n2628_19;
	wire [2:0] w_n2628_20;
	wire [2:0] w_n2628_21;
	wire [2:0] w_n2628_22;
	wire [2:0] w_n2628_23;
	wire [2:0] w_n2628_24;
	wire [2:0] w_n2628_25;
	wire [2:0] w_n2628_26;
	wire [2:0] w_n2628_27;
	wire [2:0] w_n2628_28;
	wire [2:0] w_n2628_29;
	wire [2:0] w_n2628_30;
	wire [2:0] w_n2628_31;
	wire [2:0] w_n2628_32;
	wire [2:0] w_n2628_33;
	wire [2:0] w_n2628_34;
	wire [2:0] w_n2628_35;
	wire [2:0] w_n2628_36;
	wire [2:0] w_n2628_37;
	wire [2:0] w_n2628_38;
	wire [2:0] w_n2628_39;
	wire [2:0] w_n2628_40;
	wire [2:0] w_n2628_41;
	wire [2:0] w_n2628_42;
	wire [2:0] w_n2628_43;
	wire [2:0] w_n2628_44;
	wire [2:0] w_n2628_45;
	wire [2:0] w_n2628_46;
	wire [2:0] w_n2628_47;
	wire [2:0] w_n2628_48;
	wire [2:0] w_n2628_49;
	wire [2:0] w_n2628_50;
	wire [2:0] w_n2628_51;
	wire [2:0] w_n2628_52;
	wire [2:0] w_n2628_53;
	wire [2:0] w_n2628_54;
	wire [2:0] w_n2628_55;
	wire [2:0] w_n2628_56;
	wire [2:0] w_n2628_57;
	wire [2:0] w_n2628_58;
	wire [2:0] w_n2628_59;
	wire [2:0] w_n2628_60;
	wire [2:0] w_n2628_61;
	wire [2:0] w_n2628_62;
	wire [2:0] w_n2628_63;
	wire [1:0] w_n2628_64;
	wire [2:0] w_n2658_0;
	wire [1:0] w_n2661_0;
	wire [2:0] w_n2783_0;
	wire [2:0] w_n2783_1;
	wire [2:0] w_n2783_2;
	wire [2:0] w_n2783_3;
	wire [2:0] w_n2783_4;
	wire [2:0] w_n2783_5;
	wire [2:0] w_n2783_6;
	wire [2:0] w_n2783_7;
	wire [2:0] w_n2783_8;
	wire [2:0] w_n2783_9;
	wire [2:0] w_n2783_10;
	wire [2:0] w_n2783_11;
	wire [2:0] w_n2783_12;
	wire [2:0] w_n2783_13;
	wire [2:0] w_n2783_14;
	wire [2:0] w_n2783_15;
	wire [2:0] w_n2783_16;
	wire [2:0] w_n2783_17;
	wire [2:0] w_n2783_18;
	wire [2:0] w_n2783_19;
	wire [2:0] w_n2783_20;
	wire [2:0] w_n2783_21;
	wire [2:0] w_n2783_22;
	wire [2:0] w_n2783_23;
	wire [2:0] w_n2783_24;
	wire [2:0] w_n2783_25;
	wire [2:0] w_n2783_26;
	wire [2:0] w_n2783_27;
	wire [2:0] w_n2783_28;
	wire [2:0] w_n2783_29;
	wire [2:0] w_n2783_30;
	wire [2:0] w_n2783_31;
	wire [2:0] w_n2783_32;
	wire [2:0] w_n2783_33;
	wire [2:0] w_n2783_34;
	wire [2:0] w_n2783_35;
	wire [2:0] w_n2783_36;
	wire [2:0] w_n2783_37;
	wire [2:0] w_n2783_38;
	wire [2:0] w_n2783_39;
	wire [2:0] w_n2783_40;
	wire [2:0] w_n2783_41;
	wire [2:0] w_n2783_42;
	wire [2:0] w_n2783_43;
	wire [2:0] w_n2783_44;
	wire [2:0] w_n2783_45;
	wire [2:0] w_n2783_46;
	wire [2:0] w_n2783_47;
	wire [2:0] w_n2783_48;
	wire [2:0] w_n2783_49;
	wire [2:0] w_n2783_50;
	wire [2:0] w_n2783_51;
	wire [2:0] w_n2783_52;
	wire [2:0] w_n2783_53;
	wire [2:0] w_n2783_54;
	wire [2:0] w_n2783_55;
	wire [2:0] w_n2783_56;
	wire [2:0] w_n2783_57;
	wire [2:0] w_n2783_58;
	wire [2:0] w_n2783_59;
	wire [2:0] w_n2783_60;
	wire [2:0] w_n2783_61;
	wire [2:0] w_n2783_62;
	wire [2:0] w_n2783_63;
	wire [2:0] w_n2783_64;
	wire [1:0] w_n2785_0;
	wire [1:0] w_n2786_0;
	wire [2:0] w_n2789_0;
	wire [1:0] w_n2790_0;
	wire [2:0] w_n2793_0;
	wire [1:0] w_n2796_0;
	wire [1:0] w_n2797_0;
	wire [1:0] w_n2798_0;
	wire [1:0] w_n2800_0;
	wire [2:0] w_n2804_0;
	wire [1:0] w_n2807_0;
	wire [1:0] w_n2808_0;
	wire [1:0] w_n2809_0;
	wire [1:0] w_n2811_0;
	wire [2:0] w_n2815_0;
	wire [1:0] w_n2818_0;
	wire [1:0] w_n2819_0;
	wire [1:0] w_n2820_0;
	wire [1:0] w_n2822_0;
	wire [2:0] w_n2826_0;
	wire [1:0] w_n2829_0;
	wire [1:0] w_n2830_0;
	wire [1:0] w_n2831_0;
	wire [1:0] w_n2833_0;
	wire [2:0] w_n2837_0;
	wire [1:0] w_n2840_0;
	wire [1:0] w_n2841_0;
	wire [1:0] w_n2842_0;
	wire [1:0] w_n2844_0;
	wire [2:0] w_n2848_0;
	wire [1:0] w_n2851_0;
	wire [1:0] w_n2852_0;
	wire [1:0] w_n2853_0;
	wire [1:0] w_n2857_0;
	wire [1:0] w_n2858_0;
	wire [2:0] w_n2861_0;
	wire [1:0] w_n2862_0;
	wire [2:0] w_n2865_0;
	wire [1:0] w_n2868_0;
	wire [1:0] w_n2869_0;
	wire [1:0] w_n2870_0;
	wire [1:0] w_n2872_0;
	wire [2:0] w_n2876_0;
	wire [1:0] w_n2879_0;
	wire [1:0] w_n2880_0;
	wire [1:0] w_n2881_0;
	wire [1:0] w_n2883_0;
	wire [2:0] w_n2887_0;
	wire [1:0] w_n2890_0;
	wire [1:0] w_n2891_0;
	wire [1:0] w_n2892_0;
	wire [2:0] w_n2896_0;
	wire [2:0] w_n2899_0;
	wire [1:0] w_n2899_1;
	wire [1:0] w_n2900_0;
	wire [1:0] w_n2903_0;
	wire [1:0] w_n2904_0;
	wire [2:0] w_n2907_0;
	wire [1:0] w_n2908_0;
	wire [1:0] w_n2909_0;
	wire [1:0] w_n2912_0;
	wire [1:0] w_n2913_0;
	wire [2:0] w_n2916_0;
	wire [1:0] w_n2917_0;
	wire [1:0] w_n2920_0;
	wire [1:0] w_n2921_0;
	wire [2:0] w_n2924_0;
	wire [1:0] w_n2925_0;
	wire [2:0] w_n2928_0;
	wire [1:0] w_n2931_0;
	wire [1:0] w_n2932_0;
	wire [1:0] w_n2933_0;
	wire [1:0] w_n2935_0;
	wire [2:0] w_n2939_0;
	wire [1:0] w_n2942_0;
	wire [1:0] w_n2943_0;
	wire [1:0] w_n2944_0;
	wire [1:0] w_n2946_0;
	wire [2:0] w_n2950_0;
	wire [1:0] w_n2953_0;
	wire [1:0] w_n2954_0;
	wire [1:0] w_n2955_0;
	wire [1:0] w_n2957_0;
	wire [2:0] w_n2961_0;
	wire [1:0] w_n2964_0;
	wire [1:0] w_n2965_0;
	wire [1:0] w_n2966_0;
	wire [1:0] w_n2968_0;
	wire [2:0] w_n2972_0;
	wire [1:0] w_n2975_0;
	wire [1:0] w_n2976_0;
	wire [1:0] w_n2977_0;
	wire [1:0] w_n2979_0;
	wire [2:0] w_n2983_0;
	wire [2:0] w_n2986_0;
	wire [1:0] w_n2989_0;
	wire [1:0] w_n2990_0;
	wire [1:0] w_n2991_0;
	wire [1:0] w_n2993_0;
	wire [2:0] w_n2997_0;
	wire [2:0] w_n3001_0;
	wire [1:0] w_n3005_0;
	wire [1:0] w_n3006_0;
	wire [2:0] w_n3009_0;
	wire [1:0] w_n3010_0;
	wire [1:0] w_n3011_0;
	wire [1:0] w_n3014_0;
	wire [2:0] w_n3017_0;
	wire [1:0] w_n3018_0;
	wire [2:0] w_n3021_0;
	wire [1:0] w_n3025_0;
	wire [1:0] w_n3028_0;
	wire [1:0] w_n3037_0;
	wire [2:0] w_n3040_0;
	wire [1:0] w_n3040_1;
	wire [1:0] w_n3044_0;
	wire [2:0] w_n3047_0;
	wire [1:0] w_n3047_1;
	wire [1:0] w_n3053_0;
	wire [1:0] w_n3054_0;
	wire [2:0] w_n3057_0;
	wire [1:0] w_n3058_0;
	wire [1:0] w_n3061_0;
	wire [1:0] w_n3064_0;
	wire [2:0] w_n3067_0;
	wire [1:0] w_n3067_1;
	wire [1:0] w_n3068_0;
	wire [1:0] w_n3086_0;
	wire [1:0] w_n3090_0;
	wire [2:0] w_n3095_0;
	wire [1:0] w_n3098_0;
	wire [1:0] w_n3099_0;
	wire [1:0] w_n3100_0;
	wire [1:0] w_n3107_0;
	wire [2:0] w_n3119_0;
	wire [1:0] w_n3122_0;
	wire [1:0] w_n3123_0;
	wire [1:0] w_n3126_0;
	wire [1:0] w_n3130_0;
	wire [2:0] w_n3148_0;
	wire [1:0] w_n3151_0;
	wire [1:0] w_n3152_0;
	wire [1:0] w_n3155_0;
	wire [1:0] w_n3159_0;
	wire [1:0] w_n3160_0;
	wire [2:0] w_n3163_0;
	wire [1:0] w_n3167_0;
	wire [1:0] w_n3168_0;
	wire [2:0] w_n3171_0;
	wire [1:0] w_n3172_0;
	wire [2:0] w_n3175_0;
	wire [1:0] w_n3178_0;
	wire [1:0] w_n3179_0;
	wire [1:0] w_n3182_0;
	wire [1:0] w_n3186_0;
	wire [1:0] w_n3187_0;
	wire [2:0] w_n3190_0;
	wire [1:0] w_n3191_0;
	wire [1:0] w_n3194_0;
	wire [1:0] w_n3195_0;
	wire [2:0] w_n3198_0;
	wire [2:0] w_n3202_0;
	wire [1:0] w_n3205_0;
	wire [1:0] w_n3206_0;
	wire [1:0] w_n3209_0;
	wire [2:0] w_n3213_0;
	wire [1:0] w_n3216_0;
	wire [1:0] w_n3217_0;
	wire [1:0] w_n3222_0;
	wire [1:0] w_n3223_0;
	wire [2:0] w_n3226_0;
	wire [1:0] w_n3227_0;
	wire [1:0] w_n3233_0;
	wire [1:0] w_n3255_0;
	wire [1:0] w_n3259_0;
	wire [1:0] w_n3260_0;
	wire [2:0] w_n3263_0;
	wire [1:0] w_n3267_0;
	wire [1:0] w_n3268_0;
	wire [2:0] w_n3271_0;
	wire [1:0] w_n3272_0;
	wire [2:0] w_n3275_0;
	wire [1:0] w_n3278_0;
	wire [1:0] w_n3279_0;
	wire [1:0] w_n3282_0;
	wire [1:0] w_n3285_0;
	wire [1:0] w_n3286_0;
	wire [2:0] w_n3289_0;
	wire [1:0] w_n3293_0;
	wire [1:0] w_n3294_0;
	wire [2:0] w_n3297_0;
	wire [1:0] w_n3299_0;
	wire [1:0] w_n3302_0;
	wire [1:0] w_n3303_0;
	wire [2:0] w_n3306_0;
	wire [1:0] w_n3307_0;
	wire [1:0] w_n3310_0;
	wire [1:0] w_n3311_0;
	wire [2:0] w_n3314_0;
	wire [1:0] w_n3318_0;
	wire [1:0] w_n3319_0;
	wire [2:0] w_n3322_0;
	wire [1:0] w_n3323_0;
	wire [1:0] w_n3327_0;
	wire [1:0] w_n3348_0;
	wire [1:0] w_n3352_0;
	wire [1:0] w_n3353_0;
	wire [2:0] w_n3356_0;
	wire [1:0] w_n3357_0;
	wire [1:0] w_n3360_0;
	wire [1:0] w_n3361_0;
	wire [2:0] w_n3364_0;
	wire [2:0] w_n3368_0;
	wire [1:0] w_n3371_0;
	wire [1:0] w_n3372_0;
	wire [1:0] w_n3375_0;
	wire [1:0] w_n3378_0;
	wire [1:0] w_n3379_0;
	wire [2:0] w_n3382_0;
	wire [1:0] w_n3384_0;
	wire [1:0] w_n3387_0;
	wire [1:0] w_n3388_0;
	wire [1:0] w_n3391_0;
	wire [1:0] w_n3392_0;
	wire [1:0] w_n3395_0;
	wire [1:0] w_n3398_0;
	wire [1:0] w_n3399_0;
	wire [2:0] w_n3402_0;
	wire [2:0] w_n3406_0;
	wire [1:0] w_n3409_0;
	wire [1:0] w_n3410_0;
	wire [1:0] w_n3412_0;
	wire [2:0] w_n3415_0;
	wire [1:0] w_n3418_0;
	wire [1:0] w_n3419_0;
	wire [1:0] w_n3423_0;
	wire [1:0] w_n3444_0;
	wire [1:0] w_n3448_0;
	wire [1:0] w_n3449_0;
	wire [2:0] w_n3452_0;
	wire [1:0] w_n3456_0;
	wire [1:0] w_n3457_0;
	wire [2:0] w_n3460_0;
	wire [1:0] w_n3461_0;
	wire [2:0] w_n3464_0;
	wire [1:0] w_n3467_0;
	wire [1:0] w_n3468_0;
	wire [1:0] w_n3471_0;
	wire [1:0] w_n3474_0;
	wire [1:0] w_n3475_0;
	wire [2:0] w_n3478_0;
	wire [1:0] w_n3482_0;
	wire [1:0] w_n3483_0;
	wire [2:0] w_n3486_0;
	wire [1:0] w_n3488_0;
	wire [1:0] w_n3491_0;
	wire [1:0] w_n3492_0;
	wire [2:0] w_n3495_0;
	wire [1:0] w_n3496_0;
	wire [1:0] w_n3499_0;
	wire [1:0] w_n3500_0;
	wire [2:0] w_n3503_0;
	wire [1:0] w_n3507_0;
	wire [1:0] w_n3508_0;
	wire [2:0] w_n3511_0;
	wire [1:0] w_n3512_0;
	wire [1:0] w_n3516_0;
	wire [1:0] w_n3537_0;
	wire [1:0] w_n3541_0;
	wire [1:0] w_n3542_0;
	wire [2:0] w_n3545_0;
	wire [2:0] w_n3549_0;
	wire [1:0] w_n3552_0;
	wire [1:0] w_n3553_0;
	wire [1:0] w_n3555_0;
	wire [1:0] w_n3558_0;
	wire [1:0] w_n3559_0;
	wire [2:0] w_n3562_0;
	wire [1:0] w_n3563_0;
	wire [2:0] w_n3566_0;
	wire [1:0] w_n3569_0;
	wire [1:0] w_n3570_0;
	wire [1:0] w_n3573_0;
	wire [1:0] w_n3583_0;
	wire [1:0] w_n3587_0;
	wire [1:0] w_n3588_0;
	wire [2:0] w_n3591_0;
	wire [1:0] w_n3595_0;
	wire [1:0] w_n3596_0;
	wire [2:0] w_n3599_0;
	wire [1:0] w_n3603_0;
	wire [1:0] w_n3604_0;
	wire [2:0] w_n3607_0;
	wire [1:0] w_n3608_0;
	wire [2:0] w_n3611_0;
	wire [1:0] w_n3614_0;
	wire [1:0] w_n3615_0;
	wire [1:0] w_n3618_0;
	wire [1:0] w_n3619_0;
	wire [1:0] w_n3629_0;
	wire [1:0] w_n3633_0;
	wire [1:0] w_n3634_0;
	wire [2:0] w_n3637_0;
	wire [2:0] w_n3641_0;
	wire [1:0] w_n3644_0;
	wire [1:0] w_n3645_0;
	wire [1:0] w_n3647_0;
	wire [1:0] w_n3650_0;
	wire [1:0] w_n3651_0;
	wire [2:0] w_n3654_0;
	wire [1:0] w_n3655_0;
	wire [2:0] w_n3658_0;
	wire [1:0] w_n3661_0;
	wire [1:0] w_n3662_0;
	wire [1:0] w_n3665_0;
	wire [1:0] w_n3675_0;
	wire [1:0] w_n3679_0;
	wire [1:0] w_n3680_0;
	wire [2:0] w_n3683_0;
	wire [1:0] w_n3687_0;
	wire [1:0] w_n3688_0;
	wire [2:0] w_n3691_0;
	wire [1:0] w_n3695_0;
	wire [1:0] w_n3696_0;
	wire [2:0] w_n3699_0;
	wire [1:0] w_n3700_0;
	wire [2:0] w_n3703_0;
	wire [1:0] w_n3706_0;
	wire [1:0] w_n3707_0;
	wire [1:0] w_n3710_0;
	wire [1:0] w_n3711_0;
	wire [1:0] w_n3721_0;
	wire [1:0] w_n3725_0;
	wire [1:0] w_n3726_0;
	wire [2:0] w_n3729_0;
	wire [2:0] w_n3733_0;
	wire [1:0] w_n3736_0;
	wire [1:0] w_n3737_0;
	wire [1:0] w_n3739_0;
	wire [1:0] w_n3742_0;
	wire [1:0] w_n3743_0;
	wire [2:0] w_n3746_0;
	wire [1:0] w_n3747_0;
	wire [2:0] w_n3750_0;
	wire [1:0] w_n3753_0;
	wire [1:0] w_n3754_0;
	wire [1:0] w_n3757_0;
	wire [1:0] w_n3767_0;
	wire [1:0] w_n3771_0;
	wire [1:0] w_n3772_0;
	wire [2:0] w_n3775_0;
	wire [1:0] w_n3779_0;
	wire [1:0] w_n3780_0;
	wire [2:0] w_n3783_0;
	wire [1:0] w_n3787_0;
	wire [1:0] w_n3788_0;
	wire [2:0] w_n3791_0;
	wire [1:0] w_n3792_0;
	wire [2:0] w_n3795_0;
	wire [1:0] w_n3798_0;
	wire [1:0] w_n3799_0;
	wire [1:0] w_n3802_0;
	wire [1:0] w_n3803_0;
	wire [1:0] w_n3813_0;
	wire [1:0] w_n3817_0;
	wire [1:0] w_n3818_0;
	wire [2:0] w_n3821_0;
	wire [2:0] w_n3825_0;
	wire [1:0] w_n3828_0;
	wire [1:0] w_n3829_0;
	wire [1:0] w_n3831_0;
	wire [1:0] w_n3834_0;
	wire [1:0] w_n3835_0;
	wire [2:0] w_n3838_0;
	wire [1:0] w_n3839_0;
	wire [2:0] w_n3842_0;
	wire [1:0] w_n3845_0;
	wire [1:0] w_n3846_0;
	wire [1:0] w_n3849_0;
	wire [1:0] w_n3859_0;
	wire [1:0] w_n3863_0;
	wire [1:0] w_n3864_0;
	wire [2:0] w_n3867_0;
	wire [1:0] w_n3871_0;
	wire [1:0] w_n3872_0;
	wire [2:0] w_n3875_0;
	wire [1:0] w_n3879_0;
	wire [1:0] w_n3880_0;
	wire [2:0] w_n3883_0;
	wire [1:0] w_n3884_0;
	wire [2:0] w_n3887_0;
	wire [1:0] w_n3890_0;
	wire [1:0] w_n3891_0;
	wire [1:0] w_n3894_0;
	wire [1:0] w_n3895_0;
	wire [1:0] w_n3905_0;
	wire [1:0] w_n3909_0;
	wire [1:0] w_n3910_0;
	wire [2:0] w_n3913_0;
	wire [2:0] w_n3917_0;
	wire [1:0] w_n3920_0;
	wire [1:0] w_n3921_0;
	wire [1:0] w_n3923_0;
	wire [1:0] w_n3926_0;
	wire [1:0] w_n3927_0;
	wire [2:0] w_n3930_0;
	wire [1:0] w_n3931_0;
	wire [2:0] w_n3934_0;
	wire [1:0] w_n3937_0;
	wire [1:0] w_n3938_0;
	wire [1:0] w_n3941_0;
	wire [1:0] w_n3951_0;
	wire [1:0] w_n3955_0;
	wire [1:0] w_n3956_0;
	wire [2:0] w_n3959_0;
	wire [1:0] w_n3963_0;
	wire [1:0] w_n3964_0;
	wire [2:0] w_n3967_0;
	wire [1:0] w_n3971_0;
	wire [1:0] w_n3972_0;
	wire [2:0] w_n3975_0;
	wire [1:0] w_n3976_0;
	wire [2:0] w_n3979_0;
	wire [1:0] w_n3982_0;
	wire [1:0] w_n3983_0;
	wire [1:0] w_n3986_0;
	wire [1:0] w_n3987_0;
	wire [1:0] w_n3997_0;
	wire [1:0] w_n4001_0;
	wire [1:0] w_n4002_0;
	wire [2:0] w_n4005_0;
	wire [2:0] w_n4009_0;
	wire [1:0] w_n4012_0;
	wire [1:0] w_n4013_0;
	wire [1:0] w_n4015_0;
	wire [1:0] w_n4018_0;
	wire [1:0] w_n4019_0;
	wire [2:0] w_n4022_0;
	wire [1:0] w_n4023_0;
	wire [2:0] w_n4026_0;
	wire [1:0] w_n4029_0;
	wire [1:0] w_n4030_0;
	wire [1:0] w_n4033_0;
	wire [1:0] w_n4043_0;
	wire [1:0] w_n4047_0;
	wire [1:0] w_n4048_0;
	wire [2:0] w_n4051_0;
	wire [1:0] w_n4055_0;
	wire [1:0] w_n4056_0;
	wire [2:0] w_n4059_0;
	wire [1:0] w_n4063_0;
	wire [1:0] w_n4064_0;
	wire [2:0] w_n4067_0;
	wire [1:0] w_n4068_0;
	wire [2:0] w_n4071_0;
	wire [1:0] w_n4074_0;
	wire [1:0] w_n4075_0;
	wire [1:0] w_n4078_0;
	wire [1:0] w_n4079_0;
	wire [1:0] w_n4089_0;
	wire [1:0] w_n4093_0;
	wire [1:0] w_n4094_0;
	wire [2:0] w_n4097_0;
	wire [2:0] w_n4101_0;
	wire [1:0] w_n4104_0;
	wire [1:0] w_n4105_0;
	wire [1:0] w_n4107_0;
	wire [1:0] w_n4110_0;
	wire [1:0] w_n4111_0;
	wire [2:0] w_n4114_0;
	wire [1:0] w_n4115_0;
	wire [2:0] w_n4118_0;
	wire [1:0] w_n4121_0;
	wire [1:0] w_n4122_0;
	wire [1:0] w_n4125_0;
	wire [1:0] w_n4135_0;
	wire [1:0] w_n4139_0;
	wire [1:0] w_n4140_0;
	wire [2:0] w_n4143_0;
	wire [1:0] w_n4147_0;
	wire [1:0] w_n4148_0;
	wire [2:0] w_n4151_0;
	wire [1:0] w_n4155_0;
	wire [1:0] w_n4156_0;
	wire [2:0] w_n4159_0;
	wire [1:0] w_n4160_0;
	wire [2:0] w_n4163_0;
	wire [1:0] w_n4166_0;
	wire [1:0] w_n4167_0;
	wire [1:0] w_n4170_0;
	wire [1:0] w_n4171_0;
	wire [1:0] w_n4181_0;
	wire [1:0] w_n4185_0;
	wire [1:0] w_n4186_0;
	wire [2:0] w_n4189_0;
	wire [2:0] w_n4193_0;
	wire [1:0] w_n4196_0;
	wire [1:0] w_n4197_0;
	wire [1:0] w_n4199_0;
	wire [1:0] w_n4202_0;
	wire [1:0] w_n4203_0;
	wire [2:0] w_n4206_0;
	wire [1:0] w_n4207_0;
	wire [2:0] w_n4210_0;
	wire [1:0] w_n4213_0;
	wire [1:0] w_n4214_0;
	wire [1:0] w_n4217_0;
	wire [1:0] w_n4227_0;
	wire [1:0] w_n4231_0;
	wire [1:0] w_n4232_0;
	wire [2:0] w_n4235_0;
	wire [1:0] w_n4239_0;
	wire [1:0] w_n4240_0;
	wire [2:0] w_n4243_0;
	wire [1:0] w_n4245_0;
	wire [1:0] w_n4246_0;
	wire [1:0] w_n4247_0;
	wire [2:0] w_n4248_0;
	wire [1:0] w_n4249_0;
	wire [1:0] w_n4252_0;
	wire [1:0] w_n4253_0;
	wire [2:0] w_n4256_0;
	wire [1:0] w_n4259_0;
	wire [1:0] w_n4269_0;
	wire [1:0] w_n4274_0;
	wire [1:0] w_n4290_0;
	wire [2:0] w_n4293_0;
	wire [1:0] w_n4298_0;
	wire [1:0] w_n4308_0;
	wire [1:0] w_n4309_0;
	wire [1:0] w_n4313_0;
	wire [1:0] w_n4314_0;
	wire [1:0] w_n4324_0;
	wire [1:0] w_n4344_0;
	wire [2:0] w_n4452_0;
	wire [2:0] w_n4452_1;
	wire [2:0] w_n4452_2;
	wire [2:0] w_n4452_3;
	wire [2:0] w_n4452_4;
	wire [2:0] w_n4452_5;
	wire [2:0] w_n4452_6;
	wire [2:0] w_n4452_7;
	wire [2:0] w_n4452_8;
	wire [2:0] w_n4452_9;
	wire [2:0] w_n4452_10;
	wire [2:0] w_n4452_11;
	wire [2:0] w_n4452_12;
	wire [2:0] w_n4452_13;
	wire [2:0] w_n4452_14;
	wire [2:0] w_n4452_15;
	wire [2:0] w_n4452_16;
	wire [2:0] w_n4452_17;
	wire [2:0] w_n4452_18;
	wire [2:0] w_n4452_19;
	wire [2:0] w_n4452_20;
	wire [2:0] w_n4452_21;
	wire [2:0] w_n4452_22;
	wire [2:0] w_n4452_23;
	wire [2:0] w_n4452_24;
	wire [2:0] w_n4452_25;
	wire [2:0] w_n4452_26;
	wire [2:0] w_n4452_27;
	wire [2:0] w_n4452_28;
	wire [2:0] w_n4452_29;
	wire [2:0] w_n4452_30;
	wire [2:0] w_n4452_31;
	wire [2:0] w_n4452_32;
	wire [2:0] w_n4452_33;
	wire [2:0] w_n4452_34;
	wire [2:0] w_n4452_35;
	wire [2:0] w_n4452_36;
	wire [2:0] w_n4452_37;
	wire [2:0] w_n4452_38;
	wire [2:0] w_n4452_39;
	wire [2:0] w_n4452_40;
	wire [2:0] w_n4452_41;
	wire [2:0] w_n4452_42;
	wire [2:0] w_n4452_43;
	wire [2:0] w_n4452_44;
	wire [2:0] w_n4452_45;
	wire [2:0] w_n4452_46;
	wire [2:0] w_n4452_47;
	wire [2:0] w_n4452_48;
	wire [2:0] w_n4452_49;
	wire [2:0] w_n4452_50;
	wire [2:0] w_n4452_51;
	wire [2:0] w_n4452_52;
	wire [2:0] w_n4452_53;
	wire [2:0] w_n4452_54;
	wire [2:0] w_n4452_55;
	wire [2:0] w_n4452_56;
	wire [2:0] w_n4452_57;
	wire [2:0] w_n4452_58;
	wire [2:0] w_n4452_59;
	wire [2:0] w_n4452_60;
	wire [2:0] w_n4452_61;
	wire [2:0] w_n4452_62;
	wire [1:0] w_n4452_63;
	jnot g0000(.din(w_in230_0[2]),.dout(n642),.clk(gclk));
	jand g0001(.dina(w_in330_0[2]),.dinb(n642),.dout(n643),.clk(gclk));
	jnot g0002(.din(w_n643_0[1]),.dout(n644),.clk(gclk));
	jnot g0003(.din(w_in329_0[2]),.dout(n645),.clk(gclk));
	jand g0004(.dina(n645),.dinb(w_in229_0[2]),.dout(n646),.clk(gclk));
	jnot g0005(.din(w_in229_0[1]),.dout(n647),.clk(gclk));
	jand g0006(.dina(w_in329_0[1]),.dinb(n647),.dout(n648),.clk(gclk));
	jnot g0007(.din(w_n648_0[1]),.dout(n649),.clk(gclk));
	jnot g0008(.din(w_in328_0[2]),.dout(n650),.clk(gclk));
	jand g0009(.dina(n650),.dinb(w_in228_0[2]),.dout(n651),.clk(gclk));
	jnot g0010(.din(w_in228_0[1]),.dout(n652),.clk(gclk));
	jand g0011(.dina(w_in328_0[1]),.dinb(n652),.dout(n653),.clk(gclk));
	jnot g0012(.din(w_n653_0[1]),.dout(n654),.clk(gclk));
	jnot g0013(.din(w_in327_0[2]),.dout(n655),.clk(gclk));
	jand g0014(.dina(n655),.dinb(w_in227_0[2]),.dout(n656),.clk(gclk));
	jnot g0015(.din(w_in227_0[1]),.dout(n657),.clk(gclk));
	jand g0016(.dina(w_in327_0[1]),.dinb(n657),.dout(n658),.clk(gclk));
	jnot g0017(.din(w_n658_0[1]),.dout(n659),.clk(gclk));
	jnot g0018(.din(w_in326_0[2]),.dout(n660),.clk(gclk));
	jand g0019(.dina(n660),.dinb(w_in226_0[2]),.dout(n661),.clk(gclk));
	jnot g0020(.din(w_in226_0[1]),.dout(n662),.clk(gclk));
	jand g0021(.dina(w_in326_0[1]),.dinb(n662),.dout(n663),.clk(gclk));
	jnot g0022(.din(w_n663_0[1]),.dout(n664),.clk(gclk));
	jnot g0023(.din(w_in325_0[2]),.dout(n665),.clk(gclk));
	jand g0024(.dina(n665),.dinb(w_in225_0[2]),.dout(n666),.clk(gclk));
	jnot g0025(.din(w_in225_0[1]),.dout(n667),.clk(gclk));
	jand g0026(.dina(w_in325_0[1]),.dinb(n667),.dout(n668),.clk(gclk));
	jnot g0027(.din(w_n668_0[1]),.dout(n669),.clk(gclk));
	jnot g0028(.din(w_in324_0[2]),.dout(n670),.clk(gclk));
	jand g0029(.dina(n670),.dinb(w_in224_0[2]),.dout(n671),.clk(gclk));
	jnot g0030(.din(w_in224_0[1]),.dout(n672),.clk(gclk));
	jand g0031(.dina(w_in324_0[1]),.dinb(n672),.dout(n673),.clk(gclk));
	jnot g0032(.din(w_n673_0[1]),.dout(n674),.clk(gclk));
	jnot g0033(.din(w_in323_0[2]),.dout(n675),.clk(gclk));
	jand g0034(.dina(n675),.dinb(w_in223_0[2]),.dout(n676),.clk(gclk));
	jnot g0035(.din(w_in223_0[1]),.dout(n677),.clk(gclk));
	jand g0036(.dina(w_in323_0[1]),.dinb(n677),.dout(n678),.clk(gclk));
	jnot g0037(.din(w_n678_0[1]),.dout(n679),.clk(gclk));
	jnot g0038(.din(w_in322_0[2]),.dout(n680),.clk(gclk));
	jand g0039(.dina(n680),.dinb(w_in222_0[2]),.dout(n681),.clk(gclk));
	jnot g0040(.din(w_in222_0[1]),.dout(n682),.clk(gclk));
	jand g0041(.dina(w_in322_0[1]),.dinb(n682),.dout(n683),.clk(gclk));
	jnot g0042(.din(w_n683_0[1]),.dout(n684),.clk(gclk));
	jnot g0043(.din(w_in321_0[2]),.dout(n685),.clk(gclk));
	jand g0044(.dina(n685),.dinb(w_in221_0[2]),.dout(n686),.clk(gclk));
	jnot g0045(.din(w_in221_0[1]),.dout(n687),.clk(gclk));
	jand g0046(.dina(w_in321_0[1]),.dinb(n687),.dout(n688),.clk(gclk));
	jnot g0047(.din(w_n688_0[1]),.dout(n689),.clk(gclk));
	jnot g0048(.din(w_in320_0[2]),.dout(n690),.clk(gclk));
	jand g0049(.dina(n690),.dinb(w_in220_0[2]),.dout(n691),.clk(gclk));
	jnot g0050(.din(w_in220_0[1]),.dout(n692),.clk(gclk));
	jand g0051(.dina(w_in320_0[1]),.dinb(n692),.dout(n693),.clk(gclk));
	jnot g0052(.din(w_n693_0[1]),.dout(n694),.clk(gclk));
	jnot g0053(.din(w_in319_0[2]),.dout(n695),.clk(gclk));
	jand g0054(.dina(n695),.dinb(w_in219_0[2]),.dout(n696),.clk(gclk));
	jnot g0055(.din(w_in219_0[1]),.dout(n697),.clk(gclk));
	jand g0056(.dina(w_in319_0[1]),.dinb(n697),.dout(n698),.clk(gclk));
	jnot g0057(.din(w_n698_0[1]),.dout(n699),.clk(gclk));
	jnot g0058(.din(w_in318_0[2]),.dout(n700),.clk(gclk));
	jand g0059(.dina(n700),.dinb(w_in218_0[2]),.dout(n701),.clk(gclk));
	jnot g0060(.din(w_in218_0[1]),.dout(n702),.clk(gclk));
	jand g0061(.dina(w_in318_0[1]),.dinb(n702),.dout(n703),.clk(gclk));
	jnot g0062(.din(w_n703_0[1]),.dout(n704),.clk(gclk));
	jnot g0063(.din(w_in317_0[2]),.dout(n705),.clk(gclk));
	jand g0064(.dina(n705),.dinb(w_in217_0[2]),.dout(n706),.clk(gclk));
	jnot g0065(.din(w_in217_0[1]),.dout(n707),.clk(gclk));
	jand g0066(.dina(w_in317_0[1]),.dinb(n707),.dout(n708),.clk(gclk));
	jnot g0067(.din(w_n708_0[1]),.dout(n709),.clk(gclk));
	jnot g0068(.din(w_in316_0[2]),.dout(n710),.clk(gclk));
	jand g0069(.dina(n710),.dinb(w_in216_0[2]),.dout(n711),.clk(gclk));
	jnot g0070(.din(w_in216_0[1]),.dout(n712),.clk(gclk));
	jand g0071(.dina(w_in316_0[1]),.dinb(n712),.dout(n713),.clk(gclk));
	jnot g0072(.din(w_n713_0[1]),.dout(n714),.clk(gclk));
	jnot g0073(.din(w_in315_0[2]),.dout(n715),.clk(gclk));
	jand g0074(.dina(n715),.dinb(w_in215_0[2]),.dout(n716),.clk(gclk));
	jnot g0075(.din(w_in215_0[1]),.dout(n717),.clk(gclk));
	jand g0076(.dina(w_in315_0[1]),.dinb(n717),.dout(n718),.clk(gclk));
	jnot g0077(.din(w_n718_0[1]),.dout(n719),.clk(gclk));
	jnot g0078(.din(w_in314_0[2]),.dout(n720),.clk(gclk));
	jand g0079(.dina(n720),.dinb(w_in214_0[2]),.dout(n721),.clk(gclk));
	jnot g0080(.din(w_in214_0[1]),.dout(n722),.clk(gclk));
	jand g0081(.dina(w_in314_0[1]),.dinb(n722),.dout(n723),.clk(gclk));
	jnot g0082(.din(w_n723_0[1]),.dout(n724),.clk(gclk));
	jnot g0083(.din(w_in313_0[2]),.dout(n725),.clk(gclk));
	jand g0084(.dina(n725),.dinb(w_in213_0[2]),.dout(n726),.clk(gclk));
	jnot g0085(.din(w_in213_0[1]),.dout(n727),.clk(gclk));
	jand g0086(.dina(w_in313_0[1]),.dinb(n727),.dout(n728),.clk(gclk));
	jnot g0087(.din(w_n728_0[1]),.dout(n729),.clk(gclk));
	jnot g0088(.din(w_in312_0[2]),.dout(n730),.clk(gclk));
	jand g0089(.dina(n730),.dinb(w_in212_0[2]),.dout(n731),.clk(gclk));
	jnot g0090(.din(w_in212_0[1]),.dout(n732),.clk(gclk));
	jand g0091(.dina(w_in312_0[1]),.dinb(n732),.dout(n733),.clk(gclk));
	jnot g0092(.din(w_n733_0[1]),.dout(n734),.clk(gclk));
	jnot g0093(.din(w_in311_0[2]),.dout(n735),.clk(gclk));
	jand g0094(.dina(n735),.dinb(w_in211_0[2]),.dout(n736),.clk(gclk));
	jnot g0095(.din(w_in211_0[1]),.dout(n737),.clk(gclk));
	jand g0096(.dina(w_in311_0[1]),.dinb(n737),.dout(n738),.clk(gclk));
	jnot g0097(.din(w_n738_0[1]),.dout(n739),.clk(gclk));
	jnot g0098(.din(w_in310_0[2]),.dout(n740),.clk(gclk));
	jand g0099(.dina(n740),.dinb(w_in210_0[2]),.dout(n741),.clk(gclk));
	jnot g0100(.din(w_in210_0[1]),.dout(n742),.clk(gclk));
	jand g0101(.dina(w_in310_0[1]),.dinb(n742),.dout(n743),.clk(gclk));
	jnot g0102(.din(w_n743_0[1]),.dout(n744),.clk(gclk));
	jnot g0103(.din(w_in39_0[2]),.dout(n745),.clk(gclk));
	jand g0104(.dina(n745),.dinb(w_in29_0[2]),.dout(n746),.clk(gclk));
	jnot g0105(.din(w_in29_0[1]),.dout(n747),.clk(gclk));
	jand g0106(.dina(w_in39_0[1]),.dinb(n747),.dout(n748),.clk(gclk));
	jnot g0107(.din(w_n748_0[1]),.dout(n749),.clk(gclk));
	jnot g0108(.din(w_in38_0[2]),.dout(n750),.clk(gclk));
	jand g0109(.dina(n750),.dinb(w_in28_0[2]),.dout(n751),.clk(gclk));
	jnot g0110(.din(w_in28_0[1]),.dout(n752),.clk(gclk));
	jand g0111(.dina(w_in38_0[1]),.dinb(n752),.dout(n753),.clk(gclk));
	jnot g0112(.din(w_n753_0[1]),.dout(n754),.clk(gclk));
	jnot g0113(.din(w_in37_0[2]),.dout(n755),.clk(gclk));
	jand g0114(.dina(n755),.dinb(w_in27_0[2]),.dout(n756),.clk(gclk));
	jnot g0115(.din(w_in27_0[1]),.dout(n757),.clk(gclk));
	jand g0116(.dina(w_in37_0[1]),.dinb(n757),.dout(n758),.clk(gclk));
	jnot g0117(.din(w_n758_0[1]),.dout(n759),.clk(gclk));
	jnot g0118(.din(w_in36_0[2]),.dout(n760),.clk(gclk));
	jand g0119(.dina(n760),.dinb(w_in26_0[2]),.dout(n761),.clk(gclk));
	jnot g0120(.din(w_in26_0[1]),.dout(n762),.clk(gclk));
	jand g0121(.dina(w_in36_0[1]),.dinb(n762),.dout(n763),.clk(gclk));
	jnot g0122(.din(w_n763_0[1]),.dout(n764),.clk(gclk));
	jnot g0123(.din(w_in35_0[2]),.dout(n765),.clk(gclk));
	jand g0124(.dina(n765),.dinb(w_in25_0[2]),.dout(n766),.clk(gclk));
	jnot g0125(.din(w_in25_0[1]),.dout(n767),.clk(gclk));
	jand g0126(.dina(w_in35_0[1]),.dinb(n767),.dout(n768),.clk(gclk));
	jnot g0127(.din(w_n768_0[1]),.dout(n769),.clk(gclk));
	jnot g0128(.din(w_in34_0[2]),.dout(n770),.clk(gclk));
	jand g0129(.dina(n770),.dinb(w_in24_0[2]),.dout(n771),.clk(gclk));
	jnot g0130(.din(w_in24_0[1]),.dout(n772),.clk(gclk));
	jand g0131(.dina(w_in34_0[1]),.dinb(n772),.dout(n773),.clk(gclk));
	jnot g0132(.din(w_n773_0[1]),.dout(n774),.clk(gclk));
	jnot g0133(.din(w_in33_0[2]),.dout(n775),.clk(gclk));
	jand g0134(.dina(n775),.dinb(w_in23_0[2]),.dout(n776),.clk(gclk));
	jnot g0135(.din(w_in23_0[1]),.dout(n777),.clk(gclk));
	jand g0136(.dina(w_in33_0[1]),.dinb(n777),.dout(n778),.clk(gclk));
	jnot g0137(.din(w_n778_0[1]),.dout(n779),.clk(gclk));
	jnot g0138(.din(w_in32_0[2]),.dout(n780),.clk(gclk));
	jand g0139(.dina(w_n780_0[1]),.dinb(w_in22_0[2]),.dout(n781),.clk(gclk));
	jnot g0140(.din(w_in22_0[1]),.dout(n782),.clk(gclk));
	jand g0141(.dina(w_in32_0[1]),.dinb(w_n782_0[1]),.dout(n783),.clk(gclk));
	jnot g0142(.din(w_n783_0[1]),.dout(n784),.clk(gclk));
	jnot g0143(.din(w_in31_1[1]),.dout(n785),.clk(gclk));
	jand g0144(.dina(w_n785_0[1]),.dinb(w_in21_1[1]),.dout(n786),.clk(gclk));
	jor g0145(.dina(w_n785_0[0]),.dinb(w_in21_1[0]),.dout(n787),.clk(gclk));
	jnot g0146(.din(w_in30_0[2]),.dout(n788),.clk(gclk));
	jand g0147(.dina(w_n788_0[1]),.dinb(w_in20_0[2]),.dout(n789),.clk(gclk));
	jand g0148(.dina(n789),.dinb(n787),.dout(n790),.clk(gclk));
	jor g0149(.dina(n790),.dinb(n786),.dout(n791),.clk(gclk));
	jand g0150(.dina(n791),.dinb(n784),.dout(n792),.clk(gclk));
	jor g0151(.dina(n792),.dinb(w_n781_0[1]),.dout(n793),.clk(gclk));
	jand g0152(.dina(n793),.dinb(n779),.dout(n794),.clk(gclk));
	jor g0153(.dina(n794),.dinb(w_n776_0[1]),.dout(n795),.clk(gclk));
	jand g0154(.dina(n795),.dinb(n774),.dout(n796),.clk(gclk));
	jor g0155(.dina(n796),.dinb(w_n771_0[1]),.dout(n797),.clk(gclk));
	jand g0156(.dina(n797),.dinb(n769),.dout(n798),.clk(gclk));
	jor g0157(.dina(n798),.dinb(w_n766_0[1]),.dout(n799),.clk(gclk));
	jand g0158(.dina(n799),.dinb(n764),.dout(n800),.clk(gclk));
	jor g0159(.dina(n800),.dinb(w_n761_0[1]),.dout(n801),.clk(gclk));
	jand g0160(.dina(n801),.dinb(n759),.dout(n802),.clk(gclk));
	jor g0161(.dina(n802),.dinb(w_n756_0[1]),.dout(n803),.clk(gclk));
	jand g0162(.dina(n803),.dinb(n754),.dout(n804),.clk(gclk));
	jor g0163(.dina(n804),.dinb(w_n751_0[1]),.dout(n805),.clk(gclk));
	jand g0164(.dina(n805),.dinb(n749),.dout(n806),.clk(gclk));
	jor g0165(.dina(n806),.dinb(w_n746_0[1]),.dout(n807),.clk(gclk));
	jand g0166(.dina(n807),.dinb(n744),.dout(n808),.clk(gclk));
	jor g0167(.dina(n808),.dinb(w_n741_0[1]),.dout(n809),.clk(gclk));
	jand g0168(.dina(n809),.dinb(n739),.dout(n810),.clk(gclk));
	jor g0169(.dina(n810),.dinb(w_n736_0[1]),.dout(n811),.clk(gclk));
	jand g0170(.dina(n811),.dinb(n734),.dout(n812),.clk(gclk));
	jor g0171(.dina(n812),.dinb(w_n731_0[1]),.dout(n813),.clk(gclk));
	jand g0172(.dina(n813),.dinb(n729),.dout(n814),.clk(gclk));
	jor g0173(.dina(n814),.dinb(w_n726_0[1]),.dout(n815),.clk(gclk));
	jand g0174(.dina(n815),.dinb(n724),.dout(n816),.clk(gclk));
	jor g0175(.dina(n816),.dinb(w_n721_0[1]),.dout(n817),.clk(gclk));
	jand g0176(.dina(n817),.dinb(n719),.dout(n818),.clk(gclk));
	jor g0177(.dina(n818),.dinb(w_n716_0[1]),.dout(n819),.clk(gclk));
	jand g0178(.dina(n819),.dinb(n714),.dout(n820),.clk(gclk));
	jor g0179(.dina(n820),.dinb(w_n711_0[1]),.dout(n821),.clk(gclk));
	jand g0180(.dina(n821),.dinb(n709),.dout(n822),.clk(gclk));
	jor g0181(.dina(n822),.dinb(w_n706_0[1]),.dout(n823),.clk(gclk));
	jand g0182(.dina(n823),.dinb(n704),.dout(n824),.clk(gclk));
	jor g0183(.dina(n824),.dinb(w_n701_0[1]),.dout(n825),.clk(gclk));
	jand g0184(.dina(n825),.dinb(n699),.dout(n826),.clk(gclk));
	jor g0185(.dina(n826),.dinb(w_n696_0[1]),.dout(n827),.clk(gclk));
	jand g0186(.dina(n827),.dinb(n694),.dout(n828),.clk(gclk));
	jor g0187(.dina(n828),.dinb(w_n691_0[1]),.dout(n829),.clk(gclk));
	jand g0188(.dina(n829),.dinb(n689),.dout(n830),.clk(gclk));
	jor g0189(.dina(n830),.dinb(w_n686_0[1]),.dout(n831),.clk(gclk));
	jand g0190(.dina(n831),.dinb(n684),.dout(n832),.clk(gclk));
	jor g0191(.dina(n832),.dinb(w_n681_0[1]),.dout(n833),.clk(gclk));
	jand g0192(.dina(n833),.dinb(n679),.dout(n834),.clk(gclk));
	jor g0193(.dina(n834),.dinb(w_n676_0[1]),.dout(n835),.clk(gclk));
	jand g0194(.dina(n835),.dinb(n674),.dout(n836),.clk(gclk));
	jor g0195(.dina(n836),.dinb(w_n671_0[1]),.dout(n837),.clk(gclk));
	jand g0196(.dina(n837),.dinb(n669),.dout(n838),.clk(gclk));
	jor g0197(.dina(n838),.dinb(w_n666_0[1]),.dout(n839),.clk(gclk));
	jand g0198(.dina(n839),.dinb(n664),.dout(n840),.clk(gclk));
	jor g0199(.dina(n840),.dinb(w_n661_0[1]),.dout(n841),.clk(gclk));
	jand g0200(.dina(n841),.dinb(n659),.dout(n842),.clk(gclk));
	jor g0201(.dina(n842),.dinb(w_n656_0[1]),.dout(n843),.clk(gclk));
	jand g0202(.dina(n843),.dinb(n654),.dout(n844),.clk(gclk));
	jor g0203(.dina(n844),.dinb(w_n651_0[1]),.dout(n845),.clk(gclk));
	jand g0204(.dina(n845),.dinb(n649),.dout(n846),.clk(gclk));
	jor g0205(.dina(n846),.dinb(w_n646_0[1]),.dout(n847),.clk(gclk));
	jand g0206(.dina(n847),.dinb(n644),.dout(n848),.clk(gclk));
	jnot g0207(.din(w_in330_0[1]),.dout(n849),.clk(gclk));
	jand g0208(.dina(n849),.dinb(w_in230_0[1]),.dout(n850),.clk(gclk));
	jnot g0209(.din(w_in331_0[2]),.dout(n851),.clk(gclk));
	jand g0210(.dina(n851),.dinb(w_in231_0[2]),.dout(n852),.clk(gclk));
	jor g0211(.dina(n852),.dinb(n850),.dout(n853),.clk(gclk));
	jor g0212(.dina(w_n853_0[1]),.dinb(n848),.dout(n854),.clk(gclk));
	jnot g0213(.din(w_in237_0[2]),.dout(n855),.clk(gclk));
	jand g0214(.dina(w_in337_0[2]),.dinb(n855),.dout(n856),.clk(gclk));
	jnot g0215(.din(w_in239_0[2]),.dout(n857),.clk(gclk));
	jand g0216(.dina(w_in339_0[2]),.dinb(n857),.dout(n858),.clk(gclk));
	jnot g0217(.din(w_in238_0[2]),.dout(n859),.clk(gclk));
	jand g0218(.dina(w_in338_0[2]),.dinb(n859),.dout(n860),.clk(gclk));
	jor g0219(.dina(n860),.dinb(w_n858_0[1]),.dout(n861),.clk(gclk));
	jor g0220(.dina(n861),.dinb(n856),.dout(n862),.clk(gclk));
	jnot g0221(.din(w_in235_0[2]),.dout(n863),.clk(gclk));
	jand g0222(.dina(w_in335_0[2]),.dinb(n863),.dout(n864),.clk(gclk));
	jnot g0223(.din(w_in234_0[2]),.dout(n865),.clk(gclk));
	jand g0224(.dina(w_in334_0[2]),.dinb(n865),.dout(n866),.clk(gclk));
	jor g0225(.dina(n866),.dinb(n864),.dout(n867),.clk(gclk));
	jnot g0226(.din(w_in232_0[2]),.dout(n868),.clk(gclk));
	jand g0227(.dina(w_in332_0[2]),.dinb(n868),.dout(n869),.clk(gclk));
	jnot g0228(.din(w_in233_0[2]),.dout(n870),.clk(gclk));
	jand g0229(.dina(w_in333_0[2]),.dinb(n870),.dout(n871),.clk(gclk));
	jor g0230(.dina(w_n871_0[1]),.dinb(n869),.dout(n872),.clk(gclk));
	jnot g0231(.din(w_in236_0[2]),.dout(n873),.clk(gclk));
	jand g0232(.dina(w_in336_0[2]),.dinb(n873),.dout(n874),.clk(gclk));
	jnot g0233(.din(w_in231_0[1]),.dout(n875),.clk(gclk));
	jand g0234(.dina(w_in331_0[1]),.dinb(n875),.dout(n876),.clk(gclk));
	jor g0235(.dina(n876),.dinb(w_n874_0[1]),.dout(n877),.clk(gclk));
	jor g0236(.dina(n877),.dinb(n872),.dout(n878),.clk(gclk));
	jor g0237(.dina(n878),.dinb(w_n867_0[1]),.dout(n879),.clk(gclk));
	jor g0238(.dina(n879),.dinb(w_n862_0[1]),.dout(n880),.clk(gclk));
	jnot g0239(.din(w_n880_0[1]),.dout(n881),.clk(gclk));
	jand g0240(.dina(n881),.dinb(n854),.dout(n882),.clk(gclk));
	jnot g0241(.din(w_n862_0[0]),.dout(n883),.clk(gclk));
	jnot g0242(.din(w_n874_0[0]),.dout(n884),.clk(gclk));
	jnot g0243(.din(w_in335_0[1]),.dout(n885),.clk(gclk));
	jand g0244(.dina(n885),.dinb(w_in235_0[1]),.dout(n886),.clk(gclk));
	jnot g0245(.din(w_n867_0[0]),.dout(n887),.clk(gclk));
	jnot g0246(.din(w_n871_0[0]),.dout(n888),.clk(gclk));
	jnot g0247(.din(w_in332_0[1]),.dout(n889),.clk(gclk));
	jand g0248(.dina(n889),.dinb(w_in232_0[1]),.dout(n890),.clk(gclk));
	jand g0249(.dina(n890),.dinb(n888),.dout(n891),.clk(gclk));
	jnot g0250(.din(w_in333_0[1]),.dout(n892),.clk(gclk));
	jand g0251(.dina(n892),.dinb(w_in233_0[1]),.dout(n893),.clk(gclk));
	jnot g0252(.din(w_in334_0[1]),.dout(n894),.clk(gclk));
	jand g0253(.dina(n894),.dinb(w_in234_0[1]),.dout(n895),.clk(gclk));
	jor g0254(.dina(n895),.dinb(n893),.dout(n896),.clk(gclk));
	jor g0255(.dina(n896),.dinb(n891),.dout(n897),.clk(gclk));
	jand g0256(.dina(n897),.dinb(n887),.dout(n898),.clk(gclk));
	jor g0257(.dina(n898),.dinb(n886),.dout(n899),.clk(gclk));
	jand g0258(.dina(n899),.dinb(n884),.dout(n900),.clk(gclk));
	jnot g0259(.din(w_in336_0[1]),.dout(n901),.clk(gclk));
	jand g0260(.dina(n901),.dinb(w_in236_0[1]),.dout(n902),.clk(gclk));
	jnot g0261(.din(w_in337_0[1]),.dout(n903),.clk(gclk));
	jand g0262(.dina(n903),.dinb(w_in237_0[1]),.dout(n904),.clk(gclk));
	jor g0263(.dina(n904),.dinb(n902),.dout(n905),.clk(gclk));
	jor g0264(.dina(n905),.dinb(n900),.dout(n906),.clk(gclk));
	jand g0265(.dina(n906),.dinb(n883),.dout(n907),.clk(gclk));
	jnot g0266(.din(w_n858_0[0]),.dout(n908),.clk(gclk));
	jnot g0267(.din(w_in338_0[1]),.dout(n909),.clk(gclk));
	jand g0268(.dina(n909),.dinb(w_in238_0[1]),.dout(n910),.clk(gclk));
	jand g0269(.dina(n910),.dinb(n908),.dout(n911),.clk(gclk));
	jnot g0270(.din(w_in339_0[1]),.dout(n912),.clk(gclk));
	jand g0271(.dina(n912),.dinb(w_in239_0[1]),.dout(n913),.clk(gclk));
	jor g0272(.dina(n913),.dinb(n911),.dout(n914),.clk(gclk));
	jor g0273(.dina(n914),.dinb(n907),.dout(n915),.clk(gclk));
	jor g0274(.dina(w_n915_0[1]),.dinb(n882),.dout(n916),.clk(gclk));
	jnot g0275(.din(w_in245_0[2]),.dout(n917),.clk(gclk));
	jand g0276(.dina(w_in345_0[2]),.dinb(n917),.dout(n918),.clk(gclk));
	jnot g0277(.din(w_in247_0[2]),.dout(n919),.clk(gclk));
	jand g0278(.dina(w_in347_0[2]),.dinb(n919),.dout(n920),.clk(gclk));
	jnot g0279(.din(w_in246_0[2]),.dout(n921),.clk(gclk));
	jand g0280(.dina(w_in346_0[2]),.dinb(n921),.dout(n922),.clk(gclk));
	jor g0281(.dina(n922),.dinb(w_n920_0[1]),.dout(n923),.clk(gclk));
	jor g0282(.dina(n923),.dinb(n918),.dout(n924),.clk(gclk));
	jnot g0283(.din(w_in243_0[2]),.dout(n925),.clk(gclk));
	jand g0284(.dina(w_in343_0[2]),.dinb(n925),.dout(n926),.clk(gclk));
	jnot g0285(.din(w_in242_0[2]),.dout(n927),.clk(gclk));
	jand g0286(.dina(w_in342_0[2]),.dinb(n927),.dout(n928),.clk(gclk));
	jor g0287(.dina(n928),.dinb(n926),.dout(n929),.clk(gclk));
	jnot g0288(.din(w_in244_0[2]),.dout(n930),.clk(gclk));
	jand g0289(.dina(w_in344_0[2]),.dinb(n930),.dout(n931),.clk(gclk));
	jnot g0290(.din(w_in240_0[2]),.dout(n932),.clk(gclk));
	jand g0291(.dina(w_in340_0[2]),.dinb(n932),.dout(n933),.clk(gclk));
	jnot g0292(.din(w_in241_0[2]),.dout(n934),.clk(gclk));
	jand g0293(.dina(w_in341_0[2]),.dinb(n934),.dout(n935),.clk(gclk));
	jor g0294(.dina(w_n935_0[1]),.dinb(n933),.dout(n936),.clk(gclk));
	jor g0295(.dina(n936),.dinb(w_n931_0[1]),.dout(n937),.clk(gclk));
	jor g0296(.dina(n937),.dinb(w_n929_0[1]),.dout(n938),.clk(gclk));
	jor g0297(.dina(n938),.dinb(w_n924_0[1]),.dout(n939),.clk(gclk));
	jnot g0298(.din(w_n939_0[1]),.dout(n940),.clk(gclk));
	jand g0299(.dina(n940),.dinb(n916),.dout(n941),.clk(gclk));
	jnot g0300(.din(w_n924_0[0]),.dout(n942),.clk(gclk));
	jnot g0301(.din(w_n931_0[0]),.dout(n943),.clk(gclk));
	jnot g0302(.din(w_in343_0[1]),.dout(n944),.clk(gclk));
	jand g0303(.dina(n944),.dinb(w_in243_0[1]),.dout(n945),.clk(gclk));
	jnot g0304(.din(w_n929_0[0]),.dout(n946),.clk(gclk));
	jnot g0305(.din(w_n935_0[0]),.dout(n947),.clk(gclk));
	jnot g0306(.din(w_in340_0[1]),.dout(n948),.clk(gclk));
	jand g0307(.dina(n948),.dinb(w_in240_0[1]),.dout(n949),.clk(gclk));
	jand g0308(.dina(n949),.dinb(n947),.dout(n950),.clk(gclk));
	jnot g0309(.din(w_in341_0[1]),.dout(n951),.clk(gclk));
	jand g0310(.dina(n951),.dinb(w_in241_0[1]),.dout(n952),.clk(gclk));
	jnot g0311(.din(w_in342_0[1]),.dout(n953),.clk(gclk));
	jand g0312(.dina(n953),.dinb(w_in242_0[1]),.dout(n954),.clk(gclk));
	jor g0313(.dina(n954),.dinb(n952),.dout(n955),.clk(gclk));
	jor g0314(.dina(n955),.dinb(n950),.dout(n956),.clk(gclk));
	jand g0315(.dina(n956),.dinb(n946),.dout(n957),.clk(gclk));
	jor g0316(.dina(n957),.dinb(n945),.dout(n958),.clk(gclk));
	jand g0317(.dina(n958),.dinb(n943),.dout(n959),.clk(gclk));
	jnot g0318(.din(w_in344_0[1]),.dout(n960),.clk(gclk));
	jand g0319(.dina(n960),.dinb(w_in244_0[1]),.dout(n961),.clk(gclk));
	jnot g0320(.din(w_in345_0[1]),.dout(n962),.clk(gclk));
	jand g0321(.dina(n962),.dinb(w_in245_0[1]),.dout(n963),.clk(gclk));
	jor g0322(.dina(n963),.dinb(n961),.dout(n964),.clk(gclk));
	jor g0323(.dina(n964),.dinb(n959),.dout(n965),.clk(gclk));
	jand g0324(.dina(n965),.dinb(n942),.dout(n966),.clk(gclk));
	jnot g0325(.din(w_n920_0[0]),.dout(n967),.clk(gclk));
	jnot g0326(.din(w_in346_0[1]),.dout(n968),.clk(gclk));
	jand g0327(.dina(n968),.dinb(w_in246_0[1]),.dout(n969),.clk(gclk));
	jand g0328(.dina(n969),.dinb(n967),.dout(n970),.clk(gclk));
	jnot g0329(.din(w_in347_0[1]),.dout(n971),.clk(gclk));
	jand g0330(.dina(n971),.dinb(w_in247_0[1]),.dout(n972),.clk(gclk));
	jor g0331(.dina(n972),.dinb(n970),.dout(n973),.clk(gclk));
	jor g0332(.dina(n973),.dinb(n966),.dout(n974),.clk(gclk));
	jor g0333(.dina(w_n974_0[1]),.dinb(n941),.dout(n975),.clk(gclk));
	jnot g0334(.din(w_in352_0[1]),.dout(n976),.clk(gclk));
	jnot g0335(.din(w_in253_0[2]),.dout(n977),.clk(gclk));
	jand g0336(.dina(w_in353_0[2]),.dinb(n977),.dout(n978),.clk(gclk));
	jnot g0337(.din(n978),.dout(n979),.clk(gclk));
	jand g0338(.dina(w_n979_0[1]),.dinb(n976),.dout(n980),.clk(gclk));
	jand g0339(.dina(w_n979_0[0]),.dinb(w_in252_0[2]),.dout(n981),.clk(gclk));
	jor g0340(.dina(n981),.dinb(w_n980_0[1]),.dout(n982),.clk(gclk));
	jnot g0341(.din(w_n982_0[1]),.dout(n983),.clk(gclk));
	jnot g0342(.din(w_in255_0[2]),.dout(n984),.clk(gclk));
	jand g0343(.dina(w_in355_0[2]),.dinb(n984),.dout(n985),.clk(gclk));
	jnot g0344(.din(w_in254_0[2]),.dout(n986),.clk(gclk));
	jand g0345(.dina(w_in354_0[2]),.dinb(n986),.dout(n987),.clk(gclk));
	jor g0346(.dina(n987),.dinb(n985),.dout(n988),.clk(gclk));
	jnot g0347(.din(w_in251_0[2]),.dout(n989),.clk(gclk));
	jand g0348(.dina(w_in351_0[2]),.dinb(n989),.dout(n990),.clk(gclk));
	jnot g0349(.din(w_in250_0[2]),.dout(n991),.clk(gclk));
	jand g0350(.dina(w_in350_0[2]),.dinb(n991),.dout(n992),.clk(gclk));
	jor g0351(.dina(n992),.dinb(n990),.dout(n993),.clk(gclk));
	jnot g0352(.din(w_in248_0[2]),.dout(n994),.clk(gclk));
	jand g0353(.dina(w_in348_0[2]),.dinb(n994),.dout(n995),.clk(gclk));
	jnot g0354(.din(w_in249_0[2]),.dout(n996),.clk(gclk));
	jand g0355(.dina(w_in349_0[2]),.dinb(n996),.dout(n997),.clk(gclk));
	jor g0356(.dina(w_n997_0[1]),.dinb(n995),.dout(n998),.clk(gclk));
	jor g0357(.dina(n998),.dinb(w_n993_0[1]),.dout(n999),.clk(gclk));
	jor g0358(.dina(n999),.dinb(w_n988_0[1]),.dout(n1000),.clk(gclk));
	jor g0359(.dina(n1000),.dinb(n983),.dout(n1001),.clk(gclk));
	jnot g0360(.din(w_n1001_0[1]),.dout(n1002),.clk(gclk));
	jand g0361(.dina(n1002),.dinb(n975),.dout(n1003),.clk(gclk));
	jnot g0362(.din(w_in355_0[1]),.dout(n1004),.clk(gclk));
	jand g0363(.dina(n1004),.dinb(w_in255_0[1]),.dout(n1005),.clk(gclk));
	jnot g0364(.din(w_n988_0[0]),.dout(n1006),.clk(gclk));
	jnot g0365(.din(w_in351_0[1]),.dout(n1007),.clk(gclk));
	jand g0366(.dina(n1007),.dinb(w_in251_0[1]),.dout(n1008),.clk(gclk));
	jnot g0367(.din(w_n993_0[0]),.dout(n1009),.clk(gclk));
	jnot g0368(.din(w_n997_0[0]),.dout(n1010),.clk(gclk));
	jnot g0369(.din(w_in348_0[1]),.dout(n1011),.clk(gclk));
	jand g0370(.dina(n1011),.dinb(w_in248_0[1]),.dout(n1012),.clk(gclk));
	jand g0371(.dina(n1012),.dinb(n1010),.dout(n1013),.clk(gclk));
	jnot g0372(.din(w_in349_0[1]),.dout(n1014),.clk(gclk));
	jand g0373(.dina(n1014),.dinb(w_in249_0[1]),.dout(n1015),.clk(gclk));
	jnot g0374(.din(w_in350_0[1]),.dout(n1016),.clk(gclk));
	jand g0375(.dina(n1016),.dinb(w_in250_0[1]),.dout(n1017),.clk(gclk));
	jor g0376(.dina(n1017),.dinb(n1015),.dout(n1018),.clk(gclk));
	jor g0377(.dina(n1018),.dinb(n1013),.dout(n1019),.clk(gclk));
	jand g0378(.dina(n1019),.dinb(n1009),.dout(n1020),.clk(gclk));
	jor g0379(.dina(n1020),.dinb(n1008),.dout(n1021),.clk(gclk));
	jand g0380(.dina(n1021),.dinb(w_n982_0[0]),.dout(n1022),.clk(gclk));
	jand g0381(.dina(w_n980_0[0]),.dinb(w_in252_0[1]),.dout(n1023),.clk(gclk));
	jnot g0382(.din(w_in353_0[1]),.dout(n1024),.clk(gclk));
	jand g0383(.dina(n1024),.dinb(w_in253_0[1]),.dout(n1025),.clk(gclk));
	jnot g0384(.din(w_in354_0[1]),.dout(n1026),.clk(gclk));
	jand g0385(.dina(n1026),.dinb(w_in254_0[1]),.dout(n1027),.clk(gclk));
	jor g0386(.dina(n1027),.dinb(n1025),.dout(n1028),.clk(gclk));
	jor g0387(.dina(n1028),.dinb(n1023),.dout(n1029),.clk(gclk));
	jor g0388(.dina(n1029),.dinb(n1022),.dout(n1030),.clk(gclk));
	jand g0389(.dina(n1030),.dinb(n1006),.dout(n1031),.clk(gclk));
	jor g0390(.dina(n1031),.dinb(n1005),.dout(n1032),.clk(gclk));
	jor g0391(.dina(w_n1032_0[1]),.dinb(n1003),.dout(n1033),.clk(gclk));
	jnot g0392(.din(w_in261_0[2]),.dout(n1034),.clk(gclk));
	jand g0393(.dina(w_in361_0[2]),.dinb(n1034),.dout(n1035),.clk(gclk));
	jnot g0394(.din(w_in263_0[2]),.dout(n1036),.clk(gclk));
	jand g0395(.dina(w_in363_0[2]),.dinb(n1036),.dout(n1037),.clk(gclk));
	jnot g0396(.din(w_in262_0[2]),.dout(n1038),.clk(gclk));
	jand g0397(.dina(w_in362_0[2]),.dinb(n1038),.dout(n1039),.clk(gclk));
	jor g0398(.dina(n1039),.dinb(w_n1037_0[1]),.dout(n1040),.clk(gclk));
	jor g0399(.dina(n1040),.dinb(n1035),.dout(n1041),.clk(gclk));
	jnot g0400(.din(w_in259_0[2]),.dout(n1042),.clk(gclk));
	jand g0401(.dina(w_in359_0[2]),.dinb(n1042),.dout(n1043),.clk(gclk));
	jnot g0402(.din(w_in258_0[2]),.dout(n1044),.clk(gclk));
	jand g0403(.dina(w_in358_0[2]),.dinb(n1044),.dout(n1045),.clk(gclk));
	jor g0404(.dina(n1045),.dinb(n1043),.dout(n1046),.clk(gclk));
	jnot g0405(.din(w_in260_0[2]),.dout(n1047),.clk(gclk));
	jand g0406(.dina(w_in360_0[2]),.dinb(n1047),.dout(n1048),.clk(gclk));
	jnot g0407(.din(w_in256_0[2]),.dout(n1049),.clk(gclk));
	jand g0408(.dina(w_in356_0[2]),.dinb(n1049),.dout(n1050),.clk(gclk));
	jnot g0409(.din(w_in257_0[2]),.dout(n1051),.clk(gclk));
	jand g0410(.dina(w_in357_0[2]),.dinb(n1051),.dout(n1052),.clk(gclk));
	jor g0411(.dina(w_n1052_0[1]),.dinb(n1050),.dout(n1053),.clk(gclk));
	jor g0412(.dina(n1053),.dinb(w_n1048_0[1]),.dout(n1054),.clk(gclk));
	jor g0413(.dina(n1054),.dinb(w_n1046_0[1]),.dout(n1055),.clk(gclk));
	jor g0414(.dina(n1055),.dinb(w_n1041_0[1]),.dout(n1056),.clk(gclk));
	jnot g0415(.din(w_n1056_0[1]),.dout(n1057),.clk(gclk));
	jand g0416(.dina(n1057),.dinb(n1033),.dout(n1058),.clk(gclk));
	jnot g0417(.din(w_n1041_0[0]),.dout(n1059),.clk(gclk));
	jnot g0418(.din(w_n1048_0[0]),.dout(n1060),.clk(gclk));
	jnot g0419(.din(w_in359_0[1]),.dout(n1061),.clk(gclk));
	jand g0420(.dina(n1061),.dinb(w_in259_0[1]),.dout(n1062),.clk(gclk));
	jnot g0421(.din(w_n1046_0[0]),.dout(n1063),.clk(gclk));
	jnot g0422(.din(w_n1052_0[0]),.dout(n1064),.clk(gclk));
	jnot g0423(.din(w_in356_0[1]),.dout(n1065),.clk(gclk));
	jand g0424(.dina(n1065),.dinb(w_in256_0[1]),.dout(n1066),.clk(gclk));
	jand g0425(.dina(n1066),.dinb(n1064),.dout(n1067),.clk(gclk));
	jnot g0426(.din(w_in357_0[1]),.dout(n1068),.clk(gclk));
	jand g0427(.dina(n1068),.dinb(w_in257_0[1]),.dout(n1069),.clk(gclk));
	jnot g0428(.din(w_in358_0[1]),.dout(n1070),.clk(gclk));
	jand g0429(.dina(n1070),.dinb(w_in258_0[1]),.dout(n1071),.clk(gclk));
	jor g0430(.dina(n1071),.dinb(n1069),.dout(n1072),.clk(gclk));
	jor g0431(.dina(n1072),.dinb(n1067),.dout(n1073),.clk(gclk));
	jand g0432(.dina(n1073),.dinb(n1063),.dout(n1074),.clk(gclk));
	jor g0433(.dina(n1074),.dinb(n1062),.dout(n1075),.clk(gclk));
	jand g0434(.dina(n1075),.dinb(n1060),.dout(n1076),.clk(gclk));
	jnot g0435(.din(w_in360_0[1]),.dout(n1077),.clk(gclk));
	jand g0436(.dina(n1077),.dinb(w_in260_0[1]),.dout(n1078),.clk(gclk));
	jnot g0437(.din(w_in361_0[1]),.dout(n1079),.clk(gclk));
	jand g0438(.dina(n1079),.dinb(w_in261_0[1]),.dout(n1080),.clk(gclk));
	jor g0439(.dina(n1080),.dinb(n1078),.dout(n1081),.clk(gclk));
	jor g0440(.dina(n1081),.dinb(n1076),.dout(n1082),.clk(gclk));
	jand g0441(.dina(n1082),.dinb(n1059),.dout(n1083),.clk(gclk));
	jnot g0442(.din(w_n1037_0[0]),.dout(n1084),.clk(gclk));
	jnot g0443(.din(w_in362_0[1]),.dout(n1085),.clk(gclk));
	jand g0444(.dina(n1085),.dinb(w_in262_0[1]),.dout(n1086),.clk(gclk));
	jand g0445(.dina(n1086),.dinb(n1084),.dout(n1087),.clk(gclk));
	jnot g0446(.din(w_in363_0[1]),.dout(n1088),.clk(gclk));
	jand g0447(.dina(n1088),.dinb(w_in263_0[1]),.dout(n1089),.clk(gclk));
	jor g0448(.dina(n1089),.dinb(n1087),.dout(n1090),.clk(gclk));
	jor g0449(.dina(n1090),.dinb(n1083),.dout(n1091),.clk(gclk));
	jor g0450(.dina(w_n1091_0[1]),.dinb(n1058),.dout(n1092),.clk(gclk));
	jnot g0451(.din(w_in267_0[2]),.dout(n1093),.clk(gclk));
	jand g0452(.dina(w_in367_0[2]),.dinb(n1093),.dout(n1094),.clk(gclk));
	jnot g0453(.din(w_in266_0[2]),.dout(n1095),.clk(gclk));
	jand g0454(.dina(w_in366_0[2]),.dinb(n1095),.dout(n1096),.clk(gclk));
	jor g0455(.dina(n1096),.dinb(n1094),.dout(n1097),.clk(gclk));
	jnot g0456(.din(w_in265_0[2]),.dout(n1098),.clk(gclk));
	jand g0457(.dina(w_in365_0[2]),.dinb(n1098),.dout(n1099),.clk(gclk));
	jnot g0458(.din(w_in264_0[2]),.dout(n1100),.clk(gclk));
	jand g0459(.dina(w_in364_0[2]),.dinb(n1100),.dout(n1101),.clk(gclk));
	jor g0460(.dina(n1101),.dinb(w_n1099_0[1]),.dout(n1102),.clk(gclk));
	jor g0461(.dina(n1102),.dinb(w_n1097_0[1]),.dout(n1103),.clk(gclk));
	jnot g0462(.din(w_n1103_0[1]),.dout(n1104),.clk(gclk));
	jand g0463(.dina(n1104),.dinb(n1092),.dout(n1105),.clk(gclk));
	jnot g0464(.din(w_in367_0[1]),.dout(n1106),.clk(gclk));
	jand g0465(.dina(n1106),.dinb(w_in267_0[1]),.dout(n1107),.clk(gclk));
	jnot g0466(.din(w_n1097_0[0]),.dout(n1108),.clk(gclk));
	jnot g0467(.din(w_n1099_0[0]),.dout(n1109),.clk(gclk));
	jnot g0468(.din(w_in364_0[1]),.dout(n1110),.clk(gclk));
	jand g0469(.dina(n1110),.dinb(w_in264_0[1]),.dout(n1111),.clk(gclk));
	jand g0470(.dina(n1111),.dinb(n1109),.dout(n1112),.clk(gclk));
	jnot g0471(.din(w_in365_0[1]),.dout(n1113),.clk(gclk));
	jand g0472(.dina(n1113),.dinb(w_in265_0[1]),.dout(n1114),.clk(gclk));
	jnot g0473(.din(w_in366_0[1]),.dout(n1115),.clk(gclk));
	jand g0474(.dina(n1115),.dinb(w_in266_0[1]),.dout(n1116),.clk(gclk));
	jor g0475(.dina(n1116),.dinb(n1114),.dout(n1117),.clk(gclk));
	jor g0476(.dina(n1117),.dinb(n1112),.dout(n1118),.clk(gclk));
	jand g0477(.dina(n1118),.dinb(n1108),.dout(n1119),.clk(gclk));
	jor g0478(.dina(n1119),.dinb(n1107),.dout(n1120),.clk(gclk));
	jor g0479(.dina(w_n1120_0[1]),.dinb(n1105),.dout(n1121),.clk(gclk));
	jnot g0480(.din(w_in268_0[2]),.dout(n1122),.clk(gclk));
	jand g0481(.dina(w_in368_0[2]),.dinb(n1122),.dout(n1123),.clk(gclk));
	jnot g0482(.din(w_in269_0[2]),.dout(n1124),.clk(gclk));
	jand g0483(.dina(w_in369_0[2]),.dinb(n1124),.dout(n1125),.clk(gclk));
	jnot g0484(.din(w_in271_0[2]),.dout(n1126),.clk(gclk));
	jand g0485(.dina(w_in371_0[2]),.dinb(n1126),.dout(n1127),.clk(gclk));
	jnot g0486(.din(w_in270_0[2]),.dout(n1128),.clk(gclk));
	jand g0487(.dina(w_in370_0[2]),.dinb(n1128),.dout(n1129),.clk(gclk));
	jor g0488(.dina(n1129),.dinb(w_n1127_0[1]),.dout(n1130),.clk(gclk));
	jor g0489(.dina(n1130),.dinb(n1125),.dout(n1131),.clk(gclk));
	jor g0490(.dina(w_n1131_0[1]),.dinb(n1123),.dout(n1132),.clk(gclk));
	jnot g0491(.din(w_n1132_0[1]),.dout(n1133),.clk(gclk));
	jand g0492(.dina(n1133),.dinb(n1121),.dout(n1134),.clk(gclk));
	jnot g0493(.din(w_n1131_0[0]),.dout(n1135),.clk(gclk));
	jnot g0494(.din(w_in369_0[1]),.dout(n1136),.clk(gclk));
	jand g0495(.dina(n1136),.dinb(w_in269_0[1]),.dout(n1137),.clk(gclk));
	jnot g0496(.din(w_in368_0[1]),.dout(n1138),.clk(gclk));
	jand g0497(.dina(n1138),.dinb(w_in268_0[1]),.dout(n1139),.clk(gclk));
	jor g0498(.dina(n1139),.dinb(n1137),.dout(n1140),.clk(gclk));
	jand g0499(.dina(n1140),.dinb(n1135),.dout(n1141),.clk(gclk));
	jnot g0500(.din(w_in371_0[1]),.dout(n1142),.clk(gclk));
	jand g0501(.dina(n1142),.dinb(w_in271_0[1]),.dout(n1143),.clk(gclk));
	jnot g0502(.din(w_n1127_0[0]),.dout(n1144),.clk(gclk));
	jnot g0503(.din(w_in370_0[1]),.dout(n1145),.clk(gclk));
	jand g0504(.dina(n1145),.dinb(w_in270_0[1]),.dout(n1146),.clk(gclk));
	jand g0505(.dina(n1146),.dinb(n1144),.dout(n1147),.clk(gclk));
	jor g0506(.dina(n1147),.dinb(n1143),.dout(n1148),.clk(gclk));
	jor g0507(.dina(n1148),.dinb(n1141),.dout(n1149),.clk(gclk));
	jor g0508(.dina(w_n1149_0[1]),.dinb(n1134),.dout(n1150),.clk(gclk));
	jnot g0509(.din(w_in275_0[2]),.dout(n1151),.clk(gclk));
	jand g0510(.dina(w_in375_0[2]),.dinb(n1151),.dout(n1152),.clk(gclk));
	jnot g0511(.din(w_in274_0[2]),.dout(n1153),.clk(gclk));
	jand g0512(.dina(w_in374_0[2]),.dinb(n1153),.dout(n1154),.clk(gclk));
	jor g0513(.dina(n1154),.dinb(n1152),.dout(n1155),.clk(gclk));
	jnot g0514(.din(w_in273_0[2]),.dout(n1156),.clk(gclk));
	jand g0515(.dina(w_in373_0[2]),.dinb(n1156),.dout(n1157),.clk(gclk));
	jnot g0516(.din(w_in272_0[2]),.dout(n1158),.clk(gclk));
	jand g0517(.dina(w_in372_0[2]),.dinb(n1158),.dout(n1159),.clk(gclk));
	jor g0518(.dina(n1159),.dinb(w_n1157_0[1]),.dout(n1160),.clk(gclk));
	jor g0519(.dina(n1160),.dinb(w_n1155_0[1]),.dout(n1161),.clk(gclk));
	jnot g0520(.din(w_n1161_0[1]),.dout(n1162),.clk(gclk));
	jand g0521(.dina(n1162),.dinb(n1150),.dout(n1163),.clk(gclk));
	jnot g0522(.din(w_in375_0[1]),.dout(n1164),.clk(gclk));
	jand g0523(.dina(n1164),.dinb(w_in275_0[1]),.dout(n1165),.clk(gclk));
	jnot g0524(.din(w_n1155_0[0]),.dout(n1166),.clk(gclk));
	jnot g0525(.din(w_n1157_0[0]),.dout(n1167),.clk(gclk));
	jnot g0526(.din(w_in372_0[1]),.dout(n1168),.clk(gclk));
	jand g0527(.dina(n1168),.dinb(w_in272_0[1]),.dout(n1169),.clk(gclk));
	jand g0528(.dina(n1169),.dinb(n1167),.dout(n1170),.clk(gclk));
	jnot g0529(.din(w_in373_0[1]),.dout(n1171),.clk(gclk));
	jand g0530(.dina(n1171),.dinb(w_in273_0[1]),.dout(n1172),.clk(gclk));
	jnot g0531(.din(w_in374_0[1]),.dout(n1173),.clk(gclk));
	jand g0532(.dina(n1173),.dinb(w_in274_0[1]),.dout(n1174),.clk(gclk));
	jor g0533(.dina(n1174),.dinb(n1172),.dout(n1175),.clk(gclk));
	jor g0534(.dina(n1175),.dinb(n1170),.dout(n1176),.clk(gclk));
	jand g0535(.dina(n1176),.dinb(n1166),.dout(n1177),.clk(gclk));
	jor g0536(.dina(n1177),.dinb(n1165),.dout(n1178),.clk(gclk));
	jor g0537(.dina(w_n1178_0[1]),.dinb(n1163),.dout(n1179),.clk(gclk));
	jnot g0538(.din(w_in276_0[2]),.dout(n1180),.clk(gclk));
	jand g0539(.dina(w_in376_0[2]),.dinb(n1180),.dout(n1181),.clk(gclk));
	jnot g0540(.din(w_in277_0[2]),.dout(n1182),.clk(gclk));
	jand g0541(.dina(w_in377_0[2]),.dinb(n1182),.dout(n1183),.clk(gclk));
	jnot g0542(.din(w_in279_0[2]),.dout(n1184),.clk(gclk));
	jand g0543(.dina(w_in379_0[2]),.dinb(n1184),.dout(n1185),.clk(gclk));
	jnot g0544(.din(w_in278_0[2]),.dout(n1186),.clk(gclk));
	jand g0545(.dina(w_in378_0[2]),.dinb(n1186),.dout(n1187),.clk(gclk));
	jor g0546(.dina(n1187),.dinb(w_n1185_0[1]),.dout(n1188),.clk(gclk));
	jor g0547(.dina(n1188),.dinb(n1183),.dout(n1189),.clk(gclk));
	jor g0548(.dina(w_n1189_0[1]),.dinb(n1181),.dout(n1190),.clk(gclk));
	jnot g0549(.din(w_n1190_0[1]),.dout(n1191),.clk(gclk));
	jand g0550(.dina(n1191),.dinb(n1179),.dout(n1192),.clk(gclk));
	jnot g0551(.din(w_n1189_0[0]),.dout(n1193),.clk(gclk));
	jnot g0552(.din(w_in377_0[1]),.dout(n1194),.clk(gclk));
	jand g0553(.dina(n1194),.dinb(w_in277_0[1]),.dout(n1195),.clk(gclk));
	jnot g0554(.din(w_in376_0[1]),.dout(n1196),.clk(gclk));
	jand g0555(.dina(n1196),.dinb(w_in276_0[1]),.dout(n1197),.clk(gclk));
	jor g0556(.dina(n1197),.dinb(n1195),.dout(n1198),.clk(gclk));
	jand g0557(.dina(n1198),.dinb(n1193),.dout(n1199),.clk(gclk));
	jnot g0558(.din(w_in379_0[1]),.dout(n1200),.clk(gclk));
	jand g0559(.dina(n1200),.dinb(w_in279_0[1]),.dout(n1201),.clk(gclk));
	jnot g0560(.din(w_n1185_0[0]),.dout(n1202),.clk(gclk));
	jnot g0561(.din(w_in378_0[1]),.dout(n1203),.clk(gclk));
	jand g0562(.dina(n1203),.dinb(w_in278_0[1]),.dout(n1204),.clk(gclk));
	jand g0563(.dina(n1204),.dinb(n1202),.dout(n1205),.clk(gclk));
	jor g0564(.dina(n1205),.dinb(n1201),.dout(n1206),.clk(gclk));
	jor g0565(.dina(n1206),.dinb(n1199),.dout(n1207),.clk(gclk));
	jor g0566(.dina(w_n1207_0[1]),.dinb(n1192),.dout(n1208),.clk(gclk));
	jnot g0567(.din(w_in283_0[2]),.dout(n1209),.clk(gclk));
	jand g0568(.dina(w_in383_0[2]),.dinb(n1209),.dout(n1210),.clk(gclk));
	jnot g0569(.din(w_in282_0[2]),.dout(n1211),.clk(gclk));
	jand g0570(.dina(w_in382_0[2]),.dinb(n1211),.dout(n1212),.clk(gclk));
	jor g0571(.dina(n1212),.dinb(n1210),.dout(n1213),.clk(gclk));
	jnot g0572(.din(w_in281_0[2]),.dout(n1214),.clk(gclk));
	jand g0573(.dina(w_in381_0[2]),.dinb(n1214),.dout(n1215),.clk(gclk));
	jnot g0574(.din(w_in280_0[2]),.dout(n1216),.clk(gclk));
	jand g0575(.dina(w_in380_0[2]),.dinb(n1216),.dout(n1217),.clk(gclk));
	jor g0576(.dina(n1217),.dinb(w_n1215_0[1]),.dout(n1218),.clk(gclk));
	jor g0577(.dina(n1218),.dinb(w_n1213_0[1]),.dout(n1219),.clk(gclk));
	jnot g0578(.din(w_n1219_0[1]),.dout(n1220),.clk(gclk));
	jand g0579(.dina(n1220),.dinb(n1208),.dout(n1221),.clk(gclk));
	jnot g0580(.din(w_in383_0[1]),.dout(n1222),.clk(gclk));
	jand g0581(.dina(n1222),.dinb(w_in283_0[1]),.dout(n1223),.clk(gclk));
	jnot g0582(.din(w_n1213_0[0]),.dout(n1224),.clk(gclk));
	jnot g0583(.din(w_n1215_0[0]),.dout(n1225),.clk(gclk));
	jnot g0584(.din(w_in380_0[1]),.dout(n1226),.clk(gclk));
	jand g0585(.dina(n1226),.dinb(w_in280_0[1]),.dout(n1227),.clk(gclk));
	jand g0586(.dina(n1227),.dinb(n1225),.dout(n1228),.clk(gclk));
	jnot g0587(.din(w_in381_0[1]),.dout(n1229),.clk(gclk));
	jand g0588(.dina(n1229),.dinb(w_in281_0[1]),.dout(n1230),.clk(gclk));
	jnot g0589(.din(w_in382_0[1]),.dout(n1231),.clk(gclk));
	jand g0590(.dina(n1231),.dinb(w_in282_0[1]),.dout(n1232),.clk(gclk));
	jor g0591(.dina(n1232),.dinb(n1230),.dout(n1233),.clk(gclk));
	jor g0592(.dina(n1233),.dinb(n1228),.dout(n1234),.clk(gclk));
	jand g0593(.dina(n1234),.dinb(n1224),.dout(n1235),.clk(gclk));
	jor g0594(.dina(n1235),.dinb(n1223),.dout(n1236),.clk(gclk));
	jor g0595(.dina(w_n1236_0[1]),.dinb(n1221),.dout(n1237),.clk(gclk));
	jnot g0596(.din(w_in284_0[2]),.dout(n1238),.clk(gclk));
	jand g0597(.dina(w_in384_0[2]),.dinb(n1238),.dout(n1239),.clk(gclk));
	jnot g0598(.din(w_in285_0[2]),.dout(n1240),.clk(gclk));
	jand g0599(.dina(w_in385_0[2]),.dinb(n1240),.dout(n1241),.clk(gclk));
	jnot g0600(.din(w_in287_0[2]),.dout(n1242),.clk(gclk));
	jand g0601(.dina(w_in387_0[2]),.dinb(n1242),.dout(n1243),.clk(gclk));
	jnot g0602(.din(w_in286_0[2]),.dout(n1244),.clk(gclk));
	jand g0603(.dina(w_in386_0[2]),.dinb(n1244),.dout(n1245),.clk(gclk));
	jor g0604(.dina(n1245),.dinb(w_n1243_0[1]),.dout(n1246),.clk(gclk));
	jor g0605(.dina(n1246),.dinb(n1241),.dout(n1247),.clk(gclk));
	jor g0606(.dina(w_n1247_0[1]),.dinb(n1239),.dout(n1248),.clk(gclk));
	jnot g0607(.din(w_n1248_0[1]),.dout(n1249),.clk(gclk));
	jand g0608(.dina(n1249),.dinb(n1237),.dout(n1250),.clk(gclk));
	jnot g0609(.din(w_n1247_0[0]),.dout(n1251),.clk(gclk));
	jnot g0610(.din(w_in385_0[1]),.dout(n1252),.clk(gclk));
	jand g0611(.dina(n1252),.dinb(w_in285_0[1]),.dout(n1253),.clk(gclk));
	jnot g0612(.din(w_in384_0[1]),.dout(n1254),.clk(gclk));
	jand g0613(.dina(n1254),.dinb(w_in284_0[1]),.dout(n1255),.clk(gclk));
	jor g0614(.dina(n1255),.dinb(n1253),.dout(n1256),.clk(gclk));
	jand g0615(.dina(n1256),.dinb(n1251),.dout(n1257),.clk(gclk));
	jnot g0616(.din(w_in387_0[1]),.dout(n1258),.clk(gclk));
	jand g0617(.dina(n1258),.dinb(w_in287_0[1]),.dout(n1259),.clk(gclk));
	jnot g0618(.din(w_n1243_0[0]),.dout(n1260),.clk(gclk));
	jnot g0619(.din(w_in386_0[1]),.dout(n1261),.clk(gclk));
	jand g0620(.dina(n1261),.dinb(w_in286_0[1]),.dout(n1262),.clk(gclk));
	jand g0621(.dina(n1262),.dinb(n1260),.dout(n1263),.clk(gclk));
	jor g0622(.dina(n1263),.dinb(n1259),.dout(n1264),.clk(gclk));
	jor g0623(.dina(n1264),.dinb(n1257),.dout(n1265),.clk(gclk));
	jor g0624(.dina(w_n1265_0[1]),.dinb(n1250),.dout(n1266),.clk(gclk));
	jnot g0625(.din(w_in291_0[2]),.dout(n1267),.clk(gclk));
	jand g0626(.dina(w_in391_0[2]),.dinb(n1267),.dout(n1268),.clk(gclk));
	jnot g0627(.din(w_in290_0[2]),.dout(n1269),.clk(gclk));
	jand g0628(.dina(w_in390_0[2]),.dinb(n1269),.dout(n1270),.clk(gclk));
	jor g0629(.dina(n1270),.dinb(n1268),.dout(n1271),.clk(gclk));
	jnot g0630(.din(w_in289_0[2]),.dout(n1272),.clk(gclk));
	jand g0631(.dina(w_in389_0[2]),.dinb(n1272),.dout(n1273),.clk(gclk));
	jnot g0632(.din(w_in288_0[2]),.dout(n1274),.clk(gclk));
	jand g0633(.dina(w_in388_0[2]),.dinb(n1274),.dout(n1275),.clk(gclk));
	jor g0634(.dina(n1275),.dinb(w_n1273_0[1]),.dout(n1276),.clk(gclk));
	jor g0635(.dina(n1276),.dinb(w_n1271_0[1]),.dout(n1277),.clk(gclk));
	jnot g0636(.din(w_n1277_0[1]),.dout(n1278),.clk(gclk));
	jand g0637(.dina(n1278),.dinb(n1266),.dout(n1279),.clk(gclk));
	jnot g0638(.din(w_in391_0[1]),.dout(n1280),.clk(gclk));
	jand g0639(.dina(n1280),.dinb(w_in291_0[1]),.dout(n1281),.clk(gclk));
	jnot g0640(.din(w_n1271_0[0]),.dout(n1282),.clk(gclk));
	jnot g0641(.din(w_n1273_0[0]),.dout(n1283),.clk(gclk));
	jnot g0642(.din(w_in388_0[1]),.dout(n1284),.clk(gclk));
	jand g0643(.dina(n1284),.dinb(w_in288_0[1]),.dout(n1285),.clk(gclk));
	jand g0644(.dina(n1285),.dinb(n1283),.dout(n1286),.clk(gclk));
	jnot g0645(.din(w_in389_0[1]),.dout(n1287),.clk(gclk));
	jand g0646(.dina(n1287),.dinb(w_in289_0[1]),.dout(n1288),.clk(gclk));
	jnot g0647(.din(w_in390_0[1]),.dout(n1289),.clk(gclk));
	jand g0648(.dina(n1289),.dinb(w_in290_0[1]),.dout(n1290),.clk(gclk));
	jor g0649(.dina(n1290),.dinb(n1288),.dout(n1291),.clk(gclk));
	jor g0650(.dina(n1291),.dinb(n1286),.dout(n1292),.clk(gclk));
	jand g0651(.dina(n1292),.dinb(n1282),.dout(n1293),.clk(gclk));
	jor g0652(.dina(n1293),.dinb(n1281),.dout(n1294),.clk(gclk));
	jor g0653(.dina(w_n1294_0[1]),.dinb(n1279),.dout(n1295),.clk(gclk));
	jnot g0654(.din(w_in292_0[2]),.dout(n1296),.clk(gclk));
	jand g0655(.dina(w_in392_0[2]),.dinb(n1296),.dout(n1297),.clk(gclk));
	jnot g0656(.din(w_in293_0[2]),.dout(n1298),.clk(gclk));
	jand g0657(.dina(w_in393_0[2]),.dinb(n1298),.dout(n1299),.clk(gclk));
	jnot g0658(.din(w_in295_0[2]),.dout(n1300),.clk(gclk));
	jand g0659(.dina(w_in395_0[2]),.dinb(n1300),.dout(n1301),.clk(gclk));
	jnot g0660(.din(w_in294_0[2]),.dout(n1302),.clk(gclk));
	jand g0661(.dina(w_in394_0[2]),.dinb(n1302),.dout(n1303),.clk(gclk));
	jor g0662(.dina(n1303),.dinb(w_n1301_0[1]),.dout(n1304),.clk(gclk));
	jor g0663(.dina(n1304),.dinb(n1299),.dout(n1305),.clk(gclk));
	jor g0664(.dina(w_n1305_0[1]),.dinb(n1297),.dout(n1306),.clk(gclk));
	jnot g0665(.din(w_n1306_0[1]),.dout(n1307),.clk(gclk));
	jand g0666(.dina(n1307),.dinb(n1295),.dout(n1308),.clk(gclk));
	jnot g0667(.din(w_n1305_0[0]),.dout(n1309),.clk(gclk));
	jnot g0668(.din(w_in393_0[1]),.dout(n1310),.clk(gclk));
	jand g0669(.dina(n1310),.dinb(w_in293_0[1]),.dout(n1311),.clk(gclk));
	jnot g0670(.din(w_in392_0[1]),.dout(n1312),.clk(gclk));
	jand g0671(.dina(n1312),.dinb(w_in292_0[1]),.dout(n1313),.clk(gclk));
	jor g0672(.dina(n1313),.dinb(n1311),.dout(n1314),.clk(gclk));
	jand g0673(.dina(n1314),.dinb(n1309),.dout(n1315),.clk(gclk));
	jnot g0674(.din(w_in395_0[1]),.dout(n1316),.clk(gclk));
	jand g0675(.dina(n1316),.dinb(w_in295_0[1]),.dout(n1317),.clk(gclk));
	jnot g0676(.din(w_n1301_0[0]),.dout(n1318),.clk(gclk));
	jnot g0677(.din(w_in394_0[1]),.dout(n1319),.clk(gclk));
	jand g0678(.dina(n1319),.dinb(w_in294_0[1]),.dout(n1320),.clk(gclk));
	jand g0679(.dina(n1320),.dinb(n1318),.dout(n1321),.clk(gclk));
	jor g0680(.dina(n1321),.dinb(n1317),.dout(n1322),.clk(gclk));
	jor g0681(.dina(n1322),.dinb(n1315),.dout(n1323),.clk(gclk));
	jor g0682(.dina(w_n1323_0[1]),.dinb(n1308),.dout(n1324),.clk(gclk));
	jnot g0683(.din(w_in299_0[2]),.dout(n1325),.clk(gclk));
	jand g0684(.dina(w_in399_0[2]),.dinb(n1325),.dout(n1326),.clk(gclk));
	jnot g0685(.din(w_in298_0[2]),.dout(n1327),.clk(gclk));
	jand g0686(.dina(w_in398_0[2]),.dinb(n1327),.dout(n1328),.clk(gclk));
	jor g0687(.dina(n1328),.dinb(n1326),.dout(n1329),.clk(gclk));
	jnot g0688(.din(w_in297_0[2]),.dout(n1330),.clk(gclk));
	jand g0689(.dina(w_in397_0[2]),.dinb(n1330),.dout(n1331),.clk(gclk));
	jnot g0690(.din(w_in296_0[2]),.dout(n1332),.clk(gclk));
	jand g0691(.dina(w_in396_0[2]),.dinb(n1332),.dout(n1333),.clk(gclk));
	jor g0692(.dina(n1333),.dinb(w_n1331_0[1]),.dout(n1334),.clk(gclk));
	jor g0693(.dina(n1334),.dinb(w_n1329_0[1]),.dout(n1335),.clk(gclk));
	jnot g0694(.din(w_n1335_0[1]),.dout(n1336),.clk(gclk));
	jand g0695(.dina(n1336),.dinb(n1324),.dout(n1337),.clk(gclk));
	jnot g0696(.din(w_in399_0[1]),.dout(n1338),.clk(gclk));
	jand g0697(.dina(n1338),.dinb(w_in299_0[1]),.dout(n1339),.clk(gclk));
	jnot g0698(.din(w_n1329_0[0]),.dout(n1340),.clk(gclk));
	jnot g0699(.din(w_n1331_0[0]),.dout(n1341),.clk(gclk));
	jnot g0700(.din(w_in396_0[1]),.dout(n1342),.clk(gclk));
	jand g0701(.dina(n1342),.dinb(w_in296_0[1]),.dout(n1343),.clk(gclk));
	jand g0702(.dina(n1343),.dinb(n1341),.dout(n1344),.clk(gclk));
	jnot g0703(.din(w_in397_0[1]),.dout(n1345),.clk(gclk));
	jand g0704(.dina(n1345),.dinb(w_in297_0[1]),.dout(n1346),.clk(gclk));
	jnot g0705(.din(w_in398_0[1]),.dout(n1347),.clk(gclk));
	jand g0706(.dina(n1347),.dinb(w_in298_0[1]),.dout(n1348),.clk(gclk));
	jor g0707(.dina(n1348),.dinb(n1346),.dout(n1349),.clk(gclk));
	jor g0708(.dina(n1349),.dinb(n1344),.dout(n1350),.clk(gclk));
	jand g0709(.dina(n1350),.dinb(n1340),.dout(n1351),.clk(gclk));
	jor g0710(.dina(n1351),.dinb(n1339),.dout(n1352),.clk(gclk));
	jor g0711(.dina(w_n1352_0[1]),.dinb(n1337),.dout(n1353),.clk(gclk));
	jnot g0712(.din(w_in2100_0[2]),.dout(n1354),.clk(gclk));
	jand g0713(.dina(w_in3100_0[2]),.dinb(n1354),.dout(n1355),.clk(gclk));
	jnot g0714(.din(w_in2101_0[2]),.dout(n1356),.clk(gclk));
	jand g0715(.dina(w_in3101_0[2]),.dinb(n1356),.dout(n1357),.clk(gclk));
	jnot g0716(.din(w_in2103_0[2]),.dout(n1358),.clk(gclk));
	jand g0717(.dina(w_in3103_0[2]),.dinb(n1358),.dout(n1359),.clk(gclk));
	jnot g0718(.din(w_in2102_0[2]),.dout(n1360),.clk(gclk));
	jand g0719(.dina(w_in3102_0[2]),.dinb(n1360),.dout(n1361),.clk(gclk));
	jor g0720(.dina(n1361),.dinb(w_n1359_0[1]),.dout(n1362),.clk(gclk));
	jor g0721(.dina(n1362),.dinb(n1357),.dout(n1363),.clk(gclk));
	jor g0722(.dina(w_n1363_0[1]),.dinb(n1355),.dout(n1364),.clk(gclk));
	jnot g0723(.din(w_n1364_0[1]),.dout(n1365),.clk(gclk));
	jand g0724(.dina(n1365),.dinb(n1353),.dout(n1366),.clk(gclk));
	jnot g0725(.din(w_n1363_0[0]),.dout(n1367),.clk(gclk));
	jnot g0726(.din(w_in3101_0[1]),.dout(n1368),.clk(gclk));
	jand g0727(.dina(n1368),.dinb(w_in2101_0[1]),.dout(n1369),.clk(gclk));
	jnot g0728(.din(w_in3100_0[1]),.dout(n1370),.clk(gclk));
	jand g0729(.dina(n1370),.dinb(w_in2100_0[1]),.dout(n1371),.clk(gclk));
	jor g0730(.dina(n1371),.dinb(n1369),.dout(n1372),.clk(gclk));
	jand g0731(.dina(n1372),.dinb(n1367),.dout(n1373),.clk(gclk));
	jnot g0732(.din(w_in3103_0[1]),.dout(n1374),.clk(gclk));
	jand g0733(.dina(n1374),.dinb(w_in2103_0[1]),.dout(n1375),.clk(gclk));
	jnot g0734(.din(w_n1359_0[0]),.dout(n1376),.clk(gclk));
	jnot g0735(.din(w_in3102_0[1]),.dout(n1377),.clk(gclk));
	jand g0736(.dina(n1377),.dinb(w_in2102_0[1]),.dout(n1378),.clk(gclk));
	jand g0737(.dina(n1378),.dinb(n1376),.dout(n1379),.clk(gclk));
	jor g0738(.dina(n1379),.dinb(n1375),.dout(n1380),.clk(gclk));
	jor g0739(.dina(n1380),.dinb(n1373),.dout(n1381),.clk(gclk));
	jor g0740(.dina(w_n1381_0[1]),.dinb(n1366),.dout(n1382),.clk(gclk));
	jnot g0741(.din(w_in2107_0[2]),.dout(n1383),.clk(gclk));
	jand g0742(.dina(w_in3107_0[2]),.dinb(n1383),.dout(n1384),.clk(gclk));
	jnot g0743(.din(w_in2106_0[2]),.dout(n1385),.clk(gclk));
	jand g0744(.dina(w_in3106_0[2]),.dinb(n1385),.dout(n1386),.clk(gclk));
	jor g0745(.dina(n1386),.dinb(n1384),.dout(n1387),.clk(gclk));
	jnot g0746(.din(w_in2105_0[2]),.dout(n1388),.clk(gclk));
	jand g0747(.dina(w_in3105_0[2]),.dinb(n1388),.dout(n1389),.clk(gclk));
	jnot g0748(.din(w_in2104_0[2]),.dout(n1390),.clk(gclk));
	jand g0749(.dina(w_in3104_0[2]),.dinb(n1390),.dout(n1391),.clk(gclk));
	jor g0750(.dina(n1391),.dinb(w_n1389_0[1]),.dout(n1392),.clk(gclk));
	jor g0751(.dina(n1392),.dinb(w_n1387_0[1]),.dout(n1393),.clk(gclk));
	jnot g0752(.din(w_n1393_0[1]),.dout(n1394),.clk(gclk));
	jand g0753(.dina(n1394),.dinb(n1382),.dout(n1395),.clk(gclk));
	jnot g0754(.din(w_in3107_0[1]),.dout(n1396),.clk(gclk));
	jand g0755(.dina(n1396),.dinb(w_in2107_0[1]),.dout(n1397),.clk(gclk));
	jnot g0756(.din(w_n1387_0[0]),.dout(n1398),.clk(gclk));
	jnot g0757(.din(w_n1389_0[0]),.dout(n1399),.clk(gclk));
	jnot g0758(.din(w_in3104_0[1]),.dout(n1400),.clk(gclk));
	jand g0759(.dina(n1400),.dinb(w_in2104_0[1]),.dout(n1401),.clk(gclk));
	jand g0760(.dina(n1401),.dinb(n1399),.dout(n1402),.clk(gclk));
	jnot g0761(.din(w_in3105_0[1]),.dout(n1403),.clk(gclk));
	jand g0762(.dina(n1403),.dinb(w_in2105_0[1]),.dout(n1404),.clk(gclk));
	jnot g0763(.din(w_in3106_0[1]),.dout(n1405),.clk(gclk));
	jand g0764(.dina(n1405),.dinb(w_in2106_0[1]),.dout(n1406),.clk(gclk));
	jor g0765(.dina(n1406),.dinb(n1404),.dout(n1407),.clk(gclk));
	jor g0766(.dina(n1407),.dinb(n1402),.dout(n1408),.clk(gclk));
	jand g0767(.dina(n1408),.dinb(n1398),.dout(n1409),.clk(gclk));
	jor g0768(.dina(n1409),.dinb(n1397),.dout(n1410),.clk(gclk));
	jor g0769(.dina(w_n1410_0[1]),.dinb(n1395),.dout(n1411),.clk(gclk));
	jnot g0770(.din(w_in2108_0[2]),.dout(n1412),.clk(gclk));
	jand g0771(.dina(w_in3108_0[2]),.dinb(n1412),.dout(n1413),.clk(gclk));
	jnot g0772(.din(w_in2109_0[2]),.dout(n1414),.clk(gclk));
	jand g0773(.dina(w_in3109_0[2]),.dinb(n1414),.dout(n1415),.clk(gclk));
	jnot g0774(.din(w_in2111_0[2]),.dout(n1416),.clk(gclk));
	jand g0775(.dina(w_in3111_0[2]),.dinb(n1416),.dout(n1417),.clk(gclk));
	jnot g0776(.din(w_in2110_0[2]),.dout(n1418),.clk(gclk));
	jand g0777(.dina(w_in3110_0[2]),.dinb(n1418),.dout(n1419),.clk(gclk));
	jor g0778(.dina(n1419),.dinb(w_n1417_0[1]),.dout(n1420),.clk(gclk));
	jor g0779(.dina(n1420),.dinb(n1415),.dout(n1421),.clk(gclk));
	jor g0780(.dina(w_n1421_0[1]),.dinb(n1413),.dout(n1422),.clk(gclk));
	jnot g0781(.din(w_n1422_0[1]),.dout(n1423),.clk(gclk));
	jand g0782(.dina(n1423),.dinb(n1411),.dout(n1424),.clk(gclk));
	jnot g0783(.din(w_n1421_0[0]),.dout(n1425),.clk(gclk));
	jnot g0784(.din(w_in3109_0[1]),.dout(n1426),.clk(gclk));
	jand g0785(.dina(n1426),.dinb(w_in2109_0[1]),.dout(n1427),.clk(gclk));
	jnot g0786(.din(w_in3108_0[1]),.dout(n1428),.clk(gclk));
	jand g0787(.dina(n1428),.dinb(w_in2108_0[1]),.dout(n1429),.clk(gclk));
	jor g0788(.dina(n1429),.dinb(n1427),.dout(n1430),.clk(gclk));
	jand g0789(.dina(n1430),.dinb(n1425),.dout(n1431),.clk(gclk));
	jnot g0790(.din(w_in3111_0[1]),.dout(n1432),.clk(gclk));
	jand g0791(.dina(n1432),.dinb(w_in2111_0[1]),.dout(n1433),.clk(gclk));
	jnot g0792(.din(w_n1417_0[0]),.dout(n1434),.clk(gclk));
	jnot g0793(.din(w_in3110_0[1]),.dout(n1435),.clk(gclk));
	jand g0794(.dina(n1435),.dinb(w_in2110_0[1]),.dout(n1436),.clk(gclk));
	jand g0795(.dina(n1436),.dinb(n1434),.dout(n1437),.clk(gclk));
	jor g0796(.dina(n1437),.dinb(n1433),.dout(n1438),.clk(gclk));
	jor g0797(.dina(n1438),.dinb(n1431),.dout(n1439),.clk(gclk));
	jor g0798(.dina(w_n1439_0[1]),.dinb(n1424),.dout(n1440),.clk(gclk));
	jnot g0799(.din(w_in2115_0[2]),.dout(n1441),.clk(gclk));
	jand g0800(.dina(w_in3115_0[2]),.dinb(n1441),.dout(n1442),.clk(gclk));
	jnot g0801(.din(w_in2114_0[2]),.dout(n1443),.clk(gclk));
	jand g0802(.dina(w_in3114_0[2]),.dinb(n1443),.dout(n1444),.clk(gclk));
	jor g0803(.dina(n1444),.dinb(n1442),.dout(n1445),.clk(gclk));
	jnot g0804(.din(w_in2113_0[2]),.dout(n1446),.clk(gclk));
	jand g0805(.dina(w_in3113_0[2]),.dinb(n1446),.dout(n1447),.clk(gclk));
	jnot g0806(.din(w_in2112_0[2]),.dout(n1448),.clk(gclk));
	jand g0807(.dina(w_in3112_0[2]),.dinb(n1448),.dout(n1449),.clk(gclk));
	jor g0808(.dina(n1449),.dinb(w_n1447_0[1]),.dout(n1450),.clk(gclk));
	jor g0809(.dina(n1450),.dinb(w_n1445_0[1]),.dout(n1451),.clk(gclk));
	jnot g0810(.din(w_n1451_0[1]),.dout(n1452),.clk(gclk));
	jand g0811(.dina(n1452),.dinb(n1440),.dout(n1453),.clk(gclk));
	jnot g0812(.din(w_in3115_0[1]),.dout(n1454),.clk(gclk));
	jand g0813(.dina(n1454),.dinb(w_in2115_0[1]),.dout(n1455),.clk(gclk));
	jnot g0814(.din(w_n1445_0[0]),.dout(n1456),.clk(gclk));
	jnot g0815(.din(w_n1447_0[0]),.dout(n1457),.clk(gclk));
	jnot g0816(.din(w_in3112_0[1]),.dout(n1458),.clk(gclk));
	jand g0817(.dina(n1458),.dinb(w_in2112_0[1]),.dout(n1459),.clk(gclk));
	jand g0818(.dina(n1459),.dinb(n1457),.dout(n1460),.clk(gclk));
	jnot g0819(.din(w_in3113_0[1]),.dout(n1461),.clk(gclk));
	jand g0820(.dina(n1461),.dinb(w_in2113_0[1]),.dout(n1462),.clk(gclk));
	jnot g0821(.din(w_in3114_0[1]),.dout(n1463),.clk(gclk));
	jand g0822(.dina(n1463),.dinb(w_in2114_0[1]),.dout(n1464),.clk(gclk));
	jor g0823(.dina(n1464),.dinb(n1462),.dout(n1465),.clk(gclk));
	jor g0824(.dina(n1465),.dinb(n1460),.dout(n1466),.clk(gclk));
	jand g0825(.dina(n1466),.dinb(n1456),.dout(n1467),.clk(gclk));
	jor g0826(.dina(n1467),.dinb(n1455),.dout(n1468),.clk(gclk));
	jor g0827(.dina(w_n1468_0[1]),.dinb(n1453),.dout(n1469),.clk(gclk));
	jnot g0828(.din(w_in2116_0[2]),.dout(n1470),.clk(gclk));
	jand g0829(.dina(w_in3116_0[2]),.dinb(n1470),.dout(n1471),.clk(gclk));
	jnot g0830(.din(w_in2117_0[2]),.dout(n1472),.clk(gclk));
	jand g0831(.dina(w_in3117_0[2]),.dinb(n1472),.dout(n1473),.clk(gclk));
	jnot g0832(.din(w_in2119_0[2]),.dout(n1474),.clk(gclk));
	jand g0833(.dina(w_in3119_0[2]),.dinb(n1474),.dout(n1475),.clk(gclk));
	jnot g0834(.din(w_in2118_0[2]),.dout(n1476),.clk(gclk));
	jand g0835(.dina(w_in3118_0[2]),.dinb(n1476),.dout(n1477),.clk(gclk));
	jor g0836(.dina(n1477),.dinb(w_n1475_0[1]),.dout(n1478),.clk(gclk));
	jor g0837(.dina(n1478),.dinb(n1473),.dout(n1479),.clk(gclk));
	jor g0838(.dina(w_n1479_0[1]),.dinb(n1471),.dout(n1480),.clk(gclk));
	jnot g0839(.din(w_n1480_0[1]),.dout(n1481),.clk(gclk));
	jand g0840(.dina(n1481),.dinb(n1469),.dout(n1482),.clk(gclk));
	jnot g0841(.din(w_n1479_0[0]),.dout(n1483),.clk(gclk));
	jnot g0842(.din(w_in3117_0[1]),.dout(n1484),.clk(gclk));
	jand g0843(.dina(n1484),.dinb(w_in2117_0[1]),.dout(n1485),.clk(gclk));
	jnot g0844(.din(w_in3116_0[1]),.dout(n1486),.clk(gclk));
	jand g0845(.dina(n1486),.dinb(w_in2116_0[1]),.dout(n1487),.clk(gclk));
	jor g0846(.dina(n1487),.dinb(n1485),.dout(n1488),.clk(gclk));
	jand g0847(.dina(n1488),.dinb(n1483),.dout(n1489),.clk(gclk));
	jnot g0848(.din(w_in3119_0[1]),.dout(n1490),.clk(gclk));
	jand g0849(.dina(n1490),.dinb(w_in2119_0[1]),.dout(n1491),.clk(gclk));
	jnot g0850(.din(w_n1475_0[0]),.dout(n1492),.clk(gclk));
	jnot g0851(.din(w_in3118_0[1]),.dout(n1493),.clk(gclk));
	jand g0852(.dina(n1493),.dinb(w_in2118_0[1]),.dout(n1494),.clk(gclk));
	jand g0853(.dina(n1494),.dinb(n1492),.dout(n1495),.clk(gclk));
	jor g0854(.dina(n1495),.dinb(n1491),.dout(n1496),.clk(gclk));
	jor g0855(.dina(n1496),.dinb(n1489),.dout(n1497),.clk(gclk));
	jor g0856(.dina(w_n1497_0[1]),.dinb(n1482),.dout(n1498),.clk(gclk));
	jnot g0857(.din(w_in2123_0[2]),.dout(n1499),.clk(gclk));
	jand g0858(.dina(w_in3123_0[2]),.dinb(n1499),.dout(n1500),.clk(gclk));
	jnot g0859(.din(w_in2122_0[2]),.dout(n1501),.clk(gclk));
	jand g0860(.dina(w_in3122_0[2]),.dinb(n1501),.dout(n1502),.clk(gclk));
	jor g0861(.dina(n1502),.dinb(n1500),.dout(n1503),.clk(gclk));
	jnot g0862(.din(w_in2121_0[2]),.dout(n1504),.clk(gclk));
	jand g0863(.dina(w_in3121_0[2]),.dinb(n1504),.dout(n1505),.clk(gclk));
	jnot g0864(.din(w_in2120_0[2]),.dout(n1506),.clk(gclk));
	jand g0865(.dina(w_in3120_0[2]),.dinb(n1506),.dout(n1507),.clk(gclk));
	jor g0866(.dina(n1507),.dinb(w_n1505_0[1]),.dout(n1508),.clk(gclk));
	jor g0867(.dina(n1508),.dinb(w_n1503_0[1]),.dout(n1509),.clk(gclk));
	jnot g0868(.din(w_n1509_0[1]),.dout(n1510),.clk(gclk));
	jand g0869(.dina(n1510),.dinb(n1498),.dout(n1511),.clk(gclk));
	jnot g0870(.din(w_in3123_0[1]),.dout(n1512),.clk(gclk));
	jand g0871(.dina(n1512),.dinb(w_in2123_0[1]),.dout(n1513),.clk(gclk));
	jnot g0872(.din(w_n1503_0[0]),.dout(n1514),.clk(gclk));
	jnot g0873(.din(w_n1505_0[0]),.dout(n1515),.clk(gclk));
	jnot g0874(.din(w_in3120_0[1]),.dout(n1516),.clk(gclk));
	jand g0875(.dina(n1516),.dinb(w_in2120_0[1]),.dout(n1517),.clk(gclk));
	jand g0876(.dina(n1517),.dinb(n1515),.dout(n1518),.clk(gclk));
	jnot g0877(.din(w_in3121_0[1]),.dout(n1519),.clk(gclk));
	jand g0878(.dina(n1519),.dinb(w_in2121_0[1]),.dout(n1520),.clk(gclk));
	jnot g0879(.din(w_in3122_0[1]),.dout(n1521),.clk(gclk));
	jand g0880(.dina(n1521),.dinb(w_in2122_0[1]),.dout(n1522),.clk(gclk));
	jor g0881(.dina(n1522),.dinb(n1520),.dout(n1523),.clk(gclk));
	jor g0882(.dina(n1523),.dinb(n1518),.dout(n1524),.clk(gclk));
	jand g0883(.dina(n1524),.dinb(n1514),.dout(n1525),.clk(gclk));
	jor g0884(.dina(n1525),.dinb(n1513),.dout(n1526),.clk(gclk));
	jor g0885(.dina(w_n1526_0[1]),.dinb(n1511),.dout(n1527),.clk(gclk));
	jnot g0886(.din(w_in2126_0[2]),.dout(n1528),.clk(gclk));
	jand g0887(.dina(w_in3126_0[2]),.dinb(n1528),.dout(n1529),.clk(gclk));
	jnot g0888(.din(w_in2125_0[2]),.dout(n1530),.clk(gclk));
	jand g0889(.dina(w_in3125_0[2]),.dinb(n1530),.dout(n1531),.clk(gclk));
	jor g0890(.dina(n1531),.dinb(n1529),.dout(n1532),.clk(gclk));
	jnot g0891(.din(w_in3127_0[2]),.dout(n1533),.clk(gclk));
	jand g0892(.dina(n1533),.dinb(w_in2127_0[2]),.dout(n1534),.clk(gclk));
	jnot g0893(.din(w_in2124_0[2]),.dout(n1535),.clk(gclk));
	jand g0894(.dina(w_in3124_0[2]),.dinb(n1535),.dout(n1536),.clk(gclk));
	jor g0895(.dina(n1536),.dinb(w_n1534_0[1]),.dout(n1537),.clk(gclk));
	jor g0896(.dina(n1537),.dinb(w_n1532_0[1]),.dout(n1538),.clk(gclk));
	jnot g0897(.din(w_n1538_0[1]),.dout(n1539),.clk(gclk));
	jand g0898(.dina(n1539),.dinb(n1527),.dout(n1540),.clk(gclk));
	jnot g0899(.din(w_n1534_0[0]),.dout(n1541),.clk(gclk));
	jnot g0900(.din(w_n1532_0[0]),.dout(n1542),.clk(gclk));
	jnot g0901(.din(w_in3124_0[1]),.dout(n1543),.clk(gclk));
	jand g0902(.dina(n1543),.dinb(w_in2124_0[1]),.dout(n1544),.clk(gclk));
	jnot g0903(.din(w_in3125_0[1]),.dout(n1545),.clk(gclk));
	jand g0904(.dina(n1545),.dinb(w_in2125_0[1]),.dout(n1546),.clk(gclk));
	jor g0905(.dina(n1546),.dinb(n1544),.dout(n1547),.clk(gclk));
	jand g0906(.dina(n1547),.dinb(n1542),.dout(n1548),.clk(gclk));
	jnot g0907(.din(w_in3126_0[1]),.dout(n1549),.clk(gclk));
	jand g0908(.dina(n1549),.dinb(w_in2126_0[1]),.dout(n1550),.clk(gclk));
	jor g0909(.dina(n1550),.dinb(n1548),.dout(n1551),.clk(gclk));
	jand g0910(.dina(n1551),.dinb(n1541),.dout(n1552),.clk(gclk));
	jnot g0911(.din(w_in2127_0[1]),.dout(n1553),.clk(gclk));
	jand g0912(.dina(w_in3127_0[1]),.dinb(n1553),.dout(n1554),.clk(gclk));
	jor g0913(.dina(n1554),.dinb(n1552),.dout(n1555),.clk(gclk));
	jor g0914(.dina(w_n1555_0[1]),.dinb(n1540),.dout(n1556),.clk(gclk));
	jand g0915(.dina(w_n1556_63[2]),.dinb(w_in20_0[1]),.dout(n1557),.clk(gclk));
	jnot g0916(.din(w_n646_0[0]),.dout(n1558),.clk(gclk));
	jnot g0917(.din(w_n651_0[0]),.dout(n1559),.clk(gclk));
	jnot g0918(.din(w_n656_0[0]),.dout(n1560),.clk(gclk));
	jnot g0919(.din(w_n661_0[0]),.dout(n1561),.clk(gclk));
	jnot g0920(.din(w_n666_0[0]),.dout(n1562),.clk(gclk));
	jnot g0921(.din(w_n671_0[0]),.dout(n1563),.clk(gclk));
	jnot g0922(.din(w_n676_0[0]),.dout(n1564),.clk(gclk));
	jnot g0923(.din(w_n681_0[0]),.dout(n1565),.clk(gclk));
	jnot g0924(.din(w_n686_0[0]),.dout(n1566),.clk(gclk));
	jnot g0925(.din(w_n691_0[0]),.dout(n1567),.clk(gclk));
	jnot g0926(.din(w_n696_0[0]),.dout(n1568),.clk(gclk));
	jnot g0927(.din(w_n701_0[0]),.dout(n1569),.clk(gclk));
	jnot g0928(.din(w_n706_0[0]),.dout(n1570),.clk(gclk));
	jnot g0929(.din(w_n711_0[0]),.dout(n1571),.clk(gclk));
	jnot g0930(.din(w_n716_0[0]),.dout(n1572),.clk(gclk));
	jnot g0931(.din(w_n721_0[0]),.dout(n1573),.clk(gclk));
	jnot g0932(.din(w_n726_0[0]),.dout(n1574),.clk(gclk));
	jnot g0933(.din(w_n731_0[0]),.dout(n1575),.clk(gclk));
	jnot g0934(.din(w_n736_0[0]),.dout(n1576),.clk(gclk));
	jnot g0935(.din(w_n741_0[0]),.dout(n1577),.clk(gclk));
	jnot g0936(.din(w_n746_0[0]),.dout(n1578),.clk(gclk));
	jnot g0937(.din(w_n751_0[0]),.dout(n1579),.clk(gclk));
	jnot g0938(.din(w_n756_0[0]),.dout(n1580),.clk(gclk));
	jnot g0939(.din(w_n761_0[0]),.dout(n1581),.clk(gclk));
	jnot g0940(.din(w_n766_0[0]),.dout(n1582),.clk(gclk));
	jnot g0941(.din(w_n771_0[0]),.dout(n1583),.clk(gclk));
	jnot g0942(.din(w_n776_0[0]),.dout(n1584),.clk(gclk));
	jnot g0943(.din(w_n781_0[0]),.dout(n1585),.clk(gclk));
	jnot g0944(.din(w_in21_0[2]),.dout(n1586),.clk(gclk));
	jor g0945(.dina(w_in31_1[0]),.dinb(w_n1586_0[1]),.dout(n1587),.clk(gclk));
	jand g0946(.dina(w_in31_0[2]),.dinb(w_n1586_0[0]),.dout(n1588),.clk(gclk));
	jnot g0947(.din(w_in20_0[0]),.dout(n1589),.clk(gclk));
	jor g0948(.dina(w_in30_0[1]),.dinb(w_n1589_0[1]),.dout(n1590),.clk(gclk));
	jor g0949(.dina(n1590),.dinb(n1588),.dout(n1591),.clk(gclk));
	jand g0950(.dina(n1591),.dinb(n1587),.dout(n1592),.clk(gclk));
	jor g0951(.dina(n1592),.dinb(w_n783_0[0]),.dout(n1593),.clk(gclk));
	jand g0952(.dina(n1593),.dinb(n1585),.dout(n1594),.clk(gclk));
	jor g0953(.dina(n1594),.dinb(w_n778_0[0]),.dout(n1595),.clk(gclk));
	jand g0954(.dina(n1595),.dinb(n1584),.dout(n1596),.clk(gclk));
	jor g0955(.dina(n1596),.dinb(w_n773_0[0]),.dout(n1597),.clk(gclk));
	jand g0956(.dina(n1597),.dinb(n1583),.dout(n1598),.clk(gclk));
	jor g0957(.dina(n1598),.dinb(w_n768_0[0]),.dout(n1599),.clk(gclk));
	jand g0958(.dina(n1599),.dinb(n1582),.dout(n1600),.clk(gclk));
	jor g0959(.dina(n1600),.dinb(w_n763_0[0]),.dout(n1601),.clk(gclk));
	jand g0960(.dina(n1601),.dinb(n1581),.dout(n1602),.clk(gclk));
	jor g0961(.dina(n1602),.dinb(w_n758_0[0]),.dout(n1603),.clk(gclk));
	jand g0962(.dina(n1603),.dinb(n1580),.dout(n1604),.clk(gclk));
	jor g0963(.dina(n1604),.dinb(w_n753_0[0]),.dout(n1605),.clk(gclk));
	jand g0964(.dina(n1605),.dinb(n1579),.dout(n1606),.clk(gclk));
	jor g0965(.dina(n1606),.dinb(w_n748_0[0]),.dout(n1607),.clk(gclk));
	jand g0966(.dina(n1607),.dinb(n1578),.dout(n1608),.clk(gclk));
	jor g0967(.dina(n1608),.dinb(w_n743_0[0]),.dout(n1609),.clk(gclk));
	jand g0968(.dina(n1609),.dinb(n1577),.dout(n1610),.clk(gclk));
	jor g0969(.dina(n1610),.dinb(w_n738_0[0]),.dout(n1611),.clk(gclk));
	jand g0970(.dina(n1611),.dinb(n1576),.dout(n1612),.clk(gclk));
	jor g0971(.dina(n1612),.dinb(w_n733_0[0]),.dout(n1613),.clk(gclk));
	jand g0972(.dina(n1613),.dinb(n1575),.dout(n1614),.clk(gclk));
	jor g0973(.dina(n1614),.dinb(w_n728_0[0]),.dout(n1615),.clk(gclk));
	jand g0974(.dina(n1615),.dinb(n1574),.dout(n1616),.clk(gclk));
	jor g0975(.dina(n1616),.dinb(w_n723_0[0]),.dout(n1617),.clk(gclk));
	jand g0976(.dina(n1617),.dinb(n1573),.dout(n1618),.clk(gclk));
	jor g0977(.dina(n1618),.dinb(w_n718_0[0]),.dout(n1619),.clk(gclk));
	jand g0978(.dina(n1619),.dinb(n1572),.dout(n1620),.clk(gclk));
	jor g0979(.dina(n1620),.dinb(w_n713_0[0]),.dout(n1621),.clk(gclk));
	jand g0980(.dina(n1621),.dinb(n1571),.dout(n1622),.clk(gclk));
	jor g0981(.dina(n1622),.dinb(w_n708_0[0]),.dout(n1623),.clk(gclk));
	jand g0982(.dina(n1623),.dinb(n1570),.dout(n1624),.clk(gclk));
	jor g0983(.dina(n1624),.dinb(w_n703_0[0]),.dout(n1625),.clk(gclk));
	jand g0984(.dina(n1625),.dinb(n1569),.dout(n1626),.clk(gclk));
	jor g0985(.dina(n1626),.dinb(w_n698_0[0]),.dout(n1627),.clk(gclk));
	jand g0986(.dina(n1627),.dinb(n1568),.dout(n1628),.clk(gclk));
	jor g0987(.dina(n1628),.dinb(w_n693_0[0]),.dout(n1629),.clk(gclk));
	jand g0988(.dina(n1629),.dinb(n1567),.dout(n1630),.clk(gclk));
	jor g0989(.dina(n1630),.dinb(w_n688_0[0]),.dout(n1631),.clk(gclk));
	jand g0990(.dina(n1631),.dinb(n1566),.dout(n1632),.clk(gclk));
	jor g0991(.dina(n1632),.dinb(w_n683_0[0]),.dout(n1633),.clk(gclk));
	jand g0992(.dina(n1633),.dinb(n1565),.dout(n1634),.clk(gclk));
	jor g0993(.dina(n1634),.dinb(w_n678_0[0]),.dout(n1635),.clk(gclk));
	jand g0994(.dina(n1635),.dinb(n1564),.dout(n1636),.clk(gclk));
	jor g0995(.dina(n1636),.dinb(w_n673_0[0]),.dout(n1637),.clk(gclk));
	jand g0996(.dina(n1637),.dinb(n1563),.dout(n1638),.clk(gclk));
	jor g0997(.dina(n1638),.dinb(w_n668_0[0]),.dout(n1639),.clk(gclk));
	jand g0998(.dina(n1639),.dinb(n1562),.dout(n1640),.clk(gclk));
	jor g0999(.dina(n1640),.dinb(w_n663_0[0]),.dout(n1641),.clk(gclk));
	jand g1000(.dina(n1641),.dinb(n1561),.dout(n1642),.clk(gclk));
	jor g1001(.dina(n1642),.dinb(w_n658_0[0]),.dout(n1643),.clk(gclk));
	jand g1002(.dina(n1643),.dinb(n1560),.dout(n1644),.clk(gclk));
	jor g1003(.dina(n1644),.dinb(w_n653_0[0]),.dout(n1645),.clk(gclk));
	jand g1004(.dina(n1645),.dinb(n1559),.dout(n1646),.clk(gclk));
	jor g1005(.dina(n1646),.dinb(w_n648_0[0]),.dout(n1647),.clk(gclk));
	jand g1006(.dina(n1647),.dinb(n1558),.dout(n1648),.clk(gclk));
	jor g1007(.dina(n1648),.dinb(w_n643_0[0]),.dout(n1649),.clk(gclk));
	jnot g1008(.din(w_n853_0[0]),.dout(n1650),.clk(gclk));
	jand g1009(.dina(n1650),.dinb(n1649),.dout(n1651),.clk(gclk));
	jor g1010(.dina(w_n880_0[0]),.dinb(n1651),.dout(n1652),.clk(gclk));
	jnot g1011(.din(w_n915_0[0]),.dout(n1653),.clk(gclk));
	jand g1012(.dina(n1653),.dinb(n1652),.dout(n1654),.clk(gclk));
	jor g1013(.dina(w_n939_0[0]),.dinb(n1654),.dout(n1655),.clk(gclk));
	jnot g1014(.din(w_n974_0[0]),.dout(n1656),.clk(gclk));
	jand g1015(.dina(n1656),.dinb(n1655),.dout(n1657),.clk(gclk));
	jor g1016(.dina(w_n1001_0[0]),.dinb(n1657),.dout(n1658),.clk(gclk));
	jnot g1017(.din(w_n1032_0[0]),.dout(n1659),.clk(gclk));
	jand g1018(.dina(n1659),.dinb(n1658),.dout(n1660),.clk(gclk));
	jor g1019(.dina(w_n1056_0[0]),.dinb(n1660),.dout(n1661),.clk(gclk));
	jnot g1020(.din(w_n1091_0[0]),.dout(n1662),.clk(gclk));
	jand g1021(.dina(n1662),.dinb(n1661),.dout(n1663),.clk(gclk));
	jor g1022(.dina(w_n1103_0[0]),.dinb(n1663),.dout(n1664),.clk(gclk));
	jnot g1023(.din(w_n1120_0[0]),.dout(n1665),.clk(gclk));
	jand g1024(.dina(n1665),.dinb(n1664),.dout(n1666),.clk(gclk));
	jor g1025(.dina(w_n1132_0[0]),.dinb(n1666),.dout(n1667),.clk(gclk));
	jnot g1026(.din(w_n1149_0[0]),.dout(n1668),.clk(gclk));
	jand g1027(.dina(n1668),.dinb(n1667),.dout(n1669),.clk(gclk));
	jor g1028(.dina(w_n1161_0[0]),.dinb(n1669),.dout(n1670),.clk(gclk));
	jnot g1029(.din(w_n1178_0[0]),.dout(n1671),.clk(gclk));
	jand g1030(.dina(n1671),.dinb(n1670),.dout(n1672),.clk(gclk));
	jor g1031(.dina(w_n1190_0[0]),.dinb(n1672),.dout(n1673),.clk(gclk));
	jnot g1032(.din(w_n1207_0[0]),.dout(n1674),.clk(gclk));
	jand g1033(.dina(n1674),.dinb(n1673),.dout(n1675),.clk(gclk));
	jor g1034(.dina(w_n1219_0[0]),.dinb(n1675),.dout(n1676),.clk(gclk));
	jnot g1035(.din(w_n1236_0[0]),.dout(n1677),.clk(gclk));
	jand g1036(.dina(n1677),.dinb(n1676),.dout(n1678),.clk(gclk));
	jor g1037(.dina(w_n1248_0[0]),.dinb(n1678),.dout(n1679),.clk(gclk));
	jnot g1038(.din(w_n1265_0[0]),.dout(n1680),.clk(gclk));
	jand g1039(.dina(n1680),.dinb(n1679),.dout(n1681),.clk(gclk));
	jor g1040(.dina(w_n1277_0[0]),.dinb(n1681),.dout(n1682),.clk(gclk));
	jnot g1041(.din(w_n1294_0[0]),.dout(n1683),.clk(gclk));
	jand g1042(.dina(n1683),.dinb(n1682),.dout(n1684),.clk(gclk));
	jor g1043(.dina(w_n1306_0[0]),.dinb(n1684),.dout(n1685),.clk(gclk));
	jnot g1044(.din(w_n1323_0[0]),.dout(n1686),.clk(gclk));
	jand g1045(.dina(n1686),.dinb(n1685),.dout(n1687),.clk(gclk));
	jor g1046(.dina(w_n1335_0[0]),.dinb(n1687),.dout(n1688),.clk(gclk));
	jnot g1047(.din(w_n1352_0[0]),.dout(n1689),.clk(gclk));
	jand g1048(.dina(n1689),.dinb(n1688),.dout(n1690),.clk(gclk));
	jor g1049(.dina(w_n1364_0[0]),.dinb(n1690),.dout(n1691),.clk(gclk));
	jnot g1050(.din(w_n1381_0[0]),.dout(n1692),.clk(gclk));
	jand g1051(.dina(n1692),.dinb(n1691),.dout(n1693),.clk(gclk));
	jor g1052(.dina(w_n1393_0[0]),.dinb(n1693),.dout(n1694),.clk(gclk));
	jnot g1053(.din(w_n1410_0[0]),.dout(n1695),.clk(gclk));
	jand g1054(.dina(n1695),.dinb(n1694),.dout(n1696),.clk(gclk));
	jor g1055(.dina(w_n1422_0[0]),.dinb(n1696),.dout(n1697),.clk(gclk));
	jnot g1056(.din(w_n1439_0[0]),.dout(n1698),.clk(gclk));
	jand g1057(.dina(n1698),.dinb(n1697),.dout(n1699),.clk(gclk));
	jor g1058(.dina(w_n1451_0[0]),.dinb(n1699),.dout(n1700),.clk(gclk));
	jnot g1059(.din(w_n1468_0[0]),.dout(n1701),.clk(gclk));
	jand g1060(.dina(n1701),.dinb(n1700),.dout(n1702),.clk(gclk));
	jor g1061(.dina(w_n1480_0[0]),.dinb(n1702),.dout(n1703),.clk(gclk));
	jnot g1062(.din(w_n1497_0[0]),.dout(n1704),.clk(gclk));
	jand g1063(.dina(n1704),.dinb(n1703),.dout(n1705),.clk(gclk));
	jor g1064(.dina(w_n1509_0[0]),.dinb(n1705),.dout(n1706),.clk(gclk));
	jnot g1065(.din(w_n1526_0[0]),.dout(n1707),.clk(gclk));
	jand g1066(.dina(n1707),.dinb(n1706),.dout(n1708),.clk(gclk));
	jor g1067(.dina(w_n1538_0[0]),.dinb(n1708),.dout(n1709),.clk(gclk));
	jnot g1068(.din(w_n1555_0[0]),.dout(n1710),.clk(gclk));
	jand g1069(.dina(n1710),.dinb(n1709),.dout(n1711),.clk(gclk));
	jand g1070(.dina(w_n1711_64[1]),.dinb(w_in30_0[0]),.dout(n1712),.clk(gclk));
	jor g1071(.dina(n1712),.dinb(n1557),.dout(n1713),.clk(gclk));
	jnot g1072(.din(w_in030_0[2]),.dout(n1714),.clk(gclk));
	jand g1073(.dina(w_in130_0[2]),.dinb(n1714),.dout(n1715),.clk(gclk));
	jnot g1074(.din(w_n1715_0[1]),.dout(n1716),.clk(gclk));
	jnot g1075(.din(w_in129_0[2]),.dout(n1717),.clk(gclk));
	jand g1076(.dina(n1717),.dinb(w_in029_0[2]),.dout(n1718),.clk(gclk));
	jnot g1077(.din(w_in029_0[1]),.dout(n1719),.clk(gclk));
	jand g1078(.dina(w_in129_0[1]),.dinb(n1719),.dout(n1720),.clk(gclk));
	jnot g1079(.din(w_n1720_0[1]),.dout(n1721),.clk(gclk));
	jnot g1080(.din(w_in128_0[2]),.dout(n1722),.clk(gclk));
	jand g1081(.dina(n1722),.dinb(w_in028_0[2]),.dout(n1723),.clk(gclk));
	jnot g1082(.din(w_in028_0[1]),.dout(n1724),.clk(gclk));
	jand g1083(.dina(w_in128_0[1]),.dinb(n1724),.dout(n1725),.clk(gclk));
	jnot g1084(.din(w_n1725_0[1]),.dout(n1726),.clk(gclk));
	jnot g1085(.din(w_in127_0[2]),.dout(n1727),.clk(gclk));
	jand g1086(.dina(n1727),.dinb(w_in027_0[2]),.dout(n1728),.clk(gclk));
	jnot g1087(.din(w_in027_0[1]),.dout(n1729),.clk(gclk));
	jand g1088(.dina(w_in127_0[1]),.dinb(n1729),.dout(n1730),.clk(gclk));
	jnot g1089(.din(w_n1730_0[1]),.dout(n1731),.clk(gclk));
	jnot g1090(.din(w_in126_0[2]),.dout(n1732),.clk(gclk));
	jand g1091(.dina(n1732),.dinb(w_in026_0[2]),.dout(n1733),.clk(gclk));
	jnot g1092(.din(w_in026_0[1]),.dout(n1734),.clk(gclk));
	jand g1093(.dina(w_in126_0[1]),.dinb(n1734),.dout(n1735),.clk(gclk));
	jnot g1094(.din(w_n1735_0[1]),.dout(n1736),.clk(gclk));
	jnot g1095(.din(w_in125_0[2]),.dout(n1737),.clk(gclk));
	jand g1096(.dina(n1737),.dinb(w_in025_0[2]),.dout(n1738),.clk(gclk));
	jnot g1097(.din(w_in025_0[1]),.dout(n1739),.clk(gclk));
	jand g1098(.dina(w_in125_0[1]),.dinb(n1739),.dout(n1740),.clk(gclk));
	jnot g1099(.din(w_n1740_0[1]),.dout(n1741),.clk(gclk));
	jnot g1100(.din(w_in124_0[2]),.dout(n1742),.clk(gclk));
	jand g1101(.dina(n1742),.dinb(w_in024_0[2]),.dout(n1743),.clk(gclk));
	jnot g1102(.din(w_in024_0[1]),.dout(n1744),.clk(gclk));
	jand g1103(.dina(w_in124_0[1]),.dinb(n1744),.dout(n1745),.clk(gclk));
	jnot g1104(.din(w_n1745_0[1]),.dout(n1746),.clk(gclk));
	jnot g1105(.din(w_in123_0[2]),.dout(n1747),.clk(gclk));
	jand g1106(.dina(n1747),.dinb(w_in023_0[2]),.dout(n1748),.clk(gclk));
	jnot g1107(.din(w_in023_0[1]),.dout(n1749),.clk(gclk));
	jand g1108(.dina(w_in123_0[1]),.dinb(n1749),.dout(n1750),.clk(gclk));
	jnot g1109(.din(w_n1750_0[1]),.dout(n1751),.clk(gclk));
	jnot g1110(.din(w_in122_0[2]),.dout(n1752),.clk(gclk));
	jand g1111(.dina(n1752),.dinb(w_in022_0[2]),.dout(n1753),.clk(gclk));
	jnot g1112(.din(w_in022_0[1]),.dout(n1754),.clk(gclk));
	jand g1113(.dina(w_in122_0[1]),.dinb(n1754),.dout(n1755),.clk(gclk));
	jnot g1114(.din(w_n1755_0[1]),.dout(n1756),.clk(gclk));
	jnot g1115(.din(w_in121_0[2]),.dout(n1757),.clk(gclk));
	jand g1116(.dina(n1757),.dinb(w_in021_0[2]),.dout(n1758),.clk(gclk));
	jnot g1117(.din(w_in021_0[1]),.dout(n1759),.clk(gclk));
	jand g1118(.dina(w_in121_0[1]),.dinb(n1759),.dout(n1760),.clk(gclk));
	jnot g1119(.din(w_n1760_0[1]),.dout(n1761),.clk(gclk));
	jnot g1120(.din(w_in120_0[2]),.dout(n1762),.clk(gclk));
	jand g1121(.dina(n1762),.dinb(w_in020_0[2]),.dout(n1763),.clk(gclk));
	jnot g1122(.din(w_in020_0[1]),.dout(n1764),.clk(gclk));
	jand g1123(.dina(w_in120_0[1]),.dinb(n1764),.dout(n1765),.clk(gclk));
	jnot g1124(.din(w_n1765_0[1]),.dout(n1766),.clk(gclk));
	jnot g1125(.din(w_in119_0[2]),.dout(n1767),.clk(gclk));
	jand g1126(.dina(n1767),.dinb(w_in019_0[2]),.dout(n1768),.clk(gclk));
	jnot g1127(.din(w_in019_0[1]),.dout(n1769),.clk(gclk));
	jand g1128(.dina(w_in119_0[1]),.dinb(n1769),.dout(n1770),.clk(gclk));
	jnot g1129(.din(w_n1770_0[1]),.dout(n1771),.clk(gclk));
	jnot g1130(.din(w_in118_0[2]),.dout(n1772),.clk(gclk));
	jand g1131(.dina(n1772),.dinb(w_in018_0[2]),.dout(n1773),.clk(gclk));
	jnot g1132(.din(w_in018_0[1]),.dout(n1774),.clk(gclk));
	jand g1133(.dina(w_in118_0[1]),.dinb(n1774),.dout(n1775),.clk(gclk));
	jnot g1134(.din(w_n1775_0[1]),.dout(n1776),.clk(gclk));
	jnot g1135(.din(w_in117_0[2]),.dout(n1777),.clk(gclk));
	jand g1136(.dina(n1777),.dinb(w_in017_0[2]),.dout(n1778),.clk(gclk));
	jnot g1137(.din(w_in017_0[1]),.dout(n1779),.clk(gclk));
	jand g1138(.dina(w_in117_0[1]),.dinb(n1779),.dout(n1780),.clk(gclk));
	jnot g1139(.din(w_n1780_0[1]),.dout(n1781),.clk(gclk));
	jnot g1140(.din(w_in116_0[2]),.dout(n1782),.clk(gclk));
	jand g1141(.dina(n1782),.dinb(w_in016_0[2]),.dout(n1783),.clk(gclk));
	jnot g1142(.din(w_in016_0[1]),.dout(n1784),.clk(gclk));
	jand g1143(.dina(w_in116_0[1]),.dinb(n1784),.dout(n1785),.clk(gclk));
	jnot g1144(.din(w_n1785_0[1]),.dout(n1786),.clk(gclk));
	jnot g1145(.din(w_in115_0[2]),.dout(n1787),.clk(gclk));
	jand g1146(.dina(n1787),.dinb(w_in015_0[2]),.dout(n1788),.clk(gclk));
	jnot g1147(.din(w_in015_0[1]),.dout(n1789),.clk(gclk));
	jand g1148(.dina(w_in115_0[1]),.dinb(n1789),.dout(n1790),.clk(gclk));
	jnot g1149(.din(w_n1790_0[1]),.dout(n1791),.clk(gclk));
	jnot g1150(.din(w_in114_0[2]),.dout(n1792),.clk(gclk));
	jand g1151(.dina(n1792),.dinb(w_in014_0[2]),.dout(n1793),.clk(gclk));
	jnot g1152(.din(w_in014_0[1]),.dout(n1794),.clk(gclk));
	jand g1153(.dina(w_in114_0[1]),.dinb(n1794),.dout(n1795),.clk(gclk));
	jnot g1154(.din(w_n1795_0[1]),.dout(n1796),.clk(gclk));
	jnot g1155(.din(w_in113_0[2]),.dout(n1797),.clk(gclk));
	jand g1156(.dina(n1797),.dinb(w_in013_0[2]),.dout(n1798),.clk(gclk));
	jnot g1157(.din(w_in013_0[1]),.dout(n1799),.clk(gclk));
	jand g1158(.dina(w_in113_0[1]),.dinb(n1799),.dout(n1800),.clk(gclk));
	jnot g1159(.din(w_n1800_0[1]),.dout(n1801),.clk(gclk));
	jnot g1160(.din(w_in112_0[2]),.dout(n1802),.clk(gclk));
	jand g1161(.dina(n1802),.dinb(w_in012_0[2]),.dout(n1803),.clk(gclk));
	jnot g1162(.din(w_in012_0[1]),.dout(n1804),.clk(gclk));
	jand g1163(.dina(w_in112_0[1]),.dinb(n1804),.dout(n1805),.clk(gclk));
	jnot g1164(.din(w_n1805_0[1]),.dout(n1806),.clk(gclk));
	jnot g1165(.din(w_in111_0[2]),.dout(n1807),.clk(gclk));
	jand g1166(.dina(n1807),.dinb(w_in011_0[2]),.dout(n1808),.clk(gclk));
	jnot g1167(.din(w_in011_0[1]),.dout(n1809),.clk(gclk));
	jand g1168(.dina(w_in111_0[1]),.dinb(n1809),.dout(n1810),.clk(gclk));
	jnot g1169(.din(w_n1810_0[1]),.dout(n1811),.clk(gclk));
	jnot g1170(.din(w_in110_0[2]),.dout(n1812),.clk(gclk));
	jand g1171(.dina(n1812),.dinb(w_in010_0[2]),.dout(n1813),.clk(gclk));
	jnot g1172(.din(w_in010_0[1]),.dout(n1814),.clk(gclk));
	jand g1173(.dina(w_in110_0[1]),.dinb(n1814),.dout(n1815),.clk(gclk));
	jnot g1174(.din(w_n1815_0[1]),.dout(n1816),.clk(gclk));
	jnot g1175(.din(w_in19_0[2]),.dout(n1817),.clk(gclk));
	jand g1176(.dina(n1817),.dinb(w_in09_0[2]),.dout(n1818),.clk(gclk));
	jnot g1177(.din(w_in09_0[1]),.dout(n1819),.clk(gclk));
	jand g1178(.dina(w_in19_0[1]),.dinb(n1819),.dout(n1820),.clk(gclk));
	jnot g1179(.din(w_n1820_0[1]),.dout(n1821),.clk(gclk));
	jnot g1180(.din(w_in18_0[2]),.dout(n1822),.clk(gclk));
	jand g1181(.dina(n1822),.dinb(w_in08_0[2]),.dout(n1823),.clk(gclk));
	jnot g1182(.din(w_in08_0[1]),.dout(n1824),.clk(gclk));
	jand g1183(.dina(w_in18_0[1]),.dinb(n1824),.dout(n1825),.clk(gclk));
	jnot g1184(.din(w_n1825_0[1]),.dout(n1826),.clk(gclk));
	jnot g1185(.din(w_in17_0[2]),.dout(n1827),.clk(gclk));
	jand g1186(.dina(n1827),.dinb(w_in07_0[2]),.dout(n1828),.clk(gclk));
	jnot g1187(.din(w_in07_0[1]),.dout(n1829),.clk(gclk));
	jand g1188(.dina(w_in17_0[1]),.dinb(n1829),.dout(n1830),.clk(gclk));
	jnot g1189(.din(w_n1830_0[1]),.dout(n1831),.clk(gclk));
	jnot g1190(.din(w_in16_0[2]),.dout(n1832),.clk(gclk));
	jand g1191(.dina(n1832),.dinb(w_in06_0[2]),.dout(n1833),.clk(gclk));
	jnot g1192(.din(w_in06_0[1]),.dout(n1834),.clk(gclk));
	jand g1193(.dina(w_in16_0[1]),.dinb(n1834),.dout(n1835),.clk(gclk));
	jnot g1194(.din(w_n1835_0[1]),.dout(n1836),.clk(gclk));
	jnot g1195(.din(w_in15_0[2]),.dout(n1837),.clk(gclk));
	jand g1196(.dina(n1837),.dinb(w_in05_0[2]),.dout(n1838),.clk(gclk));
	jnot g1197(.din(w_in05_0[1]),.dout(n1839),.clk(gclk));
	jand g1198(.dina(w_in15_0[1]),.dinb(n1839),.dout(n1840),.clk(gclk));
	jnot g1199(.din(w_n1840_0[1]),.dout(n1841),.clk(gclk));
	jnot g1200(.din(w_in14_0[2]),.dout(n1842),.clk(gclk));
	jand g1201(.dina(n1842),.dinb(w_in04_0[2]),.dout(n1843),.clk(gclk));
	jnot g1202(.din(w_in04_0[1]),.dout(n1844),.clk(gclk));
	jand g1203(.dina(w_in14_0[1]),.dinb(n1844),.dout(n1845),.clk(gclk));
	jnot g1204(.din(w_n1845_0[1]),.dout(n1846),.clk(gclk));
	jnot g1205(.din(w_in13_0[2]),.dout(n1847),.clk(gclk));
	jand g1206(.dina(n1847),.dinb(w_in03_0[2]),.dout(n1848),.clk(gclk));
	jnot g1207(.din(w_in03_0[1]),.dout(n1849),.clk(gclk));
	jand g1208(.dina(w_in13_0[1]),.dinb(n1849),.dout(n1850),.clk(gclk));
	jnot g1209(.din(w_n1850_0[1]),.dout(n1851),.clk(gclk));
	jnot g1210(.din(w_in12_0[2]),.dout(n1852),.clk(gclk));
	jand g1211(.dina(w_n1852_0[1]),.dinb(w_in02_0[2]),.dout(n1853),.clk(gclk));
	jnot g1212(.din(w_in02_0[1]),.dout(n1854),.clk(gclk));
	jand g1213(.dina(w_in12_0[1]),.dinb(w_n1854_0[1]),.dout(n1855),.clk(gclk));
	jnot g1214(.din(w_n1855_0[1]),.dout(n1856),.clk(gclk));
	jnot g1215(.din(w_in11_1[1]),.dout(n1857),.clk(gclk));
	jand g1216(.dina(w_n1857_0[2]),.dinb(w_in01_1[1]),.dout(n1858),.clk(gclk));
	jor g1217(.dina(w_n1857_0[1]),.dinb(w_in01_1[0]),.dout(n1859),.clk(gclk));
	jnot g1218(.din(w_in10_0[2]),.dout(n1860),.clk(gclk));
	jand g1219(.dina(w_n1860_0[1]),.dinb(w_in00_0[2]),.dout(n1861),.clk(gclk));
	jand g1220(.dina(n1861),.dinb(n1859),.dout(n1862),.clk(gclk));
	jor g1221(.dina(n1862),.dinb(n1858),.dout(n1863),.clk(gclk));
	jand g1222(.dina(n1863),.dinb(n1856),.dout(n1864),.clk(gclk));
	jor g1223(.dina(n1864),.dinb(w_n1853_0[1]),.dout(n1865),.clk(gclk));
	jand g1224(.dina(n1865),.dinb(n1851),.dout(n1866),.clk(gclk));
	jor g1225(.dina(n1866),.dinb(w_n1848_0[1]),.dout(n1867),.clk(gclk));
	jand g1226(.dina(n1867),.dinb(n1846),.dout(n1868),.clk(gclk));
	jor g1227(.dina(n1868),.dinb(w_n1843_0[1]),.dout(n1869),.clk(gclk));
	jand g1228(.dina(n1869),.dinb(n1841),.dout(n1870),.clk(gclk));
	jor g1229(.dina(n1870),.dinb(w_n1838_0[1]),.dout(n1871),.clk(gclk));
	jand g1230(.dina(n1871),.dinb(n1836),.dout(n1872),.clk(gclk));
	jor g1231(.dina(n1872),.dinb(w_n1833_0[1]),.dout(n1873),.clk(gclk));
	jand g1232(.dina(n1873),.dinb(n1831),.dout(n1874),.clk(gclk));
	jor g1233(.dina(n1874),.dinb(w_n1828_0[1]),.dout(n1875),.clk(gclk));
	jand g1234(.dina(n1875),.dinb(n1826),.dout(n1876),.clk(gclk));
	jor g1235(.dina(n1876),.dinb(w_n1823_0[1]),.dout(n1877),.clk(gclk));
	jand g1236(.dina(n1877),.dinb(n1821),.dout(n1878),.clk(gclk));
	jor g1237(.dina(n1878),.dinb(w_n1818_0[1]),.dout(n1879),.clk(gclk));
	jand g1238(.dina(n1879),.dinb(n1816),.dout(n1880),.clk(gclk));
	jor g1239(.dina(n1880),.dinb(w_n1813_0[1]),.dout(n1881),.clk(gclk));
	jand g1240(.dina(n1881),.dinb(n1811),.dout(n1882),.clk(gclk));
	jor g1241(.dina(n1882),.dinb(w_n1808_0[1]),.dout(n1883),.clk(gclk));
	jand g1242(.dina(n1883),.dinb(n1806),.dout(n1884),.clk(gclk));
	jor g1243(.dina(n1884),.dinb(w_n1803_0[1]),.dout(n1885),.clk(gclk));
	jand g1244(.dina(n1885),.dinb(n1801),.dout(n1886),.clk(gclk));
	jor g1245(.dina(n1886),.dinb(w_n1798_0[1]),.dout(n1887),.clk(gclk));
	jand g1246(.dina(n1887),.dinb(n1796),.dout(n1888),.clk(gclk));
	jor g1247(.dina(n1888),.dinb(w_n1793_0[1]),.dout(n1889),.clk(gclk));
	jand g1248(.dina(n1889),.dinb(n1791),.dout(n1890),.clk(gclk));
	jor g1249(.dina(n1890),.dinb(w_n1788_0[1]),.dout(n1891),.clk(gclk));
	jand g1250(.dina(n1891),.dinb(n1786),.dout(n1892),.clk(gclk));
	jor g1251(.dina(n1892),.dinb(w_n1783_0[1]),.dout(n1893),.clk(gclk));
	jand g1252(.dina(n1893),.dinb(n1781),.dout(n1894),.clk(gclk));
	jor g1253(.dina(n1894),.dinb(w_n1778_0[1]),.dout(n1895),.clk(gclk));
	jand g1254(.dina(n1895),.dinb(n1776),.dout(n1896),.clk(gclk));
	jor g1255(.dina(n1896),.dinb(w_n1773_0[1]),.dout(n1897),.clk(gclk));
	jand g1256(.dina(n1897),.dinb(n1771),.dout(n1898),.clk(gclk));
	jor g1257(.dina(n1898),.dinb(w_n1768_0[1]),.dout(n1899),.clk(gclk));
	jand g1258(.dina(n1899),.dinb(n1766),.dout(n1900),.clk(gclk));
	jor g1259(.dina(n1900),.dinb(w_n1763_0[1]),.dout(n1901),.clk(gclk));
	jand g1260(.dina(n1901),.dinb(n1761),.dout(n1902),.clk(gclk));
	jor g1261(.dina(n1902),.dinb(w_n1758_0[1]),.dout(n1903),.clk(gclk));
	jand g1262(.dina(n1903),.dinb(n1756),.dout(n1904),.clk(gclk));
	jor g1263(.dina(n1904),.dinb(w_n1753_0[1]),.dout(n1905),.clk(gclk));
	jand g1264(.dina(n1905),.dinb(n1751),.dout(n1906),.clk(gclk));
	jor g1265(.dina(n1906),.dinb(w_n1748_0[1]),.dout(n1907),.clk(gclk));
	jand g1266(.dina(n1907),.dinb(n1746),.dout(n1908),.clk(gclk));
	jor g1267(.dina(n1908),.dinb(w_n1743_0[1]),.dout(n1909),.clk(gclk));
	jand g1268(.dina(n1909),.dinb(n1741),.dout(n1910),.clk(gclk));
	jor g1269(.dina(n1910),.dinb(w_n1738_0[1]),.dout(n1911),.clk(gclk));
	jand g1270(.dina(n1911),.dinb(n1736),.dout(n1912),.clk(gclk));
	jor g1271(.dina(n1912),.dinb(w_n1733_0[1]),.dout(n1913),.clk(gclk));
	jand g1272(.dina(n1913),.dinb(n1731),.dout(n1914),.clk(gclk));
	jor g1273(.dina(n1914),.dinb(w_n1728_0[1]),.dout(n1915),.clk(gclk));
	jand g1274(.dina(n1915),.dinb(n1726),.dout(n1916),.clk(gclk));
	jor g1275(.dina(n1916),.dinb(w_n1723_0[1]),.dout(n1917),.clk(gclk));
	jand g1276(.dina(n1917),.dinb(n1721),.dout(n1918),.clk(gclk));
	jor g1277(.dina(n1918),.dinb(w_n1718_0[1]),.dout(n1919),.clk(gclk));
	jand g1278(.dina(n1919),.dinb(n1716),.dout(n1920),.clk(gclk));
	jnot g1279(.din(w_in130_0[1]),.dout(n1921),.clk(gclk));
	jand g1280(.dina(n1921),.dinb(w_in030_0[1]),.dout(n1922),.clk(gclk));
	jnot g1281(.din(w_in131_0[2]),.dout(n1923),.clk(gclk));
	jand g1282(.dina(n1923),.dinb(w_in031_0[2]),.dout(n1924),.clk(gclk));
	jor g1283(.dina(n1924),.dinb(n1922),.dout(n1925),.clk(gclk));
	jor g1284(.dina(w_n1925_0[1]),.dinb(n1920),.dout(n1926),.clk(gclk));
	jnot g1285(.din(w_in037_0[2]),.dout(n1927),.clk(gclk));
	jand g1286(.dina(w_in137_0[2]),.dinb(n1927),.dout(n1928),.clk(gclk));
	jnot g1287(.din(w_in039_0[2]),.dout(n1929),.clk(gclk));
	jand g1288(.dina(w_in139_0[2]),.dinb(n1929),.dout(n1930),.clk(gclk));
	jnot g1289(.din(w_in038_0[2]),.dout(n1931),.clk(gclk));
	jand g1290(.dina(w_in138_0[2]),.dinb(n1931),.dout(n1932),.clk(gclk));
	jor g1291(.dina(n1932),.dinb(w_n1930_0[1]),.dout(n1933),.clk(gclk));
	jor g1292(.dina(n1933),.dinb(n1928),.dout(n1934),.clk(gclk));
	jnot g1293(.din(w_in035_0[2]),.dout(n1935),.clk(gclk));
	jand g1294(.dina(w_in135_0[2]),.dinb(n1935),.dout(n1936),.clk(gclk));
	jnot g1295(.din(w_in034_0[2]),.dout(n1937),.clk(gclk));
	jand g1296(.dina(w_in134_0[2]),.dinb(n1937),.dout(n1938),.clk(gclk));
	jor g1297(.dina(n1938),.dinb(n1936),.dout(n1939),.clk(gclk));
	jnot g1298(.din(w_in032_0[2]),.dout(n1940),.clk(gclk));
	jand g1299(.dina(w_in132_0[2]),.dinb(n1940),.dout(n1941),.clk(gclk));
	jnot g1300(.din(w_in033_0[2]),.dout(n1942),.clk(gclk));
	jand g1301(.dina(w_in133_0[2]),.dinb(n1942),.dout(n1943),.clk(gclk));
	jor g1302(.dina(w_n1943_0[1]),.dinb(n1941),.dout(n1944),.clk(gclk));
	jnot g1303(.din(w_in036_0[2]),.dout(n1945),.clk(gclk));
	jand g1304(.dina(w_in136_0[2]),.dinb(n1945),.dout(n1946),.clk(gclk));
	jnot g1305(.din(w_in031_0[1]),.dout(n1947),.clk(gclk));
	jand g1306(.dina(w_in131_0[1]),.dinb(n1947),.dout(n1948),.clk(gclk));
	jor g1307(.dina(n1948),.dinb(w_n1946_0[1]),.dout(n1949),.clk(gclk));
	jor g1308(.dina(n1949),.dinb(n1944),.dout(n1950),.clk(gclk));
	jor g1309(.dina(n1950),.dinb(w_n1939_0[1]),.dout(n1951),.clk(gclk));
	jor g1310(.dina(n1951),.dinb(w_n1934_0[1]),.dout(n1952),.clk(gclk));
	jnot g1311(.din(w_n1952_0[1]),.dout(n1953),.clk(gclk));
	jand g1312(.dina(n1953),.dinb(n1926),.dout(n1954),.clk(gclk));
	jnot g1313(.din(w_n1934_0[0]),.dout(n1955),.clk(gclk));
	jnot g1314(.din(w_n1946_0[0]),.dout(n1956),.clk(gclk));
	jnot g1315(.din(w_in135_0[1]),.dout(n1957),.clk(gclk));
	jand g1316(.dina(n1957),.dinb(w_in035_0[1]),.dout(n1958),.clk(gclk));
	jnot g1317(.din(w_n1939_0[0]),.dout(n1959),.clk(gclk));
	jnot g1318(.din(w_n1943_0[0]),.dout(n1960),.clk(gclk));
	jnot g1319(.din(w_in132_0[1]),.dout(n1961),.clk(gclk));
	jand g1320(.dina(n1961),.dinb(w_in032_0[1]),.dout(n1962),.clk(gclk));
	jand g1321(.dina(n1962),.dinb(n1960),.dout(n1963),.clk(gclk));
	jnot g1322(.din(w_in133_0[1]),.dout(n1964),.clk(gclk));
	jand g1323(.dina(n1964),.dinb(w_in033_0[1]),.dout(n1965),.clk(gclk));
	jnot g1324(.din(w_in134_0[1]),.dout(n1966),.clk(gclk));
	jand g1325(.dina(n1966),.dinb(w_in034_0[1]),.dout(n1967),.clk(gclk));
	jor g1326(.dina(n1967),.dinb(n1965),.dout(n1968),.clk(gclk));
	jor g1327(.dina(n1968),.dinb(n1963),.dout(n1969),.clk(gclk));
	jand g1328(.dina(n1969),.dinb(n1959),.dout(n1970),.clk(gclk));
	jor g1329(.dina(n1970),.dinb(n1958),.dout(n1971),.clk(gclk));
	jand g1330(.dina(n1971),.dinb(n1956),.dout(n1972),.clk(gclk));
	jnot g1331(.din(w_in136_0[1]),.dout(n1973),.clk(gclk));
	jand g1332(.dina(n1973),.dinb(w_in036_0[1]),.dout(n1974),.clk(gclk));
	jnot g1333(.din(w_in137_0[1]),.dout(n1975),.clk(gclk));
	jand g1334(.dina(n1975),.dinb(w_in037_0[1]),.dout(n1976),.clk(gclk));
	jor g1335(.dina(n1976),.dinb(n1974),.dout(n1977),.clk(gclk));
	jor g1336(.dina(n1977),.dinb(n1972),.dout(n1978),.clk(gclk));
	jand g1337(.dina(n1978),.dinb(n1955),.dout(n1979),.clk(gclk));
	jnot g1338(.din(w_n1930_0[0]),.dout(n1980),.clk(gclk));
	jnot g1339(.din(w_in138_0[1]),.dout(n1981),.clk(gclk));
	jand g1340(.dina(n1981),.dinb(w_in038_0[1]),.dout(n1982),.clk(gclk));
	jand g1341(.dina(n1982),.dinb(n1980),.dout(n1983),.clk(gclk));
	jnot g1342(.din(w_in139_0[1]),.dout(n1984),.clk(gclk));
	jand g1343(.dina(n1984),.dinb(w_in039_0[1]),.dout(n1985),.clk(gclk));
	jor g1344(.dina(n1985),.dinb(n1983),.dout(n1986),.clk(gclk));
	jor g1345(.dina(n1986),.dinb(n1979),.dout(n1987),.clk(gclk));
	jor g1346(.dina(w_n1987_0[1]),.dinb(n1954),.dout(n1988),.clk(gclk));
	jnot g1347(.din(w_in045_0[2]),.dout(n1989),.clk(gclk));
	jand g1348(.dina(w_in145_0[2]),.dinb(n1989),.dout(n1990),.clk(gclk));
	jnot g1349(.din(w_in047_0[2]),.dout(n1991),.clk(gclk));
	jand g1350(.dina(w_in147_0[2]),.dinb(n1991),.dout(n1992),.clk(gclk));
	jnot g1351(.din(w_in046_0[2]),.dout(n1993),.clk(gclk));
	jand g1352(.dina(w_in146_0[2]),.dinb(n1993),.dout(n1994),.clk(gclk));
	jor g1353(.dina(n1994),.dinb(w_n1992_0[1]),.dout(n1995),.clk(gclk));
	jor g1354(.dina(n1995),.dinb(n1990),.dout(n1996),.clk(gclk));
	jnot g1355(.din(w_in043_0[2]),.dout(n1997),.clk(gclk));
	jand g1356(.dina(w_in143_0[2]),.dinb(n1997),.dout(n1998),.clk(gclk));
	jnot g1357(.din(w_in042_0[2]),.dout(n1999),.clk(gclk));
	jand g1358(.dina(w_in142_0[2]),.dinb(n1999),.dout(n2000),.clk(gclk));
	jor g1359(.dina(n2000),.dinb(n1998),.dout(n2001),.clk(gclk));
	jnot g1360(.din(w_in044_0[2]),.dout(n2002),.clk(gclk));
	jand g1361(.dina(w_in144_0[2]),.dinb(n2002),.dout(n2003),.clk(gclk));
	jnot g1362(.din(w_in040_0[2]),.dout(n2004),.clk(gclk));
	jand g1363(.dina(w_in140_0[2]),.dinb(n2004),.dout(n2005),.clk(gclk));
	jnot g1364(.din(w_in041_0[2]),.dout(n2006),.clk(gclk));
	jand g1365(.dina(w_in141_0[2]),.dinb(n2006),.dout(n2007),.clk(gclk));
	jor g1366(.dina(w_n2007_0[1]),.dinb(n2005),.dout(n2008),.clk(gclk));
	jor g1367(.dina(n2008),.dinb(w_n2003_0[1]),.dout(n2009),.clk(gclk));
	jor g1368(.dina(n2009),.dinb(w_n2001_0[1]),.dout(n2010),.clk(gclk));
	jor g1369(.dina(n2010),.dinb(w_n1996_0[1]),.dout(n2011),.clk(gclk));
	jnot g1370(.din(w_n2011_0[1]),.dout(n2012),.clk(gclk));
	jand g1371(.dina(n2012),.dinb(n1988),.dout(n2013),.clk(gclk));
	jnot g1372(.din(w_n1996_0[0]),.dout(n2014),.clk(gclk));
	jnot g1373(.din(w_n2003_0[0]),.dout(n2015),.clk(gclk));
	jnot g1374(.din(w_in143_0[1]),.dout(n2016),.clk(gclk));
	jand g1375(.dina(n2016),.dinb(w_in043_0[1]),.dout(n2017),.clk(gclk));
	jnot g1376(.din(w_n2001_0[0]),.dout(n2018),.clk(gclk));
	jnot g1377(.din(w_n2007_0[0]),.dout(n2019),.clk(gclk));
	jnot g1378(.din(w_in140_0[1]),.dout(n2020),.clk(gclk));
	jand g1379(.dina(n2020),.dinb(w_in040_0[1]),.dout(n2021),.clk(gclk));
	jand g1380(.dina(n2021),.dinb(n2019),.dout(n2022),.clk(gclk));
	jnot g1381(.din(w_in141_0[1]),.dout(n2023),.clk(gclk));
	jand g1382(.dina(n2023),.dinb(w_in041_0[1]),.dout(n2024),.clk(gclk));
	jnot g1383(.din(w_in142_0[1]),.dout(n2025),.clk(gclk));
	jand g1384(.dina(n2025),.dinb(w_in042_0[1]),.dout(n2026),.clk(gclk));
	jor g1385(.dina(n2026),.dinb(n2024),.dout(n2027),.clk(gclk));
	jor g1386(.dina(n2027),.dinb(n2022),.dout(n2028),.clk(gclk));
	jand g1387(.dina(n2028),.dinb(n2018),.dout(n2029),.clk(gclk));
	jor g1388(.dina(n2029),.dinb(n2017),.dout(n2030),.clk(gclk));
	jand g1389(.dina(n2030),.dinb(n2015),.dout(n2031),.clk(gclk));
	jnot g1390(.din(w_in144_0[1]),.dout(n2032),.clk(gclk));
	jand g1391(.dina(n2032),.dinb(w_in044_0[1]),.dout(n2033),.clk(gclk));
	jnot g1392(.din(w_in145_0[1]),.dout(n2034),.clk(gclk));
	jand g1393(.dina(n2034),.dinb(w_in045_0[1]),.dout(n2035),.clk(gclk));
	jor g1394(.dina(n2035),.dinb(n2033),.dout(n2036),.clk(gclk));
	jor g1395(.dina(n2036),.dinb(n2031),.dout(n2037),.clk(gclk));
	jand g1396(.dina(n2037),.dinb(n2014),.dout(n2038),.clk(gclk));
	jnot g1397(.din(w_n1992_0[0]),.dout(n2039),.clk(gclk));
	jnot g1398(.din(w_in146_0[1]),.dout(n2040),.clk(gclk));
	jand g1399(.dina(n2040),.dinb(w_in046_0[1]),.dout(n2041),.clk(gclk));
	jand g1400(.dina(n2041),.dinb(n2039),.dout(n2042),.clk(gclk));
	jnot g1401(.din(w_in147_0[1]),.dout(n2043),.clk(gclk));
	jand g1402(.dina(n2043),.dinb(w_in047_0[1]),.dout(n2044),.clk(gclk));
	jor g1403(.dina(n2044),.dinb(n2042),.dout(n2045),.clk(gclk));
	jor g1404(.dina(n2045),.dinb(n2038),.dout(n2046),.clk(gclk));
	jor g1405(.dina(w_n2046_0[1]),.dinb(n2013),.dout(n2047),.clk(gclk));
	jnot g1406(.din(w_in152_0[1]),.dout(n2048),.clk(gclk));
	jnot g1407(.din(w_in053_0[2]),.dout(n2049),.clk(gclk));
	jand g1408(.dina(w_in153_0[2]),.dinb(n2049),.dout(n2050),.clk(gclk));
	jnot g1409(.din(n2050),.dout(n2051),.clk(gclk));
	jand g1410(.dina(w_n2051_0[1]),.dinb(n2048),.dout(n2052),.clk(gclk));
	jand g1411(.dina(w_n2051_0[0]),.dinb(w_in052_0[2]),.dout(n2053),.clk(gclk));
	jor g1412(.dina(n2053),.dinb(w_n2052_0[1]),.dout(n2054),.clk(gclk));
	jnot g1413(.din(w_n2054_0[1]),.dout(n2055),.clk(gclk));
	jnot g1414(.din(w_in055_0[2]),.dout(n2056),.clk(gclk));
	jand g1415(.dina(w_in155_0[2]),.dinb(n2056),.dout(n2057),.clk(gclk));
	jnot g1416(.din(w_in054_0[2]),.dout(n2058),.clk(gclk));
	jand g1417(.dina(w_in154_0[2]),.dinb(n2058),.dout(n2059),.clk(gclk));
	jor g1418(.dina(n2059),.dinb(n2057),.dout(n2060),.clk(gclk));
	jnot g1419(.din(w_in051_0[2]),.dout(n2061),.clk(gclk));
	jand g1420(.dina(w_in151_0[2]),.dinb(n2061),.dout(n2062),.clk(gclk));
	jnot g1421(.din(w_in050_0[2]),.dout(n2063),.clk(gclk));
	jand g1422(.dina(w_in150_0[2]),.dinb(n2063),.dout(n2064),.clk(gclk));
	jor g1423(.dina(n2064),.dinb(n2062),.dout(n2065),.clk(gclk));
	jnot g1424(.din(w_in048_0[2]),.dout(n2066),.clk(gclk));
	jand g1425(.dina(w_in148_0[2]),.dinb(n2066),.dout(n2067),.clk(gclk));
	jnot g1426(.din(w_in049_0[2]),.dout(n2068),.clk(gclk));
	jand g1427(.dina(w_in149_0[2]),.dinb(n2068),.dout(n2069),.clk(gclk));
	jor g1428(.dina(w_n2069_0[1]),.dinb(n2067),.dout(n2070),.clk(gclk));
	jor g1429(.dina(n2070),.dinb(w_n2065_0[1]),.dout(n2071),.clk(gclk));
	jor g1430(.dina(n2071),.dinb(w_n2060_0[1]),.dout(n2072),.clk(gclk));
	jor g1431(.dina(n2072),.dinb(n2055),.dout(n2073),.clk(gclk));
	jnot g1432(.din(w_n2073_0[1]),.dout(n2074),.clk(gclk));
	jand g1433(.dina(n2074),.dinb(n2047),.dout(n2075),.clk(gclk));
	jnot g1434(.din(w_in155_0[1]),.dout(n2076),.clk(gclk));
	jand g1435(.dina(n2076),.dinb(w_in055_0[1]),.dout(n2077),.clk(gclk));
	jnot g1436(.din(w_n2060_0[0]),.dout(n2078),.clk(gclk));
	jnot g1437(.din(w_in151_0[1]),.dout(n2079),.clk(gclk));
	jand g1438(.dina(n2079),.dinb(w_in051_0[1]),.dout(n2080),.clk(gclk));
	jnot g1439(.din(w_n2065_0[0]),.dout(n2081),.clk(gclk));
	jnot g1440(.din(w_n2069_0[0]),.dout(n2082),.clk(gclk));
	jnot g1441(.din(w_in148_0[1]),.dout(n2083),.clk(gclk));
	jand g1442(.dina(n2083),.dinb(w_in048_0[1]),.dout(n2084),.clk(gclk));
	jand g1443(.dina(n2084),.dinb(n2082),.dout(n2085),.clk(gclk));
	jnot g1444(.din(w_in149_0[1]),.dout(n2086),.clk(gclk));
	jand g1445(.dina(n2086),.dinb(w_in049_0[1]),.dout(n2087),.clk(gclk));
	jnot g1446(.din(w_in150_0[1]),.dout(n2088),.clk(gclk));
	jand g1447(.dina(n2088),.dinb(w_in050_0[1]),.dout(n2089),.clk(gclk));
	jor g1448(.dina(n2089),.dinb(n2087),.dout(n2090),.clk(gclk));
	jor g1449(.dina(n2090),.dinb(n2085),.dout(n2091),.clk(gclk));
	jand g1450(.dina(n2091),.dinb(n2081),.dout(n2092),.clk(gclk));
	jor g1451(.dina(n2092),.dinb(n2080),.dout(n2093),.clk(gclk));
	jand g1452(.dina(n2093),.dinb(w_n2054_0[0]),.dout(n2094),.clk(gclk));
	jand g1453(.dina(w_n2052_0[0]),.dinb(w_in052_0[1]),.dout(n2095),.clk(gclk));
	jnot g1454(.din(w_in153_0[1]),.dout(n2096),.clk(gclk));
	jand g1455(.dina(n2096),.dinb(w_in053_0[1]),.dout(n2097),.clk(gclk));
	jnot g1456(.din(w_in154_0[1]),.dout(n2098),.clk(gclk));
	jand g1457(.dina(n2098),.dinb(w_in054_0[1]),.dout(n2099),.clk(gclk));
	jor g1458(.dina(n2099),.dinb(n2097),.dout(n2100),.clk(gclk));
	jor g1459(.dina(n2100),.dinb(n2095),.dout(n2101),.clk(gclk));
	jor g1460(.dina(n2101),.dinb(n2094),.dout(n2102),.clk(gclk));
	jand g1461(.dina(n2102),.dinb(n2078),.dout(n2103),.clk(gclk));
	jor g1462(.dina(n2103),.dinb(n2077),.dout(n2104),.clk(gclk));
	jor g1463(.dina(w_n2104_0[1]),.dinb(n2075),.dout(n2105),.clk(gclk));
	jnot g1464(.din(w_in061_0[2]),.dout(n2106),.clk(gclk));
	jand g1465(.dina(w_in161_0[2]),.dinb(n2106),.dout(n2107),.clk(gclk));
	jnot g1466(.din(w_in063_0[2]),.dout(n2108),.clk(gclk));
	jand g1467(.dina(w_in163_0[2]),.dinb(n2108),.dout(n2109),.clk(gclk));
	jnot g1468(.din(w_in062_0[2]),.dout(n2110),.clk(gclk));
	jand g1469(.dina(w_in162_0[2]),.dinb(n2110),.dout(n2111),.clk(gclk));
	jor g1470(.dina(n2111),.dinb(w_n2109_0[1]),.dout(n2112),.clk(gclk));
	jor g1471(.dina(n2112),.dinb(n2107),.dout(n2113),.clk(gclk));
	jnot g1472(.din(w_in059_0[2]),.dout(n2114),.clk(gclk));
	jand g1473(.dina(w_in159_0[2]),.dinb(n2114),.dout(n2115),.clk(gclk));
	jnot g1474(.din(w_in058_0[2]),.dout(n2116),.clk(gclk));
	jand g1475(.dina(w_in158_0[2]),.dinb(n2116),.dout(n2117),.clk(gclk));
	jor g1476(.dina(n2117),.dinb(n2115),.dout(n2118),.clk(gclk));
	jnot g1477(.din(w_in060_0[2]),.dout(n2119),.clk(gclk));
	jand g1478(.dina(w_in160_0[2]),.dinb(n2119),.dout(n2120),.clk(gclk));
	jnot g1479(.din(w_in056_0[2]),.dout(n2121),.clk(gclk));
	jand g1480(.dina(w_in156_0[2]),.dinb(n2121),.dout(n2122),.clk(gclk));
	jnot g1481(.din(w_in057_0[2]),.dout(n2123),.clk(gclk));
	jand g1482(.dina(w_in157_0[2]),.dinb(n2123),.dout(n2124),.clk(gclk));
	jor g1483(.dina(w_n2124_0[1]),.dinb(n2122),.dout(n2125),.clk(gclk));
	jor g1484(.dina(n2125),.dinb(w_n2120_0[1]),.dout(n2126),.clk(gclk));
	jor g1485(.dina(n2126),.dinb(w_n2118_0[1]),.dout(n2127),.clk(gclk));
	jor g1486(.dina(n2127),.dinb(w_n2113_0[1]),.dout(n2128),.clk(gclk));
	jnot g1487(.din(w_n2128_0[1]),.dout(n2129),.clk(gclk));
	jand g1488(.dina(n2129),.dinb(n2105),.dout(n2130),.clk(gclk));
	jnot g1489(.din(w_n2113_0[0]),.dout(n2131),.clk(gclk));
	jnot g1490(.din(w_n2120_0[0]),.dout(n2132),.clk(gclk));
	jnot g1491(.din(w_in159_0[1]),.dout(n2133),.clk(gclk));
	jand g1492(.dina(n2133),.dinb(w_in059_0[1]),.dout(n2134),.clk(gclk));
	jnot g1493(.din(w_n2118_0[0]),.dout(n2135),.clk(gclk));
	jnot g1494(.din(w_n2124_0[0]),.dout(n2136),.clk(gclk));
	jnot g1495(.din(w_in156_0[1]),.dout(n2137),.clk(gclk));
	jand g1496(.dina(n2137),.dinb(w_in056_0[1]),.dout(n2138),.clk(gclk));
	jand g1497(.dina(n2138),.dinb(n2136),.dout(n2139),.clk(gclk));
	jnot g1498(.din(w_in157_0[1]),.dout(n2140),.clk(gclk));
	jand g1499(.dina(n2140),.dinb(w_in057_0[1]),.dout(n2141),.clk(gclk));
	jnot g1500(.din(w_in158_0[1]),.dout(n2142),.clk(gclk));
	jand g1501(.dina(n2142),.dinb(w_in058_0[1]),.dout(n2143),.clk(gclk));
	jor g1502(.dina(n2143),.dinb(n2141),.dout(n2144),.clk(gclk));
	jor g1503(.dina(n2144),.dinb(n2139),.dout(n2145),.clk(gclk));
	jand g1504(.dina(n2145),.dinb(n2135),.dout(n2146),.clk(gclk));
	jor g1505(.dina(n2146),.dinb(n2134),.dout(n2147),.clk(gclk));
	jand g1506(.dina(n2147),.dinb(n2132),.dout(n2148),.clk(gclk));
	jnot g1507(.din(w_in160_0[1]),.dout(n2149),.clk(gclk));
	jand g1508(.dina(n2149),.dinb(w_in060_0[1]),.dout(n2150),.clk(gclk));
	jnot g1509(.din(w_in161_0[1]),.dout(n2151),.clk(gclk));
	jand g1510(.dina(n2151),.dinb(w_in061_0[1]),.dout(n2152),.clk(gclk));
	jor g1511(.dina(n2152),.dinb(n2150),.dout(n2153),.clk(gclk));
	jor g1512(.dina(n2153),.dinb(n2148),.dout(n2154),.clk(gclk));
	jand g1513(.dina(n2154),.dinb(n2131),.dout(n2155),.clk(gclk));
	jnot g1514(.din(w_n2109_0[0]),.dout(n2156),.clk(gclk));
	jnot g1515(.din(w_in162_0[1]),.dout(n2157),.clk(gclk));
	jand g1516(.dina(n2157),.dinb(w_in062_0[1]),.dout(n2158),.clk(gclk));
	jand g1517(.dina(n2158),.dinb(n2156),.dout(n2159),.clk(gclk));
	jnot g1518(.din(w_in163_0[1]),.dout(n2160),.clk(gclk));
	jand g1519(.dina(n2160),.dinb(w_in063_0[1]),.dout(n2161),.clk(gclk));
	jor g1520(.dina(n2161),.dinb(n2159),.dout(n2162),.clk(gclk));
	jor g1521(.dina(n2162),.dinb(n2155),.dout(n2163),.clk(gclk));
	jor g1522(.dina(w_n2163_0[1]),.dinb(n2130),.dout(n2164),.clk(gclk));
	jnot g1523(.din(w_in067_0[2]),.dout(n2165),.clk(gclk));
	jand g1524(.dina(w_in167_0[2]),.dinb(n2165),.dout(n2166),.clk(gclk));
	jnot g1525(.din(w_in066_0[2]),.dout(n2167),.clk(gclk));
	jand g1526(.dina(w_in166_0[2]),.dinb(n2167),.dout(n2168),.clk(gclk));
	jor g1527(.dina(n2168),.dinb(n2166),.dout(n2169),.clk(gclk));
	jnot g1528(.din(w_in065_0[2]),.dout(n2170),.clk(gclk));
	jand g1529(.dina(w_in165_0[2]),.dinb(n2170),.dout(n2171),.clk(gclk));
	jnot g1530(.din(w_in064_0[2]),.dout(n2172),.clk(gclk));
	jand g1531(.dina(w_in164_0[2]),.dinb(n2172),.dout(n2173),.clk(gclk));
	jor g1532(.dina(n2173),.dinb(w_n2171_0[1]),.dout(n2174),.clk(gclk));
	jor g1533(.dina(n2174),.dinb(w_n2169_0[1]),.dout(n2175),.clk(gclk));
	jnot g1534(.din(w_n2175_0[1]),.dout(n2176),.clk(gclk));
	jand g1535(.dina(n2176),.dinb(n2164),.dout(n2177),.clk(gclk));
	jnot g1536(.din(w_in167_0[1]),.dout(n2178),.clk(gclk));
	jand g1537(.dina(n2178),.dinb(w_in067_0[1]),.dout(n2179),.clk(gclk));
	jnot g1538(.din(w_n2169_0[0]),.dout(n2180),.clk(gclk));
	jnot g1539(.din(w_n2171_0[0]),.dout(n2181),.clk(gclk));
	jnot g1540(.din(w_in164_0[1]),.dout(n2182),.clk(gclk));
	jand g1541(.dina(n2182),.dinb(w_in064_0[1]),.dout(n2183),.clk(gclk));
	jand g1542(.dina(n2183),.dinb(n2181),.dout(n2184),.clk(gclk));
	jnot g1543(.din(w_in165_0[1]),.dout(n2185),.clk(gclk));
	jand g1544(.dina(n2185),.dinb(w_in065_0[1]),.dout(n2186),.clk(gclk));
	jnot g1545(.din(w_in166_0[1]),.dout(n2187),.clk(gclk));
	jand g1546(.dina(n2187),.dinb(w_in066_0[1]),.dout(n2188),.clk(gclk));
	jor g1547(.dina(n2188),.dinb(n2186),.dout(n2189),.clk(gclk));
	jor g1548(.dina(n2189),.dinb(n2184),.dout(n2190),.clk(gclk));
	jand g1549(.dina(n2190),.dinb(n2180),.dout(n2191),.clk(gclk));
	jor g1550(.dina(n2191),.dinb(n2179),.dout(n2192),.clk(gclk));
	jor g1551(.dina(w_n2192_0[1]),.dinb(n2177),.dout(n2193),.clk(gclk));
	jnot g1552(.din(w_in068_0[2]),.dout(n2194),.clk(gclk));
	jand g1553(.dina(w_in168_0[2]),.dinb(n2194),.dout(n2195),.clk(gclk));
	jnot g1554(.din(w_in069_0[2]),.dout(n2196),.clk(gclk));
	jand g1555(.dina(w_in169_0[2]),.dinb(n2196),.dout(n2197),.clk(gclk));
	jnot g1556(.din(w_in071_0[2]),.dout(n2198),.clk(gclk));
	jand g1557(.dina(w_in171_0[2]),.dinb(n2198),.dout(n2199),.clk(gclk));
	jnot g1558(.din(w_in070_0[2]),.dout(n2200),.clk(gclk));
	jand g1559(.dina(w_in170_0[2]),.dinb(n2200),.dout(n2201),.clk(gclk));
	jor g1560(.dina(n2201),.dinb(w_n2199_0[1]),.dout(n2202),.clk(gclk));
	jor g1561(.dina(n2202),.dinb(n2197),.dout(n2203),.clk(gclk));
	jor g1562(.dina(w_n2203_0[1]),.dinb(n2195),.dout(n2204),.clk(gclk));
	jnot g1563(.din(w_n2204_0[1]),.dout(n2205),.clk(gclk));
	jand g1564(.dina(n2205),.dinb(n2193),.dout(n2206),.clk(gclk));
	jnot g1565(.din(w_n2203_0[0]),.dout(n2207),.clk(gclk));
	jnot g1566(.din(w_in169_0[1]),.dout(n2208),.clk(gclk));
	jand g1567(.dina(n2208),.dinb(w_in069_0[1]),.dout(n2209),.clk(gclk));
	jnot g1568(.din(w_in168_0[1]),.dout(n2210),.clk(gclk));
	jand g1569(.dina(n2210),.dinb(w_in068_0[1]),.dout(n2211),.clk(gclk));
	jor g1570(.dina(n2211),.dinb(n2209),.dout(n2212),.clk(gclk));
	jand g1571(.dina(n2212),.dinb(n2207),.dout(n2213),.clk(gclk));
	jnot g1572(.din(w_in171_0[1]),.dout(n2214),.clk(gclk));
	jand g1573(.dina(n2214),.dinb(w_in071_0[1]),.dout(n2215),.clk(gclk));
	jnot g1574(.din(w_n2199_0[0]),.dout(n2216),.clk(gclk));
	jnot g1575(.din(w_in170_0[1]),.dout(n2217),.clk(gclk));
	jand g1576(.dina(n2217),.dinb(w_in070_0[1]),.dout(n2218),.clk(gclk));
	jand g1577(.dina(n2218),.dinb(n2216),.dout(n2219),.clk(gclk));
	jor g1578(.dina(n2219),.dinb(n2215),.dout(n2220),.clk(gclk));
	jor g1579(.dina(n2220),.dinb(n2213),.dout(n2221),.clk(gclk));
	jor g1580(.dina(w_n2221_0[1]),.dinb(n2206),.dout(n2222),.clk(gclk));
	jnot g1581(.din(w_in075_0[2]),.dout(n2223),.clk(gclk));
	jand g1582(.dina(w_in175_0[2]),.dinb(n2223),.dout(n2224),.clk(gclk));
	jnot g1583(.din(w_in074_0[2]),.dout(n2225),.clk(gclk));
	jand g1584(.dina(w_in174_0[2]),.dinb(n2225),.dout(n2226),.clk(gclk));
	jor g1585(.dina(n2226),.dinb(n2224),.dout(n2227),.clk(gclk));
	jnot g1586(.din(w_in073_0[2]),.dout(n2228),.clk(gclk));
	jand g1587(.dina(w_in173_0[2]),.dinb(n2228),.dout(n2229),.clk(gclk));
	jnot g1588(.din(w_in072_0[2]),.dout(n2230),.clk(gclk));
	jand g1589(.dina(w_in172_0[2]),.dinb(n2230),.dout(n2231),.clk(gclk));
	jor g1590(.dina(n2231),.dinb(w_n2229_0[1]),.dout(n2232),.clk(gclk));
	jor g1591(.dina(n2232),.dinb(w_n2227_0[1]),.dout(n2233),.clk(gclk));
	jnot g1592(.din(w_n2233_0[1]),.dout(n2234),.clk(gclk));
	jand g1593(.dina(n2234),.dinb(n2222),.dout(n2235),.clk(gclk));
	jnot g1594(.din(w_in175_0[1]),.dout(n2236),.clk(gclk));
	jand g1595(.dina(n2236),.dinb(w_in075_0[1]),.dout(n2237),.clk(gclk));
	jnot g1596(.din(w_n2227_0[0]),.dout(n2238),.clk(gclk));
	jnot g1597(.din(w_n2229_0[0]),.dout(n2239),.clk(gclk));
	jnot g1598(.din(w_in172_0[1]),.dout(n2240),.clk(gclk));
	jand g1599(.dina(n2240),.dinb(w_in072_0[1]),.dout(n2241),.clk(gclk));
	jand g1600(.dina(n2241),.dinb(n2239),.dout(n2242),.clk(gclk));
	jnot g1601(.din(w_in173_0[1]),.dout(n2243),.clk(gclk));
	jand g1602(.dina(n2243),.dinb(w_in073_0[1]),.dout(n2244),.clk(gclk));
	jnot g1603(.din(w_in174_0[1]),.dout(n2245),.clk(gclk));
	jand g1604(.dina(n2245),.dinb(w_in074_0[1]),.dout(n2246),.clk(gclk));
	jor g1605(.dina(n2246),.dinb(n2244),.dout(n2247),.clk(gclk));
	jor g1606(.dina(n2247),.dinb(n2242),.dout(n2248),.clk(gclk));
	jand g1607(.dina(n2248),.dinb(n2238),.dout(n2249),.clk(gclk));
	jor g1608(.dina(n2249),.dinb(n2237),.dout(n2250),.clk(gclk));
	jor g1609(.dina(w_n2250_0[1]),.dinb(n2235),.dout(n2251),.clk(gclk));
	jnot g1610(.din(w_in076_0[2]),.dout(n2252),.clk(gclk));
	jand g1611(.dina(w_in176_0[2]),.dinb(n2252),.dout(n2253),.clk(gclk));
	jnot g1612(.din(w_in077_0[2]),.dout(n2254),.clk(gclk));
	jand g1613(.dina(w_in177_0[2]),.dinb(n2254),.dout(n2255),.clk(gclk));
	jnot g1614(.din(w_in079_0[2]),.dout(n2256),.clk(gclk));
	jand g1615(.dina(w_in179_0[2]),.dinb(n2256),.dout(n2257),.clk(gclk));
	jnot g1616(.din(w_in078_0[2]),.dout(n2258),.clk(gclk));
	jand g1617(.dina(w_in178_0[2]),.dinb(n2258),.dout(n2259),.clk(gclk));
	jor g1618(.dina(n2259),.dinb(w_n2257_0[1]),.dout(n2260),.clk(gclk));
	jor g1619(.dina(n2260),.dinb(n2255),.dout(n2261),.clk(gclk));
	jor g1620(.dina(w_n2261_0[1]),.dinb(n2253),.dout(n2262),.clk(gclk));
	jnot g1621(.din(w_n2262_0[1]),.dout(n2263),.clk(gclk));
	jand g1622(.dina(n2263),.dinb(n2251),.dout(n2264),.clk(gclk));
	jnot g1623(.din(w_n2261_0[0]),.dout(n2265),.clk(gclk));
	jnot g1624(.din(w_in177_0[1]),.dout(n2266),.clk(gclk));
	jand g1625(.dina(n2266),.dinb(w_in077_0[1]),.dout(n2267),.clk(gclk));
	jnot g1626(.din(w_in176_0[1]),.dout(n2268),.clk(gclk));
	jand g1627(.dina(n2268),.dinb(w_in076_0[1]),.dout(n2269),.clk(gclk));
	jor g1628(.dina(n2269),.dinb(n2267),.dout(n2270),.clk(gclk));
	jand g1629(.dina(n2270),.dinb(n2265),.dout(n2271),.clk(gclk));
	jnot g1630(.din(w_in179_0[1]),.dout(n2272),.clk(gclk));
	jand g1631(.dina(n2272),.dinb(w_in079_0[1]),.dout(n2273),.clk(gclk));
	jnot g1632(.din(w_n2257_0[0]),.dout(n2274),.clk(gclk));
	jnot g1633(.din(w_in178_0[1]),.dout(n2275),.clk(gclk));
	jand g1634(.dina(n2275),.dinb(w_in078_0[1]),.dout(n2276),.clk(gclk));
	jand g1635(.dina(n2276),.dinb(n2274),.dout(n2277),.clk(gclk));
	jor g1636(.dina(n2277),.dinb(n2273),.dout(n2278),.clk(gclk));
	jor g1637(.dina(n2278),.dinb(n2271),.dout(n2279),.clk(gclk));
	jor g1638(.dina(w_n2279_0[1]),.dinb(n2264),.dout(n2280),.clk(gclk));
	jnot g1639(.din(w_in083_0[2]),.dout(n2281),.clk(gclk));
	jand g1640(.dina(w_in183_0[2]),.dinb(n2281),.dout(n2282),.clk(gclk));
	jnot g1641(.din(w_in082_0[2]),.dout(n2283),.clk(gclk));
	jand g1642(.dina(w_in182_0[2]),.dinb(n2283),.dout(n2284),.clk(gclk));
	jor g1643(.dina(n2284),.dinb(n2282),.dout(n2285),.clk(gclk));
	jnot g1644(.din(w_in081_0[2]),.dout(n2286),.clk(gclk));
	jand g1645(.dina(w_in181_0[2]),.dinb(n2286),.dout(n2287),.clk(gclk));
	jnot g1646(.din(w_in080_0[2]),.dout(n2288),.clk(gclk));
	jand g1647(.dina(w_in180_0[2]),.dinb(n2288),.dout(n2289),.clk(gclk));
	jor g1648(.dina(n2289),.dinb(w_n2287_0[1]),.dout(n2290),.clk(gclk));
	jor g1649(.dina(n2290),.dinb(w_n2285_0[1]),.dout(n2291),.clk(gclk));
	jnot g1650(.din(w_n2291_0[1]),.dout(n2292),.clk(gclk));
	jand g1651(.dina(n2292),.dinb(n2280),.dout(n2293),.clk(gclk));
	jnot g1652(.din(w_in183_0[1]),.dout(n2294),.clk(gclk));
	jand g1653(.dina(n2294),.dinb(w_in083_0[1]),.dout(n2295),.clk(gclk));
	jnot g1654(.din(w_n2285_0[0]),.dout(n2296),.clk(gclk));
	jnot g1655(.din(w_n2287_0[0]),.dout(n2297),.clk(gclk));
	jnot g1656(.din(w_in180_0[1]),.dout(n2298),.clk(gclk));
	jand g1657(.dina(n2298),.dinb(w_in080_0[1]),.dout(n2299),.clk(gclk));
	jand g1658(.dina(n2299),.dinb(n2297),.dout(n2300),.clk(gclk));
	jnot g1659(.din(w_in181_0[1]),.dout(n2301),.clk(gclk));
	jand g1660(.dina(n2301),.dinb(w_in081_0[1]),.dout(n2302),.clk(gclk));
	jnot g1661(.din(w_in182_0[1]),.dout(n2303),.clk(gclk));
	jand g1662(.dina(n2303),.dinb(w_in082_0[1]),.dout(n2304),.clk(gclk));
	jor g1663(.dina(n2304),.dinb(n2302),.dout(n2305),.clk(gclk));
	jor g1664(.dina(n2305),.dinb(n2300),.dout(n2306),.clk(gclk));
	jand g1665(.dina(n2306),.dinb(n2296),.dout(n2307),.clk(gclk));
	jor g1666(.dina(n2307),.dinb(n2295),.dout(n2308),.clk(gclk));
	jor g1667(.dina(w_n2308_0[1]),.dinb(n2293),.dout(n2309),.clk(gclk));
	jnot g1668(.din(w_in084_0[2]),.dout(n2310),.clk(gclk));
	jand g1669(.dina(w_in184_0[2]),.dinb(n2310),.dout(n2311),.clk(gclk));
	jnot g1670(.din(w_in085_0[2]),.dout(n2312),.clk(gclk));
	jand g1671(.dina(w_in185_0[2]),.dinb(n2312),.dout(n2313),.clk(gclk));
	jnot g1672(.din(w_in087_0[2]),.dout(n2314),.clk(gclk));
	jand g1673(.dina(w_in187_0[2]),.dinb(n2314),.dout(n2315),.clk(gclk));
	jnot g1674(.din(w_in086_0[2]),.dout(n2316),.clk(gclk));
	jand g1675(.dina(w_in186_0[2]),.dinb(n2316),.dout(n2317),.clk(gclk));
	jor g1676(.dina(n2317),.dinb(w_n2315_0[1]),.dout(n2318),.clk(gclk));
	jor g1677(.dina(n2318),.dinb(n2313),.dout(n2319),.clk(gclk));
	jor g1678(.dina(w_n2319_0[1]),.dinb(n2311),.dout(n2320),.clk(gclk));
	jnot g1679(.din(w_n2320_0[1]),.dout(n2321),.clk(gclk));
	jand g1680(.dina(n2321),.dinb(n2309),.dout(n2322),.clk(gclk));
	jnot g1681(.din(w_n2319_0[0]),.dout(n2323),.clk(gclk));
	jnot g1682(.din(w_in185_0[1]),.dout(n2324),.clk(gclk));
	jand g1683(.dina(n2324),.dinb(w_in085_0[1]),.dout(n2325),.clk(gclk));
	jnot g1684(.din(w_in184_0[1]),.dout(n2326),.clk(gclk));
	jand g1685(.dina(n2326),.dinb(w_in084_0[1]),.dout(n2327),.clk(gclk));
	jor g1686(.dina(n2327),.dinb(n2325),.dout(n2328),.clk(gclk));
	jand g1687(.dina(n2328),.dinb(n2323),.dout(n2329),.clk(gclk));
	jnot g1688(.din(w_in187_0[1]),.dout(n2330),.clk(gclk));
	jand g1689(.dina(n2330),.dinb(w_in087_0[1]),.dout(n2331),.clk(gclk));
	jnot g1690(.din(w_n2315_0[0]),.dout(n2332),.clk(gclk));
	jnot g1691(.din(w_in186_0[1]),.dout(n2333),.clk(gclk));
	jand g1692(.dina(n2333),.dinb(w_in086_0[1]),.dout(n2334),.clk(gclk));
	jand g1693(.dina(n2334),.dinb(n2332),.dout(n2335),.clk(gclk));
	jor g1694(.dina(n2335),.dinb(n2331),.dout(n2336),.clk(gclk));
	jor g1695(.dina(n2336),.dinb(n2329),.dout(n2337),.clk(gclk));
	jor g1696(.dina(w_n2337_0[1]),.dinb(n2322),.dout(n2338),.clk(gclk));
	jnot g1697(.din(w_in091_0[2]),.dout(n2339),.clk(gclk));
	jand g1698(.dina(w_in191_0[2]),.dinb(n2339),.dout(n2340),.clk(gclk));
	jnot g1699(.din(w_in090_0[2]),.dout(n2341),.clk(gclk));
	jand g1700(.dina(w_in190_0[2]),.dinb(n2341),.dout(n2342),.clk(gclk));
	jor g1701(.dina(n2342),.dinb(n2340),.dout(n2343),.clk(gclk));
	jnot g1702(.din(w_in089_0[2]),.dout(n2344),.clk(gclk));
	jand g1703(.dina(w_in189_0[2]),.dinb(n2344),.dout(n2345),.clk(gclk));
	jnot g1704(.din(w_in088_0[2]),.dout(n2346),.clk(gclk));
	jand g1705(.dina(w_in188_0[2]),.dinb(n2346),.dout(n2347),.clk(gclk));
	jor g1706(.dina(n2347),.dinb(w_n2345_0[1]),.dout(n2348),.clk(gclk));
	jor g1707(.dina(n2348),.dinb(w_n2343_0[1]),.dout(n2349),.clk(gclk));
	jnot g1708(.din(w_n2349_0[1]),.dout(n2350),.clk(gclk));
	jand g1709(.dina(n2350),.dinb(n2338),.dout(n2351),.clk(gclk));
	jnot g1710(.din(w_in191_0[1]),.dout(n2352),.clk(gclk));
	jand g1711(.dina(n2352),.dinb(w_in091_0[1]),.dout(n2353),.clk(gclk));
	jnot g1712(.din(w_n2343_0[0]),.dout(n2354),.clk(gclk));
	jnot g1713(.din(w_n2345_0[0]),.dout(n2355),.clk(gclk));
	jnot g1714(.din(w_in188_0[1]),.dout(n2356),.clk(gclk));
	jand g1715(.dina(n2356),.dinb(w_in088_0[1]),.dout(n2357),.clk(gclk));
	jand g1716(.dina(n2357),.dinb(n2355),.dout(n2358),.clk(gclk));
	jnot g1717(.din(w_in189_0[1]),.dout(n2359),.clk(gclk));
	jand g1718(.dina(n2359),.dinb(w_in089_0[1]),.dout(n2360),.clk(gclk));
	jnot g1719(.din(w_in190_0[1]),.dout(n2361),.clk(gclk));
	jand g1720(.dina(n2361),.dinb(w_in090_0[1]),.dout(n2362),.clk(gclk));
	jor g1721(.dina(n2362),.dinb(n2360),.dout(n2363),.clk(gclk));
	jor g1722(.dina(n2363),.dinb(n2358),.dout(n2364),.clk(gclk));
	jand g1723(.dina(n2364),.dinb(n2354),.dout(n2365),.clk(gclk));
	jor g1724(.dina(n2365),.dinb(n2353),.dout(n2366),.clk(gclk));
	jor g1725(.dina(w_n2366_0[1]),.dinb(n2351),.dout(n2367),.clk(gclk));
	jnot g1726(.din(w_in092_0[2]),.dout(n2368),.clk(gclk));
	jand g1727(.dina(w_in192_0[2]),.dinb(n2368),.dout(n2369),.clk(gclk));
	jnot g1728(.din(w_in093_0[2]),.dout(n2370),.clk(gclk));
	jand g1729(.dina(w_in193_0[2]),.dinb(n2370),.dout(n2371),.clk(gclk));
	jnot g1730(.din(w_in095_0[2]),.dout(n2372),.clk(gclk));
	jand g1731(.dina(w_in195_0[2]),.dinb(n2372),.dout(n2373),.clk(gclk));
	jnot g1732(.din(w_in094_0[2]),.dout(n2374),.clk(gclk));
	jand g1733(.dina(w_in194_0[2]),.dinb(n2374),.dout(n2375),.clk(gclk));
	jor g1734(.dina(n2375),.dinb(w_n2373_0[1]),.dout(n2376),.clk(gclk));
	jor g1735(.dina(n2376),.dinb(n2371),.dout(n2377),.clk(gclk));
	jor g1736(.dina(w_n2377_0[1]),.dinb(n2369),.dout(n2378),.clk(gclk));
	jnot g1737(.din(w_n2378_0[1]),.dout(n2379),.clk(gclk));
	jand g1738(.dina(n2379),.dinb(n2367),.dout(n2380),.clk(gclk));
	jnot g1739(.din(w_n2377_0[0]),.dout(n2381),.clk(gclk));
	jnot g1740(.din(w_in193_0[1]),.dout(n2382),.clk(gclk));
	jand g1741(.dina(n2382),.dinb(w_in093_0[1]),.dout(n2383),.clk(gclk));
	jnot g1742(.din(w_in192_0[1]),.dout(n2384),.clk(gclk));
	jand g1743(.dina(n2384),.dinb(w_in092_0[1]),.dout(n2385),.clk(gclk));
	jor g1744(.dina(n2385),.dinb(n2383),.dout(n2386),.clk(gclk));
	jand g1745(.dina(n2386),.dinb(n2381),.dout(n2387),.clk(gclk));
	jnot g1746(.din(w_in195_0[1]),.dout(n2388),.clk(gclk));
	jand g1747(.dina(n2388),.dinb(w_in095_0[1]),.dout(n2389),.clk(gclk));
	jnot g1748(.din(w_n2373_0[0]),.dout(n2390),.clk(gclk));
	jnot g1749(.din(w_in194_0[1]),.dout(n2391),.clk(gclk));
	jand g1750(.dina(n2391),.dinb(w_in094_0[1]),.dout(n2392),.clk(gclk));
	jand g1751(.dina(n2392),.dinb(n2390),.dout(n2393),.clk(gclk));
	jor g1752(.dina(n2393),.dinb(n2389),.dout(n2394),.clk(gclk));
	jor g1753(.dina(n2394),.dinb(n2387),.dout(n2395),.clk(gclk));
	jor g1754(.dina(w_n2395_0[1]),.dinb(n2380),.dout(n2396),.clk(gclk));
	jnot g1755(.din(w_in099_0[2]),.dout(n2397),.clk(gclk));
	jand g1756(.dina(w_in199_0[2]),.dinb(n2397),.dout(n2398),.clk(gclk));
	jnot g1757(.din(w_in098_0[2]),.dout(n2399),.clk(gclk));
	jand g1758(.dina(w_in198_0[2]),.dinb(n2399),.dout(n2400),.clk(gclk));
	jor g1759(.dina(n2400),.dinb(n2398),.dout(n2401),.clk(gclk));
	jnot g1760(.din(w_in097_0[2]),.dout(n2402),.clk(gclk));
	jand g1761(.dina(w_in197_0[2]),.dinb(n2402),.dout(n2403),.clk(gclk));
	jnot g1762(.din(w_in096_0[2]),.dout(n2404),.clk(gclk));
	jand g1763(.dina(w_in196_0[2]),.dinb(n2404),.dout(n2405),.clk(gclk));
	jor g1764(.dina(n2405),.dinb(w_n2403_0[1]),.dout(n2406),.clk(gclk));
	jor g1765(.dina(n2406),.dinb(w_n2401_0[1]),.dout(n2407),.clk(gclk));
	jnot g1766(.din(w_n2407_0[1]),.dout(n2408),.clk(gclk));
	jand g1767(.dina(n2408),.dinb(n2396),.dout(n2409),.clk(gclk));
	jnot g1768(.din(w_in199_0[1]),.dout(n2410),.clk(gclk));
	jand g1769(.dina(n2410),.dinb(w_in099_0[1]),.dout(n2411),.clk(gclk));
	jnot g1770(.din(w_n2401_0[0]),.dout(n2412),.clk(gclk));
	jnot g1771(.din(w_n2403_0[0]),.dout(n2413),.clk(gclk));
	jnot g1772(.din(w_in196_0[1]),.dout(n2414),.clk(gclk));
	jand g1773(.dina(n2414),.dinb(w_in096_0[1]),.dout(n2415),.clk(gclk));
	jand g1774(.dina(n2415),.dinb(n2413),.dout(n2416),.clk(gclk));
	jnot g1775(.din(w_in197_0[1]),.dout(n2417),.clk(gclk));
	jand g1776(.dina(n2417),.dinb(w_in097_0[1]),.dout(n2418),.clk(gclk));
	jnot g1777(.din(w_in198_0[1]),.dout(n2419),.clk(gclk));
	jand g1778(.dina(n2419),.dinb(w_in098_0[1]),.dout(n2420),.clk(gclk));
	jor g1779(.dina(n2420),.dinb(n2418),.dout(n2421),.clk(gclk));
	jor g1780(.dina(n2421),.dinb(n2416),.dout(n2422),.clk(gclk));
	jand g1781(.dina(n2422),.dinb(n2412),.dout(n2423),.clk(gclk));
	jor g1782(.dina(n2423),.dinb(n2411),.dout(n2424),.clk(gclk));
	jor g1783(.dina(w_n2424_0[1]),.dinb(n2409),.dout(n2425),.clk(gclk));
	jnot g1784(.din(w_in0100_0[2]),.dout(n2426),.clk(gclk));
	jand g1785(.dina(w_in1100_0[2]),.dinb(n2426),.dout(n2427),.clk(gclk));
	jnot g1786(.din(w_in0101_0[2]),.dout(n2428),.clk(gclk));
	jand g1787(.dina(w_in1101_0[2]),.dinb(n2428),.dout(n2429),.clk(gclk));
	jnot g1788(.din(w_in0103_0[2]),.dout(n2430),.clk(gclk));
	jand g1789(.dina(w_in1103_0[2]),.dinb(n2430),.dout(n2431),.clk(gclk));
	jnot g1790(.din(w_in0102_0[2]),.dout(n2432),.clk(gclk));
	jand g1791(.dina(w_in1102_0[2]),.dinb(n2432),.dout(n2433),.clk(gclk));
	jor g1792(.dina(n2433),.dinb(w_n2431_0[1]),.dout(n2434),.clk(gclk));
	jor g1793(.dina(n2434),.dinb(n2429),.dout(n2435),.clk(gclk));
	jor g1794(.dina(w_n2435_0[1]),.dinb(n2427),.dout(n2436),.clk(gclk));
	jnot g1795(.din(w_n2436_0[1]),.dout(n2437),.clk(gclk));
	jand g1796(.dina(n2437),.dinb(n2425),.dout(n2438),.clk(gclk));
	jnot g1797(.din(w_n2435_0[0]),.dout(n2439),.clk(gclk));
	jnot g1798(.din(w_in1101_0[1]),.dout(n2440),.clk(gclk));
	jand g1799(.dina(n2440),.dinb(w_in0101_0[1]),.dout(n2441),.clk(gclk));
	jnot g1800(.din(w_in1100_0[1]),.dout(n2442),.clk(gclk));
	jand g1801(.dina(n2442),.dinb(w_in0100_0[1]),.dout(n2443),.clk(gclk));
	jor g1802(.dina(n2443),.dinb(n2441),.dout(n2444),.clk(gclk));
	jand g1803(.dina(n2444),.dinb(n2439),.dout(n2445),.clk(gclk));
	jnot g1804(.din(w_in1103_0[1]),.dout(n2446),.clk(gclk));
	jand g1805(.dina(n2446),.dinb(w_in0103_0[1]),.dout(n2447),.clk(gclk));
	jnot g1806(.din(w_n2431_0[0]),.dout(n2448),.clk(gclk));
	jnot g1807(.din(w_in1102_0[1]),.dout(n2449),.clk(gclk));
	jand g1808(.dina(n2449),.dinb(w_in0102_0[1]),.dout(n2450),.clk(gclk));
	jand g1809(.dina(n2450),.dinb(n2448),.dout(n2451),.clk(gclk));
	jor g1810(.dina(n2451),.dinb(n2447),.dout(n2452),.clk(gclk));
	jor g1811(.dina(n2452),.dinb(n2445),.dout(n2453),.clk(gclk));
	jor g1812(.dina(w_n2453_0[1]),.dinb(n2438),.dout(n2454),.clk(gclk));
	jnot g1813(.din(w_in0107_0[2]),.dout(n2455),.clk(gclk));
	jand g1814(.dina(w_in1107_0[2]),.dinb(n2455),.dout(n2456),.clk(gclk));
	jnot g1815(.din(w_in0106_0[2]),.dout(n2457),.clk(gclk));
	jand g1816(.dina(w_in1106_0[2]),.dinb(n2457),.dout(n2458),.clk(gclk));
	jor g1817(.dina(n2458),.dinb(n2456),.dout(n2459),.clk(gclk));
	jnot g1818(.din(w_in0105_0[2]),.dout(n2460),.clk(gclk));
	jand g1819(.dina(w_in1105_0[2]),.dinb(n2460),.dout(n2461),.clk(gclk));
	jnot g1820(.din(w_in0104_0[2]),.dout(n2462),.clk(gclk));
	jand g1821(.dina(w_in1104_0[2]),.dinb(n2462),.dout(n2463),.clk(gclk));
	jor g1822(.dina(n2463),.dinb(w_n2461_0[1]),.dout(n2464),.clk(gclk));
	jor g1823(.dina(n2464),.dinb(w_n2459_0[1]),.dout(n2465),.clk(gclk));
	jnot g1824(.din(w_n2465_0[1]),.dout(n2466),.clk(gclk));
	jand g1825(.dina(n2466),.dinb(n2454),.dout(n2467),.clk(gclk));
	jnot g1826(.din(w_in1107_0[1]),.dout(n2468),.clk(gclk));
	jand g1827(.dina(n2468),.dinb(w_in0107_0[1]),.dout(n2469),.clk(gclk));
	jnot g1828(.din(w_n2459_0[0]),.dout(n2470),.clk(gclk));
	jnot g1829(.din(w_n2461_0[0]),.dout(n2471),.clk(gclk));
	jnot g1830(.din(w_in1104_0[1]),.dout(n2472),.clk(gclk));
	jand g1831(.dina(n2472),.dinb(w_in0104_0[1]),.dout(n2473),.clk(gclk));
	jand g1832(.dina(n2473),.dinb(n2471),.dout(n2474),.clk(gclk));
	jnot g1833(.din(w_in1105_0[1]),.dout(n2475),.clk(gclk));
	jand g1834(.dina(n2475),.dinb(w_in0105_0[1]),.dout(n2476),.clk(gclk));
	jnot g1835(.din(w_in1106_0[1]),.dout(n2477),.clk(gclk));
	jand g1836(.dina(n2477),.dinb(w_in0106_0[1]),.dout(n2478),.clk(gclk));
	jor g1837(.dina(n2478),.dinb(n2476),.dout(n2479),.clk(gclk));
	jor g1838(.dina(n2479),.dinb(n2474),.dout(n2480),.clk(gclk));
	jand g1839(.dina(n2480),.dinb(n2470),.dout(n2481),.clk(gclk));
	jor g1840(.dina(n2481),.dinb(n2469),.dout(n2482),.clk(gclk));
	jor g1841(.dina(w_n2482_0[1]),.dinb(n2467),.dout(n2483),.clk(gclk));
	jnot g1842(.din(w_in0108_0[2]),.dout(n2484),.clk(gclk));
	jand g1843(.dina(w_in1108_0[2]),.dinb(n2484),.dout(n2485),.clk(gclk));
	jnot g1844(.din(w_in0109_0[2]),.dout(n2486),.clk(gclk));
	jand g1845(.dina(w_in1109_0[2]),.dinb(n2486),.dout(n2487),.clk(gclk));
	jnot g1846(.din(w_in0111_0[2]),.dout(n2488),.clk(gclk));
	jand g1847(.dina(w_in1111_0[2]),.dinb(n2488),.dout(n2489),.clk(gclk));
	jnot g1848(.din(w_in0110_0[2]),.dout(n2490),.clk(gclk));
	jand g1849(.dina(w_in1110_0[2]),.dinb(n2490),.dout(n2491),.clk(gclk));
	jor g1850(.dina(n2491),.dinb(w_n2489_0[1]),.dout(n2492),.clk(gclk));
	jor g1851(.dina(n2492),.dinb(n2487),.dout(n2493),.clk(gclk));
	jor g1852(.dina(w_n2493_0[1]),.dinb(n2485),.dout(n2494),.clk(gclk));
	jnot g1853(.din(w_n2494_0[1]),.dout(n2495),.clk(gclk));
	jand g1854(.dina(n2495),.dinb(n2483),.dout(n2496),.clk(gclk));
	jnot g1855(.din(w_n2493_0[0]),.dout(n2497),.clk(gclk));
	jnot g1856(.din(w_in1109_0[1]),.dout(n2498),.clk(gclk));
	jand g1857(.dina(n2498),.dinb(w_in0109_0[1]),.dout(n2499),.clk(gclk));
	jnot g1858(.din(w_in1108_0[1]),.dout(n2500),.clk(gclk));
	jand g1859(.dina(n2500),.dinb(w_in0108_0[1]),.dout(n2501),.clk(gclk));
	jor g1860(.dina(n2501),.dinb(n2499),.dout(n2502),.clk(gclk));
	jand g1861(.dina(n2502),.dinb(n2497),.dout(n2503),.clk(gclk));
	jnot g1862(.din(w_in1111_0[1]),.dout(n2504),.clk(gclk));
	jand g1863(.dina(n2504),.dinb(w_in0111_0[1]),.dout(n2505),.clk(gclk));
	jnot g1864(.din(w_n2489_0[0]),.dout(n2506),.clk(gclk));
	jnot g1865(.din(w_in1110_0[1]),.dout(n2507),.clk(gclk));
	jand g1866(.dina(n2507),.dinb(w_in0110_0[1]),.dout(n2508),.clk(gclk));
	jand g1867(.dina(n2508),.dinb(n2506),.dout(n2509),.clk(gclk));
	jor g1868(.dina(n2509),.dinb(n2505),.dout(n2510),.clk(gclk));
	jor g1869(.dina(n2510),.dinb(n2503),.dout(n2511),.clk(gclk));
	jor g1870(.dina(w_n2511_0[1]),.dinb(n2496),.dout(n2512),.clk(gclk));
	jnot g1871(.din(w_in0115_0[2]),.dout(n2513),.clk(gclk));
	jand g1872(.dina(w_in1115_0[2]),.dinb(n2513),.dout(n2514),.clk(gclk));
	jnot g1873(.din(w_in0114_0[2]),.dout(n2515),.clk(gclk));
	jand g1874(.dina(w_in1114_0[2]),.dinb(n2515),.dout(n2516),.clk(gclk));
	jor g1875(.dina(n2516),.dinb(n2514),.dout(n2517),.clk(gclk));
	jnot g1876(.din(w_in0113_0[2]),.dout(n2518),.clk(gclk));
	jand g1877(.dina(w_in1113_0[2]),.dinb(n2518),.dout(n2519),.clk(gclk));
	jnot g1878(.din(w_in0112_0[2]),.dout(n2520),.clk(gclk));
	jand g1879(.dina(w_in1112_0[2]),.dinb(n2520),.dout(n2521),.clk(gclk));
	jor g1880(.dina(n2521),.dinb(w_n2519_0[1]),.dout(n2522),.clk(gclk));
	jor g1881(.dina(n2522),.dinb(w_n2517_0[1]),.dout(n2523),.clk(gclk));
	jnot g1882(.din(w_n2523_0[1]),.dout(n2524),.clk(gclk));
	jand g1883(.dina(n2524),.dinb(n2512),.dout(n2525),.clk(gclk));
	jnot g1884(.din(w_in1115_0[1]),.dout(n2526),.clk(gclk));
	jand g1885(.dina(n2526),.dinb(w_in0115_0[1]),.dout(n2527),.clk(gclk));
	jnot g1886(.din(w_n2517_0[0]),.dout(n2528),.clk(gclk));
	jnot g1887(.din(w_n2519_0[0]),.dout(n2529),.clk(gclk));
	jnot g1888(.din(w_in1112_0[1]),.dout(n2530),.clk(gclk));
	jand g1889(.dina(n2530),.dinb(w_in0112_0[1]),.dout(n2531),.clk(gclk));
	jand g1890(.dina(n2531),.dinb(n2529),.dout(n2532),.clk(gclk));
	jnot g1891(.din(w_in1113_0[1]),.dout(n2533),.clk(gclk));
	jand g1892(.dina(n2533),.dinb(w_in0113_0[1]),.dout(n2534),.clk(gclk));
	jnot g1893(.din(w_in1114_0[1]),.dout(n2535),.clk(gclk));
	jand g1894(.dina(n2535),.dinb(w_in0114_0[1]),.dout(n2536),.clk(gclk));
	jor g1895(.dina(n2536),.dinb(n2534),.dout(n2537),.clk(gclk));
	jor g1896(.dina(n2537),.dinb(n2532),.dout(n2538),.clk(gclk));
	jand g1897(.dina(n2538),.dinb(n2528),.dout(n2539),.clk(gclk));
	jor g1898(.dina(n2539),.dinb(n2527),.dout(n2540),.clk(gclk));
	jor g1899(.dina(w_n2540_0[1]),.dinb(n2525),.dout(n2541),.clk(gclk));
	jnot g1900(.din(w_in0116_0[2]),.dout(n2542),.clk(gclk));
	jand g1901(.dina(w_in1116_0[2]),.dinb(n2542),.dout(n2543),.clk(gclk));
	jnot g1902(.din(w_in0117_0[2]),.dout(n2544),.clk(gclk));
	jand g1903(.dina(w_in1117_0[2]),.dinb(n2544),.dout(n2545),.clk(gclk));
	jnot g1904(.din(w_in0119_0[2]),.dout(n2546),.clk(gclk));
	jand g1905(.dina(w_in1119_0[2]),.dinb(n2546),.dout(n2547),.clk(gclk));
	jnot g1906(.din(w_in0118_0[2]),.dout(n2548),.clk(gclk));
	jand g1907(.dina(w_in1118_0[2]),.dinb(n2548),.dout(n2549),.clk(gclk));
	jor g1908(.dina(n2549),.dinb(w_n2547_0[1]),.dout(n2550),.clk(gclk));
	jor g1909(.dina(n2550),.dinb(n2545),.dout(n2551),.clk(gclk));
	jor g1910(.dina(w_n2551_0[1]),.dinb(n2543),.dout(n2552),.clk(gclk));
	jnot g1911(.din(w_n2552_0[1]),.dout(n2553),.clk(gclk));
	jand g1912(.dina(n2553),.dinb(n2541),.dout(n2554),.clk(gclk));
	jnot g1913(.din(w_n2551_0[0]),.dout(n2555),.clk(gclk));
	jnot g1914(.din(w_in1117_0[1]),.dout(n2556),.clk(gclk));
	jand g1915(.dina(n2556),.dinb(w_in0117_0[1]),.dout(n2557),.clk(gclk));
	jnot g1916(.din(w_in1116_0[1]),.dout(n2558),.clk(gclk));
	jand g1917(.dina(n2558),.dinb(w_in0116_0[1]),.dout(n2559),.clk(gclk));
	jor g1918(.dina(n2559),.dinb(n2557),.dout(n2560),.clk(gclk));
	jand g1919(.dina(n2560),.dinb(n2555),.dout(n2561),.clk(gclk));
	jnot g1920(.din(w_in1119_0[1]),.dout(n2562),.clk(gclk));
	jand g1921(.dina(n2562),.dinb(w_in0119_0[1]),.dout(n2563),.clk(gclk));
	jnot g1922(.din(w_n2547_0[0]),.dout(n2564),.clk(gclk));
	jnot g1923(.din(w_in1118_0[1]),.dout(n2565),.clk(gclk));
	jand g1924(.dina(n2565),.dinb(w_in0118_0[1]),.dout(n2566),.clk(gclk));
	jand g1925(.dina(n2566),.dinb(n2564),.dout(n2567),.clk(gclk));
	jor g1926(.dina(n2567),.dinb(n2563),.dout(n2568),.clk(gclk));
	jor g1927(.dina(n2568),.dinb(n2561),.dout(n2569),.clk(gclk));
	jor g1928(.dina(w_n2569_0[1]),.dinb(n2554),.dout(n2570),.clk(gclk));
	jnot g1929(.din(w_in0123_0[2]),.dout(n2571),.clk(gclk));
	jand g1930(.dina(w_in1123_0[2]),.dinb(n2571),.dout(n2572),.clk(gclk));
	jnot g1931(.din(w_in0122_0[2]),.dout(n2573),.clk(gclk));
	jand g1932(.dina(w_in1122_0[2]),.dinb(n2573),.dout(n2574),.clk(gclk));
	jor g1933(.dina(n2574),.dinb(n2572),.dout(n2575),.clk(gclk));
	jnot g1934(.din(w_in0121_0[2]),.dout(n2576),.clk(gclk));
	jand g1935(.dina(w_in1121_0[2]),.dinb(n2576),.dout(n2577),.clk(gclk));
	jnot g1936(.din(w_in0120_0[2]),.dout(n2578),.clk(gclk));
	jand g1937(.dina(w_in1120_0[2]),.dinb(n2578),.dout(n2579),.clk(gclk));
	jor g1938(.dina(n2579),.dinb(w_n2577_0[1]),.dout(n2580),.clk(gclk));
	jor g1939(.dina(n2580),.dinb(w_n2575_0[1]),.dout(n2581),.clk(gclk));
	jnot g1940(.din(w_n2581_0[1]),.dout(n2582),.clk(gclk));
	jand g1941(.dina(n2582),.dinb(n2570),.dout(n2583),.clk(gclk));
	jnot g1942(.din(w_in1123_0[1]),.dout(n2584),.clk(gclk));
	jand g1943(.dina(n2584),.dinb(w_in0123_0[1]),.dout(n2585),.clk(gclk));
	jnot g1944(.din(w_n2575_0[0]),.dout(n2586),.clk(gclk));
	jnot g1945(.din(w_n2577_0[0]),.dout(n2587),.clk(gclk));
	jnot g1946(.din(w_in1120_0[1]),.dout(n2588),.clk(gclk));
	jand g1947(.dina(n2588),.dinb(w_in0120_0[1]),.dout(n2589),.clk(gclk));
	jand g1948(.dina(n2589),.dinb(n2587),.dout(n2590),.clk(gclk));
	jnot g1949(.din(w_in1121_0[1]),.dout(n2591),.clk(gclk));
	jand g1950(.dina(n2591),.dinb(w_in0121_0[1]),.dout(n2592),.clk(gclk));
	jnot g1951(.din(w_in1122_0[1]),.dout(n2593),.clk(gclk));
	jand g1952(.dina(n2593),.dinb(w_in0122_0[1]),.dout(n2594),.clk(gclk));
	jor g1953(.dina(n2594),.dinb(n2592),.dout(n2595),.clk(gclk));
	jor g1954(.dina(n2595),.dinb(n2590),.dout(n2596),.clk(gclk));
	jand g1955(.dina(n2596),.dinb(n2586),.dout(n2597),.clk(gclk));
	jor g1956(.dina(n2597),.dinb(n2585),.dout(n2598),.clk(gclk));
	jor g1957(.dina(w_n2598_0[1]),.dinb(n2583),.dout(n2599),.clk(gclk));
	jnot g1958(.din(w_in0126_0[2]),.dout(n2600),.clk(gclk));
	jand g1959(.dina(w_in1126_0[2]),.dinb(n2600),.dout(n2601),.clk(gclk));
	jnot g1960(.din(w_in0125_0[2]),.dout(n2602),.clk(gclk));
	jand g1961(.dina(w_in1125_0[2]),.dinb(n2602),.dout(n2603),.clk(gclk));
	jor g1962(.dina(n2603),.dinb(n2601),.dout(n2604),.clk(gclk));
	jnot g1963(.din(w_in1127_0[2]),.dout(n2605),.clk(gclk));
	jand g1964(.dina(n2605),.dinb(w_in0127_0[2]),.dout(n2606),.clk(gclk));
	jnot g1965(.din(w_in0124_0[2]),.dout(n2607),.clk(gclk));
	jand g1966(.dina(w_in1124_0[2]),.dinb(n2607),.dout(n2608),.clk(gclk));
	jor g1967(.dina(n2608),.dinb(w_n2606_0[1]),.dout(n2609),.clk(gclk));
	jor g1968(.dina(n2609),.dinb(w_n2604_0[1]),.dout(n2610),.clk(gclk));
	jnot g1969(.din(w_n2610_0[1]),.dout(n2611),.clk(gclk));
	jand g1970(.dina(n2611),.dinb(n2599),.dout(n2612),.clk(gclk));
	jnot g1971(.din(w_n2606_0[0]),.dout(n2613),.clk(gclk));
	jnot g1972(.din(w_n2604_0[0]),.dout(n2614),.clk(gclk));
	jnot g1973(.din(w_in1124_0[1]),.dout(n2615),.clk(gclk));
	jand g1974(.dina(n2615),.dinb(w_in0124_0[1]),.dout(n2616),.clk(gclk));
	jnot g1975(.din(w_in1125_0[1]),.dout(n2617),.clk(gclk));
	jand g1976(.dina(n2617),.dinb(w_in0125_0[1]),.dout(n2618),.clk(gclk));
	jor g1977(.dina(n2618),.dinb(n2616),.dout(n2619),.clk(gclk));
	jand g1978(.dina(n2619),.dinb(n2614),.dout(n2620),.clk(gclk));
	jnot g1979(.din(w_in1126_0[1]),.dout(n2621),.clk(gclk));
	jand g1980(.dina(n2621),.dinb(w_in0126_0[1]),.dout(n2622),.clk(gclk));
	jor g1981(.dina(n2622),.dinb(n2620),.dout(n2623),.clk(gclk));
	jand g1982(.dina(n2623),.dinb(n2613),.dout(n2624),.clk(gclk));
	jnot g1983(.din(w_in0127_0[1]),.dout(n2625),.clk(gclk));
	jand g1984(.dina(w_in1127_0[1]),.dinb(n2625),.dout(n2626),.clk(gclk));
	jor g1985(.dina(n2626),.dinb(n2624),.dout(n2627),.clk(gclk));
	jor g1986(.dina(w_n2627_0[1]),.dinb(n2612),.dout(n2628),.clk(gclk));
	jand g1987(.dina(w_n2628_64[1]),.dinb(w_in030_0[0]),.dout(n2629),.clk(gclk));
	jnot g1988(.din(w_n1718_0[0]),.dout(n2630),.clk(gclk));
	jnot g1989(.din(w_n1723_0[0]),.dout(n2631),.clk(gclk));
	jnot g1990(.din(w_n1728_0[0]),.dout(n2632),.clk(gclk));
	jnot g1991(.din(w_n1733_0[0]),.dout(n2633),.clk(gclk));
	jnot g1992(.din(w_n1738_0[0]),.dout(n2634),.clk(gclk));
	jnot g1993(.din(w_n1743_0[0]),.dout(n2635),.clk(gclk));
	jnot g1994(.din(w_n1748_0[0]),.dout(n2636),.clk(gclk));
	jnot g1995(.din(w_n1753_0[0]),.dout(n2637),.clk(gclk));
	jnot g1996(.din(w_n1758_0[0]),.dout(n2638),.clk(gclk));
	jnot g1997(.din(w_n1763_0[0]),.dout(n2639),.clk(gclk));
	jnot g1998(.din(w_n1768_0[0]),.dout(n2640),.clk(gclk));
	jnot g1999(.din(w_n1773_0[0]),.dout(n2641),.clk(gclk));
	jnot g2000(.din(w_n1778_0[0]),.dout(n2642),.clk(gclk));
	jnot g2001(.din(w_n1783_0[0]),.dout(n2643),.clk(gclk));
	jnot g2002(.din(w_n1788_0[0]),.dout(n2644),.clk(gclk));
	jnot g2003(.din(w_n1793_0[0]),.dout(n2645),.clk(gclk));
	jnot g2004(.din(w_n1798_0[0]),.dout(n2646),.clk(gclk));
	jnot g2005(.din(w_n1803_0[0]),.dout(n2647),.clk(gclk));
	jnot g2006(.din(w_n1808_0[0]),.dout(n2648),.clk(gclk));
	jnot g2007(.din(w_n1813_0[0]),.dout(n2649),.clk(gclk));
	jnot g2008(.din(w_n1818_0[0]),.dout(n2650),.clk(gclk));
	jnot g2009(.din(w_n1823_0[0]),.dout(n2651),.clk(gclk));
	jnot g2010(.din(w_n1828_0[0]),.dout(n2652),.clk(gclk));
	jnot g2011(.din(w_n1833_0[0]),.dout(n2653),.clk(gclk));
	jnot g2012(.din(w_n1838_0[0]),.dout(n2654),.clk(gclk));
	jnot g2013(.din(w_n1843_0[0]),.dout(n2655),.clk(gclk));
	jnot g2014(.din(w_n1848_0[0]),.dout(n2656),.clk(gclk));
	jnot g2015(.din(w_n1853_0[0]),.dout(n2657),.clk(gclk));
	jnot g2016(.din(w_in01_0[2]),.dout(n2658),.clk(gclk));
	jor g2017(.dina(w_in11_1[0]),.dinb(w_n2658_0[2]),.dout(n2659),.clk(gclk));
	jand g2018(.dina(w_in11_0[2]),.dinb(w_n2658_0[1]),.dout(n2660),.clk(gclk));
	jnot g2019(.din(w_in00_0[1]),.dout(n2661),.clk(gclk));
	jor g2020(.dina(w_in10_0[1]),.dinb(w_n2661_0[1]),.dout(n2662),.clk(gclk));
	jor g2021(.dina(n2662),.dinb(n2660),.dout(n2663),.clk(gclk));
	jand g2022(.dina(n2663),.dinb(n2659),.dout(n2664),.clk(gclk));
	jor g2023(.dina(n2664),.dinb(w_n1855_0[0]),.dout(n2665),.clk(gclk));
	jand g2024(.dina(n2665),.dinb(n2657),.dout(n2666),.clk(gclk));
	jor g2025(.dina(n2666),.dinb(w_n1850_0[0]),.dout(n2667),.clk(gclk));
	jand g2026(.dina(n2667),.dinb(n2656),.dout(n2668),.clk(gclk));
	jor g2027(.dina(n2668),.dinb(w_n1845_0[0]),.dout(n2669),.clk(gclk));
	jand g2028(.dina(n2669),.dinb(n2655),.dout(n2670),.clk(gclk));
	jor g2029(.dina(n2670),.dinb(w_n1840_0[0]),.dout(n2671),.clk(gclk));
	jand g2030(.dina(n2671),.dinb(n2654),.dout(n2672),.clk(gclk));
	jor g2031(.dina(n2672),.dinb(w_n1835_0[0]),.dout(n2673),.clk(gclk));
	jand g2032(.dina(n2673),.dinb(n2653),.dout(n2674),.clk(gclk));
	jor g2033(.dina(n2674),.dinb(w_n1830_0[0]),.dout(n2675),.clk(gclk));
	jand g2034(.dina(n2675),.dinb(n2652),.dout(n2676),.clk(gclk));
	jor g2035(.dina(n2676),.dinb(w_n1825_0[0]),.dout(n2677),.clk(gclk));
	jand g2036(.dina(n2677),.dinb(n2651),.dout(n2678),.clk(gclk));
	jor g2037(.dina(n2678),.dinb(w_n1820_0[0]),.dout(n2679),.clk(gclk));
	jand g2038(.dina(n2679),.dinb(n2650),.dout(n2680),.clk(gclk));
	jor g2039(.dina(n2680),.dinb(w_n1815_0[0]),.dout(n2681),.clk(gclk));
	jand g2040(.dina(n2681),.dinb(n2649),.dout(n2682),.clk(gclk));
	jor g2041(.dina(n2682),.dinb(w_n1810_0[0]),.dout(n2683),.clk(gclk));
	jand g2042(.dina(n2683),.dinb(n2648),.dout(n2684),.clk(gclk));
	jor g2043(.dina(n2684),.dinb(w_n1805_0[0]),.dout(n2685),.clk(gclk));
	jand g2044(.dina(n2685),.dinb(n2647),.dout(n2686),.clk(gclk));
	jor g2045(.dina(n2686),.dinb(w_n1800_0[0]),.dout(n2687),.clk(gclk));
	jand g2046(.dina(n2687),.dinb(n2646),.dout(n2688),.clk(gclk));
	jor g2047(.dina(n2688),.dinb(w_n1795_0[0]),.dout(n2689),.clk(gclk));
	jand g2048(.dina(n2689),.dinb(n2645),.dout(n2690),.clk(gclk));
	jor g2049(.dina(n2690),.dinb(w_n1790_0[0]),.dout(n2691),.clk(gclk));
	jand g2050(.dina(n2691),.dinb(n2644),.dout(n2692),.clk(gclk));
	jor g2051(.dina(n2692),.dinb(w_n1785_0[0]),.dout(n2693),.clk(gclk));
	jand g2052(.dina(n2693),.dinb(n2643),.dout(n2694),.clk(gclk));
	jor g2053(.dina(n2694),.dinb(w_n1780_0[0]),.dout(n2695),.clk(gclk));
	jand g2054(.dina(n2695),.dinb(n2642),.dout(n2696),.clk(gclk));
	jor g2055(.dina(n2696),.dinb(w_n1775_0[0]),.dout(n2697),.clk(gclk));
	jand g2056(.dina(n2697),.dinb(n2641),.dout(n2698),.clk(gclk));
	jor g2057(.dina(n2698),.dinb(w_n1770_0[0]),.dout(n2699),.clk(gclk));
	jand g2058(.dina(n2699),.dinb(n2640),.dout(n2700),.clk(gclk));
	jor g2059(.dina(n2700),.dinb(w_n1765_0[0]),.dout(n2701),.clk(gclk));
	jand g2060(.dina(n2701),.dinb(n2639),.dout(n2702),.clk(gclk));
	jor g2061(.dina(n2702),.dinb(w_n1760_0[0]),.dout(n2703),.clk(gclk));
	jand g2062(.dina(n2703),.dinb(n2638),.dout(n2704),.clk(gclk));
	jor g2063(.dina(n2704),.dinb(w_n1755_0[0]),.dout(n2705),.clk(gclk));
	jand g2064(.dina(n2705),.dinb(n2637),.dout(n2706),.clk(gclk));
	jor g2065(.dina(n2706),.dinb(w_n1750_0[0]),.dout(n2707),.clk(gclk));
	jand g2066(.dina(n2707),.dinb(n2636),.dout(n2708),.clk(gclk));
	jor g2067(.dina(n2708),.dinb(w_n1745_0[0]),.dout(n2709),.clk(gclk));
	jand g2068(.dina(n2709),.dinb(n2635),.dout(n2710),.clk(gclk));
	jor g2069(.dina(n2710),.dinb(w_n1740_0[0]),.dout(n2711),.clk(gclk));
	jand g2070(.dina(n2711),.dinb(n2634),.dout(n2712),.clk(gclk));
	jor g2071(.dina(n2712),.dinb(w_n1735_0[0]),.dout(n2713),.clk(gclk));
	jand g2072(.dina(n2713),.dinb(n2633),.dout(n2714),.clk(gclk));
	jor g2073(.dina(n2714),.dinb(w_n1730_0[0]),.dout(n2715),.clk(gclk));
	jand g2074(.dina(n2715),.dinb(n2632),.dout(n2716),.clk(gclk));
	jor g2075(.dina(n2716),.dinb(w_n1725_0[0]),.dout(n2717),.clk(gclk));
	jand g2076(.dina(n2717),.dinb(n2631),.dout(n2718),.clk(gclk));
	jor g2077(.dina(n2718),.dinb(w_n1720_0[0]),.dout(n2719),.clk(gclk));
	jand g2078(.dina(n2719),.dinb(n2630),.dout(n2720),.clk(gclk));
	jor g2079(.dina(n2720),.dinb(w_n1715_0[0]),.dout(n2721),.clk(gclk));
	jnot g2080(.din(w_n1925_0[0]),.dout(n2722),.clk(gclk));
	jand g2081(.dina(n2722),.dinb(n2721),.dout(n2723),.clk(gclk));
	jor g2082(.dina(w_n1952_0[0]),.dinb(n2723),.dout(n2724),.clk(gclk));
	jnot g2083(.din(w_n1987_0[0]),.dout(n2725),.clk(gclk));
	jand g2084(.dina(n2725),.dinb(n2724),.dout(n2726),.clk(gclk));
	jor g2085(.dina(w_n2011_0[0]),.dinb(n2726),.dout(n2727),.clk(gclk));
	jnot g2086(.din(w_n2046_0[0]),.dout(n2728),.clk(gclk));
	jand g2087(.dina(n2728),.dinb(n2727),.dout(n2729),.clk(gclk));
	jor g2088(.dina(w_n2073_0[0]),.dinb(n2729),.dout(n2730),.clk(gclk));
	jnot g2089(.din(w_n2104_0[0]),.dout(n2731),.clk(gclk));
	jand g2090(.dina(n2731),.dinb(n2730),.dout(n2732),.clk(gclk));
	jor g2091(.dina(w_n2128_0[0]),.dinb(n2732),.dout(n2733),.clk(gclk));
	jnot g2092(.din(w_n2163_0[0]),.dout(n2734),.clk(gclk));
	jand g2093(.dina(n2734),.dinb(n2733),.dout(n2735),.clk(gclk));
	jor g2094(.dina(w_n2175_0[0]),.dinb(n2735),.dout(n2736),.clk(gclk));
	jnot g2095(.din(w_n2192_0[0]),.dout(n2737),.clk(gclk));
	jand g2096(.dina(n2737),.dinb(n2736),.dout(n2738),.clk(gclk));
	jor g2097(.dina(w_n2204_0[0]),.dinb(n2738),.dout(n2739),.clk(gclk));
	jnot g2098(.din(w_n2221_0[0]),.dout(n2740),.clk(gclk));
	jand g2099(.dina(n2740),.dinb(n2739),.dout(n2741),.clk(gclk));
	jor g2100(.dina(w_n2233_0[0]),.dinb(n2741),.dout(n2742),.clk(gclk));
	jnot g2101(.din(w_n2250_0[0]),.dout(n2743),.clk(gclk));
	jand g2102(.dina(n2743),.dinb(n2742),.dout(n2744),.clk(gclk));
	jor g2103(.dina(w_n2262_0[0]),.dinb(n2744),.dout(n2745),.clk(gclk));
	jnot g2104(.din(w_n2279_0[0]),.dout(n2746),.clk(gclk));
	jand g2105(.dina(n2746),.dinb(n2745),.dout(n2747),.clk(gclk));
	jor g2106(.dina(w_n2291_0[0]),.dinb(n2747),.dout(n2748),.clk(gclk));
	jnot g2107(.din(w_n2308_0[0]),.dout(n2749),.clk(gclk));
	jand g2108(.dina(n2749),.dinb(n2748),.dout(n2750),.clk(gclk));
	jor g2109(.dina(w_n2320_0[0]),.dinb(n2750),.dout(n2751),.clk(gclk));
	jnot g2110(.din(w_n2337_0[0]),.dout(n2752),.clk(gclk));
	jand g2111(.dina(n2752),.dinb(n2751),.dout(n2753),.clk(gclk));
	jor g2112(.dina(w_n2349_0[0]),.dinb(n2753),.dout(n2754),.clk(gclk));
	jnot g2113(.din(w_n2366_0[0]),.dout(n2755),.clk(gclk));
	jand g2114(.dina(n2755),.dinb(n2754),.dout(n2756),.clk(gclk));
	jor g2115(.dina(w_n2378_0[0]),.dinb(n2756),.dout(n2757),.clk(gclk));
	jnot g2116(.din(w_n2395_0[0]),.dout(n2758),.clk(gclk));
	jand g2117(.dina(n2758),.dinb(n2757),.dout(n2759),.clk(gclk));
	jor g2118(.dina(w_n2407_0[0]),.dinb(n2759),.dout(n2760),.clk(gclk));
	jnot g2119(.din(w_n2424_0[0]),.dout(n2761),.clk(gclk));
	jand g2120(.dina(n2761),.dinb(n2760),.dout(n2762),.clk(gclk));
	jor g2121(.dina(w_n2436_0[0]),.dinb(n2762),.dout(n2763),.clk(gclk));
	jnot g2122(.din(w_n2453_0[0]),.dout(n2764),.clk(gclk));
	jand g2123(.dina(n2764),.dinb(n2763),.dout(n2765),.clk(gclk));
	jor g2124(.dina(w_n2465_0[0]),.dinb(n2765),.dout(n2766),.clk(gclk));
	jnot g2125(.din(w_n2482_0[0]),.dout(n2767),.clk(gclk));
	jand g2126(.dina(n2767),.dinb(n2766),.dout(n2768),.clk(gclk));
	jor g2127(.dina(w_n2494_0[0]),.dinb(n2768),.dout(n2769),.clk(gclk));
	jnot g2128(.din(w_n2511_0[0]),.dout(n2770),.clk(gclk));
	jand g2129(.dina(n2770),.dinb(n2769),.dout(n2771),.clk(gclk));
	jor g2130(.dina(w_n2523_0[0]),.dinb(n2771),.dout(n2772),.clk(gclk));
	jnot g2131(.din(w_n2540_0[0]),.dout(n2773),.clk(gclk));
	jand g2132(.dina(n2773),.dinb(n2772),.dout(n2774),.clk(gclk));
	jor g2133(.dina(w_n2552_0[0]),.dinb(n2774),.dout(n2775),.clk(gclk));
	jnot g2134(.din(w_n2569_0[0]),.dout(n2776),.clk(gclk));
	jand g2135(.dina(n2776),.dinb(n2775),.dout(n2777),.clk(gclk));
	jor g2136(.dina(w_n2581_0[0]),.dinb(n2777),.dout(n2778),.clk(gclk));
	jnot g2137(.din(w_n2598_0[0]),.dout(n2779),.clk(gclk));
	jand g2138(.dina(n2779),.dinb(n2778),.dout(n2780),.clk(gclk));
	jor g2139(.dina(w_n2610_0[0]),.dinb(n2780),.dout(n2781),.clk(gclk));
	jnot g2140(.din(w_n2627_0[0]),.dout(n2782),.clk(gclk));
	jand g2141(.dina(n2782),.dinb(n2781),.dout(n2783),.clk(gclk));
	jand g2142(.dina(w_n2783_64[2]),.dinb(w_in130_0[0]),.dout(n2784),.clk(gclk));
	jor g2143(.dina(n2784),.dinb(n2629),.dout(n2785),.clk(gclk));
	jnot g2144(.din(w_n2785_0[1]),.dout(n2786),.clk(gclk));
	jand g2145(.dina(w_n1556_63[1]),.dinb(w_in230_0[0]),.dout(n2787),.clk(gclk));
	jand g2146(.dina(w_n1711_64[0]),.dinb(w_in330_0[0]),.dout(n2788),.clk(gclk));
	jor g2147(.dina(n2788),.dinb(n2787),.dout(n2789),.clk(gclk));
	jand g2148(.dina(w_n2789_0[2]),.dinb(w_n2786_0[1]),.dout(n2790),.clk(gclk));
	jand g2149(.dina(w_n2628_64[0]),.dinb(w_in029_0[0]),.dout(n2791),.clk(gclk));
	jand g2150(.dina(w_n2783_64[1]),.dinb(w_in129_0[0]),.dout(n2792),.clk(gclk));
	jor g2151(.dina(n2792),.dinb(n2791),.dout(n2793),.clk(gclk));
	jand g2152(.dina(w_n1556_63[0]),.dinb(w_in229_0[0]),.dout(n2794),.clk(gclk));
	jand g2153(.dina(w_n1711_63[2]),.dinb(w_in329_0[0]),.dout(n2795),.clk(gclk));
	jor g2154(.dina(n2795),.dinb(n2794),.dout(n2796),.clk(gclk));
	jnot g2155(.din(w_n2796_0[1]),.dout(n2797),.clk(gclk));
	jand g2156(.dina(w_n2797_0[1]),.dinb(w_n2793_0[2]),.dout(n2798),.clk(gclk));
	jnot g2157(.din(w_n2798_0[1]),.dout(n2799),.clk(gclk));
	jor g2158(.dina(w_n2797_0[0]),.dinb(w_n2793_0[1]),.dout(n2800),.clk(gclk));
	jnot g2159(.din(w_n2800_0[1]),.dout(n2801),.clk(gclk));
	jand g2160(.dina(w_n2628_63[2]),.dinb(w_in028_0[0]),.dout(n2802),.clk(gclk));
	jand g2161(.dina(w_n2783_64[0]),.dinb(w_in128_0[0]),.dout(n2803),.clk(gclk));
	jor g2162(.dina(n2803),.dinb(n2802),.dout(n2804),.clk(gclk));
	jand g2163(.dina(w_n1556_62[2]),.dinb(w_in228_0[0]),.dout(n2805),.clk(gclk));
	jand g2164(.dina(w_n1711_63[1]),.dinb(w_in328_0[0]),.dout(n2806),.clk(gclk));
	jor g2165(.dina(n2806),.dinb(n2805),.dout(n2807),.clk(gclk));
	jnot g2166(.din(w_n2807_0[1]),.dout(n2808),.clk(gclk));
	jand g2167(.dina(w_n2808_0[1]),.dinb(w_n2804_0[2]),.dout(n2809),.clk(gclk));
	jnot g2168(.din(w_n2809_0[1]),.dout(n2810),.clk(gclk));
	jor g2169(.dina(w_n2808_0[0]),.dinb(w_n2804_0[1]),.dout(n2811),.clk(gclk));
	jnot g2170(.din(w_n2811_0[1]),.dout(n2812),.clk(gclk));
	jand g2171(.dina(w_n2628_63[1]),.dinb(w_in027_0[0]),.dout(n2813),.clk(gclk));
	jand g2172(.dina(w_n2783_63[2]),.dinb(w_in127_0[0]),.dout(n2814),.clk(gclk));
	jor g2173(.dina(n2814),.dinb(n2813),.dout(n2815),.clk(gclk));
	jand g2174(.dina(w_n1556_62[1]),.dinb(w_in227_0[0]),.dout(n2816),.clk(gclk));
	jand g2175(.dina(w_n1711_63[0]),.dinb(w_in327_0[0]),.dout(n2817),.clk(gclk));
	jor g2176(.dina(n2817),.dinb(n2816),.dout(n2818),.clk(gclk));
	jnot g2177(.din(w_n2818_0[1]),.dout(n2819),.clk(gclk));
	jand g2178(.dina(w_n2819_0[1]),.dinb(w_n2815_0[2]),.dout(n2820),.clk(gclk));
	jnot g2179(.din(w_n2820_0[1]),.dout(n2821),.clk(gclk));
	jor g2180(.dina(w_n2819_0[0]),.dinb(w_n2815_0[1]),.dout(n2822),.clk(gclk));
	jnot g2181(.din(w_n2822_0[1]),.dout(n2823),.clk(gclk));
	jand g2182(.dina(w_n2628_63[0]),.dinb(w_in026_0[0]),.dout(n2824),.clk(gclk));
	jand g2183(.dina(w_n2783_63[1]),.dinb(w_in126_0[0]),.dout(n2825),.clk(gclk));
	jor g2184(.dina(n2825),.dinb(n2824),.dout(n2826),.clk(gclk));
	jand g2185(.dina(w_n1556_62[0]),.dinb(w_in226_0[0]),.dout(n2827),.clk(gclk));
	jand g2186(.dina(w_n1711_62[2]),.dinb(w_in326_0[0]),.dout(n2828),.clk(gclk));
	jor g2187(.dina(n2828),.dinb(n2827),.dout(n2829),.clk(gclk));
	jnot g2188(.din(w_n2829_0[1]),.dout(n2830),.clk(gclk));
	jand g2189(.dina(w_n2830_0[1]),.dinb(w_n2826_0[2]),.dout(n2831),.clk(gclk));
	jnot g2190(.din(w_n2831_0[1]),.dout(n2832),.clk(gclk));
	jor g2191(.dina(w_n2830_0[0]),.dinb(w_n2826_0[1]),.dout(n2833),.clk(gclk));
	jnot g2192(.din(w_n2833_0[1]),.dout(n2834),.clk(gclk));
	jand g2193(.dina(w_n2628_62[2]),.dinb(w_in025_0[0]),.dout(n2835),.clk(gclk));
	jand g2194(.dina(w_n2783_63[0]),.dinb(w_in125_0[0]),.dout(n2836),.clk(gclk));
	jor g2195(.dina(n2836),.dinb(n2835),.dout(n2837),.clk(gclk));
	jand g2196(.dina(w_n1556_61[2]),.dinb(w_in225_0[0]),.dout(n2838),.clk(gclk));
	jand g2197(.dina(w_n1711_62[1]),.dinb(w_in325_0[0]),.dout(n2839),.clk(gclk));
	jor g2198(.dina(n2839),.dinb(n2838),.dout(n2840),.clk(gclk));
	jnot g2199(.din(w_n2840_0[1]),.dout(n2841),.clk(gclk));
	jand g2200(.dina(w_n2841_0[1]),.dinb(w_n2837_0[2]),.dout(n2842),.clk(gclk));
	jnot g2201(.din(w_n2842_0[1]),.dout(n2843),.clk(gclk));
	jor g2202(.dina(w_n2841_0[0]),.dinb(w_n2837_0[1]),.dout(n2844),.clk(gclk));
	jnot g2203(.din(w_n2844_0[1]),.dout(n2845),.clk(gclk));
	jand g2204(.dina(w_n2628_62[1]),.dinb(w_in024_0[0]),.dout(n2846),.clk(gclk));
	jand g2205(.dina(w_n2783_62[2]),.dinb(w_in124_0[0]),.dout(n2847),.clk(gclk));
	jor g2206(.dina(n2847),.dinb(n2846),.dout(n2848),.clk(gclk));
	jand g2207(.dina(w_n1556_61[1]),.dinb(w_in224_0[0]),.dout(n2849),.clk(gclk));
	jand g2208(.dina(w_n1711_62[0]),.dinb(w_in324_0[0]),.dout(n2850),.clk(gclk));
	jor g2209(.dina(n2850),.dinb(n2849),.dout(n2851),.clk(gclk));
	jnot g2210(.din(w_n2851_0[1]),.dout(n2852),.clk(gclk));
	jand g2211(.dina(w_n2852_0[1]),.dinb(w_n2848_0[2]),.dout(n2853),.clk(gclk));
	jnot g2212(.din(w_n2853_0[1]),.dout(n2854),.clk(gclk));
	jand g2213(.dina(w_n2628_62[0]),.dinb(w_in022_0[0]),.dout(n2855),.clk(gclk));
	jand g2214(.dina(w_n2783_62[1]),.dinb(w_in122_0[0]),.dout(n2856),.clk(gclk));
	jor g2215(.dina(n2856),.dinb(n2855),.dout(n2857),.clk(gclk));
	jnot g2216(.din(w_n2857_0[1]),.dout(n2858),.clk(gclk));
	jand g2217(.dina(w_n1556_61[0]),.dinb(w_in222_0[0]),.dout(n2859),.clk(gclk));
	jand g2218(.dina(w_n1711_61[2]),.dinb(w_in322_0[0]),.dout(n2860),.clk(gclk));
	jor g2219(.dina(n2860),.dinb(n2859),.dout(n2861),.clk(gclk));
	jand g2220(.dina(w_n2861_0[2]),.dinb(w_n2858_0[1]),.dout(n2862),.clk(gclk));
	jand g2221(.dina(w_n2628_61[2]),.dinb(w_in021_0[0]),.dout(n2863),.clk(gclk));
	jand g2222(.dina(w_n2783_62[0]),.dinb(w_in121_0[0]),.dout(n2864),.clk(gclk));
	jor g2223(.dina(n2864),.dinb(n2863),.dout(n2865),.clk(gclk));
	jand g2224(.dina(w_n1556_60[2]),.dinb(w_in221_0[0]),.dout(n2866),.clk(gclk));
	jand g2225(.dina(w_n1711_61[1]),.dinb(w_in321_0[0]),.dout(n2867),.clk(gclk));
	jor g2226(.dina(n2867),.dinb(n2866),.dout(n2868),.clk(gclk));
	jnot g2227(.din(w_n2868_0[1]),.dout(n2869),.clk(gclk));
	jand g2228(.dina(w_n2869_0[1]),.dinb(w_n2865_0[2]),.dout(n2870),.clk(gclk));
	jnot g2229(.din(w_n2870_0[1]),.dout(n2871),.clk(gclk));
	jor g2230(.dina(w_n2869_0[0]),.dinb(w_n2865_0[1]),.dout(n2872),.clk(gclk));
	jnot g2231(.din(w_n2872_0[1]),.dout(n2873),.clk(gclk));
	jand g2232(.dina(w_n2628_61[1]),.dinb(w_in020_0[0]),.dout(n2874),.clk(gclk));
	jand g2233(.dina(w_n2783_61[2]),.dinb(w_in120_0[0]),.dout(n2875),.clk(gclk));
	jor g2234(.dina(n2875),.dinb(n2874),.dout(n2876),.clk(gclk));
	jand g2235(.dina(w_n1556_60[1]),.dinb(w_in220_0[0]),.dout(n2877),.clk(gclk));
	jand g2236(.dina(w_n1711_61[0]),.dinb(w_in320_0[0]),.dout(n2878),.clk(gclk));
	jor g2237(.dina(n2878),.dinb(n2877),.dout(n2879),.clk(gclk));
	jnot g2238(.din(w_n2879_0[1]),.dout(n2880),.clk(gclk));
	jand g2239(.dina(w_n2880_0[1]),.dinb(w_n2876_0[2]),.dout(n2881),.clk(gclk));
	jnot g2240(.din(w_n2881_0[1]),.dout(n2882),.clk(gclk));
	jor g2241(.dina(w_n2880_0[0]),.dinb(w_n2876_0[1]),.dout(n2883),.clk(gclk));
	jnot g2242(.din(w_n2883_0[1]),.dout(n2884),.clk(gclk));
	jand g2243(.dina(w_n2628_61[0]),.dinb(w_in019_0[0]),.dout(n2885),.clk(gclk));
	jand g2244(.dina(w_n2783_61[1]),.dinb(w_in119_0[0]),.dout(n2886),.clk(gclk));
	jor g2245(.dina(n2886),.dinb(n2885),.dout(n2887),.clk(gclk));
	jand g2246(.dina(w_n1556_60[0]),.dinb(w_in219_0[0]),.dout(n2888),.clk(gclk));
	jand g2247(.dina(w_n1711_60[2]),.dinb(w_in319_0[0]),.dout(n2889),.clk(gclk));
	jor g2248(.dina(n2889),.dinb(n2888),.dout(n2890),.clk(gclk));
	jnot g2249(.din(w_n2890_0[1]),.dout(n2891),.clk(gclk));
	jand g2250(.dina(w_n2891_0[1]),.dinb(w_n2887_0[2]),.dout(n2892),.clk(gclk));
	jnot g2251(.din(w_n2892_0[1]),.dout(n2893),.clk(gclk));
	jand g2252(.dina(w_n1556_59[2]),.dinb(w_in217_0[0]),.dout(n2894),.clk(gclk));
	jand g2253(.dina(w_n1711_60[1]),.dinb(w_in317_0[0]),.dout(n2895),.clk(gclk));
	jor g2254(.dina(n2895),.dinb(n2894),.dout(n2896),.clk(gclk));
	jand g2255(.dina(w_n2628_60[2]),.dinb(w_in017_0[0]),.dout(n2897),.clk(gclk));
	jand g2256(.dina(w_n2783_61[0]),.dinb(w_in117_0[0]),.dout(n2898),.clk(gclk));
	jor g2257(.dina(n2898),.dinb(n2897),.dout(n2899),.clk(gclk));
	jnot g2258(.din(w_n2899_1[1]),.dout(n2900),.clk(gclk));
	jand g2259(.dina(w_n2628_60[1]),.dinb(w_in016_0[0]),.dout(n2901),.clk(gclk));
	jand g2260(.dina(w_n2783_60[2]),.dinb(w_in116_0[0]),.dout(n2902),.clk(gclk));
	jor g2261(.dina(n2902),.dinb(n2901),.dout(n2903),.clk(gclk));
	jnot g2262(.din(w_n2903_0[1]),.dout(n2904),.clk(gclk));
	jand g2263(.dina(w_n1556_59[1]),.dinb(w_in216_0[0]),.dout(n2905),.clk(gclk));
	jand g2264(.dina(w_n1711_60[0]),.dinb(w_in316_0[0]),.dout(n2906),.clk(gclk));
	jor g2265(.dina(n2906),.dinb(n2905),.dout(n2907),.clk(gclk));
	jand g2266(.dina(w_n2907_0[2]),.dinb(w_n2904_0[1]),.dout(n2908),.clk(gclk));
	jor g2267(.dina(w_n2907_0[1]),.dinb(w_n2904_0[0]),.dout(n2909),.clk(gclk));
	jand g2268(.dina(w_n2628_60[0]),.dinb(w_in015_0[0]),.dout(n2910),.clk(gclk));
	jand g2269(.dina(w_n2783_60[1]),.dinb(w_in115_0[0]),.dout(n2911),.clk(gclk));
	jor g2270(.dina(n2911),.dinb(n2910),.dout(n2912),.clk(gclk));
	jnot g2271(.din(w_n2912_0[1]),.dout(n2913),.clk(gclk));
	jand g2272(.dina(w_n1556_59[0]),.dinb(w_in215_0[0]),.dout(n2914),.clk(gclk));
	jand g2273(.dina(w_n1711_59[2]),.dinb(w_in315_0[0]),.dout(n2915),.clk(gclk));
	jor g2274(.dina(n2915),.dinb(n2914),.dout(n2916),.clk(gclk));
	jand g2275(.dina(w_n2916_0[2]),.dinb(w_n2913_0[1]),.dout(n2917),.clk(gclk));
	jand g2276(.dina(w_n2628_59[2]),.dinb(w_in014_0[0]),.dout(n2918),.clk(gclk));
	jand g2277(.dina(w_n2783_60[0]),.dinb(w_in114_0[0]),.dout(n2919),.clk(gclk));
	jor g2278(.dina(n2919),.dinb(n2918),.dout(n2920),.clk(gclk));
	jnot g2279(.din(w_n2920_0[1]),.dout(n2921),.clk(gclk));
	jand g2280(.dina(w_n1556_58[2]),.dinb(w_in214_0[0]),.dout(n2922),.clk(gclk));
	jand g2281(.dina(w_n1711_59[1]),.dinb(w_in314_0[0]),.dout(n2923),.clk(gclk));
	jor g2282(.dina(n2923),.dinb(n2922),.dout(n2924),.clk(gclk));
	jand g2283(.dina(w_n2924_0[2]),.dinb(w_n2921_0[1]),.dout(n2925),.clk(gclk));
	jand g2284(.dina(w_n2628_59[1]),.dinb(w_in013_0[0]),.dout(n2926),.clk(gclk));
	jand g2285(.dina(w_n2783_59[2]),.dinb(w_in113_0[0]),.dout(n2927),.clk(gclk));
	jor g2286(.dina(n2927),.dinb(n2926),.dout(n2928),.clk(gclk));
	jand g2287(.dina(w_n1556_58[1]),.dinb(w_in213_0[0]),.dout(n2929),.clk(gclk));
	jand g2288(.dina(w_n1711_59[0]),.dinb(w_in313_0[0]),.dout(n2930),.clk(gclk));
	jor g2289(.dina(n2930),.dinb(n2929),.dout(n2931),.clk(gclk));
	jnot g2290(.din(w_n2931_0[1]),.dout(n2932),.clk(gclk));
	jand g2291(.dina(w_n2932_0[1]),.dinb(w_n2928_0[2]),.dout(n2933),.clk(gclk));
	jnot g2292(.din(w_n2933_0[1]),.dout(n2934),.clk(gclk));
	jor g2293(.dina(w_n2932_0[0]),.dinb(w_n2928_0[1]),.dout(n2935),.clk(gclk));
	jnot g2294(.din(w_n2935_0[1]),.dout(n2936),.clk(gclk));
	jand g2295(.dina(w_n2628_59[0]),.dinb(w_in012_0[0]),.dout(n2937),.clk(gclk));
	jand g2296(.dina(w_n2783_59[1]),.dinb(w_in112_0[0]),.dout(n2938),.clk(gclk));
	jor g2297(.dina(n2938),.dinb(n2937),.dout(n2939),.clk(gclk));
	jand g2298(.dina(w_n1556_58[0]),.dinb(w_in212_0[0]),.dout(n2940),.clk(gclk));
	jand g2299(.dina(w_n1711_58[2]),.dinb(w_in312_0[0]),.dout(n2941),.clk(gclk));
	jor g2300(.dina(n2941),.dinb(n2940),.dout(n2942),.clk(gclk));
	jnot g2301(.din(w_n2942_0[1]),.dout(n2943),.clk(gclk));
	jand g2302(.dina(w_n2943_0[1]),.dinb(w_n2939_0[2]),.dout(n2944),.clk(gclk));
	jnot g2303(.din(w_n2944_0[1]),.dout(n2945),.clk(gclk));
	jor g2304(.dina(w_n2943_0[0]),.dinb(w_n2939_0[1]),.dout(n2946),.clk(gclk));
	jnot g2305(.din(w_n2946_0[1]),.dout(n2947),.clk(gclk));
	jand g2306(.dina(w_n2628_58[2]),.dinb(w_in011_0[0]),.dout(n2948),.clk(gclk));
	jand g2307(.dina(w_n2783_59[0]),.dinb(w_in111_0[0]),.dout(n2949),.clk(gclk));
	jor g2308(.dina(n2949),.dinb(n2948),.dout(n2950),.clk(gclk));
	jand g2309(.dina(w_n1556_57[2]),.dinb(w_in211_0[0]),.dout(n2951),.clk(gclk));
	jand g2310(.dina(w_n1711_58[1]),.dinb(w_in311_0[0]),.dout(n2952),.clk(gclk));
	jor g2311(.dina(n2952),.dinb(n2951),.dout(n2953),.clk(gclk));
	jnot g2312(.din(w_n2953_0[1]),.dout(n2954),.clk(gclk));
	jand g2313(.dina(w_n2954_0[1]),.dinb(w_n2950_0[2]),.dout(n2955),.clk(gclk));
	jnot g2314(.din(w_n2955_0[1]),.dout(n2956),.clk(gclk));
	jor g2315(.dina(w_n2954_0[0]),.dinb(w_n2950_0[1]),.dout(n2957),.clk(gclk));
	jnot g2316(.din(w_n2957_0[1]),.dout(n2958),.clk(gclk));
	jand g2317(.dina(w_n2628_58[1]),.dinb(w_in010_0[0]),.dout(n2959),.clk(gclk));
	jand g2318(.dina(w_n2783_58[2]),.dinb(w_in110_0[0]),.dout(n2960),.clk(gclk));
	jor g2319(.dina(n2960),.dinb(n2959),.dout(n2961),.clk(gclk));
	jand g2320(.dina(w_n1556_57[1]),.dinb(w_in210_0[0]),.dout(n2962),.clk(gclk));
	jand g2321(.dina(w_n1711_58[0]),.dinb(w_in310_0[0]),.dout(n2963),.clk(gclk));
	jor g2322(.dina(n2963),.dinb(n2962),.dout(n2964),.clk(gclk));
	jnot g2323(.din(w_n2964_0[1]),.dout(n2965),.clk(gclk));
	jand g2324(.dina(w_n2965_0[1]),.dinb(w_n2961_0[2]),.dout(n2966),.clk(gclk));
	jnot g2325(.din(w_n2966_0[1]),.dout(n2967),.clk(gclk));
	jor g2326(.dina(w_n2965_0[0]),.dinb(w_n2961_0[1]),.dout(n2968),.clk(gclk));
	jnot g2327(.din(w_n2968_0[1]),.dout(n2969),.clk(gclk));
	jand g2328(.dina(w_n2628_58[0]),.dinb(w_in09_0[0]),.dout(n2970),.clk(gclk));
	jand g2329(.dina(w_n2783_58[1]),.dinb(w_in19_0[0]),.dout(n2971),.clk(gclk));
	jor g2330(.dina(n2971),.dinb(n2970),.dout(n2972),.clk(gclk));
	jand g2331(.dina(w_n1556_57[0]),.dinb(w_in29_0[0]),.dout(n2973),.clk(gclk));
	jand g2332(.dina(w_n1711_57[2]),.dinb(w_in39_0[0]),.dout(n2974),.clk(gclk));
	jor g2333(.dina(n2974),.dinb(n2973),.dout(n2975),.clk(gclk));
	jnot g2334(.din(w_n2975_0[1]),.dout(n2976),.clk(gclk));
	jand g2335(.dina(w_n2976_0[1]),.dinb(w_n2972_0[2]),.dout(n2977),.clk(gclk));
	jnot g2336(.din(w_n2977_0[1]),.dout(n2978),.clk(gclk));
	jor g2337(.dina(w_n2976_0[0]),.dinb(w_n2972_0[1]),.dout(n2979),.clk(gclk));
	jnot g2338(.din(w_n2979_0[1]),.dout(n2980),.clk(gclk));
	jand g2339(.dina(w_n1556_56[2]),.dinb(w_in28_0[0]),.dout(n2981),.clk(gclk));
	jand g2340(.dina(w_n1711_57[1]),.dinb(w_in38_0[0]),.dout(n2982),.clk(gclk));
	jor g2341(.dina(n2982),.dinb(n2981),.dout(n2983),.clk(gclk));
	jand g2342(.dina(w_n2628_57[2]),.dinb(w_in07_0[0]),.dout(n2984),.clk(gclk));
	jand g2343(.dina(w_n2783_58[0]),.dinb(w_in17_0[0]),.dout(n2985),.clk(gclk));
	jor g2344(.dina(n2985),.dinb(n2984),.dout(n2986),.clk(gclk));
	jand g2345(.dina(w_n1556_56[1]),.dinb(w_in27_0[0]),.dout(n2987),.clk(gclk));
	jand g2346(.dina(w_n1711_57[0]),.dinb(w_in37_0[0]),.dout(n2988),.clk(gclk));
	jor g2347(.dina(n2988),.dinb(n2987),.dout(n2989),.clk(gclk));
	jnot g2348(.din(w_n2989_0[1]),.dout(n2990),.clk(gclk));
	jand g2349(.dina(w_n2990_0[1]),.dinb(w_n2986_0[2]),.dout(n2991),.clk(gclk));
	jnot g2350(.din(w_n2991_0[1]),.dout(n2992),.clk(gclk));
	jor g2351(.dina(w_n2990_0[0]),.dinb(w_n2986_0[1]),.dout(n2993),.clk(gclk));
	jnot g2352(.din(w_n2993_0[1]),.dout(n2994),.clk(gclk));
	jand g2353(.dina(w_n2628_57[1]),.dinb(w_in05_0[0]),.dout(n2995),.clk(gclk));
	jand g2354(.dina(w_n2783_57[2]),.dinb(w_in15_0[0]),.dout(n2996),.clk(gclk));
	jor g2355(.dina(n2996),.dinb(n2995),.dout(n2997),.clk(gclk));
	jnot g2356(.din(w_n2997_0[2]),.dout(n2998),.clk(gclk));
	jand g2357(.dina(w_n2628_57[0]),.dinb(w_in04_0[0]),.dout(n2999),.clk(gclk));
	jand g2358(.dina(w_n2783_57[1]),.dinb(w_in14_0[0]),.dout(n3000),.clk(gclk));
	jor g2359(.dina(n3000),.dinb(n2999),.dout(n3001),.clk(gclk));
	jnot g2360(.din(w_n3001_0[2]),.dout(n3002),.clk(gclk));
	jand g2361(.dina(w_n2628_56[2]),.dinb(w_in03_0[0]),.dout(n3003),.clk(gclk));
	jand g2362(.dina(w_n2783_57[0]),.dinb(w_in13_0[0]),.dout(n3004),.clk(gclk));
	jor g2363(.dina(n3004),.dinb(n3003),.dout(n3005),.clk(gclk));
	jnot g2364(.din(w_n3005_0[1]),.dout(n3006),.clk(gclk));
	jand g2365(.dina(w_n1556_56[0]),.dinb(w_in23_0[0]),.dout(n3007),.clk(gclk));
	jand g2366(.dina(w_n1711_56[2]),.dinb(w_in33_0[0]),.dout(n3008),.clk(gclk));
	jor g2367(.dina(n3008),.dinb(n3007),.dout(n3009),.clk(gclk));
	jand g2368(.dina(w_n3009_0[2]),.dinb(w_n3006_0[1]),.dout(n3010),.clk(gclk));
	jor g2369(.dina(w_n3009_0[1]),.dinb(w_n3006_0[0]),.dout(n3011),.clk(gclk));
	jor g2370(.dina(w_n2783_56[2]),.dinb(w_n1854_0[0]),.dout(n3012),.clk(gclk));
	jor g2371(.dina(w_n2628_56[1]),.dinb(w_n1852_0[0]),.dout(n3013),.clk(gclk));
	jand g2372(.dina(n3013),.dinb(n3012),.dout(n3014),.clk(gclk));
	jand g2373(.dina(w_n1556_55[2]),.dinb(w_in22_0[0]),.dout(n3015),.clk(gclk));
	jand g2374(.dina(w_n1711_56[1]),.dinb(w_in32_0[0]),.dout(n3016),.clk(gclk));
	jor g2375(.dina(n3016),.dinb(n3015),.dout(n3017),.clk(gclk));
	jand g2376(.dina(w_n3017_0[2]),.dinb(w_n3014_0[1]),.dout(n3018),.clk(gclk));
	jand g2377(.dina(w_n1556_55[1]),.dinb(w_in21_0[1]),.dout(n3019),.clk(gclk));
	jand g2378(.dina(w_n1711_56[0]),.dinb(w_in31_0[1]),.dout(n3020),.clk(gclk));
	jor g2379(.dina(n3020),.dinb(n3019),.dout(n3021),.clk(gclk));
	jor g2380(.dina(w_n2783_56[1]),.dinb(w_n2661_0[0]),.dout(n3022),.clk(gclk));
	jor g2381(.dina(w_n2628_56[0]),.dinb(w_n1860_0[0]),.dout(n3023),.clk(gclk));
	jand g2382(.dina(n3023),.dinb(n3022),.dout(n3024),.clk(gclk));
	jor g2383(.dina(n3024),.dinb(w_n1713_0[1]),.dout(n3025),.clk(gclk));
	jor g2384(.dina(w_n2783_56[0]),.dinb(w_n2658_0[0]),.dout(n3026),.clk(gclk));
	jor g2385(.dina(w_n2628_55[2]),.dinb(w_n1857_0[0]),.dout(n3027),.clk(gclk));
	jand g2386(.dina(n3027),.dinb(n3026),.dout(n3028),.clk(gclk));
	jand g2387(.dina(w_n3028_0[1]),.dinb(w_n3025_0[1]),.dout(n3029),.clk(gclk));
	jor g2388(.dina(n3029),.dinb(w_n3021_0[2]),.dout(n3030),.clk(gclk));
	jor g2389(.dina(w_n3017_0[1]),.dinb(w_n3014_0[0]),.dout(n3031),.clk(gclk));
	jor g2390(.dina(w_n3028_0[0]),.dinb(w_n3025_0[0]),.dout(n3032),.clk(gclk));
	jand g2391(.dina(n3032),.dinb(n3031),.dout(n3033),.clk(gclk));
	jand g2392(.dina(n3033),.dinb(n3030),.dout(n3034),.clk(gclk));
	jor g2393(.dina(n3034),.dinb(w_n3018_0[1]),.dout(n3035),.clk(gclk));
	jand g2394(.dina(n3035),.dinb(w_n3011_0[1]),.dout(n3036),.clk(gclk));
	jor g2395(.dina(n3036),.dinb(w_n3010_0[1]),.dout(n3037),.clk(gclk));
	jand g2396(.dina(w_n1556_55[0]),.dinb(w_in24_0[0]),.dout(n3038),.clk(gclk));
	jand g2397(.dina(w_n1711_55[2]),.dinb(w_in34_0[0]),.dout(n3039),.clk(gclk));
	jor g2398(.dina(n3039),.dinb(n3038),.dout(n3040),.clk(gclk));
	jor g2399(.dina(w_n3040_1[1]),.dinb(w_n3037_0[1]),.dout(n3041),.clk(gclk));
	jand g2400(.dina(n3041),.dinb(n3002),.dout(n3042),.clk(gclk));
	jand g2401(.dina(w_n3040_1[0]),.dinb(w_n3037_0[0]),.dout(n3043),.clk(gclk));
	jor g2402(.dina(n3043),.dinb(n3042),.dout(n3044),.clk(gclk));
	jand g2403(.dina(w_n1556_54[2]),.dinb(w_in25_0[0]),.dout(n3045),.clk(gclk));
	jand g2404(.dina(w_n1711_55[1]),.dinb(w_in35_0[0]),.dout(n3046),.clk(gclk));
	jor g2405(.dina(n3046),.dinb(n3045),.dout(n3047),.clk(gclk));
	jor g2406(.dina(w_n3047_1[1]),.dinb(w_n3044_0[1]),.dout(n3048),.clk(gclk));
	jand g2407(.dina(n3048),.dinb(n2998),.dout(n3049),.clk(gclk));
	jand g2408(.dina(w_n3047_1[0]),.dinb(w_n3044_0[0]),.dout(n3050),.clk(gclk));
	jand g2409(.dina(w_n2628_55[1]),.dinb(w_in06_0[0]),.dout(n3051),.clk(gclk));
	jand g2410(.dina(w_n2783_55[2]),.dinb(w_in16_0[0]),.dout(n3052),.clk(gclk));
	jor g2411(.dina(n3052),.dinb(n3051),.dout(n3053),.clk(gclk));
	jnot g2412(.din(w_n3053_0[1]),.dout(n3054),.clk(gclk));
	jand g2413(.dina(w_n1556_54[1]),.dinb(w_in26_0[0]),.dout(n3055),.clk(gclk));
	jand g2414(.dina(w_n1711_55[0]),.dinb(w_in36_0[0]),.dout(n3056),.clk(gclk));
	jor g2415(.dina(n3056),.dinb(n3055),.dout(n3057),.clk(gclk));
	jand g2416(.dina(w_n3057_0[2]),.dinb(w_n3054_0[1]),.dout(n3058),.clk(gclk));
	jor g2417(.dina(w_n3058_0[1]),.dinb(n3050),.dout(n3059),.clk(gclk));
	jor g2418(.dina(n3059),.dinb(n3049),.dout(n3060),.clk(gclk));
	jor g2419(.dina(w_n3057_0[1]),.dinb(w_n3054_0[0]),.dout(n3061),.clk(gclk));
	jand g2420(.dina(w_n3061_0[1]),.dinb(n3060),.dout(n3062),.clk(gclk));
	jor g2421(.dina(n3062),.dinb(n2994),.dout(n3063),.clk(gclk));
	jand g2422(.dina(n3063),.dinb(n2992),.dout(n3064),.clk(gclk));
	jand g2423(.dina(w_n2628_55[0]),.dinb(w_in08_0[0]),.dout(n3065),.clk(gclk));
	jand g2424(.dina(w_n2783_55[1]),.dinb(w_in18_0[0]),.dout(n3066),.clk(gclk));
	jor g2425(.dina(n3066),.dinb(n3065),.dout(n3067),.clk(gclk));
	jnot g2426(.din(w_n3067_1[1]),.dout(n3068),.clk(gclk));
	jand g2427(.dina(w_n3068_0[1]),.dinb(w_n3064_0[1]),.dout(n3069),.clk(gclk));
	jor g2428(.dina(n3069),.dinb(w_n2983_0[2]),.dout(n3070),.clk(gclk));
	jor g2429(.dina(w_n3068_0[0]),.dinb(w_n3064_0[0]),.dout(n3071),.clk(gclk));
	jand g2430(.dina(n3071),.dinb(n3070),.dout(n3072),.clk(gclk));
	jor g2431(.dina(n3072),.dinb(n2980),.dout(n3073),.clk(gclk));
	jand g2432(.dina(n3073),.dinb(n2978),.dout(n3074),.clk(gclk));
	jor g2433(.dina(n3074),.dinb(n2969),.dout(n3075),.clk(gclk));
	jand g2434(.dina(n3075),.dinb(n2967),.dout(n3076),.clk(gclk));
	jor g2435(.dina(n3076),.dinb(n2958),.dout(n3077),.clk(gclk));
	jand g2436(.dina(n3077),.dinb(n2956),.dout(n3078),.clk(gclk));
	jor g2437(.dina(n3078),.dinb(n2947),.dout(n3079),.clk(gclk));
	jand g2438(.dina(n3079),.dinb(n2945),.dout(n3080),.clk(gclk));
	jor g2439(.dina(n3080),.dinb(n2936),.dout(n3081),.clk(gclk));
	jand g2440(.dina(n3081),.dinb(n2934),.dout(n3082),.clk(gclk));
	jor g2441(.dina(n3082),.dinb(w_n2925_0[1]),.dout(n3083),.clk(gclk));
	jor g2442(.dina(w_n2924_0[1]),.dinb(w_n2921_0[0]),.dout(n3084),.clk(gclk));
	jor g2443(.dina(w_n2916_0[1]),.dinb(w_n2913_0[0]),.dout(n3085),.clk(gclk));
	jand g2444(.dina(n3085),.dinb(n3084),.dout(n3086),.clk(gclk));
	jand g2445(.dina(w_n3086_0[1]),.dinb(n3083),.dout(n3087),.clk(gclk));
	jor g2446(.dina(n3087),.dinb(w_n2917_0[1]),.dout(n3088),.clk(gclk));
	jand g2447(.dina(n3088),.dinb(w_n2909_0[1]),.dout(n3089),.clk(gclk));
	jor g2448(.dina(n3089),.dinb(w_n2908_0[1]),.dout(n3090),.clk(gclk));
	jand g2449(.dina(w_n3090_0[1]),.dinb(w_n2900_0[1]),.dout(n3091),.clk(gclk));
	jor g2450(.dina(n3091),.dinb(w_n2896_0[2]),.dout(n3092),.clk(gclk));
	jand g2451(.dina(w_n2628_54[2]),.dinb(w_in018_0[0]),.dout(n3093),.clk(gclk));
	jand g2452(.dina(w_n2783_55[0]),.dinb(w_in118_0[0]),.dout(n3094),.clk(gclk));
	jor g2453(.dina(n3094),.dinb(n3093),.dout(n3095),.clk(gclk));
	jand g2454(.dina(w_n1556_54[0]),.dinb(w_in218_0[0]),.dout(n3096),.clk(gclk));
	jand g2455(.dina(w_n1711_54[2]),.dinb(w_in318_0[0]),.dout(n3097),.clk(gclk));
	jor g2456(.dina(n3097),.dinb(n3096),.dout(n3098),.clk(gclk));
	jnot g2457(.din(w_n3098_0[1]),.dout(n3099),.clk(gclk));
	jand g2458(.dina(w_n3099_0[1]),.dinb(w_n3095_0[2]),.dout(n3100),.clk(gclk));
	jnot g2459(.din(w_n3100_0[1]),.dout(n3101),.clk(gclk));
	jor g2460(.dina(w_n3090_0[0]),.dinb(w_n2900_0[0]),.dout(n3102),.clk(gclk));
	jand g2461(.dina(n3102),.dinb(n3101),.dout(n3103),.clk(gclk));
	jand g2462(.dina(n3103),.dinb(n3092),.dout(n3104),.clk(gclk));
	jor g2463(.dina(w_n2891_0[0]),.dinb(w_n2887_0[1]),.dout(n3105),.clk(gclk));
	jor g2464(.dina(w_n3099_0[0]),.dinb(w_n3095_0[1]),.dout(n3106),.clk(gclk));
	jand g2465(.dina(n3106),.dinb(n3105),.dout(n3107),.clk(gclk));
	jnot g2466(.din(w_n3107_0[1]),.dout(n3108),.clk(gclk));
	jor g2467(.dina(n3108),.dinb(n3104),.dout(n3109),.clk(gclk));
	jand g2468(.dina(n3109),.dinb(n2893),.dout(n3110),.clk(gclk));
	jor g2469(.dina(n3110),.dinb(n2884),.dout(n3111),.clk(gclk));
	jand g2470(.dina(n3111),.dinb(n2882),.dout(n3112),.clk(gclk));
	jor g2471(.dina(n3112),.dinb(n2873),.dout(n3113),.clk(gclk));
	jand g2472(.dina(n3113),.dinb(n2871),.dout(n3114),.clk(gclk));
	jor g2473(.dina(n3114),.dinb(w_n2862_0[1]),.dout(n3115),.clk(gclk));
	jor g2474(.dina(w_n2861_0[1]),.dinb(w_n2858_0[0]),.dout(n3116),.clk(gclk));
	jand g2475(.dina(w_n2628_54[1]),.dinb(w_in023_0[0]),.dout(n3117),.clk(gclk));
	jand g2476(.dina(w_n2783_54[2]),.dinb(w_in123_0[0]),.dout(n3118),.clk(gclk));
	jor g2477(.dina(n3118),.dinb(n3117),.dout(n3119),.clk(gclk));
	jand g2478(.dina(w_n1556_53[2]),.dinb(w_in223_0[0]),.dout(n3120),.clk(gclk));
	jand g2479(.dina(w_n1711_54[1]),.dinb(w_in323_0[0]),.dout(n3121),.clk(gclk));
	jor g2480(.dina(n3121),.dinb(n3120),.dout(n3122),.clk(gclk));
	jnot g2481(.din(w_n3122_0[1]),.dout(n3123),.clk(gclk));
	jand g2482(.dina(w_n3123_0[1]),.dinb(w_n3119_0[2]),.dout(n3124),.clk(gclk));
	jnot g2483(.din(n3124),.dout(n3125),.clk(gclk));
	jand g2484(.dina(n3125),.dinb(n3116),.dout(n3126),.clk(gclk));
	jand g2485(.dina(w_n3126_0[1]),.dinb(n3115),.dout(n3127),.clk(gclk));
	jor g2486(.dina(w_n3123_0[0]),.dinb(w_n3119_0[1]),.dout(n3128),.clk(gclk));
	jor g2487(.dina(w_n2852_0[0]),.dinb(w_n2848_0[1]),.dout(n3129),.clk(gclk));
	jand g2488(.dina(n3129),.dinb(n3128),.dout(n3130),.clk(gclk));
	jnot g2489(.din(w_n3130_0[1]),.dout(n3131),.clk(gclk));
	jor g2490(.dina(n3131),.dinb(n3127),.dout(n3132),.clk(gclk));
	jand g2491(.dina(n3132),.dinb(n2854),.dout(n3133),.clk(gclk));
	jor g2492(.dina(n3133),.dinb(n2845),.dout(n3134),.clk(gclk));
	jand g2493(.dina(n3134),.dinb(n2843),.dout(n3135),.clk(gclk));
	jor g2494(.dina(n3135),.dinb(n2834),.dout(n3136),.clk(gclk));
	jand g2495(.dina(n3136),.dinb(n2832),.dout(n3137),.clk(gclk));
	jor g2496(.dina(n3137),.dinb(n2823),.dout(n3138),.clk(gclk));
	jand g2497(.dina(n3138),.dinb(n2821),.dout(n3139),.clk(gclk));
	jor g2498(.dina(n3139),.dinb(n2812),.dout(n3140),.clk(gclk));
	jand g2499(.dina(n3140),.dinb(n2810),.dout(n3141),.clk(gclk));
	jor g2500(.dina(n3141),.dinb(n2801),.dout(n3142),.clk(gclk));
	jand g2501(.dina(n3142),.dinb(n2799),.dout(n3143),.clk(gclk));
	jor g2502(.dina(n3143),.dinb(w_n2790_0[1]),.dout(n3144),.clk(gclk));
	jor g2503(.dina(w_n2789_0[1]),.dinb(w_n2786_0[0]),.dout(n3145),.clk(gclk));
	jand g2504(.dina(w_n2628_54[0]),.dinb(w_in031_0[0]),.dout(n3146),.clk(gclk));
	jand g2505(.dina(w_n2783_54[1]),.dinb(w_in131_0[0]),.dout(n3147),.clk(gclk));
	jor g2506(.dina(n3147),.dinb(n3146),.dout(n3148),.clk(gclk));
	jand g2507(.dina(w_n1556_53[1]),.dinb(w_in231_0[0]),.dout(n3149),.clk(gclk));
	jand g2508(.dina(w_n1711_54[0]),.dinb(w_in331_0[0]),.dout(n3150),.clk(gclk));
	jor g2509(.dina(n3150),.dinb(n3149),.dout(n3151),.clk(gclk));
	jnot g2510(.din(w_n3151_0[1]),.dout(n3152),.clk(gclk));
	jand g2511(.dina(w_n3152_0[1]),.dinb(w_n3148_0[2]),.dout(n3153),.clk(gclk));
	jnot g2512(.din(n3153),.dout(n3154),.clk(gclk));
	jand g2513(.dina(n3154),.dinb(n3145),.dout(n3155),.clk(gclk));
	jand g2514(.dina(w_n3155_0[1]),.dinb(n3144),.dout(n3156),.clk(gclk));
	jand g2515(.dina(w_n2628_53[2]),.dinb(w_in037_0[0]),.dout(n3157),.clk(gclk));
	jand g2516(.dina(w_n2783_54[0]),.dinb(w_in137_0[0]),.dout(n3158),.clk(gclk));
	jor g2517(.dina(n3158),.dinb(n3157),.dout(n3159),.clk(gclk));
	jnot g2518(.din(w_n3159_0[1]),.dout(n3160),.clk(gclk));
	jand g2519(.dina(w_n1556_53[0]),.dinb(w_in237_0[0]),.dout(n3161),.clk(gclk));
	jand g2520(.dina(w_n1711_53[2]),.dinb(w_in337_0[0]),.dout(n3162),.clk(gclk));
	jor g2521(.dina(n3162),.dinb(n3161),.dout(n3163),.clk(gclk));
	jand g2522(.dina(w_n3163_0[2]),.dinb(w_n3160_0[1]),.dout(n3164),.clk(gclk));
	jand g2523(.dina(w_n2628_53[1]),.dinb(w_in039_0[0]),.dout(n3165),.clk(gclk));
	jand g2524(.dina(w_n2783_53[2]),.dinb(w_in139_0[0]),.dout(n3166),.clk(gclk));
	jor g2525(.dina(n3166),.dinb(n3165),.dout(n3167),.clk(gclk));
	jnot g2526(.din(w_n3167_0[1]),.dout(n3168),.clk(gclk));
	jand g2527(.dina(w_n1556_52[2]),.dinb(w_in239_0[0]),.dout(n3169),.clk(gclk));
	jand g2528(.dina(w_n1711_53[1]),.dinb(w_in339_0[0]),.dout(n3170),.clk(gclk));
	jor g2529(.dina(n3170),.dinb(n3169),.dout(n3171),.clk(gclk));
	jand g2530(.dina(w_n3171_0[2]),.dinb(w_n3168_0[1]),.dout(n3172),.clk(gclk));
	jand g2531(.dina(w_n1556_52[1]),.dinb(w_in238_0[0]),.dout(n3173),.clk(gclk));
	jand g2532(.dina(w_n1711_53[0]),.dinb(w_in338_0[0]),.dout(n3174),.clk(gclk));
	jor g2533(.dina(n3174),.dinb(n3173),.dout(n3175),.clk(gclk));
	jand g2534(.dina(w_n2628_53[0]),.dinb(w_in038_0[0]),.dout(n3176),.clk(gclk));
	jand g2535(.dina(w_n2783_53[1]),.dinb(w_in138_0[0]),.dout(n3177),.clk(gclk));
	jor g2536(.dina(n3177),.dinb(n3176),.dout(n3178),.clk(gclk));
	jnot g2537(.din(w_n3178_0[1]),.dout(n3179),.clk(gclk));
	jand g2538(.dina(w_n3179_0[1]),.dinb(w_n3175_0[2]),.dout(n3180),.clk(gclk));
	jor g2539(.dina(n3180),.dinb(w_n3172_0[1]),.dout(n3181),.clk(gclk));
	jor g2540(.dina(n3181),.dinb(n3164),.dout(n3182),.clk(gclk));
	jnot g2541(.din(w_n3182_0[1]),.dout(n3183),.clk(gclk));
	jand g2542(.dina(w_n2628_52[2]),.dinb(w_in035_0[0]),.dout(n3184),.clk(gclk));
	jand g2543(.dina(w_n2783_53[0]),.dinb(w_in135_0[0]),.dout(n3185),.clk(gclk));
	jor g2544(.dina(n3185),.dinb(n3184),.dout(n3186),.clk(gclk));
	jnot g2545(.din(w_n3186_0[1]),.dout(n3187),.clk(gclk));
	jand g2546(.dina(w_n1556_52[0]),.dinb(w_in235_0[0]),.dout(n3188),.clk(gclk));
	jand g2547(.dina(w_n1711_52[2]),.dinb(w_in335_0[0]),.dout(n3189),.clk(gclk));
	jor g2548(.dina(n3189),.dinb(n3188),.dout(n3190),.clk(gclk));
	jand g2549(.dina(w_n3190_0[2]),.dinb(w_n3187_0[1]),.dout(n3191),.clk(gclk));
	jand g2550(.dina(w_n2628_52[1]),.dinb(w_in033_0[0]),.dout(n3192),.clk(gclk));
	jand g2551(.dina(w_n2783_52[2]),.dinb(w_in133_0[0]),.dout(n3193),.clk(gclk));
	jor g2552(.dina(n3193),.dinb(n3192),.dout(n3194),.clk(gclk));
	jnot g2553(.din(w_n3194_0[1]),.dout(n3195),.clk(gclk));
	jand g2554(.dina(w_n1556_51[2]),.dinb(w_in233_0[0]),.dout(n3196),.clk(gclk));
	jand g2555(.dina(w_n1711_52[1]),.dinb(w_in333_0[0]),.dout(n3197),.clk(gclk));
	jor g2556(.dina(n3197),.dinb(n3196),.dout(n3198),.clk(gclk));
	jand g2557(.dina(w_n3198_0[2]),.dinb(w_n3195_0[1]),.dout(n3199),.clk(gclk));
	jand g2558(.dina(w_n1556_51[1]),.dinb(w_in234_0[0]),.dout(n3200),.clk(gclk));
	jand g2559(.dina(w_n1711_52[0]),.dinb(w_in334_0[0]),.dout(n3201),.clk(gclk));
	jor g2560(.dina(n3201),.dinb(n3200),.dout(n3202),.clk(gclk));
	jand g2561(.dina(w_n2628_52[0]),.dinb(w_in034_0[0]),.dout(n3203),.clk(gclk));
	jand g2562(.dina(w_n2783_52[1]),.dinb(w_in134_0[0]),.dout(n3204),.clk(gclk));
	jor g2563(.dina(n3204),.dinb(n3203),.dout(n3205),.clk(gclk));
	jnot g2564(.din(w_n3205_0[1]),.dout(n3206),.clk(gclk));
	jand g2565(.dina(w_n3206_0[1]),.dinb(w_n3202_0[2]),.dout(n3207),.clk(gclk));
	jor g2566(.dina(n3207),.dinb(n3199),.dout(n3208),.clk(gclk));
	jor g2567(.dina(n3208),.dinb(w_n3191_0[1]),.dout(n3209),.clk(gclk));
	jnot g2568(.din(w_n3209_0[1]),.dout(n3210),.clk(gclk));
	jand g2569(.dina(w_n1556_51[0]),.dinb(w_in232_0[0]),.dout(n3211),.clk(gclk));
	jand g2570(.dina(w_n1711_51[2]),.dinb(w_in332_0[0]),.dout(n3212),.clk(gclk));
	jor g2571(.dina(n3212),.dinb(n3211),.dout(n3213),.clk(gclk));
	jand g2572(.dina(w_n2628_51[2]),.dinb(w_in032_0[0]),.dout(n3214),.clk(gclk));
	jand g2573(.dina(w_n2783_52[0]),.dinb(w_in132_0[0]),.dout(n3215),.clk(gclk));
	jor g2574(.dina(n3215),.dinb(n3214),.dout(n3216),.clk(gclk));
	jnot g2575(.din(w_n3216_0[1]),.dout(n3217),.clk(gclk));
	jand g2576(.dina(w_n3217_0[1]),.dinb(w_n3213_0[2]),.dout(n3218),.clk(gclk));
	jnot g2577(.din(n3218),.dout(n3219),.clk(gclk));
	jand g2578(.dina(w_n2628_51[1]),.dinb(w_in036_0[0]),.dout(n3220),.clk(gclk));
	jand g2579(.dina(w_n2783_51[2]),.dinb(w_in136_0[0]),.dout(n3221),.clk(gclk));
	jor g2580(.dina(n3221),.dinb(n3220),.dout(n3222),.clk(gclk));
	jnot g2581(.din(w_n3222_0[1]),.dout(n3223),.clk(gclk));
	jand g2582(.dina(w_n1556_50[2]),.dinb(w_in236_0[0]),.dout(n3224),.clk(gclk));
	jand g2583(.dina(w_n1711_51[1]),.dinb(w_in336_0[0]),.dout(n3225),.clk(gclk));
	jor g2584(.dina(n3225),.dinb(n3224),.dout(n3226),.clk(gclk));
	jand g2585(.dina(w_n3226_0[2]),.dinb(w_n3223_0[1]),.dout(n3227),.clk(gclk));
	jnot g2586(.din(w_n3227_0[1]),.dout(n3228),.clk(gclk));
	jor g2587(.dina(w_n3152_0[0]),.dinb(w_n3148_0[1]),.dout(n3229),.clk(gclk));
	jand g2588(.dina(n3229),.dinb(n3228),.dout(n3230),.clk(gclk));
	jand g2589(.dina(n3230),.dinb(n3219),.dout(n3231),.clk(gclk));
	jand g2590(.dina(n3231),.dinb(n3210),.dout(n3232),.clk(gclk));
	jand g2591(.dina(n3232),.dinb(n3183),.dout(n3233),.clk(gclk));
	jnot g2592(.din(w_n3233_0[1]),.dout(n3234),.clk(gclk));
	jor g2593(.dina(n3234),.dinb(n3156),.dout(n3235),.clk(gclk));
	jor g2594(.dina(w_n3217_0[0]),.dinb(w_n3213_0[1]),.dout(n3236),.clk(gclk));
	jor g2595(.dina(w_n3198_0[1]),.dinb(w_n3195_0[0]),.dout(n3237),.clk(gclk));
	jand g2596(.dina(n3237),.dinb(n3236),.dout(n3238),.clk(gclk));
	jor g2597(.dina(n3238),.dinb(w_n3209_0[0]),.dout(n3239),.clk(gclk));
	jor g2598(.dina(w_n3206_0[0]),.dinb(w_n3202_0[1]),.dout(n3240),.clk(gclk));
	jor g2599(.dina(n3240),.dinb(w_n3191_0[0]),.dout(n3241),.clk(gclk));
	jor g2600(.dina(w_n3190_0[1]),.dinb(w_n3187_0[0]),.dout(n3242),.clk(gclk));
	jand g2601(.dina(n3242),.dinb(n3241),.dout(n3243),.clk(gclk));
	jand g2602(.dina(n3243),.dinb(n3239),.dout(n3244),.clk(gclk));
	jor g2603(.dina(n3244),.dinb(w_n3227_0[0]),.dout(n3245),.clk(gclk));
	jor g2604(.dina(w_n3226_0[1]),.dinb(w_n3223_0[0]),.dout(n3246),.clk(gclk));
	jor g2605(.dina(w_n3163_0[1]),.dinb(w_n3160_0[0]),.dout(n3247),.clk(gclk));
	jand g2606(.dina(n3247),.dinb(n3246),.dout(n3248),.clk(gclk));
	jand g2607(.dina(n3248),.dinb(n3245),.dout(n3249),.clk(gclk));
	jor g2608(.dina(n3249),.dinb(w_n3182_0[0]),.dout(n3250),.clk(gclk));
	jor g2609(.dina(w_n3179_0[0]),.dinb(w_n3175_0[1]),.dout(n3251),.clk(gclk));
	jor g2610(.dina(n3251),.dinb(w_n3172_0[0]),.dout(n3252),.clk(gclk));
	jor g2611(.dina(w_n3171_0[1]),.dinb(w_n3168_0[0]),.dout(n3253),.clk(gclk));
	jand g2612(.dina(n3253),.dinb(n3252),.dout(n3254),.clk(gclk));
	jand g2613(.dina(n3254),.dinb(n3250),.dout(n3255),.clk(gclk));
	jand g2614(.dina(w_n3255_0[1]),.dinb(n3235),.dout(n3256),.clk(gclk));
	jand g2615(.dina(w_n2628_51[0]),.dinb(w_in045_0[0]),.dout(n3257),.clk(gclk));
	jand g2616(.dina(w_n2783_51[1]),.dinb(w_in145_0[0]),.dout(n3258),.clk(gclk));
	jor g2617(.dina(n3258),.dinb(n3257),.dout(n3259),.clk(gclk));
	jnot g2618(.din(w_n3259_0[1]),.dout(n3260),.clk(gclk));
	jand g2619(.dina(w_n1556_50[1]),.dinb(w_in245_0[0]),.dout(n3261),.clk(gclk));
	jand g2620(.dina(w_n1711_51[0]),.dinb(w_in345_0[0]),.dout(n3262),.clk(gclk));
	jor g2621(.dina(n3262),.dinb(n3261),.dout(n3263),.clk(gclk));
	jand g2622(.dina(w_n3263_0[2]),.dinb(w_n3260_0[1]),.dout(n3264),.clk(gclk));
	jand g2623(.dina(w_n2628_50[2]),.dinb(w_in047_0[0]),.dout(n3265),.clk(gclk));
	jand g2624(.dina(w_n2783_51[0]),.dinb(w_in147_0[0]),.dout(n3266),.clk(gclk));
	jor g2625(.dina(n3266),.dinb(n3265),.dout(n3267),.clk(gclk));
	jnot g2626(.din(w_n3267_0[1]),.dout(n3268),.clk(gclk));
	jand g2627(.dina(w_n1556_50[0]),.dinb(w_in247_0[0]),.dout(n3269),.clk(gclk));
	jand g2628(.dina(w_n1711_50[2]),.dinb(w_in347_0[0]),.dout(n3270),.clk(gclk));
	jor g2629(.dina(n3270),.dinb(n3269),.dout(n3271),.clk(gclk));
	jand g2630(.dina(w_n3271_0[2]),.dinb(w_n3268_0[1]),.dout(n3272),.clk(gclk));
	jand g2631(.dina(w_n1556_49[2]),.dinb(w_in246_0[0]),.dout(n3273),.clk(gclk));
	jand g2632(.dina(w_n1711_50[1]),.dinb(w_in346_0[0]),.dout(n3274),.clk(gclk));
	jor g2633(.dina(n3274),.dinb(n3273),.dout(n3275),.clk(gclk));
	jand g2634(.dina(w_n2628_50[1]),.dinb(w_in046_0[0]),.dout(n3276),.clk(gclk));
	jand g2635(.dina(w_n2783_50[2]),.dinb(w_in146_0[0]),.dout(n3277),.clk(gclk));
	jor g2636(.dina(n3277),.dinb(n3276),.dout(n3278),.clk(gclk));
	jnot g2637(.din(w_n3278_0[1]),.dout(n3279),.clk(gclk));
	jand g2638(.dina(w_n3279_0[1]),.dinb(w_n3275_0[2]),.dout(n3280),.clk(gclk));
	jor g2639(.dina(n3280),.dinb(w_n3272_0[1]),.dout(n3281),.clk(gclk));
	jor g2640(.dina(n3281),.dinb(n3264),.dout(n3282),.clk(gclk));
	jand g2641(.dina(w_n2628_50[0]),.dinb(w_in043_0[0]),.dout(n3283),.clk(gclk));
	jand g2642(.dina(w_n2783_50[1]),.dinb(w_in143_0[0]),.dout(n3284),.clk(gclk));
	jor g2643(.dina(n3284),.dinb(n3283),.dout(n3285),.clk(gclk));
	jnot g2644(.din(w_n3285_0[1]),.dout(n3286),.clk(gclk));
	jand g2645(.dina(w_n1556_49[1]),.dinb(w_in243_0[0]),.dout(n3287),.clk(gclk));
	jand g2646(.dina(w_n1711_50[0]),.dinb(w_in343_0[0]),.dout(n3288),.clk(gclk));
	jor g2647(.dina(n3288),.dinb(n3287),.dout(n3289),.clk(gclk));
	jand g2648(.dina(w_n3289_0[2]),.dinb(w_n3286_0[1]),.dout(n3290),.clk(gclk));
	jand g2649(.dina(w_n2628_49[2]),.dinb(w_in042_0[0]),.dout(n3291),.clk(gclk));
	jand g2650(.dina(w_n2783_50[0]),.dinb(w_in142_0[0]),.dout(n3292),.clk(gclk));
	jor g2651(.dina(n3292),.dinb(n3291),.dout(n3293),.clk(gclk));
	jnot g2652(.din(w_n3293_0[1]),.dout(n3294),.clk(gclk));
	jand g2653(.dina(w_n1556_49[0]),.dinb(w_in242_0[0]),.dout(n3295),.clk(gclk));
	jand g2654(.dina(w_n1711_49[2]),.dinb(w_in342_0[0]),.dout(n3296),.clk(gclk));
	jor g2655(.dina(n3296),.dinb(n3295),.dout(n3297),.clk(gclk));
	jand g2656(.dina(w_n3297_0[2]),.dinb(w_n3294_0[1]),.dout(n3298),.clk(gclk));
	jor g2657(.dina(n3298),.dinb(n3290),.dout(n3299),.clk(gclk));
	jand g2658(.dina(w_n2628_49[1]),.dinb(w_in044_0[0]),.dout(n3300),.clk(gclk));
	jand g2659(.dina(w_n2783_49[2]),.dinb(w_in144_0[0]),.dout(n3301),.clk(gclk));
	jor g2660(.dina(n3301),.dinb(n3300),.dout(n3302),.clk(gclk));
	jnot g2661(.din(w_n3302_0[1]),.dout(n3303),.clk(gclk));
	jand g2662(.dina(w_n1556_48[2]),.dinb(w_in244_0[0]),.dout(n3304),.clk(gclk));
	jand g2663(.dina(w_n1711_49[1]),.dinb(w_in344_0[0]),.dout(n3305),.clk(gclk));
	jor g2664(.dina(n3305),.dinb(n3304),.dout(n3306),.clk(gclk));
	jand g2665(.dina(w_n3306_0[2]),.dinb(w_n3303_0[1]),.dout(n3307),.clk(gclk));
	jand g2666(.dina(w_n2628_49[0]),.dinb(w_in040_0[0]),.dout(n3308),.clk(gclk));
	jand g2667(.dina(w_n2783_49[1]),.dinb(w_in140_0[0]),.dout(n3309),.clk(gclk));
	jor g2668(.dina(n3309),.dinb(n3308),.dout(n3310),.clk(gclk));
	jnot g2669(.din(w_n3310_0[1]),.dout(n3311),.clk(gclk));
	jand g2670(.dina(w_n1556_48[1]),.dinb(w_in240_0[0]),.dout(n3312),.clk(gclk));
	jand g2671(.dina(w_n1711_49[0]),.dinb(w_in340_0[0]),.dout(n3313),.clk(gclk));
	jor g2672(.dina(n3313),.dinb(n3312),.dout(n3314),.clk(gclk));
	jand g2673(.dina(w_n3314_0[2]),.dinb(w_n3311_0[1]),.dout(n3315),.clk(gclk));
	jand g2674(.dina(w_n2628_48[2]),.dinb(w_in041_0[0]),.dout(n3316),.clk(gclk));
	jand g2675(.dina(w_n2783_49[0]),.dinb(w_in141_0[0]),.dout(n3317),.clk(gclk));
	jor g2676(.dina(n3317),.dinb(n3316),.dout(n3318),.clk(gclk));
	jnot g2677(.din(w_n3318_0[1]),.dout(n3319),.clk(gclk));
	jand g2678(.dina(w_n1556_48[0]),.dinb(w_in241_0[0]),.dout(n3320),.clk(gclk));
	jand g2679(.dina(w_n1711_48[2]),.dinb(w_in341_0[0]),.dout(n3321),.clk(gclk));
	jor g2680(.dina(n3321),.dinb(n3320),.dout(n3322),.clk(gclk));
	jand g2681(.dina(w_n3322_0[2]),.dinb(w_n3319_0[1]),.dout(n3323),.clk(gclk));
	jor g2682(.dina(w_n3323_0[1]),.dinb(n3315),.dout(n3324),.clk(gclk));
	jor g2683(.dina(n3324),.dinb(w_n3307_0[1]),.dout(n3325),.clk(gclk));
	jor g2684(.dina(n3325),.dinb(w_n3299_0[1]),.dout(n3326),.clk(gclk));
	jor g2685(.dina(n3326),.dinb(w_n3282_0[1]),.dout(n3327),.clk(gclk));
	jor g2686(.dina(w_n3327_0[1]),.dinb(n3256),.dout(n3328),.clk(gclk));
	jor g2687(.dina(w_n3289_0[1]),.dinb(w_n3286_0[0]),.dout(n3329),.clk(gclk));
	jor g2688(.dina(w_n3314_0[1]),.dinb(w_n3311_0[0]),.dout(n3330),.clk(gclk));
	jor g2689(.dina(n3330),.dinb(w_n3323_0[0]),.dout(n3331),.clk(gclk));
	jor g2690(.dina(w_n3322_0[1]),.dinb(w_n3319_0[0]),.dout(n3332),.clk(gclk));
	jor g2691(.dina(w_n3297_0[1]),.dinb(w_n3294_0[0]),.dout(n3333),.clk(gclk));
	jand g2692(.dina(n3333),.dinb(n3332),.dout(n3334),.clk(gclk));
	jand g2693(.dina(n3334),.dinb(n3331),.dout(n3335),.clk(gclk));
	jor g2694(.dina(n3335),.dinb(w_n3299_0[0]),.dout(n3336),.clk(gclk));
	jand g2695(.dina(n3336),.dinb(n3329),.dout(n3337),.clk(gclk));
	jor g2696(.dina(n3337),.dinb(w_n3307_0[0]),.dout(n3338),.clk(gclk));
	jor g2697(.dina(w_n3306_0[1]),.dinb(w_n3303_0[0]),.dout(n3339),.clk(gclk));
	jor g2698(.dina(w_n3263_0[1]),.dinb(w_n3260_0[0]),.dout(n3340),.clk(gclk));
	jand g2699(.dina(n3340),.dinb(n3339),.dout(n3341),.clk(gclk));
	jand g2700(.dina(n3341),.dinb(n3338),.dout(n3342),.clk(gclk));
	jor g2701(.dina(n3342),.dinb(w_n3282_0[0]),.dout(n3343),.clk(gclk));
	jor g2702(.dina(w_n3279_0[0]),.dinb(w_n3275_0[1]),.dout(n3344),.clk(gclk));
	jor g2703(.dina(n3344),.dinb(w_n3272_0[0]),.dout(n3345),.clk(gclk));
	jor g2704(.dina(w_n3271_0[1]),.dinb(w_n3268_0[0]),.dout(n3346),.clk(gclk));
	jand g2705(.dina(n3346),.dinb(n3345),.dout(n3347),.clk(gclk));
	jand g2706(.dina(n3347),.dinb(n3343),.dout(n3348),.clk(gclk));
	jand g2707(.dina(w_n3348_0[1]),.dinb(n3328),.dout(n3349),.clk(gclk));
	jand g2708(.dina(w_n2628_48[1]),.dinb(w_in051_0[0]),.dout(n3350),.clk(gclk));
	jand g2709(.dina(w_n2783_48[2]),.dinb(w_in151_0[0]),.dout(n3351),.clk(gclk));
	jor g2710(.dina(n3351),.dinb(n3350),.dout(n3352),.clk(gclk));
	jnot g2711(.din(w_n3352_0[1]),.dout(n3353),.clk(gclk));
	jand g2712(.dina(w_n1556_47[2]),.dinb(w_in251_0[0]),.dout(n3354),.clk(gclk));
	jand g2713(.dina(w_n1711_48[1]),.dinb(w_in351_0[0]),.dout(n3355),.clk(gclk));
	jor g2714(.dina(n3355),.dinb(n3354),.dout(n3356),.clk(gclk));
	jand g2715(.dina(w_n3356_0[2]),.dinb(w_n3353_0[1]),.dout(n3357),.clk(gclk));
	jand g2716(.dina(w_n2628_48[0]),.dinb(w_in049_0[0]),.dout(n3358),.clk(gclk));
	jand g2717(.dina(w_n2783_48[1]),.dinb(w_in149_0[0]),.dout(n3359),.clk(gclk));
	jor g2718(.dina(n3359),.dinb(n3358),.dout(n3360),.clk(gclk));
	jnot g2719(.din(w_n3360_0[1]),.dout(n3361),.clk(gclk));
	jand g2720(.dina(w_n1556_47[1]),.dinb(w_in249_0[0]),.dout(n3362),.clk(gclk));
	jand g2721(.dina(w_n1711_48[0]),.dinb(w_in349_0[0]),.dout(n3363),.clk(gclk));
	jor g2722(.dina(n3363),.dinb(n3362),.dout(n3364),.clk(gclk));
	jand g2723(.dina(w_n3364_0[2]),.dinb(w_n3361_0[1]),.dout(n3365),.clk(gclk));
	jand g2724(.dina(w_n1556_47[0]),.dinb(w_in250_0[0]),.dout(n3366),.clk(gclk));
	jand g2725(.dina(w_n1711_47[2]),.dinb(w_in350_0[0]),.dout(n3367),.clk(gclk));
	jor g2726(.dina(n3367),.dinb(n3366),.dout(n3368),.clk(gclk));
	jand g2727(.dina(w_n2628_47[2]),.dinb(w_in050_0[0]),.dout(n3369),.clk(gclk));
	jand g2728(.dina(w_n2783_48[0]),.dinb(w_in150_0[0]),.dout(n3370),.clk(gclk));
	jor g2729(.dina(n3370),.dinb(n3369),.dout(n3371),.clk(gclk));
	jnot g2730(.din(w_n3371_0[1]),.dout(n3372),.clk(gclk));
	jand g2731(.dina(w_n3372_0[1]),.dinb(w_n3368_0[2]),.dout(n3373),.clk(gclk));
	jor g2732(.dina(n3373),.dinb(n3365),.dout(n3374),.clk(gclk));
	jor g2733(.dina(n3374),.dinb(w_n3357_0[1]),.dout(n3375),.clk(gclk));
	jand g2734(.dina(w_n2628_47[1]),.dinb(w_in053_0[0]),.dout(n3376),.clk(gclk));
	jand g2735(.dina(w_n2783_47[2]),.dinb(w_in153_0[0]),.dout(n3377),.clk(gclk));
	jor g2736(.dina(n3377),.dinb(n3376),.dout(n3378),.clk(gclk));
	jnot g2737(.din(w_n3378_0[1]),.dout(n3379),.clk(gclk));
	jand g2738(.dina(w_n1556_46[2]),.dinb(w_in253_0[0]),.dout(n3380),.clk(gclk));
	jand g2739(.dina(w_n1711_47[1]),.dinb(w_in353_0[0]),.dout(n3381),.clk(gclk));
	jor g2740(.dina(n3381),.dinb(n3380),.dout(n3382),.clk(gclk));
	jand g2741(.dina(w_n3382_0[2]),.dinb(w_n3379_0[1]),.dout(n3383),.clk(gclk));
	jnot g2742(.din(n3383),.dout(n3384),.clk(gclk));
	jand g2743(.dina(w_n2628_47[0]),.dinb(w_in052_0[0]),.dout(n3385),.clk(gclk));
	jand g2744(.dina(w_n2783_47[1]),.dinb(w_in152_0[0]),.dout(n3386),.clk(gclk));
	jor g2745(.dina(n3386),.dinb(n3385),.dout(n3387),.clk(gclk));
	jand g2746(.dina(w_n3387_0[1]),.dinb(w_n3384_0[1]),.dout(n3388),.clk(gclk));
	jand g2747(.dina(w_n1556_46[1]),.dinb(w_in252_0[0]),.dout(n3389),.clk(gclk));
	jand g2748(.dina(w_n1711_47[0]),.dinb(w_in352_0[0]),.dout(n3390),.clk(gclk));
	jor g2749(.dina(n3390),.dinb(n3389),.dout(n3391),.clk(gclk));
	jnot g2750(.din(w_n3391_0[1]),.dout(n3392),.clk(gclk));
	jand g2751(.dina(w_n3392_0[1]),.dinb(w_n3384_0[0]),.dout(n3393),.clk(gclk));
	jor g2752(.dina(n3393),.dinb(w_n3388_0[1]),.dout(n3394),.clk(gclk));
	jnot g2753(.din(n3394),.dout(n3395),.clk(gclk));
	jand g2754(.dina(w_n2628_46[2]),.dinb(w_in055_0[0]),.dout(n3396),.clk(gclk));
	jand g2755(.dina(w_n2783_47[0]),.dinb(w_in155_0[0]),.dout(n3397),.clk(gclk));
	jor g2756(.dina(n3397),.dinb(n3396),.dout(n3398),.clk(gclk));
	jnot g2757(.din(w_n3398_0[1]),.dout(n3399),.clk(gclk));
	jand g2758(.dina(w_n1556_46[0]),.dinb(w_in255_0[0]),.dout(n3400),.clk(gclk));
	jand g2759(.dina(w_n1711_46[2]),.dinb(w_in355_0[0]),.dout(n3401),.clk(gclk));
	jor g2760(.dina(n3401),.dinb(n3400),.dout(n3402),.clk(gclk));
	jand g2761(.dina(w_n3402_0[2]),.dinb(w_n3399_0[1]),.dout(n3403),.clk(gclk));
	jand g2762(.dina(w_n1556_45[2]),.dinb(w_in254_0[0]),.dout(n3404),.clk(gclk));
	jand g2763(.dina(w_n1711_46[1]),.dinb(w_in354_0[0]),.dout(n3405),.clk(gclk));
	jor g2764(.dina(n3405),.dinb(n3404),.dout(n3406),.clk(gclk));
	jand g2765(.dina(w_n2628_46[1]),.dinb(w_in054_0[0]),.dout(n3407),.clk(gclk));
	jand g2766(.dina(w_n2783_46[2]),.dinb(w_in154_0[0]),.dout(n3408),.clk(gclk));
	jor g2767(.dina(n3408),.dinb(n3407),.dout(n3409),.clk(gclk));
	jnot g2768(.din(w_n3409_0[1]),.dout(n3410),.clk(gclk));
	jand g2769(.dina(w_n3410_0[1]),.dinb(w_n3406_0[2]),.dout(n3411),.clk(gclk));
	jor g2770(.dina(n3411),.dinb(n3403),.dout(n3412),.clk(gclk));
	jand g2771(.dina(w_n1556_45[1]),.dinb(w_in248_0[0]),.dout(n3413),.clk(gclk));
	jand g2772(.dina(w_n1711_46[0]),.dinb(w_in348_0[0]),.dout(n3414),.clk(gclk));
	jor g2773(.dina(n3414),.dinb(n3413),.dout(n3415),.clk(gclk));
	jand g2774(.dina(w_n2628_46[0]),.dinb(w_in048_0[0]),.dout(n3416),.clk(gclk));
	jand g2775(.dina(w_n2783_46[1]),.dinb(w_in148_0[0]),.dout(n3417),.clk(gclk));
	jor g2776(.dina(n3417),.dinb(n3416),.dout(n3418),.clk(gclk));
	jnot g2777(.din(w_n3418_0[1]),.dout(n3419),.clk(gclk));
	jand g2778(.dina(w_n3419_0[1]),.dinb(w_n3415_0[2]),.dout(n3420),.clk(gclk));
	jor g2779(.dina(n3420),.dinb(w_n3412_0[1]),.dout(n3421),.clk(gclk));
	jor g2780(.dina(n3421),.dinb(w_n3395_0[1]),.dout(n3422),.clk(gclk));
	jor g2781(.dina(n3422),.dinb(w_n3375_0[1]),.dout(n3423),.clk(gclk));
	jor g2782(.dina(w_n3423_0[1]),.dinb(n3349),.dout(n3424),.clk(gclk));
	jor g2783(.dina(w_n3402_0[1]),.dinb(w_n3399_0[0]),.dout(n3425),.clk(gclk));
	jor g2784(.dina(w_n3419_0[0]),.dinb(w_n3415_0[1]),.dout(n3426),.clk(gclk));
	jor g2785(.dina(w_n3364_0[1]),.dinb(w_n3361_0[0]),.dout(n3427),.clk(gclk));
	jand g2786(.dina(n3427),.dinb(n3426),.dout(n3428),.clk(gclk));
	jor g2787(.dina(n3428),.dinb(w_n3375_0[0]),.dout(n3429),.clk(gclk));
	jor g2788(.dina(w_n3372_0[0]),.dinb(w_n3368_0[1]),.dout(n3430),.clk(gclk));
	jor g2789(.dina(n3430),.dinb(w_n3357_0[0]),.dout(n3431),.clk(gclk));
	jor g2790(.dina(w_n3356_0[1]),.dinb(w_n3353_0[0]),.dout(n3432),.clk(gclk));
	jand g2791(.dina(n3432),.dinb(n3431),.dout(n3433),.clk(gclk));
	jand g2792(.dina(n3433),.dinb(n3429),.dout(n3434),.clk(gclk));
	jor g2793(.dina(n3434),.dinb(w_n3395_0[0]),.dout(n3435),.clk(gclk));
	jand g2794(.dina(w_n3392_0[0]),.dinb(w_n3388_0[0]),.dout(n3436),.clk(gclk));
	jnot g2795(.din(n3436),.dout(n3437),.clk(gclk));
	jor g2796(.dina(w_n3382_0[1]),.dinb(w_n3379_0[0]),.dout(n3438),.clk(gclk));
	jor g2797(.dina(w_n3410_0[0]),.dinb(w_n3406_0[1]),.dout(n3439),.clk(gclk));
	jand g2798(.dina(n3439),.dinb(n3438),.dout(n3440),.clk(gclk));
	jand g2799(.dina(n3440),.dinb(n3437),.dout(n3441),.clk(gclk));
	jand g2800(.dina(n3441),.dinb(n3435),.dout(n3442),.clk(gclk));
	jor g2801(.dina(n3442),.dinb(w_n3412_0[0]),.dout(n3443),.clk(gclk));
	jand g2802(.dina(n3443),.dinb(n3425),.dout(n3444),.clk(gclk));
	jand g2803(.dina(w_n3444_0[1]),.dinb(n3424),.dout(n3445),.clk(gclk));
	jand g2804(.dina(w_n2628_45[2]),.dinb(w_in061_0[0]),.dout(n3446),.clk(gclk));
	jand g2805(.dina(w_n2783_46[0]),.dinb(w_in161_0[0]),.dout(n3447),.clk(gclk));
	jor g2806(.dina(n3447),.dinb(n3446),.dout(n3448),.clk(gclk));
	jnot g2807(.din(w_n3448_0[1]),.dout(n3449),.clk(gclk));
	jand g2808(.dina(w_n1556_45[0]),.dinb(w_in261_0[0]),.dout(n3450),.clk(gclk));
	jand g2809(.dina(w_n1711_45[2]),.dinb(w_in361_0[0]),.dout(n3451),.clk(gclk));
	jor g2810(.dina(n3451),.dinb(n3450),.dout(n3452),.clk(gclk));
	jand g2811(.dina(w_n3452_0[2]),.dinb(w_n3449_0[1]),.dout(n3453),.clk(gclk));
	jand g2812(.dina(w_n2628_45[1]),.dinb(w_in063_0[0]),.dout(n3454),.clk(gclk));
	jand g2813(.dina(w_n2783_45[2]),.dinb(w_in163_0[0]),.dout(n3455),.clk(gclk));
	jor g2814(.dina(n3455),.dinb(n3454),.dout(n3456),.clk(gclk));
	jnot g2815(.din(w_n3456_0[1]),.dout(n3457),.clk(gclk));
	jand g2816(.dina(w_n1556_44[2]),.dinb(w_in263_0[0]),.dout(n3458),.clk(gclk));
	jand g2817(.dina(w_n1711_45[1]),.dinb(w_in363_0[0]),.dout(n3459),.clk(gclk));
	jor g2818(.dina(n3459),.dinb(n3458),.dout(n3460),.clk(gclk));
	jand g2819(.dina(w_n3460_0[2]),.dinb(w_n3457_0[1]),.dout(n3461),.clk(gclk));
	jand g2820(.dina(w_n1556_44[1]),.dinb(w_in262_0[0]),.dout(n3462),.clk(gclk));
	jand g2821(.dina(w_n1711_45[0]),.dinb(w_in362_0[0]),.dout(n3463),.clk(gclk));
	jor g2822(.dina(n3463),.dinb(n3462),.dout(n3464),.clk(gclk));
	jand g2823(.dina(w_n2628_45[0]),.dinb(w_in062_0[0]),.dout(n3465),.clk(gclk));
	jand g2824(.dina(w_n2783_45[1]),.dinb(w_in162_0[0]),.dout(n3466),.clk(gclk));
	jor g2825(.dina(n3466),.dinb(n3465),.dout(n3467),.clk(gclk));
	jnot g2826(.din(w_n3467_0[1]),.dout(n3468),.clk(gclk));
	jand g2827(.dina(w_n3468_0[1]),.dinb(w_n3464_0[2]),.dout(n3469),.clk(gclk));
	jor g2828(.dina(n3469),.dinb(w_n3461_0[1]),.dout(n3470),.clk(gclk));
	jor g2829(.dina(n3470),.dinb(n3453),.dout(n3471),.clk(gclk));
	jand g2830(.dina(w_n2628_44[2]),.dinb(w_in059_0[0]),.dout(n3472),.clk(gclk));
	jand g2831(.dina(w_n2783_45[0]),.dinb(w_in159_0[0]),.dout(n3473),.clk(gclk));
	jor g2832(.dina(n3473),.dinb(n3472),.dout(n3474),.clk(gclk));
	jnot g2833(.din(w_n3474_0[1]),.dout(n3475),.clk(gclk));
	jand g2834(.dina(w_n1556_44[0]),.dinb(w_in259_0[0]),.dout(n3476),.clk(gclk));
	jand g2835(.dina(w_n1711_44[2]),.dinb(w_in359_0[0]),.dout(n3477),.clk(gclk));
	jor g2836(.dina(n3477),.dinb(n3476),.dout(n3478),.clk(gclk));
	jand g2837(.dina(w_n3478_0[2]),.dinb(w_n3475_0[1]),.dout(n3479),.clk(gclk));
	jand g2838(.dina(w_n2628_44[1]),.dinb(w_in058_0[0]),.dout(n3480),.clk(gclk));
	jand g2839(.dina(w_n2783_44[2]),.dinb(w_in158_0[0]),.dout(n3481),.clk(gclk));
	jor g2840(.dina(n3481),.dinb(n3480),.dout(n3482),.clk(gclk));
	jnot g2841(.din(w_n3482_0[1]),.dout(n3483),.clk(gclk));
	jand g2842(.dina(w_n1556_43[2]),.dinb(w_in258_0[0]),.dout(n3484),.clk(gclk));
	jand g2843(.dina(w_n1711_44[1]),.dinb(w_in358_0[0]),.dout(n3485),.clk(gclk));
	jor g2844(.dina(n3485),.dinb(n3484),.dout(n3486),.clk(gclk));
	jand g2845(.dina(w_n3486_0[2]),.dinb(w_n3483_0[1]),.dout(n3487),.clk(gclk));
	jor g2846(.dina(n3487),.dinb(n3479),.dout(n3488),.clk(gclk));
	jand g2847(.dina(w_n2628_44[0]),.dinb(w_in060_0[0]),.dout(n3489),.clk(gclk));
	jand g2848(.dina(w_n2783_44[1]),.dinb(w_in160_0[0]),.dout(n3490),.clk(gclk));
	jor g2849(.dina(n3490),.dinb(n3489),.dout(n3491),.clk(gclk));
	jnot g2850(.din(w_n3491_0[1]),.dout(n3492),.clk(gclk));
	jand g2851(.dina(w_n1556_43[1]),.dinb(w_in260_0[0]),.dout(n3493),.clk(gclk));
	jand g2852(.dina(w_n1711_44[0]),.dinb(w_in360_0[0]),.dout(n3494),.clk(gclk));
	jor g2853(.dina(n3494),.dinb(n3493),.dout(n3495),.clk(gclk));
	jand g2854(.dina(w_n3495_0[2]),.dinb(w_n3492_0[1]),.dout(n3496),.clk(gclk));
	jand g2855(.dina(w_n2628_43[2]),.dinb(w_in056_0[0]),.dout(n3497),.clk(gclk));
	jand g2856(.dina(w_n2783_44[0]),.dinb(w_in156_0[0]),.dout(n3498),.clk(gclk));
	jor g2857(.dina(n3498),.dinb(n3497),.dout(n3499),.clk(gclk));
	jnot g2858(.din(w_n3499_0[1]),.dout(n3500),.clk(gclk));
	jand g2859(.dina(w_n1556_43[0]),.dinb(w_in256_0[0]),.dout(n3501),.clk(gclk));
	jand g2860(.dina(w_n1711_43[2]),.dinb(w_in356_0[0]),.dout(n3502),.clk(gclk));
	jor g2861(.dina(n3502),.dinb(n3501),.dout(n3503),.clk(gclk));
	jand g2862(.dina(w_n3503_0[2]),.dinb(w_n3500_0[1]),.dout(n3504),.clk(gclk));
	jand g2863(.dina(w_n2628_43[1]),.dinb(w_in057_0[0]),.dout(n3505),.clk(gclk));
	jand g2864(.dina(w_n2783_43[2]),.dinb(w_in157_0[0]),.dout(n3506),.clk(gclk));
	jor g2865(.dina(n3506),.dinb(n3505),.dout(n3507),.clk(gclk));
	jnot g2866(.din(w_n3507_0[1]),.dout(n3508),.clk(gclk));
	jand g2867(.dina(w_n1556_42[2]),.dinb(w_in257_0[0]),.dout(n3509),.clk(gclk));
	jand g2868(.dina(w_n1711_43[1]),.dinb(w_in357_0[0]),.dout(n3510),.clk(gclk));
	jor g2869(.dina(n3510),.dinb(n3509),.dout(n3511),.clk(gclk));
	jand g2870(.dina(w_n3511_0[2]),.dinb(w_n3508_0[1]),.dout(n3512),.clk(gclk));
	jor g2871(.dina(w_n3512_0[1]),.dinb(n3504),.dout(n3513),.clk(gclk));
	jor g2872(.dina(n3513),.dinb(w_n3496_0[1]),.dout(n3514),.clk(gclk));
	jor g2873(.dina(n3514),.dinb(w_n3488_0[1]),.dout(n3515),.clk(gclk));
	jor g2874(.dina(n3515),.dinb(w_n3471_0[1]),.dout(n3516),.clk(gclk));
	jor g2875(.dina(w_n3516_0[1]),.dinb(n3445),.dout(n3517),.clk(gclk));
	jor g2876(.dina(w_n3478_0[1]),.dinb(w_n3475_0[0]),.dout(n3518),.clk(gclk));
	jor g2877(.dina(w_n3503_0[1]),.dinb(w_n3500_0[0]),.dout(n3519),.clk(gclk));
	jor g2878(.dina(n3519),.dinb(w_n3512_0[0]),.dout(n3520),.clk(gclk));
	jor g2879(.dina(w_n3511_0[1]),.dinb(w_n3508_0[0]),.dout(n3521),.clk(gclk));
	jor g2880(.dina(w_n3486_0[1]),.dinb(w_n3483_0[0]),.dout(n3522),.clk(gclk));
	jand g2881(.dina(n3522),.dinb(n3521),.dout(n3523),.clk(gclk));
	jand g2882(.dina(n3523),.dinb(n3520),.dout(n3524),.clk(gclk));
	jor g2883(.dina(n3524),.dinb(w_n3488_0[0]),.dout(n3525),.clk(gclk));
	jand g2884(.dina(n3525),.dinb(n3518),.dout(n3526),.clk(gclk));
	jor g2885(.dina(n3526),.dinb(w_n3496_0[0]),.dout(n3527),.clk(gclk));
	jor g2886(.dina(w_n3495_0[1]),.dinb(w_n3492_0[0]),.dout(n3528),.clk(gclk));
	jor g2887(.dina(w_n3452_0[1]),.dinb(w_n3449_0[0]),.dout(n3529),.clk(gclk));
	jand g2888(.dina(n3529),.dinb(n3528),.dout(n3530),.clk(gclk));
	jand g2889(.dina(n3530),.dinb(n3527),.dout(n3531),.clk(gclk));
	jor g2890(.dina(n3531),.dinb(w_n3471_0[0]),.dout(n3532),.clk(gclk));
	jor g2891(.dina(w_n3468_0[0]),.dinb(w_n3464_0[1]),.dout(n3533),.clk(gclk));
	jor g2892(.dina(n3533),.dinb(w_n3461_0[0]),.dout(n3534),.clk(gclk));
	jor g2893(.dina(w_n3460_0[1]),.dinb(w_n3457_0[0]),.dout(n3535),.clk(gclk));
	jand g2894(.dina(n3535),.dinb(n3534),.dout(n3536),.clk(gclk));
	jand g2895(.dina(n3536),.dinb(n3532),.dout(n3537),.clk(gclk));
	jand g2896(.dina(w_n3537_0[1]),.dinb(n3517),.dout(n3538),.clk(gclk));
	jand g2897(.dina(w_n2628_43[0]),.dinb(w_in067_0[0]),.dout(n3539),.clk(gclk));
	jand g2898(.dina(w_n2783_43[1]),.dinb(w_in167_0[0]),.dout(n3540),.clk(gclk));
	jor g2899(.dina(n3540),.dinb(n3539),.dout(n3541),.clk(gclk));
	jnot g2900(.din(w_n3541_0[1]),.dout(n3542),.clk(gclk));
	jand g2901(.dina(w_n1556_42[1]),.dinb(w_in267_0[0]),.dout(n3543),.clk(gclk));
	jand g2902(.dina(w_n1711_43[0]),.dinb(w_in367_0[0]),.dout(n3544),.clk(gclk));
	jor g2903(.dina(n3544),.dinb(n3543),.dout(n3545),.clk(gclk));
	jand g2904(.dina(w_n3545_0[2]),.dinb(w_n3542_0[1]),.dout(n3546),.clk(gclk));
	jand g2905(.dina(w_n1556_42[0]),.dinb(w_in266_0[0]),.dout(n3547),.clk(gclk));
	jand g2906(.dina(w_n1711_42[2]),.dinb(w_in366_0[0]),.dout(n3548),.clk(gclk));
	jor g2907(.dina(n3548),.dinb(n3547),.dout(n3549),.clk(gclk));
	jand g2908(.dina(w_n2628_42[2]),.dinb(w_in066_0[0]),.dout(n3550),.clk(gclk));
	jand g2909(.dina(w_n2783_43[0]),.dinb(w_in166_0[0]),.dout(n3551),.clk(gclk));
	jor g2910(.dina(n3551),.dinb(n3550),.dout(n3552),.clk(gclk));
	jnot g2911(.din(w_n3552_0[1]),.dout(n3553),.clk(gclk));
	jand g2912(.dina(w_n3553_0[1]),.dinb(w_n3549_0[2]),.dout(n3554),.clk(gclk));
	jor g2913(.dina(n3554),.dinb(n3546),.dout(n3555),.clk(gclk));
	jand g2914(.dina(w_n2628_42[1]),.dinb(w_in065_0[0]),.dout(n3556),.clk(gclk));
	jand g2915(.dina(w_n2783_42[2]),.dinb(w_in165_0[0]),.dout(n3557),.clk(gclk));
	jor g2916(.dina(n3557),.dinb(n3556),.dout(n3558),.clk(gclk));
	jnot g2917(.din(w_n3558_0[1]),.dout(n3559),.clk(gclk));
	jand g2918(.dina(w_n1556_41[2]),.dinb(w_in265_0[0]),.dout(n3560),.clk(gclk));
	jand g2919(.dina(w_n1711_42[1]),.dinb(w_in365_0[0]),.dout(n3561),.clk(gclk));
	jor g2920(.dina(n3561),.dinb(n3560),.dout(n3562),.clk(gclk));
	jand g2921(.dina(w_n3562_0[2]),.dinb(w_n3559_0[1]),.dout(n3563),.clk(gclk));
	jand g2922(.dina(w_n1556_41[1]),.dinb(w_in264_0[0]),.dout(n3564),.clk(gclk));
	jand g2923(.dina(w_n1711_42[0]),.dinb(w_in364_0[0]),.dout(n3565),.clk(gclk));
	jor g2924(.dina(n3565),.dinb(n3564),.dout(n3566),.clk(gclk));
	jand g2925(.dina(w_n2628_42[0]),.dinb(w_in064_0[0]),.dout(n3567),.clk(gclk));
	jand g2926(.dina(w_n2783_42[1]),.dinb(w_in164_0[0]),.dout(n3568),.clk(gclk));
	jor g2927(.dina(n3568),.dinb(n3567),.dout(n3569),.clk(gclk));
	jnot g2928(.din(w_n3569_0[1]),.dout(n3570),.clk(gclk));
	jand g2929(.dina(w_n3570_0[1]),.dinb(w_n3566_0[2]),.dout(n3571),.clk(gclk));
	jor g2930(.dina(n3571),.dinb(w_n3563_0[1]),.dout(n3572),.clk(gclk));
	jor g2931(.dina(n3572),.dinb(w_n3555_0[1]),.dout(n3573),.clk(gclk));
	jor g2932(.dina(w_n3573_0[1]),.dinb(n3538),.dout(n3574),.clk(gclk));
	jor g2933(.dina(w_n3545_0[1]),.dinb(w_n3542_0[0]),.dout(n3575),.clk(gclk));
	jor g2934(.dina(w_n3570_0[0]),.dinb(w_n3566_0[1]),.dout(n3576),.clk(gclk));
	jor g2935(.dina(n3576),.dinb(w_n3563_0[0]),.dout(n3577),.clk(gclk));
	jor g2936(.dina(w_n3562_0[1]),.dinb(w_n3559_0[0]),.dout(n3578),.clk(gclk));
	jor g2937(.dina(w_n3553_0[0]),.dinb(w_n3549_0[1]),.dout(n3579),.clk(gclk));
	jand g2938(.dina(n3579),.dinb(n3578),.dout(n3580),.clk(gclk));
	jand g2939(.dina(n3580),.dinb(n3577),.dout(n3581),.clk(gclk));
	jor g2940(.dina(n3581),.dinb(w_n3555_0[0]),.dout(n3582),.clk(gclk));
	jand g2941(.dina(n3582),.dinb(n3575),.dout(n3583),.clk(gclk));
	jand g2942(.dina(w_n3583_0[1]),.dinb(n3574),.dout(n3584),.clk(gclk));
	jand g2943(.dina(w_n2628_41[2]),.dinb(w_in068_0[0]),.dout(n3585),.clk(gclk));
	jand g2944(.dina(w_n2783_42[0]),.dinb(w_in168_0[0]),.dout(n3586),.clk(gclk));
	jor g2945(.dina(n3586),.dinb(n3585),.dout(n3587),.clk(gclk));
	jnot g2946(.din(w_n3587_0[1]),.dout(n3588),.clk(gclk));
	jand g2947(.dina(w_n1556_41[0]),.dinb(w_in268_0[0]),.dout(n3589),.clk(gclk));
	jand g2948(.dina(w_n1711_41[2]),.dinb(w_in368_0[0]),.dout(n3590),.clk(gclk));
	jor g2949(.dina(n3590),.dinb(n3589),.dout(n3591),.clk(gclk));
	jand g2950(.dina(w_n3591_0[2]),.dinb(w_n3588_0[1]),.dout(n3592),.clk(gclk));
	jand g2951(.dina(w_n2628_41[1]),.dinb(w_in069_0[0]),.dout(n3593),.clk(gclk));
	jand g2952(.dina(w_n2783_41[2]),.dinb(w_in169_0[0]),.dout(n3594),.clk(gclk));
	jor g2953(.dina(n3594),.dinb(n3593),.dout(n3595),.clk(gclk));
	jnot g2954(.din(w_n3595_0[1]),.dout(n3596),.clk(gclk));
	jand g2955(.dina(w_n1556_40[2]),.dinb(w_in269_0[0]),.dout(n3597),.clk(gclk));
	jand g2956(.dina(w_n1711_41[1]),.dinb(w_in369_0[0]),.dout(n3598),.clk(gclk));
	jor g2957(.dina(n3598),.dinb(n3597),.dout(n3599),.clk(gclk));
	jand g2958(.dina(w_n3599_0[2]),.dinb(w_n3596_0[1]),.dout(n3600),.clk(gclk));
	jand g2959(.dina(w_n2628_41[0]),.dinb(w_in071_0[0]),.dout(n3601),.clk(gclk));
	jand g2960(.dina(w_n2783_41[1]),.dinb(w_in171_0[0]),.dout(n3602),.clk(gclk));
	jor g2961(.dina(n3602),.dinb(n3601),.dout(n3603),.clk(gclk));
	jnot g2962(.din(w_n3603_0[1]),.dout(n3604),.clk(gclk));
	jand g2963(.dina(w_n1556_40[1]),.dinb(w_in271_0[0]),.dout(n3605),.clk(gclk));
	jand g2964(.dina(w_n1711_41[0]),.dinb(w_in371_0[0]),.dout(n3606),.clk(gclk));
	jor g2965(.dina(n3606),.dinb(n3605),.dout(n3607),.clk(gclk));
	jand g2966(.dina(w_n3607_0[2]),.dinb(w_n3604_0[1]),.dout(n3608),.clk(gclk));
	jand g2967(.dina(w_n1556_40[0]),.dinb(w_in270_0[0]),.dout(n3609),.clk(gclk));
	jand g2968(.dina(w_n1711_40[2]),.dinb(w_in370_0[0]),.dout(n3610),.clk(gclk));
	jor g2969(.dina(n3610),.dinb(n3609),.dout(n3611),.clk(gclk));
	jand g2970(.dina(w_n2628_40[2]),.dinb(w_in070_0[0]),.dout(n3612),.clk(gclk));
	jand g2971(.dina(w_n2783_41[0]),.dinb(w_in170_0[0]),.dout(n3613),.clk(gclk));
	jor g2972(.dina(n3613),.dinb(n3612),.dout(n3614),.clk(gclk));
	jnot g2973(.din(w_n3614_0[1]),.dout(n3615),.clk(gclk));
	jand g2974(.dina(w_n3615_0[1]),.dinb(w_n3611_0[2]),.dout(n3616),.clk(gclk));
	jor g2975(.dina(n3616),.dinb(w_n3608_0[1]),.dout(n3617),.clk(gclk));
	jor g2976(.dina(n3617),.dinb(n3600),.dout(n3618),.clk(gclk));
	jor g2977(.dina(w_n3618_0[1]),.dinb(n3592),.dout(n3619),.clk(gclk));
	jor g2978(.dina(w_n3619_0[1]),.dinb(n3584),.dout(n3620),.clk(gclk));
	jor g2979(.dina(w_n3599_0[1]),.dinb(w_n3596_0[0]),.dout(n3621),.clk(gclk));
	jor g2980(.dina(w_n3591_0[1]),.dinb(w_n3588_0[0]),.dout(n3622),.clk(gclk));
	jand g2981(.dina(n3622),.dinb(n3621),.dout(n3623),.clk(gclk));
	jor g2982(.dina(n3623),.dinb(w_n3618_0[0]),.dout(n3624),.clk(gclk));
	jor g2983(.dina(w_n3607_0[1]),.dinb(w_n3604_0[0]),.dout(n3625),.clk(gclk));
	jor g2984(.dina(w_n3615_0[0]),.dinb(w_n3611_0[1]),.dout(n3626),.clk(gclk));
	jor g2985(.dina(n3626),.dinb(w_n3608_0[0]),.dout(n3627),.clk(gclk));
	jand g2986(.dina(n3627),.dinb(n3625),.dout(n3628),.clk(gclk));
	jand g2987(.dina(n3628),.dinb(n3624),.dout(n3629),.clk(gclk));
	jand g2988(.dina(w_n3629_0[1]),.dinb(n3620),.dout(n3630),.clk(gclk));
	jand g2989(.dina(w_n2628_40[1]),.dinb(w_in075_0[0]),.dout(n3631),.clk(gclk));
	jand g2990(.dina(w_n2783_40[2]),.dinb(w_in175_0[0]),.dout(n3632),.clk(gclk));
	jor g2991(.dina(n3632),.dinb(n3631),.dout(n3633),.clk(gclk));
	jnot g2992(.din(w_n3633_0[1]),.dout(n3634),.clk(gclk));
	jand g2993(.dina(w_n1556_39[2]),.dinb(w_in275_0[0]),.dout(n3635),.clk(gclk));
	jand g2994(.dina(w_n1711_40[1]),.dinb(w_in375_0[0]),.dout(n3636),.clk(gclk));
	jor g2995(.dina(n3636),.dinb(n3635),.dout(n3637),.clk(gclk));
	jand g2996(.dina(w_n3637_0[2]),.dinb(w_n3634_0[1]),.dout(n3638),.clk(gclk));
	jand g2997(.dina(w_n1556_39[1]),.dinb(w_in274_0[0]),.dout(n3639),.clk(gclk));
	jand g2998(.dina(w_n1711_40[0]),.dinb(w_in374_0[0]),.dout(n3640),.clk(gclk));
	jor g2999(.dina(n3640),.dinb(n3639),.dout(n3641),.clk(gclk));
	jand g3000(.dina(w_n2628_40[0]),.dinb(w_in074_0[0]),.dout(n3642),.clk(gclk));
	jand g3001(.dina(w_n2783_40[1]),.dinb(w_in174_0[0]),.dout(n3643),.clk(gclk));
	jor g3002(.dina(n3643),.dinb(n3642),.dout(n3644),.clk(gclk));
	jnot g3003(.din(w_n3644_0[1]),.dout(n3645),.clk(gclk));
	jand g3004(.dina(w_n3645_0[1]),.dinb(w_n3641_0[2]),.dout(n3646),.clk(gclk));
	jor g3005(.dina(n3646),.dinb(n3638),.dout(n3647),.clk(gclk));
	jand g3006(.dina(w_n2628_39[2]),.dinb(w_in073_0[0]),.dout(n3648),.clk(gclk));
	jand g3007(.dina(w_n2783_40[0]),.dinb(w_in173_0[0]),.dout(n3649),.clk(gclk));
	jor g3008(.dina(n3649),.dinb(n3648),.dout(n3650),.clk(gclk));
	jnot g3009(.din(w_n3650_0[1]),.dout(n3651),.clk(gclk));
	jand g3010(.dina(w_n1556_39[0]),.dinb(w_in273_0[0]),.dout(n3652),.clk(gclk));
	jand g3011(.dina(w_n1711_39[2]),.dinb(w_in373_0[0]),.dout(n3653),.clk(gclk));
	jor g3012(.dina(n3653),.dinb(n3652),.dout(n3654),.clk(gclk));
	jand g3013(.dina(w_n3654_0[2]),.dinb(w_n3651_0[1]),.dout(n3655),.clk(gclk));
	jand g3014(.dina(w_n1556_38[2]),.dinb(w_in272_0[0]),.dout(n3656),.clk(gclk));
	jand g3015(.dina(w_n1711_39[1]),.dinb(w_in372_0[0]),.dout(n3657),.clk(gclk));
	jor g3016(.dina(n3657),.dinb(n3656),.dout(n3658),.clk(gclk));
	jand g3017(.dina(w_n2628_39[1]),.dinb(w_in072_0[0]),.dout(n3659),.clk(gclk));
	jand g3018(.dina(w_n2783_39[2]),.dinb(w_in172_0[0]),.dout(n3660),.clk(gclk));
	jor g3019(.dina(n3660),.dinb(n3659),.dout(n3661),.clk(gclk));
	jnot g3020(.din(w_n3661_0[1]),.dout(n3662),.clk(gclk));
	jand g3021(.dina(w_n3662_0[1]),.dinb(w_n3658_0[2]),.dout(n3663),.clk(gclk));
	jor g3022(.dina(n3663),.dinb(w_n3655_0[1]),.dout(n3664),.clk(gclk));
	jor g3023(.dina(n3664),.dinb(w_n3647_0[1]),.dout(n3665),.clk(gclk));
	jor g3024(.dina(w_n3665_0[1]),.dinb(n3630),.dout(n3666),.clk(gclk));
	jor g3025(.dina(w_n3637_0[1]),.dinb(w_n3634_0[0]),.dout(n3667),.clk(gclk));
	jor g3026(.dina(w_n3662_0[0]),.dinb(w_n3658_0[1]),.dout(n3668),.clk(gclk));
	jor g3027(.dina(n3668),.dinb(w_n3655_0[0]),.dout(n3669),.clk(gclk));
	jor g3028(.dina(w_n3654_0[1]),.dinb(w_n3651_0[0]),.dout(n3670),.clk(gclk));
	jor g3029(.dina(w_n3645_0[0]),.dinb(w_n3641_0[1]),.dout(n3671),.clk(gclk));
	jand g3030(.dina(n3671),.dinb(n3670),.dout(n3672),.clk(gclk));
	jand g3031(.dina(n3672),.dinb(n3669),.dout(n3673),.clk(gclk));
	jor g3032(.dina(n3673),.dinb(w_n3647_0[0]),.dout(n3674),.clk(gclk));
	jand g3033(.dina(n3674),.dinb(n3667),.dout(n3675),.clk(gclk));
	jand g3034(.dina(w_n3675_0[1]),.dinb(n3666),.dout(n3676),.clk(gclk));
	jand g3035(.dina(w_n2628_39[0]),.dinb(w_in076_0[0]),.dout(n3677),.clk(gclk));
	jand g3036(.dina(w_n2783_39[1]),.dinb(w_in176_0[0]),.dout(n3678),.clk(gclk));
	jor g3037(.dina(n3678),.dinb(n3677),.dout(n3679),.clk(gclk));
	jnot g3038(.din(w_n3679_0[1]),.dout(n3680),.clk(gclk));
	jand g3039(.dina(w_n1556_38[1]),.dinb(w_in276_0[0]),.dout(n3681),.clk(gclk));
	jand g3040(.dina(w_n1711_39[0]),.dinb(w_in376_0[0]),.dout(n3682),.clk(gclk));
	jor g3041(.dina(n3682),.dinb(n3681),.dout(n3683),.clk(gclk));
	jand g3042(.dina(w_n3683_0[2]),.dinb(w_n3680_0[1]),.dout(n3684),.clk(gclk));
	jand g3043(.dina(w_n2628_38[2]),.dinb(w_in077_0[0]),.dout(n3685),.clk(gclk));
	jand g3044(.dina(w_n2783_39[0]),.dinb(w_in177_0[0]),.dout(n3686),.clk(gclk));
	jor g3045(.dina(n3686),.dinb(n3685),.dout(n3687),.clk(gclk));
	jnot g3046(.din(w_n3687_0[1]),.dout(n3688),.clk(gclk));
	jand g3047(.dina(w_n1556_38[0]),.dinb(w_in277_0[0]),.dout(n3689),.clk(gclk));
	jand g3048(.dina(w_n1711_38[2]),.dinb(w_in377_0[0]),.dout(n3690),.clk(gclk));
	jor g3049(.dina(n3690),.dinb(n3689),.dout(n3691),.clk(gclk));
	jand g3050(.dina(w_n3691_0[2]),.dinb(w_n3688_0[1]),.dout(n3692),.clk(gclk));
	jand g3051(.dina(w_n2628_38[1]),.dinb(w_in079_0[0]),.dout(n3693),.clk(gclk));
	jand g3052(.dina(w_n2783_38[2]),.dinb(w_in179_0[0]),.dout(n3694),.clk(gclk));
	jor g3053(.dina(n3694),.dinb(n3693),.dout(n3695),.clk(gclk));
	jnot g3054(.din(w_n3695_0[1]),.dout(n3696),.clk(gclk));
	jand g3055(.dina(w_n1556_37[2]),.dinb(w_in279_0[0]),.dout(n3697),.clk(gclk));
	jand g3056(.dina(w_n1711_38[1]),.dinb(w_in379_0[0]),.dout(n3698),.clk(gclk));
	jor g3057(.dina(n3698),.dinb(n3697),.dout(n3699),.clk(gclk));
	jand g3058(.dina(w_n3699_0[2]),.dinb(w_n3696_0[1]),.dout(n3700),.clk(gclk));
	jand g3059(.dina(w_n1556_37[1]),.dinb(w_in278_0[0]),.dout(n3701),.clk(gclk));
	jand g3060(.dina(w_n1711_38[0]),.dinb(w_in378_0[0]),.dout(n3702),.clk(gclk));
	jor g3061(.dina(n3702),.dinb(n3701),.dout(n3703),.clk(gclk));
	jand g3062(.dina(w_n2628_38[0]),.dinb(w_in078_0[0]),.dout(n3704),.clk(gclk));
	jand g3063(.dina(w_n2783_38[1]),.dinb(w_in178_0[0]),.dout(n3705),.clk(gclk));
	jor g3064(.dina(n3705),.dinb(n3704),.dout(n3706),.clk(gclk));
	jnot g3065(.din(w_n3706_0[1]),.dout(n3707),.clk(gclk));
	jand g3066(.dina(w_n3707_0[1]),.dinb(w_n3703_0[2]),.dout(n3708),.clk(gclk));
	jor g3067(.dina(n3708),.dinb(w_n3700_0[1]),.dout(n3709),.clk(gclk));
	jor g3068(.dina(n3709),.dinb(n3692),.dout(n3710),.clk(gclk));
	jor g3069(.dina(w_n3710_0[1]),.dinb(n3684),.dout(n3711),.clk(gclk));
	jor g3070(.dina(w_n3711_0[1]),.dinb(n3676),.dout(n3712),.clk(gclk));
	jor g3071(.dina(w_n3691_0[1]),.dinb(w_n3688_0[0]),.dout(n3713),.clk(gclk));
	jor g3072(.dina(w_n3683_0[1]),.dinb(w_n3680_0[0]),.dout(n3714),.clk(gclk));
	jand g3073(.dina(n3714),.dinb(n3713),.dout(n3715),.clk(gclk));
	jor g3074(.dina(n3715),.dinb(w_n3710_0[0]),.dout(n3716),.clk(gclk));
	jor g3075(.dina(w_n3699_0[1]),.dinb(w_n3696_0[0]),.dout(n3717),.clk(gclk));
	jor g3076(.dina(w_n3707_0[0]),.dinb(w_n3703_0[1]),.dout(n3718),.clk(gclk));
	jor g3077(.dina(n3718),.dinb(w_n3700_0[0]),.dout(n3719),.clk(gclk));
	jand g3078(.dina(n3719),.dinb(n3717),.dout(n3720),.clk(gclk));
	jand g3079(.dina(n3720),.dinb(n3716),.dout(n3721),.clk(gclk));
	jand g3080(.dina(w_n3721_0[1]),.dinb(n3712),.dout(n3722),.clk(gclk));
	jand g3081(.dina(w_n2628_37[2]),.dinb(w_in083_0[0]),.dout(n3723),.clk(gclk));
	jand g3082(.dina(w_n2783_38[0]),.dinb(w_in183_0[0]),.dout(n3724),.clk(gclk));
	jor g3083(.dina(n3724),.dinb(n3723),.dout(n3725),.clk(gclk));
	jnot g3084(.din(w_n3725_0[1]),.dout(n3726),.clk(gclk));
	jand g3085(.dina(w_n1556_37[0]),.dinb(w_in283_0[0]),.dout(n3727),.clk(gclk));
	jand g3086(.dina(w_n1711_37[2]),.dinb(w_in383_0[0]),.dout(n3728),.clk(gclk));
	jor g3087(.dina(n3728),.dinb(n3727),.dout(n3729),.clk(gclk));
	jand g3088(.dina(w_n3729_0[2]),.dinb(w_n3726_0[1]),.dout(n3730),.clk(gclk));
	jand g3089(.dina(w_n1556_36[2]),.dinb(w_in282_0[0]),.dout(n3731),.clk(gclk));
	jand g3090(.dina(w_n1711_37[1]),.dinb(w_in382_0[0]),.dout(n3732),.clk(gclk));
	jor g3091(.dina(n3732),.dinb(n3731),.dout(n3733),.clk(gclk));
	jand g3092(.dina(w_n2628_37[1]),.dinb(w_in082_0[0]),.dout(n3734),.clk(gclk));
	jand g3093(.dina(w_n2783_37[2]),.dinb(w_in182_0[0]),.dout(n3735),.clk(gclk));
	jor g3094(.dina(n3735),.dinb(n3734),.dout(n3736),.clk(gclk));
	jnot g3095(.din(w_n3736_0[1]),.dout(n3737),.clk(gclk));
	jand g3096(.dina(w_n3737_0[1]),.dinb(w_n3733_0[2]),.dout(n3738),.clk(gclk));
	jor g3097(.dina(n3738),.dinb(n3730),.dout(n3739),.clk(gclk));
	jand g3098(.dina(w_n2628_37[0]),.dinb(w_in081_0[0]),.dout(n3740),.clk(gclk));
	jand g3099(.dina(w_n2783_37[1]),.dinb(w_in181_0[0]),.dout(n3741),.clk(gclk));
	jor g3100(.dina(n3741),.dinb(n3740),.dout(n3742),.clk(gclk));
	jnot g3101(.din(w_n3742_0[1]),.dout(n3743),.clk(gclk));
	jand g3102(.dina(w_n1556_36[1]),.dinb(w_in281_0[0]),.dout(n3744),.clk(gclk));
	jand g3103(.dina(w_n1711_37[0]),.dinb(w_in381_0[0]),.dout(n3745),.clk(gclk));
	jor g3104(.dina(n3745),.dinb(n3744),.dout(n3746),.clk(gclk));
	jand g3105(.dina(w_n3746_0[2]),.dinb(w_n3743_0[1]),.dout(n3747),.clk(gclk));
	jand g3106(.dina(w_n1556_36[0]),.dinb(w_in280_0[0]),.dout(n3748),.clk(gclk));
	jand g3107(.dina(w_n1711_36[2]),.dinb(w_in380_0[0]),.dout(n3749),.clk(gclk));
	jor g3108(.dina(n3749),.dinb(n3748),.dout(n3750),.clk(gclk));
	jand g3109(.dina(w_n2628_36[2]),.dinb(w_in080_0[0]),.dout(n3751),.clk(gclk));
	jand g3110(.dina(w_n2783_37[0]),.dinb(w_in180_0[0]),.dout(n3752),.clk(gclk));
	jor g3111(.dina(n3752),.dinb(n3751),.dout(n3753),.clk(gclk));
	jnot g3112(.din(w_n3753_0[1]),.dout(n3754),.clk(gclk));
	jand g3113(.dina(w_n3754_0[1]),.dinb(w_n3750_0[2]),.dout(n3755),.clk(gclk));
	jor g3114(.dina(n3755),.dinb(w_n3747_0[1]),.dout(n3756),.clk(gclk));
	jor g3115(.dina(n3756),.dinb(w_n3739_0[1]),.dout(n3757),.clk(gclk));
	jor g3116(.dina(w_n3757_0[1]),.dinb(n3722),.dout(n3758),.clk(gclk));
	jor g3117(.dina(w_n3729_0[1]),.dinb(w_n3726_0[0]),.dout(n3759),.clk(gclk));
	jor g3118(.dina(w_n3754_0[0]),.dinb(w_n3750_0[1]),.dout(n3760),.clk(gclk));
	jor g3119(.dina(n3760),.dinb(w_n3747_0[0]),.dout(n3761),.clk(gclk));
	jor g3120(.dina(w_n3746_0[1]),.dinb(w_n3743_0[0]),.dout(n3762),.clk(gclk));
	jor g3121(.dina(w_n3737_0[0]),.dinb(w_n3733_0[1]),.dout(n3763),.clk(gclk));
	jand g3122(.dina(n3763),.dinb(n3762),.dout(n3764),.clk(gclk));
	jand g3123(.dina(n3764),.dinb(n3761),.dout(n3765),.clk(gclk));
	jor g3124(.dina(n3765),.dinb(w_n3739_0[0]),.dout(n3766),.clk(gclk));
	jand g3125(.dina(n3766),.dinb(n3759),.dout(n3767),.clk(gclk));
	jand g3126(.dina(w_n3767_0[1]),.dinb(n3758),.dout(n3768),.clk(gclk));
	jand g3127(.dina(w_n2628_36[1]),.dinb(w_in084_0[0]),.dout(n3769),.clk(gclk));
	jand g3128(.dina(w_n2783_36[2]),.dinb(w_in184_0[0]),.dout(n3770),.clk(gclk));
	jor g3129(.dina(n3770),.dinb(n3769),.dout(n3771),.clk(gclk));
	jnot g3130(.din(w_n3771_0[1]),.dout(n3772),.clk(gclk));
	jand g3131(.dina(w_n1556_35[2]),.dinb(w_in284_0[0]),.dout(n3773),.clk(gclk));
	jand g3132(.dina(w_n1711_36[1]),.dinb(w_in384_0[0]),.dout(n3774),.clk(gclk));
	jor g3133(.dina(n3774),.dinb(n3773),.dout(n3775),.clk(gclk));
	jand g3134(.dina(w_n3775_0[2]),.dinb(w_n3772_0[1]),.dout(n3776),.clk(gclk));
	jand g3135(.dina(w_n2628_36[0]),.dinb(w_in085_0[0]),.dout(n3777),.clk(gclk));
	jand g3136(.dina(w_n2783_36[1]),.dinb(w_in185_0[0]),.dout(n3778),.clk(gclk));
	jor g3137(.dina(n3778),.dinb(n3777),.dout(n3779),.clk(gclk));
	jnot g3138(.din(w_n3779_0[1]),.dout(n3780),.clk(gclk));
	jand g3139(.dina(w_n1556_35[1]),.dinb(w_in285_0[0]),.dout(n3781),.clk(gclk));
	jand g3140(.dina(w_n1711_36[0]),.dinb(w_in385_0[0]),.dout(n3782),.clk(gclk));
	jor g3141(.dina(n3782),.dinb(n3781),.dout(n3783),.clk(gclk));
	jand g3142(.dina(w_n3783_0[2]),.dinb(w_n3780_0[1]),.dout(n3784),.clk(gclk));
	jand g3143(.dina(w_n2628_35[2]),.dinb(w_in087_0[0]),.dout(n3785),.clk(gclk));
	jand g3144(.dina(w_n2783_36[0]),.dinb(w_in187_0[0]),.dout(n3786),.clk(gclk));
	jor g3145(.dina(n3786),.dinb(n3785),.dout(n3787),.clk(gclk));
	jnot g3146(.din(w_n3787_0[1]),.dout(n3788),.clk(gclk));
	jand g3147(.dina(w_n1556_35[0]),.dinb(w_in287_0[0]),.dout(n3789),.clk(gclk));
	jand g3148(.dina(w_n1711_35[2]),.dinb(w_in387_0[0]),.dout(n3790),.clk(gclk));
	jor g3149(.dina(n3790),.dinb(n3789),.dout(n3791),.clk(gclk));
	jand g3150(.dina(w_n3791_0[2]),.dinb(w_n3788_0[1]),.dout(n3792),.clk(gclk));
	jand g3151(.dina(w_n1556_34[2]),.dinb(w_in286_0[0]),.dout(n3793),.clk(gclk));
	jand g3152(.dina(w_n1711_35[1]),.dinb(w_in386_0[0]),.dout(n3794),.clk(gclk));
	jor g3153(.dina(n3794),.dinb(n3793),.dout(n3795),.clk(gclk));
	jand g3154(.dina(w_n2628_35[1]),.dinb(w_in086_0[0]),.dout(n3796),.clk(gclk));
	jand g3155(.dina(w_n2783_35[2]),.dinb(w_in186_0[0]),.dout(n3797),.clk(gclk));
	jor g3156(.dina(n3797),.dinb(n3796),.dout(n3798),.clk(gclk));
	jnot g3157(.din(w_n3798_0[1]),.dout(n3799),.clk(gclk));
	jand g3158(.dina(w_n3799_0[1]),.dinb(w_n3795_0[2]),.dout(n3800),.clk(gclk));
	jor g3159(.dina(n3800),.dinb(w_n3792_0[1]),.dout(n3801),.clk(gclk));
	jor g3160(.dina(n3801),.dinb(n3784),.dout(n3802),.clk(gclk));
	jor g3161(.dina(w_n3802_0[1]),.dinb(n3776),.dout(n3803),.clk(gclk));
	jor g3162(.dina(w_n3803_0[1]),.dinb(n3768),.dout(n3804),.clk(gclk));
	jor g3163(.dina(w_n3783_0[1]),.dinb(w_n3780_0[0]),.dout(n3805),.clk(gclk));
	jor g3164(.dina(w_n3775_0[1]),.dinb(w_n3772_0[0]),.dout(n3806),.clk(gclk));
	jand g3165(.dina(n3806),.dinb(n3805),.dout(n3807),.clk(gclk));
	jor g3166(.dina(n3807),.dinb(w_n3802_0[0]),.dout(n3808),.clk(gclk));
	jor g3167(.dina(w_n3791_0[1]),.dinb(w_n3788_0[0]),.dout(n3809),.clk(gclk));
	jor g3168(.dina(w_n3799_0[0]),.dinb(w_n3795_0[1]),.dout(n3810),.clk(gclk));
	jor g3169(.dina(n3810),.dinb(w_n3792_0[0]),.dout(n3811),.clk(gclk));
	jand g3170(.dina(n3811),.dinb(n3809),.dout(n3812),.clk(gclk));
	jand g3171(.dina(n3812),.dinb(n3808),.dout(n3813),.clk(gclk));
	jand g3172(.dina(w_n3813_0[1]),.dinb(n3804),.dout(n3814),.clk(gclk));
	jand g3173(.dina(w_n2628_35[0]),.dinb(w_in091_0[0]),.dout(n3815),.clk(gclk));
	jand g3174(.dina(w_n2783_35[1]),.dinb(w_in191_0[0]),.dout(n3816),.clk(gclk));
	jor g3175(.dina(n3816),.dinb(n3815),.dout(n3817),.clk(gclk));
	jnot g3176(.din(w_n3817_0[1]),.dout(n3818),.clk(gclk));
	jand g3177(.dina(w_n1556_34[1]),.dinb(w_in291_0[0]),.dout(n3819),.clk(gclk));
	jand g3178(.dina(w_n1711_35[0]),.dinb(w_in391_0[0]),.dout(n3820),.clk(gclk));
	jor g3179(.dina(n3820),.dinb(n3819),.dout(n3821),.clk(gclk));
	jand g3180(.dina(w_n3821_0[2]),.dinb(w_n3818_0[1]),.dout(n3822),.clk(gclk));
	jand g3181(.dina(w_n1556_34[0]),.dinb(w_in290_0[0]),.dout(n3823),.clk(gclk));
	jand g3182(.dina(w_n1711_34[2]),.dinb(w_in390_0[0]),.dout(n3824),.clk(gclk));
	jor g3183(.dina(n3824),.dinb(n3823),.dout(n3825),.clk(gclk));
	jand g3184(.dina(w_n2628_34[2]),.dinb(w_in090_0[0]),.dout(n3826),.clk(gclk));
	jand g3185(.dina(w_n2783_35[0]),.dinb(w_in190_0[0]),.dout(n3827),.clk(gclk));
	jor g3186(.dina(n3827),.dinb(n3826),.dout(n3828),.clk(gclk));
	jnot g3187(.din(w_n3828_0[1]),.dout(n3829),.clk(gclk));
	jand g3188(.dina(w_n3829_0[1]),.dinb(w_n3825_0[2]),.dout(n3830),.clk(gclk));
	jor g3189(.dina(n3830),.dinb(n3822),.dout(n3831),.clk(gclk));
	jand g3190(.dina(w_n2628_34[1]),.dinb(w_in089_0[0]),.dout(n3832),.clk(gclk));
	jand g3191(.dina(w_n2783_34[2]),.dinb(w_in189_0[0]),.dout(n3833),.clk(gclk));
	jor g3192(.dina(n3833),.dinb(n3832),.dout(n3834),.clk(gclk));
	jnot g3193(.din(w_n3834_0[1]),.dout(n3835),.clk(gclk));
	jand g3194(.dina(w_n1556_33[2]),.dinb(w_in289_0[0]),.dout(n3836),.clk(gclk));
	jand g3195(.dina(w_n1711_34[1]),.dinb(w_in389_0[0]),.dout(n3837),.clk(gclk));
	jor g3196(.dina(n3837),.dinb(n3836),.dout(n3838),.clk(gclk));
	jand g3197(.dina(w_n3838_0[2]),.dinb(w_n3835_0[1]),.dout(n3839),.clk(gclk));
	jand g3198(.dina(w_n1556_33[1]),.dinb(w_in288_0[0]),.dout(n3840),.clk(gclk));
	jand g3199(.dina(w_n1711_34[0]),.dinb(w_in388_0[0]),.dout(n3841),.clk(gclk));
	jor g3200(.dina(n3841),.dinb(n3840),.dout(n3842),.clk(gclk));
	jand g3201(.dina(w_n2628_34[0]),.dinb(w_in088_0[0]),.dout(n3843),.clk(gclk));
	jand g3202(.dina(w_n2783_34[1]),.dinb(w_in188_0[0]),.dout(n3844),.clk(gclk));
	jor g3203(.dina(n3844),.dinb(n3843),.dout(n3845),.clk(gclk));
	jnot g3204(.din(w_n3845_0[1]),.dout(n3846),.clk(gclk));
	jand g3205(.dina(w_n3846_0[1]),.dinb(w_n3842_0[2]),.dout(n3847),.clk(gclk));
	jor g3206(.dina(n3847),.dinb(w_n3839_0[1]),.dout(n3848),.clk(gclk));
	jor g3207(.dina(n3848),.dinb(w_n3831_0[1]),.dout(n3849),.clk(gclk));
	jor g3208(.dina(w_n3849_0[1]),.dinb(n3814),.dout(n3850),.clk(gclk));
	jor g3209(.dina(w_n3821_0[1]),.dinb(w_n3818_0[0]),.dout(n3851),.clk(gclk));
	jor g3210(.dina(w_n3846_0[0]),.dinb(w_n3842_0[1]),.dout(n3852),.clk(gclk));
	jor g3211(.dina(n3852),.dinb(w_n3839_0[0]),.dout(n3853),.clk(gclk));
	jor g3212(.dina(w_n3838_0[1]),.dinb(w_n3835_0[0]),.dout(n3854),.clk(gclk));
	jor g3213(.dina(w_n3829_0[0]),.dinb(w_n3825_0[1]),.dout(n3855),.clk(gclk));
	jand g3214(.dina(n3855),.dinb(n3854),.dout(n3856),.clk(gclk));
	jand g3215(.dina(n3856),.dinb(n3853),.dout(n3857),.clk(gclk));
	jor g3216(.dina(n3857),.dinb(w_n3831_0[0]),.dout(n3858),.clk(gclk));
	jand g3217(.dina(n3858),.dinb(n3851),.dout(n3859),.clk(gclk));
	jand g3218(.dina(w_n3859_0[1]),.dinb(n3850),.dout(n3860),.clk(gclk));
	jand g3219(.dina(w_n2628_33[2]),.dinb(w_in092_0[0]),.dout(n3861),.clk(gclk));
	jand g3220(.dina(w_n2783_34[0]),.dinb(w_in192_0[0]),.dout(n3862),.clk(gclk));
	jor g3221(.dina(n3862),.dinb(n3861),.dout(n3863),.clk(gclk));
	jnot g3222(.din(w_n3863_0[1]),.dout(n3864),.clk(gclk));
	jand g3223(.dina(w_n1556_33[0]),.dinb(w_in292_0[0]),.dout(n3865),.clk(gclk));
	jand g3224(.dina(w_n1711_33[2]),.dinb(w_in392_0[0]),.dout(n3866),.clk(gclk));
	jor g3225(.dina(n3866),.dinb(n3865),.dout(n3867),.clk(gclk));
	jand g3226(.dina(w_n3867_0[2]),.dinb(w_n3864_0[1]),.dout(n3868),.clk(gclk));
	jand g3227(.dina(w_n2628_33[1]),.dinb(w_in093_0[0]),.dout(n3869),.clk(gclk));
	jand g3228(.dina(w_n2783_33[2]),.dinb(w_in193_0[0]),.dout(n3870),.clk(gclk));
	jor g3229(.dina(n3870),.dinb(n3869),.dout(n3871),.clk(gclk));
	jnot g3230(.din(w_n3871_0[1]),.dout(n3872),.clk(gclk));
	jand g3231(.dina(w_n1556_32[2]),.dinb(w_in293_0[0]),.dout(n3873),.clk(gclk));
	jand g3232(.dina(w_n1711_33[1]),.dinb(w_in393_0[0]),.dout(n3874),.clk(gclk));
	jor g3233(.dina(n3874),.dinb(n3873),.dout(n3875),.clk(gclk));
	jand g3234(.dina(w_n3875_0[2]),.dinb(w_n3872_0[1]),.dout(n3876),.clk(gclk));
	jand g3235(.dina(w_n2628_33[0]),.dinb(w_in095_0[0]),.dout(n3877),.clk(gclk));
	jand g3236(.dina(w_n2783_33[1]),.dinb(w_in195_0[0]),.dout(n3878),.clk(gclk));
	jor g3237(.dina(n3878),.dinb(n3877),.dout(n3879),.clk(gclk));
	jnot g3238(.din(w_n3879_0[1]),.dout(n3880),.clk(gclk));
	jand g3239(.dina(w_n1556_32[1]),.dinb(w_in295_0[0]),.dout(n3881),.clk(gclk));
	jand g3240(.dina(w_n1711_33[0]),.dinb(w_in395_0[0]),.dout(n3882),.clk(gclk));
	jor g3241(.dina(n3882),.dinb(n3881),.dout(n3883),.clk(gclk));
	jand g3242(.dina(w_n3883_0[2]),.dinb(w_n3880_0[1]),.dout(n3884),.clk(gclk));
	jand g3243(.dina(w_n1556_32[0]),.dinb(w_in294_0[0]),.dout(n3885),.clk(gclk));
	jand g3244(.dina(w_n1711_32[2]),.dinb(w_in394_0[0]),.dout(n3886),.clk(gclk));
	jor g3245(.dina(n3886),.dinb(n3885),.dout(n3887),.clk(gclk));
	jand g3246(.dina(w_n2628_32[2]),.dinb(w_in094_0[0]),.dout(n3888),.clk(gclk));
	jand g3247(.dina(w_n2783_33[0]),.dinb(w_in194_0[0]),.dout(n3889),.clk(gclk));
	jor g3248(.dina(n3889),.dinb(n3888),.dout(n3890),.clk(gclk));
	jnot g3249(.din(w_n3890_0[1]),.dout(n3891),.clk(gclk));
	jand g3250(.dina(w_n3891_0[1]),.dinb(w_n3887_0[2]),.dout(n3892),.clk(gclk));
	jor g3251(.dina(n3892),.dinb(w_n3884_0[1]),.dout(n3893),.clk(gclk));
	jor g3252(.dina(n3893),.dinb(n3876),.dout(n3894),.clk(gclk));
	jor g3253(.dina(w_n3894_0[1]),.dinb(n3868),.dout(n3895),.clk(gclk));
	jor g3254(.dina(w_n3895_0[1]),.dinb(n3860),.dout(n3896),.clk(gclk));
	jor g3255(.dina(w_n3875_0[1]),.dinb(w_n3872_0[0]),.dout(n3897),.clk(gclk));
	jor g3256(.dina(w_n3867_0[1]),.dinb(w_n3864_0[0]),.dout(n3898),.clk(gclk));
	jand g3257(.dina(n3898),.dinb(n3897),.dout(n3899),.clk(gclk));
	jor g3258(.dina(n3899),.dinb(w_n3894_0[0]),.dout(n3900),.clk(gclk));
	jor g3259(.dina(w_n3883_0[1]),.dinb(w_n3880_0[0]),.dout(n3901),.clk(gclk));
	jor g3260(.dina(w_n3891_0[0]),.dinb(w_n3887_0[1]),.dout(n3902),.clk(gclk));
	jor g3261(.dina(n3902),.dinb(w_n3884_0[0]),.dout(n3903),.clk(gclk));
	jand g3262(.dina(n3903),.dinb(n3901),.dout(n3904),.clk(gclk));
	jand g3263(.dina(n3904),.dinb(n3900),.dout(n3905),.clk(gclk));
	jand g3264(.dina(w_n3905_0[1]),.dinb(n3896),.dout(n3906),.clk(gclk));
	jand g3265(.dina(w_n2628_32[1]),.dinb(w_in099_0[0]),.dout(n3907),.clk(gclk));
	jand g3266(.dina(w_n2783_32[2]),.dinb(w_in199_0[0]),.dout(n3908),.clk(gclk));
	jor g3267(.dina(n3908),.dinb(n3907),.dout(n3909),.clk(gclk));
	jnot g3268(.din(w_n3909_0[1]),.dout(n3910),.clk(gclk));
	jand g3269(.dina(w_n1556_31[2]),.dinb(w_in299_0[0]),.dout(n3911),.clk(gclk));
	jand g3270(.dina(w_n1711_32[1]),.dinb(w_in399_0[0]),.dout(n3912),.clk(gclk));
	jor g3271(.dina(n3912),.dinb(n3911),.dout(n3913),.clk(gclk));
	jand g3272(.dina(w_n3913_0[2]),.dinb(w_n3910_0[1]),.dout(n3914),.clk(gclk));
	jand g3273(.dina(w_n1556_31[1]),.dinb(w_in298_0[0]),.dout(n3915),.clk(gclk));
	jand g3274(.dina(w_n1711_32[0]),.dinb(w_in398_0[0]),.dout(n3916),.clk(gclk));
	jor g3275(.dina(n3916),.dinb(n3915),.dout(n3917),.clk(gclk));
	jand g3276(.dina(w_n2628_32[0]),.dinb(w_in098_0[0]),.dout(n3918),.clk(gclk));
	jand g3277(.dina(w_n2783_32[1]),.dinb(w_in198_0[0]),.dout(n3919),.clk(gclk));
	jor g3278(.dina(n3919),.dinb(n3918),.dout(n3920),.clk(gclk));
	jnot g3279(.din(w_n3920_0[1]),.dout(n3921),.clk(gclk));
	jand g3280(.dina(w_n3921_0[1]),.dinb(w_n3917_0[2]),.dout(n3922),.clk(gclk));
	jor g3281(.dina(n3922),.dinb(n3914),.dout(n3923),.clk(gclk));
	jand g3282(.dina(w_n2628_31[2]),.dinb(w_in097_0[0]),.dout(n3924),.clk(gclk));
	jand g3283(.dina(w_n2783_32[0]),.dinb(w_in197_0[0]),.dout(n3925),.clk(gclk));
	jor g3284(.dina(n3925),.dinb(n3924),.dout(n3926),.clk(gclk));
	jnot g3285(.din(w_n3926_0[1]),.dout(n3927),.clk(gclk));
	jand g3286(.dina(w_n1556_31[0]),.dinb(w_in297_0[0]),.dout(n3928),.clk(gclk));
	jand g3287(.dina(w_n1711_31[2]),.dinb(w_in397_0[0]),.dout(n3929),.clk(gclk));
	jor g3288(.dina(n3929),.dinb(n3928),.dout(n3930),.clk(gclk));
	jand g3289(.dina(w_n3930_0[2]),.dinb(w_n3927_0[1]),.dout(n3931),.clk(gclk));
	jand g3290(.dina(w_n1556_30[2]),.dinb(w_in296_0[0]),.dout(n3932),.clk(gclk));
	jand g3291(.dina(w_n1711_31[1]),.dinb(w_in396_0[0]),.dout(n3933),.clk(gclk));
	jor g3292(.dina(n3933),.dinb(n3932),.dout(n3934),.clk(gclk));
	jand g3293(.dina(w_n2628_31[1]),.dinb(w_in096_0[0]),.dout(n3935),.clk(gclk));
	jand g3294(.dina(w_n2783_31[2]),.dinb(w_in196_0[0]),.dout(n3936),.clk(gclk));
	jor g3295(.dina(n3936),.dinb(n3935),.dout(n3937),.clk(gclk));
	jnot g3296(.din(w_n3937_0[1]),.dout(n3938),.clk(gclk));
	jand g3297(.dina(w_n3938_0[1]),.dinb(w_n3934_0[2]),.dout(n3939),.clk(gclk));
	jor g3298(.dina(n3939),.dinb(w_n3931_0[1]),.dout(n3940),.clk(gclk));
	jor g3299(.dina(n3940),.dinb(w_n3923_0[1]),.dout(n3941),.clk(gclk));
	jor g3300(.dina(w_n3941_0[1]),.dinb(n3906),.dout(n3942),.clk(gclk));
	jor g3301(.dina(w_n3913_0[1]),.dinb(w_n3910_0[0]),.dout(n3943),.clk(gclk));
	jor g3302(.dina(w_n3938_0[0]),.dinb(w_n3934_0[1]),.dout(n3944),.clk(gclk));
	jor g3303(.dina(n3944),.dinb(w_n3931_0[0]),.dout(n3945),.clk(gclk));
	jor g3304(.dina(w_n3930_0[1]),.dinb(w_n3927_0[0]),.dout(n3946),.clk(gclk));
	jor g3305(.dina(w_n3921_0[0]),.dinb(w_n3917_0[1]),.dout(n3947),.clk(gclk));
	jand g3306(.dina(n3947),.dinb(n3946),.dout(n3948),.clk(gclk));
	jand g3307(.dina(n3948),.dinb(n3945),.dout(n3949),.clk(gclk));
	jor g3308(.dina(n3949),.dinb(w_n3923_0[0]),.dout(n3950),.clk(gclk));
	jand g3309(.dina(n3950),.dinb(n3943),.dout(n3951),.clk(gclk));
	jand g3310(.dina(w_n3951_0[1]),.dinb(n3942),.dout(n3952),.clk(gclk));
	jand g3311(.dina(w_n2628_31[0]),.dinb(w_in0100_0[0]),.dout(n3953),.clk(gclk));
	jand g3312(.dina(w_n2783_31[1]),.dinb(w_in1100_0[0]),.dout(n3954),.clk(gclk));
	jor g3313(.dina(n3954),.dinb(n3953),.dout(n3955),.clk(gclk));
	jnot g3314(.din(w_n3955_0[1]),.dout(n3956),.clk(gclk));
	jand g3315(.dina(w_n1556_30[1]),.dinb(w_in2100_0[0]),.dout(n3957),.clk(gclk));
	jand g3316(.dina(w_n1711_31[0]),.dinb(w_in3100_0[0]),.dout(n3958),.clk(gclk));
	jor g3317(.dina(n3958),.dinb(n3957),.dout(n3959),.clk(gclk));
	jand g3318(.dina(w_n3959_0[2]),.dinb(w_n3956_0[1]),.dout(n3960),.clk(gclk));
	jand g3319(.dina(w_n2628_30[2]),.dinb(w_in0101_0[0]),.dout(n3961),.clk(gclk));
	jand g3320(.dina(w_n2783_31[0]),.dinb(w_in1101_0[0]),.dout(n3962),.clk(gclk));
	jor g3321(.dina(n3962),.dinb(n3961),.dout(n3963),.clk(gclk));
	jnot g3322(.din(w_n3963_0[1]),.dout(n3964),.clk(gclk));
	jand g3323(.dina(w_n1556_30[0]),.dinb(w_in2101_0[0]),.dout(n3965),.clk(gclk));
	jand g3324(.dina(w_n1711_30[2]),.dinb(w_in3101_0[0]),.dout(n3966),.clk(gclk));
	jor g3325(.dina(n3966),.dinb(n3965),.dout(n3967),.clk(gclk));
	jand g3326(.dina(w_n3967_0[2]),.dinb(w_n3964_0[1]),.dout(n3968),.clk(gclk));
	jand g3327(.dina(w_n2628_30[1]),.dinb(w_in0103_0[0]),.dout(n3969),.clk(gclk));
	jand g3328(.dina(w_n2783_30[2]),.dinb(w_in1103_0[0]),.dout(n3970),.clk(gclk));
	jor g3329(.dina(n3970),.dinb(n3969),.dout(n3971),.clk(gclk));
	jnot g3330(.din(w_n3971_0[1]),.dout(n3972),.clk(gclk));
	jand g3331(.dina(w_n1556_29[2]),.dinb(w_in2103_0[0]),.dout(n3973),.clk(gclk));
	jand g3332(.dina(w_n1711_30[1]),.dinb(w_in3103_0[0]),.dout(n3974),.clk(gclk));
	jor g3333(.dina(n3974),.dinb(n3973),.dout(n3975),.clk(gclk));
	jand g3334(.dina(w_n3975_0[2]),.dinb(w_n3972_0[1]),.dout(n3976),.clk(gclk));
	jand g3335(.dina(w_n1556_29[1]),.dinb(w_in2102_0[0]),.dout(n3977),.clk(gclk));
	jand g3336(.dina(w_n1711_30[0]),.dinb(w_in3102_0[0]),.dout(n3978),.clk(gclk));
	jor g3337(.dina(n3978),.dinb(n3977),.dout(n3979),.clk(gclk));
	jand g3338(.dina(w_n2628_30[0]),.dinb(w_in0102_0[0]),.dout(n3980),.clk(gclk));
	jand g3339(.dina(w_n2783_30[1]),.dinb(w_in1102_0[0]),.dout(n3981),.clk(gclk));
	jor g3340(.dina(n3981),.dinb(n3980),.dout(n3982),.clk(gclk));
	jnot g3341(.din(w_n3982_0[1]),.dout(n3983),.clk(gclk));
	jand g3342(.dina(w_n3983_0[1]),.dinb(w_n3979_0[2]),.dout(n3984),.clk(gclk));
	jor g3343(.dina(n3984),.dinb(w_n3976_0[1]),.dout(n3985),.clk(gclk));
	jor g3344(.dina(n3985),.dinb(n3968),.dout(n3986),.clk(gclk));
	jor g3345(.dina(w_n3986_0[1]),.dinb(n3960),.dout(n3987),.clk(gclk));
	jor g3346(.dina(w_n3987_0[1]),.dinb(n3952),.dout(n3988),.clk(gclk));
	jor g3347(.dina(w_n3967_0[1]),.dinb(w_n3964_0[0]),.dout(n3989),.clk(gclk));
	jor g3348(.dina(w_n3959_0[1]),.dinb(w_n3956_0[0]),.dout(n3990),.clk(gclk));
	jand g3349(.dina(n3990),.dinb(n3989),.dout(n3991),.clk(gclk));
	jor g3350(.dina(n3991),.dinb(w_n3986_0[0]),.dout(n3992),.clk(gclk));
	jor g3351(.dina(w_n3975_0[1]),.dinb(w_n3972_0[0]),.dout(n3993),.clk(gclk));
	jor g3352(.dina(w_n3983_0[0]),.dinb(w_n3979_0[1]),.dout(n3994),.clk(gclk));
	jor g3353(.dina(n3994),.dinb(w_n3976_0[0]),.dout(n3995),.clk(gclk));
	jand g3354(.dina(n3995),.dinb(n3993),.dout(n3996),.clk(gclk));
	jand g3355(.dina(n3996),.dinb(n3992),.dout(n3997),.clk(gclk));
	jand g3356(.dina(w_n3997_0[1]),.dinb(n3988),.dout(n3998),.clk(gclk));
	jand g3357(.dina(w_n2628_29[2]),.dinb(w_in0107_0[0]),.dout(n3999),.clk(gclk));
	jand g3358(.dina(w_n2783_30[0]),.dinb(w_in1107_0[0]),.dout(n4000),.clk(gclk));
	jor g3359(.dina(n4000),.dinb(n3999),.dout(n4001),.clk(gclk));
	jnot g3360(.din(w_n4001_0[1]),.dout(n4002),.clk(gclk));
	jand g3361(.dina(w_n1556_29[0]),.dinb(w_in2107_0[0]),.dout(n4003),.clk(gclk));
	jand g3362(.dina(w_n1711_29[2]),.dinb(w_in3107_0[0]),.dout(n4004),.clk(gclk));
	jor g3363(.dina(n4004),.dinb(n4003),.dout(n4005),.clk(gclk));
	jand g3364(.dina(w_n4005_0[2]),.dinb(w_n4002_0[1]),.dout(n4006),.clk(gclk));
	jand g3365(.dina(w_n1556_28[2]),.dinb(w_in2106_0[0]),.dout(n4007),.clk(gclk));
	jand g3366(.dina(w_n1711_29[1]),.dinb(w_in3106_0[0]),.dout(n4008),.clk(gclk));
	jor g3367(.dina(n4008),.dinb(n4007),.dout(n4009),.clk(gclk));
	jand g3368(.dina(w_n2628_29[1]),.dinb(w_in0106_0[0]),.dout(n4010),.clk(gclk));
	jand g3369(.dina(w_n2783_29[2]),.dinb(w_in1106_0[0]),.dout(n4011),.clk(gclk));
	jor g3370(.dina(n4011),.dinb(n4010),.dout(n4012),.clk(gclk));
	jnot g3371(.din(w_n4012_0[1]),.dout(n4013),.clk(gclk));
	jand g3372(.dina(w_n4013_0[1]),.dinb(w_n4009_0[2]),.dout(n4014),.clk(gclk));
	jor g3373(.dina(n4014),.dinb(n4006),.dout(n4015),.clk(gclk));
	jand g3374(.dina(w_n2628_29[0]),.dinb(w_in0105_0[0]),.dout(n4016),.clk(gclk));
	jand g3375(.dina(w_n2783_29[1]),.dinb(w_in1105_0[0]),.dout(n4017),.clk(gclk));
	jor g3376(.dina(n4017),.dinb(n4016),.dout(n4018),.clk(gclk));
	jnot g3377(.din(w_n4018_0[1]),.dout(n4019),.clk(gclk));
	jand g3378(.dina(w_n1556_28[1]),.dinb(w_in2105_0[0]),.dout(n4020),.clk(gclk));
	jand g3379(.dina(w_n1711_29[0]),.dinb(w_in3105_0[0]),.dout(n4021),.clk(gclk));
	jor g3380(.dina(n4021),.dinb(n4020),.dout(n4022),.clk(gclk));
	jand g3381(.dina(w_n4022_0[2]),.dinb(w_n4019_0[1]),.dout(n4023),.clk(gclk));
	jand g3382(.dina(w_n1556_28[0]),.dinb(w_in2104_0[0]),.dout(n4024),.clk(gclk));
	jand g3383(.dina(w_n1711_28[2]),.dinb(w_in3104_0[0]),.dout(n4025),.clk(gclk));
	jor g3384(.dina(n4025),.dinb(n4024),.dout(n4026),.clk(gclk));
	jand g3385(.dina(w_n2628_28[2]),.dinb(w_in0104_0[0]),.dout(n4027),.clk(gclk));
	jand g3386(.dina(w_n2783_29[0]),.dinb(w_in1104_0[0]),.dout(n4028),.clk(gclk));
	jor g3387(.dina(n4028),.dinb(n4027),.dout(n4029),.clk(gclk));
	jnot g3388(.din(w_n4029_0[1]),.dout(n4030),.clk(gclk));
	jand g3389(.dina(w_n4030_0[1]),.dinb(w_n4026_0[2]),.dout(n4031),.clk(gclk));
	jor g3390(.dina(n4031),.dinb(w_n4023_0[1]),.dout(n4032),.clk(gclk));
	jor g3391(.dina(n4032),.dinb(w_n4015_0[1]),.dout(n4033),.clk(gclk));
	jor g3392(.dina(w_n4033_0[1]),.dinb(n3998),.dout(n4034),.clk(gclk));
	jor g3393(.dina(w_n4005_0[1]),.dinb(w_n4002_0[0]),.dout(n4035),.clk(gclk));
	jor g3394(.dina(w_n4030_0[0]),.dinb(w_n4026_0[1]),.dout(n4036),.clk(gclk));
	jor g3395(.dina(n4036),.dinb(w_n4023_0[0]),.dout(n4037),.clk(gclk));
	jor g3396(.dina(w_n4022_0[1]),.dinb(w_n4019_0[0]),.dout(n4038),.clk(gclk));
	jor g3397(.dina(w_n4013_0[0]),.dinb(w_n4009_0[1]),.dout(n4039),.clk(gclk));
	jand g3398(.dina(n4039),.dinb(n4038),.dout(n4040),.clk(gclk));
	jand g3399(.dina(n4040),.dinb(n4037),.dout(n4041),.clk(gclk));
	jor g3400(.dina(n4041),.dinb(w_n4015_0[0]),.dout(n4042),.clk(gclk));
	jand g3401(.dina(n4042),.dinb(n4035),.dout(n4043),.clk(gclk));
	jand g3402(.dina(w_n4043_0[1]),.dinb(n4034),.dout(n4044),.clk(gclk));
	jand g3403(.dina(w_n2628_28[1]),.dinb(w_in0108_0[0]),.dout(n4045),.clk(gclk));
	jand g3404(.dina(w_n2783_28[2]),.dinb(w_in1108_0[0]),.dout(n4046),.clk(gclk));
	jor g3405(.dina(n4046),.dinb(n4045),.dout(n4047),.clk(gclk));
	jnot g3406(.din(w_n4047_0[1]),.dout(n4048),.clk(gclk));
	jand g3407(.dina(w_n1556_27[2]),.dinb(w_in2108_0[0]),.dout(n4049),.clk(gclk));
	jand g3408(.dina(w_n1711_28[1]),.dinb(w_in3108_0[0]),.dout(n4050),.clk(gclk));
	jor g3409(.dina(n4050),.dinb(n4049),.dout(n4051),.clk(gclk));
	jand g3410(.dina(w_n4051_0[2]),.dinb(w_n4048_0[1]),.dout(n4052),.clk(gclk));
	jand g3411(.dina(w_n2628_28[0]),.dinb(w_in0109_0[0]),.dout(n4053),.clk(gclk));
	jand g3412(.dina(w_n2783_28[1]),.dinb(w_in1109_0[0]),.dout(n4054),.clk(gclk));
	jor g3413(.dina(n4054),.dinb(n4053),.dout(n4055),.clk(gclk));
	jnot g3414(.din(w_n4055_0[1]),.dout(n4056),.clk(gclk));
	jand g3415(.dina(w_n1556_27[1]),.dinb(w_in2109_0[0]),.dout(n4057),.clk(gclk));
	jand g3416(.dina(w_n1711_28[0]),.dinb(w_in3109_0[0]),.dout(n4058),.clk(gclk));
	jor g3417(.dina(n4058),.dinb(n4057),.dout(n4059),.clk(gclk));
	jand g3418(.dina(w_n4059_0[2]),.dinb(w_n4056_0[1]),.dout(n4060),.clk(gclk));
	jand g3419(.dina(w_n2628_27[2]),.dinb(w_in0111_0[0]),.dout(n4061),.clk(gclk));
	jand g3420(.dina(w_n2783_28[0]),.dinb(w_in1111_0[0]),.dout(n4062),.clk(gclk));
	jor g3421(.dina(n4062),.dinb(n4061),.dout(n4063),.clk(gclk));
	jnot g3422(.din(w_n4063_0[1]),.dout(n4064),.clk(gclk));
	jand g3423(.dina(w_n1556_27[0]),.dinb(w_in2111_0[0]),.dout(n4065),.clk(gclk));
	jand g3424(.dina(w_n1711_27[2]),.dinb(w_in3111_0[0]),.dout(n4066),.clk(gclk));
	jor g3425(.dina(n4066),.dinb(n4065),.dout(n4067),.clk(gclk));
	jand g3426(.dina(w_n4067_0[2]),.dinb(w_n4064_0[1]),.dout(n4068),.clk(gclk));
	jand g3427(.dina(w_n1556_26[2]),.dinb(w_in2110_0[0]),.dout(n4069),.clk(gclk));
	jand g3428(.dina(w_n1711_27[1]),.dinb(w_in3110_0[0]),.dout(n4070),.clk(gclk));
	jor g3429(.dina(n4070),.dinb(n4069),.dout(n4071),.clk(gclk));
	jand g3430(.dina(w_n2628_27[1]),.dinb(w_in0110_0[0]),.dout(n4072),.clk(gclk));
	jand g3431(.dina(w_n2783_27[2]),.dinb(w_in1110_0[0]),.dout(n4073),.clk(gclk));
	jor g3432(.dina(n4073),.dinb(n4072),.dout(n4074),.clk(gclk));
	jnot g3433(.din(w_n4074_0[1]),.dout(n4075),.clk(gclk));
	jand g3434(.dina(w_n4075_0[1]),.dinb(w_n4071_0[2]),.dout(n4076),.clk(gclk));
	jor g3435(.dina(n4076),.dinb(w_n4068_0[1]),.dout(n4077),.clk(gclk));
	jor g3436(.dina(n4077),.dinb(n4060),.dout(n4078),.clk(gclk));
	jor g3437(.dina(w_n4078_0[1]),.dinb(n4052),.dout(n4079),.clk(gclk));
	jor g3438(.dina(w_n4079_0[1]),.dinb(n4044),.dout(n4080),.clk(gclk));
	jor g3439(.dina(w_n4059_0[1]),.dinb(w_n4056_0[0]),.dout(n4081),.clk(gclk));
	jor g3440(.dina(w_n4051_0[1]),.dinb(w_n4048_0[0]),.dout(n4082),.clk(gclk));
	jand g3441(.dina(n4082),.dinb(n4081),.dout(n4083),.clk(gclk));
	jor g3442(.dina(n4083),.dinb(w_n4078_0[0]),.dout(n4084),.clk(gclk));
	jor g3443(.dina(w_n4067_0[1]),.dinb(w_n4064_0[0]),.dout(n4085),.clk(gclk));
	jor g3444(.dina(w_n4075_0[0]),.dinb(w_n4071_0[1]),.dout(n4086),.clk(gclk));
	jor g3445(.dina(n4086),.dinb(w_n4068_0[0]),.dout(n4087),.clk(gclk));
	jand g3446(.dina(n4087),.dinb(n4085),.dout(n4088),.clk(gclk));
	jand g3447(.dina(n4088),.dinb(n4084),.dout(n4089),.clk(gclk));
	jand g3448(.dina(w_n4089_0[1]),.dinb(n4080),.dout(n4090),.clk(gclk));
	jand g3449(.dina(w_n2628_27[0]),.dinb(w_in0115_0[0]),.dout(n4091),.clk(gclk));
	jand g3450(.dina(w_n2783_27[1]),.dinb(w_in1115_0[0]),.dout(n4092),.clk(gclk));
	jor g3451(.dina(n4092),.dinb(n4091),.dout(n4093),.clk(gclk));
	jnot g3452(.din(w_n4093_0[1]),.dout(n4094),.clk(gclk));
	jand g3453(.dina(w_n1556_26[1]),.dinb(w_in2115_0[0]),.dout(n4095),.clk(gclk));
	jand g3454(.dina(w_n1711_27[0]),.dinb(w_in3115_0[0]),.dout(n4096),.clk(gclk));
	jor g3455(.dina(n4096),.dinb(n4095),.dout(n4097),.clk(gclk));
	jand g3456(.dina(w_n4097_0[2]),.dinb(w_n4094_0[1]),.dout(n4098),.clk(gclk));
	jand g3457(.dina(w_n1556_26[0]),.dinb(w_in2114_0[0]),.dout(n4099),.clk(gclk));
	jand g3458(.dina(w_n1711_26[2]),.dinb(w_in3114_0[0]),.dout(n4100),.clk(gclk));
	jor g3459(.dina(n4100),.dinb(n4099),.dout(n4101),.clk(gclk));
	jand g3460(.dina(w_n2628_26[2]),.dinb(w_in0114_0[0]),.dout(n4102),.clk(gclk));
	jand g3461(.dina(w_n2783_27[0]),.dinb(w_in1114_0[0]),.dout(n4103),.clk(gclk));
	jor g3462(.dina(n4103),.dinb(n4102),.dout(n4104),.clk(gclk));
	jnot g3463(.din(w_n4104_0[1]),.dout(n4105),.clk(gclk));
	jand g3464(.dina(w_n4105_0[1]),.dinb(w_n4101_0[2]),.dout(n4106),.clk(gclk));
	jor g3465(.dina(n4106),.dinb(n4098),.dout(n4107),.clk(gclk));
	jand g3466(.dina(w_n2628_26[1]),.dinb(w_in0113_0[0]),.dout(n4108),.clk(gclk));
	jand g3467(.dina(w_n2783_26[2]),.dinb(w_in1113_0[0]),.dout(n4109),.clk(gclk));
	jor g3468(.dina(n4109),.dinb(n4108),.dout(n4110),.clk(gclk));
	jnot g3469(.din(w_n4110_0[1]),.dout(n4111),.clk(gclk));
	jand g3470(.dina(w_n1556_25[2]),.dinb(w_in2113_0[0]),.dout(n4112),.clk(gclk));
	jand g3471(.dina(w_n1711_26[1]),.dinb(w_in3113_0[0]),.dout(n4113),.clk(gclk));
	jor g3472(.dina(n4113),.dinb(n4112),.dout(n4114),.clk(gclk));
	jand g3473(.dina(w_n4114_0[2]),.dinb(w_n4111_0[1]),.dout(n4115),.clk(gclk));
	jand g3474(.dina(w_n1556_25[1]),.dinb(w_in2112_0[0]),.dout(n4116),.clk(gclk));
	jand g3475(.dina(w_n1711_26[0]),.dinb(w_in3112_0[0]),.dout(n4117),.clk(gclk));
	jor g3476(.dina(n4117),.dinb(n4116),.dout(n4118),.clk(gclk));
	jand g3477(.dina(w_n2628_26[0]),.dinb(w_in0112_0[0]),.dout(n4119),.clk(gclk));
	jand g3478(.dina(w_n2783_26[1]),.dinb(w_in1112_0[0]),.dout(n4120),.clk(gclk));
	jor g3479(.dina(n4120),.dinb(n4119),.dout(n4121),.clk(gclk));
	jnot g3480(.din(w_n4121_0[1]),.dout(n4122),.clk(gclk));
	jand g3481(.dina(w_n4122_0[1]),.dinb(w_n4118_0[2]),.dout(n4123),.clk(gclk));
	jor g3482(.dina(n4123),.dinb(w_n4115_0[1]),.dout(n4124),.clk(gclk));
	jor g3483(.dina(n4124),.dinb(w_n4107_0[1]),.dout(n4125),.clk(gclk));
	jor g3484(.dina(w_n4125_0[1]),.dinb(n4090),.dout(n4126),.clk(gclk));
	jor g3485(.dina(w_n4097_0[1]),.dinb(w_n4094_0[0]),.dout(n4127),.clk(gclk));
	jor g3486(.dina(w_n4122_0[0]),.dinb(w_n4118_0[1]),.dout(n4128),.clk(gclk));
	jor g3487(.dina(n4128),.dinb(w_n4115_0[0]),.dout(n4129),.clk(gclk));
	jor g3488(.dina(w_n4114_0[1]),.dinb(w_n4111_0[0]),.dout(n4130),.clk(gclk));
	jor g3489(.dina(w_n4105_0[0]),.dinb(w_n4101_0[1]),.dout(n4131),.clk(gclk));
	jand g3490(.dina(n4131),.dinb(n4130),.dout(n4132),.clk(gclk));
	jand g3491(.dina(n4132),.dinb(n4129),.dout(n4133),.clk(gclk));
	jor g3492(.dina(n4133),.dinb(w_n4107_0[0]),.dout(n4134),.clk(gclk));
	jand g3493(.dina(n4134),.dinb(n4127),.dout(n4135),.clk(gclk));
	jand g3494(.dina(w_n4135_0[1]),.dinb(n4126),.dout(n4136),.clk(gclk));
	jand g3495(.dina(w_n2628_25[2]),.dinb(w_in0116_0[0]),.dout(n4137),.clk(gclk));
	jand g3496(.dina(w_n2783_26[0]),.dinb(w_in1116_0[0]),.dout(n4138),.clk(gclk));
	jor g3497(.dina(n4138),.dinb(n4137),.dout(n4139),.clk(gclk));
	jnot g3498(.din(w_n4139_0[1]),.dout(n4140),.clk(gclk));
	jand g3499(.dina(w_n1556_25[0]),.dinb(w_in2116_0[0]),.dout(n4141),.clk(gclk));
	jand g3500(.dina(w_n1711_25[2]),.dinb(w_in3116_0[0]),.dout(n4142),.clk(gclk));
	jor g3501(.dina(n4142),.dinb(n4141),.dout(n4143),.clk(gclk));
	jand g3502(.dina(w_n4143_0[2]),.dinb(w_n4140_0[1]),.dout(n4144),.clk(gclk));
	jand g3503(.dina(w_n2628_25[1]),.dinb(w_in0117_0[0]),.dout(n4145),.clk(gclk));
	jand g3504(.dina(w_n2783_25[2]),.dinb(w_in1117_0[0]),.dout(n4146),.clk(gclk));
	jor g3505(.dina(n4146),.dinb(n4145),.dout(n4147),.clk(gclk));
	jnot g3506(.din(w_n4147_0[1]),.dout(n4148),.clk(gclk));
	jand g3507(.dina(w_n1556_24[2]),.dinb(w_in2117_0[0]),.dout(n4149),.clk(gclk));
	jand g3508(.dina(w_n1711_25[1]),.dinb(w_in3117_0[0]),.dout(n4150),.clk(gclk));
	jor g3509(.dina(n4150),.dinb(n4149),.dout(n4151),.clk(gclk));
	jand g3510(.dina(w_n4151_0[2]),.dinb(w_n4148_0[1]),.dout(n4152),.clk(gclk));
	jand g3511(.dina(w_n2628_25[0]),.dinb(w_in0119_0[0]),.dout(n4153),.clk(gclk));
	jand g3512(.dina(w_n2783_25[1]),.dinb(w_in1119_0[0]),.dout(n4154),.clk(gclk));
	jor g3513(.dina(n4154),.dinb(n4153),.dout(n4155),.clk(gclk));
	jnot g3514(.din(w_n4155_0[1]),.dout(n4156),.clk(gclk));
	jand g3515(.dina(w_n1556_24[1]),.dinb(w_in2119_0[0]),.dout(n4157),.clk(gclk));
	jand g3516(.dina(w_n1711_25[0]),.dinb(w_in3119_0[0]),.dout(n4158),.clk(gclk));
	jor g3517(.dina(n4158),.dinb(n4157),.dout(n4159),.clk(gclk));
	jand g3518(.dina(w_n4159_0[2]),.dinb(w_n4156_0[1]),.dout(n4160),.clk(gclk));
	jand g3519(.dina(w_n1556_24[0]),.dinb(w_in2118_0[0]),.dout(n4161),.clk(gclk));
	jand g3520(.dina(w_n1711_24[2]),.dinb(w_in3118_0[0]),.dout(n4162),.clk(gclk));
	jor g3521(.dina(n4162),.dinb(n4161),.dout(n4163),.clk(gclk));
	jand g3522(.dina(w_n2628_24[2]),.dinb(w_in0118_0[0]),.dout(n4164),.clk(gclk));
	jand g3523(.dina(w_n2783_25[0]),.dinb(w_in1118_0[0]),.dout(n4165),.clk(gclk));
	jor g3524(.dina(n4165),.dinb(n4164),.dout(n4166),.clk(gclk));
	jnot g3525(.din(w_n4166_0[1]),.dout(n4167),.clk(gclk));
	jand g3526(.dina(w_n4167_0[1]),.dinb(w_n4163_0[2]),.dout(n4168),.clk(gclk));
	jor g3527(.dina(n4168),.dinb(w_n4160_0[1]),.dout(n4169),.clk(gclk));
	jor g3528(.dina(n4169),.dinb(n4152),.dout(n4170),.clk(gclk));
	jor g3529(.dina(w_n4170_0[1]),.dinb(n4144),.dout(n4171),.clk(gclk));
	jor g3530(.dina(w_n4171_0[1]),.dinb(n4136),.dout(n4172),.clk(gclk));
	jor g3531(.dina(w_n4151_0[1]),.dinb(w_n4148_0[0]),.dout(n4173),.clk(gclk));
	jor g3532(.dina(w_n4143_0[1]),.dinb(w_n4140_0[0]),.dout(n4174),.clk(gclk));
	jand g3533(.dina(n4174),.dinb(n4173),.dout(n4175),.clk(gclk));
	jor g3534(.dina(n4175),.dinb(w_n4170_0[0]),.dout(n4176),.clk(gclk));
	jor g3535(.dina(w_n4159_0[1]),.dinb(w_n4156_0[0]),.dout(n4177),.clk(gclk));
	jor g3536(.dina(w_n4167_0[0]),.dinb(w_n4163_0[1]),.dout(n4178),.clk(gclk));
	jor g3537(.dina(n4178),.dinb(w_n4160_0[0]),.dout(n4179),.clk(gclk));
	jand g3538(.dina(n4179),.dinb(n4177),.dout(n4180),.clk(gclk));
	jand g3539(.dina(n4180),.dinb(n4176),.dout(n4181),.clk(gclk));
	jand g3540(.dina(w_n4181_0[1]),.dinb(n4172),.dout(n4182),.clk(gclk));
	jand g3541(.dina(w_n2628_24[1]),.dinb(w_in0123_0[0]),.dout(n4183),.clk(gclk));
	jand g3542(.dina(w_n2783_24[2]),.dinb(w_in1123_0[0]),.dout(n4184),.clk(gclk));
	jor g3543(.dina(n4184),.dinb(n4183),.dout(n4185),.clk(gclk));
	jnot g3544(.din(w_n4185_0[1]),.dout(n4186),.clk(gclk));
	jand g3545(.dina(w_n1556_23[2]),.dinb(w_in2123_0[0]),.dout(n4187),.clk(gclk));
	jand g3546(.dina(w_n1711_24[1]),.dinb(w_in3123_0[0]),.dout(n4188),.clk(gclk));
	jor g3547(.dina(n4188),.dinb(n4187),.dout(n4189),.clk(gclk));
	jand g3548(.dina(w_n4189_0[2]),.dinb(w_n4186_0[1]),.dout(n4190),.clk(gclk));
	jand g3549(.dina(w_n1556_23[1]),.dinb(w_in2122_0[0]),.dout(n4191),.clk(gclk));
	jand g3550(.dina(w_n1711_24[0]),.dinb(w_in3122_0[0]),.dout(n4192),.clk(gclk));
	jor g3551(.dina(n4192),.dinb(n4191),.dout(n4193),.clk(gclk));
	jand g3552(.dina(w_n2628_24[0]),.dinb(w_in0122_0[0]),.dout(n4194),.clk(gclk));
	jand g3553(.dina(w_n2783_24[1]),.dinb(w_in1122_0[0]),.dout(n4195),.clk(gclk));
	jor g3554(.dina(n4195),.dinb(n4194),.dout(n4196),.clk(gclk));
	jnot g3555(.din(w_n4196_0[1]),.dout(n4197),.clk(gclk));
	jand g3556(.dina(w_n4197_0[1]),.dinb(w_n4193_0[2]),.dout(n4198),.clk(gclk));
	jor g3557(.dina(n4198),.dinb(n4190),.dout(n4199),.clk(gclk));
	jand g3558(.dina(w_n2628_23[2]),.dinb(w_in0121_0[0]),.dout(n4200),.clk(gclk));
	jand g3559(.dina(w_n2783_24[0]),.dinb(w_in1121_0[0]),.dout(n4201),.clk(gclk));
	jor g3560(.dina(n4201),.dinb(n4200),.dout(n4202),.clk(gclk));
	jnot g3561(.din(w_n4202_0[1]),.dout(n4203),.clk(gclk));
	jand g3562(.dina(w_n1556_23[0]),.dinb(w_in2121_0[0]),.dout(n4204),.clk(gclk));
	jand g3563(.dina(w_n1711_23[2]),.dinb(w_in3121_0[0]),.dout(n4205),.clk(gclk));
	jor g3564(.dina(n4205),.dinb(n4204),.dout(n4206),.clk(gclk));
	jand g3565(.dina(w_n4206_0[2]),.dinb(w_n4203_0[1]),.dout(n4207),.clk(gclk));
	jand g3566(.dina(w_n1556_22[2]),.dinb(w_in2120_0[0]),.dout(n4208),.clk(gclk));
	jand g3567(.dina(w_n1711_23[1]),.dinb(w_in3120_0[0]),.dout(n4209),.clk(gclk));
	jor g3568(.dina(n4209),.dinb(n4208),.dout(n4210),.clk(gclk));
	jand g3569(.dina(w_n2628_23[1]),.dinb(w_in0120_0[0]),.dout(n4211),.clk(gclk));
	jand g3570(.dina(w_n2783_23[2]),.dinb(w_in1120_0[0]),.dout(n4212),.clk(gclk));
	jor g3571(.dina(n4212),.dinb(n4211),.dout(n4213),.clk(gclk));
	jnot g3572(.din(w_n4213_0[1]),.dout(n4214),.clk(gclk));
	jand g3573(.dina(w_n4214_0[1]),.dinb(w_n4210_0[2]),.dout(n4215),.clk(gclk));
	jor g3574(.dina(n4215),.dinb(w_n4207_0[1]),.dout(n4216),.clk(gclk));
	jor g3575(.dina(n4216),.dinb(w_n4199_0[1]),.dout(n4217),.clk(gclk));
	jor g3576(.dina(w_n4217_0[1]),.dinb(n4182),.dout(n4218),.clk(gclk));
	jor g3577(.dina(w_n4189_0[1]),.dinb(w_n4186_0[0]),.dout(n4219),.clk(gclk));
	jor g3578(.dina(w_n4214_0[0]),.dinb(w_n4210_0[1]),.dout(n4220),.clk(gclk));
	jor g3579(.dina(n4220),.dinb(w_n4207_0[0]),.dout(n4221),.clk(gclk));
	jor g3580(.dina(w_n4206_0[1]),.dinb(w_n4203_0[0]),.dout(n4222),.clk(gclk));
	jor g3581(.dina(w_n4197_0[0]),.dinb(w_n4193_0[1]),.dout(n4223),.clk(gclk));
	jand g3582(.dina(n4223),.dinb(n4222),.dout(n4224),.clk(gclk));
	jand g3583(.dina(n4224),.dinb(n4221),.dout(n4225),.clk(gclk));
	jor g3584(.dina(n4225),.dinb(w_n4199_0[0]),.dout(n4226),.clk(gclk));
	jand g3585(.dina(n4226),.dinb(n4219),.dout(n4227),.clk(gclk));
	jand g3586(.dina(w_n4227_0[1]),.dinb(n4218),.dout(n4228),.clk(gclk));
	jand g3587(.dina(w_n2628_23[0]),.dinb(w_in0126_0[0]),.dout(n4229),.clk(gclk));
	jand g3588(.dina(w_n2783_23[1]),.dinb(w_in1126_0[0]),.dout(n4230),.clk(gclk));
	jor g3589(.dina(n4230),.dinb(n4229),.dout(n4231),.clk(gclk));
	jnot g3590(.din(w_n4231_0[1]),.dout(n4232),.clk(gclk));
	jand g3591(.dina(w_n1556_22[1]),.dinb(w_in2126_0[0]),.dout(n4233),.clk(gclk));
	jand g3592(.dina(w_n1711_23[0]),.dinb(w_in3126_0[0]),.dout(n4234),.clk(gclk));
	jor g3593(.dina(n4234),.dinb(n4233),.dout(n4235),.clk(gclk));
	jand g3594(.dina(w_n4235_0[2]),.dinb(w_n4232_0[1]),.dout(n4236),.clk(gclk));
	jand g3595(.dina(w_n2628_22[2]),.dinb(w_in0125_0[0]),.dout(n4237),.clk(gclk));
	jand g3596(.dina(w_n2783_23[0]),.dinb(w_in1125_0[0]),.dout(n4238),.clk(gclk));
	jor g3597(.dina(n4238),.dinb(n4237),.dout(n4239),.clk(gclk));
	jnot g3598(.din(w_n4239_0[1]),.dout(n4240),.clk(gclk));
	jand g3599(.dina(w_n1556_22[0]),.dinb(w_in2125_0[0]),.dout(n4241),.clk(gclk));
	jand g3600(.dina(w_n1711_22[2]),.dinb(w_in3125_0[0]),.dout(n4242),.clk(gclk));
	jor g3601(.dina(n4242),.dinb(n4241),.dout(n4243),.clk(gclk));
	jand g3602(.dina(w_n4243_0[2]),.dinb(w_n4240_0[1]),.dout(n4244),.clk(gclk));
	jor g3603(.dina(n4244),.dinb(n4236),.dout(n4245),.clk(gclk));
	jand g3604(.dina(w_in3127_0[0]),.dinb(w_in2127_0[0]),.dout(n4246),.clk(gclk));
	jnot g3605(.din(w_n4246_0[1]),.dout(n4247),.clk(gclk));
	jand g3606(.dina(w_in1127_0[0]),.dinb(w_in0127_0[0]),.dout(n4248),.clk(gclk));
	jand g3607(.dina(w_n4248_0[2]),.dinb(w_n4247_0[1]),.dout(n4249),.clk(gclk));
	jand g3608(.dina(w_n2628_22[1]),.dinb(w_in0124_0[0]),.dout(n4250),.clk(gclk));
	jand g3609(.dina(w_n2783_22[2]),.dinb(w_in1124_0[0]),.dout(n4251),.clk(gclk));
	jor g3610(.dina(n4251),.dinb(n4250),.dout(n4252),.clk(gclk));
	jnot g3611(.din(w_n4252_0[1]),.dout(n4253),.clk(gclk));
	jand g3612(.dina(w_n1556_21[2]),.dinb(w_in2124_0[0]),.dout(n4254),.clk(gclk));
	jand g3613(.dina(w_n1711_22[1]),.dinb(w_in3124_0[0]),.dout(n4255),.clk(gclk));
	jor g3614(.dina(n4255),.dinb(n4254),.dout(n4256),.clk(gclk));
	jand g3615(.dina(w_n4256_0[2]),.dinb(w_n4253_0[1]),.dout(n4257),.clk(gclk));
	jor g3616(.dina(n4257),.dinb(w_n4249_0[1]),.dout(n4258),.clk(gclk));
	jor g3617(.dina(n4258),.dinb(w_n4245_0[1]),.dout(n4259),.clk(gclk));
	jor g3618(.dina(w_n4259_0[1]),.dinb(n4228),.dout(n4260),.clk(gclk));
	jor g3619(.dina(w_n4256_0[1]),.dinb(w_n4253_0[0]),.dout(n4261),.clk(gclk));
	jor g3620(.dina(w_n4243_0[1]),.dinb(w_n4240_0[0]),.dout(n4262),.clk(gclk));
	jand g3621(.dina(n4262),.dinb(n4261),.dout(n4263),.clk(gclk));
	jor g3622(.dina(n4263),.dinb(w_n4245_0[0]),.dout(n4264),.clk(gclk));
	jor g3623(.dina(w_n4248_0[1]),.dinb(w_n4247_0[0]),.dout(n4265),.clk(gclk));
	jor g3624(.dina(w_n4235_0[1]),.dinb(w_n4232_0[0]),.dout(n4266),.clk(gclk));
	jand g3625(.dina(n4266),.dinb(n4265),.dout(n4267),.clk(gclk));
	jand g3626(.dina(n4267),.dinb(n4264),.dout(n4268),.clk(gclk));
	jor g3627(.dina(n4268),.dinb(w_n4249_0[0]),.dout(n4269),.clk(gclk));
	jand g3628(.dina(w_n4269_0[1]),.dinb(n4260),.dout(address[1]),.clk(gclk));
	jand g3629(.dina(w_address1_63[1]),.dinb(w_n1713_0[0]),.dout(n4271),.clk(gclk));
	jand g3630(.dina(w_n2628_22[0]),.dinb(w_in00_0[0]),.dout(n4272),.clk(gclk));
	jand g3631(.dina(w_n2783_22[1]),.dinb(w_in10_0[0]),.dout(n4273),.clk(gclk));
	jor g3632(.dina(n4273),.dinb(n4272),.dout(n4274),.clk(gclk));
	jnot g3633(.din(w_n2790_0[0]),.dout(n4275),.clk(gclk));
	jnot g3634(.din(w_n2862_0[0]),.dout(n4276),.clk(gclk));
	jnot g3635(.din(w_n2896_0[1]),.dout(n4277),.clk(gclk));
	jnot g3636(.din(w_n2908_0[0]),.dout(n4278),.clk(gclk));
	jnot g3637(.din(w_n2909_0[0]),.dout(n4279),.clk(gclk));
	jnot g3638(.din(w_n2917_0[0]),.dout(n4280),.clk(gclk));
	jnot g3639(.din(w_n2925_0[0]),.dout(n4281),.clk(gclk));
	jnot g3640(.din(w_n2983_0[1]),.dout(n4282),.clk(gclk));
	jnot g3641(.din(w_n3010_0[0]),.dout(n4283),.clk(gclk));
	jnot g3642(.din(w_n3011_0[0]),.dout(n4284),.clk(gclk));
	jnot g3643(.din(w_n3018_0[0]),.dout(n4285),.clk(gclk));
	jnot g3644(.din(w_n3021_0[1]),.dout(n4286),.clk(gclk));
	jor g3645(.dina(w_n1711_22[0]),.dinb(w_n1589_0[0]),.dout(n4287),.clk(gclk));
	jor g3646(.dina(w_n1556_21[1]),.dinb(w_n788_0[0]),.dout(n4288),.clk(gclk));
	jand g3647(.dina(n4288),.dinb(n4287),.dout(n4289),.clk(gclk));
	jand g3648(.dina(w_n4274_0[1]),.dinb(n4289),.dout(n4290),.clk(gclk));
	jand g3649(.dina(w_n2628_21[2]),.dinb(w_in01_0[1]),.dout(n4291),.clk(gclk));
	jand g3650(.dina(w_n2783_22[0]),.dinb(w_in11_0[1]),.dout(n4292),.clk(gclk));
	jor g3651(.dina(n4292),.dinb(n4291),.dout(n4293),.clk(gclk));
	jor g3652(.dina(w_n4293_0[2]),.dinb(w_n4290_0[1]),.dout(n4294),.clk(gclk));
	jand g3653(.dina(n4294),.dinb(n4286),.dout(n4295),.clk(gclk));
	jand g3654(.dina(w_n2628_21[1]),.dinb(w_in02_0[0]),.dout(n4296),.clk(gclk));
	jand g3655(.dina(w_n2783_21[2]),.dinb(w_in12_0[0]),.dout(n4297),.clk(gclk));
	jor g3656(.dina(n4297),.dinb(n4296),.dout(n4298),.clk(gclk));
	jor g3657(.dina(w_n1711_21[2]),.dinb(w_n782_0[0]),.dout(n4299),.clk(gclk));
	jor g3658(.dina(w_n1556_21[0]),.dinb(w_n780_0[0]),.dout(n4300),.clk(gclk));
	jand g3659(.dina(n4300),.dinb(n4299),.dout(n4301),.clk(gclk));
	jand g3660(.dina(n4301),.dinb(w_n4298_0[1]),.dout(n4302),.clk(gclk));
	jand g3661(.dina(w_n4293_0[1]),.dinb(w_n4290_0[0]),.dout(n4303),.clk(gclk));
	jor g3662(.dina(n4303),.dinb(n4302),.dout(n4304),.clk(gclk));
	jor g3663(.dina(n4304),.dinb(n4295),.dout(n4305),.clk(gclk));
	jand g3664(.dina(n4305),.dinb(n4285),.dout(n4306),.clk(gclk));
	jor g3665(.dina(n4306),.dinb(n4284),.dout(n4307),.clk(gclk));
	jand g3666(.dina(n4307),.dinb(n4283),.dout(n4308),.clk(gclk));
	jnot g3667(.din(w_n3040_0[2]),.dout(n4309),.clk(gclk));
	jand g3668(.dina(w_n4309_0[1]),.dinb(w_n4308_0[1]),.dout(n4310),.clk(gclk));
	jor g3669(.dina(n4310),.dinb(w_n3001_0[1]),.dout(n4311),.clk(gclk));
	jor g3670(.dina(w_n4309_0[0]),.dinb(w_n4308_0[0]),.dout(n4312),.clk(gclk));
	jand g3671(.dina(n4312),.dinb(n4311),.dout(n4313),.clk(gclk));
	jnot g3672(.din(w_n3047_0[2]),.dout(n4314),.clk(gclk));
	jand g3673(.dina(w_n4314_0[1]),.dinb(w_n4313_0[1]),.dout(n4315),.clk(gclk));
	jor g3674(.dina(n4315),.dinb(w_n2997_0[1]),.dout(n4316),.clk(gclk));
	jor g3675(.dina(w_n4314_0[0]),.dinb(w_n4313_0[0]),.dout(n4317),.clk(gclk));
	jnot g3676(.din(w_n3058_0[0]),.dout(n4318),.clk(gclk));
	jand g3677(.dina(n4318),.dinb(n4317),.dout(n4319),.clk(gclk));
	jand g3678(.dina(n4319),.dinb(n4316),.dout(n4320),.clk(gclk));
	jnot g3679(.din(w_n3061_0[0]),.dout(n4321),.clk(gclk));
	jor g3680(.dina(n4321),.dinb(n4320),.dout(n4322),.clk(gclk));
	jand g3681(.dina(n4322),.dinb(w_n2993_0[0]),.dout(n4323),.clk(gclk));
	jor g3682(.dina(n4323),.dinb(w_n2991_0[0]),.dout(n4324),.clk(gclk));
	jor g3683(.dina(w_n3067_1[0]),.dinb(w_n4324_0[1]),.dout(n4325),.clk(gclk));
	jand g3684(.dina(n4325),.dinb(n4282),.dout(n4326),.clk(gclk));
	jand g3685(.dina(w_n3067_0[2]),.dinb(w_n4324_0[0]),.dout(n4327),.clk(gclk));
	jor g3686(.dina(n4327),.dinb(n4326),.dout(n4328),.clk(gclk));
	jand g3687(.dina(n4328),.dinb(w_n2979_0[0]),.dout(n4329),.clk(gclk));
	jor g3688(.dina(n4329),.dinb(w_n2977_0[0]),.dout(n4330),.clk(gclk));
	jand g3689(.dina(n4330),.dinb(w_n2968_0[0]),.dout(n4331),.clk(gclk));
	jor g3690(.dina(n4331),.dinb(w_n2966_0[0]),.dout(n4332),.clk(gclk));
	jand g3691(.dina(n4332),.dinb(w_n2957_0[0]),.dout(n4333),.clk(gclk));
	jor g3692(.dina(n4333),.dinb(w_n2955_0[0]),.dout(n4334),.clk(gclk));
	jand g3693(.dina(n4334),.dinb(w_n2946_0[0]),.dout(n4335),.clk(gclk));
	jor g3694(.dina(n4335),.dinb(w_n2944_0[0]),.dout(n4336),.clk(gclk));
	jand g3695(.dina(n4336),.dinb(w_n2935_0[0]),.dout(n4337),.clk(gclk));
	jor g3696(.dina(n4337),.dinb(w_n2933_0[0]),.dout(n4338),.clk(gclk));
	jand g3697(.dina(n4338),.dinb(n4281),.dout(n4339),.clk(gclk));
	jnot g3698(.din(w_n3086_0[0]),.dout(n4340),.clk(gclk));
	jor g3699(.dina(n4340),.dinb(n4339),.dout(n4341),.clk(gclk));
	jand g3700(.dina(n4341),.dinb(n4280),.dout(n4342),.clk(gclk));
	jor g3701(.dina(n4342),.dinb(n4279),.dout(n4343),.clk(gclk));
	jand g3702(.dina(n4343),.dinb(n4278),.dout(n4344),.clk(gclk));
	jor g3703(.dina(w_n4344_0[1]),.dinb(w_n2899_1[0]),.dout(n4345),.clk(gclk));
	jand g3704(.dina(n4345),.dinb(n4277),.dout(n4346),.clk(gclk));
	jand g3705(.dina(w_n4344_0[0]),.dinb(w_n2899_0[2]),.dout(n4347),.clk(gclk));
	jor g3706(.dina(n4347),.dinb(w_n3100_0[0]),.dout(n4348),.clk(gclk));
	jor g3707(.dina(n4348),.dinb(n4346),.dout(n4349),.clk(gclk));
	jand g3708(.dina(w_n3107_0[0]),.dinb(n4349),.dout(n4350),.clk(gclk));
	jor g3709(.dina(n4350),.dinb(w_n2892_0[0]),.dout(n4351),.clk(gclk));
	jand g3710(.dina(n4351),.dinb(w_n2883_0[0]),.dout(n4352),.clk(gclk));
	jor g3711(.dina(n4352),.dinb(w_n2881_0[0]),.dout(n4353),.clk(gclk));
	jand g3712(.dina(n4353),.dinb(w_n2872_0[0]),.dout(n4354),.clk(gclk));
	jor g3713(.dina(n4354),.dinb(w_n2870_0[0]),.dout(n4355),.clk(gclk));
	jand g3714(.dina(n4355),.dinb(n4276),.dout(n4356),.clk(gclk));
	jnot g3715(.din(w_n3126_0[0]),.dout(n4357),.clk(gclk));
	jor g3716(.dina(n4357),.dinb(n4356),.dout(n4358),.clk(gclk));
	jand g3717(.dina(w_n3130_0[0]),.dinb(n4358),.dout(n4359),.clk(gclk));
	jor g3718(.dina(n4359),.dinb(w_n2853_0[0]),.dout(n4360),.clk(gclk));
	jand g3719(.dina(n4360),.dinb(w_n2844_0[0]),.dout(n4361),.clk(gclk));
	jor g3720(.dina(n4361),.dinb(w_n2842_0[0]),.dout(n4362),.clk(gclk));
	jand g3721(.dina(n4362),.dinb(w_n2833_0[0]),.dout(n4363),.clk(gclk));
	jor g3722(.dina(n4363),.dinb(w_n2831_0[0]),.dout(n4364),.clk(gclk));
	jand g3723(.dina(n4364),.dinb(w_n2822_0[0]),.dout(n4365),.clk(gclk));
	jor g3724(.dina(n4365),.dinb(w_n2820_0[0]),.dout(n4366),.clk(gclk));
	jand g3725(.dina(n4366),.dinb(w_n2811_0[0]),.dout(n4367),.clk(gclk));
	jor g3726(.dina(n4367),.dinb(w_n2809_0[0]),.dout(n4368),.clk(gclk));
	jand g3727(.dina(n4368),.dinb(w_n2800_0[0]),.dout(n4369),.clk(gclk));
	jor g3728(.dina(n4369),.dinb(w_n2798_0[0]),.dout(n4370),.clk(gclk));
	jand g3729(.dina(n4370),.dinb(n4275),.dout(n4371),.clk(gclk));
	jnot g3730(.din(w_n3155_0[0]),.dout(n4372),.clk(gclk));
	jor g3731(.dina(n4372),.dinb(n4371),.dout(n4373),.clk(gclk));
	jand g3732(.dina(w_n3233_0[0]),.dinb(n4373),.dout(n4374),.clk(gclk));
	jnot g3733(.din(w_n3255_0[0]),.dout(n4375),.clk(gclk));
	jor g3734(.dina(n4375),.dinb(n4374),.dout(n4376),.clk(gclk));
	jnot g3735(.din(w_n3327_0[0]),.dout(n4377),.clk(gclk));
	jand g3736(.dina(n4377),.dinb(n4376),.dout(n4378),.clk(gclk));
	jnot g3737(.din(w_n3348_0[0]),.dout(n4379),.clk(gclk));
	jor g3738(.dina(n4379),.dinb(n4378),.dout(n4380),.clk(gclk));
	jnot g3739(.din(w_n3423_0[0]),.dout(n4381),.clk(gclk));
	jand g3740(.dina(n4381),.dinb(n4380),.dout(n4382),.clk(gclk));
	jnot g3741(.din(w_n3444_0[0]),.dout(n4383),.clk(gclk));
	jor g3742(.dina(n4383),.dinb(n4382),.dout(n4384),.clk(gclk));
	jnot g3743(.din(w_n3516_0[0]),.dout(n4385),.clk(gclk));
	jand g3744(.dina(n4385),.dinb(n4384),.dout(n4386),.clk(gclk));
	jnot g3745(.din(w_n3537_0[0]),.dout(n4387),.clk(gclk));
	jor g3746(.dina(n4387),.dinb(n4386),.dout(n4388),.clk(gclk));
	jnot g3747(.din(w_n3573_0[0]),.dout(n4389),.clk(gclk));
	jand g3748(.dina(n4389),.dinb(n4388),.dout(n4390),.clk(gclk));
	jnot g3749(.din(w_n3583_0[0]),.dout(n4391),.clk(gclk));
	jor g3750(.dina(n4391),.dinb(n4390),.dout(n4392),.clk(gclk));
	jnot g3751(.din(w_n3619_0[0]),.dout(n4393),.clk(gclk));
	jand g3752(.dina(n4393),.dinb(n4392),.dout(n4394),.clk(gclk));
	jnot g3753(.din(w_n3629_0[0]),.dout(n4395),.clk(gclk));
	jor g3754(.dina(n4395),.dinb(n4394),.dout(n4396),.clk(gclk));
	jnot g3755(.din(w_n3665_0[0]),.dout(n4397),.clk(gclk));
	jand g3756(.dina(n4397),.dinb(n4396),.dout(n4398),.clk(gclk));
	jnot g3757(.din(w_n3675_0[0]),.dout(n4399),.clk(gclk));
	jor g3758(.dina(n4399),.dinb(n4398),.dout(n4400),.clk(gclk));
	jnot g3759(.din(w_n3711_0[0]),.dout(n4401),.clk(gclk));
	jand g3760(.dina(n4401),.dinb(n4400),.dout(n4402),.clk(gclk));
	jnot g3761(.din(w_n3721_0[0]),.dout(n4403),.clk(gclk));
	jor g3762(.dina(n4403),.dinb(n4402),.dout(n4404),.clk(gclk));
	jnot g3763(.din(w_n3757_0[0]),.dout(n4405),.clk(gclk));
	jand g3764(.dina(n4405),.dinb(n4404),.dout(n4406),.clk(gclk));
	jnot g3765(.din(w_n3767_0[0]),.dout(n4407),.clk(gclk));
	jor g3766(.dina(n4407),.dinb(n4406),.dout(n4408),.clk(gclk));
	jnot g3767(.din(w_n3803_0[0]),.dout(n4409),.clk(gclk));
	jand g3768(.dina(n4409),.dinb(n4408),.dout(n4410),.clk(gclk));
	jnot g3769(.din(w_n3813_0[0]),.dout(n4411),.clk(gclk));
	jor g3770(.dina(n4411),.dinb(n4410),.dout(n4412),.clk(gclk));
	jnot g3771(.din(w_n3849_0[0]),.dout(n4413),.clk(gclk));
	jand g3772(.dina(n4413),.dinb(n4412),.dout(n4414),.clk(gclk));
	jnot g3773(.din(w_n3859_0[0]),.dout(n4415),.clk(gclk));
	jor g3774(.dina(n4415),.dinb(n4414),.dout(n4416),.clk(gclk));
	jnot g3775(.din(w_n3895_0[0]),.dout(n4417),.clk(gclk));
	jand g3776(.dina(n4417),.dinb(n4416),.dout(n4418),.clk(gclk));
	jnot g3777(.din(w_n3905_0[0]),.dout(n4419),.clk(gclk));
	jor g3778(.dina(n4419),.dinb(n4418),.dout(n4420),.clk(gclk));
	jnot g3779(.din(w_n3941_0[0]),.dout(n4421),.clk(gclk));
	jand g3780(.dina(n4421),.dinb(n4420),.dout(n4422),.clk(gclk));
	jnot g3781(.din(w_n3951_0[0]),.dout(n4423),.clk(gclk));
	jor g3782(.dina(n4423),.dinb(n4422),.dout(n4424),.clk(gclk));
	jnot g3783(.din(w_n3987_0[0]),.dout(n4425),.clk(gclk));
	jand g3784(.dina(n4425),.dinb(n4424),.dout(n4426),.clk(gclk));
	jnot g3785(.din(w_n3997_0[0]),.dout(n4427),.clk(gclk));
	jor g3786(.dina(n4427),.dinb(n4426),.dout(n4428),.clk(gclk));
	jnot g3787(.din(w_n4033_0[0]),.dout(n4429),.clk(gclk));
	jand g3788(.dina(n4429),.dinb(n4428),.dout(n4430),.clk(gclk));
	jnot g3789(.din(w_n4043_0[0]),.dout(n4431),.clk(gclk));
	jor g3790(.dina(n4431),.dinb(n4430),.dout(n4432),.clk(gclk));
	jnot g3791(.din(w_n4079_0[0]),.dout(n4433),.clk(gclk));
	jand g3792(.dina(n4433),.dinb(n4432),.dout(n4434),.clk(gclk));
	jnot g3793(.din(w_n4089_0[0]),.dout(n4435),.clk(gclk));
	jor g3794(.dina(n4435),.dinb(n4434),.dout(n4436),.clk(gclk));
	jnot g3795(.din(w_n4125_0[0]),.dout(n4437),.clk(gclk));
	jand g3796(.dina(n4437),.dinb(n4436),.dout(n4438),.clk(gclk));
	jnot g3797(.din(w_n4135_0[0]),.dout(n4439),.clk(gclk));
	jor g3798(.dina(n4439),.dinb(n4438),.dout(n4440),.clk(gclk));
	jnot g3799(.din(w_n4171_0[0]),.dout(n4441),.clk(gclk));
	jand g3800(.dina(n4441),.dinb(n4440),.dout(n4442),.clk(gclk));
	jnot g3801(.din(w_n4181_0[0]),.dout(n4443),.clk(gclk));
	jor g3802(.dina(n4443),.dinb(n4442),.dout(n4444),.clk(gclk));
	jnot g3803(.din(w_n4217_0[0]),.dout(n4445),.clk(gclk));
	jand g3804(.dina(n4445),.dinb(n4444),.dout(n4446),.clk(gclk));
	jnot g3805(.din(w_n4227_0[0]),.dout(n4447),.clk(gclk));
	jor g3806(.dina(n4447),.dinb(n4446),.dout(n4448),.clk(gclk));
	jnot g3807(.din(w_n4259_0[0]),.dout(n4449),.clk(gclk));
	jand g3808(.dina(n4449),.dinb(n4448),.dout(n4450),.clk(gclk));
	jnot g3809(.din(w_n4269_0[0]),.dout(n4451),.clk(gclk));
	jor g3810(.dina(n4451),.dinb(n4450),.dout(n4452),.clk(gclk));
	jand g3811(.dina(w_n4452_63[1]),.dinb(w_n4274_0[0]),.dout(n4453),.clk(gclk));
	jor g3812(.dina(n4453),.dinb(n4271),.dout(result[0]),.clk(gclk));
	jor g3813(.dina(w_address1_63[0]),.dinb(w_n4293_0[0]),.dout(n4455),.clk(gclk));
	jor g3814(.dina(w_n4452_63[0]),.dinb(w_n3021_0[0]),.dout(n4456),.clk(gclk));
	jand g3815(.dina(n4456),.dinb(n4455),.dout(result[1]),.clk(gclk));
	jor g3816(.dina(w_address1_62[2]),.dinb(w_n4298_0[0]),.dout(n4458),.clk(gclk));
	jor g3817(.dina(w_n4452_62[2]),.dinb(w_n3017_0[0]),.dout(n4459),.clk(gclk));
	jand g3818(.dina(n4459),.dinb(n4458),.dout(result[2]),.clk(gclk));
	jor g3819(.dina(w_address1_62[1]),.dinb(w_n3005_0[0]),.dout(n4461),.clk(gclk));
	jor g3820(.dina(w_n4452_62[1]),.dinb(w_n3009_0[0]),.dout(n4462),.clk(gclk));
	jand g3821(.dina(n4462),.dinb(n4461),.dout(result[3]),.clk(gclk));
	jand g3822(.dina(w_address1_62[0]),.dinb(w_n3040_0[1]),.dout(n4464),.clk(gclk));
	jand g3823(.dina(w_n4452_62[0]),.dinb(w_n3001_0[0]),.dout(n4465),.clk(gclk));
	jor g3824(.dina(n4465),.dinb(n4464),.dout(result[4]),.clk(gclk));
	jand g3825(.dina(w_address1_61[2]),.dinb(w_n3047_0[1]),.dout(n4467),.clk(gclk));
	jand g3826(.dina(w_n4452_61[2]),.dinb(w_n2997_0[0]),.dout(n4468),.clk(gclk));
	jor g3827(.dina(n4468),.dinb(n4467),.dout(result[5]),.clk(gclk));
	jand g3828(.dina(w_address1_61[1]),.dinb(w_n3057_0[0]),.dout(n4470),.clk(gclk));
	jand g3829(.dina(w_n4452_61[1]),.dinb(w_n3053_0[0]),.dout(n4471),.clk(gclk));
	jor g3830(.dina(n4471),.dinb(n4470),.dout(result[6]),.clk(gclk));
	jor g3831(.dina(w_address1_61[0]),.dinb(w_n2986_0[0]),.dout(n4473),.clk(gclk));
	jor g3832(.dina(w_n4452_61[0]),.dinb(w_n2989_0[0]),.dout(n4474),.clk(gclk));
	jand g3833(.dina(n4474),.dinb(n4473),.dout(result[7]),.clk(gclk));
	jand g3834(.dina(w_address1_60[2]),.dinb(w_n2983_0[0]),.dout(n4476),.clk(gclk));
	jand g3835(.dina(w_n4452_60[2]),.dinb(w_n3067_0[1]),.dout(n4477),.clk(gclk));
	jor g3836(.dina(n4477),.dinb(n4476),.dout(result[8]),.clk(gclk));
	jor g3837(.dina(w_address1_60[1]),.dinb(w_n2972_0[0]),.dout(n4479),.clk(gclk));
	jor g3838(.dina(w_n4452_60[1]),.dinb(w_n2975_0[0]),.dout(n4480),.clk(gclk));
	jand g3839(.dina(n4480),.dinb(n4479),.dout(result[9]),.clk(gclk));
	jor g3840(.dina(w_address1_60[0]),.dinb(w_n2961_0[0]),.dout(n4482),.clk(gclk));
	jor g3841(.dina(w_n4452_60[0]),.dinb(w_n2964_0[0]),.dout(n4483),.clk(gclk));
	jand g3842(.dina(n4483),.dinb(n4482),.dout(result[10]),.clk(gclk));
	jor g3843(.dina(w_address1_59[2]),.dinb(w_n2950_0[0]),.dout(n4485),.clk(gclk));
	jor g3844(.dina(w_n4452_59[2]),.dinb(w_n2953_0[0]),.dout(n4486),.clk(gclk));
	jand g3845(.dina(n4486),.dinb(n4485),.dout(result[11]),.clk(gclk));
	jor g3846(.dina(w_address1_59[1]),.dinb(w_n2939_0[0]),.dout(n4488),.clk(gclk));
	jor g3847(.dina(w_n4452_59[1]),.dinb(w_n2942_0[0]),.dout(n4489),.clk(gclk));
	jand g3848(.dina(n4489),.dinb(n4488),.dout(result[12]),.clk(gclk));
	jor g3849(.dina(w_address1_59[0]),.dinb(w_n2928_0[0]),.dout(n4491),.clk(gclk));
	jor g3850(.dina(w_n4452_59[0]),.dinb(w_n2931_0[0]),.dout(n4492),.clk(gclk));
	jand g3851(.dina(n4492),.dinb(n4491),.dout(result[13]),.clk(gclk));
	jor g3852(.dina(w_address1_58[2]),.dinb(w_n2920_0[0]),.dout(n4494),.clk(gclk));
	jor g3853(.dina(w_n4452_58[2]),.dinb(w_n2924_0[0]),.dout(n4495),.clk(gclk));
	jand g3854(.dina(n4495),.dinb(n4494),.dout(result[14]),.clk(gclk));
	jor g3855(.dina(w_address1_58[1]),.dinb(w_n2912_0[0]),.dout(n4497),.clk(gclk));
	jor g3856(.dina(w_n4452_58[1]),.dinb(w_n2916_0[0]),.dout(n4498),.clk(gclk));
	jand g3857(.dina(n4498),.dinb(n4497),.dout(result[15]),.clk(gclk));
	jor g3858(.dina(w_address1_58[0]),.dinb(w_n2903_0[0]),.dout(n4500),.clk(gclk));
	jor g3859(.dina(w_n4452_58[0]),.dinb(w_n2907_0[0]),.dout(n4501),.clk(gclk));
	jand g3860(.dina(n4501),.dinb(n4500),.dout(result[16]),.clk(gclk));
	jor g3861(.dina(w_address1_57[2]),.dinb(w_n2899_0[1]),.dout(n4503),.clk(gclk));
	jor g3862(.dina(w_n4452_57[2]),.dinb(w_n2896_0[0]),.dout(n4504),.clk(gclk));
	jand g3863(.dina(n4504),.dinb(n4503),.dout(result[17]),.clk(gclk));
	jor g3864(.dina(w_address1_57[1]),.dinb(w_n3095_0[0]),.dout(n4506),.clk(gclk));
	jor g3865(.dina(w_n4452_57[1]),.dinb(w_n3098_0[0]),.dout(n4507),.clk(gclk));
	jand g3866(.dina(n4507),.dinb(n4506),.dout(result[18]),.clk(gclk));
	jor g3867(.dina(w_address1_57[0]),.dinb(w_n2887_0[0]),.dout(n4509),.clk(gclk));
	jor g3868(.dina(w_n4452_57[0]),.dinb(w_n2890_0[0]),.dout(n4510),.clk(gclk));
	jand g3869(.dina(n4510),.dinb(n4509),.dout(result[19]),.clk(gclk));
	jor g3870(.dina(w_address1_56[2]),.dinb(w_n2876_0[0]),.dout(n4512),.clk(gclk));
	jor g3871(.dina(w_n4452_56[2]),.dinb(w_n2879_0[0]),.dout(n4513),.clk(gclk));
	jand g3872(.dina(n4513),.dinb(n4512),.dout(result[20]),.clk(gclk));
	jor g3873(.dina(w_address1_56[1]),.dinb(w_n2865_0[0]),.dout(n4515),.clk(gclk));
	jor g3874(.dina(w_n4452_56[1]),.dinb(w_n2868_0[0]),.dout(n4516),.clk(gclk));
	jand g3875(.dina(n4516),.dinb(n4515),.dout(result[21]),.clk(gclk));
	jor g3876(.dina(w_address1_56[0]),.dinb(w_n2857_0[0]),.dout(n4518),.clk(gclk));
	jor g3877(.dina(w_n4452_56[0]),.dinb(w_n2861_0[0]),.dout(n4519),.clk(gclk));
	jand g3878(.dina(n4519),.dinb(n4518),.dout(result[22]),.clk(gclk));
	jor g3879(.dina(w_address1_55[2]),.dinb(w_n3119_0[0]),.dout(n4521),.clk(gclk));
	jor g3880(.dina(w_n4452_55[2]),.dinb(w_n3122_0[0]),.dout(n4522),.clk(gclk));
	jand g3881(.dina(n4522),.dinb(n4521),.dout(result[23]),.clk(gclk));
	jor g3882(.dina(w_address1_55[1]),.dinb(w_n2848_0[0]),.dout(n4524),.clk(gclk));
	jor g3883(.dina(w_n4452_55[1]),.dinb(w_n2851_0[0]),.dout(n4525),.clk(gclk));
	jand g3884(.dina(n4525),.dinb(n4524),.dout(result[24]),.clk(gclk));
	jor g3885(.dina(w_address1_55[0]),.dinb(w_n2837_0[0]),.dout(n4527),.clk(gclk));
	jor g3886(.dina(w_n4452_55[0]),.dinb(w_n2840_0[0]),.dout(n4528),.clk(gclk));
	jand g3887(.dina(n4528),.dinb(n4527),.dout(result[25]),.clk(gclk));
	jor g3888(.dina(w_address1_54[2]),.dinb(w_n2826_0[0]),.dout(n4530),.clk(gclk));
	jor g3889(.dina(w_n4452_54[2]),.dinb(w_n2829_0[0]),.dout(n4531),.clk(gclk));
	jand g3890(.dina(n4531),.dinb(n4530),.dout(result[26]),.clk(gclk));
	jor g3891(.dina(w_address1_54[1]),.dinb(w_n2815_0[0]),.dout(n4533),.clk(gclk));
	jor g3892(.dina(w_n4452_54[1]),.dinb(w_n2818_0[0]),.dout(n4534),.clk(gclk));
	jand g3893(.dina(n4534),.dinb(n4533),.dout(result[27]),.clk(gclk));
	jor g3894(.dina(w_address1_54[0]),.dinb(w_n2804_0[0]),.dout(n4536),.clk(gclk));
	jor g3895(.dina(w_n4452_54[0]),.dinb(w_n2807_0[0]),.dout(n4537),.clk(gclk));
	jand g3896(.dina(n4537),.dinb(n4536),.dout(result[28]),.clk(gclk));
	jor g3897(.dina(w_address1_53[2]),.dinb(w_n2793_0[0]),.dout(n4539),.clk(gclk));
	jor g3898(.dina(w_n4452_53[2]),.dinb(w_n2796_0[0]),.dout(n4540),.clk(gclk));
	jand g3899(.dina(n4540),.dinb(n4539),.dout(result[29]),.clk(gclk));
	jor g3900(.dina(w_address1_53[1]),.dinb(w_n2785_0[0]),.dout(n4542),.clk(gclk));
	jor g3901(.dina(w_n4452_53[1]),.dinb(w_n2789_0[0]),.dout(n4543),.clk(gclk));
	jand g3902(.dina(n4543),.dinb(n4542),.dout(result[30]),.clk(gclk));
	jor g3903(.dina(w_address1_53[0]),.dinb(w_n3148_0[0]),.dout(n4545),.clk(gclk));
	jor g3904(.dina(w_n4452_53[0]),.dinb(w_n3151_0[0]),.dout(n4546),.clk(gclk));
	jand g3905(.dina(n4546),.dinb(n4545),.dout(result[31]),.clk(gclk));
	jor g3906(.dina(w_address1_52[2]),.dinb(w_n3216_0[0]),.dout(n4548),.clk(gclk));
	jor g3907(.dina(w_n4452_52[2]),.dinb(w_n3213_0[0]),.dout(n4549),.clk(gclk));
	jand g3908(.dina(n4549),.dinb(n4548),.dout(result[32]),.clk(gclk));
	jor g3909(.dina(w_address1_52[1]),.dinb(w_n3194_0[0]),.dout(n4551),.clk(gclk));
	jor g3910(.dina(w_n4452_52[1]),.dinb(w_n3198_0[0]),.dout(n4552),.clk(gclk));
	jand g3911(.dina(n4552),.dinb(n4551),.dout(result[33]),.clk(gclk));
	jor g3912(.dina(w_address1_52[0]),.dinb(w_n3205_0[0]),.dout(n4554),.clk(gclk));
	jor g3913(.dina(w_n4452_52[0]),.dinb(w_n3202_0[0]),.dout(n4555),.clk(gclk));
	jand g3914(.dina(n4555),.dinb(n4554),.dout(result[34]),.clk(gclk));
	jor g3915(.dina(w_address1_51[2]),.dinb(w_n3186_0[0]),.dout(n4557),.clk(gclk));
	jor g3916(.dina(w_n4452_51[2]),.dinb(w_n3190_0[0]),.dout(n4558),.clk(gclk));
	jand g3917(.dina(n4558),.dinb(n4557),.dout(result[35]),.clk(gclk));
	jor g3918(.dina(w_address1_51[1]),.dinb(w_n3222_0[0]),.dout(n4560),.clk(gclk));
	jor g3919(.dina(w_n4452_51[1]),.dinb(w_n3226_0[0]),.dout(n4561),.clk(gclk));
	jand g3920(.dina(n4561),.dinb(n4560),.dout(result[36]),.clk(gclk));
	jor g3921(.dina(w_address1_51[0]),.dinb(w_n3159_0[0]),.dout(n4563),.clk(gclk));
	jor g3922(.dina(w_n4452_51[0]),.dinb(w_n3163_0[0]),.dout(n4564),.clk(gclk));
	jand g3923(.dina(n4564),.dinb(n4563),.dout(result[37]),.clk(gclk));
	jor g3924(.dina(w_address1_50[2]),.dinb(w_n3178_0[0]),.dout(n4566),.clk(gclk));
	jor g3925(.dina(w_n4452_50[2]),.dinb(w_n3175_0[0]),.dout(n4567),.clk(gclk));
	jand g3926(.dina(n4567),.dinb(n4566),.dout(result[38]),.clk(gclk));
	jor g3927(.dina(w_address1_50[1]),.dinb(w_n3167_0[0]),.dout(n4569),.clk(gclk));
	jor g3928(.dina(w_n4452_50[1]),.dinb(w_n3171_0[0]),.dout(n4570),.clk(gclk));
	jand g3929(.dina(n4570),.dinb(n4569),.dout(result[39]),.clk(gclk));
	jor g3930(.dina(w_address1_50[0]),.dinb(w_n3310_0[0]),.dout(n4572),.clk(gclk));
	jor g3931(.dina(w_n4452_50[0]),.dinb(w_n3314_0[0]),.dout(n4573),.clk(gclk));
	jand g3932(.dina(n4573),.dinb(n4572),.dout(result[40]),.clk(gclk));
	jor g3933(.dina(w_address1_49[2]),.dinb(w_n3318_0[0]),.dout(n4575),.clk(gclk));
	jor g3934(.dina(w_n4452_49[2]),.dinb(w_n3322_0[0]),.dout(n4576),.clk(gclk));
	jand g3935(.dina(n4576),.dinb(n4575),.dout(result[41]),.clk(gclk));
	jor g3936(.dina(w_address1_49[1]),.dinb(w_n3293_0[0]),.dout(n4578),.clk(gclk));
	jor g3937(.dina(w_n4452_49[1]),.dinb(w_n3297_0[0]),.dout(n4579),.clk(gclk));
	jand g3938(.dina(n4579),.dinb(n4578),.dout(result[42]),.clk(gclk));
	jor g3939(.dina(w_address1_49[0]),.dinb(w_n3285_0[0]),.dout(n4581),.clk(gclk));
	jor g3940(.dina(w_n4452_49[0]),.dinb(w_n3289_0[0]),.dout(n4582),.clk(gclk));
	jand g3941(.dina(n4582),.dinb(n4581),.dout(result[43]),.clk(gclk));
	jor g3942(.dina(w_address1_48[2]),.dinb(w_n3302_0[0]),.dout(n4584),.clk(gclk));
	jor g3943(.dina(w_n4452_48[2]),.dinb(w_n3306_0[0]),.dout(n4585),.clk(gclk));
	jand g3944(.dina(n4585),.dinb(n4584),.dout(result[44]),.clk(gclk));
	jor g3945(.dina(w_address1_48[1]),.dinb(w_n3259_0[0]),.dout(n4587),.clk(gclk));
	jor g3946(.dina(w_n4452_48[1]),.dinb(w_n3263_0[0]),.dout(n4588),.clk(gclk));
	jand g3947(.dina(n4588),.dinb(n4587),.dout(result[45]),.clk(gclk));
	jor g3948(.dina(w_address1_48[0]),.dinb(w_n3278_0[0]),.dout(n4590),.clk(gclk));
	jor g3949(.dina(w_n4452_48[0]),.dinb(w_n3275_0[0]),.dout(n4591),.clk(gclk));
	jand g3950(.dina(n4591),.dinb(n4590),.dout(result[46]),.clk(gclk));
	jor g3951(.dina(w_address1_47[2]),.dinb(w_n3267_0[0]),.dout(n4593),.clk(gclk));
	jor g3952(.dina(w_n4452_47[2]),.dinb(w_n3271_0[0]),.dout(n4594),.clk(gclk));
	jand g3953(.dina(n4594),.dinb(n4593),.dout(result[47]),.clk(gclk));
	jor g3954(.dina(w_address1_47[1]),.dinb(w_n3418_0[0]),.dout(n4596),.clk(gclk));
	jor g3955(.dina(w_n4452_47[1]),.dinb(w_n3415_0[0]),.dout(n4597),.clk(gclk));
	jand g3956(.dina(n4597),.dinb(n4596),.dout(result[48]),.clk(gclk));
	jor g3957(.dina(w_address1_47[0]),.dinb(w_n3360_0[0]),.dout(n4599),.clk(gclk));
	jor g3958(.dina(w_n4452_47[0]),.dinb(w_n3364_0[0]),.dout(n4600),.clk(gclk));
	jand g3959(.dina(n4600),.dinb(n4599),.dout(result[49]),.clk(gclk));
	jor g3960(.dina(w_address1_46[2]),.dinb(w_n3371_0[0]),.dout(n4602),.clk(gclk));
	jor g3961(.dina(w_n4452_46[2]),.dinb(w_n3368_0[0]),.dout(n4603),.clk(gclk));
	jand g3962(.dina(n4603),.dinb(n4602),.dout(result[50]),.clk(gclk));
	jor g3963(.dina(w_address1_46[1]),.dinb(w_n3352_0[0]),.dout(n4605),.clk(gclk));
	jor g3964(.dina(w_n4452_46[1]),.dinb(w_n3356_0[0]),.dout(n4606),.clk(gclk));
	jand g3965(.dina(n4606),.dinb(n4605),.dout(result[51]),.clk(gclk));
	jor g3966(.dina(w_address1_46[0]),.dinb(w_n3387_0[0]),.dout(n4608),.clk(gclk));
	jor g3967(.dina(w_n4452_46[0]),.dinb(w_n3391_0[0]),.dout(n4609),.clk(gclk));
	jand g3968(.dina(n4609),.dinb(n4608),.dout(result[52]),.clk(gclk));
	jor g3969(.dina(w_address1_45[2]),.dinb(w_n3378_0[0]),.dout(n4611),.clk(gclk));
	jor g3970(.dina(w_n4452_45[2]),.dinb(w_n3382_0[0]),.dout(n4612),.clk(gclk));
	jand g3971(.dina(n4612),.dinb(n4611),.dout(result[53]),.clk(gclk));
	jor g3972(.dina(w_address1_45[1]),.dinb(w_n3409_0[0]),.dout(n4614),.clk(gclk));
	jor g3973(.dina(w_n4452_45[1]),.dinb(w_n3406_0[0]),.dout(n4615),.clk(gclk));
	jand g3974(.dina(n4615),.dinb(n4614),.dout(result[54]),.clk(gclk));
	jor g3975(.dina(w_address1_45[0]),.dinb(w_n3398_0[0]),.dout(n4617),.clk(gclk));
	jor g3976(.dina(w_n4452_45[0]),.dinb(w_n3402_0[0]),.dout(n4618),.clk(gclk));
	jand g3977(.dina(n4618),.dinb(n4617),.dout(result[55]),.clk(gclk));
	jor g3978(.dina(w_address1_44[2]),.dinb(w_n3499_0[0]),.dout(n4620),.clk(gclk));
	jor g3979(.dina(w_n4452_44[2]),.dinb(w_n3503_0[0]),.dout(n4621),.clk(gclk));
	jand g3980(.dina(n4621),.dinb(n4620),.dout(result[56]),.clk(gclk));
	jor g3981(.dina(w_address1_44[1]),.dinb(w_n3507_0[0]),.dout(n4623),.clk(gclk));
	jor g3982(.dina(w_n4452_44[1]),.dinb(w_n3511_0[0]),.dout(n4624),.clk(gclk));
	jand g3983(.dina(n4624),.dinb(n4623),.dout(result[57]),.clk(gclk));
	jor g3984(.dina(w_address1_44[0]),.dinb(w_n3482_0[0]),.dout(n4626),.clk(gclk));
	jor g3985(.dina(w_n4452_44[0]),.dinb(w_n3486_0[0]),.dout(n4627),.clk(gclk));
	jand g3986(.dina(n4627),.dinb(n4626),.dout(result[58]),.clk(gclk));
	jor g3987(.dina(w_address1_43[2]),.dinb(w_n3474_0[0]),.dout(n4629),.clk(gclk));
	jor g3988(.dina(w_n4452_43[2]),.dinb(w_n3478_0[0]),.dout(n4630),.clk(gclk));
	jand g3989(.dina(n4630),.dinb(n4629),.dout(result[59]),.clk(gclk));
	jor g3990(.dina(w_address1_43[1]),.dinb(w_n3491_0[0]),.dout(n4632),.clk(gclk));
	jor g3991(.dina(w_n4452_43[1]),.dinb(w_n3495_0[0]),.dout(n4633),.clk(gclk));
	jand g3992(.dina(n4633),.dinb(n4632),.dout(result[60]),.clk(gclk));
	jor g3993(.dina(w_address1_43[0]),.dinb(w_n3448_0[0]),.dout(n4635),.clk(gclk));
	jor g3994(.dina(w_n4452_43[0]),.dinb(w_n3452_0[0]),.dout(n4636),.clk(gclk));
	jand g3995(.dina(n4636),.dinb(n4635),.dout(result[61]),.clk(gclk));
	jor g3996(.dina(w_address1_42[2]),.dinb(w_n3467_0[0]),.dout(n4638),.clk(gclk));
	jor g3997(.dina(w_n4452_42[2]),.dinb(w_n3464_0[0]),.dout(n4639),.clk(gclk));
	jand g3998(.dina(n4639),.dinb(n4638),.dout(result[62]),.clk(gclk));
	jor g3999(.dina(w_address1_42[1]),.dinb(w_n3456_0[0]),.dout(n4641),.clk(gclk));
	jor g4000(.dina(w_n4452_42[1]),.dinb(w_n3460_0[0]),.dout(n4642),.clk(gclk));
	jand g4001(.dina(n4642),.dinb(n4641),.dout(result[63]),.clk(gclk));
	jor g4002(.dina(w_address1_42[0]),.dinb(w_n3569_0[0]),.dout(n4644),.clk(gclk));
	jor g4003(.dina(w_n4452_42[0]),.dinb(w_n3566_0[0]),.dout(n4645),.clk(gclk));
	jand g4004(.dina(n4645),.dinb(n4644),.dout(result[64]),.clk(gclk));
	jor g4005(.dina(w_address1_41[2]),.dinb(w_n3558_0[0]),.dout(n4647),.clk(gclk));
	jor g4006(.dina(w_n4452_41[2]),.dinb(w_n3562_0[0]),.dout(n4648),.clk(gclk));
	jand g4007(.dina(n4648),.dinb(n4647),.dout(result[65]),.clk(gclk));
	jor g4008(.dina(w_address1_41[1]),.dinb(w_n3552_0[0]),.dout(n4650),.clk(gclk));
	jor g4009(.dina(w_n4452_41[1]),.dinb(w_n3549_0[0]),.dout(n4651),.clk(gclk));
	jand g4010(.dina(n4651),.dinb(n4650),.dout(result[66]),.clk(gclk));
	jor g4011(.dina(w_address1_41[0]),.dinb(w_n3541_0[0]),.dout(n4653),.clk(gclk));
	jor g4012(.dina(w_n4452_41[0]),.dinb(w_n3545_0[0]),.dout(n4654),.clk(gclk));
	jand g4013(.dina(n4654),.dinb(n4653),.dout(result[67]),.clk(gclk));
	jor g4014(.dina(w_address1_40[2]),.dinb(w_n3587_0[0]),.dout(n4656),.clk(gclk));
	jor g4015(.dina(w_n4452_40[2]),.dinb(w_n3591_0[0]),.dout(n4657),.clk(gclk));
	jand g4016(.dina(n4657),.dinb(n4656),.dout(result[68]),.clk(gclk));
	jor g4017(.dina(w_address1_40[1]),.dinb(w_n3595_0[0]),.dout(n4659),.clk(gclk));
	jor g4018(.dina(w_n4452_40[1]),.dinb(w_n3599_0[0]),.dout(n4660),.clk(gclk));
	jand g4019(.dina(n4660),.dinb(n4659),.dout(result[69]),.clk(gclk));
	jor g4020(.dina(w_address1_40[0]),.dinb(w_n3614_0[0]),.dout(n4662),.clk(gclk));
	jor g4021(.dina(w_n4452_40[0]),.dinb(w_n3611_0[0]),.dout(n4663),.clk(gclk));
	jand g4022(.dina(n4663),.dinb(n4662),.dout(result[70]),.clk(gclk));
	jor g4023(.dina(w_address1_39[2]),.dinb(w_n3603_0[0]),.dout(n4665),.clk(gclk));
	jor g4024(.dina(w_n4452_39[2]),.dinb(w_n3607_0[0]),.dout(n4666),.clk(gclk));
	jand g4025(.dina(n4666),.dinb(n4665),.dout(result[71]),.clk(gclk));
	jor g4026(.dina(w_address1_39[1]),.dinb(w_n3661_0[0]),.dout(n4668),.clk(gclk));
	jor g4027(.dina(w_n4452_39[1]),.dinb(w_n3658_0[0]),.dout(n4669),.clk(gclk));
	jand g4028(.dina(n4669),.dinb(n4668),.dout(result[72]),.clk(gclk));
	jor g4029(.dina(w_address1_39[0]),.dinb(w_n3650_0[0]),.dout(n4671),.clk(gclk));
	jor g4030(.dina(w_n4452_39[0]),.dinb(w_n3654_0[0]),.dout(n4672),.clk(gclk));
	jand g4031(.dina(n4672),.dinb(n4671),.dout(result[73]),.clk(gclk));
	jor g4032(.dina(w_address1_38[2]),.dinb(w_n3644_0[0]),.dout(n4674),.clk(gclk));
	jor g4033(.dina(w_n4452_38[2]),.dinb(w_n3641_0[0]),.dout(n4675),.clk(gclk));
	jand g4034(.dina(n4675),.dinb(n4674),.dout(result[74]),.clk(gclk));
	jor g4035(.dina(w_address1_38[1]),.dinb(w_n3633_0[0]),.dout(n4677),.clk(gclk));
	jor g4036(.dina(w_n4452_38[1]),.dinb(w_n3637_0[0]),.dout(n4678),.clk(gclk));
	jand g4037(.dina(n4678),.dinb(n4677),.dout(result[75]),.clk(gclk));
	jor g4038(.dina(w_address1_38[0]),.dinb(w_n3679_0[0]),.dout(n4680),.clk(gclk));
	jor g4039(.dina(w_n4452_38[0]),.dinb(w_n3683_0[0]),.dout(n4681),.clk(gclk));
	jand g4040(.dina(n4681),.dinb(n4680),.dout(result[76]),.clk(gclk));
	jor g4041(.dina(w_address1_37[2]),.dinb(w_n3687_0[0]),.dout(n4683),.clk(gclk));
	jor g4042(.dina(w_n4452_37[2]),.dinb(w_n3691_0[0]),.dout(n4684),.clk(gclk));
	jand g4043(.dina(n4684),.dinb(n4683),.dout(result[77]),.clk(gclk));
	jor g4044(.dina(w_address1_37[1]),.dinb(w_n3706_0[0]),.dout(n4686),.clk(gclk));
	jor g4045(.dina(w_n4452_37[1]),.dinb(w_n3703_0[0]),.dout(n4687),.clk(gclk));
	jand g4046(.dina(n4687),.dinb(n4686),.dout(result[78]),.clk(gclk));
	jor g4047(.dina(w_address1_37[0]),.dinb(w_n3695_0[0]),.dout(n4689),.clk(gclk));
	jor g4048(.dina(w_n4452_37[0]),.dinb(w_n3699_0[0]),.dout(n4690),.clk(gclk));
	jand g4049(.dina(n4690),.dinb(n4689),.dout(result[79]),.clk(gclk));
	jor g4050(.dina(w_address1_36[2]),.dinb(w_n3753_0[0]),.dout(n4692),.clk(gclk));
	jor g4051(.dina(w_n4452_36[2]),.dinb(w_n3750_0[0]),.dout(n4693),.clk(gclk));
	jand g4052(.dina(n4693),.dinb(n4692),.dout(result[80]),.clk(gclk));
	jor g4053(.dina(w_address1_36[1]),.dinb(w_n3742_0[0]),.dout(n4695),.clk(gclk));
	jor g4054(.dina(w_n4452_36[1]),.dinb(w_n3746_0[0]),.dout(n4696),.clk(gclk));
	jand g4055(.dina(n4696),.dinb(n4695),.dout(result[81]),.clk(gclk));
	jor g4056(.dina(w_address1_36[0]),.dinb(w_n3736_0[0]),.dout(n4698),.clk(gclk));
	jor g4057(.dina(w_n4452_36[0]),.dinb(w_n3733_0[0]),.dout(n4699),.clk(gclk));
	jand g4058(.dina(n4699),.dinb(n4698),.dout(result[82]),.clk(gclk));
	jor g4059(.dina(w_address1_35[2]),.dinb(w_n3725_0[0]),.dout(n4701),.clk(gclk));
	jor g4060(.dina(w_n4452_35[2]),.dinb(w_n3729_0[0]),.dout(n4702),.clk(gclk));
	jand g4061(.dina(n4702),.dinb(n4701),.dout(result[83]),.clk(gclk));
	jor g4062(.dina(w_address1_35[1]),.dinb(w_n3771_0[0]),.dout(n4704),.clk(gclk));
	jor g4063(.dina(w_n4452_35[1]),.dinb(w_n3775_0[0]),.dout(n4705),.clk(gclk));
	jand g4064(.dina(n4705),.dinb(n4704),.dout(result[84]),.clk(gclk));
	jor g4065(.dina(w_address1_35[0]),.dinb(w_n3779_0[0]),.dout(n4707),.clk(gclk));
	jor g4066(.dina(w_n4452_35[0]),.dinb(w_n3783_0[0]),.dout(n4708),.clk(gclk));
	jand g4067(.dina(n4708),.dinb(n4707),.dout(result[85]),.clk(gclk));
	jor g4068(.dina(w_address1_34[2]),.dinb(w_n3798_0[0]),.dout(n4710),.clk(gclk));
	jor g4069(.dina(w_n4452_34[2]),.dinb(w_n3795_0[0]),.dout(n4711),.clk(gclk));
	jand g4070(.dina(n4711),.dinb(n4710),.dout(result[86]),.clk(gclk));
	jor g4071(.dina(w_address1_34[1]),.dinb(w_n3787_0[0]),.dout(n4713),.clk(gclk));
	jor g4072(.dina(w_n4452_34[1]),.dinb(w_n3791_0[0]),.dout(n4714),.clk(gclk));
	jand g4073(.dina(n4714),.dinb(n4713),.dout(result[87]),.clk(gclk));
	jor g4074(.dina(w_address1_34[0]),.dinb(w_n3845_0[0]),.dout(n4716),.clk(gclk));
	jor g4075(.dina(w_n4452_34[0]),.dinb(w_n3842_0[0]),.dout(n4717),.clk(gclk));
	jand g4076(.dina(n4717),.dinb(n4716),.dout(result[88]),.clk(gclk));
	jor g4077(.dina(w_address1_33[2]),.dinb(w_n3834_0[0]),.dout(n4719),.clk(gclk));
	jor g4078(.dina(w_n4452_33[2]),.dinb(w_n3838_0[0]),.dout(n4720),.clk(gclk));
	jand g4079(.dina(n4720),.dinb(n4719),.dout(result[89]),.clk(gclk));
	jor g4080(.dina(w_address1_33[1]),.dinb(w_n3828_0[0]),.dout(n4722),.clk(gclk));
	jor g4081(.dina(w_n4452_33[1]),.dinb(w_n3825_0[0]),.dout(n4723),.clk(gclk));
	jand g4082(.dina(n4723),.dinb(n4722),.dout(result[90]),.clk(gclk));
	jor g4083(.dina(w_address1_33[0]),.dinb(w_n3817_0[0]),.dout(n4725),.clk(gclk));
	jor g4084(.dina(w_n4452_33[0]),.dinb(w_n3821_0[0]),.dout(n4726),.clk(gclk));
	jand g4085(.dina(n4726),.dinb(n4725),.dout(result[91]),.clk(gclk));
	jor g4086(.dina(w_address1_32[2]),.dinb(w_n3863_0[0]),.dout(n4728),.clk(gclk));
	jor g4087(.dina(w_n4452_32[2]),.dinb(w_n3867_0[0]),.dout(n4729),.clk(gclk));
	jand g4088(.dina(n4729),.dinb(n4728),.dout(result[92]),.clk(gclk));
	jor g4089(.dina(w_address1_32[1]),.dinb(w_n3871_0[0]),.dout(n4731),.clk(gclk));
	jor g4090(.dina(w_n4452_32[1]),.dinb(w_n3875_0[0]),.dout(n4732),.clk(gclk));
	jand g4091(.dina(n4732),.dinb(n4731),.dout(result[93]),.clk(gclk));
	jor g4092(.dina(w_address1_32[0]),.dinb(w_n3890_0[0]),.dout(n4734),.clk(gclk));
	jor g4093(.dina(w_n4452_32[0]),.dinb(w_n3887_0[0]),.dout(n4735),.clk(gclk));
	jand g4094(.dina(n4735),.dinb(n4734),.dout(result[94]),.clk(gclk));
	jor g4095(.dina(w_address1_31[2]),.dinb(w_n3879_0[0]),.dout(n4737),.clk(gclk));
	jor g4096(.dina(w_n4452_31[2]),.dinb(w_n3883_0[0]),.dout(n4738),.clk(gclk));
	jand g4097(.dina(n4738),.dinb(n4737),.dout(result[95]),.clk(gclk));
	jor g4098(.dina(w_address1_31[1]),.dinb(w_n3937_0[0]),.dout(n4740),.clk(gclk));
	jor g4099(.dina(w_n4452_31[1]),.dinb(w_n3934_0[0]),.dout(n4741),.clk(gclk));
	jand g4100(.dina(n4741),.dinb(n4740),.dout(result[96]),.clk(gclk));
	jor g4101(.dina(w_address1_31[0]),.dinb(w_n3926_0[0]),.dout(n4743),.clk(gclk));
	jor g4102(.dina(w_n4452_31[0]),.dinb(w_n3930_0[0]),.dout(n4744),.clk(gclk));
	jand g4103(.dina(n4744),.dinb(n4743),.dout(result[97]),.clk(gclk));
	jor g4104(.dina(w_address1_30[2]),.dinb(w_n3920_0[0]),.dout(n4746),.clk(gclk));
	jor g4105(.dina(w_n4452_30[2]),.dinb(w_n3917_0[0]),.dout(n4747),.clk(gclk));
	jand g4106(.dina(n4747),.dinb(n4746),.dout(result[98]),.clk(gclk));
	jor g4107(.dina(w_address1_30[1]),.dinb(w_n3909_0[0]),.dout(n4749),.clk(gclk));
	jor g4108(.dina(w_n4452_30[1]),.dinb(w_n3913_0[0]),.dout(n4750),.clk(gclk));
	jand g4109(.dina(n4750),.dinb(n4749),.dout(result[99]),.clk(gclk));
	jor g4110(.dina(w_address1_30[0]),.dinb(w_n3955_0[0]),.dout(n4752),.clk(gclk));
	jor g4111(.dina(w_n4452_30[0]),.dinb(w_n3959_0[0]),.dout(n4753),.clk(gclk));
	jand g4112(.dina(n4753),.dinb(n4752),.dout(result[100]),.clk(gclk));
	jor g4113(.dina(w_address1_29[2]),.dinb(w_n3963_0[0]),.dout(n4755),.clk(gclk));
	jor g4114(.dina(w_n4452_29[2]),.dinb(w_n3967_0[0]),.dout(n4756),.clk(gclk));
	jand g4115(.dina(n4756),.dinb(n4755),.dout(result[101]),.clk(gclk));
	jor g4116(.dina(w_address1_29[1]),.dinb(w_n3982_0[0]),.dout(n4758),.clk(gclk));
	jor g4117(.dina(w_n4452_29[1]),.dinb(w_n3979_0[0]),.dout(n4759),.clk(gclk));
	jand g4118(.dina(n4759),.dinb(n4758),.dout(result[102]),.clk(gclk));
	jor g4119(.dina(w_address1_29[0]),.dinb(w_n3971_0[0]),.dout(n4761),.clk(gclk));
	jor g4120(.dina(w_n4452_29[0]),.dinb(w_n3975_0[0]),.dout(n4762),.clk(gclk));
	jand g4121(.dina(n4762),.dinb(n4761),.dout(result[103]),.clk(gclk));
	jor g4122(.dina(w_address1_28[2]),.dinb(w_n4029_0[0]),.dout(n4764),.clk(gclk));
	jor g4123(.dina(w_n4452_28[2]),.dinb(w_n4026_0[0]),.dout(n4765),.clk(gclk));
	jand g4124(.dina(n4765),.dinb(n4764),.dout(result[104]),.clk(gclk));
	jor g4125(.dina(w_address1_28[1]),.dinb(w_n4018_0[0]),.dout(n4767),.clk(gclk));
	jor g4126(.dina(w_n4452_28[1]),.dinb(w_n4022_0[0]),.dout(n4768),.clk(gclk));
	jand g4127(.dina(n4768),.dinb(n4767),.dout(result[105]),.clk(gclk));
	jor g4128(.dina(w_address1_28[0]),.dinb(w_n4012_0[0]),.dout(n4770),.clk(gclk));
	jor g4129(.dina(w_n4452_28[0]),.dinb(w_n4009_0[0]),.dout(n4771),.clk(gclk));
	jand g4130(.dina(n4771),.dinb(n4770),.dout(result[106]),.clk(gclk));
	jor g4131(.dina(w_address1_27[2]),.dinb(w_n4001_0[0]),.dout(n4773),.clk(gclk));
	jor g4132(.dina(w_n4452_27[2]),.dinb(w_n4005_0[0]),.dout(n4774),.clk(gclk));
	jand g4133(.dina(n4774),.dinb(n4773),.dout(result[107]),.clk(gclk));
	jor g4134(.dina(w_address1_27[1]),.dinb(w_n4047_0[0]),.dout(n4776),.clk(gclk));
	jor g4135(.dina(w_n4452_27[1]),.dinb(w_n4051_0[0]),.dout(n4777),.clk(gclk));
	jand g4136(.dina(n4777),.dinb(n4776),.dout(result[108]),.clk(gclk));
	jor g4137(.dina(w_address1_27[0]),.dinb(w_n4055_0[0]),.dout(n4779),.clk(gclk));
	jor g4138(.dina(w_n4452_27[0]),.dinb(w_n4059_0[0]),.dout(n4780),.clk(gclk));
	jand g4139(.dina(n4780),.dinb(n4779),.dout(result[109]),.clk(gclk));
	jor g4140(.dina(w_address1_26[2]),.dinb(w_n4074_0[0]),.dout(n4782),.clk(gclk));
	jor g4141(.dina(w_n4452_26[2]),.dinb(w_n4071_0[0]),.dout(n4783),.clk(gclk));
	jand g4142(.dina(n4783),.dinb(n4782),.dout(result[110]),.clk(gclk));
	jor g4143(.dina(w_address1_26[1]),.dinb(w_n4063_0[0]),.dout(n4785),.clk(gclk));
	jor g4144(.dina(w_n4452_26[1]),.dinb(w_n4067_0[0]),.dout(n4786),.clk(gclk));
	jand g4145(.dina(n4786),.dinb(n4785),.dout(result[111]),.clk(gclk));
	jor g4146(.dina(w_address1_26[0]),.dinb(w_n4121_0[0]),.dout(n4788),.clk(gclk));
	jor g4147(.dina(w_n4452_26[0]),.dinb(w_n4118_0[0]),.dout(n4789),.clk(gclk));
	jand g4148(.dina(n4789),.dinb(n4788),.dout(result[112]),.clk(gclk));
	jor g4149(.dina(w_address1_25[2]),.dinb(w_n4110_0[0]),.dout(n4791),.clk(gclk));
	jor g4150(.dina(w_n4452_25[2]),.dinb(w_n4114_0[0]),.dout(n4792),.clk(gclk));
	jand g4151(.dina(n4792),.dinb(n4791),.dout(result[113]),.clk(gclk));
	jor g4152(.dina(w_address1_25[1]),.dinb(w_n4104_0[0]),.dout(n4794),.clk(gclk));
	jor g4153(.dina(w_n4452_25[1]),.dinb(w_n4101_0[0]),.dout(n4795),.clk(gclk));
	jand g4154(.dina(n4795),.dinb(n4794),.dout(result[114]),.clk(gclk));
	jor g4155(.dina(w_address1_25[0]),.dinb(w_n4093_0[0]),.dout(n4797),.clk(gclk));
	jor g4156(.dina(w_n4452_25[0]),.dinb(w_n4097_0[0]),.dout(n4798),.clk(gclk));
	jand g4157(.dina(n4798),.dinb(n4797),.dout(result[115]),.clk(gclk));
	jor g4158(.dina(w_address1_24[2]),.dinb(w_n4139_0[0]),.dout(n4800),.clk(gclk));
	jor g4159(.dina(w_n4452_24[2]),.dinb(w_n4143_0[0]),.dout(n4801),.clk(gclk));
	jand g4160(.dina(n4801),.dinb(n4800),.dout(result[116]),.clk(gclk));
	jor g4161(.dina(w_address1_24[1]),.dinb(w_n4147_0[0]),.dout(n4803),.clk(gclk));
	jor g4162(.dina(w_n4452_24[1]),.dinb(w_n4151_0[0]),.dout(n4804),.clk(gclk));
	jand g4163(.dina(n4804),.dinb(n4803),.dout(result[117]),.clk(gclk));
	jor g4164(.dina(w_address1_24[0]),.dinb(w_n4166_0[0]),.dout(n4806),.clk(gclk));
	jor g4165(.dina(w_n4452_24[0]),.dinb(w_n4163_0[0]),.dout(n4807),.clk(gclk));
	jand g4166(.dina(n4807),.dinb(n4806),.dout(result[118]),.clk(gclk));
	jor g4167(.dina(w_address1_23[2]),.dinb(w_n4155_0[0]),.dout(n4809),.clk(gclk));
	jor g4168(.dina(w_n4452_23[2]),.dinb(w_n4159_0[0]),.dout(n4810),.clk(gclk));
	jand g4169(.dina(n4810),.dinb(n4809),.dout(result[119]),.clk(gclk));
	jor g4170(.dina(w_address1_23[1]),.dinb(w_n4213_0[0]),.dout(n4812),.clk(gclk));
	jor g4171(.dina(w_n4452_23[1]),.dinb(w_n4210_0[0]),.dout(n4813),.clk(gclk));
	jand g4172(.dina(n4813),.dinb(n4812),.dout(result[120]),.clk(gclk));
	jor g4173(.dina(w_address1_23[0]),.dinb(w_n4202_0[0]),.dout(n4815),.clk(gclk));
	jor g4174(.dina(w_n4452_23[0]),.dinb(w_n4206_0[0]),.dout(n4816),.clk(gclk));
	jand g4175(.dina(n4816),.dinb(n4815),.dout(result[121]),.clk(gclk));
	jor g4176(.dina(w_address1_22[2]),.dinb(w_n4196_0[0]),.dout(n4818),.clk(gclk));
	jor g4177(.dina(w_n4452_22[2]),.dinb(w_n4193_0[0]),.dout(n4819),.clk(gclk));
	jand g4178(.dina(n4819),.dinb(n4818),.dout(result[122]),.clk(gclk));
	jor g4179(.dina(w_address1_22[1]),.dinb(w_n4185_0[0]),.dout(n4821),.clk(gclk));
	jor g4180(.dina(w_n4452_22[1]),.dinb(w_n4189_0[0]),.dout(n4822),.clk(gclk));
	jand g4181(.dina(n4822),.dinb(n4821),.dout(result[123]),.clk(gclk));
	jor g4182(.dina(w_address1_22[0]),.dinb(w_n4252_0[0]),.dout(n4824),.clk(gclk));
	jor g4183(.dina(w_n4452_22[0]),.dinb(w_n4256_0[0]),.dout(n4825),.clk(gclk));
	jand g4184(.dina(n4825),.dinb(n4824),.dout(result[124]),.clk(gclk));
	jor g4185(.dina(w_address1_21[2]),.dinb(w_n4239_0[0]),.dout(n4827),.clk(gclk));
	jor g4186(.dina(w_n4452_21[2]),.dinb(w_n4243_0[0]),.dout(n4828),.clk(gclk));
	jand g4187(.dina(n4828),.dinb(n4827),.dout(result[125]),.clk(gclk));
	jor g4188(.dina(w_address1_21[1]),.dinb(w_n4231_0[0]),.dout(n4830),.clk(gclk));
	jor g4189(.dina(w_n4452_21[1]),.dinb(w_n4235_0[0]),.dout(n4831),.clk(gclk));
	jand g4190(.dina(n4831),.dinb(n4830),.dout(result[126]),.clk(gclk));
	jand g4191(.dina(w_n4248_0[0]),.dinb(w_n4246_0[0]),.dout(result[127]),.clk(gclk));
	jor g4192(.dina(w_address1_21[0]),.dinb(w_n2783_21[1]),.dout(n4834),.clk(gclk));
	jor g4193(.dina(w_n4452_21[0]),.dinb(w_n1711_21[1]),.dout(n4835),.clk(gclk));
	jand g4194(.dina(n4835),.dinb(n4834),.dout(address_fa_1),.clk(gclk));
	jspl3 jspl3_w_in00_0(.douta(w_in00_0[0]),.doutb(w_in00_0[1]),.doutc(w_in00_0[2]),.din(in0[0]));
	jspl3 jspl3_w_in01_0(.douta(w_in01_0[0]),.doutb(w_in01_0[1]),.doutc(w_in01_0[2]),.din(in0[1]));
	jspl jspl_w_in01_1(.douta(w_in01_1[0]),.doutb(w_in01_1[1]),.din(w_in01_0[0]));
	jspl3 jspl3_w_in02_0(.douta(w_in02_0[0]),.doutb(w_in02_0[1]),.doutc(w_in02_0[2]),.din(in0[2]));
	jspl3 jspl3_w_in03_0(.douta(w_in03_0[0]),.doutb(w_in03_0[1]),.doutc(w_in03_0[2]),.din(in0[3]));
	jspl3 jspl3_w_in04_0(.douta(w_in04_0[0]),.doutb(w_in04_0[1]),.doutc(w_in04_0[2]),.din(in0[4]));
	jspl3 jspl3_w_in05_0(.douta(w_in05_0[0]),.doutb(w_in05_0[1]),.doutc(w_in05_0[2]),.din(in0[5]));
	jspl3 jspl3_w_in06_0(.douta(w_in06_0[0]),.doutb(w_in06_0[1]),.doutc(w_in06_0[2]),.din(in0[6]));
	jspl3 jspl3_w_in07_0(.douta(w_in07_0[0]),.doutb(w_in07_0[1]),.doutc(w_in07_0[2]),.din(in0[7]));
	jspl3 jspl3_w_in08_0(.douta(w_in08_0[0]),.doutb(w_in08_0[1]),.doutc(w_in08_0[2]),.din(in0[8]));
	jspl3 jspl3_w_in09_0(.douta(w_in09_0[0]),.doutb(w_in09_0[1]),.doutc(w_in09_0[2]),.din(in0[9]));
	jspl3 jspl3_w_in010_0(.douta(w_in010_0[0]),.doutb(w_in010_0[1]),.doutc(w_in010_0[2]),.din(in0[10]));
	jspl3 jspl3_w_in011_0(.douta(w_in011_0[0]),.doutb(w_in011_0[1]),.doutc(w_in011_0[2]),.din(in0[11]));
	jspl3 jspl3_w_in012_0(.douta(w_in012_0[0]),.doutb(w_in012_0[1]),.doutc(w_in012_0[2]),.din(in0[12]));
	jspl3 jspl3_w_in013_0(.douta(w_in013_0[0]),.doutb(w_in013_0[1]),.doutc(w_in013_0[2]),.din(in0[13]));
	jspl3 jspl3_w_in014_0(.douta(w_in014_0[0]),.doutb(w_in014_0[1]),.doutc(w_in014_0[2]),.din(in0[14]));
	jspl3 jspl3_w_in015_0(.douta(w_in015_0[0]),.doutb(w_in015_0[1]),.doutc(w_in015_0[2]),.din(in0[15]));
	jspl3 jspl3_w_in016_0(.douta(w_in016_0[0]),.doutb(w_in016_0[1]),.doutc(w_in016_0[2]),.din(in0[16]));
	jspl3 jspl3_w_in017_0(.douta(w_in017_0[0]),.doutb(w_in017_0[1]),.doutc(w_in017_0[2]),.din(in0[17]));
	jspl3 jspl3_w_in018_0(.douta(w_in018_0[0]),.doutb(w_in018_0[1]),.doutc(w_in018_0[2]),.din(in0[18]));
	jspl3 jspl3_w_in019_0(.douta(w_in019_0[0]),.doutb(w_in019_0[1]),.doutc(w_in019_0[2]),.din(in0[19]));
	jspl3 jspl3_w_in020_0(.douta(w_in020_0[0]),.doutb(w_in020_0[1]),.doutc(w_in020_0[2]),.din(in0[20]));
	jspl3 jspl3_w_in021_0(.douta(w_in021_0[0]),.doutb(w_in021_0[1]),.doutc(w_in021_0[2]),.din(in0[21]));
	jspl3 jspl3_w_in022_0(.douta(w_in022_0[0]),.doutb(w_in022_0[1]),.doutc(w_in022_0[2]),.din(in0[22]));
	jspl3 jspl3_w_in023_0(.douta(w_in023_0[0]),.doutb(w_in023_0[1]),.doutc(w_in023_0[2]),.din(in0[23]));
	jspl3 jspl3_w_in024_0(.douta(w_in024_0[0]),.doutb(w_in024_0[1]),.doutc(w_in024_0[2]),.din(in0[24]));
	jspl3 jspl3_w_in025_0(.douta(w_in025_0[0]),.doutb(w_in025_0[1]),.doutc(w_in025_0[2]),.din(in0[25]));
	jspl3 jspl3_w_in026_0(.douta(w_in026_0[0]),.doutb(w_in026_0[1]),.doutc(w_in026_0[2]),.din(in0[26]));
	jspl3 jspl3_w_in027_0(.douta(w_in027_0[0]),.doutb(w_in027_0[1]),.doutc(w_in027_0[2]),.din(in0[27]));
	jspl3 jspl3_w_in028_0(.douta(w_in028_0[0]),.doutb(w_in028_0[1]),.doutc(w_in028_0[2]),.din(in0[28]));
	jspl3 jspl3_w_in029_0(.douta(w_in029_0[0]),.doutb(w_in029_0[1]),.doutc(w_in029_0[2]),.din(in0[29]));
	jspl3 jspl3_w_in030_0(.douta(w_in030_0[0]),.doutb(w_in030_0[1]),.doutc(w_in030_0[2]),.din(in0[30]));
	jspl3 jspl3_w_in031_0(.douta(w_in031_0[0]),.doutb(w_in031_0[1]),.doutc(w_in031_0[2]),.din(in0[31]));
	jspl3 jspl3_w_in032_0(.douta(w_in032_0[0]),.doutb(w_in032_0[1]),.doutc(w_in032_0[2]),.din(in0[32]));
	jspl3 jspl3_w_in033_0(.douta(w_in033_0[0]),.doutb(w_in033_0[1]),.doutc(w_in033_0[2]),.din(in0[33]));
	jspl3 jspl3_w_in034_0(.douta(w_in034_0[0]),.doutb(w_in034_0[1]),.doutc(w_in034_0[2]),.din(in0[34]));
	jspl3 jspl3_w_in035_0(.douta(w_in035_0[0]),.doutb(w_in035_0[1]),.doutc(w_in035_0[2]),.din(in0[35]));
	jspl3 jspl3_w_in036_0(.douta(w_in036_0[0]),.doutb(w_in036_0[1]),.doutc(w_in036_0[2]),.din(in0[36]));
	jspl3 jspl3_w_in037_0(.douta(w_in037_0[0]),.doutb(w_in037_0[1]),.doutc(w_in037_0[2]),.din(in0[37]));
	jspl3 jspl3_w_in038_0(.douta(w_in038_0[0]),.doutb(w_in038_0[1]),.doutc(w_in038_0[2]),.din(in0[38]));
	jspl3 jspl3_w_in039_0(.douta(w_in039_0[0]),.doutb(w_in039_0[1]),.doutc(w_in039_0[2]),.din(in0[39]));
	jspl3 jspl3_w_in040_0(.douta(w_in040_0[0]),.doutb(w_in040_0[1]),.doutc(w_in040_0[2]),.din(in0[40]));
	jspl3 jspl3_w_in041_0(.douta(w_in041_0[0]),.doutb(w_in041_0[1]),.doutc(w_in041_0[2]),.din(in0[41]));
	jspl3 jspl3_w_in042_0(.douta(w_in042_0[0]),.doutb(w_in042_0[1]),.doutc(w_in042_0[2]),.din(in0[42]));
	jspl3 jspl3_w_in043_0(.douta(w_in043_0[0]),.doutb(w_in043_0[1]),.doutc(w_in043_0[2]),.din(in0[43]));
	jspl3 jspl3_w_in044_0(.douta(w_in044_0[0]),.doutb(w_in044_0[1]),.doutc(w_in044_0[2]),.din(in0[44]));
	jspl3 jspl3_w_in045_0(.douta(w_in045_0[0]),.doutb(w_in045_0[1]),.doutc(w_in045_0[2]),.din(in0[45]));
	jspl3 jspl3_w_in046_0(.douta(w_in046_0[0]),.doutb(w_in046_0[1]),.doutc(w_in046_0[2]),.din(in0[46]));
	jspl3 jspl3_w_in047_0(.douta(w_in047_0[0]),.doutb(w_in047_0[1]),.doutc(w_in047_0[2]),.din(in0[47]));
	jspl3 jspl3_w_in048_0(.douta(w_in048_0[0]),.doutb(w_in048_0[1]),.doutc(w_in048_0[2]),.din(in0[48]));
	jspl3 jspl3_w_in049_0(.douta(w_in049_0[0]),.doutb(w_in049_0[1]),.doutc(w_in049_0[2]),.din(in0[49]));
	jspl3 jspl3_w_in050_0(.douta(w_in050_0[0]),.doutb(w_in050_0[1]),.doutc(w_in050_0[2]),.din(in0[50]));
	jspl3 jspl3_w_in051_0(.douta(w_in051_0[0]),.doutb(w_in051_0[1]),.doutc(w_in051_0[2]),.din(in0[51]));
	jspl3 jspl3_w_in052_0(.douta(w_in052_0[0]),.doutb(w_in052_0[1]),.doutc(w_in052_0[2]),.din(in0[52]));
	jspl3 jspl3_w_in053_0(.douta(w_in053_0[0]),.doutb(w_in053_0[1]),.doutc(w_in053_0[2]),.din(in0[53]));
	jspl3 jspl3_w_in054_0(.douta(w_in054_0[0]),.doutb(w_in054_0[1]),.doutc(w_in054_0[2]),.din(in0[54]));
	jspl3 jspl3_w_in055_0(.douta(w_in055_0[0]),.doutb(w_in055_0[1]),.doutc(w_in055_0[2]),.din(in0[55]));
	jspl3 jspl3_w_in056_0(.douta(w_in056_0[0]),.doutb(w_in056_0[1]),.doutc(w_in056_0[2]),.din(in0[56]));
	jspl3 jspl3_w_in057_0(.douta(w_in057_0[0]),.doutb(w_in057_0[1]),.doutc(w_in057_0[2]),.din(in0[57]));
	jspl3 jspl3_w_in058_0(.douta(w_in058_0[0]),.doutb(w_in058_0[1]),.doutc(w_in058_0[2]),.din(in0[58]));
	jspl3 jspl3_w_in059_0(.douta(w_in059_0[0]),.doutb(w_in059_0[1]),.doutc(w_in059_0[2]),.din(in0[59]));
	jspl3 jspl3_w_in060_0(.douta(w_in060_0[0]),.doutb(w_in060_0[1]),.doutc(w_in060_0[2]),.din(in0[60]));
	jspl3 jspl3_w_in061_0(.douta(w_in061_0[0]),.doutb(w_in061_0[1]),.doutc(w_in061_0[2]),.din(in0[61]));
	jspl3 jspl3_w_in062_0(.douta(w_in062_0[0]),.doutb(w_in062_0[1]),.doutc(w_in062_0[2]),.din(in0[62]));
	jspl3 jspl3_w_in063_0(.douta(w_in063_0[0]),.doutb(w_in063_0[1]),.doutc(w_in063_0[2]),.din(in0[63]));
	jspl3 jspl3_w_in064_0(.douta(w_in064_0[0]),.doutb(w_in064_0[1]),.doutc(w_in064_0[2]),.din(in0[64]));
	jspl3 jspl3_w_in065_0(.douta(w_in065_0[0]),.doutb(w_in065_0[1]),.doutc(w_in065_0[2]),.din(in0[65]));
	jspl3 jspl3_w_in066_0(.douta(w_in066_0[0]),.doutb(w_in066_0[1]),.doutc(w_in066_0[2]),.din(in0[66]));
	jspl3 jspl3_w_in067_0(.douta(w_in067_0[0]),.doutb(w_in067_0[1]),.doutc(w_in067_0[2]),.din(in0[67]));
	jspl3 jspl3_w_in068_0(.douta(w_in068_0[0]),.doutb(w_in068_0[1]),.doutc(w_in068_0[2]),.din(in0[68]));
	jspl3 jspl3_w_in069_0(.douta(w_in069_0[0]),.doutb(w_in069_0[1]),.doutc(w_in069_0[2]),.din(in0[69]));
	jspl3 jspl3_w_in070_0(.douta(w_in070_0[0]),.doutb(w_in070_0[1]),.doutc(w_in070_0[2]),.din(in0[70]));
	jspl3 jspl3_w_in071_0(.douta(w_in071_0[0]),.doutb(w_in071_0[1]),.doutc(w_in071_0[2]),.din(in0[71]));
	jspl3 jspl3_w_in072_0(.douta(w_in072_0[0]),.doutb(w_in072_0[1]),.doutc(w_in072_0[2]),.din(in0[72]));
	jspl3 jspl3_w_in073_0(.douta(w_in073_0[0]),.doutb(w_in073_0[1]),.doutc(w_in073_0[2]),.din(in0[73]));
	jspl3 jspl3_w_in074_0(.douta(w_in074_0[0]),.doutb(w_in074_0[1]),.doutc(w_in074_0[2]),.din(in0[74]));
	jspl3 jspl3_w_in075_0(.douta(w_in075_0[0]),.doutb(w_in075_0[1]),.doutc(w_in075_0[2]),.din(in0[75]));
	jspl3 jspl3_w_in076_0(.douta(w_in076_0[0]),.doutb(w_in076_0[1]),.doutc(w_in076_0[2]),.din(in0[76]));
	jspl3 jspl3_w_in077_0(.douta(w_in077_0[0]),.doutb(w_in077_0[1]),.doutc(w_in077_0[2]),.din(in0[77]));
	jspl3 jspl3_w_in078_0(.douta(w_in078_0[0]),.doutb(w_in078_0[1]),.doutc(w_in078_0[2]),.din(in0[78]));
	jspl3 jspl3_w_in079_0(.douta(w_in079_0[0]),.doutb(w_in079_0[1]),.doutc(w_in079_0[2]),.din(in0[79]));
	jspl3 jspl3_w_in080_0(.douta(w_in080_0[0]),.doutb(w_in080_0[1]),.doutc(w_in080_0[2]),.din(in0[80]));
	jspl3 jspl3_w_in081_0(.douta(w_in081_0[0]),.doutb(w_in081_0[1]),.doutc(w_in081_0[2]),.din(in0[81]));
	jspl3 jspl3_w_in082_0(.douta(w_in082_0[0]),.doutb(w_in082_0[1]),.doutc(w_in082_0[2]),.din(in0[82]));
	jspl3 jspl3_w_in083_0(.douta(w_in083_0[0]),.doutb(w_in083_0[1]),.doutc(w_in083_0[2]),.din(in0[83]));
	jspl3 jspl3_w_in084_0(.douta(w_in084_0[0]),.doutb(w_in084_0[1]),.doutc(w_in084_0[2]),.din(in0[84]));
	jspl3 jspl3_w_in085_0(.douta(w_in085_0[0]),.doutb(w_in085_0[1]),.doutc(w_in085_0[2]),.din(in0[85]));
	jspl3 jspl3_w_in086_0(.douta(w_in086_0[0]),.doutb(w_in086_0[1]),.doutc(w_in086_0[2]),.din(in0[86]));
	jspl3 jspl3_w_in087_0(.douta(w_in087_0[0]),.doutb(w_in087_0[1]),.doutc(w_in087_0[2]),.din(in0[87]));
	jspl3 jspl3_w_in088_0(.douta(w_in088_0[0]),.doutb(w_in088_0[1]),.doutc(w_in088_0[2]),.din(in0[88]));
	jspl3 jspl3_w_in089_0(.douta(w_in089_0[0]),.doutb(w_in089_0[1]),.doutc(w_in089_0[2]),.din(in0[89]));
	jspl3 jspl3_w_in090_0(.douta(w_in090_0[0]),.doutb(w_in090_0[1]),.doutc(w_in090_0[2]),.din(in0[90]));
	jspl3 jspl3_w_in091_0(.douta(w_in091_0[0]),.doutb(w_in091_0[1]),.doutc(w_in091_0[2]),.din(in0[91]));
	jspl3 jspl3_w_in092_0(.douta(w_in092_0[0]),.doutb(w_in092_0[1]),.doutc(w_in092_0[2]),.din(in0[92]));
	jspl3 jspl3_w_in093_0(.douta(w_in093_0[0]),.doutb(w_in093_0[1]),.doutc(w_in093_0[2]),.din(in0[93]));
	jspl3 jspl3_w_in094_0(.douta(w_in094_0[0]),.doutb(w_in094_0[1]),.doutc(w_in094_0[2]),.din(in0[94]));
	jspl3 jspl3_w_in095_0(.douta(w_in095_0[0]),.doutb(w_in095_0[1]),.doutc(w_in095_0[2]),.din(in0[95]));
	jspl3 jspl3_w_in096_0(.douta(w_in096_0[0]),.doutb(w_in096_0[1]),.doutc(w_in096_0[2]),.din(in0[96]));
	jspl3 jspl3_w_in097_0(.douta(w_in097_0[0]),.doutb(w_in097_0[1]),.doutc(w_in097_0[2]),.din(in0[97]));
	jspl3 jspl3_w_in098_0(.douta(w_in098_0[0]),.doutb(w_in098_0[1]),.doutc(w_in098_0[2]),.din(in0[98]));
	jspl3 jspl3_w_in099_0(.douta(w_in099_0[0]),.doutb(w_in099_0[1]),.doutc(w_in099_0[2]),.din(in0[99]));
	jspl3 jspl3_w_in0100_0(.douta(w_in0100_0[0]),.doutb(w_in0100_0[1]),.doutc(w_in0100_0[2]),.din(in0[100]));
	jspl3 jspl3_w_in0101_0(.douta(w_in0101_0[0]),.doutb(w_in0101_0[1]),.doutc(w_in0101_0[2]),.din(in0[101]));
	jspl3 jspl3_w_in0102_0(.douta(w_in0102_0[0]),.doutb(w_in0102_0[1]),.doutc(w_in0102_0[2]),.din(in0[102]));
	jspl3 jspl3_w_in0103_0(.douta(w_in0103_0[0]),.doutb(w_in0103_0[1]),.doutc(w_in0103_0[2]),.din(in0[103]));
	jspl3 jspl3_w_in0104_0(.douta(w_in0104_0[0]),.doutb(w_in0104_0[1]),.doutc(w_in0104_0[2]),.din(in0[104]));
	jspl3 jspl3_w_in0105_0(.douta(w_in0105_0[0]),.doutb(w_in0105_0[1]),.doutc(w_in0105_0[2]),.din(in0[105]));
	jspl3 jspl3_w_in0106_0(.douta(w_in0106_0[0]),.doutb(w_in0106_0[1]),.doutc(w_in0106_0[2]),.din(in0[106]));
	jspl3 jspl3_w_in0107_0(.douta(w_in0107_0[0]),.doutb(w_in0107_0[1]),.doutc(w_in0107_0[2]),.din(in0[107]));
	jspl3 jspl3_w_in0108_0(.douta(w_in0108_0[0]),.doutb(w_in0108_0[1]),.doutc(w_in0108_0[2]),.din(in0[108]));
	jspl3 jspl3_w_in0109_0(.douta(w_in0109_0[0]),.doutb(w_in0109_0[1]),.doutc(w_in0109_0[2]),.din(in0[109]));
	jspl3 jspl3_w_in0110_0(.douta(w_in0110_0[0]),.doutb(w_in0110_0[1]),.doutc(w_in0110_0[2]),.din(in0[110]));
	jspl3 jspl3_w_in0111_0(.douta(w_in0111_0[0]),.doutb(w_in0111_0[1]),.doutc(w_in0111_0[2]),.din(in0[111]));
	jspl3 jspl3_w_in0112_0(.douta(w_in0112_0[0]),.doutb(w_in0112_0[1]),.doutc(w_in0112_0[2]),.din(in0[112]));
	jspl3 jspl3_w_in0113_0(.douta(w_in0113_0[0]),.doutb(w_in0113_0[1]),.doutc(w_in0113_0[2]),.din(in0[113]));
	jspl3 jspl3_w_in0114_0(.douta(w_in0114_0[0]),.doutb(w_in0114_0[1]),.doutc(w_in0114_0[2]),.din(in0[114]));
	jspl3 jspl3_w_in0115_0(.douta(w_in0115_0[0]),.doutb(w_in0115_0[1]),.doutc(w_in0115_0[2]),.din(in0[115]));
	jspl3 jspl3_w_in0116_0(.douta(w_in0116_0[0]),.doutb(w_in0116_0[1]),.doutc(w_in0116_0[2]),.din(in0[116]));
	jspl3 jspl3_w_in0117_0(.douta(w_in0117_0[0]),.doutb(w_in0117_0[1]),.doutc(w_in0117_0[2]),.din(in0[117]));
	jspl3 jspl3_w_in0118_0(.douta(w_in0118_0[0]),.doutb(w_in0118_0[1]),.doutc(w_in0118_0[2]),.din(in0[118]));
	jspl3 jspl3_w_in0119_0(.douta(w_in0119_0[0]),.doutb(w_in0119_0[1]),.doutc(w_in0119_0[2]),.din(in0[119]));
	jspl3 jspl3_w_in0120_0(.douta(w_in0120_0[0]),.doutb(w_in0120_0[1]),.doutc(w_in0120_0[2]),.din(in0[120]));
	jspl3 jspl3_w_in0121_0(.douta(w_in0121_0[0]),.doutb(w_in0121_0[1]),.doutc(w_in0121_0[2]),.din(in0[121]));
	jspl3 jspl3_w_in0122_0(.douta(w_in0122_0[0]),.doutb(w_in0122_0[1]),.doutc(w_in0122_0[2]),.din(in0[122]));
	jspl3 jspl3_w_in0123_0(.douta(w_in0123_0[0]),.doutb(w_in0123_0[1]),.doutc(w_in0123_0[2]),.din(in0[123]));
	jspl3 jspl3_w_in0124_0(.douta(w_in0124_0[0]),.doutb(w_in0124_0[1]),.doutc(w_in0124_0[2]),.din(in0[124]));
	jspl3 jspl3_w_in0125_0(.douta(w_in0125_0[0]),.doutb(w_in0125_0[1]),.doutc(w_in0125_0[2]),.din(in0[125]));
	jspl3 jspl3_w_in0126_0(.douta(w_in0126_0[0]),.doutb(w_in0126_0[1]),.doutc(w_in0126_0[2]),.din(in0[126]));
	jspl3 jspl3_w_in0127_0(.douta(w_in0127_0[0]),.doutb(w_in0127_0[1]),.doutc(w_in0127_0[2]),.din(in0[127]));
	jspl3 jspl3_w_in10_0(.douta(w_in10_0[0]),.doutb(w_in10_0[1]),.doutc(w_in10_0[2]),.din(in1[0]));
	jspl3 jspl3_w_in11_0(.douta(w_in11_0[0]),.doutb(w_in11_0[1]),.doutc(w_in11_0[2]),.din(in1[1]));
	jspl jspl_w_in11_1(.douta(w_in11_1[0]),.doutb(w_in11_1[1]),.din(w_in11_0[0]));
	jspl3 jspl3_w_in12_0(.douta(w_in12_0[0]),.doutb(w_in12_0[1]),.doutc(w_in12_0[2]),.din(in1[2]));
	jspl3 jspl3_w_in13_0(.douta(w_in13_0[0]),.doutb(w_in13_0[1]),.doutc(w_in13_0[2]),.din(in1[3]));
	jspl3 jspl3_w_in14_0(.douta(w_in14_0[0]),.doutb(w_in14_0[1]),.doutc(w_in14_0[2]),.din(in1[4]));
	jspl3 jspl3_w_in15_0(.douta(w_in15_0[0]),.doutb(w_in15_0[1]),.doutc(w_in15_0[2]),.din(in1[5]));
	jspl3 jspl3_w_in16_0(.douta(w_in16_0[0]),.doutb(w_in16_0[1]),.doutc(w_in16_0[2]),.din(in1[6]));
	jspl3 jspl3_w_in17_0(.douta(w_in17_0[0]),.doutb(w_in17_0[1]),.doutc(w_in17_0[2]),.din(in1[7]));
	jspl3 jspl3_w_in18_0(.douta(w_in18_0[0]),.doutb(w_in18_0[1]),.doutc(w_in18_0[2]),.din(in1[8]));
	jspl3 jspl3_w_in19_0(.douta(w_in19_0[0]),.doutb(w_in19_0[1]),.doutc(w_in19_0[2]),.din(in1[9]));
	jspl3 jspl3_w_in110_0(.douta(w_in110_0[0]),.doutb(w_in110_0[1]),.doutc(w_in110_0[2]),.din(in1[10]));
	jspl3 jspl3_w_in111_0(.douta(w_in111_0[0]),.doutb(w_in111_0[1]),.doutc(w_in111_0[2]),.din(in1[11]));
	jspl3 jspl3_w_in112_0(.douta(w_in112_0[0]),.doutb(w_in112_0[1]),.doutc(w_in112_0[2]),.din(in1[12]));
	jspl3 jspl3_w_in113_0(.douta(w_in113_0[0]),.doutb(w_in113_0[1]),.doutc(w_in113_0[2]),.din(in1[13]));
	jspl3 jspl3_w_in114_0(.douta(w_in114_0[0]),.doutb(w_in114_0[1]),.doutc(w_in114_0[2]),.din(in1[14]));
	jspl3 jspl3_w_in115_0(.douta(w_in115_0[0]),.doutb(w_in115_0[1]),.doutc(w_in115_0[2]),.din(in1[15]));
	jspl3 jspl3_w_in116_0(.douta(w_in116_0[0]),.doutb(w_in116_0[1]),.doutc(w_in116_0[2]),.din(in1[16]));
	jspl3 jspl3_w_in117_0(.douta(w_in117_0[0]),.doutb(w_in117_0[1]),.doutc(w_in117_0[2]),.din(in1[17]));
	jspl3 jspl3_w_in118_0(.douta(w_in118_0[0]),.doutb(w_in118_0[1]),.doutc(w_in118_0[2]),.din(in1[18]));
	jspl3 jspl3_w_in119_0(.douta(w_in119_0[0]),.doutb(w_in119_0[1]),.doutc(w_in119_0[2]),.din(in1[19]));
	jspl3 jspl3_w_in120_0(.douta(w_in120_0[0]),.doutb(w_in120_0[1]),.doutc(w_in120_0[2]),.din(in1[20]));
	jspl3 jspl3_w_in121_0(.douta(w_in121_0[0]),.doutb(w_in121_0[1]),.doutc(w_in121_0[2]),.din(in1[21]));
	jspl3 jspl3_w_in122_0(.douta(w_in122_0[0]),.doutb(w_in122_0[1]),.doutc(w_in122_0[2]),.din(in1[22]));
	jspl3 jspl3_w_in123_0(.douta(w_in123_0[0]),.doutb(w_in123_0[1]),.doutc(w_in123_0[2]),.din(in1[23]));
	jspl3 jspl3_w_in124_0(.douta(w_in124_0[0]),.doutb(w_in124_0[1]),.doutc(w_in124_0[2]),.din(in1[24]));
	jspl3 jspl3_w_in125_0(.douta(w_in125_0[0]),.doutb(w_in125_0[1]),.doutc(w_in125_0[2]),.din(in1[25]));
	jspl3 jspl3_w_in126_0(.douta(w_in126_0[0]),.doutb(w_in126_0[1]),.doutc(w_in126_0[2]),.din(in1[26]));
	jspl3 jspl3_w_in127_0(.douta(w_in127_0[0]),.doutb(w_in127_0[1]),.doutc(w_in127_0[2]),.din(in1[27]));
	jspl3 jspl3_w_in128_0(.douta(w_in128_0[0]),.doutb(w_in128_0[1]),.doutc(w_in128_0[2]),.din(in1[28]));
	jspl3 jspl3_w_in129_0(.douta(w_in129_0[0]),.doutb(w_in129_0[1]),.doutc(w_in129_0[2]),.din(in1[29]));
	jspl3 jspl3_w_in130_0(.douta(w_in130_0[0]),.doutb(w_in130_0[1]),.doutc(w_in130_0[2]),.din(in1[30]));
	jspl3 jspl3_w_in131_0(.douta(w_in131_0[0]),.doutb(w_in131_0[1]),.doutc(w_in131_0[2]),.din(in1[31]));
	jspl3 jspl3_w_in132_0(.douta(w_in132_0[0]),.doutb(w_in132_0[1]),.doutc(w_in132_0[2]),.din(in1[32]));
	jspl3 jspl3_w_in133_0(.douta(w_in133_0[0]),.doutb(w_in133_0[1]),.doutc(w_in133_0[2]),.din(in1[33]));
	jspl3 jspl3_w_in134_0(.douta(w_in134_0[0]),.doutb(w_in134_0[1]),.doutc(w_in134_0[2]),.din(in1[34]));
	jspl3 jspl3_w_in135_0(.douta(w_in135_0[0]),.doutb(w_in135_0[1]),.doutc(w_in135_0[2]),.din(in1[35]));
	jspl3 jspl3_w_in136_0(.douta(w_in136_0[0]),.doutb(w_in136_0[1]),.doutc(w_in136_0[2]),.din(in1[36]));
	jspl3 jspl3_w_in137_0(.douta(w_in137_0[0]),.doutb(w_in137_0[1]),.doutc(w_in137_0[2]),.din(in1[37]));
	jspl3 jspl3_w_in138_0(.douta(w_in138_0[0]),.doutb(w_in138_0[1]),.doutc(w_in138_0[2]),.din(in1[38]));
	jspl3 jspl3_w_in139_0(.douta(w_in139_0[0]),.doutb(w_in139_0[1]),.doutc(w_in139_0[2]),.din(in1[39]));
	jspl3 jspl3_w_in140_0(.douta(w_in140_0[0]),.doutb(w_in140_0[1]),.doutc(w_in140_0[2]),.din(in1[40]));
	jspl3 jspl3_w_in141_0(.douta(w_in141_0[0]),.doutb(w_in141_0[1]),.doutc(w_in141_0[2]),.din(in1[41]));
	jspl3 jspl3_w_in142_0(.douta(w_in142_0[0]),.doutb(w_in142_0[1]),.doutc(w_in142_0[2]),.din(in1[42]));
	jspl3 jspl3_w_in143_0(.douta(w_in143_0[0]),.doutb(w_in143_0[1]),.doutc(w_in143_0[2]),.din(in1[43]));
	jspl3 jspl3_w_in144_0(.douta(w_in144_0[0]),.doutb(w_in144_0[1]),.doutc(w_in144_0[2]),.din(in1[44]));
	jspl3 jspl3_w_in145_0(.douta(w_in145_0[0]),.doutb(w_in145_0[1]),.doutc(w_in145_0[2]),.din(in1[45]));
	jspl3 jspl3_w_in146_0(.douta(w_in146_0[0]),.doutb(w_in146_0[1]),.doutc(w_in146_0[2]),.din(in1[46]));
	jspl3 jspl3_w_in147_0(.douta(w_in147_0[0]),.doutb(w_in147_0[1]),.doutc(w_in147_0[2]),.din(in1[47]));
	jspl3 jspl3_w_in148_0(.douta(w_in148_0[0]),.doutb(w_in148_0[1]),.doutc(w_in148_0[2]),.din(in1[48]));
	jspl3 jspl3_w_in149_0(.douta(w_in149_0[0]),.doutb(w_in149_0[1]),.doutc(w_in149_0[2]),.din(in1[49]));
	jspl3 jspl3_w_in150_0(.douta(w_in150_0[0]),.doutb(w_in150_0[1]),.doutc(w_in150_0[2]),.din(in1[50]));
	jspl3 jspl3_w_in151_0(.douta(w_in151_0[0]),.doutb(w_in151_0[1]),.doutc(w_in151_0[2]),.din(in1[51]));
	jspl jspl_w_in152_0(.douta(w_in152_0[0]),.doutb(w_in152_0[1]),.din(in1[52]));
	jspl3 jspl3_w_in153_0(.douta(w_in153_0[0]),.doutb(w_in153_0[1]),.doutc(w_in153_0[2]),.din(in1[53]));
	jspl3 jspl3_w_in154_0(.douta(w_in154_0[0]),.doutb(w_in154_0[1]),.doutc(w_in154_0[2]),.din(in1[54]));
	jspl3 jspl3_w_in155_0(.douta(w_in155_0[0]),.doutb(w_in155_0[1]),.doutc(w_in155_0[2]),.din(in1[55]));
	jspl3 jspl3_w_in156_0(.douta(w_in156_0[0]),.doutb(w_in156_0[1]),.doutc(w_in156_0[2]),.din(in1[56]));
	jspl3 jspl3_w_in157_0(.douta(w_in157_0[0]),.doutb(w_in157_0[1]),.doutc(w_in157_0[2]),.din(in1[57]));
	jspl3 jspl3_w_in158_0(.douta(w_in158_0[0]),.doutb(w_in158_0[1]),.doutc(w_in158_0[2]),.din(in1[58]));
	jspl3 jspl3_w_in159_0(.douta(w_in159_0[0]),.doutb(w_in159_0[1]),.doutc(w_in159_0[2]),.din(in1[59]));
	jspl3 jspl3_w_in160_0(.douta(w_in160_0[0]),.doutb(w_in160_0[1]),.doutc(w_in160_0[2]),.din(in1[60]));
	jspl3 jspl3_w_in161_0(.douta(w_in161_0[0]),.doutb(w_in161_0[1]),.doutc(w_in161_0[2]),.din(in1[61]));
	jspl3 jspl3_w_in162_0(.douta(w_in162_0[0]),.doutb(w_in162_0[1]),.doutc(w_in162_0[2]),.din(in1[62]));
	jspl3 jspl3_w_in163_0(.douta(w_in163_0[0]),.doutb(w_in163_0[1]),.doutc(w_in163_0[2]),.din(in1[63]));
	jspl3 jspl3_w_in164_0(.douta(w_in164_0[0]),.doutb(w_in164_0[1]),.doutc(w_in164_0[2]),.din(in1[64]));
	jspl3 jspl3_w_in165_0(.douta(w_in165_0[0]),.doutb(w_in165_0[1]),.doutc(w_in165_0[2]),.din(in1[65]));
	jspl3 jspl3_w_in166_0(.douta(w_in166_0[0]),.doutb(w_in166_0[1]),.doutc(w_in166_0[2]),.din(in1[66]));
	jspl3 jspl3_w_in167_0(.douta(w_in167_0[0]),.doutb(w_in167_0[1]),.doutc(w_in167_0[2]),.din(in1[67]));
	jspl3 jspl3_w_in168_0(.douta(w_in168_0[0]),.doutb(w_in168_0[1]),.doutc(w_in168_0[2]),.din(in1[68]));
	jspl3 jspl3_w_in169_0(.douta(w_in169_0[0]),.doutb(w_in169_0[1]),.doutc(w_in169_0[2]),.din(in1[69]));
	jspl3 jspl3_w_in170_0(.douta(w_in170_0[0]),.doutb(w_in170_0[1]),.doutc(w_in170_0[2]),.din(in1[70]));
	jspl3 jspl3_w_in171_0(.douta(w_in171_0[0]),.doutb(w_in171_0[1]),.doutc(w_in171_0[2]),.din(in1[71]));
	jspl3 jspl3_w_in172_0(.douta(w_in172_0[0]),.doutb(w_in172_0[1]),.doutc(w_in172_0[2]),.din(in1[72]));
	jspl3 jspl3_w_in173_0(.douta(w_in173_0[0]),.doutb(w_in173_0[1]),.doutc(w_in173_0[2]),.din(in1[73]));
	jspl3 jspl3_w_in174_0(.douta(w_in174_0[0]),.doutb(w_in174_0[1]),.doutc(w_in174_0[2]),.din(in1[74]));
	jspl3 jspl3_w_in175_0(.douta(w_in175_0[0]),.doutb(w_in175_0[1]),.doutc(w_in175_0[2]),.din(in1[75]));
	jspl3 jspl3_w_in176_0(.douta(w_in176_0[0]),.doutb(w_in176_0[1]),.doutc(w_in176_0[2]),.din(in1[76]));
	jspl3 jspl3_w_in177_0(.douta(w_in177_0[0]),.doutb(w_in177_0[1]),.doutc(w_in177_0[2]),.din(in1[77]));
	jspl3 jspl3_w_in178_0(.douta(w_in178_0[0]),.doutb(w_in178_0[1]),.doutc(w_in178_0[2]),.din(in1[78]));
	jspl3 jspl3_w_in179_0(.douta(w_in179_0[0]),.doutb(w_in179_0[1]),.doutc(w_in179_0[2]),.din(in1[79]));
	jspl3 jspl3_w_in180_0(.douta(w_in180_0[0]),.doutb(w_in180_0[1]),.doutc(w_in180_0[2]),.din(in1[80]));
	jspl3 jspl3_w_in181_0(.douta(w_in181_0[0]),.doutb(w_in181_0[1]),.doutc(w_in181_0[2]),.din(in1[81]));
	jspl3 jspl3_w_in182_0(.douta(w_in182_0[0]),.doutb(w_in182_0[1]),.doutc(w_in182_0[2]),.din(in1[82]));
	jspl3 jspl3_w_in183_0(.douta(w_in183_0[0]),.doutb(w_in183_0[1]),.doutc(w_in183_0[2]),.din(in1[83]));
	jspl3 jspl3_w_in184_0(.douta(w_in184_0[0]),.doutb(w_in184_0[1]),.doutc(w_in184_0[2]),.din(in1[84]));
	jspl3 jspl3_w_in185_0(.douta(w_in185_0[0]),.doutb(w_in185_0[1]),.doutc(w_in185_0[2]),.din(in1[85]));
	jspl3 jspl3_w_in186_0(.douta(w_in186_0[0]),.doutb(w_in186_0[1]),.doutc(w_in186_0[2]),.din(in1[86]));
	jspl3 jspl3_w_in187_0(.douta(w_in187_0[0]),.doutb(w_in187_0[1]),.doutc(w_in187_0[2]),.din(in1[87]));
	jspl3 jspl3_w_in188_0(.douta(w_in188_0[0]),.doutb(w_in188_0[1]),.doutc(w_in188_0[2]),.din(in1[88]));
	jspl3 jspl3_w_in189_0(.douta(w_in189_0[0]),.doutb(w_in189_0[1]),.doutc(w_in189_0[2]),.din(in1[89]));
	jspl3 jspl3_w_in190_0(.douta(w_in190_0[0]),.doutb(w_in190_0[1]),.doutc(w_in190_0[2]),.din(in1[90]));
	jspl3 jspl3_w_in191_0(.douta(w_in191_0[0]),.doutb(w_in191_0[1]),.doutc(w_in191_0[2]),.din(in1[91]));
	jspl3 jspl3_w_in192_0(.douta(w_in192_0[0]),.doutb(w_in192_0[1]),.doutc(w_in192_0[2]),.din(in1[92]));
	jspl3 jspl3_w_in193_0(.douta(w_in193_0[0]),.doutb(w_in193_0[1]),.doutc(w_in193_0[2]),.din(in1[93]));
	jspl3 jspl3_w_in194_0(.douta(w_in194_0[0]),.doutb(w_in194_0[1]),.doutc(w_in194_0[2]),.din(in1[94]));
	jspl3 jspl3_w_in195_0(.douta(w_in195_0[0]),.doutb(w_in195_0[1]),.doutc(w_in195_0[2]),.din(in1[95]));
	jspl3 jspl3_w_in196_0(.douta(w_in196_0[0]),.doutb(w_in196_0[1]),.doutc(w_in196_0[2]),.din(in1[96]));
	jspl3 jspl3_w_in197_0(.douta(w_in197_0[0]),.doutb(w_in197_0[1]),.doutc(w_in197_0[2]),.din(in1[97]));
	jspl3 jspl3_w_in198_0(.douta(w_in198_0[0]),.doutb(w_in198_0[1]),.doutc(w_in198_0[2]),.din(in1[98]));
	jspl3 jspl3_w_in199_0(.douta(w_in199_0[0]),.doutb(w_in199_0[1]),.doutc(w_in199_0[2]),.din(in1[99]));
	jspl3 jspl3_w_in1100_0(.douta(w_in1100_0[0]),.doutb(w_in1100_0[1]),.doutc(w_in1100_0[2]),.din(in1[100]));
	jspl3 jspl3_w_in1101_0(.douta(w_in1101_0[0]),.doutb(w_in1101_0[1]),.doutc(w_in1101_0[2]),.din(in1[101]));
	jspl3 jspl3_w_in1102_0(.douta(w_in1102_0[0]),.doutb(w_in1102_0[1]),.doutc(w_in1102_0[2]),.din(in1[102]));
	jspl3 jspl3_w_in1103_0(.douta(w_in1103_0[0]),.doutb(w_in1103_0[1]),.doutc(w_in1103_0[2]),.din(in1[103]));
	jspl3 jspl3_w_in1104_0(.douta(w_in1104_0[0]),.doutb(w_in1104_0[1]),.doutc(w_in1104_0[2]),.din(in1[104]));
	jspl3 jspl3_w_in1105_0(.douta(w_in1105_0[0]),.doutb(w_in1105_0[1]),.doutc(w_in1105_0[2]),.din(in1[105]));
	jspl3 jspl3_w_in1106_0(.douta(w_in1106_0[0]),.doutb(w_in1106_0[1]),.doutc(w_in1106_0[2]),.din(in1[106]));
	jspl3 jspl3_w_in1107_0(.douta(w_in1107_0[0]),.doutb(w_in1107_0[1]),.doutc(w_in1107_0[2]),.din(in1[107]));
	jspl3 jspl3_w_in1108_0(.douta(w_in1108_0[0]),.doutb(w_in1108_0[1]),.doutc(w_in1108_0[2]),.din(in1[108]));
	jspl3 jspl3_w_in1109_0(.douta(w_in1109_0[0]),.doutb(w_in1109_0[1]),.doutc(w_in1109_0[2]),.din(in1[109]));
	jspl3 jspl3_w_in1110_0(.douta(w_in1110_0[0]),.doutb(w_in1110_0[1]),.doutc(w_in1110_0[2]),.din(in1[110]));
	jspl3 jspl3_w_in1111_0(.douta(w_in1111_0[0]),.doutb(w_in1111_0[1]),.doutc(w_in1111_0[2]),.din(in1[111]));
	jspl3 jspl3_w_in1112_0(.douta(w_in1112_0[0]),.doutb(w_in1112_0[1]),.doutc(w_in1112_0[2]),.din(in1[112]));
	jspl3 jspl3_w_in1113_0(.douta(w_in1113_0[0]),.doutb(w_in1113_0[1]),.doutc(w_in1113_0[2]),.din(in1[113]));
	jspl3 jspl3_w_in1114_0(.douta(w_in1114_0[0]),.doutb(w_in1114_0[1]),.doutc(w_in1114_0[2]),.din(in1[114]));
	jspl3 jspl3_w_in1115_0(.douta(w_in1115_0[0]),.doutb(w_in1115_0[1]),.doutc(w_in1115_0[2]),.din(in1[115]));
	jspl3 jspl3_w_in1116_0(.douta(w_in1116_0[0]),.doutb(w_in1116_0[1]),.doutc(w_in1116_0[2]),.din(in1[116]));
	jspl3 jspl3_w_in1117_0(.douta(w_in1117_0[0]),.doutb(w_in1117_0[1]),.doutc(w_in1117_0[2]),.din(in1[117]));
	jspl3 jspl3_w_in1118_0(.douta(w_in1118_0[0]),.doutb(w_in1118_0[1]),.doutc(w_in1118_0[2]),.din(in1[118]));
	jspl3 jspl3_w_in1119_0(.douta(w_in1119_0[0]),.doutb(w_in1119_0[1]),.doutc(w_in1119_0[2]),.din(in1[119]));
	jspl3 jspl3_w_in1120_0(.douta(w_in1120_0[0]),.doutb(w_in1120_0[1]),.doutc(w_in1120_0[2]),.din(in1[120]));
	jspl3 jspl3_w_in1121_0(.douta(w_in1121_0[0]),.doutb(w_in1121_0[1]),.doutc(w_in1121_0[2]),.din(in1[121]));
	jspl3 jspl3_w_in1122_0(.douta(w_in1122_0[0]),.doutb(w_in1122_0[1]),.doutc(w_in1122_0[2]),.din(in1[122]));
	jspl3 jspl3_w_in1123_0(.douta(w_in1123_0[0]),.doutb(w_in1123_0[1]),.doutc(w_in1123_0[2]),.din(in1[123]));
	jspl3 jspl3_w_in1124_0(.douta(w_in1124_0[0]),.doutb(w_in1124_0[1]),.doutc(w_in1124_0[2]),.din(in1[124]));
	jspl3 jspl3_w_in1125_0(.douta(w_in1125_0[0]),.doutb(w_in1125_0[1]),.doutc(w_in1125_0[2]),.din(in1[125]));
	jspl3 jspl3_w_in1126_0(.douta(w_in1126_0[0]),.doutb(w_in1126_0[1]),.doutc(w_in1126_0[2]),.din(in1[126]));
	jspl3 jspl3_w_in1127_0(.douta(w_in1127_0[0]),.doutb(w_in1127_0[1]),.doutc(w_in1127_0[2]),.din(in1[127]));
	jspl3 jspl3_w_in20_0(.douta(w_in20_0[0]),.doutb(w_in20_0[1]),.doutc(w_in20_0[2]),.din(in2[0]));
	jspl3 jspl3_w_in21_0(.douta(w_in21_0[0]),.doutb(w_in21_0[1]),.doutc(w_in21_0[2]),.din(in2[1]));
	jspl jspl_w_in21_1(.douta(w_in21_1[0]),.doutb(w_in21_1[1]),.din(w_in21_0[0]));
	jspl3 jspl3_w_in22_0(.douta(w_in22_0[0]),.doutb(w_in22_0[1]),.doutc(w_in22_0[2]),.din(in2[2]));
	jspl3 jspl3_w_in23_0(.douta(w_in23_0[0]),.doutb(w_in23_0[1]),.doutc(w_in23_0[2]),.din(in2[3]));
	jspl3 jspl3_w_in24_0(.douta(w_in24_0[0]),.doutb(w_in24_0[1]),.doutc(w_in24_0[2]),.din(in2[4]));
	jspl3 jspl3_w_in25_0(.douta(w_in25_0[0]),.doutb(w_in25_0[1]),.doutc(w_in25_0[2]),.din(in2[5]));
	jspl3 jspl3_w_in26_0(.douta(w_in26_0[0]),.doutb(w_in26_0[1]),.doutc(w_in26_0[2]),.din(in2[6]));
	jspl3 jspl3_w_in27_0(.douta(w_in27_0[0]),.doutb(w_in27_0[1]),.doutc(w_in27_0[2]),.din(in2[7]));
	jspl3 jspl3_w_in28_0(.douta(w_in28_0[0]),.doutb(w_in28_0[1]),.doutc(w_in28_0[2]),.din(in2[8]));
	jspl3 jspl3_w_in29_0(.douta(w_in29_0[0]),.doutb(w_in29_0[1]),.doutc(w_in29_0[2]),.din(in2[9]));
	jspl3 jspl3_w_in210_0(.douta(w_in210_0[0]),.doutb(w_in210_0[1]),.doutc(w_in210_0[2]),.din(in2[10]));
	jspl3 jspl3_w_in211_0(.douta(w_in211_0[0]),.doutb(w_in211_0[1]),.doutc(w_in211_0[2]),.din(in2[11]));
	jspl3 jspl3_w_in212_0(.douta(w_in212_0[0]),.doutb(w_in212_0[1]),.doutc(w_in212_0[2]),.din(in2[12]));
	jspl3 jspl3_w_in213_0(.douta(w_in213_0[0]),.doutb(w_in213_0[1]),.doutc(w_in213_0[2]),.din(in2[13]));
	jspl3 jspl3_w_in214_0(.douta(w_in214_0[0]),.doutb(w_in214_0[1]),.doutc(w_in214_0[2]),.din(in2[14]));
	jspl3 jspl3_w_in215_0(.douta(w_in215_0[0]),.doutb(w_in215_0[1]),.doutc(w_in215_0[2]),.din(in2[15]));
	jspl3 jspl3_w_in216_0(.douta(w_in216_0[0]),.doutb(w_in216_0[1]),.doutc(w_in216_0[2]),.din(in2[16]));
	jspl3 jspl3_w_in217_0(.douta(w_in217_0[0]),.doutb(w_in217_0[1]),.doutc(w_in217_0[2]),.din(in2[17]));
	jspl3 jspl3_w_in218_0(.douta(w_in218_0[0]),.doutb(w_in218_0[1]),.doutc(w_in218_0[2]),.din(in2[18]));
	jspl3 jspl3_w_in219_0(.douta(w_in219_0[0]),.doutb(w_in219_0[1]),.doutc(w_in219_0[2]),.din(in2[19]));
	jspl3 jspl3_w_in220_0(.douta(w_in220_0[0]),.doutb(w_in220_0[1]),.doutc(w_in220_0[2]),.din(in2[20]));
	jspl3 jspl3_w_in221_0(.douta(w_in221_0[0]),.doutb(w_in221_0[1]),.doutc(w_in221_0[2]),.din(in2[21]));
	jspl3 jspl3_w_in222_0(.douta(w_in222_0[0]),.doutb(w_in222_0[1]),.doutc(w_in222_0[2]),.din(in2[22]));
	jspl3 jspl3_w_in223_0(.douta(w_in223_0[0]),.doutb(w_in223_0[1]),.doutc(w_in223_0[2]),.din(in2[23]));
	jspl3 jspl3_w_in224_0(.douta(w_in224_0[0]),.doutb(w_in224_0[1]),.doutc(w_in224_0[2]),.din(in2[24]));
	jspl3 jspl3_w_in225_0(.douta(w_in225_0[0]),.doutb(w_in225_0[1]),.doutc(w_in225_0[2]),.din(in2[25]));
	jspl3 jspl3_w_in226_0(.douta(w_in226_0[0]),.doutb(w_in226_0[1]),.doutc(w_in226_0[2]),.din(in2[26]));
	jspl3 jspl3_w_in227_0(.douta(w_in227_0[0]),.doutb(w_in227_0[1]),.doutc(w_in227_0[2]),.din(in2[27]));
	jspl3 jspl3_w_in228_0(.douta(w_in228_0[0]),.doutb(w_in228_0[1]),.doutc(w_in228_0[2]),.din(in2[28]));
	jspl3 jspl3_w_in229_0(.douta(w_in229_0[0]),.doutb(w_in229_0[1]),.doutc(w_in229_0[2]),.din(in2[29]));
	jspl3 jspl3_w_in230_0(.douta(w_in230_0[0]),.doutb(w_in230_0[1]),.doutc(w_in230_0[2]),.din(in2[30]));
	jspl3 jspl3_w_in231_0(.douta(w_in231_0[0]),.doutb(w_in231_0[1]),.doutc(w_in231_0[2]),.din(in2[31]));
	jspl3 jspl3_w_in232_0(.douta(w_in232_0[0]),.doutb(w_in232_0[1]),.doutc(w_in232_0[2]),.din(in2[32]));
	jspl3 jspl3_w_in233_0(.douta(w_in233_0[0]),.doutb(w_in233_0[1]),.doutc(w_in233_0[2]),.din(in2[33]));
	jspl3 jspl3_w_in234_0(.douta(w_in234_0[0]),.doutb(w_in234_0[1]),.doutc(w_in234_0[2]),.din(in2[34]));
	jspl3 jspl3_w_in235_0(.douta(w_in235_0[0]),.doutb(w_in235_0[1]),.doutc(w_in235_0[2]),.din(in2[35]));
	jspl3 jspl3_w_in236_0(.douta(w_in236_0[0]),.doutb(w_in236_0[1]),.doutc(w_in236_0[2]),.din(in2[36]));
	jspl3 jspl3_w_in237_0(.douta(w_in237_0[0]),.doutb(w_in237_0[1]),.doutc(w_in237_0[2]),.din(in2[37]));
	jspl3 jspl3_w_in238_0(.douta(w_in238_0[0]),.doutb(w_in238_0[1]),.doutc(w_in238_0[2]),.din(in2[38]));
	jspl3 jspl3_w_in239_0(.douta(w_in239_0[0]),.doutb(w_in239_0[1]),.doutc(w_in239_0[2]),.din(in2[39]));
	jspl3 jspl3_w_in240_0(.douta(w_in240_0[0]),.doutb(w_in240_0[1]),.doutc(w_in240_0[2]),.din(in2[40]));
	jspl3 jspl3_w_in241_0(.douta(w_in241_0[0]),.doutb(w_in241_0[1]),.doutc(w_in241_0[2]),.din(in2[41]));
	jspl3 jspl3_w_in242_0(.douta(w_in242_0[0]),.doutb(w_in242_0[1]),.doutc(w_in242_0[2]),.din(in2[42]));
	jspl3 jspl3_w_in243_0(.douta(w_in243_0[0]),.doutb(w_in243_0[1]),.doutc(w_in243_0[2]),.din(in2[43]));
	jspl3 jspl3_w_in244_0(.douta(w_in244_0[0]),.doutb(w_in244_0[1]),.doutc(w_in244_0[2]),.din(in2[44]));
	jspl3 jspl3_w_in245_0(.douta(w_in245_0[0]),.doutb(w_in245_0[1]),.doutc(w_in245_0[2]),.din(in2[45]));
	jspl3 jspl3_w_in246_0(.douta(w_in246_0[0]),.doutb(w_in246_0[1]),.doutc(w_in246_0[2]),.din(in2[46]));
	jspl3 jspl3_w_in247_0(.douta(w_in247_0[0]),.doutb(w_in247_0[1]),.doutc(w_in247_0[2]),.din(in2[47]));
	jspl3 jspl3_w_in248_0(.douta(w_in248_0[0]),.doutb(w_in248_0[1]),.doutc(w_in248_0[2]),.din(in2[48]));
	jspl3 jspl3_w_in249_0(.douta(w_in249_0[0]),.doutb(w_in249_0[1]),.doutc(w_in249_0[2]),.din(in2[49]));
	jspl3 jspl3_w_in250_0(.douta(w_in250_0[0]),.doutb(w_in250_0[1]),.doutc(w_in250_0[2]),.din(in2[50]));
	jspl3 jspl3_w_in251_0(.douta(w_in251_0[0]),.doutb(w_in251_0[1]),.doutc(w_in251_0[2]),.din(in2[51]));
	jspl3 jspl3_w_in252_0(.douta(w_in252_0[0]),.doutb(w_in252_0[1]),.doutc(w_in252_0[2]),.din(in2[52]));
	jspl3 jspl3_w_in253_0(.douta(w_in253_0[0]),.doutb(w_in253_0[1]),.doutc(w_in253_0[2]),.din(in2[53]));
	jspl3 jspl3_w_in254_0(.douta(w_in254_0[0]),.doutb(w_in254_0[1]),.doutc(w_in254_0[2]),.din(in2[54]));
	jspl3 jspl3_w_in255_0(.douta(w_in255_0[0]),.doutb(w_in255_0[1]),.doutc(w_in255_0[2]),.din(in2[55]));
	jspl3 jspl3_w_in256_0(.douta(w_in256_0[0]),.doutb(w_in256_0[1]),.doutc(w_in256_0[2]),.din(in2[56]));
	jspl3 jspl3_w_in257_0(.douta(w_in257_0[0]),.doutb(w_in257_0[1]),.doutc(w_in257_0[2]),.din(in2[57]));
	jspl3 jspl3_w_in258_0(.douta(w_in258_0[0]),.doutb(w_in258_0[1]),.doutc(w_in258_0[2]),.din(in2[58]));
	jspl3 jspl3_w_in259_0(.douta(w_in259_0[0]),.doutb(w_in259_0[1]),.doutc(w_in259_0[2]),.din(in2[59]));
	jspl3 jspl3_w_in260_0(.douta(w_in260_0[0]),.doutb(w_in260_0[1]),.doutc(w_in260_0[2]),.din(in2[60]));
	jspl3 jspl3_w_in261_0(.douta(w_in261_0[0]),.doutb(w_in261_0[1]),.doutc(w_in261_0[2]),.din(in2[61]));
	jspl3 jspl3_w_in262_0(.douta(w_in262_0[0]),.doutb(w_in262_0[1]),.doutc(w_in262_0[2]),.din(in2[62]));
	jspl3 jspl3_w_in263_0(.douta(w_in263_0[0]),.doutb(w_in263_0[1]),.doutc(w_in263_0[2]),.din(in2[63]));
	jspl3 jspl3_w_in264_0(.douta(w_in264_0[0]),.doutb(w_in264_0[1]),.doutc(w_in264_0[2]),.din(in2[64]));
	jspl3 jspl3_w_in265_0(.douta(w_in265_0[0]),.doutb(w_in265_0[1]),.doutc(w_in265_0[2]),.din(in2[65]));
	jspl3 jspl3_w_in266_0(.douta(w_in266_0[0]),.doutb(w_in266_0[1]),.doutc(w_in266_0[2]),.din(in2[66]));
	jspl3 jspl3_w_in267_0(.douta(w_in267_0[0]),.doutb(w_in267_0[1]),.doutc(w_in267_0[2]),.din(in2[67]));
	jspl3 jspl3_w_in268_0(.douta(w_in268_0[0]),.doutb(w_in268_0[1]),.doutc(w_in268_0[2]),.din(in2[68]));
	jspl3 jspl3_w_in269_0(.douta(w_in269_0[0]),.doutb(w_in269_0[1]),.doutc(w_in269_0[2]),.din(in2[69]));
	jspl3 jspl3_w_in270_0(.douta(w_in270_0[0]),.doutb(w_in270_0[1]),.doutc(w_in270_0[2]),.din(in2[70]));
	jspl3 jspl3_w_in271_0(.douta(w_in271_0[0]),.doutb(w_in271_0[1]),.doutc(w_in271_0[2]),.din(in2[71]));
	jspl3 jspl3_w_in272_0(.douta(w_in272_0[0]),.doutb(w_in272_0[1]),.doutc(w_in272_0[2]),.din(in2[72]));
	jspl3 jspl3_w_in273_0(.douta(w_in273_0[0]),.doutb(w_in273_0[1]),.doutc(w_in273_0[2]),.din(in2[73]));
	jspl3 jspl3_w_in274_0(.douta(w_in274_0[0]),.doutb(w_in274_0[1]),.doutc(w_in274_0[2]),.din(in2[74]));
	jspl3 jspl3_w_in275_0(.douta(w_in275_0[0]),.doutb(w_in275_0[1]),.doutc(w_in275_0[2]),.din(in2[75]));
	jspl3 jspl3_w_in276_0(.douta(w_in276_0[0]),.doutb(w_in276_0[1]),.doutc(w_in276_0[2]),.din(in2[76]));
	jspl3 jspl3_w_in277_0(.douta(w_in277_0[0]),.doutb(w_in277_0[1]),.doutc(w_in277_0[2]),.din(in2[77]));
	jspl3 jspl3_w_in278_0(.douta(w_in278_0[0]),.doutb(w_in278_0[1]),.doutc(w_in278_0[2]),.din(in2[78]));
	jspl3 jspl3_w_in279_0(.douta(w_in279_0[0]),.doutb(w_in279_0[1]),.doutc(w_in279_0[2]),.din(in2[79]));
	jspl3 jspl3_w_in280_0(.douta(w_in280_0[0]),.doutb(w_in280_0[1]),.doutc(w_in280_0[2]),.din(in2[80]));
	jspl3 jspl3_w_in281_0(.douta(w_in281_0[0]),.doutb(w_in281_0[1]),.doutc(w_in281_0[2]),.din(in2[81]));
	jspl3 jspl3_w_in282_0(.douta(w_in282_0[0]),.doutb(w_in282_0[1]),.doutc(w_in282_0[2]),.din(in2[82]));
	jspl3 jspl3_w_in283_0(.douta(w_in283_0[0]),.doutb(w_in283_0[1]),.doutc(w_in283_0[2]),.din(in2[83]));
	jspl3 jspl3_w_in284_0(.douta(w_in284_0[0]),.doutb(w_in284_0[1]),.doutc(w_in284_0[2]),.din(in2[84]));
	jspl3 jspl3_w_in285_0(.douta(w_in285_0[0]),.doutb(w_in285_0[1]),.doutc(w_in285_0[2]),.din(in2[85]));
	jspl3 jspl3_w_in286_0(.douta(w_in286_0[0]),.doutb(w_in286_0[1]),.doutc(w_in286_0[2]),.din(in2[86]));
	jspl3 jspl3_w_in287_0(.douta(w_in287_0[0]),.doutb(w_in287_0[1]),.doutc(w_in287_0[2]),.din(in2[87]));
	jspl3 jspl3_w_in288_0(.douta(w_in288_0[0]),.doutb(w_in288_0[1]),.doutc(w_in288_0[2]),.din(in2[88]));
	jspl3 jspl3_w_in289_0(.douta(w_in289_0[0]),.doutb(w_in289_0[1]),.doutc(w_in289_0[2]),.din(in2[89]));
	jspl3 jspl3_w_in290_0(.douta(w_in290_0[0]),.doutb(w_in290_0[1]),.doutc(w_in290_0[2]),.din(in2[90]));
	jspl3 jspl3_w_in291_0(.douta(w_in291_0[0]),.doutb(w_in291_0[1]),.doutc(w_in291_0[2]),.din(in2[91]));
	jspl3 jspl3_w_in292_0(.douta(w_in292_0[0]),.doutb(w_in292_0[1]),.doutc(w_in292_0[2]),.din(in2[92]));
	jspl3 jspl3_w_in293_0(.douta(w_in293_0[0]),.doutb(w_in293_0[1]),.doutc(w_in293_0[2]),.din(in2[93]));
	jspl3 jspl3_w_in294_0(.douta(w_in294_0[0]),.doutb(w_in294_0[1]),.doutc(w_in294_0[2]),.din(in2[94]));
	jspl3 jspl3_w_in295_0(.douta(w_in295_0[0]),.doutb(w_in295_0[1]),.doutc(w_in295_0[2]),.din(in2[95]));
	jspl3 jspl3_w_in296_0(.douta(w_in296_0[0]),.doutb(w_in296_0[1]),.doutc(w_in296_0[2]),.din(in2[96]));
	jspl3 jspl3_w_in297_0(.douta(w_in297_0[0]),.doutb(w_in297_0[1]),.doutc(w_in297_0[2]),.din(in2[97]));
	jspl3 jspl3_w_in298_0(.douta(w_in298_0[0]),.doutb(w_in298_0[1]),.doutc(w_in298_0[2]),.din(in2[98]));
	jspl3 jspl3_w_in299_0(.douta(w_in299_0[0]),.doutb(w_in299_0[1]),.doutc(w_in299_0[2]),.din(in2[99]));
	jspl3 jspl3_w_in2100_0(.douta(w_in2100_0[0]),.doutb(w_in2100_0[1]),.doutc(w_in2100_0[2]),.din(in2[100]));
	jspl3 jspl3_w_in2101_0(.douta(w_in2101_0[0]),.doutb(w_in2101_0[1]),.doutc(w_in2101_0[2]),.din(in2[101]));
	jspl3 jspl3_w_in2102_0(.douta(w_in2102_0[0]),.doutb(w_in2102_0[1]),.doutc(w_in2102_0[2]),.din(in2[102]));
	jspl3 jspl3_w_in2103_0(.douta(w_in2103_0[0]),.doutb(w_in2103_0[1]),.doutc(w_in2103_0[2]),.din(in2[103]));
	jspl3 jspl3_w_in2104_0(.douta(w_in2104_0[0]),.doutb(w_in2104_0[1]),.doutc(w_in2104_0[2]),.din(in2[104]));
	jspl3 jspl3_w_in2105_0(.douta(w_in2105_0[0]),.doutb(w_in2105_0[1]),.doutc(w_in2105_0[2]),.din(in2[105]));
	jspl3 jspl3_w_in2106_0(.douta(w_in2106_0[0]),.doutb(w_in2106_0[1]),.doutc(w_in2106_0[2]),.din(in2[106]));
	jspl3 jspl3_w_in2107_0(.douta(w_in2107_0[0]),.doutb(w_in2107_0[1]),.doutc(w_in2107_0[2]),.din(in2[107]));
	jspl3 jspl3_w_in2108_0(.douta(w_in2108_0[0]),.doutb(w_in2108_0[1]),.doutc(w_in2108_0[2]),.din(in2[108]));
	jspl3 jspl3_w_in2109_0(.douta(w_in2109_0[0]),.doutb(w_in2109_0[1]),.doutc(w_in2109_0[2]),.din(in2[109]));
	jspl3 jspl3_w_in2110_0(.douta(w_in2110_0[0]),.doutb(w_in2110_0[1]),.doutc(w_in2110_0[2]),.din(in2[110]));
	jspl3 jspl3_w_in2111_0(.douta(w_in2111_0[0]),.doutb(w_in2111_0[1]),.doutc(w_in2111_0[2]),.din(in2[111]));
	jspl3 jspl3_w_in2112_0(.douta(w_in2112_0[0]),.doutb(w_in2112_0[1]),.doutc(w_in2112_0[2]),.din(in2[112]));
	jspl3 jspl3_w_in2113_0(.douta(w_in2113_0[0]),.doutb(w_in2113_0[1]),.doutc(w_in2113_0[2]),.din(in2[113]));
	jspl3 jspl3_w_in2114_0(.douta(w_in2114_0[0]),.doutb(w_in2114_0[1]),.doutc(w_in2114_0[2]),.din(in2[114]));
	jspl3 jspl3_w_in2115_0(.douta(w_in2115_0[0]),.doutb(w_in2115_0[1]),.doutc(w_in2115_0[2]),.din(in2[115]));
	jspl3 jspl3_w_in2116_0(.douta(w_in2116_0[0]),.doutb(w_in2116_0[1]),.doutc(w_in2116_0[2]),.din(in2[116]));
	jspl3 jspl3_w_in2117_0(.douta(w_in2117_0[0]),.doutb(w_in2117_0[1]),.doutc(w_in2117_0[2]),.din(in2[117]));
	jspl3 jspl3_w_in2118_0(.douta(w_in2118_0[0]),.doutb(w_in2118_0[1]),.doutc(w_in2118_0[2]),.din(in2[118]));
	jspl3 jspl3_w_in2119_0(.douta(w_in2119_0[0]),.doutb(w_in2119_0[1]),.doutc(w_in2119_0[2]),.din(in2[119]));
	jspl3 jspl3_w_in2120_0(.douta(w_in2120_0[0]),.doutb(w_in2120_0[1]),.doutc(w_in2120_0[2]),.din(in2[120]));
	jspl3 jspl3_w_in2121_0(.douta(w_in2121_0[0]),.doutb(w_in2121_0[1]),.doutc(w_in2121_0[2]),.din(in2[121]));
	jspl3 jspl3_w_in2122_0(.douta(w_in2122_0[0]),.doutb(w_in2122_0[1]),.doutc(w_in2122_0[2]),.din(in2[122]));
	jspl3 jspl3_w_in2123_0(.douta(w_in2123_0[0]),.doutb(w_in2123_0[1]),.doutc(w_in2123_0[2]),.din(in2[123]));
	jspl3 jspl3_w_in2124_0(.douta(w_in2124_0[0]),.doutb(w_in2124_0[1]),.doutc(w_in2124_0[2]),.din(in2[124]));
	jspl3 jspl3_w_in2125_0(.douta(w_in2125_0[0]),.doutb(w_in2125_0[1]),.doutc(w_in2125_0[2]),.din(in2[125]));
	jspl3 jspl3_w_in2126_0(.douta(w_in2126_0[0]),.doutb(w_in2126_0[1]),.doutc(w_in2126_0[2]),.din(in2[126]));
	jspl3 jspl3_w_in2127_0(.douta(w_in2127_0[0]),.doutb(w_in2127_0[1]),.doutc(w_in2127_0[2]),.din(in2[127]));
	jspl3 jspl3_w_in30_0(.douta(w_in30_0[0]),.doutb(w_in30_0[1]),.doutc(w_in30_0[2]),.din(in3[0]));
	jspl3 jspl3_w_in31_0(.douta(w_in31_0[0]),.doutb(w_in31_0[1]),.doutc(w_in31_0[2]),.din(in3[1]));
	jspl jspl_w_in31_1(.douta(w_in31_1[0]),.doutb(w_in31_1[1]),.din(w_in31_0[0]));
	jspl3 jspl3_w_in32_0(.douta(w_in32_0[0]),.doutb(w_in32_0[1]),.doutc(w_in32_0[2]),.din(in3[2]));
	jspl3 jspl3_w_in33_0(.douta(w_in33_0[0]),.doutb(w_in33_0[1]),.doutc(w_in33_0[2]),.din(in3[3]));
	jspl3 jspl3_w_in34_0(.douta(w_in34_0[0]),.doutb(w_in34_0[1]),.doutc(w_in34_0[2]),.din(in3[4]));
	jspl3 jspl3_w_in35_0(.douta(w_in35_0[0]),.doutb(w_in35_0[1]),.doutc(w_in35_0[2]),.din(in3[5]));
	jspl3 jspl3_w_in36_0(.douta(w_in36_0[0]),.doutb(w_in36_0[1]),.doutc(w_in36_0[2]),.din(in3[6]));
	jspl3 jspl3_w_in37_0(.douta(w_in37_0[0]),.doutb(w_in37_0[1]),.doutc(w_in37_0[2]),.din(in3[7]));
	jspl3 jspl3_w_in38_0(.douta(w_in38_0[0]),.doutb(w_in38_0[1]),.doutc(w_in38_0[2]),.din(in3[8]));
	jspl3 jspl3_w_in39_0(.douta(w_in39_0[0]),.doutb(w_in39_0[1]),.doutc(w_in39_0[2]),.din(in3[9]));
	jspl3 jspl3_w_in310_0(.douta(w_in310_0[0]),.doutb(w_in310_0[1]),.doutc(w_in310_0[2]),.din(in3[10]));
	jspl3 jspl3_w_in311_0(.douta(w_in311_0[0]),.doutb(w_in311_0[1]),.doutc(w_in311_0[2]),.din(in3[11]));
	jspl3 jspl3_w_in312_0(.douta(w_in312_0[0]),.doutb(w_in312_0[1]),.doutc(w_in312_0[2]),.din(in3[12]));
	jspl3 jspl3_w_in313_0(.douta(w_in313_0[0]),.doutb(w_in313_0[1]),.doutc(w_in313_0[2]),.din(in3[13]));
	jspl3 jspl3_w_in314_0(.douta(w_in314_0[0]),.doutb(w_in314_0[1]),.doutc(w_in314_0[2]),.din(in3[14]));
	jspl3 jspl3_w_in315_0(.douta(w_in315_0[0]),.doutb(w_in315_0[1]),.doutc(w_in315_0[2]),.din(in3[15]));
	jspl3 jspl3_w_in316_0(.douta(w_in316_0[0]),.doutb(w_in316_0[1]),.doutc(w_in316_0[2]),.din(in3[16]));
	jspl3 jspl3_w_in317_0(.douta(w_in317_0[0]),.doutb(w_in317_0[1]),.doutc(w_in317_0[2]),.din(in3[17]));
	jspl3 jspl3_w_in318_0(.douta(w_in318_0[0]),.doutb(w_in318_0[1]),.doutc(w_in318_0[2]),.din(in3[18]));
	jspl3 jspl3_w_in319_0(.douta(w_in319_0[0]),.doutb(w_in319_0[1]),.doutc(w_in319_0[2]),.din(in3[19]));
	jspl3 jspl3_w_in320_0(.douta(w_in320_0[0]),.doutb(w_in320_0[1]),.doutc(w_in320_0[2]),.din(in3[20]));
	jspl3 jspl3_w_in321_0(.douta(w_in321_0[0]),.doutb(w_in321_0[1]),.doutc(w_in321_0[2]),.din(in3[21]));
	jspl3 jspl3_w_in322_0(.douta(w_in322_0[0]),.doutb(w_in322_0[1]),.doutc(w_in322_0[2]),.din(in3[22]));
	jspl3 jspl3_w_in323_0(.douta(w_in323_0[0]),.doutb(w_in323_0[1]),.doutc(w_in323_0[2]),.din(in3[23]));
	jspl3 jspl3_w_in324_0(.douta(w_in324_0[0]),.doutb(w_in324_0[1]),.doutc(w_in324_0[2]),.din(in3[24]));
	jspl3 jspl3_w_in325_0(.douta(w_in325_0[0]),.doutb(w_in325_0[1]),.doutc(w_in325_0[2]),.din(in3[25]));
	jspl3 jspl3_w_in326_0(.douta(w_in326_0[0]),.doutb(w_in326_0[1]),.doutc(w_in326_0[2]),.din(in3[26]));
	jspl3 jspl3_w_in327_0(.douta(w_in327_0[0]),.doutb(w_in327_0[1]),.doutc(w_in327_0[2]),.din(in3[27]));
	jspl3 jspl3_w_in328_0(.douta(w_in328_0[0]),.doutb(w_in328_0[1]),.doutc(w_in328_0[2]),.din(in3[28]));
	jspl3 jspl3_w_in329_0(.douta(w_in329_0[0]),.doutb(w_in329_0[1]),.doutc(w_in329_0[2]),.din(in3[29]));
	jspl3 jspl3_w_in330_0(.douta(w_in330_0[0]),.doutb(w_in330_0[1]),.doutc(w_in330_0[2]),.din(in3[30]));
	jspl3 jspl3_w_in331_0(.douta(w_in331_0[0]),.doutb(w_in331_0[1]),.doutc(w_in331_0[2]),.din(in3[31]));
	jspl3 jspl3_w_in332_0(.douta(w_in332_0[0]),.doutb(w_in332_0[1]),.doutc(w_in332_0[2]),.din(in3[32]));
	jspl3 jspl3_w_in333_0(.douta(w_in333_0[0]),.doutb(w_in333_0[1]),.doutc(w_in333_0[2]),.din(in3[33]));
	jspl3 jspl3_w_in334_0(.douta(w_in334_0[0]),.doutb(w_in334_0[1]),.doutc(w_in334_0[2]),.din(in3[34]));
	jspl3 jspl3_w_in335_0(.douta(w_in335_0[0]),.doutb(w_in335_0[1]),.doutc(w_in335_0[2]),.din(in3[35]));
	jspl3 jspl3_w_in336_0(.douta(w_in336_0[0]),.doutb(w_in336_0[1]),.doutc(w_in336_0[2]),.din(in3[36]));
	jspl3 jspl3_w_in337_0(.douta(w_in337_0[0]),.doutb(w_in337_0[1]),.doutc(w_in337_0[2]),.din(in3[37]));
	jspl3 jspl3_w_in338_0(.douta(w_in338_0[0]),.doutb(w_in338_0[1]),.doutc(w_in338_0[2]),.din(in3[38]));
	jspl3 jspl3_w_in339_0(.douta(w_in339_0[0]),.doutb(w_in339_0[1]),.doutc(w_in339_0[2]),.din(in3[39]));
	jspl3 jspl3_w_in340_0(.douta(w_in340_0[0]),.doutb(w_in340_0[1]),.doutc(w_in340_0[2]),.din(in3[40]));
	jspl3 jspl3_w_in341_0(.douta(w_in341_0[0]),.doutb(w_in341_0[1]),.doutc(w_in341_0[2]),.din(in3[41]));
	jspl3 jspl3_w_in342_0(.douta(w_in342_0[0]),.doutb(w_in342_0[1]),.doutc(w_in342_0[2]),.din(in3[42]));
	jspl3 jspl3_w_in343_0(.douta(w_in343_0[0]),.doutb(w_in343_0[1]),.doutc(w_in343_0[2]),.din(in3[43]));
	jspl3 jspl3_w_in344_0(.douta(w_in344_0[0]),.doutb(w_in344_0[1]),.doutc(w_in344_0[2]),.din(in3[44]));
	jspl3 jspl3_w_in345_0(.douta(w_in345_0[0]),.doutb(w_in345_0[1]),.doutc(w_in345_0[2]),.din(in3[45]));
	jspl3 jspl3_w_in346_0(.douta(w_in346_0[0]),.doutb(w_in346_0[1]),.doutc(w_in346_0[2]),.din(in3[46]));
	jspl3 jspl3_w_in347_0(.douta(w_in347_0[0]),.doutb(w_in347_0[1]),.doutc(w_in347_0[2]),.din(in3[47]));
	jspl3 jspl3_w_in348_0(.douta(w_in348_0[0]),.doutb(w_in348_0[1]),.doutc(w_in348_0[2]),.din(in3[48]));
	jspl3 jspl3_w_in349_0(.douta(w_in349_0[0]),.doutb(w_in349_0[1]),.doutc(w_in349_0[2]),.din(in3[49]));
	jspl3 jspl3_w_in350_0(.douta(w_in350_0[0]),.doutb(w_in350_0[1]),.doutc(w_in350_0[2]),.din(in3[50]));
	jspl3 jspl3_w_in351_0(.douta(w_in351_0[0]),.doutb(w_in351_0[1]),.doutc(w_in351_0[2]),.din(in3[51]));
	jspl jspl_w_in352_0(.douta(w_in352_0[0]),.doutb(w_in352_0[1]),.din(in3[52]));
	jspl3 jspl3_w_in353_0(.douta(w_in353_0[0]),.doutb(w_in353_0[1]),.doutc(w_in353_0[2]),.din(in3[53]));
	jspl3 jspl3_w_in354_0(.douta(w_in354_0[0]),.doutb(w_in354_0[1]),.doutc(w_in354_0[2]),.din(in3[54]));
	jspl3 jspl3_w_in355_0(.douta(w_in355_0[0]),.doutb(w_in355_0[1]),.doutc(w_in355_0[2]),.din(in3[55]));
	jspl3 jspl3_w_in356_0(.douta(w_in356_0[0]),.doutb(w_in356_0[1]),.doutc(w_in356_0[2]),.din(in3[56]));
	jspl3 jspl3_w_in357_0(.douta(w_in357_0[0]),.doutb(w_in357_0[1]),.doutc(w_in357_0[2]),.din(in3[57]));
	jspl3 jspl3_w_in358_0(.douta(w_in358_0[0]),.doutb(w_in358_0[1]),.doutc(w_in358_0[2]),.din(in3[58]));
	jspl3 jspl3_w_in359_0(.douta(w_in359_0[0]),.doutb(w_in359_0[1]),.doutc(w_in359_0[2]),.din(in3[59]));
	jspl3 jspl3_w_in360_0(.douta(w_in360_0[0]),.doutb(w_in360_0[1]),.doutc(w_in360_0[2]),.din(in3[60]));
	jspl3 jspl3_w_in361_0(.douta(w_in361_0[0]),.doutb(w_in361_0[1]),.doutc(w_in361_0[2]),.din(in3[61]));
	jspl3 jspl3_w_in362_0(.douta(w_in362_0[0]),.doutb(w_in362_0[1]),.doutc(w_in362_0[2]),.din(in3[62]));
	jspl3 jspl3_w_in363_0(.douta(w_in363_0[0]),.doutb(w_in363_0[1]),.doutc(w_in363_0[2]),.din(in3[63]));
	jspl3 jspl3_w_in364_0(.douta(w_in364_0[0]),.doutb(w_in364_0[1]),.doutc(w_in364_0[2]),.din(in3[64]));
	jspl3 jspl3_w_in365_0(.douta(w_in365_0[0]),.doutb(w_in365_0[1]),.doutc(w_in365_0[2]),.din(in3[65]));
	jspl3 jspl3_w_in366_0(.douta(w_in366_0[0]),.doutb(w_in366_0[1]),.doutc(w_in366_0[2]),.din(in3[66]));
	jspl3 jspl3_w_in367_0(.douta(w_in367_0[0]),.doutb(w_in367_0[1]),.doutc(w_in367_0[2]),.din(in3[67]));
	jspl3 jspl3_w_in368_0(.douta(w_in368_0[0]),.doutb(w_in368_0[1]),.doutc(w_in368_0[2]),.din(in3[68]));
	jspl3 jspl3_w_in369_0(.douta(w_in369_0[0]),.doutb(w_in369_0[1]),.doutc(w_in369_0[2]),.din(in3[69]));
	jspl3 jspl3_w_in370_0(.douta(w_in370_0[0]),.doutb(w_in370_0[1]),.doutc(w_in370_0[2]),.din(in3[70]));
	jspl3 jspl3_w_in371_0(.douta(w_in371_0[0]),.doutb(w_in371_0[1]),.doutc(w_in371_0[2]),.din(in3[71]));
	jspl3 jspl3_w_in372_0(.douta(w_in372_0[0]),.doutb(w_in372_0[1]),.doutc(w_in372_0[2]),.din(in3[72]));
	jspl3 jspl3_w_in373_0(.douta(w_in373_0[0]),.doutb(w_in373_0[1]),.doutc(w_in373_0[2]),.din(in3[73]));
	jspl3 jspl3_w_in374_0(.douta(w_in374_0[0]),.doutb(w_in374_0[1]),.doutc(w_in374_0[2]),.din(in3[74]));
	jspl3 jspl3_w_in375_0(.douta(w_in375_0[0]),.doutb(w_in375_0[1]),.doutc(w_in375_0[2]),.din(in3[75]));
	jspl3 jspl3_w_in376_0(.douta(w_in376_0[0]),.doutb(w_in376_0[1]),.doutc(w_in376_0[2]),.din(in3[76]));
	jspl3 jspl3_w_in377_0(.douta(w_in377_0[0]),.doutb(w_in377_0[1]),.doutc(w_in377_0[2]),.din(in3[77]));
	jspl3 jspl3_w_in378_0(.douta(w_in378_0[0]),.doutb(w_in378_0[1]),.doutc(w_in378_0[2]),.din(in3[78]));
	jspl3 jspl3_w_in379_0(.douta(w_in379_0[0]),.doutb(w_in379_0[1]),.doutc(w_in379_0[2]),.din(in3[79]));
	jspl3 jspl3_w_in380_0(.douta(w_in380_0[0]),.doutb(w_in380_0[1]),.doutc(w_in380_0[2]),.din(in3[80]));
	jspl3 jspl3_w_in381_0(.douta(w_in381_0[0]),.doutb(w_in381_0[1]),.doutc(w_in381_0[2]),.din(in3[81]));
	jspl3 jspl3_w_in382_0(.douta(w_in382_0[0]),.doutb(w_in382_0[1]),.doutc(w_in382_0[2]),.din(in3[82]));
	jspl3 jspl3_w_in383_0(.douta(w_in383_0[0]),.doutb(w_in383_0[1]),.doutc(w_in383_0[2]),.din(in3[83]));
	jspl3 jspl3_w_in384_0(.douta(w_in384_0[0]),.doutb(w_in384_0[1]),.doutc(w_in384_0[2]),.din(in3[84]));
	jspl3 jspl3_w_in385_0(.douta(w_in385_0[0]),.doutb(w_in385_0[1]),.doutc(w_in385_0[2]),.din(in3[85]));
	jspl3 jspl3_w_in386_0(.douta(w_in386_0[0]),.doutb(w_in386_0[1]),.doutc(w_in386_0[2]),.din(in3[86]));
	jspl3 jspl3_w_in387_0(.douta(w_in387_0[0]),.doutb(w_in387_0[1]),.doutc(w_in387_0[2]),.din(in3[87]));
	jspl3 jspl3_w_in388_0(.douta(w_in388_0[0]),.doutb(w_in388_0[1]),.doutc(w_in388_0[2]),.din(in3[88]));
	jspl3 jspl3_w_in389_0(.douta(w_in389_0[0]),.doutb(w_in389_0[1]),.doutc(w_in389_0[2]),.din(in3[89]));
	jspl3 jspl3_w_in390_0(.douta(w_in390_0[0]),.doutb(w_in390_0[1]),.doutc(w_in390_0[2]),.din(in3[90]));
	jspl3 jspl3_w_in391_0(.douta(w_in391_0[0]),.doutb(w_in391_0[1]),.doutc(w_in391_0[2]),.din(in3[91]));
	jspl3 jspl3_w_in392_0(.douta(w_in392_0[0]),.doutb(w_in392_0[1]),.doutc(w_in392_0[2]),.din(in3[92]));
	jspl3 jspl3_w_in393_0(.douta(w_in393_0[0]),.doutb(w_in393_0[1]),.doutc(w_in393_0[2]),.din(in3[93]));
	jspl3 jspl3_w_in394_0(.douta(w_in394_0[0]),.doutb(w_in394_0[1]),.doutc(w_in394_0[2]),.din(in3[94]));
	jspl3 jspl3_w_in395_0(.douta(w_in395_0[0]),.doutb(w_in395_0[1]),.doutc(w_in395_0[2]),.din(in3[95]));
	jspl3 jspl3_w_in396_0(.douta(w_in396_0[0]),.doutb(w_in396_0[1]),.doutc(w_in396_0[2]),.din(in3[96]));
	jspl3 jspl3_w_in397_0(.douta(w_in397_0[0]),.doutb(w_in397_0[1]),.doutc(w_in397_0[2]),.din(in3[97]));
	jspl3 jspl3_w_in398_0(.douta(w_in398_0[0]),.doutb(w_in398_0[1]),.doutc(w_in398_0[2]),.din(in3[98]));
	jspl3 jspl3_w_in399_0(.douta(w_in399_0[0]),.doutb(w_in399_0[1]),.doutc(w_in399_0[2]),.din(in3[99]));
	jspl3 jspl3_w_in3100_0(.douta(w_in3100_0[0]),.doutb(w_in3100_0[1]),.doutc(w_in3100_0[2]),.din(in3[100]));
	jspl3 jspl3_w_in3101_0(.douta(w_in3101_0[0]),.doutb(w_in3101_0[1]),.doutc(w_in3101_0[2]),.din(in3[101]));
	jspl3 jspl3_w_in3102_0(.douta(w_in3102_0[0]),.doutb(w_in3102_0[1]),.doutc(w_in3102_0[2]),.din(in3[102]));
	jspl3 jspl3_w_in3103_0(.douta(w_in3103_0[0]),.doutb(w_in3103_0[1]),.doutc(w_in3103_0[2]),.din(in3[103]));
	jspl3 jspl3_w_in3104_0(.douta(w_in3104_0[0]),.doutb(w_in3104_0[1]),.doutc(w_in3104_0[2]),.din(in3[104]));
	jspl3 jspl3_w_in3105_0(.douta(w_in3105_0[0]),.doutb(w_in3105_0[1]),.doutc(w_in3105_0[2]),.din(in3[105]));
	jspl3 jspl3_w_in3106_0(.douta(w_in3106_0[0]),.doutb(w_in3106_0[1]),.doutc(w_in3106_0[2]),.din(in3[106]));
	jspl3 jspl3_w_in3107_0(.douta(w_in3107_0[0]),.doutb(w_in3107_0[1]),.doutc(w_in3107_0[2]),.din(in3[107]));
	jspl3 jspl3_w_in3108_0(.douta(w_in3108_0[0]),.doutb(w_in3108_0[1]),.doutc(w_in3108_0[2]),.din(in3[108]));
	jspl3 jspl3_w_in3109_0(.douta(w_in3109_0[0]),.doutb(w_in3109_0[1]),.doutc(w_in3109_0[2]),.din(in3[109]));
	jspl3 jspl3_w_in3110_0(.douta(w_in3110_0[0]),.doutb(w_in3110_0[1]),.doutc(w_in3110_0[2]),.din(in3[110]));
	jspl3 jspl3_w_in3111_0(.douta(w_in3111_0[0]),.doutb(w_in3111_0[1]),.doutc(w_in3111_0[2]),.din(in3[111]));
	jspl3 jspl3_w_in3112_0(.douta(w_in3112_0[0]),.doutb(w_in3112_0[1]),.doutc(w_in3112_0[2]),.din(in3[112]));
	jspl3 jspl3_w_in3113_0(.douta(w_in3113_0[0]),.doutb(w_in3113_0[1]),.doutc(w_in3113_0[2]),.din(in3[113]));
	jspl3 jspl3_w_in3114_0(.douta(w_in3114_0[0]),.doutb(w_in3114_0[1]),.doutc(w_in3114_0[2]),.din(in3[114]));
	jspl3 jspl3_w_in3115_0(.douta(w_in3115_0[0]),.doutb(w_in3115_0[1]),.doutc(w_in3115_0[2]),.din(in3[115]));
	jspl3 jspl3_w_in3116_0(.douta(w_in3116_0[0]),.doutb(w_in3116_0[1]),.doutc(w_in3116_0[2]),.din(in3[116]));
	jspl3 jspl3_w_in3117_0(.douta(w_in3117_0[0]),.doutb(w_in3117_0[1]),.doutc(w_in3117_0[2]),.din(in3[117]));
	jspl3 jspl3_w_in3118_0(.douta(w_in3118_0[0]),.doutb(w_in3118_0[1]),.doutc(w_in3118_0[2]),.din(in3[118]));
	jspl3 jspl3_w_in3119_0(.douta(w_in3119_0[0]),.doutb(w_in3119_0[1]),.doutc(w_in3119_0[2]),.din(in3[119]));
	jspl3 jspl3_w_in3120_0(.douta(w_in3120_0[0]),.doutb(w_in3120_0[1]),.doutc(w_in3120_0[2]),.din(in3[120]));
	jspl3 jspl3_w_in3121_0(.douta(w_in3121_0[0]),.doutb(w_in3121_0[1]),.doutc(w_in3121_0[2]),.din(in3[121]));
	jspl3 jspl3_w_in3122_0(.douta(w_in3122_0[0]),.doutb(w_in3122_0[1]),.doutc(w_in3122_0[2]),.din(in3[122]));
	jspl3 jspl3_w_in3123_0(.douta(w_in3123_0[0]),.doutb(w_in3123_0[1]),.doutc(w_in3123_0[2]),.din(in3[123]));
	jspl3 jspl3_w_in3124_0(.douta(w_in3124_0[0]),.doutb(w_in3124_0[1]),.doutc(w_in3124_0[2]),.din(in3[124]));
	jspl3 jspl3_w_in3125_0(.douta(w_in3125_0[0]),.doutb(w_in3125_0[1]),.doutc(w_in3125_0[2]),.din(in3[125]));
	jspl3 jspl3_w_in3126_0(.douta(w_in3126_0[0]),.doutb(w_in3126_0[1]),.doutc(w_in3126_0[2]),.din(in3[126]));
	jspl3 jspl3_w_in3127_0(.douta(w_in3127_0[0]),.doutb(w_in3127_0[1]),.doutc(w_in3127_0[2]),.din(in3[127]));
	jspl3 jspl3_w_address1_0(.douta(w_address1_0[0]),.doutb(w_address1_0[1]),.doutc(w_address1_0[2]),.din(address_fa_1));
	jspl3 jspl3_w_address1_1(.douta(w_address1_1[0]),.doutb(w_address1_1[1]),.doutc(w_address1_1[2]),.din(w_address1_0[0]));
	jspl3 jspl3_w_address1_2(.douta(w_address1_2[0]),.doutb(w_address1_2[1]),.doutc(w_address1_2[2]),.din(w_address1_0[1]));
	jspl3 jspl3_w_address1_3(.douta(w_address1_3[0]),.doutb(w_address1_3[1]),.doutc(w_address1_3[2]),.din(w_address1_0[2]));
	jspl3 jspl3_w_address1_4(.douta(w_address1_4[0]),.doutb(w_address1_4[1]),.doutc(w_address1_4[2]),.din(w_address1_1[0]));
	jspl3 jspl3_w_address1_5(.douta(w_address1_5[0]),.doutb(w_address1_5[1]),.doutc(w_address1_5[2]),.din(w_address1_1[1]));
	jspl3 jspl3_w_address1_6(.douta(w_address1_6[0]),.doutb(w_address1_6[1]),.doutc(w_address1_6[2]),.din(w_address1_1[2]));
	jspl3 jspl3_w_address1_7(.douta(w_address1_7[0]),.doutb(w_address1_7[1]),.doutc(w_address1_7[2]),.din(w_address1_2[0]));
	jspl3 jspl3_w_address1_8(.douta(w_address1_8[0]),.doutb(w_address1_8[1]),.doutc(w_address1_8[2]),.din(w_address1_2[1]));
	jspl3 jspl3_w_address1_9(.douta(w_address1_9[0]),.doutb(w_address1_9[1]),.doutc(w_address1_9[2]),.din(w_address1_2[2]));
	jspl3 jspl3_w_address1_10(.douta(w_address1_10[0]),.doutb(w_address1_10[1]),.doutc(w_address1_10[2]),.din(w_address1_3[0]));
	jspl3 jspl3_w_address1_11(.douta(w_address1_11[0]),.doutb(w_address1_11[1]),.doutc(w_address1_11[2]),.din(w_address1_3[1]));
	jspl3 jspl3_w_address1_12(.douta(w_address1_12[0]),.doutb(w_address1_12[1]),.doutc(w_address1_12[2]),.din(w_address1_3[2]));
	jspl3 jspl3_w_address1_13(.douta(w_address1_13[0]),.doutb(w_address1_13[1]),.doutc(w_address1_13[2]),.din(w_address1_4[0]));
	jspl3 jspl3_w_address1_14(.douta(w_address1_14[0]),.doutb(w_address1_14[1]),.doutc(w_address1_14[2]),.din(w_address1_4[1]));
	jspl3 jspl3_w_address1_15(.douta(w_address1_15[0]),.doutb(w_address1_15[1]),.doutc(w_address1_15[2]),.din(w_address1_4[2]));
	jspl3 jspl3_w_address1_16(.douta(w_address1_16[0]),.doutb(w_address1_16[1]),.doutc(w_address1_16[2]),.din(w_address1_5[0]));
	jspl3 jspl3_w_address1_17(.douta(w_address1_17[0]),.doutb(w_address1_17[1]),.doutc(w_address1_17[2]),.din(w_address1_5[1]));
	jspl3 jspl3_w_address1_18(.douta(w_address1_18[0]),.doutb(w_address1_18[1]),.doutc(w_address1_18[2]),.din(w_address1_5[2]));
	jspl3 jspl3_w_address1_19(.douta(w_address1_19[0]),.doutb(w_address1_19[1]),.doutc(w_address1_19[2]),.din(w_address1_6[0]));
	jspl3 jspl3_w_address1_20(.douta(w_address1_20[0]),.doutb(w_address1_20[1]),.doutc(w_address1_20[2]),.din(w_address1_6[1]));
	jspl3 jspl3_w_address1_21(.douta(w_address1_21[0]),.doutb(w_address1_21[1]),.doutc(w_address1_21[2]),.din(w_address1_6[2]));
	jspl3 jspl3_w_address1_22(.douta(w_address1_22[0]),.doutb(w_address1_22[1]),.doutc(w_address1_22[2]),.din(w_address1_7[0]));
	jspl3 jspl3_w_address1_23(.douta(w_address1_23[0]),.doutb(w_address1_23[1]),.doutc(w_address1_23[2]),.din(w_address1_7[1]));
	jspl3 jspl3_w_address1_24(.douta(w_address1_24[0]),.doutb(w_address1_24[1]),.doutc(w_address1_24[2]),.din(w_address1_7[2]));
	jspl3 jspl3_w_address1_25(.douta(w_address1_25[0]),.doutb(w_address1_25[1]),.doutc(w_address1_25[2]),.din(w_address1_8[0]));
	jspl3 jspl3_w_address1_26(.douta(w_address1_26[0]),.doutb(w_address1_26[1]),.doutc(w_address1_26[2]),.din(w_address1_8[1]));
	jspl3 jspl3_w_address1_27(.douta(w_address1_27[0]),.doutb(w_address1_27[1]),.doutc(w_address1_27[2]),.din(w_address1_8[2]));
	jspl3 jspl3_w_address1_28(.douta(w_address1_28[0]),.doutb(w_address1_28[1]),.doutc(w_address1_28[2]),.din(w_address1_9[0]));
	jspl3 jspl3_w_address1_29(.douta(w_address1_29[0]),.doutb(w_address1_29[1]),.doutc(w_address1_29[2]),.din(w_address1_9[1]));
	jspl3 jspl3_w_address1_30(.douta(w_address1_30[0]),.doutb(w_address1_30[1]),.doutc(w_address1_30[2]),.din(w_address1_9[2]));
	jspl3 jspl3_w_address1_31(.douta(w_address1_31[0]),.doutb(w_address1_31[1]),.doutc(w_address1_31[2]),.din(w_address1_10[0]));
	jspl3 jspl3_w_address1_32(.douta(w_address1_32[0]),.doutb(w_address1_32[1]),.doutc(w_address1_32[2]),.din(w_address1_10[1]));
	jspl3 jspl3_w_address1_33(.douta(w_address1_33[0]),.doutb(w_address1_33[1]),.doutc(w_address1_33[2]),.din(w_address1_10[2]));
	jspl3 jspl3_w_address1_34(.douta(w_address1_34[0]),.doutb(w_address1_34[1]),.doutc(w_address1_34[2]),.din(w_address1_11[0]));
	jspl3 jspl3_w_address1_35(.douta(w_address1_35[0]),.doutb(w_address1_35[1]),.doutc(w_address1_35[2]),.din(w_address1_11[1]));
	jspl3 jspl3_w_address1_36(.douta(w_address1_36[0]),.doutb(w_address1_36[1]),.doutc(w_address1_36[2]),.din(w_address1_11[2]));
	jspl3 jspl3_w_address1_37(.douta(w_address1_37[0]),.doutb(w_address1_37[1]),.doutc(w_address1_37[2]),.din(w_address1_12[0]));
	jspl3 jspl3_w_address1_38(.douta(w_address1_38[0]),.doutb(w_address1_38[1]),.doutc(w_address1_38[2]),.din(w_address1_12[1]));
	jspl3 jspl3_w_address1_39(.douta(w_address1_39[0]),.doutb(w_address1_39[1]),.doutc(w_address1_39[2]),.din(w_address1_12[2]));
	jspl3 jspl3_w_address1_40(.douta(w_address1_40[0]),.doutb(w_address1_40[1]),.doutc(w_address1_40[2]),.din(w_address1_13[0]));
	jspl3 jspl3_w_address1_41(.douta(w_address1_41[0]),.doutb(w_address1_41[1]),.doutc(w_address1_41[2]),.din(w_address1_13[1]));
	jspl3 jspl3_w_address1_42(.douta(w_address1_42[0]),.doutb(w_address1_42[1]),.doutc(w_address1_42[2]),.din(w_address1_13[2]));
	jspl3 jspl3_w_address1_43(.douta(w_address1_43[0]),.doutb(w_address1_43[1]),.doutc(w_address1_43[2]),.din(w_address1_14[0]));
	jspl3 jspl3_w_address1_44(.douta(w_address1_44[0]),.doutb(w_address1_44[1]),.doutc(w_address1_44[2]),.din(w_address1_14[1]));
	jspl3 jspl3_w_address1_45(.douta(w_address1_45[0]),.doutb(w_address1_45[1]),.doutc(w_address1_45[2]),.din(w_address1_14[2]));
	jspl3 jspl3_w_address1_46(.douta(w_address1_46[0]),.doutb(w_address1_46[1]),.doutc(w_address1_46[2]),.din(w_address1_15[0]));
	jspl3 jspl3_w_address1_47(.douta(w_address1_47[0]),.doutb(w_address1_47[1]),.doutc(w_address1_47[2]),.din(w_address1_15[1]));
	jspl3 jspl3_w_address1_48(.douta(w_address1_48[0]),.doutb(w_address1_48[1]),.doutc(w_address1_48[2]),.din(w_address1_15[2]));
	jspl3 jspl3_w_address1_49(.douta(w_address1_49[0]),.doutb(w_address1_49[1]),.doutc(w_address1_49[2]),.din(w_address1_16[0]));
	jspl3 jspl3_w_address1_50(.douta(w_address1_50[0]),.doutb(w_address1_50[1]),.doutc(w_address1_50[2]),.din(w_address1_16[1]));
	jspl3 jspl3_w_address1_51(.douta(w_address1_51[0]),.doutb(w_address1_51[1]),.doutc(w_address1_51[2]),.din(w_address1_16[2]));
	jspl3 jspl3_w_address1_52(.douta(w_address1_52[0]),.doutb(w_address1_52[1]),.doutc(w_address1_52[2]),.din(w_address1_17[0]));
	jspl3 jspl3_w_address1_53(.douta(w_address1_53[0]),.doutb(w_address1_53[1]),.doutc(w_address1_53[2]),.din(w_address1_17[1]));
	jspl3 jspl3_w_address1_54(.douta(w_address1_54[0]),.doutb(w_address1_54[1]),.doutc(w_address1_54[2]),.din(w_address1_17[2]));
	jspl3 jspl3_w_address1_55(.douta(w_address1_55[0]),.doutb(w_address1_55[1]),.doutc(w_address1_55[2]),.din(w_address1_18[0]));
	jspl3 jspl3_w_address1_56(.douta(w_address1_56[0]),.doutb(w_address1_56[1]),.doutc(w_address1_56[2]),.din(w_address1_18[1]));
	jspl3 jspl3_w_address1_57(.douta(w_address1_57[0]),.doutb(w_address1_57[1]),.doutc(w_address1_57[2]),.din(w_address1_18[2]));
	jspl3 jspl3_w_address1_58(.douta(w_address1_58[0]),.doutb(w_address1_58[1]),.doutc(w_address1_58[2]),.din(w_address1_19[0]));
	jspl3 jspl3_w_address1_59(.douta(w_address1_59[0]),.doutb(w_address1_59[1]),.doutc(w_address1_59[2]),.din(w_address1_19[1]));
	jspl3 jspl3_w_address1_60(.douta(w_address1_60[0]),.doutb(w_address1_60[1]),.doutc(w_address1_60[2]),.din(w_address1_19[2]));
	jspl3 jspl3_w_address1_61(.douta(w_address1_61[0]),.doutb(w_address1_61[1]),.doutc(w_address1_61[2]),.din(w_address1_20[0]));
	jspl3 jspl3_w_address1_62(.douta(w_address1_62[0]),.doutb(w_address1_62[1]),.doutc(w_address1_62[2]),.din(w_address1_20[1]));
	jspl3 jspl3_w_address1_63(.douta(w_address1_63[0]),.doutb(w_address1_63[1]),.doutc(address[0]),.din(w_address1_20[2]));
	jspl jspl_w_n643_0(.douta(w_n643_0[0]),.doutb(w_n643_0[1]),.din(n643));
	jspl jspl_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.din(n646));
	jspl jspl_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.din(n648));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.din(n653));
	jspl jspl_w_n656_0(.douta(w_n656_0[0]),.doutb(w_n656_0[1]),.din(n656));
	jspl jspl_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.din(n658));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.din(n663));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n668_0(.douta(w_n668_0[0]),.doutb(w_n668_0[1]),.din(n668));
	jspl jspl_w_n671_0(.douta(w_n671_0[0]),.doutb(w_n671_0[1]),.din(n671));
	jspl jspl_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.din(n673));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n688_0(.douta(w_n688_0[0]),.doutb(w_n688_0[1]),.din(n688));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(n696));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl jspl_w_n731_0(.douta(w_n731_0[0]),.doutb(w_n731_0[1]),.din(n731));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl jspl_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.din(n743));
	jspl jspl_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.din(n746));
	jspl jspl_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.din(n748));
	jspl jspl_w_n751_0(.douta(w_n751_0[0]),.doutb(w_n751_0[1]),.din(n751));
	jspl jspl_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.din(n753));
	jspl jspl_w_n756_0(.douta(w_n756_0[0]),.doutb(w_n756_0[1]),.din(n756));
	jspl jspl_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.din(n758));
	jspl jspl_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.din(n761));
	jspl jspl_w_n763_0(.douta(w_n763_0[0]),.doutb(w_n763_0[1]),.din(n763));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(n766));
	jspl jspl_w_n768_0(.douta(w_n768_0[0]),.doutb(w_n768_0[1]),.din(n768));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n776_0(.douta(w_n776_0[0]),.doutb(w_n776_0[1]),.din(n776));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(n781));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.din(n783));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl jspl_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.din(n853));
	jspl jspl_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.din(n858));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(n915));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_n931_0[1]),.din(n931));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(n939));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.din(n980));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(n988));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.din(n1032));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(n1037));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.din(n1046));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(n1048));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(n1091));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(n1103));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(n1127));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1132_0(.douta(w_n1132_0[0]),.doutb(w_n1132_0[1]),.din(n1132));
	jspl jspl_w_n1149_0(.douta(w_n1149_0[0]),.doutb(w_n1149_0[1]),.din(n1149));
	jspl jspl_w_n1155_0(.douta(w_n1155_0[0]),.doutb(w_n1155_0[1]),.din(n1155));
	jspl jspl_w_n1157_0(.douta(w_n1157_0[0]),.doutb(w_n1157_0[1]),.din(n1157));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(n1161));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(n1178));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(n1190));
	jspl jspl_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.din(n1207));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(n1215));
	jspl jspl_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.din(n1219));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1243_0(.douta(w_n1243_0[0]),.doutb(w_n1243_0[1]),.din(n1243));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(n1247));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(n1248));
	jspl jspl_w_n1265_0(.douta(w_n1265_0[0]),.doutb(w_n1265_0[1]),.din(n1265));
	jspl jspl_w_n1271_0(.douta(w_n1271_0[0]),.doutb(w_n1271_0[1]),.din(n1271));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(n1273));
	jspl jspl_w_n1277_0(.douta(w_n1277_0[0]),.doutb(w_n1277_0[1]),.din(n1277));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_n1294_0[1]),.din(n1294));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1323_0(.douta(w_n1323_0[0]),.doutb(w_n1323_0[1]),.din(n1323));
	jspl jspl_w_n1329_0(.douta(w_n1329_0[0]),.doutb(w_n1329_0[1]),.din(n1329));
	jspl jspl_w_n1331_0(.douta(w_n1331_0[0]),.doutb(w_n1331_0[1]),.din(n1331));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(n1352));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(n1364));
	jspl jspl_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.din(n1381));
	jspl jspl_w_n1387_0(.douta(w_n1387_0[0]),.doutb(w_n1387_0[1]),.din(n1387));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1417_0(.douta(w_n1417_0[0]),.doutb(w_n1417_0[1]),.din(n1417));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1422_0(.douta(w_n1422_0[0]),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1475_0(.douta(w_n1475_0[0]),.doutb(w_n1475_0[1]),.din(n1475));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1497_0(.douta(w_n1497_0[0]),.doutb(w_n1497_0[1]),.din(n1497));
	jspl jspl_w_n1503_0(.douta(w_n1503_0[0]),.doutb(w_n1503_0[1]),.din(n1503));
	jspl jspl_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.din(n1505));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1526_0(.douta(w_n1526_0[0]),.doutb(w_n1526_0[1]),.din(n1526));
	jspl jspl_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.din(n1532));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(n1555));
	jspl3 jspl3_w_n1556_0(.douta(w_n1556_0[0]),.doutb(w_n1556_0[1]),.doutc(w_n1556_0[2]),.din(n1556));
	jspl3 jspl3_w_n1556_1(.douta(w_n1556_1[0]),.doutb(w_n1556_1[1]),.doutc(w_n1556_1[2]),.din(w_n1556_0[0]));
	jspl3 jspl3_w_n1556_2(.douta(w_n1556_2[0]),.doutb(w_n1556_2[1]),.doutc(w_n1556_2[2]),.din(w_n1556_0[1]));
	jspl3 jspl3_w_n1556_3(.douta(w_n1556_3[0]),.doutb(w_n1556_3[1]),.doutc(w_n1556_3[2]),.din(w_n1556_0[2]));
	jspl3 jspl3_w_n1556_4(.douta(w_n1556_4[0]),.doutb(w_n1556_4[1]),.doutc(w_n1556_4[2]),.din(w_n1556_1[0]));
	jspl3 jspl3_w_n1556_5(.douta(w_n1556_5[0]),.doutb(w_n1556_5[1]),.doutc(w_n1556_5[2]),.din(w_n1556_1[1]));
	jspl3 jspl3_w_n1556_6(.douta(w_n1556_6[0]),.doutb(w_n1556_6[1]),.doutc(w_n1556_6[2]),.din(w_n1556_1[2]));
	jspl3 jspl3_w_n1556_7(.douta(w_n1556_7[0]),.doutb(w_n1556_7[1]),.doutc(w_n1556_7[2]),.din(w_n1556_2[0]));
	jspl3 jspl3_w_n1556_8(.douta(w_n1556_8[0]),.doutb(w_n1556_8[1]),.doutc(w_n1556_8[2]),.din(w_n1556_2[1]));
	jspl3 jspl3_w_n1556_9(.douta(w_n1556_9[0]),.doutb(w_n1556_9[1]),.doutc(w_n1556_9[2]),.din(w_n1556_2[2]));
	jspl3 jspl3_w_n1556_10(.douta(w_n1556_10[0]),.doutb(w_n1556_10[1]),.doutc(w_n1556_10[2]),.din(w_n1556_3[0]));
	jspl3 jspl3_w_n1556_11(.douta(w_n1556_11[0]),.doutb(w_n1556_11[1]),.doutc(w_n1556_11[2]),.din(w_n1556_3[1]));
	jspl3 jspl3_w_n1556_12(.douta(w_n1556_12[0]),.doutb(w_n1556_12[1]),.doutc(w_n1556_12[2]),.din(w_n1556_3[2]));
	jspl3 jspl3_w_n1556_13(.douta(w_n1556_13[0]),.doutb(w_n1556_13[1]),.doutc(w_n1556_13[2]),.din(w_n1556_4[0]));
	jspl3 jspl3_w_n1556_14(.douta(w_n1556_14[0]),.doutb(w_n1556_14[1]),.doutc(w_n1556_14[2]),.din(w_n1556_4[1]));
	jspl3 jspl3_w_n1556_15(.douta(w_n1556_15[0]),.doutb(w_n1556_15[1]),.doutc(w_n1556_15[2]),.din(w_n1556_4[2]));
	jspl3 jspl3_w_n1556_16(.douta(w_n1556_16[0]),.doutb(w_n1556_16[1]),.doutc(w_n1556_16[2]),.din(w_n1556_5[0]));
	jspl3 jspl3_w_n1556_17(.douta(w_n1556_17[0]),.doutb(w_n1556_17[1]),.doutc(w_n1556_17[2]),.din(w_n1556_5[1]));
	jspl3 jspl3_w_n1556_18(.douta(w_n1556_18[0]),.doutb(w_n1556_18[1]),.doutc(w_n1556_18[2]),.din(w_n1556_5[2]));
	jspl3 jspl3_w_n1556_19(.douta(w_n1556_19[0]),.doutb(w_n1556_19[1]),.doutc(w_n1556_19[2]),.din(w_n1556_6[0]));
	jspl3 jspl3_w_n1556_20(.douta(w_n1556_20[0]),.doutb(w_n1556_20[1]),.doutc(w_n1556_20[2]),.din(w_n1556_6[1]));
	jspl3 jspl3_w_n1556_21(.douta(w_n1556_21[0]),.doutb(w_n1556_21[1]),.doutc(w_n1556_21[2]),.din(w_n1556_6[2]));
	jspl3 jspl3_w_n1556_22(.douta(w_n1556_22[0]),.doutb(w_n1556_22[1]),.doutc(w_n1556_22[2]),.din(w_n1556_7[0]));
	jspl3 jspl3_w_n1556_23(.douta(w_n1556_23[0]),.doutb(w_n1556_23[1]),.doutc(w_n1556_23[2]),.din(w_n1556_7[1]));
	jspl3 jspl3_w_n1556_24(.douta(w_n1556_24[0]),.doutb(w_n1556_24[1]),.doutc(w_n1556_24[2]),.din(w_n1556_7[2]));
	jspl3 jspl3_w_n1556_25(.douta(w_n1556_25[0]),.doutb(w_n1556_25[1]),.doutc(w_n1556_25[2]),.din(w_n1556_8[0]));
	jspl3 jspl3_w_n1556_26(.douta(w_n1556_26[0]),.doutb(w_n1556_26[1]),.doutc(w_n1556_26[2]),.din(w_n1556_8[1]));
	jspl3 jspl3_w_n1556_27(.douta(w_n1556_27[0]),.doutb(w_n1556_27[1]),.doutc(w_n1556_27[2]),.din(w_n1556_8[2]));
	jspl3 jspl3_w_n1556_28(.douta(w_n1556_28[0]),.doutb(w_n1556_28[1]),.doutc(w_n1556_28[2]),.din(w_n1556_9[0]));
	jspl3 jspl3_w_n1556_29(.douta(w_n1556_29[0]),.doutb(w_n1556_29[1]),.doutc(w_n1556_29[2]),.din(w_n1556_9[1]));
	jspl3 jspl3_w_n1556_30(.douta(w_n1556_30[0]),.doutb(w_n1556_30[1]),.doutc(w_n1556_30[2]),.din(w_n1556_9[2]));
	jspl3 jspl3_w_n1556_31(.douta(w_n1556_31[0]),.doutb(w_n1556_31[1]),.doutc(w_n1556_31[2]),.din(w_n1556_10[0]));
	jspl3 jspl3_w_n1556_32(.douta(w_n1556_32[0]),.doutb(w_n1556_32[1]),.doutc(w_n1556_32[2]),.din(w_n1556_10[1]));
	jspl3 jspl3_w_n1556_33(.douta(w_n1556_33[0]),.doutb(w_n1556_33[1]),.doutc(w_n1556_33[2]),.din(w_n1556_10[2]));
	jspl3 jspl3_w_n1556_34(.douta(w_n1556_34[0]),.doutb(w_n1556_34[1]),.doutc(w_n1556_34[2]),.din(w_n1556_11[0]));
	jspl3 jspl3_w_n1556_35(.douta(w_n1556_35[0]),.doutb(w_n1556_35[1]),.doutc(w_n1556_35[2]),.din(w_n1556_11[1]));
	jspl3 jspl3_w_n1556_36(.douta(w_n1556_36[0]),.doutb(w_n1556_36[1]),.doutc(w_n1556_36[2]),.din(w_n1556_11[2]));
	jspl3 jspl3_w_n1556_37(.douta(w_n1556_37[0]),.doutb(w_n1556_37[1]),.doutc(w_n1556_37[2]),.din(w_n1556_12[0]));
	jspl3 jspl3_w_n1556_38(.douta(w_n1556_38[0]),.doutb(w_n1556_38[1]),.doutc(w_n1556_38[2]),.din(w_n1556_12[1]));
	jspl3 jspl3_w_n1556_39(.douta(w_n1556_39[0]),.doutb(w_n1556_39[1]),.doutc(w_n1556_39[2]),.din(w_n1556_12[2]));
	jspl3 jspl3_w_n1556_40(.douta(w_n1556_40[0]),.doutb(w_n1556_40[1]),.doutc(w_n1556_40[2]),.din(w_n1556_13[0]));
	jspl3 jspl3_w_n1556_41(.douta(w_n1556_41[0]),.doutb(w_n1556_41[1]),.doutc(w_n1556_41[2]),.din(w_n1556_13[1]));
	jspl3 jspl3_w_n1556_42(.douta(w_n1556_42[0]),.doutb(w_n1556_42[1]),.doutc(w_n1556_42[2]),.din(w_n1556_13[2]));
	jspl3 jspl3_w_n1556_43(.douta(w_n1556_43[0]),.doutb(w_n1556_43[1]),.doutc(w_n1556_43[2]),.din(w_n1556_14[0]));
	jspl3 jspl3_w_n1556_44(.douta(w_n1556_44[0]),.doutb(w_n1556_44[1]),.doutc(w_n1556_44[2]),.din(w_n1556_14[1]));
	jspl3 jspl3_w_n1556_45(.douta(w_n1556_45[0]),.doutb(w_n1556_45[1]),.doutc(w_n1556_45[2]),.din(w_n1556_14[2]));
	jspl3 jspl3_w_n1556_46(.douta(w_n1556_46[0]),.doutb(w_n1556_46[1]),.doutc(w_n1556_46[2]),.din(w_n1556_15[0]));
	jspl3 jspl3_w_n1556_47(.douta(w_n1556_47[0]),.doutb(w_n1556_47[1]),.doutc(w_n1556_47[2]),.din(w_n1556_15[1]));
	jspl3 jspl3_w_n1556_48(.douta(w_n1556_48[0]),.doutb(w_n1556_48[1]),.doutc(w_n1556_48[2]),.din(w_n1556_15[2]));
	jspl3 jspl3_w_n1556_49(.douta(w_n1556_49[0]),.doutb(w_n1556_49[1]),.doutc(w_n1556_49[2]),.din(w_n1556_16[0]));
	jspl3 jspl3_w_n1556_50(.douta(w_n1556_50[0]),.doutb(w_n1556_50[1]),.doutc(w_n1556_50[2]),.din(w_n1556_16[1]));
	jspl3 jspl3_w_n1556_51(.douta(w_n1556_51[0]),.doutb(w_n1556_51[1]),.doutc(w_n1556_51[2]),.din(w_n1556_16[2]));
	jspl3 jspl3_w_n1556_52(.douta(w_n1556_52[0]),.doutb(w_n1556_52[1]),.doutc(w_n1556_52[2]),.din(w_n1556_17[0]));
	jspl3 jspl3_w_n1556_53(.douta(w_n1556_53[0]),.doutb(w_n1556_53[1]),.doutc(w_n1556_53[2]),.din(w_n1556_17[1]));
	jspl3 jspl3_w_n1556_54(.douta(w_n1556_54[0]),.doutb(w_n1556_54[1]),.doutc(w_n1556_54[2]),.din(w_n1556_17[2]));
	jspl3 jspl3_w_n1556_55(.douta(w_n1556_55[0]),.doutb(w_n1556_55[1]),.doutc(w_n1556_55[2]),.din(w_n1556_18[0]));
	jspl3 jspl3_w_n1556_56(.douta(w_n1556_56[0]),.doutb(w_n1556_56[1]),.doutc(w_n1556_56[2]),.din(w_n1556_18[1]));
	jspl3 jspl3_w_n1556_57(.douta(w_n1556_57[0]),.doutb(w_n1556_57[1]),.doutc(w_n1556_57[2]),.din(w_n1556_18[2]));
	jspl3 jspl3_w_n1556_58(.douta(w_n1556_58[0]),.doutb(w_n1556_58[1]),.doutc(w_n1556_58[2]),.din(w_n1556_19[0]));
	jspl3 jspl3_w_n1556_59(.douta(w_n1556_59[0]),.doutb(w_n1556_59[1]),.doutc(w_n1556_59[2]),.din(w_n1556_19[1]));
	jspl3 jspl3_w_n1556_60(.douta(w_n1556_60[0]),.doutb(w_n1556_60[1]),.doutc(w_n1556_60[2]),.din(w_n1556_19[2]));
	jspl3 jspl3_w_n1556_61(.douta(w_n1556_61[0]),.doutb(w_n1556_61[1]),.doutc(w_n1556_61[2]),.din(w_n1556_20[0]));
	jspl3 jspl3_w_n1556_62(.douta(w_n1556_62[0]),.doutb(w_n1556_62[1]),.doutc(w_n1556_62[2]),.din(w_n1556_20[1]));
	jspl3 jspl3_w_n1556_63(.douta(w_n1556_63[0]),.doutb(w_n1556_63[1]),.doutc(w_n1556_63[2]),.din(w_n1556_20[2]));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(n1586));
	jspl jspl_w_n1589_0(.douta(w_n1589_0[0]),.doutb(w_n1589_0[1]),.din(n1589));
	jspl3 jspl3_w_n1711_0(.douta(w_n1711_0[0]),.doutb(w_n1711_0[1]),.doutc(w_n1711_0[2]),.din(n1711));
	jspl3 jspl3_w_n1711_1(.douta(w_n1711_1[0]),.doutb(w_n1711_1[1]),.doutc(w_n1711_1[2]),.din(w_n1711_0[0]));
	jspl3 jspl3_w_n1711_2(.douta(w_n1711_2[0]),.doutb(w_n1711_2[1]),.doutc(w_n1711_2[2]),.din(w_n1711_0[1]));
	jspl3 jspl3_w_n1711_3(.douta(w_n1711_3[0]),.doutb(w_n1711_3[1]),.doutc(w_n1711_3[2]),.din(w_n1711_0[2]));
	jspl3 jspl3_w_n1711_4(.douta(w_n1711_4[0]),.doutb(w_n1711_4[1]),.doutc(w_n1711_4[2]),.din(w_n1711_1[0]));
	jspl3 jspl3_w_n1711_5(.douta(w_n1711_5[0]),.doutb(w_n1711_5[1]),.doutc(w_n1711_5[2]),.din(w_n1711_1[1]));
	jspl3 jspl3_w_n1711_6(.douta(w_n1711_6[0]),.doutb(w_n1711_6[1]),.doutc(w_n1711_6[2]),.din(w_n1711_1[2]));
	jspl3 jspl3_w_n1711_7(.douta(w_n1711_7[0]),.doutb(w_n1711_7[1]),.doutc(w_n1711_7[2]),.din(w_n1711_2[0]));
	jspl3 jspl3_w_n1711_8(.douta(w_n1711_8[0]),.doutb(w_n1711_8[1]),.doutc(w_n1711_8[2]),.din(w_n1711_2[1]));
	jspl3 jspl3_w_n1711_9(.douta(w_n1711_9[0]),.doutb(w_n1711_9[1]),.doutc(w_n1711_9[2]),.din(w_n1711_2[2]));
	jspl3 jspl3_w_n1711_10(.douta(w_n1711_10[0]),.doutb(w_n1711_10[1]),.doutc(w_n1711_10[2]),.din(w_n1711_3[0]));
	jspl3 jspl3_w_n1711_11(.douta(w_n1711_11[0]),.doutb(w_n1711_11[1]),.doutc(w_n1711_11[2]),.din(w_n1711_3[1]));
	jspl3 jspl3_w_n1711_12(.douta(w_n1711_12[0]),.doutb(w_n1711_12[1]),.doutc(w_n1711_12[2]),.din(w_n1711_3[2]));
	jspl3 jspl3_w_n1711_13(.douta(w_n1711_13[0]),.doutb(w_n1711_13[1]),.doutc(w_n1711_13[2]),.din(w_n1711_4[0]));
	jspl3 jspl3_w_n1711_14(.douta(w_n1711_14[0]),.doutb(w_n1711_14[1]),.doutc(w_n1711_14[2]),.din(w_n1711_4[1]));
	jspl3 jspl3_w_n1711_15(.douta(w_n1711_15[0]),.doutb(w_n1711_15[1]),.doutc(w_n1711_15[2]),.din(w_n1711_4[2]));
	jspl3 jspl3_w_n1711_16(.douta(w_n1711_16[0]),.doutb(w_n1711_16[1]),.doutc(w_n1711_16[2]),.din(w_n1711_5[0]));
	jspl3 jspl3_w_n1711_17(.douta(w_n1711_17[0]),.doutb(w_n1711_17[1]),.doutc(w_n1711_17[2]),.din(w_n1711_5[1]));
	jspl3 jspl3_w_n1711_18(.douta(w_n1711_18[0]),.doutb(w_n1711_18[1]),.doutc(w_n1711_18[2]),.din(w_n1711_5[2]));
	jspl3 jspl3_w_n1711_19(.douta(w_n1711_19[0]),.doutb(w_n1711_19[1]),.doutc(w_n1711_19[2]),.din(w_n1711_6[0]));
	jspl3 jspl3_w_n1711_20(.douta(w_n1711_20[0]),.doutb(w_n1711_20[1]),.doutc(w_n1711_20[2]),.din(w_n1711_6[1]));
	jspl3 jspl3_w_n1711_21(.douta(w_n1711_21[0]),.doutb(w_n1711_21[1]),.doutc(w_n1711_21[2]),.din(w_n1711_6[2]));
	jspl3 jspl3_w_n1711_22(.douta(w_n1711_22[0]),.doutb(w_n1711_22[1]),.doutc(w_n1711_22[2]),.din(w_n1711_7[0]));
	jspl3 jspl3_w_n1711_23(.douta(w_n1711_23[0]),.doutb(w_n1711_23[1]),.doutc(w_n1711_23[2]),.din(w_n1711_7[1]));
	jspl3 jspl3_w_n1711_24(.douta(w_n1711_24[0]),.doutb(w_n1711_24[1]),.doutc(w_n1711_24[2]),.din(w_n1711_7[2]));
	jspl3 jspl3_w_n1711_25(.douta(w_n1711_25[0]),.doutb(w_n1711_25[1]),.doutc(w_n1711_25[2]),.din(w_n1711_8[0]));
	jspl3 jspl3_w_n1711_26(.douta(w_n1711_26[0]),.doutb(w_n1711_26[1]),.doutc(w_n1711_26[2]),.din(w_n1711_8[1]));
	jspl3 jspl3_w_n1711_27(.douta(w_n1711_27[0]),.doutb(w_n1711_27[1]),.doutc(w_n1711_27[2]),.din(w_n1711_8[2]));
	jspl3 jspl3_w_n1711_28(.douta(w_n1711_28[0]),.doutb(w_n1711_28[1]),.doutc(w_n1711_28[2]),.din(w_n1711_9[0]));
	jspl3 jspl3_w_n1711_29(.douta(w_n1711_29[0]),.doutb(w_n1711_29[1]),.doutc(w_n1711_29[2]),.din(w_n1711_9[1]));
	jspl3 jspl3_w_n1711_30(.douta(w_n1711_30[0]),.doutb(w_n1711_30[1]),.doutc(w_n1711_30[2]),.din(w_n1711_9[2]));
	jspl3 jspl3_w_n1711_31(.douta(w_n1711_31[0]),.doutb(w_n1711_31[1]),.doutc(w_n1711_31[2]),.din(w_n1711_10[0]));
	jspl3 jspl3_w_n1711_32(.douta(w_n1711_32[0]),.doutb(w_n1711_32[1]),.doutc(w_n1711_32[2]),.din(w_n1711_10[1]));
	jspl3 jspl3_w_n1711_33(.douta(w_n1711_33[0]),.doutb(w_n1711_33[1]),.doutc(w_n1711_33[2]),.din(w_n1711_10[2]));
	jspl3 jspl3_w_n1711_34(.douta(w_n1711_34[0]),.doutb(w_n1711_34[1]),.doutc(w_n1711_34[2]),.din(w_n1711_11[0]));
	jspl3 jspl3_w_n1711_35(.douta(w_n1711_35[0]),.doutb(w_n1711_35[1]),.doutc(w_n1711_35[2]),.din(w_n1711_11[1]));
	jspl3 jspl3_w_n1711_36(.douta(w_n1711_36[0]),.doutb(w_n1711_36[1]),.doutc(w_n1711_36[2]),.din(w_n1711_11[2]));
	jspl3 jspl3_w_n1711_37(.douta(w_n1711_37[0]),.doutb(w_n1711_37[1]),.doutc(w_n1711_37[2]),.din(w_n1711_12[0]));
	jspl3 jspl3_w_n1711_38(.douta(w_n1711_38[0]),.doutb(w_n1711_38[1]),.doutc(w_n1711_38[2]),.din(w_n1711_12[1]));
	jspl3 jspl3_w_n1711_39(.douta(w_n1711_39[0]),.doutb(w_n1711_39[1]),.doutc(w_n1711_39[2]),.din(w_n1711_12[2]));
	jspl3 jspl3_w_n1711_40(.douta(w_n1711_40[0]),.doutb(w_n1711_40[1]),.doutc(w_n1711_40[2]),.din(w_n1711_13[0]));
	jspl3 jspl3_w_n1711_41(.douta(w_n1711_41[0]),.doutb(w_n1711_41[1]),.doutc(w_n1711_41[2]),.din(w_n1711_13[1]));
	jspl3 jspl3_w_n1711_42(.douta(w_n1711_42[0]),.doutb(w_n1711_42[1]),.doutc(w_n1711_42[2]),.din(w_n1711_13[2]));
	jspl3 jspl3_w_n1711_43(.douta(w_n1711_43[0]),.doutb(w_n1711_43[1]),.doutc(w_n1711_43[2]),.din(w_n1711_14[0]));
	jspl3 jspl3_w_n1711_44(.douta(w_n1711_44[0]),.doutb(w_n1711_44[1]),.doutc(w_n1711_44[2]),.din(w_n1711_14[1]));
	jspl3 jspl3_w_n1711_45(.douta(w_n1711_45[0]),.doutb(w_n1711_45[1]),.doutc(w_n1711_45[2]),.din(w_n1711_14[2]));
	jspl3 jspl3_w_n1711_46(.douta(w_n1711_46[0]),.doutb(w_n1711_46[1]),.doutc(w_n1711_46[2]),.din(w_n1711_15[0]));
	jspl3 jspl3_w_n1711_47(.douta(w_n1711_47[0]),.doutb(w_n1711_47[1]),.doutc(w_n1711_47[2]),.din(w_n1711_15[1]));
	jspl3 jspl3_w_n1711_48(.douta(w_n1711_48[0]),.doutb(w_n1711_48[1]),.doutc(w_n1711_48[2]),.din(w_n1711_15[2]));
	jspl3 jspl3_w_n1711_49(.douta(w_n1711_49[0]),.doutb(w_n1711_49[1]),.doutc(w_n1711_49[2]),.din(w_n1711_16[0]));
	jspl3 jspl3_w_n1711_50(.douta(w_n1711_50[0]),.doutb(w_n1711_50[1]),.doutc(w_n1711_50[2]),.din(w_n1711_16[1]));
	jspl3 jspl3_w_n1711_51(.douta(w_n1711_51[0]),.doutb(w_n1711_51[1]),.doutc(w_n1711_51[2]),.din(w_n1711_16[2]));
	jspl3 jspl3_w_n1711_52(.douta(w_n1711_52[0]),.doutb(w_n1711_52[1]),.doutc(w_n1711_52[2]),.din(w_n1711_17[0]));
	jspl3 jspl3_w_n1711_53(.douta(w_n1711_53[0]),.doutb(w_n1711_53[1]),.doutc(w_n1711_53[2]),.din(w_n1711_17[1]));
	jspl3 jspl3_w_n1711_54(.douta(w_n1711_54[0]),.doutb(w_n1711_54[1]),.doutc(w_n1711_54[2]),.din(w_n1711_17[2]));
	jspl3 jspl3_w_n1711_55(.douta(w_n1711_55[0]),.doutb(w_n1711_55[1]),.doutc(w_n1711_55[2]),.din(w_n1711_18[0]));
	jspl3 jspl3_w_n1711_56(.douta(w_n1711_56[0]),.doutb(w_n1711_56[1]),.doutc(w_n1711_56[2]),.din(w_n1711_18[1]));
	jspl3 jspl3_w_n1711_57(.douta(w_n1711_57[0]),.doutb(w_n1711_57[1]),.doutc(w_n1711_57[2]),.din(w_n1711_18[2]));
	jspl3 jspl3_w_n1711_58(.douta(w_n1711_58[0]),.doutb(w_n1711_58[1]),.doutc(w_n1711_58[2]),.din(w_n1711_19[0]));
	jspl3 jspl3_w_n1711_59(.douta(w_n1711_59[0]),.doutb(w_n1711_59[1]),.doutc(w_n1711_59[2]),.din(w_n1711_19[1]));
	jspl3 jspl3_w_n1711_60(.douta(w_n1711_60[0]),.doutb(w_n1711_60[1]),.doutc(w_n1711_60[2]),.din(w_n1711_19[2]));
	jspl3 jspl3_w_n1711_61(.douta(w_n1711_61[0]),.doutb(w_n1711_61[1]),.doutc(w_n1711_61[2]),.din(w_n1711_20[0]));
	jspl3 jspl3_w_n1711_62(.douta(w_n1711_62[0]),.doutb(w_n1711_62[1]),.doutc(w_n1711_62[2]),.din(w_n1711_20[1]));
	jspl3 jspl3_w_n1711_63(.douta(w_n1711_63[0]),.doutb(w_n1711_63[1]),.doutc(w_n1711_63[2]),.din(w_n1711_20[2]));
	jspl jspl_w_n1711_64(.douta(w_n1711_64[0]),.doutb(w_n1711_64[1]),.din(w_n1711_21[0]));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl jspl_w_n1715_0(.douta(w_n1715_0[0]),.doutb(w_n1715_0[1]),.din(n1715));
	jspl jspl_w_n1718_0(.douta(w_n1718_0[0]),.doutb(w_n1718_0[1]),.din(n1718));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1723_0(.douta(w_n1723_0[0]),.doutb(w_n1723_0[1]),.din(n1723));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_n1728_0[1]),.din(n1728));
	jspl jspl_w_n1730_0(.douta(w_n1730_0[0]),.doutb(w_n1730_0[1]),.din(n1730));
	jspl jspl_w_n1733_0(.douta(w_n1733_0[0]),.doutb(w_n1733_0[1]),.din(n1733));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(n1735));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(n1738));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(n1740));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(n1743));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(n1745));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl jspl_w_n1753_0(.douta(w_n1753_0[0]),.doutb(w_n1753_0[1]),.din(n1753));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1760_0(.douta(w_n1760_0[0]),.doutb(w_n1760_0[1]),.din(n1760));
	jspl jspl_w_n1763_0(.douta(w_n1763_0[0]),.doutb(w_n1763_0[1]),.din(n1763));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_n1768_0[1]),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(n1770));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(n1773));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(n1775));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(n1778));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1788_0(.douta(w_n1788_0[0]),.doutb(w_n1788_0[1]),.din(n1788));
	jspl jspl_w_n1790_0(.douta(w_n1790_0[0]),.doutb(w_n1790_0[1]),.din(n1790));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1795_0(.douta(w_n1795_0[0]),.doutb(w_n1795_0[1]),.din(n1795));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(n1798));
	jspl jspl_w_n1800_0(.douta(w_n1800_0[0]),.doutb(w_n1800_0[1]),.din(n1800));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_n1805_0[1]),.din(n1805));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(n1808));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1818_0(.douta(w_n1818_0[0]),.doutb(w_n1818_0[1]),.din(n1818));
	jspl jspl_w_n1820_0(.douta(w_n1820_0[0]),.doutb(w_n1820_0[1]),.din(n1820));
	jspl jspl_w_n1823_0(.douta(w_n1823_0[0]),.doutb(w_n1823_0[1]),.din(n1823));
	jspl jspl_w_n1825_0(.douta(w_n1825_0[0]),.doutb(w_n1825_0[1]),.din(n1825));
	jspl jspl_w_n1828_0(.douta(w_n1828_0[0]),.doutb(w_n1828_0[1]),.din(n1828));
	jspl jspl_w_n1830_0(.douta(w_n1830_0[0]),.doutb(w_n1830_0[1]),.din(n1830));
	jspl jspl_w_n1833_0(.douta(w_n1833_0[0]),.doutb(w_n1833_0[1]),.din(n1833));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(n1838));
	jspl jspl_w_n1840_0(.douta(w_n1840_0[0]),.doutb(w_n1840_0[1]),.din(n1840));
	jspl jspl_w_n1843_0(.douta(w_n1843_0[0]),.doutb(w_n1843_0[1]),.din(n1843));
	jspl jspl_w_n1845_0(.douta(w_n1845_0[0]),.doutb(w_n1845_0[1]),.din(n1845));
	jspl jspl_w_n1848_0(.douta(w_n1848_0[0]),.doutb(w_n1848_0[1]),.din(n1848));
	jspl jspl_w_n1850_0(.douta(w_n1850_0[0]),.doutb(w_n1850_0[1]),.din(n1850));
	jspl jspl_w_n1852_0(.douta(w_n1852_0[0]),.doutb(w_n1852_0[1]),.din(n1852));
	jspl jspl_w_n1853_0(.douta(w_n1853_0[0]),.doutb(w_n1853_0[1]),.din(n1853));
	jspl jspl_w_n1854_0(.douta(w_n1854_0[0]),.doutb(w_n1854_0[1]),.din(n1854));
	jspl jspl_w_n1855_0(.douta(w_n1855_0[0]),.doutb(w_n1855_0[1]),.din(n1855));
	jspl3 jspl3_w_n1857_0(.douta(w_n1857_0[0]),.doutb(w_n1857_0[1]),.doutc(w_n1857_0[2]),.din(n1857));
	jspl jspl_w_n1860_0(.douta(w_n1860_0[0]),.doutb(w_n1860_0[1]),.din(n1860));
	jspl jspl_w_n1925_0(.douta(w_n1925_0[0]),.doutb(w_n1925_0[1]),.din(n1925));
	jspl jspl_w_n1930_0(.douta(w_n1930_0[0]),.doutb(w_n1930_0[1]),.din(n1930));
	jspl jspl_w_n1934_0(.douta(w_n1934_0[0]),.doutb(w_n1934_0[1]),.din(n1934));
	jspl jspl_w_n1939_0(.douta(w_n1939_0[0]),.doutb(w_n1939_0[1]),.din(n1939));
	jspl jspl_w_n1943_0(.douta(w_n1943_0[0]),.doutb(w_n1943_0[1]),.din(n1943));
	jspl jspl_w_n1946_0(.douta(w_n1946_0[0]),.doutb(w_n1946_0[1]),.din(n1946));
	jspl jspl_w_n1952_0(.douta(w_n1952_0[0]),.doutb(w_n1952_0[1]),.din(n1952));
	jspl jspl_w_n1987_0(.douta(w_n1987_0[0]),.doutb(w_n1987_0[1]),.din(n1987));
	jspl jspl_w_n1992_0(.douta(w_n1992_0[0]),.doutb(w_n1992_0[1]),.din(n1992));
	jspl jspl_w_n1996_0(.douta(w_n1996_0[0]),.doutb(w_n1996_0[1]),.din(n1996));
	jspl jspl_w_n2001_0(.douta(w_n2001_0[0]),.doutb(w_n2001_0[1]),.din(n2001));
	jspl jspl_w_n2003_0(.douta(w_n2003_0[0]),.doutb(w_n2003_0[1]),.din(n2003));
	jspl jspl_w_n2007_0(.douta(w_n2007_0[0]),.doutb(w_n2007_0[1]),.din(n2007));
	jspl jspl_w_n2011_0(.douta(w_n2011_0[0]),.doutb(w_n2011_0[1]),.din(n2011));
	jspl jspl_w_n2046_0(.douta(w_n2046_0[0]),.doutb(w_n2046_0[1]),.din(n2046));
	jspl jspl_w_n2051_0(.douta(w_n2051_0[0]),.doutb(w_n2051_0[1]),.din(n2051));
	jspl jspl_w_n2052_0(.douta(w_n2052_0[0]),.doutb(w_n2052_0[1]),.din(n2052));
	jspl jspl_w_n2054_0(.douta(w_n2054_0[0]),.doutb(w_n2054_0[1]),.din(n2054));
	jspl jspl_w_n2060_0(.douta(w_n2060_0[0]),.doutb(w_n2060_0[1]),.din(n2060));
	jspl jspl_w_n2065_0(.douta(w_n2065_0[0]),.doutb(w_n2065_0[1]),.din(n2065));
	jspl jspl_w_n2069_0(.douta(w_n2069_0[0]),.doutb(w_n2069_0[1]),.din(n2069));
	jspl jspl_w_n2073_0(.douta(w_n2073_0[0]),.doutb(w_n2073_0[1]),.din(n2073));
	jspl jspl_w_n2104_0(.douta(w_n2104_0[0]),.doutb(w_n2104_0[1]),.din(n2104));
	jspl jspl_w_n2109_0(.douta(w_n2109_0[0]),.doutb(w_n2109_0[1]),.din(n2109));
	jspl jspl_w_n2113_0(.douta(w_n2113_0[0]),.doutb(w_n2113_0[1]),.din(n2113));
	jspl jspl_w_n2118_0(.douta(w_n2118_0[0]),.doutb(w_n2118_0[1]),.din(n2118));
	jspl jspl_w_n2120_0(.douta(w_n2120_0[0]),.doutb(w_n2120_0[1]),.din(n2120));
	jspl jspl_w_n2124_0(.douta(w_n2124_0[0]),.doutb(w_n2124_0[1]),.din(n2124));
	jspl jspl_w_n2128_0(.douta(w_n2128_0[0]),.doutb(w_n2128_0[1]),.din(n2128));
	jspl jspl_w_n2163_0(.douta(w_n2163_0[0]),.doutb(w_n2163_0[1]),.din(n2163));
	jspl jspl_w_n2169_0(.douta(w_n2169_0[0]),.doutb(w_n2169_0[1]),.din(n2169));
	jspl jspl_w_n2171_0(.douta(w_n2171_0[0]),.doutb(w_n2171_0[1]),.din(n2171));
	jspl jspl_w_n2175_0(.douta(w_n2175_0[0]),.doutb(w_n2175_0[1]),.din(n2175));
	jspl jspl_w_n2192_0(.douta(w_n2192_0[0]),.doutb(w_n2192_0[1]),.din(n2192));
	jspl jspl_w_n2199_0(.douta(w_n2199_0[0]),.doutb(w_n2199_0[1]),.din(n2199));
	jspl jspl_w_n2203_0(.douta(w_n2203_0[0]),.doutb(w_n2203_0[1]),.din(n2203));
	jspl jspl_w_n2204_0(.douta(w_n2204_0[0]),.doutb(w_n2204_0[1]),.din(n2204));
	jspl jspl_w_n2221_0(.douta(w_n2221_0[0]),.doutb(w_n2221_0[1]),.din(n2221));
	jspl jspl_w_n2227_0(.douta(w_n2227_0[0]),.doutb(w_n2227_0[1]),.din(n2227));
	jspl jspl_w_n2229_0(.douta(w_n2229_0[0]),.doutb(w_n2229_0[1]),.din(n2229));
	jspl jspl_w_n2233_0(.douta(w_n2233_0[0]),.doutb(w_n2233_0[1]),.din(n2233));
	jspl jspl_w_n2250_0(.douta(w_n2250_0[0]),.doutb(w_n2250_0[1]),.din(n2250));
	jspl jspl_w_n2257_0(.douta(w_n2257_0[0]),.doutb(w_n2257_0[1]),.din(n2257));
	jspl jspl_w_n2261_0(.douta(w_n2261_0[0]),.doutb(w_n2261_0[1]),.din(n2261));
	jspl jspl_w_n2262_0(.douta(w_n2262_0[0]),.doutb(w_n2262_0[1]),.din(n2262));
	jspl jspl_w_n2279_0(.douta(w_n2279_0[0]),.doutb(w_n2279_0[1]),.din(n2279));
	jspl jspl_w_n2285_0(.douta(w_n2285_0[0]),.doutb(w_n2285_0[1]),.din(n2285));
	jspl jspl_w_n2287_0(.douta(w_n2287_0[0]),.doutb(w_n2287_0[1]),.din(n2287));
	jspl jspl_w_n2291_0(.douta(w_n2291_0[0]),.doutb(w_n2291_0[1]),.din(n2291));
	jspl jspl_w_n2308_0(.douta(w_n2308_0[0]),.doutb(w_n2308_0[1]),.din(n2308));
	jspl jspl_w_n2315_0(.douta(w_n2315_0[0]),.doutb(w_n2315_0[1]),.din(n2315));
	jspl jspl_w_n2319_0(.douta(w_n2319_0[0]),.doutb(w_n2319_0[1]),.din(n2319));
	jspl jspl_w_n2320_0(.douta(w_n2320_0[0]),.doutb(w_n2320_0[1]),.din(n2320));
	jspl jspl_w_n2337_0(.douta(w_n2337_0[0]),.doutb(w_n2337_0[1]),.din(n2337));
	jspl jspl_w_n2343_0(.douta(w_n2343_0[0]),.doutb(w_n2343_0[1]),.din(n2343));
	jspl jspl_w_n2345_0(.douta(w_n2345_0[0]),.doutb(w_n2345_0[1]),.din(n2345));
	jspl jspl_w_n2349_0(.douta(w_n2349_0[0]),.doutb(w_n2349_0[1]),.din(n2349));
	jspl jspl_w_n2366_0(.douta(w_n2366_0[0]),.doutb(w_n2366_0[1]),.din(n2366));
	jspl jspl_w_n2373_0(.douta(w_n2373_0[0]),.doutb(w_n2373_0[1]),.din(n2373));
	jspl jspl_w_n2377_0(.douta(w_n2377_0[0]),.doutb(w_n2377_0[1]),.din(n2377));
	jspl jspl_w_n2378_0(.douta(w_n2378_0[0]),.doutb(w_n2378_0[1]),.din(n2378));
	jspl jspl_w_n2395_0(.douta(w_n2395_0[0]),.doutb(w_n2395_0[1]),.din(n2395));
	jspl jspl_w_n2401_0(.douta(w_n2401_0[0]),.doutb(w_n2401_0[1]),.din(n2401));
	jspl jspl_w_n2403_0(.douta(w_n2403_0[0]),.doutb(w_n2403_0[1]),.din(n2403));
	jspl jspl_w_n2407_0(.douta(w_n2407_0[0]),.doutb(w_n2407_0[1]),.din(n2407));
	jspl jspl_w_n2424_0(.douta(w_n2424_0[0]),.doutb(w_n2424_0[1]),.din(n2424));
	jspl jspl_w_n2431_0(.douta(w_n2431_0[0]),.doutb(w_n2431_0[1]),.din(n2431));
	jspl jspl_w_n2435_0(.douta(w_n2435_0[0]),.doutb(w_n2435_0[1]),.din(n2435));
	jspl jspl_w_n2436_0(.douta(w_n2436_0[0]),.doutb(w_n2436_0[1]),.din(n2436));
	jspl jspl_w_n2453_0(.douta(w_n2453_0[0]),.doutb(w_n2453_0[1]),.din(n2453));
	jspl jspl_w_n2459_0(.douta(w_n2459_0[0]),.doutb(w_n2459_0[1]),.din(n2459));
	jspl jspl_w_n2461_0(.douta(w_n2461_0[0]),.doutb(w_n2461_0[1]),.din(n2461));
	jspl jspl_w_n2465_0(.douta(w_n2465_0[0]),.doutb(w_n2465_0[1]),.din(n2465));
	jspl jspl_w_n2482_0(.douta(w_n2482_0[0]),.doutb(w_n2482_0[1]),.din(n2482));
	jspl jspl_w_n2489_0(.douta(w_n2489_0[0]),.doutb(w_n2489_0[1]),.din(n2489));
	jspl jspl_w_n2493_0(.douta(w_n2493_0[0]),.doutb(w_n2493_0[1]),.din(n2493));
	jspl jspl_w_n2494_0(.douta(w_n2494_0[0]),.doutb(w_n2494_0[1]),.din(n2494));
	jspl jspl_w_n2511_0(.douta(w_n2511_0[0]),.doutb(w_n2511_0[1]),.din(n2511));
	jspl jspl_w_n2517_0(.douta(w_n2517_0[0]),.doutb(w_n2517_0[1]),.din(n2517));
	jspl jspl_w_n2519_0(.douta(w_n2519_0[0]),.doutb(w_n2519_0[1]),.din(n2519));
	jspl jspl_w_n2523_0(.douta(w_n2523_0[0]),.doutb(w_n2523_0[1]),.din(n2523));
	jspl jspl_w_n2540_0(.douta(w_n2540_0[0]),.doutb(w_n2540_0[1]),.din(n2540));
	jspl jspl_w_n2547_0(.douta(w_n2547_0[0]),.doutb(w_n2547_0[1]),.din(n2547));
	jspl jspl_w_n2551_0(.douta(w_n2551_0[0]),.doutb(w_n2551_0[1]),.din(n2551));
	jspl jspl_w_n2552_0(.douta(w_n2552_0[0]),.doutb(w_n2552_0[1]),.din(n2552));
	jspl jspl_w_n2569_0(.douta(w_n2569_0[0]),.doutb(w_n2569_0[1]),.din(n2569));
	jspl jspl_w_n2575_0(.douta(w_n2575_0[0]),.doutb(w_n2575_0[1]),.din(n2575));
	jspl jspl_w_n2577_0(.douta(w_n2577_0[0]),.doutb(w_n2577_0[1]),.din(n2577));
	jspl jspl_w_n2581_0(.douta(w_n2581_0[0]),.doutb(w_n2581_0[1]),.din(n2581));
	jspl jspl_w_n2598_0(.douta(w_n2598_0[0]),.doutb(w_n2598_0[1]),.din(n2598));
	jspl jspl_w_n2604_0(.douta(w_n2604_0[0]),.doutb(w_n2604_0[1]),.din(n2604));
	jspl jspl_w_n2606_0(.douta(w_n2606_0[0]),.doutb(w_n2606_0[1]),.din(n2606));
	jspl jspl_w_n2610_0(.douta(w_n2610_0[0]),.doutb(w_n2610_0[1]),.din(n2610));
	jspl jspl_w_n2627_0(.douta(w_n2627_0[0]),.doutb(w_n2627_0[1]),.din(n2627));
	jspl3 jspl3_w_n2628_0(.douta(w_n2628_0[0]),.doutb(w_n2628_0[1]),.doutc(w_n2628_0[2]),.din(n2628));
	jspl3 jspl3_w_n2628_1(.douta(w_n2628_1[0]),.doutb(w_n2628_1[1]),.doutc(w_n2628_1[2]),.din(w_n2628_0[0]));
	jspl3 jspl3_w_n2628_2(.douta(w_n2628_2[0]),.doutb(w_n2628_2[1]),.doutc(w_n2628_2[2]),.din(w_n2628_0[1]));
	jspl3 jspl3_w_n2628_3(.douta(w_n2628_3[0]),.doutb(w_n2628_3[1]),.doutc(w_n2628_3[2]),.din(w_n2628_0[2]));
	jspl3 jspl3_w_n2628_4(.douta(w_n2628_4[0]),.doutb(w_n2628_4[1]),.doutc(w_n2628_4[2]),.din(w_n2628_1[0]));
	jspl3 jspl3_w_n2628_5(.douta(w_n2628_5[0]),.doutb(w_n2628_5[1]),.doutc(w_n2628_5[2]),.din(w_n2628_1[1]));
	jspl3 jspl3_w_n2628_6(.douta(w_n2628_6[0]),.doutb(w_n2628_6[1]),.doutc(w_n2628_6[2]),.din(w_n2628_1[2]));
	jspl3 jspl3_w_n2628_7(.douta(w_n2628_7[0]),.doutb(w_n2628_7[1]),.doutc(w_n2628_7[2]),.din(w_n2628_2[0]));
	jspl3 jspl3_w_n2628_8(.douta(w_n2628_8[0]),.doutb(w_n2628_8[1]),.doutc(w_n2628_8[2]),.din(w_n2628_2[1]));
	jspl3 jspl3_w_n2628_9(.douta(w_n2628_9[0]),.doutb(w_n2628_9[1]),.doutc(w_n2628_9[2]),.din(w_n2628_2[2]));
	jspl3 jspl3_w_n2628_10(.douta(w_n2628_10[0]),.doutb(w_n2628_10[1]),.doutc(w_n2628_10[2]),.din(w_n2628_3[0]));
	jspl3 jspl3_w_n2628_11(.douta(w_n2628_11[0]),.doutb(w_n2628_11[1]),.doutc(w_n2628_11[2]),.din(w_n2628_3[1]));
	jspl3 jspl3_w_n2628_12(.douta(w_n2628_12[0]),.doutb(w_n2628_12[1]),.doutc(w_n2628_12[2]),.din(w_n2628_3[2]));
	jspl3 jspl3_w_n2628_13(.douta(w_n2628_13[0]),.doutb(w_n2628_13[1]),.doutc(w_n2628_13[2]),.din(w_n2628_4[0]));
	jspl3 jspl3_w_n2628_14(.douta(w_n2628_14[0]),.doutb(w_n2628_14[1]),.doutc(w_n2628_14[2]),.din(w_n2628_4[1]));
	jspl3 jspl3_w_n2628_15(.douta(w_n2628_15[0]),.doutb(w_n2628_15[1]),.doutc(w_n2628_15[2]),.din(w_n2628_4[2]));
	jspl3 jspl3_w_n2628_16(.douta(w_n2628_16[0]),.doutb(w_n2628_16[1]),.doutc(w_n2628_16[2]),.din(w_n2628_5[0]));
	jspl3 jspl3_w_n2628_17(.douta(w_n2628_17[0]),.doutb(w_n2628_17[1]),.doutc(w_n2628_17[2]),.din(w_n2628_5[1]));
	jspl3 jspl3_w_n2628_18(.douta(w_n2628_18[0]),.doutb(w_n2628_18[1]),.doutc(w_n2628_18[2]),.din(w_n2628_5[2]));
	jspl3 jspl3_w_n2628_19(.douta(w_n2628_19[0]),.doutb(w_n2628_19[1]),.doutc(w_n2628_19[2]),.din(w_n2628_6[0]));
	jspl3 jspl3_w_n2628_20(.douta(w_n2628_20[0]),.doutb(w_n2628_20[1]),.doutc(w_n2628_20[2]),.din(w_n2628_6[1]));
	jspl3 jspl3_w_n2628_21(.douta(w_n2628_21[0]),.doutb(w_n2628_21[1]),.doutc(w_n2628_21[2]),.din(w_n2628_6[2]));
	jspl3 jspl3_w_n2628_22(.douta(w_n2628_22[0]),.doutb(w_n2628_22[1]),.doutc(w_n2628_22[2]),.din(w_n2628_7[0]));
	jspl3 jspl3_w_n2628_23(.douta(w_n2628_23[0]),.doutb(w_n2628_23[1]),.doutc(w_n2628_23[2]),.din(w_n2628_7[1]));
	jspl3 jspl3_w_n2628_24(.douta(w_n2628_24[0]),.doutb(w_n2628_24[1]),.doutc(w_n2628_24[2]),.din(w_n2628_7[2]));
	jspl3 jspl3_w_n2628_25(.douta(w_n2628_25[0]),.doutb(w_n2628_25[1]),.doutc(w_n2628_25[2]),.din(w_n2628_8[0]));
	jspl3 jspl3_w_n2628_26(.douta(w_n2628_26[0]),.doutb(w_n2628_26[1]),.doutc(w_n2628_26[2]),.din(w_n2628_8[1]));
	jspl3 jspl3_w_n2628_27(.douta(w_n2628_27[0]),.doutb(w_n2628_27[1]),.doutc(w_n2628_27[2]),.din(w_n2628_8[2]));
	jspl3 jspl3_w_n2628_28(.douta(w_n2628_28[0]),.doutb(w_n2628_28[1]),.doutc(w_n2628_28[2]),.din(w_n2628_9[0]));
	jspl3 jspl3_w_n2628_29(.douta(w_n2628_29[0]),.doutb(w_n2628_29[1]),.doutc(w_n2628_29[2]),.din(w_n2628_9[1]));
	jspl3 jspl3_w_n2628_30(.douta(w_n2628_30[0]),.doutb(w_n2628_30[1]),.doutc(w_n2628_30[2]),.din(w_n2628_9[2]));
	jspl3 jspl3_w_n2628_31(.douta(w_n2628_31[0]),.doutb(w_n2628_31[1]),.doutc(w_n2628_31[2]),.din(w_n2628_10[0]));
	jspl3 jspl3_w_n2628_32(.douta(w_n2628_32[0]),.doutb(w_n2628_32[1]),.doutc(w_n2628_32[2]),.din(w_n2628_10[1]));
	jspl3 jspl3_w_n2628_33(.douta(w_n2628_33[0]),.doutb(w_n2628_33[1]),.doutc(w_n2628_33[2]),.din(w_n2628_10[2]));
	jspl3 jspl3_w_n2628_34(.douta(w_n2628_34[0]),.doutb(w_n2628_34[1]),.doutc(w_n2628_34[2]),.din(w_n2628_11[0]));
	jspl3 jspl3_w_n2628_35(.douta(w_n2628_35[0]),.doutb(w_n2628_35[1]),.doutc(w_n2628_35[2]),.din(w_n2628_11[1]));
	jspl3 jspl3_w_n2628_36(.douta(w_n2628_36[0]),.doutb(w_n2628_36[1]),.doutc(w_n2628_36[2]),.din(w_n2628_11[2]));
	jspl3 jspl3_w_n2628_37(.douta(w_n2628_37[0]),.doutb(w_n2628_37[1]),.doutc(w_n2628_37[2]),.din(w_n2628_12[0]));
	jspl3 jspl3_w_n2628_38(.douta(w_n2628_38[0]),.doutb(w_n2628_38[1]),.doutc(w_n2628_38[2]),.din(w_n2628_12[1]));
	jspl3 jspl3_w_n2628_39(.douta(w_n2628_39[0]),.doutb(w_n2628_39[1]),.doutc(w_n2628_39[2]),.din(w_n2628_12[2]));
	jspl3 jspl3_w_n2628_40(.douta(w_n2628_40[0]),.doutb(w_n2628_40[1]),.doutc(w_n2628_40[2]),.din(w_n2628_13[0]));
	jspl3 jspl3_w_n2628_41(.douta(w_n2628_41[0]),.doutb(w_n2628_41[1]),.doutc(w_n2628_41[2]),.din(w_n2628_13[1]));
	jspl3 jspl3_w_n2628_42(.douta(w_n2628_42[0]),.doutb(w_n2628_42[1]),.doutc(w_n2628_42[2]),.din(w_n2628_13[2]));
	jspl3 jspl3_w_n2628_43(.douta(w_n2628_43[0]),.doutb(w_n2628_43[1]),.doutc(w_n2628_43[2]),.din(w_n2628_14[0]));
	jspl3 jspl3_w_n2628_44(.douta(w_n2628_44[0]),.doutb(w_n2628_44[1]),.doutc(w_n2628_44[2]),.din(w_n2628_14[1]));
	jspl3 jspl3_w_n2628_45(.douta(w_n2628_45[0]),.doutb(w_n2628_45[1]),.doutc(w_n2628_45[2]),.din(w_n2628_14[2]));
	jspl3 jspl3_w_n2628_46(.douta(w_n2628_46[0]),.doutb(w_n2628_46[1]),.doutc(w_n2628_46[2]),.din(w_n2628_15[0]));
	jspl3 jspl3_w_n2628_47(.douta(w_n2628_47[0]),.doutb(w_n2628_47[1]),.doutc(w_n2628_47[2]),.din(w_n2628_15[1]));
	jspl3 jspl3_w_n2628_48(.douta(w_n2628_48[0]),.doutb(w_n2628_48[1]),.doutc(w_n2628_48[2]),.din(w_n2628_15[2]));
	jspl3 jspl3_w_n2628_49(.douta(w_n2628_49[0]),.doutb(w_n2628_49[1]),.doutc(w_n2628_49[2]),.din(w_n2628_16[0]));
	jspl3 jspl3_w_n2628_50(.douta(w_n2628_50[0]),.doutb(w_n2628_50[1]),.doutc(w_n2628_50[2]),.din(w_n2628_16[1]));
	jspl3 jspl3_w_n2628_51(.douta(w_n2628_51[0]),.doutb(w_n2628_51[1]),.doutc(w_n2628_51[2]),.din(w_n2628_16[2]));
	jspl3 jspl3_w_n2628_52(.douta(w_n2628_52[0]),.doutb(w_n2628_52[1]),.doutc(w_n2628_52[2]),.din(w_n2628_17[0]));
	jspl3 jspl3_w_n2628_53(.douta(w_n2628_53[0]),.doutb(w_n2628_53[1]),.doutc(w_n2628_53[2]),.din(w_n2628_17[1]));
	jspl3 jspl3_w_n2628_54(.douta(w_n2628_54[0]),.doutb(w_n2628_54[1]),.doutc(w_n2628_54[2]),.din(w_n2628_17[2]));
	jspl3 jspl3_w_n2628_55(.douta(w_n2628_55[0]),.doutb(w_n2628_55[1]),.doutc(w_n2628_55[2]),.din(w_n2628_18[0]));
	jspl3 jspl3_w_n2628_56(.douta(w_n2628_56[0]),.doutb(w_n2628_56[1]),.doutc(w_n2628_56[2]),.din(w_n2628_18[1]));
	jspl3 jspl3_w_n2628_57(.douta(w_n2628_57[0]),.doutb(w_n2628_57[1]),.doutc(w_n2628_57[2]),.din(w_n2628_18[2]));
	jspl3 jspl3_w_n2628_58(.douta(w_n2628_58[0]),.doutb(w_n2628_58[1]),.doutc(w_n2628_58[2]),.din(w_n2628_19[0]));
	jspl3 jspl3_w_n2628_59(.douta(w_n2628_59[0]),.doutb(w_n2628_59[1]),.doutc(w_n2628_59[2]),.din(w_n2628_19[1]));
	jspl3 jspl3_w_n2628_60(.douta(w_n2628_60[0]),.doutb(w_n2628_60[1]),.doutc(w_n2628_60[2]),.din(w_n2628_19[2]));
	jspl3 jspl3_w_n2628_61(.douta(w_n2628_61[0]),.doutb(w_n2628_61[1]),.doutc(w_n2628_61[2]),.din(w_n2628_20[0]));
	jspl3 jspl3_w_n2628_62(.douta(w_n2628_62[0]),.doutb(w_n2628_62[1]),.doutc(w_n2628_62[2]),.din(w_n2628_20[1]));
	jspl3 jspl3_w_n2628_63(.douta(w_n2628_63[0]),.doutb(w_n2628_63[1]),.doutc(w_n2628_63[2]),.din(w_n2628_20[2]));
	jspl jspl_w_n2628_64(.douta(w_n2628_64[0]),.doutb(w_n2628_64[1]),.din(w_n2628_21[0]));
	jspl3 jspl3_w_n2658_0(.douta(w_n2658_0[0]),.doutb(w_n2658_0[1]),.doutc(w_n2658_0[2]),.din(n2658));
	jspl jspl_w_n2661_0(.douta(w_n2661_0[0]),.doutb(w_n2661_0[1]),.din(n2661));
	jspl3 jspl3_w_n2783_0(.douta(w_n2783_0[0]),.doutb(w_n2783_0[1]),.doutc(w_n2783_0[2]),.din(n2783));
	jspl3 jspl3_w_n2783_1(.douta(w_n2783_1[0]),.doutb(w_n2783_1[1]),.doutc(w_n2783_1[2]),.din(w_n2783_0[0]));
	jspl3 jspl3_w_n2783_2(.douta(w_n2783_2[0]),.doutb(w_n2783_2[1]),.doutc(w_n2783_2[2]),.din(w_n2783_0[1]));
	jspl3 jspl3_w_n2783_3(.douta(w_n2783_3[0]),.doutb(w_n2783_3[1]),.doutc(w_n2783_3[2]),.din(w_n2783_0[2]));
	jspl3 jspl3_w_n2783_4(.douta(w_n2783_4[0]),.doutb(w_n2783_4[1]),.doutc(w_n2783_4[2]),.din(w_n2783_1[0]));
	jspl3 jspl3_w_n2783_5(.douta(w_n2783_5[0]),.doutb(w_n2783_5[1]),.doutc(w_n2783_5[2]),.din(w_n2783_1[1]));
	jspl3 jspl3_w_n2783_6(.douta(w_n2783_6[0]),.doutb(w_n2783_6[1]),.doutc(w_n2783_6[2]),.din(w_n2783_1[2]));
	jspl3 jspl3_w_n2783_7(.douta(w_n2783_7[0]),.doutb(w_n2783_7[1]),.doutc(w_n2783_7[2]),.din(w_n2783_2[0]));
	jspl3 jspl3_w_n2783_8(.douta(w_n2783_8[0]),.doutb(w_n2783_8[1]),.doutc(w_n2783_8[2]),.din(w_n2783_2[1]));
	jspl3 jspl3_w_n2783_9(.douta(w_n2783_9[0]),.doutb(w_n2783_9[1]),.doutc(w_n2783_9[2]),.din(w_n2783_2[2]));
	jspl3 jspl3_w_n2783_10(.douta(w_n2783_10[0]),.doutb(w_n2783_10[1]),.doutc(w_n2783_10[2]),.din(w_n2783_3[0]));
	jspl3 jspl3_w_n2783_11(.douta(w_n2783_11[0]),.doutb(w_n2783_11[1]),.doutc(w_n2783_11[2]),.din(w_n2783_3[1]));
	jspl3 jspl3_w_n2783_12(.douta(w_n2783_12[0]),.doutb(w_n2783_12[1]),.doutc(w_n2783_12[2]),.din(w_n2783_3[2]));
	jspl3 jspl3_w_n2783_13(.douta(w_n2783_13[0]),.doutb(w_n2783_13[1]),.doutc(w_n2783_13[2]),.din(w_n2783_4[0]));
	jspl3 jspl3_w_n2783_14(.douta(w_n2783_14[0]),.doutb(w_n2783_14[1]),.doutc(w_n2783_14[2]),.din(w_n2783_4[1]));
	jspl3 jspl3_w_n2783_15(.douta(w_n2783_15[0]),.doutb(w_n2783_15[1]),.doutc(w_n2783_15[2]),.din(w_n2783_4[2]));
	jspl3 jspl3_w_n2783_16(.douta(w_n2783_16[0]),.doutb(w_n2783_16[1]),.doutc(w_n2783_16[2]),.din(w_n2783_5[0]));
	jspl3 jspl3_w_n2783_17(.douta(w_n2783_17[0]),.doutb(w_n2783_17[1]),.doutc(w_n2783_17[2]),.din(w_n2783_5[1]));
	jspl3 jspl3_w_n2783_18(.douta(w_n2783_18[0]),.doutb(w_n2783_18[1]),.doutc(w_n2783_18[2]),.din(w_n2783_5[2]));
	jspl3 jspl3_w_n2783_19(.douta(w_n2783_19[0]),.doutb(w_n2783_19[1]),.doutc(w_n2783_19[2]),.din(w_n2783_6[0]));
	jspl3 jspl3_w_n2783_20(.douta(w_n2783_20[0]),.doutb(w_n2783_20[1]),.doutc(w_n2783_20[2]),.din(w_n2783_6[1]));
	jspl3 jspl3_w_n2783_21(.douta(w_n2783_21[0]),.doutb(w_n2783_21[1]),.doutc(w_n2783_21[2]),.din(w_n2783_6[2]));
	jspl3 jspl3_w_n2783_22(.douta(w_n2783_22[0]),.doutb(w_n2783_22[1]),.doutc(w_n2783_22[2]),.din(w_n2783_7[0]));
	jspl3 jspl3_w_n2783_23(.douta(w_n2783_23[0]),.doutb(w_n2783_23[1]),.doutc(w_n2783_23[2]),.din(w_n2783_7[1]));
	jspl3 jspl3_w_n2783_24(.douta(w_n2783_24[0]),.doutb(w_n2783_24[1]),.doutc(w_n2783_24[2]),.din(w_n2783_7[2]));
	jspl3 jspl3_w_n2783_25(.douta(w_n2783_25[0]),.doutb(w_n2783_25[1]),.doutc(w_n2783_25[2]),.din(w_n2783_8[0]));
	jspl3 jspl3_w_n2783_26(.douta(w_n2783_26[0]),.doutb(w_n2783_26[1]),.doutc(w_n2783_26[2]),.din(w_n2783_8[1]));
	jspl3 jspl3_w_n2783_27(.douta(w_n2783_27[0]),.doutb(w_n2783_27[1]),.doutc(w_n2783_27[2]),.din(w_n2783_8[2]));
	jspl3 jspl3_w_n2783_28(.douta(w_n2783_28[0]),.doutb(w_n2783_28[1]),.doutc(w_n2783_28[2]),.din(w_n2783_9[0]));
	jspl3 jspl3_w_n2783_29(.douta(w_n2783_29[0]),.doutb(w_n2783_29[1]),.doutc(w_n2783_29[2]),.din(w_n2783_9[1]));
	jspl3 jspl3_w_n2783_30(.douta(w_n2783_30[0]),.doutb(w_n2783_30[1]),.doutc(w_n2783_30[2]),.din(w_n2783_9[2]));
	jspl3 jspl3_w_n2783_31(.douta(w_n2783_31[0]),.doutb(w_n2783_31[1]),.doutc(w_n2783_31[2]),.din(w_n2783_10[0]));
	jspl3 jspl3_w_n2783_32(.douta(w_n2783_32[0]),.doutb(w_n2783_32[1]),.doutc(w_n2783_32[2]),.din(w_n2783_10[1]));
	jspl3 jspl3_w_n2783_33(.douta(w_n2783_33[0]),.doutb(w_n2783_33[1]),.doutc(w_n2783_33[2]),.din(w_n2783_10[2]));
	jspl3 jspl3_w_n2783_34(.douta(w_n2783_34[0]),.doutb(w_n2783_34[1]),.doutc(w_n2783_34[2]),.din(w_n2783_11[0]));
	jspl3 jspl3_w_n2783_35(.douta(w_n2783_35[0]),.doutb(w_n2783_35[1]),.doutc(w_n2783_35[2]),.din(w_n2783_11[1]));
	jspl3 jspl3_w_n2783_36(.douta(w_n2783_36[0]),.doutb(w_n2783_36[1]),.doutc(w_n2783_36[2]),.din(w_n2783_11[2]));
	jspl3 jspl3_w_n2783_37(.douta(w_n2783_37[0]),.doutb(w_n2783_37[1]),.doutc(w_n2783_37[2]),.din(w_n2783_12[0]));
	jspl3 jspl3_w_n2783_38(.douta(w_n2783_38[0]),.doutb(w_n2783_38[1]),.doutc(w_n2783_38[2]),.din(w_n2783_12[1]));
	jspl3 jspl3_w_n2783_39(.douta(w_n2783_39[0]),.doutb(w_n2783_39[1]),.doutc(w_n2783_39[2]),.din(w_n2783_12[2]));
	jspl3 jspl3_w_n2783_40(.douta(w_n2783_40[0]),.doutb(w_n2783_40[1]),.doutc(w_n2783_40[2]),.din(w_n2783_13[0]));
	jspl3 jspl3_w_n2783_41(.douta(w_n2783_41[0]),.doutb(w_n2783_41[1]),.doutc(w_n2783_41[2]),.din(w_n2783_13[1]));
	jspl3 jspl3_w_n2783_42(.douta(w_n2783_42[0]),.doutb(w_n2783_42[1]),.doutc(w_n2783_42[2]),.din(w_n2783_13[2]));
	jspl3 jspl3_w_n2783_43(.douta(w_n2783_43[0]),.doutb(w_n2783_43[1]),.doutc(w_n2783_43[2]),.din(w_n2783_14[0]));
	jspl3 jspl3_w_n2783_44(.douta(w_n2783_44[0]),.doutb(w_n2783_44[1]),.doutc(w_n2783_44[2]),.din(w_n2783_14[1]));
	jspl3 jspl3_w_n2783_45(.douta(w_n2783_45[0]),.doutb(w_n2783_45[1]),.doutc(w_n2783_45[2]),.din(w_n2783_14[2]));
	jspl3 jspl3_w_n2783_46(.douta(w_n2783_46[0]),.doutb(w_n2783_46[1]),.doutc(w_n2783_46[2]),.din(w_n2783_15[0]));
	jspl3 jspl3_w_n2783_47(.douta(w_n2783_47[0]),.doutb(w_n2783_47[1]),.doutc(w_n2783_47[2]),.din(w_n2783_15[1]));
	jspl3 jspl3_w_n2783_48(.douta(w_n2783_48[0]),.doutb(w_n2783_48[1]),.doutc(w_n2783_48[2]),.din(w_n2783_15[2]));
	jspl3 jspl3_w_n2783_49(.douta(w_n2783_49[0]),.doutb(w_n2783_49[1]),.doutc(w_n2783_49[2]),.din(w_n2783_16[0]));
	jspl3 jspl3_w_n2783_50(.douta(w_n2783_50[0]),.doutb(w_n2783_50[1]),.doutc(w_n2783_50[2]),.din(w_n2783_16[1]));
	jspl3 jspl3_w_n2783_51(.douta(w_n2783_51[0]),.doutb(w_n2783_51[1]),.doutc(w_n2783_51[2]),.din(w_n2783_16[2]));
	jspl3 jspl3_w_n2783_52(.douta(w_n2783_52[0]),.doutb(w_n2783_52[1]),.doutc(w_n2783_52[2]),.din(w_n2783_17[0]));
	jspl3 jspl3_w_n2783_53(.douta(w_n2783_53[0]),.doutb(w_n2783_53[1]),.doutc(w_n2783_53[2]),.din(w_n2783_17[1]));
	jspl3 jspl3_w_n2783_54(.douta(w_n2783_54[0]),.doutb(w_n2783_54[1]),.doutc(w_n2783_54[2]),.din(w_n2783_17[2]));
	jspl3 jspl3_w_n2783_55(.douta(w_n2783_55[0]),.doutb(w_n2783_55[1]),.doutc(w_n2783_55[2]),.din(w_n2783_18[0]));
	jspl3 jspl3_w_n2783_56(.douta(w_n2783_56[0]),.doutb(w_n2783_56[1]),.doutc(w_n2783_56[2]),.din(w_n2783_18[1]));
	jspl3 jspl3_w_n2783_57(.douta(w_n2783_57[0]),.doutb(w_n2783_57[1]),.doutc(w_n2783_57[2]),.din(w_n2783_18[2]));
	jspl3 jspl3_w_n2783_58(.douta(w_n2783_58[0]),.doutb(w_n2783_58[1]),.doutc(w_n2783_58[2]),.din(w_n2783_19[0]));
	jspl3 jspl3_w_n2783_59(.douta(w_n2783_59[0]),.doutb(w_n2783_59[1]),.doutc(w_n2783_59[2]),.din(w_n2783_19[1]));
	jspl3 jspl3_w_n2783_60(.douta(w_n2783_60[0]),.doutb(w_n2783_60[1]),.doutc(w_n2783_60[2]),.din(w_n2783_19[2]));
	jspl3 jspl3_w_n2783_61(.douta(w_n2783_61[0]),.doutb(w_n2783_61[1]),.doutc(w_n2783_61[2]),.din(w_n2783_20[0]));
	jspl3 jspl3_w_n2783_62(.douta(w_n2783_62[0]),.doutb(w_n2783_62[1]),.doutc(w_n2783_62[2]),.din(w_n2783_20[1]));
	jspl3 jspl3_w_n2783_63(.douta(w_n2783_63[0]),.doutb(w_n2783_63[1]),.doutc(w_n2783_63[2]),.din(w_n2783_20[2]));
	jspl3 jspl3_w_n2783_64(.douta(w_n2783_64[0]),.doutb(w_n2783_64[1]),.doutc(w_n2783_64[2]),.din(w_n2783_21[0]));
	jspl jspl_w_n2785_0(.douta(w_n2785_0[0]),.doutb(w_n2785_0[1]),.din(n2785));
	jspl jspl_w_n2786_0(.douta(w_n2786_0[0]),.doutb(w_n2786_0[1]),.din(n2786));
	jspl3 jspl3_w_n2789_0(.douta(w_n2789_0[0]),.doutb(w_n2789_0[1]),.doutc(w_n2789_0[2]),.din(n2789));
	jspl jspl_w_n2790_0(.douta(w_n2790_0[0]),.doutb(w_n2790_0[1]),.din(n2790));
	jspl3 jspl3_w_n2793_0(.douta(w_n2793_0[0]),.doutb(w_n2793_0[1]),.doutc(w_n2793_0[2]),.din(n2793));
	jspl jspl_w_n2796_0(.douta(w_n2796_0[0]),.doutb(w_n2796_0[1]),.din(n2796));
	jspl jspl_w_n2797_0(.douta(w_n2797_0[0]),.doutb(w_n2797_0[1]),.din(n2797));
	jspl jspl_w_n2798_0(.douta(w_n2798_0[0]),.doutb(w_n2798_0[1]),.din(n2798));
	jspl jspl_w_n2800_0(.douta(w_n2800_0[0]),.doutb(w_n2800_0[1]),.din(n2800));
	jspl3 jspl3_w_n2804_0(.douta(w_n2804_0[0]),.doutb(w_n2804_0[1]),.doutc(w_n2804_0[2]),.din(n2804));
	jspl jspl_w_n2807_0(.douta(w_n2807_0[0]),.doutb(w_n2807_0[1]),.din(n2807));
	jspl jspl_w_n2808_0(.douta(w_n2808_0[0]),.doutb(w_n2808_0[1]),.din(n2808));
	jspl jspl_w_n2809_0(.douta(w_n2809_0[0]),.doutb(w_n2809_0[1]),.din(n2809));
	jspl jspl_w_n2811_0(.douta(w_n2811_0[0]),.doutb(w_n2811_0[1]),.din(n2811));
	jspl3 jspl3_w_n2815_0(.douta(w_n2815_0[0]),.doutb(w_n2815_0[1]),.doutc(w_n2815_0[2]),.din(n2815));
	jspl jspl_w_n2818_0(.douta(w_n2818_0[0]),.doutb(w_n2818_0[1]),.din(n2818));
	jspl jspl_w_n2819_0(.douta(w_n2819_0[0]),.doutb(w_n2819_0[1]),.din(n2819));
	jspl jspl_w_n2820_0(.douta(w_n2820_0[0]),.doutb(w_n2820_0[1]),.din(n2820));
	jspl jspl_w_n2822_0(.douta(w_n2822_0[0]),.doutb(w_n2822_0[1]),.din(n2822));
	jspl3 jspl3_w_n2826_0(.douta(w_n2826_0[0]),.doutb(w_n2826_0[1]),.doutc(w_n2826_0[2]),.din(n2826));
	jspl jspl_w_n2829_0(.douta(w_n2829_0[0]),.doutb(w_n2829_0[1]),.din(n2829));
	jspl jspl_w_n2830_0(.douta(w_n2830_0[0]),.doutb(w_n2830_0[1]),.din(n2830));
	jspl jspl_w_n2831_0(.douta(w_n2831_0[0]),.doutb(w_n2831_0[1]),.din(n2831));
	jspl jspl_w_n2833_0(.douta(w_n2833_0[0]),.doutb(w_n2833_0[1]),.din(n2833));
	jspl3 jspl3_w_n2837_0(.douta(w_n2837_0[0]),.doutb(w_n2837_0[1]),.doutc(w_n2837_0[2]),.din(n2837));
	jspl jspl_w_n2840_0(.douta(w_n2840_0[0]),.doutb(w_n2840_0[1]),.din(n2840));
	jspl jspl_w_n2841_0(.douta(w_n2841_0[0]),.doutb(w_n2841_0[1]),.din(n2841));
	jspl jspl_w_n2842_0(.douta(w_n2842_0[0]),.doutb(w_n2842_0[1]),.din(n2842));
	jspl jspl_w_n2844_0(.douta(w_n2844_0[0]),.doutb(w_n2844_0[1]),.din(n2844));
	jspl3 jspl3_w_n2848_0(.douta(w_n2848_0[0]),.doutb(w_n2848_0[1]),.doutc(w_n2848_0[2]),.din(n2848));
	jspl jspl_w_n2851_0(.douta(w_n2851_0[0]),.doutb(w_n2851_0[1]),.din(n2851));
	jspl jspl_w_n2852_0(.douta(w_n2852_0[0]),.doutb(w_n2852_0[1]),.din(n2852));
	jspl jspl_w_n2853_0(.douta(w_n2853_0[0]),.doutb(w_n2853_0[1]),.din(n2853));
	jspl jspl_w_n2857_0(.douta(w_n2857_0[0]),.doutb(w_n2857_0[1]),.din(n2857));
	jspl jspl_w_n2858_0(.douta(w_n2858_0[0]),.doutb(w_n2858_0[1]),.din(n2858));
	jspl3 jspl3_w_n2861_0(.douta(w_n2861_0[0]),.doutb(w_n2861_0[1]),.doutc(w_n2861_0[2]),.din(n2861));
	jspl jspl_w_n2862_0(.douta(w_n2862_0[0]),.doutb(w_n2862_0[1]),.din(n2862));
	jspl3 jspl3_w_n2865_0(.douta(w_n2865_0[0]),.doutb(w_n2865_0[1]),.doutc(w_n2865_0[2]),.din(n2865));
	jspl jspl_w_n2868_0(.douta(w_n2868_0[0]),.doutb(w_n2868_0[1]),.din(n2868));
	jspl jspl_w_n2869_0(.douta(w_n2869_0[0]),.doutb(w_n2869_0[1]),.din(n2869));
	jspl jspl_w_n2870_0(.douta(w_n2870_0[0]),.doutb(w_n2870_0[1]),.din(n2870));
	jspl jspl_w_n2872_0(.douta(w_n2872_0[0]),.doutb(w_n2872_0[1]),.din(n2872));
	jspl3 jspl3_w_n2876_0(.douta(w_n2876_0[0]),.doutb(w_n2876_0[1]),.doutc(w_n2876_0[2]),.din(n2876));
	jspl jspl_w_n2879_0(.douta(w_n2879_0[0]),.doutb(w_n2879_0[1]),.din(n2879));
	jspl jspl_w_n2880_0(.douta(w_n2880_0[0]),.doutb(w_n2880_0[1]),.din(n2880));
	jspl jspl_w_n2881_0(.douta(w_n2881_0[0]),.doutb(w_n2881_0[1]),.din(n2881));
	jspl jspl_w_n2883_0(.douta(w_n2883_0[0]),.doutb(w_n2883_0[1]),.din(n2883));
	jspl3 jspl3_w_n2887_0(.douta(w_n2887_0[0]),.doutb(w_n2887_0[1]),.doutc(w_n2887_0[2]),.din(n2887));
	jspl jspl_w_n2890_0(.douta(w_n2890_0[0]),.doutb(w_n2890_0[1]),.din(n2890));
	jspl jspl_w_n2891_0(.douta(w_n2891_0[0]),.doutb(w_n2891_0[1]),.din(n2891));
	jspl jspl_w_n2892_0(.douta(w_n2892_0[0]),.doutb(w_n2892_0[1]),.din(n2892));
	jspl3 jspl3_w_n2896_0(.douta(w_n2896_0[0]),.doutb(w_n2896_0[1]),.doutc(w_n2896_0[2]),.din(n2896));
	jspl3 jspl3_w_n2899_0(.douta(w_n2899_0[0]),.doutb(w_n2899_0[1]),.doutc(w_n2899_0[2]),.din(n2899));
	jspl jspl_w_n2899_1(.douta(w_n2899_1[0]),.doutb(w_n2899_1[1]),.din(w_n2899_0[0]));
	jspl jspl_w_n2900_0(.douta(w_n2900_0[0]),.doutb(w_n2900_0[1]),.din(n2900));
	jspl jspl_w_n2903_0(.douta(w_n2903_0[0]),.doutb(w_n2903_0[1]),.din(n2903));
	jspl jspl_w_n2904_0(.douta(w_n2904_0[0]),.doutb(w_n2904_0[1]),.din(n2904));
	jspl3 jspl3_w_n2907_0(.douta(w_n2907_0[0]),.doutb(w_n2907_0[1]),.doutc(w_n2907_0[2]),.din(n2907));
	jspl jspl_w_n2908_0(.douta(w_n2908_0[0]),.doutb(w_n2908_0[1]),.din(n2908));
	jspl jspl_w_n2909_0(.douta(w_n2909_0[0]),.doutb(w_n2909_0[1]),.din(n2909));
	jspl jspl_w_n2912_0(.douta(w_n2912_0[0]),.doutb(w_n2912_0[1]),.din(n2912));
	jspl jspl_w_n2913_0(.douta(w_n2913_0[0]),.doutb(w_n2913_0[1]),.din(n2913));
	jspl3 jspl3_w_n2916_0(.douta(w_n2916_0[0]),.doutb(w_n2916_0[1]),.doutc(w_n2916_0[2]),.din(n2916));
	jspl jspl_w_n2917_0(.douta(w_n2917_0[0]),.doutb(w_n2917_0[1]),.din(n2917));
	jspl jspl_w_n2920_0(.douta(w_n2920_0[0]),.doutb(w_n2920_0[1]),.din(n2920));
	jspl jspl_w_n2921_0(.douta(w_n2921_0[0]),.doutb(w_n2921_0[1]),.din(n2921));
	jspl3 jspl3_w_n2924_0(.douta(w_n2924_0[0]),.doutb(w_n2924_0[1]),.doutc(w_n2924_0[2]),.din(n2924));
	jspl jspl_w_n2925_0(.douta(w_n2925_0[0]),.doutb(w_n2925_0[1]),.din(n2925));
	jspl3 jspl3_w_n2928_0(.douta(w_n2928_0[0]),.doutb(w_n2928_0[1]),.doutc(w_n2928_0[2]),.din(n2928));
	jspl jspl_w_n2931_0(.douta(w_n2931_0[0]),.doutb(w_n2931_0[1]),.din(n2931));
	jspl jspl_w_n2932_0(.douta(w_n2932_0[0]),.doutb(w_n2932_0[1]),.din(n2932));
	jspl jspl_w_n2933_0(.douta(w_n2933_0[0]),.doutb(w_n2933_0[1]),.din(n2933));
	jspl jspl_w_n2935_0(.douta(w_n2935_0[0]),.doutb(w_n2935_0[1]),.din(n2935));
	jspl3 jspl3_w_n2939_0(.douta(w_n2939_0[0]),.doutb(w_n2939_0[1]),.doutc(w_n2939_0[2]),.din(n2939));
	jspl jspl_w_n2942_0(.douta(w_n2942_0[0]),.doutb(w_n2942_0[1]),.din(n2942));
	jspl jspl_w_n2943_0(.douta(w_n2943_0[0]),.doutb(w_n2943_0[1]),.din(n2943));
	jspl jspl_w_n2944_0(.douta(w_n2944_0[0]),.doutb(w_n2944_0[1]),.din(n2944));
	jspl jspl_w_n2946_0(.douta(w_n2946_0[0]),.doutb(w_n2946_0[1]),.din(n2946));
	jspl3 jspl3_w_n2950_0(.douta(w_n2950_0[0]),.doutb(w_n2950_0[1]),.doutc(w_n2950_0[2]),.din(n2950));
	jspl jspl_w_n2953_0(.douta(w_n2953_0[0]),.doutb(w_n2953_0[1]),.din(n2953));
	jspl jspl_w_n2954_0(.douta(w_n2954_0[0]),.doutb(w_n2954_0[1]),.din(n2954));
	jspl jspl_w_n2955_0(.douta(w_n2955_0[0]),.doutb(w_n2955_0[1]),.din(n2955));
	jspl jspl_w_n2957_0(.douta(w_n2957_0[0]),.doutb(w_n2957_0[1]),.din(n2957));
	jspl3 jspl3_w_n2961_0(.douta(w_n2961_0[0]),.doutb(w_n2961_0[1]),.doutc(w_n2961_0[2]),.din(n2961));
	jspl jspl_w_n2964_0(.douta(w_n2964_0[0]),.doutb(w_n2964_0[1]),.din(n2964));
	jspl jspl_w_n2965_0(.douta(w_n2965_0[0]),.doutb(w_n2965_0[1]),.din(n2965));
	jspl jspl_w_n2966_0(.douta(w_n2966_0[0]),.doutb(w_n2966_0[1]),.din(n2966));
	jspl jspl_w_n2968_0(.douta(w_n2968_0[0]),.doutb(w_n2968_0[1]),.din(n2968));
	jspl3 jspl3_w_n2972_0(.douta(w_n2972_0[0]),.doutb(w_n2972_0[1]),.doutc(w_n2972_0[2]),.din(n2972));
	jspl jspl_w_n2975_0(.douta(w_n2975_0[0]),.doutb(w_n2975_0[1]),.din(n2975));
	jspl jspl_w_n2976_0(.douta(w_n2976_0[0]),.doutb(w_n2976_0[1]),.din(n2976));
	jspl jspl_w_n2977_0(.douta(w_n2977_0[0]),.doutb(w_n2977_0[1]),.din(n2977));
	jspl jspl_w_n2979_0(.douta(w_n2979_0[0]),.doutb(w_n2979_0[1]),.din(n2979));
	jspl3 jspl3_w_n2983_0(.douta(w_n2983_0[0]),.doutb(w_n2983_0[1]),.doutc(w_n2983_0[2]),.din(n2983));
	jspl3 jspl3_w_n2986_0(.douta(w_n2986_0[0]),.doutb(w_n2986_0[1]),.doutc(w_n2986_0[2]),.din(n2986));
	jspl jspl_w_n2989_0(.douta(w_n2989_0[0]),.doutb(w_n2989_0[1]),.din(n2989));
	jspl jspl_w_n2990_0(.douta(w_n2990_0[0]),.doutb(w_n2990_0[1]),.din(n2990));
	jspl jspl_w_n2991_0(.douta(w_n2991_0[0]),.doutb(w_n2991_0[1]),.din(n2991));
	jspl jspl_w_n2993_0(.douta(w_n2993_0[0]),.doutb(w_n2993_0[1]),.din(n2993));
	jspl3 jspl3_w_n2997_0(.douta(w_n2997_0[0]),.doutb(w_n2997_0[1]),.doutc(w_n2997_0[2]),.din(n2997));
	jspl3 jspl3_w_n3001_0(.douta(w_n3001_0[0]),.doutb(w_n3001_0[1]),.doutc(w_n3001_0[2]),.din(n3001));
	jspl jspl_w_n3005_0(.douta(w_n3005_0[0]),.doutb(w_n3005_0[1]),.din(n3005));
	jspl jspl_w_n3006_0(.douta(w_n3006_0[0]),.doutb(w_n3006_0[1]),.din(n3006));
	jspl3 jspl3_w_n3009_0(.douta(w_n3009_0[0]),.doutb(w_n3009_0[1]),.doutc(w_n3009_0[2]),.din(n3009));
	jspl jspl_w_n3010_0(.douta(w_n3010_0[0]),.doutb(w_n3010_0[1]),.din(n3010));
	jspl jspl_w_n3011_0(.douta(w_n3011_0[0]),.doutb(w_n3011_0[1]),.din(n3011));
	jspl jspl_w_n3014_0(.douta(w_n3014_0[0]),.doutb(w_n3014_0[1]),.din(n3014));
	jspl3 jspl3_w_n3017_0(.douta(w_n3017_0[0]),.doutb(w_n3017_0[1]),.doutc(w_n3017_0[2]),.din(n3017));
	jspl jspl_w_n3018_0(.douta(w_n3018_0[0]),.doutb(w_n3018_0[1]),.din(n3018));
	jspl3 jspl3_w_n3021_0(.douta(w_n3021_0[0]),.doutb(w_n3021_0[1]),.doutc(w_n3021_0[2]),.din(n3021));
	jspl jspl_w_n3025_0(.douta(w_n3025_0[0]),.doutb(w_n3025_0[1]),.din(n3025));
	jspl jspl_w_n3028_0(.douta(w_n3028_0[0]),.doutb(w_n3028_0[1]),.din(n3028));
	jspl jspl_w_n3037_0(.douta(w_n3037_0[0]),.doutb(w_n3037_0[1]),.din(n3037));
	jspl3 jspl3_w_n3040_0(.douta(w_n3040_0[0]),.doutb(w_n3040_0[1]),.doutc(w_n3040_0[2]),.din(n3040));
	jspl jspl_w_n3040_1(.douta(w_n3040_1[0]),.doutb(w_n3040_1[1]),.din(w_n3040_0[0]));
	jspl jspl_w_n3044_0(.douta(w_n3044_0[0]),.doutb(w_n3044_0[1]),.din(n3044));
	jspl3 jspl3_w_n3047_0(.douta(w_n3047_0[0]),.doutb(w_n3047_0[1]),.doutc(w_n3047_0[2]),.din(n3047));
	jspl jspl_w_n3047_1(.douta(w_n3047_1[0]),.doutb(w_n3047_1[1]),.din(w_n3047_0[0]));
	jspl jspl_w_n3053_0(.douta(w_n3053_0[0]),.doutb(w_n3053_0[1]),.din(n3053));
	jspl jspl_w_n3054_0(.douta(w_n3054_0[0]),.doutb(w_n3054_0[1]),.din(n3054));
	jspl3 jspl3_w_n3057_0(.douta(w_n3057_0[0]),.doutb(w_n3057_0[1]),.doutc(w_n3057_0[2]),.din(n3057));
	jspl jspl_w_n3058_0(.douta(w_n3058_0[0]),.doutb(w_n3058_0[1]),.din(n3058));
	jspl jspl_w_n3061_0(.douta(w_n3061_0[0]),.doutb(w_n3061_0[1]),.din(n3061));
	jspl jspl_w_n3064_0(.douta(w_n3064_0[0]),.doutb(w_n3064_0[1]),.din(n3064));
	jspl3 jspl3_w_n3067_0(.douta(w_n3067_0[0]),.doutb(w_n3067_0[1]),.doutc(w_n3067_0[2]),.din(n3067));
	jspl jspl_w_n3067_1(.douta(w_n3067_1[0]),.doutb(w_n3067_1[1]),.din(w_n3067_0[0]));
	jspl jspl_w_n3068_0(.douta(w_n3068_0[0]),.doutb(w_n3068_0[1]),.din(n3068));
	jspl jspl_w_n3086_0(.douta(w_n3086_0[0]),.doutb(w_n3086_0[1]),.din(n3086));
	jspl jspl_w_n3090_0(.douta(w_n3090_0[0]),.doutb(w_n3090_0[1]),.din(n3090));
	jspl3 jspl3_w_n3095_0(.douta(w_n3095_0[0]),.doutb(w_n3095_0[1]),.doutc(w_n3095_0[2]),.din(n3095));
	jspl jspl_w_n3098_0(.douta(w_n3098_0[0]),.doutb(w_n3098_0[1]),.din(n3098));
	jspl jspl_w_n3099_0(.douta(w_n3099_0[0]),.doutb(w_n3099_0[1]),.din(n3099));
	jspl jspl_w_n3100_0(.douta(w_n3100_0[0]),.doutb(w_n3100_0[1]),.din(n3100));
	jspl jspl_w_n3107_0(.douta(w_n3107_0[0]),.doutb(w_n3107_0[1]),.din(n3107));
	jspl3 jspl3_w_n3119_0(.douta(w_n3119_0[0]),.doutb(w_n3119_0[1]),.doutc(w_n3119_0[2]),.din(n3119));
	jspl jspl_w_n3122_0(.douta(w_n3122_0[0]),.doutb(w_n3122_0[1]),.din(n3122));
	jspl jspl_w_n3123_0(.douta(w_n3123_0[0]),.doutb(w_n3123_0[1]),.din(n3123));
	jspl jspl_w_n3126_0(.douta(w_n3126_0[0]),.doutb(w_n3126_0[1]),.din(n3126));
	jspl jspl_w_n3130_0(.douta(w_n3130_0[0]),.doutb(w_n3130_0[1]),.din(n3130));
	jspl3 jspl3_w_n3148_0(.douta(w_n3148_0[0]),.doutb(w_n3148_0[1]),.doutc(w_n3148_0[2]),.din(n3148));
	jspl jspl_w_n3151_0(.douta(w_n3151_0[0]),.doutb(w_n3151_0[1]),.din(n3151));
	jspl jspl_w_n3152_0(.douta(w_n3152_0[0]),.doutb(w_n3152_0[1]),.din(n3152));
	jspl jspl_w_n3155_0(.douta(w_n3155_0[0]),.doutb(w_n3155_0[1]),.din(n3155));
	jspl jspl_w_n3159_0(.douta(w_n3159_0[0]),.doutb(w_n3159_0[1]),.din(n3159));
	jspl jspl_w_n3160_0(.douta(w_n3160_0[0]),.doutb(w_n3160_0[1]),.din(n3160));
	jspl3 jspl3_w_n3163_0(.douta(w_n3163_0[0]),.doutb(w_n3163_0[1]),.doutc(w_n3163_0[2]),.din(n3163));
	jspl jspl_w_n3167_0(.douta(w_n3167_0[0]),.doutb(w_n3167_0[1]),.din(n3167));
	jspl jspl_w_n3168_0(.douta(w_n3168_0[0]),.doutb(w_n3168_0[1]),.din(n3168));
	jspl3 jspl3_w_n3171_0(.douta(w_n3171_0[0]),.doutb(w_n3171_0[1]),.doutc(w_n3171_0[2]),.din(n3171));
	jspl jspl_w_n3172_0(.douta(w_n3172_0[0]),.doutb(w_n3172_0[1]),.din(n3172));
	jspl3 jspl3_w_n3175_0(.douta(w_n3175_0[0]),.doutb(w_n3175_0[1]),.doutc(w_n3175_0[2]),.din(n3175));
	jspl jspl_w_n3178_0(.douta(w_n3178_0[0]),.doutb(w_n3178_0[1]),.din(n3178));
	jspl jspl_w_n3179_0(.douta(w_n3179_0[0]),.doutb(w_n3179_0[1]),.din(n3179));
	jspl jspl_w_n3182_0(.douta(w_n3182_0[0]),.doutb(w_n3182_0[1]),.din(n3182));
	jspl jspl_w_n3186_0(.douta(w_n3186_0[0]),.doutb(w_n3186_0[1]),.din(n3186));
	jspl jspl_w_n3187_0(.douta(w_n3187_0[0]),.doutb(w_n3187_0[1]),.din(n3187));
	jspl3 jspl3_w_n3190_0(.douta(w_n3190_0[0]),.doutb(w_n3190_0[1]),.doutc(w_n3190_0[2]),.din(n3190));
	jspl jspl_w_n3191_0(.douta(w_n3191_0[0]),.doutb(w_n3191_0[1]),.din(n3191));
	jspl jspl_w_n3194_0(.douta(w_n3194_0[0]),.doutb(w_n3194_0[1]),.din(n3194));
	jspl jspl_w_n3195_0(.douta(w_n3195_0[0]),.doutb(w_n3195_0[1]),.din(n3195));
	jspl3 jspl3_w_n3198_0(.douta(w_n3198_0[0]),.doutb(w_n3198_0[1]),.doutc(w_n3198_0[2]),.din(n3198));
	jspl3 jspl3_w_n3202_0(.douta(w_n3202_0[0]),.doutb(w_n3202_0[1]),.doutc(w_n3202_0[2]),.din(n3202));
	jspl jspl_w_n3205_0(.douta(w_n3205_0[0]),.doutb(w_n3205_0[1]),.din(n3205));
	jspl jspl_w_n3206_0(.douta(w_n3206_0[0]),.doutb(w_n3206_0[1]),.din(n3206));
	jspl jspl_w_n3209_0(.douta(w_n3209_0[0]),.doutb(w_n3209_0[1]),.din(n3209));
	jspl3 jspl3_w_n3213_0(.douta(w_n3213_0[0]),.doutb(w_n3213_0[1]),.doutc(w_n3213_0[2]),.din(n3213));
	jspl jspl_w_n3216_0(.douta(w_n3216_0[0]),.doutb(w_n3216_0[1]),.din(n3216));
	jspl jspl_w_n3217_0(.douta(w_n3217_0[0]),.doutb(w_n3217_0[1]),.din(n3217));
	jspl jspl_w_n3222_0(.douta(w_n3222_0[0]),.doutb(w_n3222_0[1]),.din(n3222));
	jspl jspl_w_n3223_0(.douta(w_n3223_0[0]),.doutb(w_n3223_0[1]),.din(n3223));
	jspl3 jspl3_w_n3226_0(.douta(w_n3226_0[0]),.doutb(w_n3226_0[1]),.doutc(w_n3226_0[2]),.din(n3226));
	jspl jspl_w_n3227_0(.douta(w_n3227_0[0]),.doutb(w_n3227_0[1]),.din(n3227));
	jspl jspl_w_n3233_0(.douta(w_n3233_0[0]),.doutb(w_n3233_0[1]),.din(n3233));
	jspl jspl_w_n3255_0(.douta(w_n3255_0[0]),.doutb(w_n3255_0[1]),.din(n3255));
	jspl jspl_w_n3259_0(.douta(w_n3259_0[0]),.doutb(w_n3259_0[1]),.din(n3259));
	jspl jspl_w_n3260_0(.douta(w_n3260_0[0]),.doutb(w_n3260_0[1]),.din(n3260));
	jspl3 jspl3_w_n3263_0(.douta(w_n3263_0[0]),.doutb(w_n3263_0[1]),.doutc(w_n3263_0[2]),.din(n3263));
	jspl jspl_w_n3267_0(.douta(w_n3267_0[0]),.doutb(w_n3267_0[1]),.din(n3267));
	jspl jspl_w_n3268_0(.douta(w_n3268_0[0]),.doutb(w_n3268_0[1]),.din(n3268));
	jspl3 jspl3_w_n3271_0(.douta(w_n3271_0[0]),.doutb(w_n3271_0[1]),.doutc(w_n3271_0[2]),.din(n3271));
	jspl jspl_w_n3272_0(.douta(w_n3272_0[0]),.doutb(w_n3272_0[1]),.din(n3272));
	jspl3 jspl3_w_n3275_0(.douta(w_n3275_0[0]),.doutb(w_n3275_0[1]),.doutc(w_n3275_0[2]),.din(n3275));
	jspl jspl_w_n3278_0(.douta(w_n3278_0[0]),.doutb(w_n3278_0[1]),.din(n3278));
	jspl jspl_w_n3279_0(.douta(w_n3279_0[0]),.doutb(w_n3279_0[1]),.din(n3279));
	jspl jspl_w_n3282_0(.douta(w_n3282_0[0]),.doutb(w_n3282_0[1]),.din(n3282));
	jspl jspl_w_n3285_0(.douta(w_n3285_0[0]),.doutb(w_n3285_0[1]),.din(n3285));
	jspl jspl_w_n3286_0(.douta(w_n3286_0[0]),.doutb(w_n3286_0[1]),.din(n3286));
	jspl3 jspl3_w_n3289_0(.douta(w_n3289_0[0]),.doutb(w_n3289_0[1]),.doutc(w_n3289_0[2]),.din(n3289));
	jspl jspl_w_n3293_0(.douta(w_n3293_0[0]),.doutb(w_n3293_0[1]),.din(n3293));
	jspl jspl_w_n3294_0(.douta(w_n3294_0[0]),.doutb(w_n3294_0[1]),.din(n3294));
	jspl3 jspl3_w_n3297_0(.douta(w_n3297_0[0]),.doutb(w_n3297_0[1]),.doutc(w_n3297_0[2]),.din(n3297));
	jspl jspl_w_n3299_0(.douta(w_n3299_0[0]),.doutb(w_n3299_0[1]),.din(n3299));
	jspl jspl_w_n3302_0(.douta(w_n3302_0[0]),.doutb(w_n3302_0[1]),.din(n3302));
	jspl jspl_w_n3303_0(.douta(w_n3303_0[0]),.doutb(w_n3303_0[1]),.din(n3303));
	jspl3 jspl3_w_n3306_0(.douta(w_n3306_0[0]),.doutb(w_n3306_0[1]),.doutc(w_n3306_0[2]),.din(n3306));
	jspl jspl_w_n3307_0(.douta(w_n3307_0[0]),.doutb(w_n3307_0[1]),.din(n3307));
	jspl jspl_w_n3310_0(.douta(w_n3310_0[0]),.doutb(w_n3310_0[1]),.din(n3310));
	jspl jspl_w_n3311_0(.douta(w_n3311_0[0]),.doutb(w_n3311_0[1]),.din(n3311));
	jspl3 jspl3_w_n3314_0(.douta(w_n3314_0[0]),.doutb(w_n3314_0[1]),.doutc(w_n3314_0[2]),.din(n3314));
	jspl jspl_w_n3318_0(.douta(w_n3318_0[0]),.doutb(w_n3318_0[1]),.din(n3318));
	jspl jspl_w_n3319_0(.douta(w_n3319_0[0]),.doutb(w_n3319_0[1]),.din(n3319));
	jspl3 jspl3_w_n3322_0(.douta(w_n3322_0[0]),.doutb(w_n3322_0[1]),.doutc(w_n3322_0[2]),.din(n3322));
	jspl jspl_w_n3323_0(.douta(w_n3323_0[0]),.doutb(w_n3323_0[1]),.din(n3323));
	jspl jspl_w_n3327_0(.douta(w_n3327_0[0]),.doutb(w_n3327_0[1]),.din(n3327));
	jspl jspl_w_n3348_0(.douta(w_n3348_0[0]),.doutb(w_n3348_0[1]),.din(n3348));
	jspl jspl_w_n3352_0(.douta(w_n3352_0[0]),.doutb(w_n3352_0[1]),.din(n3352));
	jspl jspl_w_n3353_0(.douta(w_n3353_0[0]),.doutb(w_n3353_0[1]),.din(n3353));
	jspl3 jspl3_w_n3356_0(.douta(w_n3356_0[0]),.doutb(w_n3356_0[1]),.doutc(w_n3356_0[2]),.din(n3356));
	jspl jspl_w_n3357_0(.douta(w_n3357_0[0]),.doutb(w_n3357_0[1]),.din(n3357));
	jspl jspl_w_n3360_0(.douta(w_n3360_0[0]),.doutb(w_n3360_0[1]),.din(n3360));
	jspl jspl_w_n3361_0(.douta(w_n3361_0[0]),.doutb(w_n3361_0[1]),.din(n3361));
	jspl3 jspl3_w_n3364_0(.douta(w_n3364_0[0]),.doutb(w_n3364_0[1]),.doutc(w_n3364_0[2]),.din(n3364));
	jspl3 jspl3_w_n3368_0(.douta(w_n3368_0[0]),.doutb(w_n3368_0[1]),.doutc(w_n3368_0[2]),.din(n3368));
	jspl jspl_w_n3371_0(.douta(w_n3371_0[0]),.doutb(w_n3371_0[1]),.din(n3371));
	jspl jspl_w_n3372_0(.douta(w_n3372_0[0]),.doutb(w_n3372_0[1]),.din(n3372));
	jspl jspl_w_n3375_0(.douta(w_n3375_0[0]),.doutb(w_n3375_0[1]),.din(n3375));
	jspl jspl_w_n3378_0(.douta(w_n3378_0[0]),.doutb(w_n3378_0[1]),.din(n3378));
	jspl jspl_w_n3379_0(.douta(w_n3379_0[0]),.doutb(w_n3379_0[1]),.din(n3379));
	jspl3 jspl3_w_n3382_0(.douta(w_n3382_0[0]),.doutb(w_n3382_0[1]),.doutc(w_n3382_0[2]),.din(n3382));
	jspl jspl_w_n3384_0(.douta(w_n3384_0[0]),.doutb(w_n3384_0[1]),.din(n3384));
	jspl jspl_w_n3387_0(.douta(w_n3387_0[0]),.doutb(w_n3387_0[1]),.din(n3387));
	jspl jspl_w_n3388_0(.douta(w_n3388_0[0]),.doutb(w_n3388_0[1]),.din(n3388));
	jspl jspl_w_n3391_0(.douta(w_n3391_0[0]),.doutb(w_n3391_0[1]),.din(n3391));
	jspl jspl_w_n3392_0(.douta(w_n3392_0[0]),.doutb(w_n3392_0[1]),.din(n3392));
	jspl jspl_w_n3395_0(.douta(w_n3395_0[0]),.doutb(w_n3395_0[1]),.din(n3395));
	jspl jspl_w_n3398_0(.douta(w_n3398_0[0]),.doutb(w_n3398_0[1]),.din(n3398));
	jspl jspl_w_n3399_0(.douta(w_n3399_0[0]),.doutb(w_n3399_0[1]),.din(n3399));
	jspl3 jspl3_w_n3402_0(.douta(w_n3402_0[0]),.doutb(w_n3402_0[1]),.doutc(w_n3402_0[2]),.din(n3402));
	jspl3 jspl3_w_n3406_0(.douta(w_n3406_0[0]),.doutb(w_n3406_0[1]),.doutc(w_n3406_0[2]),.din(n3406));
	jspl jspl_w_n3409_0(.douta(w_n3409_0[0]),.doutb(w_n3409_0[1]),.din(n3409));
	jspl jspl_w_n3410_0(.douta(w_n3410_0[0]),.doutb(w_n3410_0[1]),.din(n3410));
	jspl jspl_w_n3412_0(.douta(w_n3412_0[0]),.doutb(w_n3412_0[1]),.din(n3412));
	jspl3 jspl3_w_n3415_0(.douta(w_n3415_0[0]),.doutb(w_n3415_0[1]),.doutc(w_n3415_0[2]),.din(n3415));
	jspl jspl_w_n3418_0(.douta(w_n3418_0[0]),.doutb(w_n3418_0[1]),.din(n3418));
	jspl jspl_w_n3419_0(.douta(w_n3419_0[0]),.doutb(w_n3419_0[1]),.din(n3419));
	jspl jspl_w_n3423_0(.douta(w_n3423_0[0]),.doutb(w_n3423_0[1]),.din(n3423));
	jspl jspl_w_n3444_0(.douta(w_n3444_0[0]),.doutb(w_n3444_0[1]),.din(n3444));
	jspl jspl_w_n3448_0(.douta(w_n3448_0[0]),.doutb(w_n3448_0[1]),.din(n3448));
	jspl jspl_w_n3449_0(.douta(w_n3449_0[0]),.doutb(w_n3449_0[1]),.din(n3449));
	jspl3 jspl3_w_n3452_0(.douta(w_n3452_0[0]),.doutb(w_n3452_0[1]),.doutc(w_n3452_0[2]),.din(n3452));
	jspl jspl_w_n3456_0(.douta(w_n3456_0[0]),.doutb(w_n3456_0[1]),.din(n3456));
	jspl jspl_w_n3457_0(.douta(w_n3457_0[0]),.doutb(w_n3457_0[1]),.din(n3457));
	jspl3 jspl3_w_n3460_0(.douta(w_n3460_0[0]),.doutb(w_n3460_0[1]),.doutc(w_n3460_0[2]),.din(n3460));
	jspl jspl_w_n3461_0(.douta(w_n3461_0[0]),.doutb(w_n3461_0[1]),.din(n3461));
	jspl3 jspl3_w_n3464_0(.douta(w_n3464_0[0]),.doutb(w_n3464_0[1]),.doutc(w_n3464_0[2]),.din(n3464));
	jspl jspl_w_n3467_0(.douta(w_n3467_0[0]),.doutb(w_n3467_0[1]),.din(n3467));
	jspl jspl_w_n3468_0(.douta(w_n3468_0[0]),.doutb(w_n3468_0[1]),.din(n3468));
	jspl jspl_w_n3471_0(.douta(w_n3471_0[0]),.doutb(w_n3471_0[1]),.din(n3471));
	jspl jspl_w_n3474_0(.douta(w_n3474_0[0]),.doutb(w_n3474_0[1]),.din(n3474));
	jspl jspl_w_n3475_0(.douta(w_n3475_0[0]),.doutb(w_n3475_0[1]),.din(n3475));
	jspl3 jspl3_w_n3478_0(.douta(w_n3478_0[0]),.doutb(w_n3478_0[1]),.doutc(w_n3478_0[2]),.din(n3478));
	jspl jspl_w_n3482_0(.douta(w_n3482_0[0]),.doutb(w_n3482_0[1]),.din(n3482));
	jspl jspl_w_n3483_0(.douta(w_n3483_0[0]),.doutb(w_n3483_0[1]),.din(n3483));
	jspl3 jspl3_w_n3486_0(.douta(w_n3486_0[0]),.doutb(w_n3486_0[1]),.doutc(w_n3486_0[2]),.din(n3486));
	jspl jspl_w_n3488_0(.douta(w_n3488_0[0]),.doutb(w_n3488_0[1]),.din(n3488));
	jspl jspl_w_n3491_0(.douta(w_n3491_0[0]),.doutb(w_n3491_0[1]),.din(n3491));
	jspl jspl_w_n3492_0(.douta(w_n3492_0[0]),.doutb(w_n3492_0[1]),.din(n3492));
	jspl3 jspl3_w_n3495_0(.douta(w_n3495_0[0]),.doutb(w_n3495_0[1]),.doutc(w_n3495_0[2]),.din(n3495));
	jspl jspl_w_n3496_0(.douta(w_n3496_0[0]),.doutb(w_n3496_0[1]),.din(n3496));
	jspl jspl_w_n3499_0(.douta(w_n3499_0[0]),.doutb(w_n3499_0[1]),.din(n3499));
	jspl jspl_w_n3500_0(.douta(w_n3500_0[0]),.doutb(w_n3500_0[1]),.din(n3500));
	jspl3 jspl3_w_n3503_0(.douta(w_n3503_0[0]),.doutb(w_n3503_0[1]),.doutc(w_n3503_0[2]),.din(n3503));
	jspl jspl_w_n3507_0(.douta(w_n3507_0[0]),.doutb(w_n3507_0[1]),.din(n3507));
	jspl jspl_w_n3508_0(.douta(w_n3508_0[0]),.doutb(w_n3508_0[1]),.din(n3508));
	jspl3 jspl3_w_n3511_0(.douta(w_n3511_0[0]),.doutb(w_n3511_0[1]),.doutc(w_n3511_0[2]),.din(n3511));
	jspl jspl_w_n3512_0(.douta(w_n3512_0[0]),.doutb(w_n3512_0[1]),.din(n3512));
	jspl jspl_w_n3516_0(.douta(w_n3516_0[0]),.doutb(w_n3516_0[1]),.din(n3516));
	jspl jspl_w_n3537_0(.douta(w_n3537_0[0]),.doutb(w_n3537_0[1]),.din(n3537));
	jspl jspl_w_n3541_0(.douta(w_n3541_0[0]),.doutb(w_n3541_0[1]),.din(n3541));
	jspl jspl_w_n3542_0(.douta(w_n3542_0[0]),.doutb(w_n3542_0[1]),.din(n3542));
	jspl3 jspl3_w_n3545_0(.douta(w_n3545_0[0]),.doutb(w_n3545_0[1]),.doutc(w_n3545_0[2]),.din(n3545));
	jspl3 jspl3_w_n3549_0(.douta(w_n3549_0[0]),.doutb(w_n3549_0[1]),.doutc(w_n3549_0[2]),.din(n3549));
	jspl jspl_w_n3552_0(.douta(w_n3552_0[0]),.doutb(w_n3552_0[1]),.din(n3552));
	jspl jspl_w_n3553_0(.douta(w_n3553_0[0]),.doutb(w_n3553_0[1]),.din(n3553));
	jspl jspl_w_n3555_0(.douta(w_n3555_0[0]),.doutb(w_n3555_0[1]),.din(n3555));
	jspl jspl_w_n3558_0(.douta(w_n3558_0[0]),.doutb(w_n3558_0[1]),.din(n3558));
	jspl jspl_w_n3559_0(.douta(w_n3559_0[0]),.doutb(w_n3559_0[1]),.din(n3559));
	jspl3 jspl3_w_n3562_0(.douta(w_n3562_0[0]),.doutb(w_n3562_0[1]),.doutc(w_n3562_0[2]),.din(n3562));
	jspl jspl_w_n3563_0(.douta(w_n3563_0[0]),.doutb(w_n3563_0[1]),.din(n3563));
	jspl3 jspl3_w_n3566_0(.douta(w_n3566_0[0]),.doutb(w_n3566_0[1]),.doutc(w_n3566_0[2]),.din(n3566));
	jspl jspl_w_n3569_0(.douta(w_n3569_0[0]),.doutb(w_n3569_0[1]),.din(n3569));
	jspl jspl_w_n3570_0(.douta(w_n3570_0[0]),.doutb(w_n3570_0[1]),.din(n3570));
	jspl jspl_w_n3573_0(.douta(w_n3573_0[0]),.doutb(w_n3573_0[1]),.din(n3573));
	jspl jspl_w_n3583_0(.douta(w_n3583_0[0]),.doutb(w_n3583_0[1]),.din(n3583));
	jspl jspl_w_n3587_0(.douta(w_n3587_0[0]),.doutb(w_n3587_0[1]),.din(n3587));
	jspl jspl_w_n3588_0(.douta(w_n3588_0[0]),.doutb(w_n3588_0[1]),.din(n3588));
	jspl3 jspl3_w_n3591_0(.douta(w_n3591_0[0]),.doutb(w_n3591_0[1]),.doutc(w_n3591_0[2]),.din(n3591));
	jspl jspl_w_n3595_0(.douta(w_n3595_0[0]),.doutb(w_n3595_0[1]),.din(n3595));
	jspl jspl_w_n3596_0(.douta(w_n3596_0[0]),.doutb(w_n3596_0[1]),.din(n3596));
	jspl3 jspl3_w_n3599_0(.douta(w_n3599_0[0]),.doutb(w_n3599_0[1]),.doutc(w_n3599_0[2]),.din(n3599));
	jspl jspl_w_n3603_0(.douta(w_n3603_0[0]),.doutb(w_n3603_0[1]),.din(n3603));
	jspl jspl_w_n3604_0(.douta(w_n3604_0[0]),.doutb(w_n3604_0[1]),.din(n3604));
	jspl3 jspl3_w_n3607_0(.douta(w_n3607_0[0]),.doutb(w_n3607_0[1]),.doutc(w_n3607_0[2]),.din(n3607));
	jspl jspl_w_n3608_0(.douta(w_n3608_0[0]),.doutb(w_n3608_0[1]),.din(n3608));
	jspl3 jspl3_w_n3611_0(.douta(w_n3611_0[0]),.doutb(w_n3611_0[1]),.doutc(w_n3611_0[2]),.din(n3611));
	jspl jspl_w_n3614_0(.douta(w_n3614_0[0]),.doutb(w_n3614_0[1]),.din(n3614));
	jspl jspl_w_n3615_0(.douta(w_n3615_0[0]),.doutb(w_n3615_0[1]),.din(n3615));
	jspl jspl_w_n3618_0(.douta(w_n3618_0[0]),.doutb(w_n3618_0[1]),.din(n3618));
	jspl jspl_w_n3619_0(.douta(w_n3619_0[0]),.doutb(w_n3619_0[1]),.din(n3619));
	jspl jspl_w_n3629_0(.douta(w_n3629_0[0]),.doutb(w_n3629_0[1]),.din(n3629));
	jspl jspl_w_n3633_0(.douta(w_n3633_0[0]),.doutb(w_n3633_0[1]),.din(n3633));
	jspl jspl_w_n3634_0(.douta(w_n3634_0[0]),.doutb(w_n3634_0[1]),.din(n3634));
	jspl3 jspl3_w_n3637_0(.douta(w_n3637_0[0]),.doutb(w_n3637_0[1]),.doutc(w_n3637_0[2]),.din(n3637));
	jspl3 jspl3_w_n3641_0(.douta(w_n3641_0[0]),.doutb(w_n3641_0[1]),.doutc(w_n3641_0[2]),.din(n3641));
	jspl jspl_w_n3644_0(.douta(w_n3644_0[0]),.doutb(w_n3644_0[1]),.din(n3644));
	jspl jspl_w_n3645_0(.douta(w_n3645_0[0]),.doutb(w_n3645_0[1]),.din(n3645));
	jspl jspl_w_n3647_0(.douta(w_n3647_0[0]),.doutb(w_n3647_0[1]),.din(n3647));
	jspl jspl_w_n3650_0(.douta(w_n3650_0[0]),.doutb(w_n3650_0[1]),.din(n3650));
	jspl jspl_w_n3651_0(.douta(w_n3651_0[0]),.doutb(w_n3651_0[1]),.din(n3651));
	jspl3 jspl3_w_n3654_0(.douta(w_n3654_0[0]),.doutb(w_n3654_0[1]),.doutc(w_n3654_0[2]),.din(n3654));
	jspl jspl_w_n3655_0(.douta(w_n3655_0[0]),.doutb(w_n3655_0[1]),.din(n3655));
	jspl3 jspl3_w_n3658_0(.douta(w_n3658_0[0]),.doutb(w_n3658_0[1]),.doutc(w_n3658_0[2]),.din(n3658));
	jspl jspl_w_n3661_0(.douta(w_n3661_0[0]),.doutb(w_n3661_0[1]),.din(n3661));
	jspl jspl_w_n3662_0(.douta(w_n3662_0[0]),.doutb(w_n3662_0[1]),.din(n3662));
	jspl jspl_w_n3665_0(.douta(w_n3665_0[0]),.doutb(w_n3665_0[1]),.din(n3665));
	jspl jspl_w_n3675_0(.douta(w_n3675_0[0]),.doutb(w_n3675_0[1]),.din(n3675));
	jspl jspl_w_n3679_0(.douta(w_n3679_0[0]),.doutb(w_n3679_0[1]),.din(n3679));
	jspl jspl_w_n3680_0(.douta(w_n3680_0[0]),.doutb(w_n3680_0[1]),.din(n3680));
	jspl3 jspl3_w_n3683_0(.douta(w_n3683_0[0]),.doutb(w_n3683_0[1]),.doutc(w_n3683_0[2]),.din(n3683));
	jspl jspl_w_n3687_0(.douta(w_n3687_0[0]),.doutb(w_n3687_0[1]),.din(n3687));
	jspl jspl_w_n3688_0(.douta(w_n3688_0[0]),.doutb(w_n3688_0[1]),.din(n3688));
	jspl3 jspl3_w_n3691_0(.douta(w_n3691_0[0]),.doutb(w_n3691_0[1]),.doutc(w_n3691_0[2]),.din(n3691));
	jspl jspl_w_n3695_0(.douta(w_n3695_0[0]),.doutb(w_n3695_0[1]),.din(n3695));
	jspl jspl_w_n3696_0(.douta(w_n3696_0[0]),.doutb(w_n3696_0[1]),.din(n3696));
	jspl3 jspl3_w_n3699_0(.douta(w_n3699_0[0]),.doutb(w_n3699_0[1]),.doutc(w_n3699_0[2]),.din(n3699));
	jspl jspl_w_n3700_0(.douta(w_n3700_0[0]),.doutb(w_n3700_0[1]),.din(n3700));
	jspl3 jspl3_w_n3703_0(.douta(w_n3703_0[0]),.doutb(w_n3703_0[1]),.doutc(w_n3703_0[2]),.din(n3703));
	jspl jspl_w_n3706_0(.douta(w_n3706_0[0]),.doutb(w_n3706_0[1]),.din(n3706));
	jspl jspl_w_n3707_0(.douta(w_n3707_0[0]),.doutb(w_n3707_0[1]),.din(n3707));
	jspl jspl_w_n3710_0(.douta(w_n3710_0[0]),.doutb(w_n3710_0[1]),.din(n3710));
	jspl jspl_w_n3711_0(.douta(w_n3711_0[0]),.doutb(w_n3711_0[1]),.din(n3711));
	jspl jspl_w_n3721_0(.douta(w_n3721_0[0]),.doutb(w_n3721_0[1]),.din(n3721));
	jspl jspl_w_n3725_0(.douta(w_n3725_0[0]),.doutb(w_n3725_0[1]),.din(n3725));
	jspl jspl_w_n3726_0(.douta(w_n3726_0[0]),.doutb(w_n3726_0[1]),.din(n3726));
	jspl3 jspl3_w_n3729_0(.douta(w_n3729_0[0]),.doutb(w_n3729_0[1]),.doutc(w_n3729_0[2]),.din(n3729));
	jspl3 jspl3_w_n3733_0(.douta(w_n3733_0[0]),.doutb(w_n3733_0[1]),.doutc(w_n3733_0[2]),.din(n3733));
	jspl jspl_w_n3736_0(.douta(w_n3736_0[0]),.doutb(w_n3736_0[1]),.din(n3736));
	jspl jspl_w_n3737_0(.douta(w_n3737_0[0]),.doutb(w_n3737_0[1]),.din(n3737));
	jspl jspl_w_n3739_0(.douta(w_n3739_0[0]),.doutb(w_n3739_0[1]),.din(n3739));
	jspl jspl_w_n3742_0(.douta(w_n3742_0[0]),.doutb(w_n3742_0[1]),.din(n3742));
	jspl jspl_w_n3743_0(.douta(w_n3743_0[0]),.doutb(w_n3743_0[1]),.din(n3743));
	jspl3 jspl3_w_n3746_0(.douta(w_n3746_0[0]),.doutb(w_n3746_0[1]),.doutc(w_n3746_0[2]),.din(n3746));
	jspl jspl_w_n3747_0(.douta(w_n3747_0[0]),.doutb(w_n3747_0[1]),.din(n3747));
	jspl3 jspl3_w_n3750_0(.douta(w_n3750_0[0]),.doutb(w_n3750_0[1]),.doutc(w_n3750_0[2]),.din(n3750));
	jspl jspl_w_n3753_0(.douta(w_n3753_0[0]),.doutb(w_n3753_0[1]),.din(n3753));
	jspl jspl_w_n3754_0(.douta(w_n3754_0[0]),.doutb(w_n3754_0[1]),.din(n3754));
	jspl jspl_w_n3757_0(.douta(w_n3757_0[0]),.doutb(w_n3757_0[1]),.din(n3757));
	jspl jspl_w_n3767_0(.douta(w_n3767_0[0]),.doutb(w_n3767_0[1]),.din(n3767));
	jspl jspl_w_n3771_0(.douta(w_n3771_0[0]),.doutb(w_n3771_0[1]),.din(n3771));
	jspl jspl_w_n3772_0(.douta(w_n3772_0[0]),.doutb(w_n3772_0[1]),.din(n3772));
	jspl3 jspl3_w_n3775_0(.douta(w_n3775_0[0]),.doutb(w_n3775_0[1]),.doutc(w_n3775_0[2]),.din(n3775));
	jspl jspl_w_n3779_0(.douta(w_n3779_0[0]),.doutb(w_n3779_0[1]),.din(n3779));
	jspl jspl_w_n3780_0(.douta(w_n3780_0[0]),.doutb(w_n3780_0[1]),.din(n3780));
	jspl3 jspl3_w_n3783_0(.douta(w_n3783_0[0]),.doutb(w_n3783_0[1]),.doutc(w_n3783_0[2]),.din(n3783));
	jspl jspl_w_n3787_0(.douta(w_n3787_0[0]),.doutb(w_n3787_0[1]),.din(n3787));
	jspl jspl_w_n3788_0(.douta(w_n3788_0[0]),.doutb(w_n3788_0[1]),.din(n3788));
	jspl3 jspl3_w_n3791_0(.douta(w_n3791_0[0]),.doutb(w_n3791_0[1]),.doutc(w_n3791_0[2]),.din(n3791));
	jspl jspl_w_n3792_0(.douta(w_n3792_0[0]),.doutb(w_n3792_0[1]),.din(n3792));
	jspl3 jspl3_w_n3795_0(.douta(w_n3795_0[0]),.doutb(w_n3795_0[1]),.doutc(w_n3795_0[2]),.din(n3795));
	jspl jspl_w_n3798_0(.douta(w_n3798_0[0]),.doutb(w_n3798_0[1]),.din(n3798));
	jspl jspl_w_n3799_0(.douta(w_n3799_0[0]),.doutb(w_n3799_0[1]),.din(n3799));
	jspl jspl_w_n3802_0(.douta(w_n3802_0[0]),.doutb(w_n3802_0[1]),.din(n3802));
	jspl jspl_w_n3803_0(.douta(w_n3803_0[0]),.doutb(w_n3803_0[1]),.din(n3803));
	jspl jspl_w_n3813_0(.douta(w_n3813_0[0]),.doutb(w_n3813_0[1]),.din(n3813));
	jspl jspl_w_n3817_0(.douta(w_n3817_0[0]),.doutb(w_n3817_0[1]),.din(n3817));
	jspl jspl_w_n3818_0(.douta(w_n3818_0[0]),.doutb(w_n3818_0[1]),.din(n3818));
	jspl3 jspl3_w_n3821_0(.douta(w_n3821_0[0]),.doutb(w_n3821_0[1]),.doutc(w_n3821_0[2]),.din(n3821));
	jspl3 jspl3_w_n3825_0(.douta(w_n3825_0[0]),.doutb(w_n3825_0[1]),.doutc(w_n3825_0[2]),.din(n3825));
	jspl jspl_w_n3828_0(.douta(w_n3828_0[0]),.doutb(w_n3828_0[1]),.din(n3828));
	jspl jspl_w_n3829_0(.douta(w_n3829_0[0]),.doutb(w_n3829_0[1]),.din(n3829));
	jspl jspl_w_n3831_0(.douta(w_n3831_0[0]),.doutb(w_n3831_0[1]),.din(n3831));
	jspl jspl_w_n3834_0(.douta(w_n3834_0[0]),.doutb(w_n3834_0[1]),.din(n3834));
	jspl jspl_w_n3835_0(.douta(w_n3835_0[0]),.doutb(w_n3835_0[1]),.din(n3835));
	jspl3 jspl3_w_n3838_0(.douta(w_n3838_0[0]),.doutb(w_n3838_0[1]),.doutc(w_n3838_0[2]),.din(n3838));
	jspl jspl_w_n3839_0(.douta(w_n3839_0[0]),.doutb(w_n3839_0[1]),.din(n3839));
	jspl3 jspl3_w_n3842_0(.douta(w_n3842_0[0]),.doutb(w_n3842_0[1]),.doutc(w_n3842_0[2]),.din(n3842));
	jspl jspl_w_n3845_0(.douta(w_n3845_0[0]),.doutb(w_n3845_0[1]),.din(n3845));
	jspl jspl_w_n3846_0(.douta(w_n3846_0[0]),.doutb(w_n3846_0[1]),.din(n3846));
	jspl jspl_w_n3849_0(.douta(w_n3849_0[0]),.doutb(w_n3849_0[1]),.din(n3849));
	jspl jspl_w_n3859_0(.douta(w_n3859_0[0]),.doutb(w_n3859_0[1]),.din(n3859));
	jspl jspl_w_n3863_0(.douta(w_n3863_0[0]),.doutb(w_n3863_0[1]),.din(n3863));
	jspl jspl_w_n3864_0(.douta(w_n3864_0[0]),.doutb(w_n3864_0[1]),.din(n3864));
	jspl3 jspl3_w_n3867_0(.douta(w_n3867_0[0]),.doutb(w_n3867_0[1]),.doutc(w_n3867_0[2]),.din(n3867));
	jspl jspl_w_n3871_0(.douta(w_n3871_0[0]),.doutb(w_n3871_0[1]),.din(n3871));
	jspl jspl_w_n3872_0(.douta(w_n3872_0[0]),.doutb(w_n3872_0[1]),.din(n3872));
	jspl3 jspl3_w_n3875_0(.douta(w_n3875_0[0]),.doutb(w_n3875_0[1]),.doutc(w_n3875_0[2]),.din(n3875));
	jspl jspl_w_n3879_0(.douta(w_n3879_0[0]),.doutb(w_n3879_0[1]),.din(n3879));
	jspl jspl_w_n3880_0(.douta(w_n3880_0[0]),.doutb(w_n3880_0[1]),.din(n3880));
	jspl3 jspl3_w_n3883_0(.douta(w_n3883_0[0]),.doutb(w_n3883_0[1]),.doutc(w_n3883_0[2]),.din(n3883));
	jspl jspl_w_n3884_0(.douta(w_n3884_0[0]),.doutb(w_n3884_0[1]),.din(n3884));
	jspl3 jspl3_w_n3887_0(.douta(w_n3887_0[0]),.doutb(w_n3887_0[1]),.doutc(w_n3887_0[2]),.din(n3887));
	jspl jspl_w_n3890_0(.douta(w_n3890_0[0]),.doutb(w_n3890_0[1]),.din(n3890));
	jspl jspl_w_n3891_0(.douta(w_n3891_0[0]),.doutb(w_n3891_0[1]),.din(n3891));
	jspl jspl_w_n3894_0(.douta(w_n3894_0[0]),.doutb(w_n3894_0[1]),.din(n3894));
	jspl jspl_w_n3895_0(.douta(w_n3895_0[0]),.doutb(w_n3895_0[1]),.din(n3895));
	jspl jspl_w_n3905_0(.douta(w_n3905_0[0]),.doutb(w_n3905_0[1]),.din(n3905));
	jspl jspl_w_n3909_0(.douta(w_n3909_0[0]),.doutb(w_n3909_0[1]),.din(n3909));
	jspl jspl_w_n3910_0(.douta(w_n3910_0[0]),.doutb(w_n3910_0[1]),.din(n3910));
	jspl3 jspl3_w_n3913_0(.douta(w_n3913_0[0]),.doutb(w_n3913_0[1]),.doutc(w_n3913_0[2]),.din(n3913));
	jspl3 jspl3_w_n3917_0(.douta(w_n3917_0[0]),.doutb(w_n3917_0[1]),.doutc(w_n3917_0[2]),.din(n3917));
	jspl jspl_w_n3920_0(.douta(w_n3920_0[0]),.doutb(w_n3920_0[1]),.din(n3920));
	jspl jspl_w_n3921_0(.douta(w_n3921_0[0]),.doutb(w_n3921_0[1]),.din(n3921));
	jspl jspl_w_n3923_0(.douta(w_n3923_0[0]),.doutb(w_n3923_0[1]),.din(n3923));
	jspl jspl_w_n3926_0(.douta(w_n3926_0[0]),.doutb(w_n3926_0[1]),.din(n3926));
	jspl jspl_w_n3927_0(.douta(w_n3927_0[0]),.doutb(w_n3927_0[1]),.din(n3927));
	jspl3 jspl3_w_n3930_0(.douta(w_n3930_0[0]),.doutb(w_n3930_0[1]),.doutc(w_n3930_0[2]),.din(n3930));
	jspl jspl_w_n3931_0(.douta(w_n3931_0[0]),.doutb(w_n3931_0[1]),.din(n3931));
	jspl3 jspl3_w_n3934_0(.douta(w_n3934_0[0]),.doutb(w_n3934_0[1]),.doutc(w_n3934_0[2]),.din(n3934));
	jspl jspl_w_n3937_0(.douta(w_n3937_0[0]),.doutb(w_n3937_0[1]),.din(n3937));
	jspl jspl_w_n3938_0(.douta(w_n3938_0[0]),.doutb(w_n3938_0[1]),.din(n3938));
	jspl jspl_w_n3941_0(.douta(w_n3941_0[0]),.doutb(w_n3941_0[1]),.din(n3941));
	jspl jspl_w_n3951_0(.douta(w_n3951_0[0]),.doutb(w_n3951_0[1]),.din(n3951));
	jspl jspl_w_n3955_0(.douta(w_n3955_0[0]),.doutb(w_n3955_0[1]),.din(n3955));
	jspl jspl_w_n3956_0(.douta(w_n3956_0[0]),.doutb(w_n3956_0[1]),.din(n3956));
	jspl3 jspl3_w_n3959_0(.douta(w_n3959_0[0]),.doutb(w_n3959_0[1]),.doutc(w_n3959_0[2]),.din(n3959));
	jspl jspl_w_n3963_0(.douta(w_n3963_0[0]),.doutb(w_n3963_0[1]),.din(n3963));
	jspl jspl_w_n3964_0(.douta(w_n3964_0[0]),.doutb(w_n3964_0[1]),.din(n3964));
	jspl3 jspl3_w_n3967_0(.douta(w_n3967_0[0]),.doutb(w_n3967_0[1]),.doutc(w_n3967_0[2]),.din(n3967));
	jspl jspl_w_n3971_0(.douta(w_n3971_0[0]),.doutb(w_n3971_0[1]),.din(n3971));
	jspl jspl_w_n3972_0(.douta(w_n3972_0[0]),.doutb(w_n3972_0[1]),.din(n3972));
	jspl3 jspl3_w_n3975_0(.douta(w_n3975_0[0]),.doutb(w_n3975_0[1]),.doutc(w_n3975_0[2]),.din(n3975));
	jspl jspl_w_n3976_0(.douta(w_n3976_0[0]),.doutb(w_n3976_0[1]),.din(n3976));
	jspl3 jspl3_w_n3979_0(.douta(w_n3979_0[0]),.doutb(w_n3979_0[1]),.doutc(w_n3979_0[2]),.din(n3979));
	jspl jspl_w_n3982_0(.douta(w_n3982_0[0]),.doutb(w_n3982_0[1]),.din(n3982));
	jspl jspl_w_n3983_0(.douta(w_n3983_0[0]),.doutb(w_n3983_0[1]),.din(n3983));
	jspl jspl_w_n3986_0(.douta(w_n3986_0[0]),.doutb(w_n3986_0[1]),.din(n3986));
	jspl jspl_w_n3987_0(.douta(w_n3987_0[0]),.doutb(w_n3987_0[1]),.din(n3987));
	jspl jspl_w_n3997_0(.douta(w_n3997_0[0]),.doutb(w_n3997_0[1]),.din(n3997));
	jspl jspl_w_n4001_0(.douta(w_n4001_0[0]),.doutb(w_n4001_0[1]),.din(n4001));
	jspl jspl_w_n4002_0(.douta(w_n4002_0[0]),.doutb(w_n4002_0[1]),.din(n4002));
	jspl3 jspl3_w_n4005_0(.douta(w_n4005_0[0]),.doutb(w_n4005_0[1]),.doutc(w_n4005_0[2]),.din(n4005));
	jspl3 jspl3_w_n4009_0(.douta(w_n4009_0[0]),.doutb(w_n4009_0[1]),.doutc(w_n4009_0[2]),.din(n4009));
	jspl jspl_w_n4012_0(.douta(w_n4012_0[0]),.doutb(w_n4012_0[1]),.din(n4012));
	jspl jspl_w_n4013_0(.douta(w_n4013_0[0]),.doutb(w_n4013_0[1]),.din(n4013));
	jspl jspl_w_n4015_0(.douta(w_n4015_0[0]),.doutb(w_n4015_0[1]),.din(n4015));
	jspl jspl_w_n4018_0(.douta(w_n4018_0[0]),.doutb(w_n4018_0[1]),.din(n4018));
	jspl jspl_w_n4019_0(.douta(w_n4019_0[0]),.doutb(w_n4019_0[1]),.din(n4019));
	jspl3 jspl3_w_n4022_0(.douta(w_n4022_0[0]),.doutb(w_n4022_0[1]),.doutc(w_n4022_0[2]),.din(n4022));
	jspl jspl_w_n4023_0(.douta(w_n4023_0[0]),.doutb(w_n4023_0[1]),.din(n4023));
	jspl3 jspl3_w_n4026_0(.douta(w_n4026_0[0]),.doutb(w_n4026_0[1]),.doutc(w_n4026_0[2]),.din(n4026));
	jspl jspl_w_n4029_0(.douta(w_n4029_0[0]),.doutb(w_n4029_0[1]),.din(n4029));
	jspl jspl_w_n4030_0(.douta(w_n4030_0[0]),.doutb(w_n4030_0[1]),.din(n4030));
	jspl jspl_w_n4033_0(.douta(w_n4033_0[0]),.doutb(w_n4033_0[1]),.din(n4033));
	jspl jspl_w_n4043_0(.douta(w_n4043_0[0]),.doutb(w_n4043_0[1]),.din(n4043));
	jspl jspl_w_n4047_0(.douta(w_n4047_0[0]),.doutb(w_n4047_0[1]),.din(n4047));
	jspl jspl_w_n4048_0(.douta(w_n4048_0[0]),.doutb(w_n4048_0[1]),.din(n4048));
	jspl3 jspl3_w_n4051_0(.douta(w_n4051_0[0]),.doutb(w_n4051_0[1]),.doutc(w_n4051_0[2]),.din(n4051));
	jspl jspl_w_n4055_0(.douta(w_n4055_0[0]),.doutb(w_n4055_0[1]),.din(n4055));
	jspl jspl_w_n4056_0(.douta(w_n4056_0[0]),.doutb(w_n4056_0[1]),.din(n4056));
	jspl3 jspl3_w_n4059_0(.douta(w_n4059_0[0]),.doutb(w_n4059_0[1]),.doutc(w_n4059_0[2]),.din(n4059));
	jspl jspl_w_n4063_0(.douta(w_n4063_0[0]),.doutb(w_n4063_0[1]),.din(n4063));
	jspl jspl_w_n4064_0(.douta(w_n4064_0[0]),.doutb(w_n4064_0[1]),.din(n4064));
	jspl3 jspl3_w_n4067_0(.douta(w_n4067_0[0]),.doutb(w_n4067_0[1]),.doutc(w_n4067_0[2]),.din(n4067));
	jspl jspl_w_n4068_0(.douta(w_n4068_0[0]),.doutb(w_n4068_0[1]),.din(n4068));
	jspl3 jspl3_w_n4071_0(.douta(w_n4071_0[0]),.doutb(w_n4071_0[1]),.doutc(w_n4071_0[2]),.din(n4071));
	jspl jspl_w_n4074_0(.douta(w_n4074_0[0]),.doutb(w_n4074_0[1]),.din(n4074));
	jspl jspl_w_n4075_0(.douta(w_n4075_0[0]),.doutb(w_n4075_0[1]),.din(n4075));
	jspl jspl_w_n4078_0(.douta(w_n4078_0[0]),.doutb(w_n4078_0[1]),.din(n4078));
	jspl jspl_w_n4079_0(.douta(w_n4079_0[0]),.doutb(w_n4079_0[1]),.din(n4079));
	jspl jspl_w_n4089_0(.douta(w_n4089_0[0]),.doutb(w_n4089_0[1]),.din(n4089));
	jspl jspl_w_n4093_0(.douta(w_n4093_0[0]),.doutb(w_n4093_0[1]),.din(n4093));
	jspl jspl_w_n4094_0(.douta(w_n4094_0[0]),.doutb(w_n4094_0[1]),.din(n4094));
	jspl3 jspl3_w_n4097_0(.douta(w_n4097_0[0]),.doutb(w_n4097_0[1]),.doutc(w_n4097_0[2]),.din(n4097));
	jspl3 jspl3_w_n4101_0(.douta(w_n4101_0[0]),.doutb(w_n4101_0[1]),.doutc(w_n4101_0[2]),.din(n4101));
	jspl jspl_w_n4104_0(.douta(w_n4104_0[0]),.doutb(w_n4104_0[1]),.din(n4104));
	jspl jspl_w_n4105_0(.douta(w_n4105_0[0]),.doutb(w_n4105_0[1]),.din(n4105));
	jspl jspl_w_n4107_0(.douta(w_n4107_0[0]),.doutb(w_n4107_0[1]),.din(n4107));
	jspl jspl_w_n4110_0(.douta(w_n4110_0[0]),.doutb(w_n4110_0[1]),.din(n4110));
	jspl jspl_w_n4111_0(.douta(w_n4111_0[0]),.doutb(w_n4111_0[1]),.din(n4111));
	jspl3 jspl3_w_n4114_0(.douta(w_n4114_0[0]),.doutb(w_n4114_0[1]),.doutc(w_n4114_0[2]),.din(n4114));
	jspl jspl_w_n4115_0(.douta(w_n4115_0[0]),.doutb(w_n4115_0[1]),.din(n4115));
	jspl3 jspl3_w_n4118_0(.douta(w_n4118_0[0]),.doutb(w_n4118_0[1]),.doutc(w_n4118_0[2]),.din(n4118));
	jspl jspl_w_n4121_0(.douta(w_n4121_0[0]),.doutb(w_n4121_0[1]),.din(n4121));
	jspl jspl_w_n4122_0(.douta(w_n4122_0[0]),.doutb(w_n4122_0[1]),.din(n4122));
	jspl jspl_w_n4125_0(.douta(w_n4125_0[0]),.doutb(w_n4125_0[1]),.din(n4125));
	jspl jspl_w_n4135_0(.douta(w_n4135_0[0]),.doutb(w_n4135_0[1]),.din(n4135));
	jspl jspl_w_n4139_0(.douta(w_n4139_0[0]),.doutb(w_n4139_0[1]),.din(n4139));
	jspl jspl_w_n4140_0(.douta(w_n4140_0[0]),.doutb(w_n4140_0[1]),.din(n4140));
	jspl3 jspl3_w_n4143_0(.douta(w_n4143_0[0]),.doutb(w_n4143_0[1]),.doutc(w_n4143_0[2]),.din(n4143));
	jspl jspl_w_n4147_0(.douta(w_n4147_0[0]),.doutb(w_n4147_0[1]),.din(n4147));
	jspl jspl_w_n4148_0(.douta(w_n4148_0[0]),.doutb(w_n4148_0[1]),.din(n4148));
	jspl3 jspl3_w_n4151_0(.douta(w_n4151_0[0]),.doutb(w_n4151_0[1]),.doutc(w_n4151_0[2]),.din(n4151));
	jspl jspl_w_n4155_0(.douta(w_n4155_0[0]),.doutb(w_n4155_0[1]),.din(n4155));
	jspl jspl_w_n4156_0(.douta(w_n4156_0[0]),.doutb(w_n4156_0[1]),.din(n4156));
	jspl3 jspl3_w_n4159_0(.douta(w_n4159_0[0]),.doutb(w_n4159_0[1]),.doutc(w_n4159_0[2]),.din(n4159));
	jspl jspl_w_n4160_0(.douta(w_n4160_0[0]),.doutb(w_n4160_0[1]),.din(n4160));
	jspl3 jspl3_w_n4163_0(.douta(w_n4163_0[0]),.doutb(w_n4163_0[1]),.doutc(w_n4163_0[2]),.din(n4163));
	jspl jspl_w_n4166_0(.douta(w_n4166_0[0]),.doutb(w_n4166_0[1]),.din(n4166));
	jspl jspl_w_n4167_0(.douta(w_n4167_0[0]),.doutb(w_n4167_0[1]),.din(n4167));
	jspl jspl_w_n4170_0(.douta(w_n4170_0[0]),.doutb(w_n4170_0[1]),.din(n4170));
	jspl jspl_w_n4171_0(.douta(w_n4171_0[0]),.doutb(w_n4171_0[1]),.din(n4171));
	jspl jspl_w_n4181_0(.douta(w_n4181_0[0]),.doutb(w_n4181_0[1]),.din(n4181));
	jspl jspl_w_n4185_0(.douta(w_n4185_0[0]),.doutb(w_n4185_0[1]),.din(n4185));
	jspl jspl_w_n4186_0(.douta(w_n4186_0[0]),.doutb(w_n4186_0[1]),.din(n4186));
	jspl3 jspl3_w_n4189_0(.douta(w_n4189_0[0]),.doutb(w_n4189_0[1]),.doutc(w_n4189_0[2]),.din(n4189));
	jspl3 jspl3_w_n4193_0(.douta(w_n4193_0[0]),.doutb(w_n4193_0[1]),.doutc(w_n4193_0[2]),.din(n4193));
	jspl jspl_w_n4196_0(.douta(w_n4196_0[0]),.doutb(w_n4196_0[1]),.din(n4196));
	jspl jspl_w_n4197_0(.douta(w_n4197_0[0]),.doutb(w_n4197_0[1]),.din(n4197));
	jspl jspl_w_n4199_0(.douta(w_n4199_0[0]),.doutb(w_n4199_0[1]),.din(n4199));
	jspl jspl_w_n4202_0(.douta(w_n4202_0[0]),.doutb(w_n4202_0[1]),.din(n4202));
	jspl jspl_w_n4203_0(.douta(w_n4203_0[0]),.doutb(w_n4203_0[1]),.din(n4203));
	jspl3 jspl3_w_n4206_0(.douta(w_n4206_0[0]),.doutb(w_n4206_0[1]),.doutc(w_n4206_0[2]),.din(n4206));
	jspl jspl_w_n4207_0(.douta(w_n4207_0[0]),.doutb(w_n4207_0[1]),.din(n4207));
	jspl3 jspl3_w_n4210_0(.douta(w_n4210_0[0]),.doutb(w_n4210_0[1]),.doutc(w_n4210_0[2]),.din(n4210));
	jspl jspl_w_n4213_0(.douta(w_n4213_0[0]),.doutb(w_n4213_0[1]),.din(n4213));
	jspl jspl_w_n4214_0(.douta(w_n4214_0[0]),.doutb(w_n4214_0[1]),.din(n4214));
	jspl jspl_w_n4217_0(.douta(w_n4217_0[0]),.doutb(w_n4217_0[1]),.din(n4217));
	jspl jspl_w_n4227_0(.douta(w_n4227_0[0]),.doutb(w_n4227_0[1]),.din(n4227));
	jspl jspl_w_n4231_0(.douta(w_n4231_0[0]),.doutb(w_n4231_0[1]),.din(n4231));
	jspl jspl_w_n4232_0(.douta(w_n4232_0[0]),.doutb(w_n4232_0[1]),.din(n4232));
	jspl3 jspl3_w_n4235_0(.douta(w_n4235_0[0]),.doutb(w_n4235_0[1]),.doutc(w_n4235_0[2]),.din(n4235));
	jspl jspl_w_n4239_0(.douta(w_n4239_0[0]),.doutb(w_n4239_0[1]),.din(n4239));
	jspl jspl_w_n4240_0(.douta(w_n4240_0[0]),.doutb(w_n4240_0[1]),.din(n4240));
	jspl3 jspl3_w_n4243_0(.douta(w_n4243_0[0]),.doutb(w_n4243_0[1]),.doutc(w_n4243_0[2]),.din(n4243));
	jspl jspl_w_n4245_0(.douta(w_n4245_0[0]),.doutb(w_n4245_0[1]),.din(n4245));
	jspl jspl_w_n4246_0(.douta(w_n4246_0[0]),.doutb(w_n4246_0[1]),.din(n4246));
	jspl jspl_w_n4247_0(.douta(w_n4247_0[0]),.doutb(w_n4247_0[1]),.din(n4247));
	jspl3 jspl3_w_n4248_0(.douta(w_n4248_0[0]),.doutb(w_n4248_0[1]),.doutc(w_n4248_0[2]),.din(n4248));
	jspl jspl_w_n4249_0(.douta(w_n4249_0[0]),.doutb(w_n4249_0[1]),.din(n4249));
	jspl jspl_w_n4252_0(.douta(w_n4252_0[0]),.doutb(w_n4252_0[1]),.din(n4252));
	jspl jspl_w_n4253_0(.douta(w_n4253_0[0]),.doutb(w_n4253_0[1]),.din(n4253));
	jspl3 jspl3_w_n4256_0(.douta(w_n4256_0[0]),.doutb(w_n4256_0[1]),.doutc(w_n4256_0[2]),.din(n4256));
	jspl jspl_w_n4259_0(.douta(w_n4259_0[0]),.doutb(w_n4259_0[1]),.din(n4259));
	jspl jspl_w_n4269_0(.douta(w_n4269_0[0]),.doutb(w_n4269_0[1]),.din(n4269));
	jspl jspl_w_n4274_0(.douta(w_n4274_0[0]),.doutb(w_n4274_0[1]),.din(n4274));
	jspl jspl_w_n4290_0(.douta(w_n4290_0[0]),.doutb(w_n4290_0[1]),.din(n4290));
	jspl3 jspl3_w_n4293_0(.douta(w_n4293_0[0]),.doutb(w_n4293_0[1]),.doutc(w_n4293_0[2]),.din(n4293));
	jspl jspl_w_n4298_0(.douta(w_n4298_0[0]),.doutb(w_n4298_0[1]),.din(n4298));
	jspl jspl_w_n4308_0(.douta(w_n4308_0[0]),.doutb(w_n4308_0[1]),.din(n4308));
	jspl jspl_w_n4309_0(.douta(w_n4309_0[0]),.doutb(w_n4309_0[1]),.din(n4309));
	jspl jspl_w_n4313_0(.douta(w_n4313_0[0]),.doutb(w_n4313_0[1]),.din(n4313));
	jspl jspl_w_n4314_0(.douta(w_n4314_0[0]),.doutb(w_n4314_0[1]),.din(n4314));
	jspl jspl_w_n4324_0(.douta(w_n4324_0[0]),.doutb(w_n4324_0[1]),.din(n4324));
	jspl jspl_w_n4344_0(.douta(w_n4344_0[0]),.doutb(w_n4344_0[1]),.din(n4344));
	jspl3 jspl3_w_n4452_0(.douta(w_n4452_0[0]),.doutb(w_n4452_0[1]),.doutc(w_n4452_0[2]),.din(n4452));
	jspl3 jspl3_w_n4452_1(.douta(w_n4452_1[0]),.doutb(w_n4452_1[1]),.doutc(w_n4452_1[2]),.din(w_n4452_0[0]));
	jspl3 jspl3_w_n4452_2(.douta(w_n4452_2[0]),.doutb(w_n4452_2[1]),.doutc(w_n4452_2[2]),.din(w_n4452_0[1]));
	jspl3 jspl3_w_n4452_3(.douta(w_n4452_3[0]),.doutb(w_n4452_3[1]),.doutc(w_n4452_3[2]),.din(w_n4452_0[2]));
	jspl3 jspl3_w_n4452_4(.douta(w_n4452_4[0]),.doutb(w_n4452_4[1]),.doutc(w_n4452_4[2]),.din(w_n4452_1[0]));
	jspl3 jspl3_w_n4452_5(.douta(w_n4452_5[0]),.doutb(w_n4452_5[1]),.doutc(w_n4452_5[2]),.din(w_n4452_1[1]));
	jspl3 jspl3_w_n4452_6(.douta(w_n4452_6[0]),.doutb(w_n4452_6[1]),.doutc(w_n4452_6[2]),.din(w_n4452_1[2]));
	jspl3 jspl3_w_n4452_7(.douta(w_n4452_7[0]),.doutb(w_n4452_7[1]),.doutc(w_n4452_7[2]),.din(w_n4452_2[0]));
	jspl3 jspl3_w_n4452_8(.douta(w_n4452_8[0]),.doutb(w_n4452_8[1]),.doutc(w_n4452_8[2]),.din(w_n4452_2[1]));
	jspl3 jspl3_w_n4452_9(.douta(w_n4452_9[0]),.doutb(w_n4452_9[1]),.doutc(w_n4452_9[2]),.din(w_n4452_2[2]));
	jspl3 jspl3_w_n4452_10(.douta(w_n4452_10[0]),.doutb(w_n4452_10[1]),.doutc(w_n4452_10[2]),.din(w_n4452_3[0]));
	jspl3 jspl3_w_n4452_11(.douta(w_n4452_11[0]),.doutb(w_n4452_11[1]),.doutc(w_n4452_11[2]),.din(w_n4452_3[1]));
	jspl3 jspl3_w_n4452_12(.douta(w_n4452_12[0]),.doutb(w_n4452_12[1]),.doutc(w_n4452_12[2]),.din(w_n4452_3[2]));
	jspl3 jspl3_w_n4452_13(.douta(w_n4452_13[0]),.doutb(w_n4452_13[1]),.doutc(w_n4452_13[2]),.din(w_n4452_4[0]));
	jspl3 jspl3_w_n4452_14(.douta(w_n4452_14[0]),.doutb(w_n4452_14[1]),.doutc(w_n4452_14[2]),.din(w_n4452_4[1]));
	jspl3 jspl3_w_n4452_15(.douta(w_n4452_15[0]),.doutb(w_n4452_15[1]),.doutc(w_n4452_15[2]),.din(w_n4452_4[2]));
	jspl3 jspl3_w_n4452_16(.douta(w_n4452_16[0]),.doutb(w_n4452_16[1]),.doutc(w_n4452_16[2]),.din(w_n4452_5[0]));
	jspl3 jspl3_w_n4452_17(.douta(w_n4452_17[0]),.doutb(w_n4452_17[1]),.doutc(w_n4452_17[2]),.din(w_n4452_5[1]));
	jspl3 jspl3_w_n4452_18(.douta(w_n4452_18[0]),.doutb(w_n4452_18[1]),.doutc(w_n4452_18[2]),.din(w_n4452_5[2]));
	jspl3 jspl3_w_n4452_19(.douta(w_n4452_19[0]),.doutb(w_n4452_19[1]),.doutc(w_n4452_19[2]),.din(w_n4452_6[0]));
	jspl3 jspl3_w_n4452_20(.douta(w_n4452_20[0]),.doutb(w_n4452_20[1]),.doutc(w_n4452_20[2]),.din(w_n4452_6[1]));
	jspl3 jspl3_w_n4452_21(.douta(w_n4452_21[0]),.doutb(w_n4452_21[1]),.doutc(w_n4452_21[2]),.din(w_n4452_6[2]));
	jspl3 jspl3_w_n4452_22(.douta(w_n4452_22[0]),.doutb(w_n4452_22[1]),.doutc(w_n4452_22[2]),.din(w_n4452_7[0]));
	jspl3 jspl3_w_n4452_23(.douta(w_n4452_23[0]),.doutb(w_n4452_23[1]),.doutc(w_n4452_23[2]),.din(w_n4452_7[1]));
	jspl3 jspl3_w_n4452_24(.douta(w_n4452_24[0]),.doutb(w_n4452_24[1]),.doutc(w_n4452_24[2]),.din(w_n4452_7[2]));
	jspl3 jspl3_w_n4452_25(.douta(w_n4452_25[0]),.doutb(w_n4452_25[1]),.doutc(w_n4452_25[2]),.din(w_n4452_8[0]));
	jspl3 jspl3_w_n4452_26(.douta(w_n4452_26[0]),.doutb(w_n4452_26[1]),.doutc(w_n4452_26[2]),.din(w_n4452_8[1]));
	jspl3 jspl3_w_n4452_27(.douta(w_n4452_27[0]),.doutb(w_n4452_27[1]),.doutc(w_n4452_27[2]),.din(w_n4452_8[2]));
	jspl3 jspl3_w_n4452_28(.douta(w_n4452_28[0]),.doutb(w_n4452_28[1]),.doutc(w_n4452_28[2]),.din(w_n4452_9[0]));
	jspl3 jspl3_w_n4452_29(.douta(w_n4452_29[0]),.doutb(w_n4452_29[1]),.doutc(w_n4452_29[2]),.din(w_n4452_9[1]));
	jspl3 jspl3_w_n4452_30(.douta(w_n4452_30[0]),.doutb(w_n4452_30[1]),.doutc(w_n4452_30[2]),.din(w_n4452_9[2]));
	jspl3 jspl3_w_n4452_31(.douta(w_n4452_31[0]),.doutb(w_n4452_31[1]),.doutc(w_n4452_31[2]),.din(w_n4452_10[0]));
	jspl3 jspl3_w_n4452_32(.douta(w_n4452_32[0]),.doutb(w_n4452_32[1]),.doutc(w_n4452_32[2]),.din(w_n4452_10[1]));
	jspl3 jspl3_w_n4452_33(.douta(w_n4452_33[0]),.doutb(w_n4452_33[1]),.doutc(w_n4452_33[2]),.din(w_n4452_10[2]));
	jspl3 jspl3_w_n4452_34(.douta(w_n4452_34[0]),.doutb(w_n4452_34[1]),.doutc(w_n4452_34[2]),.din(w_n4452_11[0]));
	jspl3 jspl3_w_n4452_35(.douta(w_n4452_35[0]),.doutb(w_n4452_35[1]),.doutc(w_n4452_35[2]),.din(w_n4452_11[1]));
	jspl3 jspl3_w_n4452_36(.douta(w_n4452_36[0]),.doutb(w_n4452_36[1]),.doutc(w_n4452_36[2]),.din(w_n4452_11[2]));
	jspl3 jspl3_w_n4452_37(.douta(w_n4452_37[0]),.doutb(w_n4452_37[1]),.doutc(w_n4452_37[2]),.din(w_n4452_12[0]));
	jspl3 jspl3_w_n4452_38(.douta(w_n4452_38[0]),.doutb(w_n4452_38[1]),.doutc(w_n4452_38[2]),.din(w_n4452_12[1]));
	jspl3 jspl3_w_n4452_39(.douta(w_n4452_39[0]),.doutb(w_n4452_39[1]),.doutc(w_n4452_39[2]),.din(w_n4452_12[2]));
	jspl3 jspl3_w_n4452_40(.douta(w_n4452_40[0]),.doutb(w_n4452_40[1]),.doutc(w_n4452_40[2]),.din(w_n4452_13[0]));
	jspl3 jspl3_w_n4452_41(.douta(w_n4452_41[0]),.doutb(w_n4452_41[1]),.doutc(w_n4452_41[2]),.din(w_n4452_13[1]));
	jspl3 jspl3_w_n4452_42(.douta(w_n4452_42[0]),.doutb(w_n4452_42[1]),.doutc(w_n4452_42[2]),.din(w_n4452_13[2]));
	jspl3 jspl3_w_n4452_43(.douta(w_n4452_43[0]),.doutb(w_n4452_43[1]),.doutc(w_n4452_43[2]),.din(w_n4452_14[0]));
	jspl3 jspl3_w_n4452_44(.douta(w_n4452_44[0]),.doutb(w_n4452_44[1]),.doutc(w_n4452_44[2]),.din(w_n4452_14[1]));
	jspl3 jspl3_w_n4452_45(.douta(w_n4452_45[0]),.doutb(w_n4452_45[1]),.doutc(w_n4452_45[2]),.din(w_n4452_14[2]));
	jspl3 jspl3_w_n4452_46(.douta(w_n4452_46[0]),.doutb(w_n4452_46[1]),.doutc(w_n4452_46[2]),.din(w_n4452_15[0]));
	jspl3 jspl3_w_n4452_47(.douta(w_n4452_47[0]),.doutb(w_n4452_47[1]),.doutc(w_n4452_47[2]),.din(w_n4452_15[1]));
	jspl3 jspl3_w_n4452_48(.douta(w_n4452_48[0]),.doutb(w_n4452_48[1]),.doutc(w_n4452_48[2]),.din(w_n4452_15[2]));
	jspl3 jspl3_w_n4452_49(.douta(w_n4452_49[0]),.doutb(w_n4452_49[1]),.doutc(w_n4452_49[2]),.din(w_n4452_16[0]));
	jspl3 jspl3_w_n4452_50(.douta(w_n4452_50[0]),.doutb(w_n4452_50[1]),.doutc(w_n4452_50[2]),.din(w_n4452_16[1]));
	jspl3 jspl3_w_n4452_51(.douta(w_n4452_51[0]),.doutb(w_n4452_51[1]),.doutc(w_n4452_51[2]),.din(w_n4452_16[2]));
	jspl3 jspl3_w_n4452_52(.douta(w_n4452_52[0]),.doutb(w_n4452_52[1]),.doutc(w_n4452_52[2]),.din(w_n4452_17[0]));
	jspl3 jspl3_w_n4452_53(.douta(w_n4452_53[0]),.doutb(w_n4452_53[1]),.doutc(w_n4452_53[2]),.din(w_n4452_17[1]));
	jspl3 jspl3_w_n4452_54(.douta(w_n4452_54[0]),.doutb(w_n4452_54[1]),.doutc(w_n4452_54[2]),.din(w_n4452_17[2]));
	jspl3 jspl3_w_n4452_55(.douta(w_n4452_55[0]),.doutb(w_n4452_55[1]),.doutc(w_n4452_55[2]),.din(w_n4452_18[0]));
	jspl3 jspl3_w_n4452_56(.douta(w_n4452_56[0]),.doutb(w_n4452_56[1]),.doutc(w_n4452_56[2]),.din(w_n4452_18[1]));
	jspl3 jspl3_w_n4452_57(.douta(w_n4452_57[0]),.doutb(w_n4452_57[1]),.doutc(w_n4452_57[2]),.din(w_n4452_18[2]));
	jspl3 jspl3_w_n4452_58(.douta(w_n4452_58[0]),.doutb(w_n4452_58[1]),.doutc(w_n4452_58[2]),.din(w_n4452_19[0]));
	jspl3 jspl3_w_n4452_59(.douta(w_n4452_59[0]),.doutb(w_n4452_59[1]),.doutc(w_n4452_59[2]),.din(w_n4452_19[1]));
	jspl3 jspl3_w_n4452_60(.douta(w_n4452_60[0]),.doutb(w_n4452_60[1]),.doutc(w_n4452_60[2]),.din(w_n4452_19[2]));
	jspl3 jspl3_w_n4452_61(.douta(w_n4452_61[0]),.doutb(w_n4452_61[1]),.doutc(w_n4452_61[2]),.din(w_n4452_20[0]));
	jspl3 jspl3_w_n4452_62(.douta(w_n4452_62[0]),.doutb(w_n4452_62[1]),.doutc(w_n4452_62[2]),.din(w_n4452_20[1]));
	jspl jspl_w_n4452_63(.douta(w_n4452_63[0]),.doutb(w_n4452_63[1]),.din(w_n4452_20[2]));
endmodule

