/*

c499:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jdff: 477
	jand: 69
	jor: 2

Summary:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jdff: 477
	jand: 69
	jor: 2
*/

module c499(gclk, Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr, God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10, God11, God12, God13, God14, God15, God16, God17, God18, God19, God20, God21, God22, God23, God24, God25, God26, God27, God28, God29, God30, God31);
	input gclk;
	input Gid0;
	input Gid1;
	input Gid2;
	input Gid3;
	input Gid4;
	input Gid5;
	input Gid6;
	input Gid7;
	input Gid8;
	input Gid9;
	input Gid10;
	input Gid11;
	input Gid12;
	input Gid13;
	input Gid14;
	input Gid15;
	input Gid16;
	input Gid17;
	input Gid18;
	input Gid19;
	input Gid20;
	input Gid21;
	input Gid22;
	input Gid23;
	input Gid24;
	input Gid25;
	input Gid26;
	input Gid27;
	input Gid28;
	input Gid29;
	input Gid30;
	input Gid31;
	input Gic0;
	input Gic1;
	input Gic2;
	input Gic3;
	input Gic4;
	input Gic5;
	input Gic6;
	input Gic7;
	input Gr;
	output God0;
	output God1;
	output God2;
	output God3;
	output God4;
	output God5;
	output God6;
	output God7;
	output God8;
	output God9;
	output God10;
	output God11;
	output God12;
	output God13;
	output God14;
	output God15;
	output God16;
	output God17;
	output God18;
	output God19;
	output God20;
	output God21;
	output God22;
	output God23;
	output God24;
	output God25;
	output God26;
	output God27;
	output God28;
	output God29;
	output God30;
	output God31;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n180;
	wire n182;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n208;
	wire n210;
	wire n212;
	wire n214;
	wire n215;
	wire n217;
	wire n219;
	wire n221;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n236;
	wire n238;
	wire n240;
	wire n242;
	wire n243;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n257;
	wire n259;
	wire n261;
	wire n263;
	wire n264;
	wire n266;
	wire n268;
	wire n270;
	wire[2:0] w_Gid0_0;
	wire[2:0] w_Gid1_0;
	wire[2:0] w_Gid2_0;
	wire[2:0] w_Gid3_0;
	wire[2:0] w_Gid4_0;
	wire[2:0] w_Gid5_0;
	wire[2:0] w_Gid6_0;
	wire[2:0] w_Gid7_0;
	wire[2:0] w_Gid8_0;
	wire[2:0] w_Gid9_0;
	wire[2:0] w_Gid10_0;
	wire[2:0] w_Gid11_0;
	wire[2:0] w_Gid12_0;
	wire[2:0] w_Gid13_0;
	wire[2:0] w_Gid14_0;
	wire[2:0] w_Gid15_0;
	wire[2:0] w_Gid16_0;
	wire[2:0] w_Gid17_0;
	wire[2:0] w_Gid18_0;
	wire[2:0] w_Gid19_0;
	wire[2:0] w_Gid20_0;
	wire[2:0] w_Gid21_0;
	wire[2:0] w_Gid22_0;
	wire[2:0] w_Gid23_0;
	wire[2:0] w_Gid24_0;
	wire[2:0] w_Gid25_0;
	wire[2:0] w_Gid26_0;
	wire[2:0] w_Gid27_0;
	wire[2:0] w_Gid28_0;
	wire[2:0] w_Gid29_0;
	wire[2:0] w_Gid30_0;
	wire[2:0] w_Gid31_0;
	wire[2:0] w_Gr_0;
	wire[2:0] w_Gr_1;
	wire[2:0] w_Gr_2;
	wire[1:0] w_Gr_3;
	wire[1:0] w_n75_0;
	wire[1:0] w_n76_0;
	wire[1:0] w_n80_0;
	wire[1:0] w_n83_0;
	wire[1:0] w_n84_0;
	wire[2:0] w_n85_0;
	wire[2:0] w_n85_1;
	wire[1:0] w_n85_2;
	wire[1:0] w_n88_0;
	wire[1:0] w_n89_0;
	wire[1:0] w_n94_0;
	wire[1:0] w_n97_0;
	wire[1:0] w_n98_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n110_0;
	wire[2:0] w_n112_0;
	wire[2:0] w_n112_1;
	wire[2:0] w_n112_2;
	wire[1:0] w_n113_0;
	wire[1:0] w_n116_0;
	wire[1:0] w_n117_0;
	wire[2:0] w_n121_0;
	wire[2:0] w_n124_0;
	wire[1:0] w_n125_0;
	wire[2:0] w_n126_0;
	wire[2:0] w_n126_1;
	wire[1:0] w_n126_2;
	wire[1:0] w_n128_0;
	wire[1:0] w_n134_0;
	wire[1:0] w_n135_0;
	wire[1:0] w_n136_0;
	wire[1:0] w_n142_0;
	wire[1:0] w_n143_0;
	wire[2:0] w_n147_0;
	wire[2:0] w_n147_1;
	wire[1:0] w_n147_2;
	wire[2:0] w_n149_0;
	wire[2:0] w_n149_1;
	wire[1:0] w_n149_2;
	wire[1:0] w_n153_0;
	wire[1:0] w_n156_0;
	wire[2:0] w_n159_0;
	wire[2:0] w_n166_0;
	wire[2:0] w_n166_1;
	wire[2:0] w_n166_2;
	wire[1:0] w_n169_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n173_0;
	wire[1:0] w_n174_0;
	wire[1:0] w_n175_0;
	wire[2:0] w_n177_0;
	wire[1:0] w_n177_1;
	wire[2:0] w_n187_0;
	wire[2:0] w_n187_1;
	wire[1:0] w_n187_2;
	wire[1:0] w_n188_0;
	wire[1:0] w_n190_0;
	wire[2:0] w_n191_0;
	wire[1:0] w_n191_1;
	wire[1:0] w_n200_0;
	wire[2:0] w_n202_0;
	wire[2:0] w_n202_1;
	wire[1:0] w_n202_2;
	wire[1:0] w_n203_0;
	wire[2:0] w_n205_0;
	wire[1:0] w_n205_1;
	wire[2:0] w_n214_0;
	wire[1:0] w_n214_1;
	wire[1:0] w_n223_0;
	wire[1:0] w_n231_0;
	wire[1:0] w_n232_0;
	wire[2:0] w_n233_0;
	wire[1:0] w_n233_1;
	wire[1:0] w_n242_0;
	wire[2:0] w_n243_0;
	wire[1:0] w_n243_1;
	wire[1:0] w_n253_0;
	wire[2:0] w_n254_0;
	wire[1:0] w_n254_1;
	wire[2:0] w_n263_0;
	wire[1:0] w_n263_1;
	wire w_dff_A_HoWUHdQH2_0;
	wire w_dff_B_pAbBgdB52_2;
	wire w_dff_B_GMpZWws20_2;
	wire w_dff_A_8ZijYjOL7_1;
	wire w_dff_B_UJm8ovED1_2;
	wire w_dff_B_kwEaaIlM6_2;
	wire w_dff_B_Aagbht658_2;
	wire w_dff_B_NNXjPwoP5_2;
	wire w_dff_B_w91MFonu0_0;
	wire w_dff_A_YtGQicij1_0;
	wire w_dff_A_ckHqjUs57_0;
	wire w_dff_A_k11gxhEr1_0;
	wire w_dff_A_txyzGUW91_0;
	wire w_dff_A_UUr1NN2G1_0;
	wire w_dff_A_SkGcpYNV2_0;
	wire w_dff_A_KRqS4puO4_0;
	wire w_dff_A_YfLut0Hh9_0;
	wire w_dff_A_fa5kmyk58_0;
	wire w_dff_A_5aPM2m0H6_0;
	wire w_dff_A_cc2FcGqv5_0;
	wire w_dff_A_BZGLh76p3_0;
	wire w_dff_A_Nz3soHCj8_0;
	wire w_dff_A_x4VMgrds9_0;
	wire w_dff_A_JbhDJidZ3_0;
	wire w_dff_A_Yk1quGHS8_0;
	wire w_dff_A_jSEIuM0S2_0;
	wire w_dff_A_y93vSQD31_0;
	wire w_dff_A_dq7HSxkn7_0;
	wire w_dff_A_G3Odxsz12_0;
	wire w_dff_B_J5qPlMcc4_1;
	wire w_dff_B_HSrG6axq3_1;
	wire w_dff_B_aHXBSO2c5_1;
	wire w_dff_A_WjkkbW1A7_0;
	wire w_dff_A_Okz3N2ZI5_0;
	wire w_dff_A_QZzevMzZ2_0;
	wire w_dff_A_dm90QVCZ2_0;
	wire w_dff_A_GLdBpa8R2_0;
	wire w_dff_B_EIVXnNwD6_2;
	wire w_dff_B_DeFoqr9n1_2;
	wire w_dff_B_jyQNsKvf0_2;
	wire w_dff_B_ECkcM7Sk3_2;
	wire w_dff_A_zbWGbccO9_0;
	wire w_dff_A_H1bURtMk2_0;
	wire w_dff_A_sKlTtmZo9_0;
	wire w_dff_A_O2hrJ8Oi5_0;
	wire w_dff_A_kouesCZ51_0;
	wire w_dff_B_jD4msZKY8_1;
	wire w_dff_B_CrkLuT4L1_1;
	wire w_dff_B_skr2rCCy2_1;
	wire w_dff_A_LsGM724X9_1;
	wire w_dff_A_aKNrtzEE3_0;
	wire w_dff_A_gAl6sXE41_0;
	wire w_dff_A_CSdkc0uV9_0;
	wire w_dff_A_AESXkZ3g1_0;
	wire w_dff_A_1oHMNMIl0_0;
	wire w_dff_A_4zMwLGa54_0;
	wire w_dff_A_lzSRPRLW0_2;
	wire w_dff_A_kRLD7ASN1_2;
	wire w_dff_A_zsyRP6U56_2;
	wire w_dff_A_euOnKGV63_2;
	wire w_dff_A_oK3Rfrt93_2;
	wire w_dff_A_d3L3hxUC9_2;
	wire w_dff_A_EsOppI9A6_0;
	wire w_dff_A_OtUZ3OQg5_0;
	wire w_dff_A_h2hSAZqx3_0;
	wire w_dff_A_gsMY22nn1_0;
	wire w_dff_A_0ElUoHYA1_0;
	wire w_dff_A_NNcyoPb40_0;
	wire w_dff_A_1Q3AdVVT1_0;
	wire w_dff_A_NHKn0XM39_0;
	wire w_dff_A_ioDMRqFO1_2;
	wire w_dff_A_h1Sv8cbK3_2;
	wire w_dff_A_lKT3LCmM4_2;
	wire w_dff_A_tGFfRfQO9_2;
	wire w_dff_A_vJhGN7vr4_2;
	wire w_dff_A_1IGmGCdt3_2;
	wire w_dff_B_OGea3b1V6_0;
	wire w_dff_A_v5AgDqSn0_1;
	wire w_dff_A_o8GW8mLm4_0;
	wire w_dff_A_Y39bNc334_0;
	wire w_dff_A_gCHxkEGT6_0;
	wire w_dff_A_0FX5yOxr7_0;
	wire w_dff_A_fWHsbvL39_0;
	wire w_dff_A_VvhUkKYo0_0;
	wire w_dff_A_zYqpquXc1_2;
	wire w_dff_A_fvWKGZ906_2;
	wire w_dff_A_PTWxl2Bg8_2;
	wire w_dff_A_w7k5JWZQ5_2;
	wire w_dff_A_GLAz6XHV1_2;
	wire w_dff_A_yqkwcKb51_2;
	wire w_dff_A_lKVvOPZU8_0;
	wire w_dff_A_Zrr6ZSQM2_0;
	wire w_dff_A_EVBvp8uP4_0;
	wire w_dff_A_ocZJeKfG0_0;
	wire w_dff_A_S6SPzRxd2_0;
	wire w_dff_A_Zltb77XP4_0;
	wire w_dff_A_e9DOuGuZ2_0;
	wire w_dff_A_Mi6puyjn1_0;
	wire w_dff_A_ncOT31789_0;
	wire w_dff_A_6kCoJHCc9_0;
	wire w_dff_A_EDN1BP2P5_2;
	wire w_dff_A_YOnhxyEB8_2;
	wire w_dff_A_t0bRbQ4e2_2;
	wire w_dff_A_RsE4UdCg0_2;
	wire w_dff_A_wLh0IS6b7_2;
	wire w_dff_A_NlFUP3rV4_2;
	wire w_dff_B_xfF7qKG06_0;
	wire w_dff_A_27tCEe9p9_0;
	wire w_dff_A_0DJYsMlD9_0;
	wire w_dff_A_BTlMwhvN4_0;
	wire w_dff_A_MqcPDGpM3_0;
	wire w_dff_A_szVXKRdS1_0;
	wire w_dff_A_XUUVkTQw2_1;
	wire w_dff_A_4x0k3mbf3_0;
	wire w_dff_A_x1O8sHmc6_0;
	wire w_dff_A_syVzu0mB6_0;
	wire w_dff_A_HuCNUgV15_0;
	wire w_dff_A_HpnwQW0I7_0;
	wire w_dff_A_deQt634Y1_0;
	wire w_dff_A_XTMqNynd8_0;
	wire w_dff_A_HSpUMFuf5_0;
	wire w_dff_A_a8ovwaJa4_0;
	wire w_dff_A_FsZ928ee4_0;
	wire w_dff_A_SgK2oljL9_0;
	wire w_dff_A_Slrt1nby0_0;
	wire w_dff_A_1weuSl5B8_0;
	wire w_dff_A_2asTmUIh8_0;
	wire w_dff_A_BM23FvwM2_0;
	wire w_dff_A_2vsEVonw8_0;
	wire w_dff_A_UpPWbCxt4_0;
	wire w_dff_A_gUAHoXEa4_0;
	wire w_dff_A_RL22MX3t8_0;
	wire w_dff_A_RDPAxx727_0;
	wire w_dff_A_0dG4O0b87_0;
	wire w_dff_A_7qfItyga7_0;
	wire w_dff_A_YlGH6HEB1_0;
	wire w_dff_A_w9If26RQ8_0;
	wire w_dff_A_ixdvjmhe7_0;
	wire w_dff_A_xpHHIJ0p7_0;
	wire w_dff_A_w8I692aC8_0;
	wire w_dff_A_ThPsk3tD9_0;
	wire w_dff_A_HP0K8dfy3_0;
	wire w_dff_A_F2RObYci4_0;
	wire w_dff_A_T2khZzMp1_0;
	wire w_dff_A_6IxBHSti0_0;
	wire w_dff_A_xgpiTuYB9_0;
	wire w_dff_A_FvW3GEIA6_0;
	wire w_dff_A_pmZLmlXD6_0;
	wire w_dff_A_p0dDEl534_0;
	wire w_dff_A_rz776DlD4_0;
	wire w_dff_A_XVn4JwNj8_0;
	wire w_dff_A_66WhRsON5_0;
	wire w_dff_A_2Yd29BnD0_0;
	wire w_dff_A_h4E10oPH3_1;
	wire w_dff_A_cHjRnBxy3_0;
	wire w_dff_A_JRTUmYCW1_0;
	wire w_dff_A_ntJ5gssM9_0;
	wire w_dff_A_meMhRixP4_0;
	wire w_dff_A_A41J6o1b2_0;
	wire w_dff_A_U8Hfjj2e2_0;
	wire w_dff_A_L4KpYBWZ2_0;
	wire w_dff_A_xqOlH3Yn3_0;
	wire w_dff_A_23xFbOV76_0;
	wire w_dff_A_45nYmdsw5_0;
	wire w_dff_A_RzDX4wxU4_0;
	wire w_dff_A_0Q5O5aZM4_0;
	wire w_dff_A_p9R3FxQu2_0;
	wire w_dff_A_cFJWuGx49_0;
	wire w_dff_A_GIYOLG237_0;
	wire w_dff_A_5rg81iup9_0;
	wire w_dff_A_eddGRi5j7_0;
	wire w_dff_A_vXhZ7gUh3_0;
	wire w_dff_A_PdSI8fnx1_0;
	wire w_dff_A_mPGuB67I3_0;
	wire w_dff_A_RfshTlXF4_0;
	wire w_dff_A_4HkAsBd42_0;
	wire w_dff_A_F4QdNfe19_0;
	wire w_dff_A_oIdDMQgo5_0;
	wire w_dff_A_FBsyP8q70_0;
	wire w_dff_A_btI128zX7_0;
	wire w_dff_A_q2l4SC2z5_0;
	wire w_dff_A_zGCazSqR4_0;
	wire w_dff_A_e4PhpqOI8_0;
	wire w_dff_A_UzWUyWuH4_0;
	wire w_dff_A_sjsJuoN04_0;
	wire w_dff_A_suIrNB7M6_0;
	wire w_dff_A_yvqttXuw3_0;
	wire w_dff_A_xd2SLPAM3_0;
	wire w_dff_A_bsMIfAdG0_0;
	wire w_dff_A_vXBOCL5A2_0;
	wire w_dff_A_rx0CEOyP5_0;
	wire w_dff_A_70Je6q9c2_0;
	wire w_dff_A_WtRxzlij2_0;
	wire w_dff_A_R5CqIMM82_0;
	wire w_dff_B_7bfFOply5_2;
	wire w_dff_B_cCHm3leD5_2;
	wire w_dff_B_lMxa1oXZ0_2;
	wire w_dff_B_q2Ij04a04_2;
	wire w_dff_A_VOw69Q4S9_0;
	wire w_dff_A_PK6uusgM9_0;
	wire w_dff_A_fOvJW4xP6_0;
	wire w_dff_A_v320Hgdd9_0;
	wire w_dff_A_o65peZUF4_0;
	wire w_dff_A_pw6h5Ib81_0;
	wire w_dff_A_u5gmwgAq8_0;
	wire w_dff_A_9TD7mNXE9_0;
	wire w_dff_A_VPJegpDt5_0;
	wire w_dff_A_tn5P6gzj0_0;
	wire w_dff_A_VbyMVxYj9_0;
	wire w_dff_A_GsIAFlQd8_0;
	wire w_dff_A_Bwilk3af1_0;
	wire w_dff_A_QzTvfGdj4_0;
	wire w_dff_A_tlxPseM01_0;
	wire w_dff_A_1zdsX12Y0_0;
	wire w_dff_A_eElExFlk9_0;
	wire w_dff_A_UPxqfPJI7_0;
	wire w_dff_A_D31qGBF63_0;
	wire w_dff_A_QrUoxd2A3_0;
	wire w_dff_A_m45EXfcm5_0;
	wire w_dff_A_I0gkpmK81_0;
	wire w_dff_A_7uLpjd9s5_0;
	wire w_dff_A_h2uxgz751_0;
	wire w_dff_A_dQ76stEf8_0;
	wire w_dff_A_pufpSbk40_0;
	wire w_dff_A_jEOMZGKt5_0;
	wire w_dff_A_JXubLcg98_0;
	wire w_dff_A_5nbRMX5v0_0;
	wire w_dff_A_whgqRjwp1_0;
	wire w_dff_A_GdoRZXIG5_0;
	wire w_dff_A_8LCjIbj19_0;
	wire w_dff_A_FWM7JK3s7_0;
	wire w_dff_A_TC7oSpl93_0;
	wire w_dff_A_e1BCPvu42_0;
	wire w_dff_A_eU6Lhmnj2_0;
	wire w_dff_A_HhPt07mp3_0;
	wire w_dff_A_f6jCHpFM7_0;
	wire w_dff_A_g8vQeElE0_0;
	wire w_dff_A_vMrH8TvP3_0;
	wire w_dff_A_cASUW5hR5_0;
	wire w_dff_A_3RA6tENn7_0;
	wire w_dff_A_EXawvFXI8_0;
	wire w_dff_A_65aplbU78_0;
	wire w_dff_A_68BJbQ8D3_0;
	wire w_dff_A_Y33yLsSb7_0;
	wire w_dff_A_B5CPzabP4_0;
	wire w_dff_A_prlhLW9Z2_0;
	wire w_dff_A_PF7j2tx89_0;
	wire w_dff_A_Ajz5gCAU9_0;
	wire w_dff_A_3hvJBpol7_0;
	wire w_dff_A_2P9YjnMl8_0;
	wire w_dff_A_NaWxm0Vu2_0;
	wire w_dff_A_UbLBlLK47_0;
	wire w_dff_A_FvYcQYev2_0;
	wire w_dff_A_g3z3w5oC1_0;
	wire w_dff_A_RhQtjhXb3_0;
	wire w_dff_A_UiipUCVH4_0;
	wire w_dff_A_8K991h965_0;
	wire w_dff_A_l8AYu8lY4_0;
	wire w_dff_A_fDsKudNf5_0;
	wire w_dff_A_vcPrUY5d1_0;
	wire w_dff_A_dtvuA91o4_0;
	wire w_dff_A_xYnyUA9b2_0;
	wire w_dff_A_nJFnqXJF3_0;
	wire w_dff_A_ZHeeBaHR4_0;
	wire w_dff_A_ZqU9HZ8v1_0;
	wire w_dff_A_DtzoR74x6_0;
	wire w_dff_A_0KiXf2cX7_0;
	wire w_dff_A_0IcjlmqK9_0;
	wire w_dff_A_OXRPh0kW4_0;
	wire w_dff_A_6mAf3AwT7_0;
	wire w_dff_A_48fX9mcn2_0;
	wire w_dff_A_3osGbBNr1_0;
	wire w_dff_A_nQCWmlJu7_0;
	wire w_dff_A_Hp5DeOLV0_0;
	wire w_dff_A_8LkhMyKa0_0;
	wire w_dff_A_4qy07Ypo5_0;
	wire w_dff_A_x97rfs7l2_0;
	wire w_dff_A_h1OxO95z7_0;
	wire w_dff_A_7ZuYobcK0_0;
	wire w_dff_A_hTRPTVZH1_0;
	wire w_dff_A_qbgQ2jDN7_0;
	wire w_dff_A_swKGAntW1_0;
	wire w_dff_A_2LDJkh3t8_0;
	wire w_dff_A_zJfUTd4q8_0;
	wire w_dff_A_ZDrkqYjG0_0;
	wire w_dff_A_0vXoOyjT0_0;
	wire w_dff_A_5Q5qA0642_0;
	wire w_dff_A_gYVOYK0p1_0;
	wire w_dff_A_UJmpBvXi7_0;
	wire w_dff_A_uDsOVl0F8_0;
	wire w_dff_A_iODDi2CH9_0;
	wire w_dff_A_gwoAee4U9_0;
	wire w_dff_A_TvXjSViK8_0;
	wire w_dff_A_IKEsPeSf3_0;
	wire w_dff_A_8WEIMdgR7_0;
	wire w_dff_A_CLwDdsUQ3_0;
	wire w_dff_A_p84QDqHd2_0;
	wire w_dff_A_IGBZRrqz4_0;
	wire w_dff_A_zj45PG1S7_0;
	wire w_dff_A_6GUgtQJS9_0;
	wire w_dff_A_tUs3HHDq8_0;
	wire w_dff_A_7i76XiWq5_0;
	wire w_dff_A_JCF0EKvh4_0;
	wire w_dff_A_luKafPcj5_0;
	wire w_dff_A_YvK4cSR30_0;
	wire w_dff_A_3vm7JMe32_0;
	wire w_dff_A_OBmMmhu55_0;
	wire w_dff_A_EuTwiRAA3_0;
	wire w_dff_A_rLjbzQKE6_0;
	wire w_dff_A_e9BCc0k89_0;
	wire w_dff_A_041ZalXw9_0;
	wire w_dff_A_fHLJIFQ38_0;
	wire w_dff_A_LwhnlwNA6_0;
	wire w_dff_A_gUwHN94g7_0;
	wire w_dff_A_KgZ5YJTo9_0;
	wire w_dff_A_Trwj7LQB3_0;
	wire w_dff_A_I4GWRoe42_0;
	wire w_dff_A_7dXePNXv4_0;
	wire w_dff_A_ciMjUmTy3_0;
	wire w_dff_A_s2YLLYJL1_0;
	wire w_dff_A_LHlD12sB5_0;
	wire w_dff_A_XBz8Iay49_0;
	wire w_dff_A_XraUgurW5_0;
	wire w_dff_A_olOnVLQo1_0;
	wire w_dff_A_52hF7bX48_0;
	wire w_dff_A_wiKkNZ6w2_0;
	wire w_dff_A_cPxyNrLc5_0;
	wire w_dff_A_trgskhLC3_0;
	wire w_dff_A_nNMzKHqI9_0;
	wire w_dff_A_MNZtudzM7_0;
	wire w_dff_A_Emcxli7F3_0;
	wire w_dff_A_4qEya7Iu6_0;
	wire w_dff_A_QMle7d0n5_0;
	wire w_dff_A_Uask23rq9_0;
	wire w_dff_A_L0dnapZQ4_0;
	wire w_dff_A_8cZ2XvID8_0;
	wire w_dff_A_dnRLACyM0_0;
	wire w_dff_A_o1k0E09P9_0;
	wire w_dff_A_4azYrVDd9_0;
	wire w_dff_A_3VzZp6fV1_0;
	wire w_dff_A_Ib0LBkQ53_0;
	wire w_dff_A_QydXU8MJ2_0;
	wire w_dff_A_x29eqbbc9_0;
	wire w_dff_A_gt2eYnkQ7_0;
	wire w_dff_A_Nui8Siru6_0;
	wire w_dff_A_rF4NN6kG4_0;
	wire w_dff_A_UaHlL3YW6_0;
	wire w_dff_A_B3s3Xmxd5_0;
	wire w_dff_A_rpyOg9iQ7_0;
	wire w_dff_A_quShtIId7_0;
	wire w_dff_A_xKTCn2ip9_0;
	wire w_dff_A_Ob44XYIB0_0;
	wire w_dff_A_JbNBaWVt4_0;
	wire w_dff_A_UgT0i45a7_0;
	wire w_dff_A_Ox8FXqk35_0;
	wire w_dff_A_gyYCP9vq7_0;
	wire w_dff_A_ZxTT2OXD6_0;
	wire w_dff_A_eez2zmGH1_0;
	wire w_dff_A_buFgwA2A6_0;
	wire w_dff_A_kPOjCu7D2_0;
	wire w_dff_A_T4fA4E962_0;
	wire w_dff_A_zDinP9BW2_0;
	wire w_dff_A_RV9iZpna7_0;
	wire w_dff_A_48nMjq3h3_0;
	wire w_dff_A_zee0PFFx7_0;
	wire w_dff_A_ImYl7bbI2_0;
	wire w_dff_A_j95C3OIv4_0;
	wire w_dff_A_oELo6KbY4_0;
	wire w_dff_A_GQuxPzKt6_0;
	wire w_dff_A_LKbD6RPp6_0;
	wire w_dff_A_pWVRce4r7_0;
	wire w_dff_A_FEmzwO6L8_0;
	wire w_dff_A_nFNYR6Rh8_0;
	wire w_dff_A_htS3z7by4_0;
	wire w_dff_A_TWSLCyWV2_0;
	wire w_dff_A_1KYJRseF7_0;
	wire w_dff_A_Pg6Sjzua4_0;
	wire w_dff_A_5m77TeH39_0;
	wire w_dff_A_pjcVxXi56_0;
	wire w_dff_A_HhRBAEDp7_0;
	wire w_dff_A_5bnA5CB90_0;
	wire w_dff_A_RtkDc7Dv4_0;
	wire w_dff_A_yIuxIPZN8_0;
	wire w_dff_A_IoQM1IDB9_0;
	wire w_dff_A_U1vFxNb61_0;
	wire w_dff_A_EnUdaxB08_0;
	wire w_dff_A_7lphQtNi1_0;
	wire w_dff_A_s506qQm57_0;
	wire w_dff_A_5G4JXHHt5_0;
	wire w_dff_A_uDLRzEar5_0;
	wire w_dff_A_JIYmvVR86_0;
	wire w_dff_A_kaxjGrzs2_0;
	wire w_dff_A_RoU1uwMN6_0;
	wire w_dff_A_lgfvsrkH8_0;
	wire w_dff_A_LYdN8MiC6_0;
	wire w_dff_A_m54Sm2SY7_0;
	wire w_dff_A_0GLQNQEO1_0;
	wire w_dff_A_IrMCqxkP2_0;
	wire w_dff_A_slFS2xON7_0;
	wire w_dff_A_eoiM19aI5_0;
	wire w_dff_A_jQXMnGLa6_0;
	wire w_dff_A_xOWaKdHa1_0;
	wire w_dff_A_CFYOo6Dg7_0;
	wire w_dff_A_b0TOLugh7_0;
	wire w_dff_A_D7URHJsV8_0;
	wire w_dff_A_e0dDOrGk2_0;
	wire w_dff_A_z1dcoJah6_0;
	wire w_dff_A_eJ6E6ibW1_0;
	wire w_dff_A_0tpNe0sL6_0;
	wire w_dff_A_HEepittY7_0;
	wire w_dff_A_7MOUxzP32_0;
	wire w_dff_A_lZWHOGJ01_0;
	wire w_dff_A_AO9QGGjU0_0;
	wire w_dff_A_rlF4guPS3_0;
	wire w_dff_A_HDG8o1MW2_0;
	wire w_dff_A_itpsinfy8_0;
	wire w_dff_A_mWAiAKq28_0;
	wire w_dff_A_Nde5DTjx7_0;
	wire w_dff_A_j2Jl1zX12_0;
	wire w_dff_A_6EMXGX7K5_0;
	wire w_dff_A_gVxcNbrD3_0;
	wire w_dff_A_PCqWS4FX8_0;
	wire w_dff_A_2PhElid30_0;
	wire w_dff_A_02ACiawp3_0;
	wire w_dff_A_ZE2YkXj61_0;
	wire w_dff_A_QNDgQq9I7_0;
	wire w_dff_A_UG1DeCEJ9_0;
	wire w_dff_A_U9iWXrnT9_0;
	wire w_dff_A_7IrYAtEj3_0;
	wire w_dff_A_MvyTxmeJ9_0;
	wire w_dff_A_UW1KUhnE1_0;
	wire w_dff_A_5Xk5mWEQ3_0;
	wire w_dff_A_2ncx7ghg9_0;
	wire w_dff_A_kQDGFQS41_0;
	wire w_dff_A_DN2GL6VX9_0;
	wire w_dff_A_r0UfnC7k9_0;
	wire w_dff_A_VV47jh2h5_0;
	wire w_dff_A_7OG5vszE2_0;
	wire w_dff_A_89jrkGWO8_0;
	wire w_dff_A_KcPfHo4i8_0;
	wire w_dff_A_26dNHKoN0_0;
	wire w_dff_A_SIUIpMYO3_0;
	wire w_dff_A_EXZ40ExW8_0;
	wire w_dff_A_zjYQiali2_0;
	wire w_dff_A_PiNvl5Oa2_0;
	wire w_dff_A_PRPEmvZp8_0;
	wire w_dff_A_RwXCACcd3_0;
	wire w_dff_A_WCpZzk0x8_0;
	wire w_dff_A_b00r57cX9_0;
	wire w_dff_A_jrTa5pKo7_0;
	wire w_dff_A_fbe2HY1E3_0;
	wire w_dff_A_oPrjtPxO0_0;
	wire w_dff_A_Lhdn5QVK2_0;
	wire w_dff_A_Rnby4Qjf5_0;
	wire w_dff_A_DUEzQ0Zt6_0;
	wire w_dff_A_59tip4um6_0;
	wire w_dff_A_JYr03RyS0_0;
	wire w_dff_A_3YAnqSFD0_0;
	wire w_dff_A_ZPhOJqXE6_0;
	wire w_dff_A_PmGAFBZK7_0;
	wire w_dff_A_VBd96eJ74_0;
	wire w_dff_A_GTlv67Vm9_2;
	wire w_dff_A_GSZfjr7J0_2;
	wire w_dff_A_uQkLPNWZ8_2;
	wire w_dff_A_55Gbgj6p6_2;
	wire w_dff_A_B8wZr4MU3_2;
	wire w_dff_A_yRU2enKl6_2;
	wire w_dff_A_Q05eg1e32_2;
	wire w_dff_A_tI95YF7r3_2;
	wire w_dff_A_M8cCqJfp6_2;
	wire w_dff_A_TN9CdVrU9_2;
	wire w_dff_A_SdT464Q11_2;
	wire w_dff_A_lnT3lzl99_2;
	wire w_dff_A_7jbkq2NO0_2;
	wire w_dff_A_EIKtJcB52_2;
	wire w_dff_A_5MddvVjy9_2;
	wire w_dff_A_64k6T4eZ6_2;
	jxor g000(.dina(w_Gid12_0[2]),.dinb(w_Gid8_0[2]),.dout(n73),.clk(gclk));
	jxor g001(.dina(w_Gid4_0[2]),.dinb(w_Gid0_0[2]),.dout(n74),.clk(gclk));
	jxor g002(.dina(n74),.dinb(n73),.dout(n75),.clk(gclk));
	jand g003(.dina(w_Gr_3[1]),.dinb(Gic0),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_n76_0[1]),.dinb(w_n75_0[1]),.dout(n77),.clk(gclk));
	jxor g005(.dina(w_Gid19_0[2]),.dinb(w_Gid18_0[2]),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_Gid17_0[2]),.dinb(w_Gid16_0[2]),.dout(n79),.clk(gclk));
	jxor g007(.dina(n79),.dinb(n78),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_Gid23_0[2]),.dinb(w_Gid22_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(w_Gid21_0[2]),.dinb(w_Gid20_0[2]),.dout(n82),.clk(gclk));
	jxor g010(.dina(n82),.dinb(n81),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_n83_0[1]),.dinb(w_n80_0[1]),.dout(n84),.clk(gclk));
	jxor g012(.dina(w_n84_0[1]),.dinb(n77),.dout(n85),.clk(gclk));
	jxor g013(.dina(w_Gid31_0[2]),.dinb(w_Gid27_0[2]),.dout(n86),.clk(gclk));
	jxor g014(.dina(w_Gid23_0[1]),.dinb(w_Gid19_0[1]),.dout(n87),.clk(gclk));
	jxor g015(.dina(n87),.dinb(n86),.dout(n88),.clk(gclk));
	jand g016(.dina(w_Gr_3[0]),.dinb(Gic7),.dout(n89),.clk(gclk));
	jnot g017(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jxor g018(.dina(n90),.dinb(w_n88_0[1]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_Gid7_0[2]),.dinb(w_Gid6_0[2]),.dout(n92),.clk(gclk));
	jxor g020(.dina(w_Gid5_0[2]),.dinb(w_Gid4_0[1]),.dout(n93),.clk(gclk));
	jxor g021(.dina(n93),.dinb(n92),.dout(n94),.clk(gclk));
	jxor g022(.dina(w_Gid15_0[2]),.dinb(w_Gid14_0[2]),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_Gid13_0[2]),.dinb(w_Gid12_0[1]),.dout(n96),.clk(gclk));
	jxor g024(.dina(n96),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_n97_0[1]),.dinb(w_n94_0[1]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_n98_0[1]),.dinb(n91),.dout(n99),.clk(gclk));
	jxor g027(.dina(w_Gid30_0[2]),.dinb(w_Gid26_0[2]),.dout(n100),.clk(gclk));
	jxor g028(.dina(w_Gid22_0[1]),.dinb(w_Gid18_0[1]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n100),.dout(n102),.clk(gclk));
	jand g030(.dina(w_Gr_2[2]),.dinb(Gic6),.dout(n103),.clk(gclk));
	jxor g031(.dina(w_dff_B_OGea3b1V6_0),.dinb(n102),.dout(n104),.clk(gclk));
	jxor g032(.dina(w_Gid3_0[2]),.dinb(w_Gid2_0[2]),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_Gid1_0[2]),.dinb(w_Gid0_0[1]),.dout(n106),.clk(gclk));
	jxor g034(.dina(n106),.dinb(n105),.dout(n107),.clk(gclk));
	jxor g035(.dina(w_Gid11_0[2]),.dinb(w_Gid10_0[2]),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_Gid9_0[2]),.dinb(w_Gid8_0[1]),.dout(n109),.clk(gclk));
	jxor g037(.dina(n109),.dinb(n108),.dout(n110),.clk(gclk));
	jxor g038(.dina(w_n110_0[1]),.dinb(w_n107_0[1]),.dout(n111),.clk(gclk));
	jxor g039(.dina(n111),.dinb(n104),.dout(n112),.clk(gclk));
	jand g040(.dina(w_n112_2[2]),.dinb(w_n99_0[1]),.dout(n113),.clk(gclk));
	jxor g041(.dina(w_Gid13_0[1]),.dinb(w_Gid9_0[1]),.dout(n114),.clk(gclk));
	jxor g042(.dina(w_Gid5_0[1]),.dinb(w_Gid1_0[1]),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jand g044(.dina(w_Gr_2[1]),.dinb(Gic1),.dout(n117),.clk(gclk));
	jxor g045(.dina(w_n117_0[1]),.dinb(w_n116_0[1]),.dout(n118),.clk(gclk));
	jxor g046(.dina(w_Gid31_0[1]),.dinb(w_Gid30_0[1]),.dout(n119),.clk(gclk));
	jxor g047(.dina(w_Gid29_0[2]),.dinb(w_Gid28_0[2]),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(n119),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_Gid27_0[1]),.dinb(w_Gid26_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_Gid25_0[2]),.dinb(w_Gid24_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(w_n124_0[2]),.dinb(w_n121_0[2]),.dout(n125),.clk(gclk));
	jxor g053(.dina(w_n125_0[1]),.dinb(n118),.dout(n126),.clk(gclk));
	jxor g054(.dina(w_n126_2[1]),.dinb(w_n85_2[1]),.dout(n127),.clk(gclk));
	jand g055(.dina(w_Gr_2[0]),.dinb(Gic3),.dout(n128),.clk(gclk));
	jnot g056(.din(w_n128_0[1]),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(w_n121_0[1]),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_Gid15_0[1]),.dinb(w_Gid11_0[1]),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_Gid7_0[1]),.dinb(w_Gid3_0[1]),.dout(n132),.clk(gclk));
	jxor g060(.dina(n132),.dinb(n131),.dout(n133),.clk(gclk));
	jxor g061(.dina(n133),.dinb(w_n83_0[0]),.dout(n134),.clk(gclk));
	jxor g062(.dina(w_n134_0[1]),.dinb(n130),.dout(n135),.clk(gclk));
	jand g063(.dina(w_Gr_1[2]),.dinb(Gic2),.dout(n136),.clk(gclk));
	jnot g064(.din(w_n136_0[1]),.dout(n137),.clk(gclk));
	jxor g065(.dina(n137),.dinb(w_n124_0[1]),.dout(n138),.clk(gclk));
	jxor g066(.dina(w_Gid14_0[1]),.dinb(w_Gid10_0[1]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_Gid6_0[1]),.dinb(w_Gid2_0[1]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g069(.dina(n141),.dinb(w_n80_0[0]),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_n142_0[1]),.dinb(n138),.dout(n143),.clk(gclk));
	jand g071(.dina(w_n143_0[1]),.dinb(w_n135_0[1]),.dout(n144),.clk(gclk));
	jand g072(.dina(n144),.dinb(n127),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_n128_0[0]),.dinb(w_n121_0[0]),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_n134_0[0]),.dinb(n146),.dout(n147),.clk(gclk));
	jxor g075(.dina(w_n136_0[0]),.dinb(w_n124_0[0]),.dout(n148),.clk(gclk));
	jxor g076(.dina(w_n142_0[0]),.dinb(n148),.dout(n149),.clk(gclk));
	jxor g077(.dina(w_n149_2[1]),.dinb(w_n147_2[1]),.dout(n150),.clk(gclk));
	jnot g078(.din(w_n76_0[0]),.dout(n151),.clk(gclk));
	jxor g079(.dina(n151),.dinb(w_n75_0[0]),.dout(n152),.clk(gclk));
	jxor g080(.dina(w_n84_0[0]),.dinb(n152),.dout(n153),.clk(gclk));
	jnot g081(.din(w_n117_0[0]),.dout(n154),.clk(gclk));
	jxor g082(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_n125_0[0]),.dinb(n155),.dout(n156),.clk(gclk));
	jand g084(.dina(w_n156_0[1]),.dinb(w_n153_0[1]),.dout(n157),.clk(gclk));
	jand g085(.dina(n157),.dinb(n150),.dout(n158),.clk(gclk));
	jor g086(.dina(n158),.dinb(n145),.dout(n159),.clk(gclk));
	jxor g087(.dina(w_Gid28_0[1]),.dinb(w_Gid24_0[1]),.dout(n160),.clk(gclk));
	jxor g088(.dina(w_Gid20_0[1]),.dinb(w_Gid16_0[1]),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(n160),.dout(n162),.clk(gclk));
	jand g090(.dina(w_Gr_1[1]),.dinb(Gic4),.dout(n163),.clk(gclk));
	jxor g091(.dina(w_dff_B_xfF7qKG06_0),.dinb(n162),.dout(n164),.clk(gclk));
	jxor g092(.dina(w_n107_0[0]),.dinb(w_n94_0[0]),.dout(n165),.clk(gclk));
	jxor g093(.dina(n165),.dinb(n164),.dout(n166),.clk(gclk));
	jxor g094(.dina(w_Gid29_0[1]),.dinb(w_Gid25_0[1]),.dout(n167),.clk(gclk));
	jxor g095(.dina(w_Gid21_0[1]),.dinb(w_Gid17_0[1]),.dout(n168),.clk(gclk));
	jxor g096(.dina(n168),.dinb(n167),.dout(n169),.clk(gclk));
	jand g097(.dina(w_Gr_1[0]),.dinb(Gic5),.dout(n170),.clk(gclk));
	jnot g098(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jxor g099(.dina(n171),.dinb(w_n169_0[1]),.dout(n172),.clk(gclk));
	jxor g100(.dina(w_n110_0[0]),.dinb(w_n97_0[0]),.dout(n173),.clk(gclk));
	jxor g101(.dina(w_n173_0[1]),.dinb(n172),.dout(n174),.clk(gclk));
	jand g102(.dina(w_n174_0[1]),.dinb(w_n166_2[2]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_0[1]),.dinb(w_n159_0[2]),.dout(n176),.clk(gclk));
	jand g104(.dina(n176),.dinb(w_n113_0[1]),.dout(n177),.clk(gclk));
	jand g105(.dina(w_n177_1[1]),.dinb(w_n85_2[0]),.dout(n178),.clk(gclk));
	jxor g106(.dina(n178),.dinb(w_Gid0_0[0]),.dout(w_dff_A_GTlv67Vm9_2),.clk(gclk));
	jand g107(.dina(w_n177_1[0]),.dinb(w_n126_2[0]),.dout(n180),.clk(gclk));
	jxor g108(.dina(n180),.dinb(w_Gid1_0[0]),.dout(w_dff_A_GSZfjr7J0_2),.clk(gclk));
	jand g109(.dina(w_n177_0[2]),.dinb(w_n149_2[0]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_Gid2_0[0]),.dout(w_dff_A_uQkLPNWZ8_2),.clk(gclk));
	jand g111(.dina(w_n177_0[1]),.dinb(w_n147_2[0]),.dout(n184),.clk(gclk));
	jxor g112(.dina(n184),.dinb(w_Gid3_0[0]),.dout(w_dff_A_55Gbgj6p6_2),.clk(gclk));
	jxor g113(.dina(w_n89_0[0]),.dinb(w_n88_0[0]),.dout(n186),.clk(gclk));
	jxor g114(.dina(w_n98_0[0]),.dinb(n186),.dout(n187),.clk(gclk));
	jnot g115(.din(w_n112_2[1]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n188_0[1]),.dinb(w_n187_2[1]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_dff_B_w91MFonu0_0),.dinb(w_n159_0[1]),.dout(n190),.clk(gclk));
	jand g118(.dina(w_n190_0[1]),.dinb(w_n175_0[0]),.dout(n191),.clk(gclk));
	jand g119(.dina(w_n191_1[1]),.dinb(w_n85_1[2]),.dout(n192),.clk(gclk));
	jxor g120(.dina(n192),.dinb(w_Gid4_0[0]),.dout(w_dff_A_B8wZr4MU3_2),.clk(gclk));
	jand g121(.dina(w_n191_1[0]),.dinb(w_n126_1[2]),.dout(n194),.clk(gclk));
	jxor g122(.dina(n194),.dinb(w_Gid5_0[0]),.dout(w_dff_A_yRU2enKl6_2),.clk(gclk));
	jand g123(.dina(w_n191_0[2]),.dinb(w_n149_1[2]),.dout(n196),.clk(gclk));
	jxor g124(.dina(n196),.dinb(w_Gid6_0[0]),.dout(w_dff_A_Q05eg1e32_2),.clk(gclk));
	jand g125(.dina(w_n191_0[1]),.dinb(w_n147_1[2]),.dout(n198),.clk(gclk));
	jxor g126(.dina(n198),.dinb(w_Gid7_0[0]),.dout(w_dff_A_tI95YF7r3_2),.clk(gclk));
	jnot g127(.din(w_n166_2[1]),.dout(n200),.clk(gclk));
	jxor g128(.dina(w_n170_0[0]),.dinb(w_n169_0[0]),.dout(n201),.clk(gclk));
	jxor g129(.dina(w_n173_0[0]),.dinb(n201),.dout(n202),.clk(gclk));
	jand g130(.dina(w_n202_2[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jand g131(.dina(w_n159_0[0]),.dinb(w_n113_0[0]),.dout(n204),.clk(gclk));
	jand g132(.dina(n204),.dinb(w_n203_0[1]),.dout(n205),.clk(gclk));
	jand g133(.dina(w_n205_1[1]),.dinb(w_n85_1[1]),.dout(n206),.clk(gclk));
	jxor g134(.dina(n206),.dinb(w_Gid8_0[0]),.dout(w_dff_A_M8cCqJfp6_2),.clk(gclk));
	jand g135(.dina(w_n205_1[0]),.dinb(w_n126_1[1]),.dout(n208),.clk(gclk));
	jxor g136(.dina(n208),.dinb(w_Gid9_0[0]),.dout(w_dff_A_TN9CdVrU9_2),.clk(gclk));
	jand g137(.dina(w_n205_0[2]),.dinb(w_n149_1[1]),.dout(n210),.clk(gclk));
	jxor g138(.dina(n210),.dinb(w_Gid10_0[0]),.dout(w_dff_A_SdT464Q11_2),.clk(gclk));
	jand g139(.dina(w_n205_0[1]),.dinb(w_n147_1[1]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_Gid11_0[0]),.dout(w_dff_A_lnT3lzl99_2),.clk(gclk));
	jand g141(.dina(w_n203_0[0]),.dinb(w_n190_0[0]),.dout(n214),.clk(gclk));
	jand g142(.dina(w_n214_1[1]),.dinb(w_n85_1[0]),.dout(n215),.clk(gclk));
	jxor g143(.dina(n215),.dinb(w_Gid12_0[0]),.dout(w_dff_A_7jbkq2NO0_2),.clk(gclk));
	jand g144(.dina(w_n214_1[0]),.dinb(w_n126_1[0]),.dout(n217),.clk(gclk));
	jxor g145(.dina(n217),.dinb(w_Gid13_0[0]),.dout(w_dff_A_EIKtJcB52_2),.clk(gclk));
	jand g146(.dina(w_n214_0[2]),.dinb(w_n149_1[0]),.dout(n219),.clk(gclk));
	jxor g147(.dina(n219),.dinb(w_Gid14_0[0]),.dout(w_dff_A_5MddvVjy9_2),.clk(gclk));
	jand g148(.dina(w_n214_0[1]),.dinb(w_n147_1[0]),.dout(n221),.clk(gclk));
	jxor g149(.dina(n221),.dinb(w_Gid15_0[0]),.dout(w_dff_A_64k6T4eZ6_2),.clk(gclk));
	jand g150(.dina(w_n149_0[2]),.dinb(w_n135_0[0]),.dout(n223),.clk(gclk));
	jand g151(.dina(w_n156_0[0]),.dinb(w_n85_0[2]),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n112_2[0]),.dinb(w_n187_2[0]),.dout(n225),.clk(gclk));
	jand g153(.dina(n225),.dinb(w_n174_0[0]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(w_n200_0[0]),.dout(n227),.clk(gclk));
	jxor g155(.dina(w_n202_2[0]),.dinb(w_n166_2[0]),.dout(n228),.clk(gclk));
	jand g156(.dina(n228),.dinb(w_n99_0[0]),.dout(n229),.clk(gclk));
	jand g157(.dina(n229),.dinb(w_n188_0[0]),.dout(n230),.clk(gclk));
	jor g158(.dina(n230),.dinb(n227),.dout(n231),.clk(gclk));
	jand g159(.dina(w_n231_0[1]),.dinb(w_dff_B_aHXBSO2c5_1),.dout(n232),.clk(gclk));
	jand g160(.dina(w_n232_0[1]),.dinb(w_n223_0[1]),.dout(n233),.clk(gclk));
	jand g161(.dina(w_n233_1[1]),.dinb(w_n166_1[2]),.dout(n234),.clk(gclk));
	jxor g162(.dina(n234),.dinb(w_Gid16_0[0]),.dout(God16),.clk(gclk));
	jand g163(.dina(w_n233_1[0]),.dinb(w_n202_1[2]),.dout(n236),.clk(gclk));
	jxor g164(.dina(n236),.dinb(w_Gid17_0[0]),.dout(God17),.clk(gclk));
	jand g165(.dina(w_n233_0[2]),.dinb(w_n112_1[2]),.dout(n238),.clk(gclk));
	jxor g166(.dina(n238),.dinb(w_Gid18_0[0]),.dout(God18),.clk(gclk));
	jand g167(.dina(w_n233_0[1]),.dinb(w_n187_1[2]),.dout(n240),.clk(gclk));
	jxor g168(.dina(n240),.dinb(w_Gid19_0[0]),.dout(God19),.clk(gclk));
	jand g169(.dina(w_n143_0[0]),.dinb(w_n147_0[2]),.dout(n242),.clk(gclk));
	jand g170(.dina(w_n232_0[0]),.dinb(w_n242_0[1]),.dout(n243),.clk(gclk));
	jand g171(.dina(w_n243_1[1]),.dinb(w_n166_1[1]),.dout(n244),.clk(gclk));
	jxor g172(.dina(n244),.dinb(w_Gid20_0[0]),.dout(God20),.clk(gclk));
	jand g173(.dina(w_n243_1[0]),.dinb(w_n202_1[1]),.dout(n246),.clk(gclk));
	jxor g174(.dina(n246),.dinb(w_Gid21_0[0]),.dout(God21),.clk(gclk));
	jand g175(.dina(w_n243_0[2]),.dinb(w_n112_1[1]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_Gid22_0[0]),.dout(God22),.clk(gclk));
	jand g177(.dina(w_n243_0[1]),.dinb(w_n187_1[1]),.dout(n250),.clk(gclk));
	jxor g178(.dina(n250),.dinb(w_Gid23_0[0]),.dout(God23),.clk(gclk));
	jand g179(.dina(w_n126_0[2]),.dinb(w_n153_0[0]),.dout(n252),.clk(gclk));
	jand g180(.dina(w_n231_0[0]),.dinb(w_dff_B_skr2rCCy2_1),.dout(n253),.clk(gclk));
	jand g181(.dina(w_n253_0[1]),.dinb(w_n223_0[0]),.dout(n254),.clk(gclk));
	jand g182(.dina(w_n254_1[1]),.dinb(w_n166_1[0]),.dout(n255),.clk(gclk));
	jxor g183(.dina(n255),.dinb(w_Gid24_0[0]),.dout(God24),.clk(gclk));
	jand g184(.dina(w_n254_1[0]),.dinb(w_n202_1[0]),.dout(n257),.clk(gclk));
	jxor g185(.dina(n257),.dinb(w_Gid25_0[0]),.dout(God25),.clk(gclk));
	jand g186(.dina(w_n254_0[2]),.dinb(w_n112_1[0]),.dout(n259),.clk(gclk));
	jxor g187(.dina(n259),.dinb(w_Gid26_0[0]),.dout(God26),.clk(gclk));
	jand g188(.dina(w_n254_0[1]),.dinb(w_n187_1[0]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_Gid27_0[0]),.dout(God27),.clk(gclk));
	jand g190(.dina(w_n253_0[0]),.dinb(w_n242_0[0]),.dout(n263),.clk(gclk));
	jand g191(.dina(w_n263_1[1]),.dinb(w_n166_0[2]),.dout(n264),.clk(gclk));
	jxor g192(.dina(n264),.dinb(w_Gid28_0[0]),.dout(God28),.clk(gclk));
	jand g193(.dina(w_n263_1[0]),.dinb(w_n202_0[2]),.dout(n266),.clk(gclk));
	jxor g194(.dina(n266),.dinb(w_Gid29_0[0]),.dout(God29),.clk(gclk));
	jand g195(.dina(w_n263_0[2]),.dinb(w_n112_0[2]),.dout(n268),.clk(gclk));
	jxor g196(.dina(n268),.dinb(w_Gid30_0[0]),.dout(God30),.clk(gclk));
	jand g197(.dina(w_n263_0[1]),.dinb(w_n187_0[2]),.dout(n270),.clk(gclk));
	jxor g198(.dina(n270),.dinb(w_Gid31_0[0]),.dout(God31),.clk(gclk));
	jspl3 jspl3_w_Gid0_0(.douta(w_dff_A_mPGuB67I3_0),.doutb(w_Gid0_0[1]),.doutc(w_Gid0_0[2]),.din(Gid0));
	jspl3 jspl3_w_Gid1_0(.douta(w_dff_A_RDPAxx727_0),.doutb(w_Gid1_0[1]),.doutc(w_Gid1_0[2]),.din(Gid1));
	jspl3 jspl3_w_Gid2_0(.douta(w_dff_A_QrUoxd2A3_0),.doutb(w_Gid2_0[1]),.doutc(w_Gid2_0[2]),.din(Gid2));
	jspl3 jspl3_w_Gid3_0(.douta(w_dff_A_Ob44XYIB0_0),.doutb(w_Gid3_0[1]),.doutc(w_Gid3_0[2]),.din(Gid3));
	jspl3 jspl3_w_Gid4_0(.douta(w_dff_A_45nYmdsw5_0),.doutb(w_Gid4_0[1]),.doutc(w_Gid4_0[2]),.din(Gid4));
	jspl3 jspl3_w_Gid5_0(.douta(w_dff_A_FsZ928ee4_0),.doutb(w_Gid5_0[1]),.doutc(w_Gid5_0[2]),.din(Gid5));
	jspl3 jspl3_w_Gid6_0(.douta(w_dff_A_tn5P6gzj0_0),.doutb(w_Gid6_0[1]),.doutc(w_Gid6_0[2]),.din(Gid6));
	jspl3 jspl3_w_Gid7_0(.douta(w_dff_A_QydXU8MJ2_0),.doutb(w_Gid7_0[1]),.doutc(w_Gid7_0[2]),.din(Gid7));
	jspl3 jspl3_w_Gid8_0(.douta(w_dff_A_R5CqIMM82_0),.doutb(w_Gid8_0[1]),.doutc(w_Gid8_0[2]),.din(Gid8));
	jspl3 jspl3_w_Gid9_0(.douta(w_dff_A_2Yd29BnD0_0),.doutb(w_Gid9_0[1]),.doutc(w_Gid9_0[2]),.din(Gid9));
	jspl3 jspl3_w_Gid10_0(.douta(w_dff_A_vMrH8TvP3_0),.doutb(w_Gid10_0[1]),.doutc(w_Gid10_0[2]),.din(Gid10));
	jspl3 jspl3_w_Gid11_0(.douta(w_dff_A_FEmzwO6L8_0),.doutb(w_Gid11_0[1]),.doutc(w_Gid11_0[2]),.din(Gid11));
	jspl3 jspl3_w_Gid12_0(.douta(w_dff_A_UzWUyWuH4_0),.doutb(w_Gid12_0[1]),.doutc(w_Gid12_0[2]),.din(Gid12));
	jspl3 jspl3_w_Gid13_0(.douta(w_dff_A_F2RObYci4_0),.doutb(w_Gid13_0[1]),.doutc(w_Gid13_0[2]),.din(Gid13));
	jspl3 jspl3_w_Gid14_0(.douta(w_dff_A_whgqRjwp1_0),.doutb(w_Gid14_0[1]),.doutc(w_Gid14_0[2]),.din(Gid14));
	jspl3 jspl3_w_Gid15_0(.douta(w_dff_A_zDinP9BW2_0),.doutb(w_Gid15_0[1]),.doutc(w_Gid15_0[2]),.din(Gid15));
	jspl3 jspl3_w_Gid16_0(.douta(w_dff_A_vcPrUY5d1_0),.doutb(w_Gid16_0[1]),.doutc(w_Gid16_0[2]),.din(Gid16));
	jspl3 jspl3_w_Gid17_0(.douta(w_dff_A_3hvJBpol7_0),.doutb(w_Gid17_0[1]),.doutc(w_Gid17_0[2]),.din(Gid17));
	jspl3 jspl3_w_Gid18_0(.douta(w_dff_A_swKGAntW1_0),.doutb(w_Gid18_0[1]),.doutc(w_Gid18_0[2]),.din(Gid18));
	jspl3 jspl3_w_Gid19_0(.douta(w_dff_A_48fX9mcn2_0),.doutb(w_Gid19_0[1]),.doutc(w_Gid19_0[2]),.din(Gid19));
	jspl3 jspl3_w_Gid20_0(.douta(w_dff_A_lgfvsrkH8_0),.doutb(w_Gid20_0[1]),.doutc(w_Gid20_0[2]),.din(Gid20));
	jspl3 jspl3_w_Gid21_0(.douta(w_dff_A_yIuxIPZN8_0),.doutb(w_Gid21_0[1]),.doutc(w_Gid21_0[2]),.din(Gid21));
	jspl3 jspl3_w_Gid22_0(.douta(w_dff_A_itpsinfy8_0),.doutb(w_Gid22_0[1]),.doutc(w_Gid22_0[2]),.din(Gid22));
	jspl3 jspl3_w_Gid23_0(.douta(w_dff_A_D7URHJsV8_0),.doutb(w_Gid23_0[1]),.doutc(w_Gid23_0[2]),.din(Gid23));
	jspl3 jspl3_w_Gid24_0(.douta(w_dff_A_YvK4cSR30_0),.doutb(w_Gid24_0[1]),.doutc(w_Gid24_0[2]),.din(Gid24));
	jspl3 jspl3_w_Gid25_0(.douta(w_dff_A_IKEsPeSf3_0),.doutb(w_Gid25_0[1]),.doutc(w_Gid25_0[2]),.din(Gid25));
	jspl3 jspl3_w_Gid26_0(.douta(w_dff_A_cPxyNrLc5_0),.doutb(w_Gid26_0[1]),.doutc(w_Gid26_0[2]),.din(Gid26));
	jspl3 jspl3_w_Gid27_0(.douta(w_dff_A_Trwj7LQB3_0),.doutb(w_Gid27_0[1]),.doutc(w_Gid27_0[2]),.din(Gid27));
	jspl3 jspl3_w_Gid28_0(.douta(w_dff_A_89jrkGWO8_0),.doutb(w_Gid28_0[1]),.doutc(w_Gid28_0[2]),.din(Gid28));
	jspl3 jspl3_w_Gid29_0(.douta(w_dff_A_U9iWXrnT9_0),.doutb(w_Gid29_0[1]),.doutc(w_Gid29_0[2]),.din(Gid29));
	jspl3 jspl3_w_Gid30_0(.douta(w_dff_A_VBd96eJ74_0),.doutb(w_Gid30_0[1]),.doutc(w_Gid30_0[2]),.din(Gid30));
	jspl3 jspl3_w_Gid31_0(.douta(w_dff_A_jrTa5pKo7_0),.doutb(w_Gid31_0[1]),.doutc(w_Gid31_0[2]),.din(Gid31));
	jspl3 jspl3_w_Gr_0(.douta(w_Gr_0[0]),.doutb(w_Gr_0[1]),.doutc(w_Gr_0[2]),.din(Gr));
	jspl3 jspl3_w_Gr_1(.douta(w_Gr_1[0]),.doutb(w_Gr_1[1]),.doutc(w_Gr_1[2]),.din(w_Gr_0[0]));
	jspl3 jspl3_w_Gr_2(.douta(w_Gr_2[0]),.doutb(w_Gr_2[1]),.doutc(w_Gr_2[2]),.din(w_Gr_0[1]));
	jspl jspl_w_Gr_3(.douta(w_Gr_3[0]),.doutb(w_Gr_3[1]),.din(w_Gr_0[2]));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_dff_A_h4E10oPH3_1),.din(n76));
	jspl jspl_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_GLdBpa8R2_0),.doutb(w_n85_0[1]),.doutc(w_n85_0[2]),.din(n85));
	jspl3 jspl3_w_n85_1(.douta(w_n85_1[0]),.doutb(w_n85_1[1]),.doutc(w_n85_1[2]),.din(w_n85_0[0]));
	jspl jspl_w_n85_2(.douta(w_dff_A_G3Odxsz12_0),.doutb(w_n85_2[1]),.din(w_n85_0[1]));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n89_0(.douta(w_dff_A_lKVvOPZU8_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_dff_A_EsOppI9A6_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_NHKn0XM39_0),.doutb(w_n112_0[1]),.doutc(w_dff_A_1IGmGCdt3_2),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_dff_A_8ZijYjOL7_1),.din(w_dff_B_kwEaaIlM6_2));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.din(n116));
	jspl jspl_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_XUUVkTQw2_1),.din(n117));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.doutc(w_n124_0[2]),.din(n124));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_szVXKRdS1_0),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl3 jspl3_w_n126_1(.douta(w_n126_1[0]),.doutb(w_n126_1[1]),.doutc(w_n126_1[2]),.din(w_n126_0[0]));
	jspl jspl_w_n126_2(.douta(w_dff_A_JbhDJidZ3_0),.doutb(w_n126_2[1]),.din(w_n126_0[1]));
	jspl jspl_w_n128_0(.douta(w_dff_A_mWAiAKq28_0),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n134_0(.douta(w_n134_0[0]),.doutb(w_n134_0[1]),.din(n134));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n136_0(.douta(w_dff_A_2LDJkh3t8_0),.doutb(w_n136_0[1]),.din(n136));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl3 jspl3_w_n147_0(.douta(w_dff_A_4qEya7Iu6_0),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n147_1(.douta(w_n147_1[0]),.doutb(w_n147_1[1]),.doutc(w_n147_1[2]),.din(w_n147_0[0]));
	jspl jspl_w_n147_2(.douta(w_dff_A_5aPM2m0H6_0),.doutb(w_n147_2[1]),.din(w_n147_0[1]));
	jspl3 jspl3_w_n149_0(.douta(w_dff_A_kouesCZ51_0),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_n149_1[1]),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_UUr1NN2G1_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl jspl_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.din(n153));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl3 jspl3_w_n166_0(.douta(w_dff_A_6kCoJHCc9_0),.doutb(w_n166_0[1]),.doutc(w_dff_A_NlFUP3rV4_2),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.doutc(w_n166_1[2]),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_n166_2[2]),.din(w_n166_0[1]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_dff_A_EVBvp8uP4_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl jspl_w_n174_0(.douta(w_dff_A_Zrr6ZSQM2_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_dff_A_HoWUHdQH2_0),.doutb(w_n175_0[1]),.din(w_dff_B_GMpZWws20_2));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl jspl_w_n177_1(.douta(w_n177_1[0]),.doutb(w_n177_1[1]),.din(w_n177_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_dff_A_VvhUkKYo0_0),.doutb(w_n187_0[1]),.doutc(w_dff_A_yqkwcKb51_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_n187_1[0]),.doutb(w_n187_1[1]),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n187_2(.douta(w_n187_2[0]),.doutb(w_dff_A_v5AgDqSn0_1),.din(w_n187_0[1]));
	jspl jspl_w_n188_0(.douta(w_dff_A_OtUZ3OQg5_0),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n191_1(.douta(w_n191_1[0]),.doutb(w_n191_1[1]),.din(w_n191_0[0]));
	jspl jspl_w_n200_0(.douta(w_dff_A_ocZJeKfG0_0),.doutb(w_n200_0[1]),.din(n200));
	jspl3 jspl3_w_n202_0(.douta(w_dff_A_4zMwLGa54_0),.doutb(w_n202_0[1]),.doutc(w_dff_A_d3L3hxUC9_2),.din(n202));
	jspl3 jspl3_w_n202_1(.douta(w_n202_1[0]),.doutb(w_n202_1[1]),.doutc(w_n202_1[2]),.din(w_n202_0[0]));
	jspl jspl_w_n202_2(.douta(w_n202_2[0]),.doutb(w_dff_A_LsGM724X9_1),.din(w_n202_0[1]));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(w_dff_B_NNXjPwoP5_2));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(n205));
	jspl jspl_w_n205_1(.douta(w_n205_1[0]),.doutb(w_n205_1[1]),.din(w_n205_0[0]));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl jspl_w_n214_1(.douta(w_n214_1[0]),.doutb(w_n214_1[1]),.din(w_n214_0[0]));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.din(w_dff_B_ECkcM7Sk3_2));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(w_dff_B_q2Ij04a04_2));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n243_1(.douta(w_n243_1[0]),.doutb(w_n243_1[1]),.din(w_n243_0[0]));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.doutc(w_n263_0[2]),.din(n263));
	jspl jspl_w_n263_1(.douta(w_n263_1[0]),.doutb(w_n263_1[1]),.din(w_n263_0[0]));
	jdff dff_A_HoWUHdQH2_0(.dout(w_n175_0[0]),.din(w_dff_A_HoWUHdQH2_0),.clk(gclk));
	jdff dff_B_pAbBgdB52_2(.din(n175),.dout(w_dff_B_pAbBgdB52_2),.clk(gclk));
	jdff dff_B_GMpZWws20_2(.din(w_dff_B_pAbBgdB52_2),.dout(w_dff_B_GMpZWws20_2),.clk(gclk));
	jdff dff_A_8ZijYjOL7_1(.dout(w_n113_0[1]),.din(w_dff_A_8ZijYjOL7_1),.clk(gclk));
	jdff dff_B_UJm8ovED1_2(.din(n113),.dout(w_dff_B_UJm8ovED1_2),.clk(gclk));
	jdff dff_B_kwEaaIlM6_2(.din(w_dff_B_UJm8ovED1_2),.dout(w_dff_B_kwEaaIlM6_2),.clk(gclk));
	jdff dff_B_Aagbht658_2(.din(n203),.dout(w_dff_B_Aagbht658_2),.clk(gclk));
	jdff dff_B_NNXjPwoP5_2(.din(w_dff_B_Aagbht658_2),.dout(w_dff_B_NNXjPwoP5_2),.clk(gclk));
	jdff dff_B_w91MFonu0_0(.din(n189),.dout(w_dff_B_w91MFonu0_0),.clk(gclk));
	jdff dff_A_YtGQicij1_0(.dout(w_n149_2[0]),.din(w_dff_A_YtGQicij1_0),.clk(gclk));
	jdff dff_A_ckHqjUs57_0(.dout(w_dff_A_YtGQicij1_0),.din(w_dff_A_ckHqjUs57_0),.clk(gclk));
	jdff dff_A_k11gxhEr1_0(.dout(w_dff_A_ckHqjUs57_0),.din(w_dff_A_k11gxhEr1_0),.clk(gclk));
	jdff dff_A_txyzGUW91_0(.dout(w_dff_A_k11gxhEr1_0),.din(w_dff_A_txyzGUW91_0),.clk(gclk));
	jdff dff_A_UUr1NN2G1_0(.dout(w_dff_A_txyzGUW91_0),.din(w_dff_A_UUr1NN2G1_0),.clk(gclk));
	jdff dff_A_SkGcpYNV2_0(.dout(w_n147_2[0]),.din(w_dff_A_SkGcpYNV2_0),.clk(gclk));
	jdff dff_A_KRqS4puO4_0(.dout(w_dff_A_SkGcpYNV2_0),.din(w_dff_A_KRqS4puO4_0),.clk(gclk));
	jdff dff_A_YfLut0Hh9_0(.dout(w_dff_A_KRqS4puO4_0),.din(w_dff_A_YfLut0Hh9_0),.clk(gclk));
	jdff dff_A_fa5kmyk58_0(.dout(w_dff_A_YfLut0Hh9_0),.din(w_dff_A_fa5kmyk58_0),.clk(gclk));
	jdff dff_A_5aPM2m0H6_0(.dout(w_dff_A_fa5kmyk58_0),.din(w_dff_A_5aPM2m0H6_0),.clk(gclk));
	jdff dff_A_cc2FcGqv5_0(.dout(w_n126_2[0]),.din(w_dff_A_cc2FcGqv5_0),.clk(gclk));
	jdff dff_A_BZGLh76p3_0(.dout(w_dff_A_cc2FcGqv5_0),.din(w_dff_A_BZGLh76p3_0),.clk(gclk));
	jdff dff_A_Nz3soHCj8_0(.dout(w_dff_A_BZGLh76p3_0),.din(w_dff_A_Nz3soHCj8_0),.clk(gclk));
	jdff dff_A_x4VMgrds9_0(.dout(w_dff_A_Nz3soHCj8_0),.din(w_dff_A_x4VMgrds9_0),.clk(gclk));
	jdff dff_A_JbhDJidZ3_0(.dout(w_dff_A_x4VMgrds9_0),.din(w_dff_A_JbhDJidZ3_0),.clk(gclk));
	jdff dff_A_Yk1quGHS8_0(.dout(w_n85_2[0]),.din(w_dff_A_Yk1quGHS8_0),.clk(gclk));
	jdff dff_A_jSEIuM0S2_0(.dout(w_dff_A_Yk1quGHS8_0),.din(w_dff_A_jSEIuM0S2_0),.clk(gclk));
	jdff dff_A_y93vSQD31_0(.dout(w_dff_A_jSEIuM0S2_0),.din(w_dff_A_y93vSQD31_0),.clk(gclk));
	jdff dff_A_dq7HSxkn7_0(.dout(w_dff_A_y93vSQD31_0),.din(w_dff_A_dq7HSxkn7_0),.clk(gclk));
	jdff dff_A_G3Odxsz12_0(.dout(w_dff_A_dq7HSxkn7_0),.din(w_dff_A_G3Odxsz12_0),.clk(gclk));
	jdff dff_B_J5qPlMcc4_1(.din(n224),.dout(w_dff_B_J5qPlMcc4_1),.clk(gclk));
	jdff dff_B_HSrG6axq3_1(.din(w_dff_B_J5qPlMcc4_1),.dout(w_dff_B_HSrG6axq3_1),.clk(gclk));
	jdff dff_B_aHXBSO2c5_1(.din(w_dff_B_HSrG6axq3_1),.dout(w_dff_B_aHXBSO2c5_1),.clk(gclk));
	jdff dff_A_WjkkbW1A7_0(.dout(w_n85_0[0]),.din(w_dff_A_WjkkbW1A7_0),.clk(gclk));
	jdff dff_A_Okz3N2ZI5_0(.dout(w_dff_A_WjkkbW1A7_0),.din(w_dff_A_Okz3N2ZI5_0),.clk(gclk));
	jdff dff_A_QZzevMzZ2_0(.dout(w_dff_A_Okz3N2ZI5_0),.din(w_dff_A_QZzevMzZ2_0),.clk(gclk));
	jdff dff_A_dm90QVCZ2_0(.dout(w_dff_A_QZzevMzZ2_0),.din(w_dff_A_dm90QVCZ2_0),.clk(gclk));
	jdff dff_A_GLdBpa8R2_0(.dout(w_dff_A_dm90QVCZ2_0),.din(w_dff_A_GLdBpa8R2_0),.clk(gclk));
	jdff dff_B_EIVXnNwD6_2(.din(n223),.dout(w_dff_B_EIVXnNwD6_2),.clk(gclk));
	jdff dff_B_DeFoqr9n1_2(.din(w_dff_B_EIVXnNwD6_2),.dout(w_dff_B_DeFoqr9n1_2),.clk(gclk));
	jdff dff_B_jyQNsKvf0_2(.din(w_dff_B_DeFoqr9n1_2),.dout(w_dff_B_jyQNsKvf0_2),.clk(gclk));
	jdff dff_B_ECkcM7Sk3_2(.din(w_dff_B_jyQNsKvf0_2),.dout(w_dff_B_ECkcM7Sk3_2),.clk(gclk));
	jdff dff_A_zbWGbccO9_0(.dout(w_n149_0[0]),.din(w_dff_A_zbWGbccO9_0),.clk(gclk));
	jdff dff_A_H1bURtMk2_0(.dout(w_dff_A_zbWGbccO9_0),.din(w_dff_A_H1bURtMk2_0),.clk(gclk));
	jdff dff_A_sKlTtmZo9_0(.dout(w_dff_A_H1bURtMk2_0),.din(w_dff_A_sKlTtmZo9_0),.clk(gclk));
	jdff dff_A_O2hrJ8Oi5_0(.dout(w_dff_A_sKlTtmZo9_0),.din(w_dff_A_O2hrJ8Oi5_0),.clk(gclk));
	jdff dff_A_kouesCZ51_0(.dout(w_dff_A_O2hrJ8Oi5_0),.din(w_dff_A_kouesCZ51_0),.clk(gclk));
	jdff dff_B_jD4msZKY8_1(.din(n252),.dout(w_dff_B_jD4msZKY8_1),.clk(gclk));
	jdff dff_B_CrkLuT4L1_1(.din(w_dff_B_jD4msZKY8_1),.dout(w_dff_B_CrkLuT4L1_1),.clk(gclk));
	jdff dff_B_skr2rCCy2_1(.din(w_dff_B_CrkLuT4L1_1),.dout(w_dff_B_skr2rCCy2_1),.clk(gclk));
	jdff dff_A_LsGM724X9_1(.dout(w_n202_2[1]),.din(w_dff_A_LsGM724X9_1),.clk(gclk));
	jdff dff_A_aKNrtzEE3_0(.dout(w_n202_0[0]),.din(w_dff_A_aKNrtzEE3_0),.clk(gclk));
	jdff dff_A_gAl6sXE41_0(.dout(w_dff_A_aKNrtzEE3_0),.din(w_dff_A_gAl6sXE41_0),.clk(gclk));
	jdff dff_A_CSdkc0uV9_0(.dout(w_dff_A_gAl6sXE41_0),.din(w_dff_A_CSdkc0uV9_0),.clk(gclk));
	jdff dff_A_AESXkZ3g1_0(.dout(w_dff_A_CSdkc0uV9_0),.din(w_dff_A_AESXkZ3g1_0),.clk(gclk));
	jdff dff_A_1oHMNMIl0_0(.dout(w_dff_A_AESXkZ3g1_0),.din(w_dff_A_1oHMNMIl0_0),.clk(gclk));
	jdff dff_A_4zMwLGa54_0(.dout(w_dff_A_1oHMNMIl0_0),.din(w_dff_A_4zMwLGa54_0),.clk(gclk));
	jdff dff_A_lzSRPRLW0_2(.dout(w_n202_0[2]),.din(w_dff_A_lzSRPRLW0_2),.clk(gclk));
	jdff dff_A_kRLD7ASN1_2(.dout(w_dff_A_lzSRPRLW0_2),.din(w_dff_A_kRLD7ASN1_2),.clk(gclk));
	jdff dff_A_zsyRP6U56_2(.dout(w_dff_A_kRLD7ASN1_2),.din(w_dff_A_zsyRP6U56_2),.clk(gclk));
	jdff dff_A_euOnKGV63_2(.dout(w_dff_A_zsyRP6U56_2),.din(w_dff_A_euOnKGV63_2),.clk(gclk));
	jdff dff_A_oK3Rfrt93_2(.dout(w_dff_A_euOnKGV63_2),.din(w_dff_A_oK3Rfrt93_2),.clk(gclk));
	jdff dff_A_d3L3hxUC9_2(.dout(w_dff_A_oK3Rfrt93_2),.din(w_dff_A_d3L3hxUC9_2),.clk(gclk));
	jdff dff_A_EsOppI9A6_0(.dout(w_n99_0[0]),.din(w_dff_A_EsOppI9A6_0),.clk(gclk));
	jdff dff_A_OtUZ3OQg5_0(.dout(w_n188_0[0]),.din(w_dff_A_OtUZ3OQg5_0),.clk(gclk));
	jdff dff_A_h2hSAZqx3_0(.dout(w_n112_0[0]),.din(w_dff_A_h2hSAZqx3_0),.clk(gclk));
	jdff dff_A_gsMY22nn1_0(.dout(w_dff_A_h2hSAZqx3_0),.din(w_dff_A_gsMY22nn1_0),.clk(gclk));
	jdff dff_A_0ElUoHYA1_0(.dout(w_dff_A_gsMY22nn1_0),.din(w_dff_A_0ElUoHYA1_0),.clk(gclk));
	jdff dff_A_NNcyoPb40_0(.dout(w_dff_A_0ElUoHYA1_0),.din(w_dff_A_NNcyoPb40_0),.clk(gclk));
	jdff dff_A_1Q3AdVVT1_0(.dout(w_dff_A_NNcyoPb40_0),.din(w_dff_A_1Q3AdVVT1_0),.clk(gclk));
	jdff dff_A_NHKn0XM39_0(.dout(w_dff_A_1Q3AdVVT1_0),.din(w_dff_A_NHKn0XM39_0),.clk(gclk));
	jdff dff_A_ioDMRqFO1_2(.dout(w_n112_0[2]),.din(w_dff_A_ioDMRqFO1_2),.clk(gclk));
	jdff dff_A_h1Sv8cbK3_2(.dout(w_dff_A_ioDMRqFO1_2),.din(w_dff_A_h1Sv8cbK3_2),.clk(gclk));
	jdff dff_A_lKT3LCmM4_2(.dout(w_dff_A_h1Sv8cbK3_2),.din(w_dff_A_lKT3LCmM4_2),.clk(gclk));
	jdff dff_A_tGFfRfQO9_2(.dout(w_dff_A_lKT3LCmM4_2),.din(w_dff_A_tGFfRfQO9_2),.clk(gclk));
	jdff dff_A_vJhGN7vr4_2(.dout(w_dff_A_tGFfRfQO9_2),.din(w_dff_A_vJhGN7vr4_2),.clk(gclk));
	jdff dff_A_1IGmGCdt3_2(.dout(w_dff_A_vJhGN7vr4_2),.din(w_dff_A_1IGmGCdt3_2),.clk(gclk));
	jdff dff_B_OGea3b1V6_0(.din(n103),.dout(w_dff_B_OGea3b1V6_0),.clk(gclk));
	jdff dff_A_v5AgDqSn0_1(.dout(w_n187_2[1]),.din(w_dff_A_v5AgDqSn0_1),.clk(gclk));
	jdff dff_A_o8GW8mLm4_0(.dout(w_n187_0[0]),.din(w_dff_A_o8GW8mLm4_0),.clk(gclk));
	jdff dff_A_Y39bNc334_0(.dout(w_dff_A_o8GW8mLm4_0),.din(w_dff_A_Y39bNc334_0),.clk(gclk));
	jdff dff_A_gCHxkEGT6_0(.dout(w_dff_A_Y39bNc334_0),.din(w_dff_A_gCHxkEGT6_0),.clk(gclk));
	jdff dff_A_0FX5yOxr7_0(.dout(w_dff_A_gCHxkEGT6_0),.din(w_dff_A_0FX5yOxr7_0),.clk(gclk));
	jdff dff_A_fWHsbvL39_0(.dout(w_dff_A_0FX5yOxr7_0),.din(w_dff_A_fWHsbvL39_0),.clk(gclk));
	jdff dff_A_VvhUkKYo0_0(.dout(w_dff_A_fWHsbvL39_0),.din(w_dff_A_VvhUkKYo0_0),.clk(gclk));
	jdff dff_A_zYqpquXc1_2(.dout(w_n187_0[2]),.din(w_dff_A_zYqpquXc1_2),.clk(gclk));
	jdff dff_A_fvWKGZ906_2(.dout(w_dff_A_zYqpquXc1_2),.din(w_dff_A_fvWKGZ906_2),.clk(gclk));
	jdff dff_A_PTWxl2Bg8_2(.dout(w_dff_A_fvWKGZ906_2),.din(w_dff_A_PTWxl2Bg8_2),.clk(gclk));
	jdff dff_A_w7k5JWZQ5_2(.dout(w_dff_A_PTWxl2Bg8_2),.din(w_dff_A_w7k5JWZQ5_2),.clk(gclk));
	jdff dff_A_GLAz6XHV1_2(.dout(w_dff_A_w7k5JWZQ5_2),.din(w_dff_A_GLAz6XHV1_2),.clk(gclk));
	jdff dff_A_yqkwcKb51_2(.dout(w_dff_A_GLAz6XHV1_2),.din(w_dff_A_yqkwcKb51_2),.clk(gclk));
	jdff dff_A_lKVvOPZU8_0(.dout(w_n89_0[0]),.din(w_dff_A_lKVvOPZU8_0),.clk(gclk));
	jdff dff_A_Zrr6ZSQM2_0(.dout(w_n174_0[0]),.din(w_dff_A_Zrr6ZSQM2_0),.clk(gclk));
	jdff dff_A_EVBvp8uP4_0(.dout(w_n170_0[0]),.din(w_dff_A_EVBvp8uP4_0),.clk(gclk));
	jdff dff_A_ocZJeKfG0_0(.dout(w_n200_0[0]),.din(w_dff_A_ocZJeKfG0_0),.clk(gclk));
	jdff dff_A_S6SPzRxd2_0(.dout(w_n166_0[0]),.din(w_dff_A_S6SPzRxd2_0),.clk(gclk));
	jdff dff_A_Zltb77XP4_0(.dout(w_dff_A_S6SPzRxd2_0),.din(w_dff_A_Zltb77XP4_0),.clk(gclk));
	jdff dff_A_e9DOuGuZ2_0(.dout(w_dff_A_Zltb77XP4_0),.din(w_dff_A_e9DOuGuZ2_0),.clk(gclk));
	jdff dff_A_Mi6puyjn1_0(.dout(w_dff_A_e9DOuGuZ2_0),.din(w_dff_A_Mi6puyjn1_0),.clk(gclk));
	jdff dff_A_ncOT31789_0(.dout(w_dff_A_Mi6puyjn1_0),.din(w_dff_A_ncOT31789_0),.clk(gclk));
	jdff dff_A_6kCoJHCc9_0(.dout(w_dff_A_ncOT31789_0),.din(w_dff_A_6kCoJHCc9_0),.clk(gclk));
	jdff dff_A_EDN1BP2P5_2(.dout(w_n166_0[2]),.din(w_dff_A_EDN1BP2P5_2),.clk(gclk));
	jdff dff_A_YOnhxyEB8_2(.dout(w_dff_A_EDN1BP2P5_2),.din(w_dff_A_YOnhxyEB8_2),.clk(gclk));
	jdff dff_A_t0bRbQ4e2_2(.dout(w_dff_A_YOnhxyEB8_2),.din(w_dff_A_t0bRbQ4e2_2),.clk(gclk));
	jdff dff_A_RsE4UdCg0_2(.dout(w_dff_A_t0bRbQ4e2_2),.din(w_dff_A_RsE4UdCg0_2),.clk(gclk));
	jdff dff_A_wLh0IS6b7_2(.dout(w_dff_A_RsE4UdCg0_2),.din(w_dff_A_wLh0IS6b7_2),.clk(gclk));
	jdff dff_A_NlFUP3rV4_2(.dout(w_dff_A_wLh0IS6b7_2),.din(w_dff_A_NlFUP3rV4_2),.clk(gclk));
	jdff dff_B_xfF7qKG06_0(.din(n163),.dout(w_dff_B_xfF7qKG06_0),.clk(gclk));
	jdff dff_A_27tCEe9p9_0(.dout(w_n126_0[0]),.din(w_dff_A_27tCEe9p9_0),.clk(gclk));
	jdff dff_A_0DJYsMlD9_0(.dout(w_dff_A_27tCEe9p9_0),.din(w_dff_A_0DJYsMlD9_0),.clk(gclk));
	jdff dff_A_BTlMwhvN4_0(.dout(w_dff_A_0DJYsMlD9_0),.din(w_dff_A_BTlMwhvN4_0),.clk(gclk));
	jdff dff_A_MqcPDGpM3_0(.dout(w_dff_A_BTlMwhvN4_0),.din(w_dff_A_MqcPDGpM3_0),.clk(gclk));
	jdff dff_A_szVXKRdS1_0(.dout(w_dff_A_MqcPDGpM3_0),.din(w_dff_A_szVXKRdS1_0),.clk(gclk));
	jdff dff_A_XUUVkTQw2_1(.dout(w_n117_0[1]),.din(w_dff_A_XUUVkTQw2_1),.clk(gclk));
	jdff dff_A_4x0k3mbf3_0(.dout(w_Gid5_0[0]),.din(w_dff_A_4x0k3mbf3_0),.clk(gclk));
	jdff dff_A_x1O8sHmc6_0(.dout(w_dff_A_4x0k3mbf3_0),.din(w_dff_A_x1O8sHmc6_0),.clk(gclk));
	jdff dff_A_syVzu0mB6_0(.dout(w_dff_A_x1O8sHmc6_0),.din(w_dff_A_syVzu0mB6_0),.clk(gclk));
	jdff dff_A_HuCNUgV15_0(.dout(w_dff_A_syVzu0mB6_0),.din(w_dff_A_HuCNUgV15_0),.clk(gclk));
	jdff dff_A_HpnwQW0I7_0(.dout(w_dff_A_HuCNUgV15_0),.din(w_dff_A_HpnwQW0I7_0),.clk(gclk));
	jdff dff_A_deQt634Y1_0(.dout(w_dff_A_HpnwQW0I7_0),.din(w_dff_A_deQt634Y1_0),.clk(gclk));
	jdff dff_A_XTMqNynd8_0(.dout(w_dff_A_deQt634Y1_0),.din(w_dff_A_XTMqNynd8_0),.clk(gclk));
	jdff dff_A_HSpUMFuf5_0(.dout(w_dff_A_XTMqNynd8_0),.din(w_dff_A_HSpUMFuf5_0),.clk(gclk));
	jdff dff_A_a8ovwaJa4_0(.dout(w_dff_A_HSpUMFuf5_0),.din(w_dff_A_a8ovwaJa4_0),.clk(gclk));
	jdff dff_A_FsZ928ee4_0(.dout(w_dff_A_a8ovwaJa4_0),.din(w_dff_A_FsZ928ee4_0),.clk(gclk));
	jdff dff_A_SgK2oljL9_0(.dout(w_Gid1_0[0]),.din(w_dff_A_SgK2oljL9_0),.clk(gclk));
	jdff dff_A_Slrt1nby0_0(.dout(w_dff_A_SgK2oljL9_0),.din(w_dff_A_Slrt1nby0_0),.clk(gclk));
	jdff dff_A_1weuSl5B8_0(.dout(w_dff_A_Slrt1nby0_0),.din(w_dff_A_1weuSl5B8_0),.clk(gclk));
	jdff dff_A_2asTmUIh8_0(.dout(w_dff_A_1weuSl5B8_0),.din(w_dff_A_2asTmUIh8_0),.clk(gclk));
	jdff dff_A_BM23FvwM2_0(.dout(w_dff_A_2asTmUIh8_0),.din(w_dff_A_BM23FvwM2_0),.clk(gclk));
	jdff dff_A_2vsEVonw8_0(.dout(w_dff_A_BM23FvwM2_0),.din(w_dff_A_2vsEVonw8_0),.clk(gclk));
	jdff dff_A_UpPWbCxt4_0(.dout(w_dff_A_2vsEVonw8_0),.din(w_dff_A_UpPWbCxt4_0),.clk(gclk));
	jdff dff_A_gUAHoXEa4_0(.dout(w_dff_A_UpPWbCxt4_0),.din(w_dff_A_gUAHoXEa4_0),.clk(gclk));
	jdff dff_A_RL22MX3t8_0(.dout(w_dff_A_gUAHoXEa4_0),.din(w_dff_A_RL22MX3t8_0),.clk(gclk));
	jdff dff_A_RDPAxx727_0(.dout(w_dff_A_RL22MX3t8_0),.din(w_dff_A_RDPAxx727_0),.clk(gclk));
	jdff dff_A_0dG4O0b87_0(.dout(w_Gid13_0[0]),.din(w_dff_A_0dG4O0b87_0),.clk(gclk));
	jdff dff_A_7qfItyga7_0(.dout(w_dff_A_0dG4O0b87_0),.din(w_dff_A_7qfItyga7_0),.clk(gclk));
	jdff dff_A_YlGH6HEB1_0(.dout(w_dff_A_7qfItyga7_0),.din(w_dff_A_YlGH6HEB1_0),.clk(gclk));
	jdff dff_A_w9If26RQ8_0(.dout(w_dff_A_YlGH6HEB1_0),.din(w_dff_A_w9If26RQ8_0),.clk(gclk));
	jdff dff_A_ixdvjmhe7_0(.dout(w_dff_A_w9If26RQ8_0),.din(w_dff_A_ixdvjmhe7_0),.clk(gclk));
	jdff dff_A_xpHHIJ0p7_0(.dout(w_dff_A_ixdvjmhe7_0),.din(w_dff_A_xpHHIJ0p7_0),.clk(gclk));
	jdff dff_A_w8I692aC8_0(.dout(w_dff_A_xpHHIJ0p7_0),.din(w_dff_A_w8I692aC8_0),.clk(gclk));
	jdff dff_A_ThPsk3tD9_0(.dout(w_dff_A_w8I692aC8_0),.din(w_dff_A_ThPsk3tD9_0),.clk(gclk));
	jdff dff_A_HP0K8dfy3_0(.dout(w_dff_A_ThPsk3tD9_0),.din(w_dff_A_HP0K8dfy3_0),.clk(gclk));
	jdff dff_A_F2RObYci4_0(.dout(w_dff_A_HP0K8dfy3_0),.din(w_dff_A_F2RObYci4_0),.clk(gclk));
	jdff dff_A_T2khZzMp1_0(.dout(w_Gid9_0[0]),.din(w_dff_A_T2khZzMp1_0),.clk(gclk));
	jdff dff_A_6IxBHSti0_0(.dout(w_dff_A_T2khZzMp1_0),.din(w_dff_A_6IxBHSti0_0),.clk(gclk));
	jdff dff_A_xgpiTuYB9_0(.dout(w_dff_A_6IxBHSti0_0),.din(w_dff_A_xgpiTuYB9_0),.clk(gclk));
	jdff dff_A_FvW3GEIA6_0(.dout(w_dff_A_xgpiTuYB9_0),.din(w_dff_A_FvW3GEIA6_0),.clk(gclk));
	jdff dff_A_pmZLmlXD6_0(.dout(w_dff_A_FvW3GEIA6_0),.din(w_dff_A_pmZLmlXD6_0),.clk(gclk));
	jdff dff_A_p0dDEl534_0(.dout(w_dff_A_pmZLmlXD6_0),.din(w_dff_A_p0dDEl534_0),.clk(gclk));
	jdff dff_A_rz776DlD4_0(.dout(w_dff_A_p0dDEl534_0),.din(w_dff_A_rz776DlD4_0),.clk(gclk));
	jdff dff_A_XVn4JwNj8_0(.dout(w_dff_A_rz776DlD4_0),.din(w_dff_A_XVn4JwNj8_0),.clk(gclk));
	jdff dff_A_66WhRsON5_0(.dout(w_dff_A_XVn4JwNj8_0),.din(w_dff_A_66WhRsON5_0),.clk(gclk));
	jdff dff_A_2Yd29BnD0_0(.dout(w_dff_A_66WhRsON5_0),.din(w_dff_A_2Yd29BnD0_0),.clk(gclk));
	jdff dff_A_h4E10oPH3_1(.dout(w_n76_0[1]),.din(w_dff_A_h4E10oPH3_1),.clk(gclk));
	jdff dff_A_cHjRnBxy3_0(.dout(w_Gid4_0[0]),.din(w_dff_A_cHjRnBxy3_0),.clk(gclk));
	jdff dff_A_JRTUmYCW1_0(.dout(w_dff_A_cHjRnBxy3_0),.din(w_dff_A_JRTUmYCW1_0),.clk(gclk));
	jdff dff_A_ntJ5gssM9_0(.dout(w_dff_A_JRTUmYCW1_0),.din(w_dff_A_ntJ5gssM9_0),.clk(gclk));
	jdff dff_A_meMhRixP4_0(.dout(w_dff_A_ntJ5gssM9_0),.din(w_dff_A_meMhRixP4_0),.clk(gclk));
	jdff dff_A_A41J6o1b2_0(.dout(w_dff_A_meMhRixP4_0),.din(w_dff_A_A41J6o1b2_0),.clk(gclk));
	jdff dff_A_U8Hfjj2e2_0(.dout(w_dff_A_A41J6o1b2_0),.din(w_dff_A_U8Hfjj2e2_0),.clk(gclk));
	jdff dff_A_L4KpYBWZ2_0(.dout(w_dff_A_U8Hfjj2e2_0),.din(w_dff_A_L4KpYBWZ2_0),.clk(gclk));
	jdff dff_A_xqOlH3Yn3_0(.dout(w_dff_A_L4KpYBWZ2_0),.din(w_dff_A_xqOlH3Yn3_0),.clk(gclk));
	jdff dff_A_23xFbOV76_0(.dout(w_dff_A_xqOlH3Yn3_0),.din(w_dff_A_23xFbOV76_0),.clk(gclk));
	jdff dff_A_45nYmdsw5_0(.dout(w_dff_A_23xFbOV76_0),.din(w_dff_A_45nYmdsw5_0),.clk(gclk));
	jdff dff_A_RzDX4wxU4_0(.dout(w_Gid0_0[0]),.din(w_dff_A_RzDX4wxU4_0),.clk(gclk));
	jdff dff_A_0Q5O5aZM4_0(.dout(w_dff_A_RzDX4wxU4_0),.din(w_dff_A_0Q5O5aZM4_0),.clk(gclk));
	jdff dff_A_p9R3FxQu2_0(.dout(w_dff_A_0Q5O5aZM4_0),.din(w_dff_A_p9R3FxQu2_0),.clk(gclk));
	jdff dff_A_cFJWuGx49_0(.dout(w_dff_A_p9R3FxQu2_0),.din(w_dff_A_cFJWuGx49_0),.clk(gclk));
	jdff dff_A_GIYOLG237_0(.dout(w_dff_A_cFJWuGx49_0),.din(w_dff_A_GIYOLG237_0),.clk(gclk));
	jdff dff_A_5rg81iup9_0(.dout(w_dff_A_GIYOLG237_0),.din(w_dff_A_5rg81iup9_0),.clk(gclk));
	jdff dff_A_eddGRi5j7_0(.dout(w_dff_A_5rg81iup9_0),.din(w_dff_A_eddGRi5j7_0),.clk(gclk));
	jdff dff_A_vXhZ7gUh3_0(.dout(w_dff_A_eddGRi5j7_0),.din(w_dff_A_vXhZ7gUh3_0),.clk(gclk));
	jdff dff_A_PdSI8fnx1_0(.dout(w_dff_A_vXhZ7gUh3_0),.din(w_dff_A_PdSI8fnx1_0),.clk(gclk));
	jdff dff_A_mPGuB67I3_0(.dout(w_dff_A_PdSI8fnx1_0),.din(w_dff_A_mPGuB67I3_0),.clk(gclk));
	jdff dff_A_RfshTlXF4_0(.dout(w_Gid12_0[0]),.din(w_dff_A_RfshTlXF4_0),.clk(gclk));
	jdff dff_A_4HkAsBd42_0(.dout(w_dff_A_RfshTlXF4_0),.din(w_dff_A_4HkAsBd42_0),.clk(gclk));
	jdff dff_A_F4QdNfe19_0(.dout(w_dff_A_4HkAsBd42_0),.din(w_dff_A_F4QdNfe19_0),.clk(gclk));
	jdff dff_A_oIdDMQgo5_0(.dout(w_dff_A_F4QdNfe19_0),.din(w_dff_A_oIdDMQgo5_0),.clk(gclk));
	jdff dff_A_FBsyP8q70_0(.dout(w_dff_A_oIdDMQgo5_0),.din(w_dff_A_FBsyP8q70_0),.clk(gclk));
	jdff dff_A_btI128zX7_0(.dout(w_dff_A_FBsyP8q70_0),.din(w_dff_A_btI128zX7_0),.clk(gclk));
	jdff dff_A_q2l4SC2z5_0(.dout(w_dff_A_btI128zX7_0),.din(w_dff_A_q2l4SC2z5_0),.clk(gclk));
	jdff dff_A_zGCazSqR4_0(.dout(w_dff_A_q2l4SC2z5_0),.din(w_dff_A_zGCazSqR4_0),.clk(gclk));
	jdff dff_A_e4PhpqOI8_0(.dout(w_dff_A_zGCazSqR4_0),.din(w_dff_A_e4PhpqOI8_0),.clk(gclk));
	jdff dff_A_UzWUyWuH4_0(.dout(w_dff_A_e4PhpqOI8_0),.din(w_dff_A_UzWUyWuH4_0),.clk(gclk));
	jdff dff_A_sjsJuoN04_0(.dout(w_Gid8_0[0]),.din(w_dff_A_sjsJuoN04_0),.clk(gclk));
	jdff dff_A_suIrNB7M6_0(.dout(w_dff_A_sjsJuoN04_0),.din(w_dff_A_suIrNB7M6_0),.clk(gclk));
	jdff dff_A_yvqttXuw3_0(.dout(w_dff_A_suIrNB7M6_0),.din(w_dff_A_yvqttXuw3_0),.clk(gclk));
	jdff dff_A_xd2SLPAM3_0(.dout(w_dff_A_yvqttXuw3_0),.din(w_dff_A_xd2SLPAM3_0),.clk(gclk));
	jdff dff_A_bsMIfAdG0_0(.dout(w_dff_A_xd2SLPAM3_0),.din(w_dff_A_bsMIfAdG0_0),.clk(gclk));
	jdff dff_A_vXBOCL5A2_0(.dout(w_dff_A_bsMIfAdG0_0),.din(w_dff_A_vXBOCL5A2_0),.clk(gclk));
	jdff dff_A_rx0CEOyP5_0(.dout(w_dff_A_vXBOCL5A2_0),.din(w_dff_A_rx0CEOyP5_0),.clk(gclk));
	jdff dff_A_70Je6q9c2_0(.dout(w_dff_A_rx0CEOyP5_0),.din(w_dff_A_70Je6q9c2_0),.clk(gclk));
	jdff dff_A_WtRxzlij2_0(.dout(w_dff_A_70Je6q9c2_0),.din(w_dff_A_WtRxzlij2_0),.clk(gclk));
	jdff dff_A_R5CqIMM82_0(.dout(w_dff_A_WtRxzlij2_0),.din(w_dff_A_R5CqIMM82_0),.clk(gclk));
	jdff dff_B_7bfFOply5_2(.din(n242),.dout(w_dff_B_7bfFOply5_2),.clk(gclk));
	jdff dff_B_cCHm3leD5_2(.din(w_dff_B_7bfFOply5_2),.dout(w_dff_B_cCHm3leD5_2),.clk(gclk));
	jdff dff_B_lMxa1oXZ0_2(.din(w_dff_B_cCHm3leD5_2),.dout(w_dff_B_lMxa1oXZ0_2),.clk(gclk));
	jdff dff_B_q2Ij04a04_2(.din(w_dff_B_lMxa1oXZ0_2),.dout(w_dff_B_q2Ij04a04_2),.clk(gclk));
	jdff dff_A_VOw69Q4S9_0(.dout(w_Gid6_0[0]),.din(w_dff_A_VOw69Q4S9_0),.clk(gclk));
	jdff dff_A_PK6uusgM9_0(.dout(w_dff_A_VOw69Q4S9_0),.din(w_dff_A_PK6uusgM9_0),.clk(gclk));
	jdff dff_A_fOvJW4xP6_0(.dout(w_dff_A_PK6uusgM9_0),.din(w_dff_A_fOvJW4xP6_0),.clk(gclk));
	jdff dff_A_v320Hgdd9_0(.dout(w_dff_A_fOvJW4xP6_0),.din(w_dff_A_v320Hgdd9_0),.clk(gclk));
	jdff dff_A_o65peZUF4_0(.dout(w_dff_A_v320Hgdd9_0),.din(w_dff_A_o65peZUF4_0),.clk(gclk));
	jdff dff_A_pw6h5Ib81_0(.dout(w_dff_A_o65peZUF4_0),.din(w_dff_A_pw6h5Ib81_0),.clk(gclk));
	jdff dff_A_u5gmwgAq8_0(.dout(w_dff_A_pw6h5Ib81_0),.din(w_dff_A_u5gmwgAq8_0),.clk(gclk));
	jdff dff_A_9TD7mNXE9_0(.dout(w_dff_A_u5gmwgAq8_0),.din(w_dff_A_9TD7mNXE9_0),.clk(gclk));
	jdff dff_A_VPJegpDt5_0(.dout(w_dff_A_9TD7mNXE9_0),.din(w_dff_A_VPJegpDt5_0),.clk(gclk));
	jdff dff_A_tn5P6gzj0_0(.dout(w_dff_A_VPJegpDt5_0),.din(w_dff_A_tn5P6gzj0_0),.clk(gclk));
	jdff dff_A_VbyMVxYj9_0(.dout(w_Gid2_0[0]),.din(w_dff_A_VbyMVxYj9_0),.clk(gclk));
	jdff dff_A_GsIAFlQd8_0(.dout(w_dff_A_VbyMVxYj9_0),.din(w_dff_A_GsIAFlQd8_0),.clk(gclk));
	jdff dff_A_Bwilk3af1_0(.dout(w_dff_A_GsIAFlQd8_0),.din(w_dff_A_Bwilk3af1_0),.clk(gclk));
	jdff dff_A_QzTvfGdj4_0(.dout(w_dff_A_Bwilk3af1_0),.din(w_dff_A_QzTvfGdj4_0),.clk(gclk));
	jdff dff_A_tlxPseM01_0(.dout(w_dff_A_QzTvfGdj4_0),.din(w_dff_A_tlxPseM01_0),.clk(gclk));
	jdff dff_A_1zdsX12Y0_0(.dout(w_dff_A_tlxPseM01_0),.din(w_dff_A_1zdsX12Y0_0),.clk(gclk));
	jdff dff_A_eElExFlk9_0(.dout(w_dff_A_1zdsX12Y0_0),.din(w_dff_A_eElExFlk9_0),.clk(gclk));
	jdff dff_A_UPxqfPJI7_0(.dout(w_dff_A_eElExFlk9_0),.din(w_dff_A_UPxqfPJI7_0),.clk(gclk));
	jdff dff_A_D31qGBF63_0(.dout(w_dff_A_UPxqfPJI7_0),.din(w_dff_A_D31qGBF63_0),.clk(gclk));
	jdff dff_A_QrUoxd2A3_0(.dout(w_dff_A_D31qGBF63_0),.din(w_dff_A_QrUoxd2A3_0),.clk(gclk));
	jdff dff_A_m45EXfcm5_0(.dout(w_Gid14_0[0]),.din(w_dff_A_m45EXfcm5_0),.clk(gclk));
	jdff dff_A_I0gkpmK81_0(.dout(w_dff_A_m45EXfcm5_0),.din(w_dff_A_I0gkpmK81_0),.clk(gclk));
	jdff dff_A_7uLpjd9s5_0(.dout(w_dff_A_I0gkpmK81_0),.din(w_dff_A_7uLpjd9s5_0),.clk(gclk));
	jdff dff_A_h2uxgz751_0(.dout(w_dff_A_7uLpjd9s5_0),.din(w_dff_A_h2uxgz751_0),.clk(gclk));
	jdff dff_A_dQ76stEf8_0(.dout(w_dff_A_h2uxgz751_0),.din(w_dff_A_dQ76stEf8_0),.clk(gclk));
	jdff dff_A_pufpSbk40_0(.dout(w_dff_A_dQ76stEf8_0),.din(w_dff_A_pufpSbk40_0),.clk(gclk));
	jdff dff_A_jEOMZGKt5_0(.dout(w_dff_A_pufpSbk40_0),.din(w_dff_A_jEOMZGKt5_0),.clk(gclk));
	jdff dff_A_JXubLcg98_0(.dout(w_dff_A_jEOMZGKt5_0),.din(w_dff_A_JXubLcg98_0),.clk(gclk));
	jdff dff_A_5nbRMX5v0_0(.dout(w_dff_A_JXubLcg98_0),.din(w_dff_A_5nbRMX5v0_0),.clk(gclk));
	jdff dff_A_whgqRjwp1_0(.dout(w_dff_A_5nbRMX5v0_0),.din(w_dff_A_whgqRjwp1_0),.clk(gclk));
	jdff dff_A_GdoRZXIG5_0(.dout(w_Gid10_0[0]),.din(w_dff_A_GdoRZXIG5_0),.clk(gclk));
	jdff dff_A_8LCjIbj19_0(.dout(w_dff_A_GdoRZXIG5_0),.din(w_dff_A_8LCjIbj19_0),.clk(gclk));
	jdff dff_A_FWM7JK3s7_0(.dout(w_dff_A_8LCjIbj19_0),.din(w_dff_A_FWM7JK3s7_0),.clk(gclk));
	jdff dff_A_TC7oSpl93_0(.dout(w_dff_A_FWM7JK3s7_0),.din(w_dff_A_TC7oSpl93_0),.clk(gclk));
	jdff dff_A_e1BCPvu42_0(.dout(w_dff_A_TC7oSpl93_0),.din(w_dff_A_e1BCPvu42_0),.clk(gclk));
	jdff dff_A_eU6Lhmnj2_0(.dout(w_dff_A_e1BCPvu42_0),.din(w_dff_A_eU6Lhmnj2_0),.clk(gclk));
	jdff dff_A_HhPt07mp3_0(.dout(w_dff_A_eU6Lhmnj2_0),.din(w_dff_A_HhPt07mp3_0),.clk(gclk));
	jdff dff_A_f6jCHpFM7_0(.dout(w_dff_A_HhPt07mp3_0),.din(w_dff_A_f6jCHpFM7_0),.clk(gclk));
	jdff dff_A_g8vQeElE0_0(.dout(w_dff_A_f6jCHpFM7_0),.din(w_dff_A_g8vQeElE0_0),.clk(gclk));
	jdff dff_A_vMrH8TvP3_0(.dout(w_dff_A_g8vQeElE0_0),.din(w_dff_A_vMrH8TvP3_0),.clk(gclk));
	jdff dff_A_cASUW5hR5_0(.dout(w_Gid17_0[0]),.din(w_dff_A_cASUW5hR5_0),.clk(gclk));
	jdff dff_A_3RA6tENn7_0(.dout(w_dff_A_cASUW5hR5_0),.din(w_dff_A_3RA6tENn7_0),.clk(gclk));
	jdff dff_A_EXawvFXI8_0(.dout(w_dff_A_3RA6tENn7_0),.din(w_dff_A_EXawvFXI8_0),.clk(gclk));
	jdff dff_A_65aplbU78_0(.dout(w_dff_A_EXawvFXI8_0),.din(w_dff_A_65aplbU78_0),.clk(gclk));
	jdff dff_A_68BJbQ8D3_0(.dout(w_dff_A_65aplbU78_0),.din(w_dff_A_68BJbQ8D3_0),.clk(gclk));
	jdff dff_A_Y33yLsSb7_0(.dout(w_dff_A_68BJbQ8D3_0),.din(w_dff_A_Y33yLsSb7_0),.clk(gclk));
	jdff dff_A_B5CPzabP4_0(.dout(w_dff_A_Y33yLsSb7_0),.din(w_dff_A_B5CPzabP4_0),.clk(gclk));
	jdff dff_A_prlhLW9Z2_0(.dout(w_dff_A_B5CPzabP4_0),.din(w_dff_A_prlhLW9Z2_0),.clk(gclk));
	jdff dff_A_PF7j2tx89_0(.dout(w_dff_A_prlhLW9Z2_0),.din(w_dff_A_PF7j2tx89_0),.clk(gclk));
	jdff dff_A_Ajz5gCAU9_0(.dout(w_dff_A_PF7j2tx89_0),.din(w_dff_A_Ajz5gCAU9_0),.clk(gclk));
	jdff dff_A_3hvJBpol7_0(.dout(w_dff_A_Ajz5gCAU9_0),.din(w_dff_A_3hvJBpol7_0),.clk(gclk));
	jdff dff_A_2P9YjnMl8_0(.dout(w_Gid16_0[0]),.din(w_dff_A_2P9YjnMl8_0),.clk(gclk));
	jdff dff_A_NaWxm0Vu2_0(.dout(w_dff_A_2P9YjnMl8_0),.din(w_dff_A_NaWxm0Vu2_0),.clk(gclk));
	jdff dff_A_UbLBlLK47_0(.dout(w_dff_A_NaWxm0Vu2_0),.din(w_dff_A_UbLBlLK47_0),.clk(gclk));
	jdff dff_A_FvYcQYev2_0(.dout(w_dff_A_UbLBlLK47_0),.din(w_dff_A_FvYcQYev2_0),.clk(gclk));
	jdff dff_A_g3z3w5oC1_0(.dout(w_dff_A_FvYcQYev2_0),.din(w_dff_A_g3z3w5oC1_0),.clk(gclk));
	jdff dff_A_RhQtjhXb3_0(.dout(w_dff_A_g3z3w5oC1_0),.din(w_dff_A_RhQtjhXb3_0),.clk(gclk));
	jdff dff_A_UiipUCVH4_0(.dout(w_dff_A_RhQtjhXb3_0),.din(w_dff_A_UiipUCVH4_0),.clk(gclk));
	jdff dff_A_8K991h965_0(.dout(w_dff_A_UiipUCVH4_0),.din(w_dff_A_8K991h965_0),.clk(gclk));
	jdff dff_A_l8AYu8lY4_0(.dout(w_dff_A_8K991h965_0),.din(w_dff_A_l8AYu8lY4_0),.clk(gclk));
	jdff dff_A_fDsKudNf5_0(.dout(w_dff_A_l8AYu8lY4_0),.din(w_dff_A_fDsKudNf5_0),.clk(gclk));
	jdff dff_A_vcPrUY5d1_0(.dout(w_dff_A_fDsKudNf5_0),.din(w_dff_A_vcPrUY5d1_0),.clk(gclk));
	jdff dff_A_dtvuA91o4_0(.dout(w_Gid19_0[0]),.din(w_dff_A_dtvuA91o4_0),.clk(gclk));
	jdff dff_A_xYnyUA9b2_0(.dout(w_dff_A_dtvuA91o4_0),.din(w_dff_A_xYnyUA9b2_0),.clk(gclk));
	jdff dff_A_nJFnqXJF3_0(.dout(w_dff_A_xYnyUA9b2_0),.din(w_dff_A_nJFnqXJF3_0),.clk(gclk));
	jdff dff_A_ZHeeBaHR4_0(.dout(w_dff_A_nJFnqXJF3_0),.din(w_dff_A_ZHeeBaHR4_0),.clk(gclk));
	jdff dff_A_ZqU9HZ8v1_0(.dout(w_dff_A_ZHeeBaHR4_0),.din(w_dff_A_ZqU9HZ8v1_0),.clk(gclk));
	jdff dff_A_DtzoR74x6_0(.dout(w_dff_A_ZqU9HZ8v1_0),.din(w_dff_A_DtzoR74x6_0),.clk(gclk));
	jdff dff_A_0KiXf2cX7_0(.dout(w_dff_A_DtzoR74x6_0),.din(w_dff_A_0KiXf2cX7_0),.clk(gclk));
	jdff dff_A_0IcjlmqK9_0(.dout(w_dff_A_0KiXf2cX7_0),.din(w_dff_A_0IcjlmqK9_0),.clk(gclk));
	jdff dff_A_OXRPh0kW4_0(.dout(w_dff_A_0IcjlmqK9_0),.din(w_dff_A_OXRPh0kW4_0),.clk(gclk));
	jdff dff_A_6mAf3AwT7_0(.dout(w_dff_A_OXRPh0kW4_0),.din(w_dff_A_6mAf3AwT7_0),.clk(gclk));
	jdff dff_A_48fX9mcn2_0(.dout(w_dff_A_6mAf3AwT7_0),.din(w_dff_A_48fX9mcn2_0),.clk(gclk));
	jdff dff_A_3osGbBNr1_0(.dout(w_Gid18_0[0]),.din(w_dff_A_3osGbBNr1_0),.clk(gclk));
	jdff dff_A_nQCWmlJu7_0(.dout(w_dff_A_3osGbBNr1_0),.din(w_dff_A_nQCWmlJu7_0),.clk(gclk));
	jdff dff_A_Hp5DeOLV0_0(.dout(w_dff_A_nQCWmlJu7_0),.din(w_dff_A_Hp5DeOLV0_0),.clk(gclk));
	jdff dff_A_8LkhMyKa0_0(.dout(w_dff_A_Hp5DeOLV0_0),.din(w_dff_A_8LkhMyKa0_0),.clk(gclk));
	jdff dff_A_4qy07Ypo5_0(.dout(w_dff_A_8LkhMyKa0_0),.din(w_dff_A_4qy07Ypo5_0),.clk(gclk));
	jdff dff_A_x97rfs7l2_0(.dout(w_dff_A_4qy07Ypo5_0),.din(w_dff_A_x97rfs7l2_0),.clk(gclk));
	jdff dff_A_h1OxO95z7_0(.dout(w_dff_A_x97rfs7l2_0),.din(w_dff_A_h1OxO95z7_0),.clk(gclk));
	jdff dff_A_7ZuYobcK0_0(.dout(w_dff_A_h1OxO95z7_0),.din(w_dff_A_7ZuYobcK0_0),.clk(gclk));
	jdff dff_A_hTRPTVZH1_0(.dout(w_dff_A_7ZuYobcK0_0),.din(w_dff_A_hTRPTVZH1_0),.clk(gclk));
	jdff dff_A_qbgQ2jDN7_0(.dout(w_dff_A_hTRPTVZH1_0),.din(w_dff_A_qbgQ2jDN7_0),.clk(gclk));
	jdff dff_A_swKGAntW1_0(.dout(w_dff_A_qbgQ2jDN7_0),.din(w_dff_A_swKGAntW1_0),.clk(gclk));
	jdff dff_A_2LDJkh3t8_0(.dout(w_n136_0[0]),.din(w_dff_A_2LDJkh3t8_0),.clk(gclk));
	jdff dff_A_zJfUTd4q8_0(.dout(w_Gid25_0[0]),.din(w_dff_A_zJfUTd4q8_0),.clk(gclk));
	jdff dff_A_ZDrkqYjG0_0(.dout(w_dff_A_zJfUTd4q8_0),.din(w_dff_A_ZDrkqYjG0_0),.clk(gclk));
	jdff dff_A_0vXoOyjT0_0(.dout(w_dff_A_ZDrkqYjG0_0),.din(w_dff_A_0vXoOyjT0_0),.clk(gclk));
	jdff dff_A_5Q5qA0642_0(.dout(w_dff_A_0vXoOyjT0_0),.din(w_dff_A_5Q5qA0642_0),.clk(gclk));
	jdff dff_A_gYVOYK0p1_0(.dout(w_dff_A_5Q5qA0642_0),.din(w_dff_A_gYVOYK0p1_0),.clk(gclk));
	jdff dff_A_UJmpBvXi7_0(.dout(w_dff_A_gYVOYK0p1_0),.din(w_dff_A_UJmpBvXi7_0),.clk(gclk));
	jdff dff_A_uDsOVl0F8_0(.dout(w_dff_A_UJmpBvXi7_0),.din(w_dff_A_uDsOVl0F8_0),.clk(gclk));
	jdff dff_A_iODDi2CH9_0(.dout(w_dff_A_uDsOVl0F8_0),.din(w_dff_A_iODDi2CH9_0),.clk(gclk));
	jdff dff_A_gwoAee4U9_0(.dout(w_dff_A_iODDi2CH9_0),.din(w_dff_A_gwoAee4U9_0),.clk(gclk));
	jdff dff_A_TvXjSViK8_0(.dout(w_dff_A_gwoAee4U9_0),.din(w_dff_A_TvXjSViK8_0),.clk(gclk));
	jdff dff_A_IKEsPeSf3_0(.dout(w_dff_A_TvXjSViK8_0),.din(w_dff_A_IKEsPeSf3_0),.clk(gclk));
	jdff dff_A_8WEIMdgR7_0(.dout(w_Gid24_0[0]),.din(w_dff_A_8WEIMdgR7_0),.clk(gclk));
	jdff dff_A_CLwDdsUQ3_0(.dout(w_dff_A_8WEIMdgR7_0),.din(w_dff_A_CLwDdsUQ3_0),.clk(gclk));
	jdff dff_A_p84QDqHd2_0(.dout(w_dff_A_CLwDdsUQ3_0),.din(w_dff_A_p84QDqHd2_0),.clk(gclk));
	jdff dff_A_IGBZRrqz4_0(.dout(w_dff_A_p84QDqHd2_0),.din(w_dff_A_IGBZRrqz4_0),.clk(gclk));
	jdff dff_A_zj45PG1S7_0(.dout(w_dff_A_IGBZRrqz4_0),.din(w_dff_A_zj45PG1S7_0),.clk(gclk));
	jdff dff_A_6GUgtQJS9_0(.dout(w_dff_A_zj45PG1S7_0),.din(w_dff_A_6GUgtQJS9_0),.clk(gclk));
	jdff dff_A_tUs3HHDq8_0(.dout(w_dff_A_6GUgtQJS9_0),.din(w_dff_A_tUs3HHDq8_0),.clk(gclk));
	jdff dff_A_7i76XiWq5_0(.dout(w_dff_A_tUs3HHDq8_0),.din(w_dff_A_7i76XiWq5_0),.clk(gclk));
	jdff dff_A_JCF0EKvh4_0(.dout(w_dff_A_7i76XiWq5_0),.din(w_dff_A_JCF0EKvh4_0),.clk(gclk));
	jdff dff_A_luKafPcj5_0(.dout(w_dff_A_JCF0EKvh4_0),.din(w_dff_A_luKafPcj5_0),.clk(gclk));
	jdff dff_A_YvK4cSR30_0(.dout(w_dff_A_luKafPcj5_0),.din(w_dff_A_YvK4cSR30_0),.clk(gclk));
	jdff dff_A_3vm7JMe32_0(.dout(w_Gid27_0[0]),.din(w_dff_A_3vm7JMe32_0),.clk(gclk));
	jdff dff_A_OBmMmhu55_0(.dout(w_dff_A_3vm7JMe32_0),.din(w_dff_A_OBmMmhu55_0),.clk(gclk));
	jdff dff_A_EuTwiRAA3_0(.dout(w_dff_A_OBmMmhu55_0),.din(w_dff_A_EuTwiRAA3_0),.clk(gclk));
	jdff dff_A_rLjbzQKE6_0(.dout(w_dff_A_EuTwiRAA3_0),.din(w_dff_A_rLjbzQKE6_0),.clk(gclk));
	jdff dff_A_e9BCc0k89_0(.dout(w_dff_A_rLjbzQKE6_0),.din(w_dff_A_e9BCc0k89_0),.clk(gclk));
	jdff dff_A_041ZalXw9_0(.dout(w_dff_A_e9BCc0k89_0),.din(w_dff_A_041ZalXw9_0),.clk(gclk));
	jdff dff_A_fHLJIFQ38_0(.dout(w_dff_A_041ZalXw9_0),.din(w_dff_A_fHLJIFQ38_0),.clk(gclk));
	jdff dff_A_LwhnlwNA6_0(.dout(w_dff_A_fHLJIFQ38_0),.din(w_dff_A_LwhnlwNA6_0),.clk(gclk));
	jdff dff_A_gUwHN94g7_0(.dout(w_dff_A_LwhnlwNA6_0),.din(w_dff_A_gUwHN94g7_0),.clk(gclk));
	jdff dff_A_KgZ5YJTo9_0(.dout(w_dff_A_gUwHN94g7_0),.din(w_dff_A_KgZ5YJTo9_0),.clk(gclk));
	jdff dff_A_Trwj7LQB3_0(.dout(w_dff_A_KgZ5YJTo9_0),.din(w_dff_A_Trwj7LQB3_0),.clk(gclk));
	jdff dff_A_I4GWRoe42_0(.dout(w_Gid26_0[0]),.din(w_dff_A_I4GWRoe42_0),.clk(gclk));
	jdff dff_A_7dXePNXv4_0(.dout(w_dff_A_I4GWRoe42_0),.din(w_dff_A_7dXePNXv4_0),.clk(gclk));
	jdff dff_A_ciMjUmTy3_0(.dout(w_dff_A_7dXePNXv4_0),.din(w_dff_A_ciMjUmTy3_0),.clk(gclk));
	jdff dff_A_s2YLLYJL1_0(.dout(w_dff_A_ciMjUmTy3_0),.din(w_dff_A_s2YLLYJL1_0),.clk(gclk));
	jdff dff_A_LHlD12sB5_0(.dout(w_dff_A_s2YLLYJL1_0),.din(w_dff_A_LHlD12sB5_0),.clk(gclk));
	jdff dff_A_XBz8Iay49_0(.dout(w_dff_A_LHlD12sB5_0),.din(w_dff_A_XBz8Iay49_0),.clk(gclk));
	jdff dff_A_XraUgurW5_0(.dout(w_dff_A_XBz8Iay49_0),.din(w_dff_A_XraUgurW5_0),.clk(gclk));
	jdff dff_A_olOnVLQo1_0(.dout(w_dff_A_XraUgurW5_0),.din(w_dff_A_olOnVLQo1_0),.clk(gclk));
	jdff dff_A_52hF7bX48_0(.dout(w_dff_A_olOnVLQo1_0),.din(w_dff_A_52hF7bX48_0),.clk(gclk));
	jdff dff_A_wiKkNZ6w2_0(.dout(w_dff_A_52hF7bX48_0),.din(w_dff_A_wiKkNZ6w2_0),.clk(gclk));
	jdff dff_A_cPxyNrLc5_0(.dout(w_dff_A_wiKkNZ6w2_0),.din(w_dff_A_cPxyNrLc5_0),.clk(gclk));
	jdff dff_A_trgskhLC3_0(.dout(w_n147_0[0]),.din(w_dff_A_trgskhLC3_0),.clk(gclk));
	jdff dff_A_nNMzKHqI9_0(.dout(w_dff_A_trgskhLC3_0),.din(w_dff_A_nNMzKHqI9_0),.clk(gclk));
	jdff dff_A_MNZtudzM7_0(.dout(w_dff_A_nNMzKHqI9_0),.din(w_dff_A_MNZtudzM7_0),.clk(gclk));
	jdff dff_A_Emcxli7F3_0(.dout(w_dff_A_MNZtudzM7_0),.din(w_dff_A_Emcxli7F3_0),.clk(gclk));
	jdff dff_A_4qEya7Iu6_0(.dout(w_dff_A_Emcxli7F3_0),.din(w_dff_A_4qEya7Iu6_0),.clk(gclk));
	jdff dff_A_QMle7d0n5_0(.dout(w_Gid7_0[0]),.din(w_dff_A_QMle7d0n5_0),.clk(gclk));
	jdff dff_A_Uask23rq9_0(.dout(w_dff_A_QMle7d0n5_0),.din(w_dff_A_Uask23rq9_0),.clk(gclk));
	jdff dff_A_L0dnapZQ4_0(.dout(w_dff_A_Uask23rq9_0),.din(w_dff_A_L0dnapZQ4_0),.clk(gclk));
	jdff dff_A_8cZ2XvID8_0(.dout(w_dff_A_L0dnapZQ4_0),.din(w_dff_A_8cZ2XvID8_0),.clk(gclk));
	jdff dff_A_dnRLACyM0_0(.dout(w_dff_A_8cZ2XvID8_0),.din(w_dff_A_dnRLACyM0_0),.clk(gclk));
	jdff dff_A_o1k0E09P9_0(.dout(w_dff_A_dnRLACyM0_0),.din(w_dff_A_o1k0E09P9_0),.clk(gclk));
	jdff dff_A_4azYrVDd9_0(.dout(w_dff_A_o1k0E09P9_0),.din(w_dff_A_4azYrVDd9_0),.clk(gclk));
	jdff dff_A_3VzZp6fV1_0(.dout(w_dff_A_4azYrVDd9_0),.din(w_dff_A_3VzZp6fV1_0),.clk(gclk));
	jdff dff_A_Ib0LBkQ53_0(.dout(w_dff_A_3VzZp6fV1_0),.din(w_dff_A_Ib0LBkQ53_0),.clk(gclk));
	jdff dff_A_QydXU8MJ2_0(.dout(w_dff_A_Ib0LBkQ53_0),.din(w_dff_A_QydXU8MJ2_0),.clk(gclk));
	jdff dff_A_x29eqbbc9_0(.dout(w_Gid3_0[0]),.din(w_dff_A_x29eqbbc9_0),.clk(gclk));
	jdff dff_A_gt2eYnkQ7_0(.dout(w_dff_A_x29eqbbc9_0),.din(w_dff_A_gt2eYnkQ7_0),.clk(gclk));
	jdff dff_A_Nui8Siru6_0(.dout(w_dff_A_gt2eYnkQ7_0),.din(w_dff_A_Nui8Siru6_0),.clk(gclk));
	jdff dff_A_rF4NN6kG4_0(.dout(w_dff_A_Nui8Siru6_0),.din(w_dff_A_rF4NN6kG4_0),.clk(gclk));
	jdff dff_A_UaHlL3YW6_0(.dout(w_dff_A_rF4NN6kG4_0),.din(w_dff_A_UaHlL3YW6_0),.clk(gclk));
	jdff dff_A_B3s3Xmxd5_0(.dout(w_dff_A_UaHlL3YW6_0),.din(w_dff_A_B3s3Xmxd5_0),.clk(gclk));
	jdff dff_A_rpyOg9iQ7_0(.dout(w_dff_A_B3s3Xmxd5_0),.din(w_dff_A_rpyOg9iQ7_0),.clk(gclk));
	jdff dff_A_quShtIId7_0(.dout(w_dff_A_rpyOg9iQ7_0),.din(w_dff_A_quShtIId7_0),.clk(gclk));
	jdff dff_A_xKTCn2ip9_0(.dout(w_dff_A_quShtIId7_0),.din(w_dff_A_xKTCn2ip9_0),.clk(gclk));
	jdff dff_A_Ob44XYIB0_0(.dout(w_dff_A_xKTCn2ip9_0),.din(w_dff_A_Ob44XYIB0_0),.clk(gclk));
	jdff dff_A_JbNBaWVt4_0(.dout(w_Gid15_0[0]),.din(w_dff_A_JbNBaWVt4_0),.clk(gclk));
	jdff dff_A_UgT0i45a7_0(.dout(w_dff_A_JbNBaWVt4_0),.din(w_dff_A_UgT0i45a7_0),.clk(gclk));
	jdff dff_A_Ox8FXqk35_0(.dout(w_dff_A_UgT0i45a7_0),.din(w_dff_A_Ox8FXqk35_0),.clk(gclk));
	jdff dff_A_gyYCP9vq7_0(.dout(w_dff_A_Ox8FXqk35_0),.din(w_dff_A_gyYCP9vq7_0),.clk(gclk));
	jdff dff_A_ZxTT2OXD6_0(.dout(w_dff_A_gyYCP9vq7_0),.din(w_dff_A_ZxTT2OXD6_0),.clk(gclk));
	jdff dff_A_eez2zmGH1_0(.dout(w_dff_A_ZxTT2OXD6_0),.din(w_dff_A_eez2zmGH1_0),.clk(gclk));
	jdff dff_A_buFgwA2A6_0(.dout(w_dff_A_eez2zmGH1_0),.din(w_dff_A_buFgwA2A6_0),.clk(gclk));
	jdff dff_A_kPOjCu7D2_0(.dout(w_dff_A_buFgwA2A6_0),.din(w_dff_A_kPOjCu7D2_0),.clk(gclk));
	jdff dff_A_T4fA4E962_0(.dout(w_dff_A_kPOjCu7D2_0),.din(w_dff_A_T4fA4E962_0),.clk(gclk));
	jdff dff_A_zDinP9BW2_0(.dout(w_dff_A_T4fA4E962_0),.din(w_dff_A_zDinP9BW2_0),.clk(gclk));
	jdff dff_A_RV9iZpna7_0(.dout(w_Gid11_0[0]),.din(w_dff_A_RV9iZpna7_0),.clk(gclk));
	jdff dff_A_48nMjq3h3_0(.dout(w_dff_A_RV9iZpna7_0),.din(w_dff_A_48nMjq3h3_0),.clk(gclk));
	jdff dff_A_zee0PFFx7_0(.dout(w_dff_A_48nMjq3h3_0),.din(w_dff_A_zee0PFFx7_0),.clk(gclk));
	jdff dff_A_ImYl7bbI2_0(.dout(w_dff_A_zee0PFFx7_0),.din(w_dff_A_ImYl7bbI2_0),.clk(gclk));
	jdff dff_A_j95C3OIv4_0(.dout(w_dff_A_ImYl7bbI2_0),.din(w_dff_A_j95C3OIv4_0),.clk(gclk));
	jdff dff_A_oELo6KbY4_0(.dout(w_dff_A_j95C3OIv4_0),.din(w_dff_A_oELo6KbY4_0),.clk(gclk));
	jdff dff_A_GQuxPzKt6_0(.dout(w_dff_A_oELo6KbY4_0),.din(w_dff_A_GQuxPzKt6_0),.clk(gclk));
	jdff dff_A_LKbD6RPp6_0(.dout(w_dff_A_GQuxPzKt6_0),.din(w_dff_A_LKbD6RPp6_0),.clk(gclk));
	jdff dff_A_pWVRce4r7_0(.dout(w_dff_A_LKbD6RPp6_0),.din(w_dff_A_pWVRce4r7_0),.clk(gclk));
	jdff dff_A_FEmzwO6L8_0(.dout(w_dff_A_pWVRce4r7_0),.din(w_dff_A_FEmzwO6L8_0),.clk(gclk));
	jdff dff_A_nFNYR6Rh8_0(.dout(w_Gid21_0[0]),.din(w_dff_A_nFNYR6Rh8_0),.clk(gclk));
	jdff dff_A_htS3z7by4_0(.dout(w_dff_A_nFNYR6Rh8_0),.din(w_dff_A_htS3z7by4_0),.clk(gclk));
	jdff dff_A_TWSLCyWV2_0(.dout(w_dff_A_htS3z7by4_0),.din(w_dff_A_TWSLCyWV2_0),.clk(gclk));
	jdff dff_A_1KYJRseF7_0(.dout(w_dff_A_TWSLCyWV2_0),.din(w_dff_A_1KYJRseF7_0),.clk(gclk));
	jdff dff_A_Pg6Sjzua4_0(.dout(w_dff_A_1KYJRseF7_0),.din(w_dff_A_Pg6Sjzua4_0),.clk(gclk));
	jdff dff_A_5m77TeH39_0(.dout(w_dff_A_Pg6Sjzua4_0),.din(w_dff_A_5m77TeH39_0),.clk(gclk));
	jdff dff_A_pjcVxXi56_0(.dout(w_dff_A_5m77TeH39_0),.din(w_dff_A_pjcVxXi56_0),.clk(gclk));
	jdff dff_A_HhRBAEDp7_0(.dout(w_dff_A_pjcVxXi56_0),.din(w_dff_A_HhRBAEDp7_0),.clk(gclk));
	jdff dff_A_5bnA5CB90_0(.dout(w_dff_A_HhRBAEDp7_0),.din(w_dff_A_5bnA5CB90_0),.clk(gclk));
	jdff dff_A_RtkDc7Dv4_0(.dout(w_dff_A_5bnA5CB90_0),.din(w_dff_A_RtkDc7Dv4_0),.clk(gclk));
	jdff dff_A_yIuxIPZN8_0(.dout(w_dff_A_RtkDc7Dv4_0),.din(w_dff_A_yIuxIPZN8_0),.clk(gclk));
	jdff dff_A_IoQM1IDB9_0(.dout(w_Gid20_0[0]),.din(w_dff_A_IoQM1IDB9_0),.clk(gclk));
	jdff dff_A_U1vFxNb61_0(.dout(w_dff_A_IoQM1IDB9_0),.din(w_dff_A_U1vFxNb61_0),.clk(gclk));
	jdff dff_A_EnUdaxB08_0(.dout(w_dff_A_U1vFxNb61_0),.din(w_dff_A_EnUdaxB08_0),.clk(gclk));
	jdff dff_A_7lphQtNi1_0(.dout(w_dff_A_EnUdaxB08_0),.din(w_dff_A_7lphQtNi1_0),.clk(gclk));
	jdff dff_A_s506qQm57_0(.dout(w_dff_A_7lphQtNi1_0),.din(w_dff_A_s506qQm57_0),.clk(gclk));
	jdff dff_A_5G4JXHHt5_0(.dout(w_dff_A_s506qQm57_0),.din(w_dff_A_5G4JXHHt5_0),.clk(gclk));
	jdff dff_A_uDLRzEar5_0(.dout(w_dff_A_5G4JXHHt5_0),.din(w_dff_A_uDLRzEar5_0),.clk(gclk));
	jdff dff_A_JIYmvVR86_0(.dout(w_dff_A_uDLRzEar5_0),.din(w_dff_A_JIYmvVR86_0),.clk(gclk));
	jdff dff_A_kaxjGrzs2_0(.dout(w_dff_A_JIYmvVR86_0),.din(w_dff_A_kaxjGrzs2_0),.clk(gclk));
	jdff dff_A_RoU1uwMN6_0(.dout(w_dff_A_kaxjGrzs2_0),.din(w_dff_A_RoU1uwMN6_0),.clk(gclk));
	jdff dff_A_lgfvsrkH8_0(.dout(w_dff_A_RoU1uwMN6_0),.din(w_dff_A_lgfvsrkH8_0),.clk(gclk));
	jdff dff_A_LYdN8MiC6_0(.dout(w_Gid23_0[0]),.din(w_dff_A_LYdN8MiC6_0),.clk(gclk));
	jdff dff_A_m54Sm2SY7_0(.dout(w_dff_A_LYdN8MiC6_0),.din(w_dff_A_m54Sm2SY7_0),.clk(gclk));
	jdff dff_A_0GLQNQEO1_0(.dout(w_dff_A_m54Sm2SY7_0),.din(w_dff_A_0GLQNQEO1_0),.clk(gclk));
	jdff dff_A_IrMCqxkP2_0(.dout(w_dff_A_0GLQNQEO1_0),.din(w_dff_A_IrMCqxkP2_0),.clk(gclk));
	jdff dff_A_slFS2xON7_0(.dout(w_dff_A_IrMCqxkP2_0),.din(w_dff_A_slFS2xON7_0),.clk(gclk));
	jdff dff_A_eoiM19aI5_0(.dout(w_dff_A_slFS2xON7_0),.din(w_dff_A_eoiM19aI5_0),.clk(gclk));
	jdff dff_A_jQXMnGLa6_0(.dout(w_dff_A_eoiM19aI5_0),.din(w_dff_A_jQXMnGLa6_0),.clk(gclk));
	jdff dff_A_xOWaKdHa1_0(.dout(w_dff_A_jQXMnGLa6_0),.din(w_dff_A_xOWaKdHa1_0),.clk(gclk));
	jdff dff_A_CFYOo6Dg7_0(.dout(w_dff_A_xOWaKdHa1_0),.din(w_dff_A_CFYOo6Dg7_0),.clk(gclk));
	jdff dff_A_b0TOLugh7_0(.dout(w_dff_A_CFYOo6Dg7_0),.din(w_dff_A_b0TOLugh7_0),.clk(gclk));
	jdff dff_A_D7URHJsV8_0(.dout(w_dff_A_b0TOLugh7_0),.din(w_dff_A_D7URHJsV8_0),.clk(gclk));
	jdff dff_A_e0dDOrGk2_0(.dout(w_Gid22_0[0]),.din(w_dff_A_e0dDOrGk2_0),.clk(gclk));
	jdff dff_A_z1dcoJah6_0(.dout(w_dff_A_e0dDOrGk2_0),.din(w_dff_A_z1dcoJah6_0),.clk(gclk));
	jdff dff_A_eJ6E6ibW1_0(.dout(w_dff_A_z1dcoJah6_0),.din(w_dff_A_eJ6E6ibW1_0),.clk(gclk));
	jdff dff_A_0tpNe0sL6_0(.dout(w_dff_A_eJ6E6ibW1_0),.din(w_dff_A_0tpNe0sL6_0),.clk(gclk));
	jdff dff_A_HEepittY7_0(.dout(w_dff_A_0tpNe0sL6_0),.din(w_dff_A_HEepittY7_0),.clk(gclk));
	jdff dff_A_7MOUxzP32_0(.dout(w_dff_A_HEepittY7_0),.din(w_dff_A_7MOUxzP32_0),.clk(gclk));
	jdff dff_A_lZWHOGJ01_0(.dout(w_dff_A_7MOUxzP32_0),.din(w_dff_A_lZWHOGJ01_0),.clk(gclk));
	jdff dff_A_AO9QGGjU0_0(.dout(w_dff_A_lZWHOGJ01_0),.din(w_dff_A_AO9QGGjU0_0),.clk(gclk));
	jdff dff_A_rlF4guPS3_0(.dout(w_dff_A_AO9QGGjU0_0),.din(w_dff_A_rlF4guPS3_0),.clk(gclk));
	jdff dff_A_HDG8o1MW2_0(.dout(w_dff_A_rlF4guPS3_0),.din(w_dff_A_HDG8o1MW2_0),.clk(gclk));
	jdff dff_A_itpsinfy8_0(.dout(w_dff_A_HDG8o1MW2_0),.din(w_dff_A_itpsinfy8_0),.clk(gclk));
	jdff dff_A_mWAiAKq28_0(.dout(w_n128_0[0]),.din(w_dff_A_mWAiAKq28_0),.clk(gclk));
	jdff dff_A_Nde5DTjx7_0(.dout(w_Gid29_0[0]),.din(w_dff_A_Nde5DTjx7_0),.clk(gclk));
	jdff dff_A_j2Jl1zX12_0(.dout(w_dff_A_Nde5DTjx7_0),.din(w_dff_A_j2Jl1zX12_0),.clk(gclk));
	jdff dff_A_6EMXGX7K5_0(.dout(w_dff_A_j2Jl1zX12_0),.din(w_dff_A_6EMXGX7K5_0),.clk(gclk));
	jdff dff_A_gVxcNbrD3_0(.dout(w_dff_A_6EMXGX7K5_0),.din(w_dff_A_gVxcNbrD3_0),.clk(gclk));
	jdff dff_A_PCqWS4FX8_0(.dout(w_dff_A_gVxcNbrD3_0),.din(w_dff_A_PCqWS4FX8_0),.clk(gclk));
	jdff dff_A_2PhElid30_0(.dout(w_dff_A_PCqWS4FX8_0),.din(w_dff_A_2PhElid30_0),.clk(gclk));
	jdff dff_A_02ACiawp3_0(.dout(w_dff_A_2PhElid30_0),.din(w_dff_A_02ACiawp3_0),.clk(gclk));
	jdff dff_A_ZE2YkXj61_0(.dout(w_dff_A_02ACiawp3_0),.din(w_dff_A_ZE2YkXj61_0),.clk(gclk));
	jdff dff_A_QNDgQq9I7_0(.dout(w_dff_A_ZE2YkXj61_0),.din(w_dff_A_QNDgQq9I7_0),.clk(gclk));
	jdff dff_A_UG1DeCEJ9_0(.dout(w_dff_A_QNDgQq9I7_0),.din(w_dff_A_UG1DeCEJ9_0),.clk(gclk));
	jdff dff_A_U9iWXrnT9_0(.dout(w_dff_A_UG1DeCEJ9_0),.din(w_dff_A_U9iWXrnT9_0),.clk(gclk));
	jdff dff_A_7IrYAtEj3_0(.dout(w_Gid28_0[0]),.din(w_dff_A_7IrYAtEj3_0),.clk(gclk));
	jdff dff_A_MvyTxmeJ9_0(.dout(w_dff_A_7IrYAtEj3_0),.din(w_dff_A_MvyTxmeJ9_0),.clk(gclk));
	jdff dff_A_UW1KUhnE1_0(.dout(w_dff_A_MvyTxmeJ9_0),.din(w_dff_A_UW1KUhnE1_0),.clk(gclk));
	jdff dff_A_5Xk5mWEQ3_0(.dout(w_dff_A_UW1KUhnE1_0),.din(w_dff_A_5Xk5mWEQ3_0),.clk(gclk));
	jdff dff_A_2ncx7ghg9_0(.dout(w_dff_A_5Xk5mWEQ3_0),.din(w_dff_A_2ncx7ghg9_0),.clk(gclk));
	jdff dff_A_kQDGFQS41_0(.dout(w_dff_A_2ncx7ghg9_0),.din(w_dff_A_kQDGFQS41_0),.clk(gclk));
	jdff dff_A_DN2GL6VX9_0(.dout(w_dff_A_kQDGFQS41_0),.din(w_dff_A_DN2GL6VX9_0),.clk(gclk));
	jdff dff_A_r0UfnC7k9_0(.dout(w_dff_A_DN2GL6VX9_0),.din(w_dff_A_r0UfnC7k9_0),.clk(gclk));
	jdff dff_A_VV47jh2h5_0(.dout(w_dff_A_r0UfnC7k9_0),.din(w_dff_A_VV47jh2h5_0),.clk(gclk));
	jdff dff_A_7OG5vszE2_0(.dout(w_dff_A_VV47jh2h5_0),.din(w_dff_A_7OG5vszE2_0),.clk(gclk));
	jdff dff_A_89jrkGWO8_0(.dout(w_dff_A_7OG5vszE2_0),.din(w_dff_A_89jrkGWO8_0),.clk(gclk));
	jdff dff_A_KcPfHo4i8_0(.dout(w_Gid31_0[0]),.din(w_dff_A_KcPfHo4i8_0),.clk(gclk));
	jdff dff_A_26dNHKoN0_0(.dout(w_dff_A_KcPfHo4i8_0),.din(w_dff_A_26dNHKoN0_0),.clk(gclk));
	jdff dff_A_SIUIpMYO3_0(.dout(w_dff_A_26dNHKoN0_0),.din(w_dff_A_SIUIpMYO3_0),.clk(gclk));
	jdff dff_A_EXZ40ExW8_0(.dout(w_dff_A_SIUIpMYO3_0),.din(w_dff_A_EXZ40ExW8_0),.clk(gclk));
	jdff dff_A_zjYQiali2_0(.dout(w_dff_A_EXZ40ExW8_0),.din(w_dff_A_zjYQiali2_0),.clk(gclk));
	jdff dff_A_PiNvl5Oa2_0(.dout(w_dff_A_zjYQiali2_0),.din(w_dff_A_PiNvl5Oa2_0),.clk(gclk));
	jdff dff_A_PRPEmvZp8_0(.dout(w_dff_A_PiNvl5Oa2_0),.din(w_dff_A_PRPEmvZp8_0),.clk(gclk));
	jdff dff_A_RwXCACcd3_0(.dout(w_dff_A_PRPEmvZp8_0),.din(w_dff_A_RwXCACcd3_0),.clk(gclk));
	jdff dff_A_WCpZzk0x8_0(.dout(w_dff_A_RwXCACcd3_0),.din(w_dff_A_WCpZzk0x8_0),.clk(gclk));
	jdff dff_A_b00r57cX9_0(.dout(w_dff_A_WCpZzk0x8_0),.din(w_dff_A_b00r57cX9_0),.clk(gclk));
	jdff dff_A_jrTa5pKo7_0(.dout(w_dff_A_b00r57cX9_0),.din(w_dff_A_jrTa5pKo7_0),.clk(gclk));
	jdff dff_A_fbe2HY1E3_0(.dout(w_Gid30_0[0]),.din(w_dff_A_fbe2HY1E3_0),.clk(gclk));
	jdff dff_A_oPrjtPxO0_0(.dout(w_dff_A_fbe2HY1E3_0),.din(w_dff_A_oPrjtPxO0_0),.clk(gclk));
	jdff dff_A_Lhdn5QVK2_0(.dout(w_dff_A_oPrjtPxO0_0),.din(w_dff_A_Lhdn5QVK2_0),.clk(gclk));
	jdff dff_A_Rnby4Qjf5_0(.dout(w_dff_A_Lhdn5QVK2_0),.din(w_dff_A_Rnby4Qjf5_0),.clk(gclk));
	jdff dff_A_DUEzQ0Zt6_0(.dout(w_dff_A_Rnby4Qjf5_0),.din(w_dff_A_DUEzQ0Zt6_0),.clk(gclk));
	jdff dff_A_59tip4um6_0(.dout(w_dff_A_DUEzQ0Zt6_0),.din(w_dff_A_59tip4um6_0),.clk(gclk));
	jdff dff_A_JYr03RyS0_0(.dout(w_dff_A_59tip4um6_0),.din(w_dff_A_JYr03RyS0_0),.clk(gclk));
	jdff dff_A_3YAnqSFD0_0(.dout(w_dff_A_JYr03RyS0_0),.din(w_dff_A_3YAnqSFD0_0),.clk(gclk));
	jdff dff_A_ZPhOJqXE6_0(.dout(w_dff_A_3YAnqSFD0_0),.din(w_dff_A_ZPhOJqXE6_0),.clk(gclk));
	jdff dff_A_PmGAFBZK7_0(.dout(w_dff_A_ZPhOJqXE6_0),.din(w_dff_A_PmGAFBZK7_0),.clk(gclk));
	jdff dff_A_VBd96eJ74_0(.dout(w_dff_A_PmGAFBZK7_0),.din(w_dff_A_VBd96eJ74_0),.clk(gclk));
	jdff dff_A_GTlv67Vm9_2(.dout(God0),.din(w_dff_A_GTlv67Vm9_2),.clk(gclk));
	jdff dff_A_GSZfjr7J0_2(.dout(God1),.din(w_dff_A_GSZfjr7J0_2),.clk(gclk));
	jdff dff_A_uQkLPNWZ8_2(.dout(God2),.din(w_dff_A_uQkLPNWZ8_2),.clk(gclk));
	jdff dff_A_55Gbgj6p6_2(.dout(God3),.din(w_dff_A_55Gbgj6p6_2),.clk(gclk));
	jdff dff_A_B8wZr4MU3_2(.dout(God4),.din(w_dff_A_B8wZr4MU3_2),.clk(gclk));
	jdff dff_A_yRU2enKl6_2(.dout(God5),.din(w_dff_A_yRU2enKl6_2),.clk(gclk));
	jdff dff_A_Q05eg1e32_2(.dout(God6),.din(w_dff_A_Q05eg1e32_2),.clk(gclk));
	jdff dff_A_tI95YF7r3_2(.dout(God7),.din(w_dff_A_tI95YF7r3_2),.clk(gclk));
	jdff dff_A_M8cCqJfp6_2(.dout(God8),.din(w_dff_A_M8cCqJfp6_2),.clk(gclk));
	jdff dff_A_TN9CdVrU9_2(.dout(God9),.din(w_dff_A_TN9CdVrU9_2),.clk(gclk));
	jdff dff_A_SdT464Q11_2(.dout(God10),.din(w_dff_A_SdT464Q11_2),.clk(gclk));
	jdff dff_A_lnT3lzl99_2(.dout(God11),.din(w_dff_A_lnT3lzl99_2),.clk(gclk));
	jdff dff_A_7jbkq2NO0_2(.dout(God12),.din(w_dff_A_7jbkq2NO0_2),.clk(gclk));
	jdff dff_A_EIKtJcB52_2(.dout(God13),.din(w_dff_A_EIKtJcB52_2),.clk(gclk));
	jdff dff_A_5MddvVjy9_2(.dout(God14),.din(w_dff_A_5MddvVjy9_2),.clk(gclk));
	jdff dff_A_64k6T4eZ6_2(.dout(God15),.din(w_dff_A_64k6T4eZ6_2),.clk(gclk));
endmodule

