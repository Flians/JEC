// Benchmark "top" written by ABC on Thu May 28 22:00:58 2020

module gf_sin ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    sin0 , sin1 , sin2 , sin3 , sin4 , sin5 , sin6 ,
    sin7 , sin8 , sin9 , sin10 , sin11 , sin12 ,
    sin13 , sin14 , sin15 , sin16 , sin17 , sin18 ,
    sin19 , sin20 , sin21 , sin22 , sin23 , sin24   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ;
  output sin0 , sin1 , sin2 , sin3 , sin4 , sin5 , sin6 ,
    sin7 , sin8 , sin9 , sin10 , sin11 , sin12 ,
    sin13 , sin14 , sin15 , sin16 , sin17 , sin18 ,
    sin19 , sin20 , sin21 , sin22 , sin23 , sin24 ;
  wire n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
    n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
    n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
    n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
    n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
    n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
    n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
    n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
    n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
    n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
    n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
    n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
    n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
    n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
    n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
    n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
    n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
    n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4214, n4215, n4216, n4219, n4220, n4221, n4222, n4223, n4224,
    n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
    n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4716, n4717, n4718, n4719, n4720,
    n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
    n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
    n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
    n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
    n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
    n5004, n5005, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5116,
    n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
    n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
    n5208, n5209, n5210, n5211, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
    n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5381,
    n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
    n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
    n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
    n5455, n5456, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
    n5498, n5499, n5500, n5501, n5502, n5503;
  jnot g0000(.din(a22 ), .dout(n49));
  jor  g0001(.dina(a1 ), .dinb(a0 ), .dout(n50));
  jor  g0002(.dina(n50), .dinb(a2 ), .dout(n51));
  jor  g0003(.dina(n51), .dinb(a3 ), .dout(n52));
  jor  g0004(.dina(n52), .dinb(a4 ), .dout(n53));
  jor  g0005(.dina(n53), .dinb(a5 ), .dout(n54));
  jor  g0006(.dina(n54), .dinb(a6 ), .dout(n55));
  jor  g0007(.dina(n55), .dinb(a7 ), .dout(n56));
  jor  g0008(.dina(n56), .dinb(a8 ), .dout(n57));
  jor  g0009(.dina(n57), .dinb(a9 ), .dout(n58));
  jor  g0010(.dina(n58), .dinb(a10 ), .dout(n59));
  jor  g0011(.dina(n59), .dinb(a11 ), .dout(n60));
  jor  g0012(.dina(n60), .dinb(a12 ), .dout(n61));
  jor  g0013(.dina(n61), .dinb(a13 ), .dout(n62));
  jor  g0014(.dina(n62), .dinb(a14 ), .dout(n63));
  jor  g0015(.dina(n63), .dinb(a15 ), .dout(n64));
  jor  g0016(.dina(n64), .dinb(a16 ), .dout(n65));
  jor  g0017(.dina(n65), .dinb(a17 ), .dout(n66));
  jor  g0018(.dina(n66), .dinb(a18 ), .dout(n67));
  jor  g0019(.dina(n67), .dinb(a19 ), .dout(n68));
  jand g0020(.dina(n68), .dinb(n49), .dout(n69));
  jxor g0021(.dina(n69), .dinb(a20 ), .dout(n70));
  jnot g0022(.din(a21 ), .dout(n71));
  jor  g0023(.dina(n68), .dinb(a20 ), .dout(n72));
  jand g0024(.dina(n72), .dinb(n49), .dout(n73));
  jxor g0025(.dina(n73), .dinb(n71), .dout(n74));
  jor  g0026(.dina(n74), .dinb(n70), .dout(n75));
  jand g0027(.dina(n63), .dinb(n49), .dout(n76));
  jxor g0028(.dina(n76), .dinb(a15 ), .dout(n77));
  jor  g0029(.dina(n77), .dinb(n75), .dout(n78));
  jnot g0030(.din(a19 ), .dout(n79));
  jand g0031(.dina(n67), .dinb(n49), .dout(n80));
  jxor g0032(.dina(n80), .dinb(n79), .dout(n81));
  jand g0033(.dina(n66), .dinb(n49), .dout(n82));
  jxor g0034(.dina(n82), .dinb(a18 ), .dout(n83));
  jnot g0035(.din(n83), .dout(n84));
  jand g0036(.dina(n84), .dinb(n81), .dout(n85));
  jand g0037(.dina(n65), .dinb(n49), .dout(n86));
  jxor g0038(.dina(n86), .dinb(a17 ), .dout(n87));
  jnot g0039(.din(n87), .dout(n88));
  jand g0040(.dina(n64), .dinb(n49), .dout(n89));
  jxor g0041(.dina(n89), .dinb(a16 ), .dout(n90));
  jand g0042(.dina(n90), .dinb(n88), .dout(n91));
  jand g0043(.dina(n91), .dinb(n85), .dout(n92));
  jnot g0044(.din(n92), .dout(n93));
  jor  g0045(.dina(n93), .dinb(n78), .dout(n94));
  jxor g0046(.dina(n80), .dinb(a19 ), .dout(n95));
  jand g0047(.dina(n83), .dinb(n95), .dout(n96));
  jand g0048(.dina(n90), .dinb(n87), .dout(n97));
  jand g0049(.dina(n97), .dinb(n96), .dout(n98));
  jnot g0050(.din(n98), .dout(n99));
  jnot g0051(.din(n77), .dout(n100));
  jor  g0052(.dina(n100), .dinb(n75), .dout(n101));
  jor  g0053(.dina(n101), .dinb(n99), .dout(n102));
  jand g0054(.dina(n102), .dinb(n94), .dout(n103));
  jnot g0055(.din(a20 ), .dout(n104));
  jxor g0056(.dina(n69), .dinb(n104), .dout(n105));
  jxor g0057(.dina(n73), .dinb(a21 ), .dout(n106));
  jor  g0058(.dina(n106), .dinb(n105), .dout(n107));
  jor  g0059(.dina(n107), .dinb(n100), .dout(n108));
  jnot g0060(.din(n90), .dout(n109));
  jand g0061(.dina(n109), .dinb(n88), .dout(n110));
  jand g0062(.dina(n83), .dinb(n81), .dout(n111));
  jand g0063(.dina(n111), .dinb(n110), .dout(n112));
  jnot g0064(.din(n112), .dout(n113));
  jor  g0065(.dina(n113), .dinb(n108), .dout(n114));
  jand g0066(.dina(n109), .dinb(n87), .dout(n115));
  jand g0067(.dina(n115), .dinb(n96), .dout(n116));
  jand g0068(.dina(n74), .dinb(n105), .dout(n117));
  jand g0069(.dina(n117), .dinb(n100), .dout(n118));
  jand g0070(.dina(n118), .dinb(n116), .dout(n119));
  jnot g0071(.din(n119), .dout(n120));
  jand g0072(.dina(n120), .dinb(n114), .dout(n121));
  jand g0073(.dina(n121), .dinb(n103), .dout(n122));
  jnot g0074(.din(n116), .dout(n123));
  jor  g0075(.dina(n123), .dinb(n108), .dout(n124));
  jor  g0076(.dina(n107), .dinb(n77), .dout(n125));
  jand g0077(.dina(n111), .dinb(n91), .dout(n126));
  jnot g0078(.din(n126), .dout(n127));
  jor  g0079(.dina(n127), .dinb(n125), .dout(n128));
  jand g0080(.dina(n128), .dinb(n124), .dout(n129));
  jand g0081(.dina(n111), .dinb(n97), .dout(n130));
  jand g0082(.dina(n130), .dinb(n117), .dout(n131));
  jand g0083(.dina(n131), .dinb(n77), .dout(n132));
  jnot g0084(.din(n132), .dout(n133));
  jor  g0085(.dina(n74), .dinb(n105), .dout(n134));
  jor  g0086(.dina(n134), .dinb(n100), .dout(n135));
  jor  g0087(.dina(n135), .dinb(n123), .dout(n136));
  jand g0088(.dina(n136), .dinb(n133), .dout(n137));
  jor  g0089(.dina(n134), .dinb(n77), .dout(n138));
  jand g0090(.dina(n84), .dinb(n95), .dout(n139));
  jand g0091(.dina(n139), .dinb(n115), .dout(n140));
  jnot g0092(.din(n140), .dout(n141));
  jor  g0093(.dina(n141), .dinb(n138), .dout(n142));
  jand g0094(.dina(n106), .dinb(n70), .dout(n143));
  jand g0095(.dina(n143), .dinb(n100), .dout(n144));
  jand g0096(.dina(n139), .dinb(n97), .dout(n145));
  jand g0097(.dina(n145), .dinb(n144), .dout(n146));
  jnot g0098(.din(n146), .dout(n147));
  jand g0099(.dina(n147), .dinb(n142), .dout(n148));
  jand g0100(.dina(n148), .dinb(n137), .dout(n149));
  jand g0101(.dina(n149), .dinb(n129), .dout(n150));
  jnot g0102(.din(n130), .dout(n151));
  jor  g0103(.dina(n135), .dinb(n151), .dout(n152));
  jand g0104(.dina(n152), .dinb(n150), .dout(n153));
  jand g0105(.dina(n143), .dinb(n77), .dout(n154));
  jand g0106(.dina(n139), .dinb(n91), .dout(n155));
  jand g0107(.dina(n155), .dinb(n154), .dout(n156));
  jnot g0108(.din(n156), .dout(n157));
  jor  g0109(.dina(n125), .dinb(n123), .dout(n158));
  jor  g0110(.dina(n123), .dinb(n75), .dout(n159));
  jor  g0111(.dina(n159), .dinb(n100), .dout(n160));
  jand g0112(.dina(n160), .dinb(n158), .dout(n161));
  jor  g0113(.dina(n138), .dinb(n151), .dout(n162));
  jand g0114(.dina(n162), .dinb(n161), .dout(n163));
  jand g0115(.dina(n163), .dinb(n157), .dout(n164));
  jnot g0116(.din(n155), .dout(n165));
  jor  g0117(.dina(n165), .dinb(n138), .dout(n166));
  jand g0118(.dina(n115), .dinb(n111), .dout(n167));
  jnot g0119(.din(n167), .dout(n168));
  jor  g0120(.dina(n168), .dinb(n138), .dout(n169));
  jand g0121(.dina(n169), .dinb(n166), .dout(n170));
  jand g0122(.dina(n96), .dinb(n91), .dout(n171));
  jand g0123(.dina(n171), .dinb(n144), .dout(n172));
  jnot g0124(.din(n172), .dout(n173));
  jand g0125(.dina(n117), .dinb(n77), .dout(n174));
  jand g0126(.dina(n174), .dinb(n167), .dout(n175));
  jnot g0127(.din(n175), .dout(n176));
  jand g0128(.dina(n176), .dinb(n173), .dout(n177));
  jand g0129(.dina(n177), .dinb(n170), .dout(n178));
  jand g0130(.dina(n178), .dinb(n164), .dout(n179));
  jand g0131(.dina(n179), .dinb(n153), .dout(n180));
  jand g0132(.dina(n180), .dinb(n122), .dout(n181));
  jor  g0133(.dina(n168), .dinb(n101), .dout(n182));
  jand g0134(.dina(n74), .dinb(n70), .dout(n183));
  jand g0135(.dina(n183), .dinb(n77), .dout(n184));
  jand g0136(.dina(n115), .dinb(n85), .dout(n185));
  jand g0137(.dina(n185), .dinb(n184), .dout(n186));
  jnot g0138(.din(n186), .dout(n187));
  jor  g0139(.dina(n138), .dinb(n127), .dout(n188));
  jand g0140(.dina(n188), .dinb(n187), .dout(n189));
  jand g0141(.dina(n189), .dinb(n182), .dout(n190));
  jor  g0142(.dina(n138), .dinb(n123), .dout(n191));
  jand g0143(.dina(n139), .dinb(n110), .dout(n192));
  jnot g0144(.din(n192), .dout(n193));
  jor  g0145(.dina(n193), .dinb(n75), .dout(n194));
  jor  g0146(.dina(n194), .dinb(n77), .dout(n195));
  jand g0147(.dina(n118), .dinb(n92), .dout(n196));
  jnot g0148(.din(n196), .dout(n197));
  jand g0149(.dina(n197), .dinb(n195), .dout(n198));
  jand g0150(.dina(n198), .dinb(n191), .dout(n199));
  jand g0151(.dina(n199), .dinb(n190), .dout(n200));
  jor  g0152(.dina(n84), .dinb(n81), .dout(n201));
  jnot g0153(.din(n110), .dout(n202));
  jor  g0154(.dina(n202), .dinb(n201), .dout(n203));
  jor  g0155(.dina(n203), .dinb(n125), .dout(n204));
  jand g0156(.dina(n140), .dinb(n154), .dout(n205));
  jnot g0157(.din(n205), .dout(n206));
  jor  g0158(.dina(n193), .dinb(n125), .dout(n207));
  jand g0159(.dina(n207), .dinb(n206), .dout(n208));
  jand g0160(.dina(n208), .dinb(n204), .dout(n209));
  jand g0161(.dina(n209), .dinb(n200), .dout(n210));
  jand g0162(.dina(n210), .dinb(n181), .dout(n211));
  jand g0163(.dina(n140), .dinb(n184), .dout(n212));
  jnot g0164(.din(n212), .dout(n213));
  jand g0165(.dina(n145), .dinb(n154), .dout(n214));
  jnot g0166(.din(n214), .dout(n215));
  jor  g0167(.dina(n106), .dinb(n70), .dout(n216));
  jor  g0168(.dina(n216), .dinb(n100), .dout(n217));
  jor  g0169(.dina(n217), .dinb(n165), .dout(n218));
  jand g0170(.dina(n218), .dinb(n215), .dout(n219));
  jand g0171(.dina(n219), .dinb(n213), .dout(n220));
  jor  g0172(.dina(n193), .dinb(n135), .dout(n221));
  jor  g0173(.dina(n159), .dinb(n77), .dout(n222));
  jand g0174(.dina(n106), .dinb(n105), .dout(n223));
  jand g0175(.dina(n77), .dinb(n223), .dout(n224));
  jand g0176(.dina(n171), .dinb(n224), .dout(n225));
  jnot g0177(.din(n225), .dout(n226));
  jand g0178(.dina(n226), .dinb(n222), .dout(n227));
  jand g0179(.dina(n227), .dinb(n221), .dout(n228));
  jand g0180(.dina(n228), .dinb(n220), .dout(n229));
  jand g0181(.dina(n97), .dinb(n85), .dout(n230));
  jnot g0182(.din(n230), .dout(n231));
  jor  g0183(.dina(n231), .dinb(n135), .dout(n232));
  jor  g0184(.dina(n138), .dinb(n93), .dout(n233));
  jand g0185(.dina(n233), .dinb(n232), .dout(n234));
  jor  g0186(.dina(n135), .dinb(n127), .dout(n235));
  jor  g0187(.dina(n168), .dinb(n135), .dout(n236));
  jand g0188(.dina(n236), .dinb(n235), .dout(n237));
  jor  g0189(.dina(n127), .dinb(n101), .dout(n238));
  jand g0190(.dina(n174), .dinb(n112), .dout(n239));
  jnot g0191(.din(n239), .dout(n240));
  jand g0192(.dina(n240), .dinb(n238), .dout(n241));
  jand g0193(.dina(n241), .dinb(n237), .dout(n242));
  jand g0194(.dina(n242), .dinb(n234), .dout(n243));
  jor  g0195(.dina(n231), .dinb(n108), .dout(n244));
  jor  g0196(.dina(n217), .dinb(n123), .dout(n245));
  jand g0197(.dina(n245), .dinb(n244), .dout(n246));
  jand g0198(.dina(n230), .dinb(n174), .dout(n247));
  jnot g0199(.din(n247), .dout(n248));
  jnot g0200(.din(n185), .dout(n249));
  jor  g0201(.dina(n249), .dinb(n217), .dout(n250));
  jand g0202(.dina(n250), .dinb(n248), .dout(n251));
  jor  g0203(.dina(n203), .dinb(n78), .dout(n252));
  jand g0204(.dina(n183), .dinb(n100), .dout(n253));
  jand g0205(.dina(n140), .dinb(n253), .dout(n254));
  jnot g0206(.din(n254), .dout(n255));
  jand g0207(.dina(n255), .dinb(n252), .dout(n256));
  jand g0208(.dina(n256), .dinb(n251), .dout(n257));
  jand g0209(.dina(n257), .dinb(n246), .dout(n258));
  jand g0210(.dina(n258), .dinb(n243), .dout(n259));
  jand g0211(.dina(n259), .dinb(n229), .dout(n260));
  jor  g0212(.dina(n217), .dinb(n127), .dout(n261));
  jand g0213(.dina(n100), .dinb(n223), .dout(n262));
  jand g0214(.dina(n110), .dinb(n85), .dout(n263));
  jand g0215(.dina(n263), .dinb(n262), .dout(n264));
  jnot g0216(.din(n264), .dout(n265));
  jand g0217(.dina(n184), .dinb(n98), .dout(n266));
  jnot g0218(.din(n266), .dout(n267));
  jnot g0219(.din(n263), .dout(n268));
  jor  g0220(.dina(n268), .dinb(n135), .dout(n269));
  jand g0221(.dina(n269), .dinb(n267), .dout(n270));
  jand g0222(.dina(n270), .dinb(n265), .dout(n271));
  jand g0223(.dina(n271), .dinb(n261), .dout(n272));
  jand g0224(.dina(n272), .dinb(n260), .dout(n273));
  jand g0225(.dina(n145), .dinb(n118), .dout(n274));
  jnot g0226(.din(n274), .dout(n275));
  jor  g0227(.dina(n165), .dinb(n108), .dout(n276));
  jand g0228(.dina(n276), .dinb(n275), .dout(n277));
  jor  g0229(.dina(n113), .dinb(n78), .dout(n278));
  jor  g0230(.dina(n203), .dinb(n134), .dout(n279));
  jor  g0231(.dina(n279), .dinb(n77), .dout(n280));
  jand g0232(.dina(n280), .dinb(n278), .dout(n281));
  jand g0233(.dina(n145), .dinb(n262), .dout(n282));
  jnot g0234(.din(n282), .dout(n283));
  jand g0235(.dina(n283), .dinb(n281), .dout(n284));
  jand g0236(.dina(n284), .dinb(n277), .dout(n285));
  jor  g0237(.dina(n279), .dinb(n100), .dout(n286));
  jand g0238(.dina(n263), .dinb(n184), .dout(n287));
  jnot g0239(.din(n287), .dout(n288));
  jnot g0240(.din(n171), .dout(n289));
  jor  g0241(.dina(n289), .dinb(n135), .dout(n290));
  jand g0242(.dina(n290), .dinb(n288), .dout(n291));
  jand g0243(.dina(n291), .dinb(n286), .dout(n292));
  jand g0244(.dina(n292), .dinb(n285), .dout(n293));
  jor  g0245(.dina(n138), .dinb(n99), .dout(n294));
  jand g0246(.dina(n140), .dinb(n223), .dout(n295));
  jand g0247(.dina(n295), .dinb(n77), .dout(n296));
  jnot g0248(.din(n296), .dout(n297));
  jand g0249(.dina(n297), .dinb(n294), .dout(n298));
  jand g0250(.dina(n154), .dinb(n92), .dout(n299));
  jnot g0251(.din(n299), .dout(n300));
  jand g0252(.dina(n145), .dinb(n183), .dout(n301));
  jand g0253(.dina(n301), .dinb(n100), .dout(n302));
  jnot g0254(.din(n302), .dout(n303));
  jand g0255(.dina(n303), .dinb(n300), .dout(n304));
  jor  g0256(.dina(n113), .dinb(n101), .dout(n305));
  jand g0257(.dina(n305), .dinb(n304), .dout(n306));
  jand g0258(.dina(n306), .dinb(n298), .dout(n307));
  jand g0259(.dina(n145), .dinb(n224), .dout(n308));
  jnot g0260(.din(n308), .dout(n309));
  jor  g0261(.dina(n289), .dinb(n125), .dout(n310));
  jand g0262(.dina(n110), .dinb(n96), .dout(n311));
  jand g0263(.dina(n311), .dinb(n224), .dout(n312));
  jnot g0264(.din(n312), .dout(n313));
  jand g0265(.dina(n230), .dinb(n144), .dout(n314));
  jnot g0266(.din(n314), .dout(n315));
  jand g0267(.dina(n315), .dinb(n313), .dout(n316));
  jand g0268(.dina(n316), .dinb(n310), .dout(n317));
  jand g0269(.dina(n317), .dinb(n309), .dout(n318));
  jand g0270(.dina(n318), .dinb(n307), .dout(n319));
  jand g0271(.dina(n319), .dinb(n293), .dout(n320));
  jor  g0272(.dina(n165), .dinb(n101), .dout(n321));
  jand g0273(.dina(n321), .dinb(n320), .dout(n322));
  jand g0274(.dina(n322), .dinb(n273), .dout(n323));
  jand g0275(.dina(n323), .dinb(n211), .dout(n324));
  jnot g0276(.din(n324), .dout(n325));
  jand g0277(.dina(n294), .dinb(n191), .dout(n326));
  jor  g0278(.dina(n289), .dinb(n108), .dout(n327));
  jand g0279(.dina(n327), .dinb(n280), .dout(n328));
  jand g0280(.dina(n328), .dinb(n326), .dout(n329));
  jand g0281(.dina(n253), .dinb(n92), .dout(n330));
  jnot g0282(.din(n330), .dout(n331));
  jor  g0283(.dina(n168), .dinb(n78), .dout(n332));
  jor  g0284(.dina(n108), .dinb(n93), .dout(n333));
  jand g0285(.dina(n333), .dinb(n332), .dout(n334));
  jand g0286(.dina(n334), .dinb(n331), .dout(n335));
  jor  g0287(.dina(n216), .dinb(n77), .dout(n336));
  jor  g0288(.dina(n168), .dinb(n336), .dout(n337));
  jand g0289(.dina(n337), .dinb(n250), .dout(n338));
  jor  g0290(.dina(n193), .dinb(n108), .dout(n339));
  jand g0291(.dina(n339), .dinb(n176), .dout(n340));
  jand g0292(.dina(n340), .dinb(n133), .dout(n341));
  jand g0293(.dina(n341), .dinb(n338), .dout(n342));
  jand g0294(.dina(n342), .dinb(n335), .dout(n343));
  jor  g0295(.dina(n203), .dinb(n108), .dout(n344));
  jand g0296(.dina(n269), .dinb(n188), .dout(n345));
  jor  g0297(.dina(n268), .dinb(n125), .dout(n346));
  jor  g0298(.dina(n268), .dinb(n138), .dout(n347));
  jand g0299(.dina(n347), .dinb(n346), .dout(n348));
  jand g0300(.dina(n348), .dinb(n345), .dout(n349));
  jand g0301(.dina(n349), .dinb(n344), .dout(n350));
  jand g0302(.dina(n305), .dinb(n238), .dout(n351));
  jand g0303(.dina(n351), .dinb(n288), .dout(n352));
  jor  g0304(.dina(n127), .dinb(n108), .dout(n353));
  jand g0305(.dina(n353), .dinb(n195), .dout(n354));
  jand g0306(.dina(n354), .dinb(n161), .dout(n355));
  jand g0307(.dina(n355), .dinb(n352), .dout(n356));
  jand g0308(.dina(n356), .dinb(n350), .dout(n357));
  jand g0309(.dina(n357), .dinb(n343), .dout(n358));
  jand g0310(.dina(n358), .dinb(n329), .dout(n359));
  jand g0311(.dina(n171), .dinb(n262), .dout(n360));
  jnot g0312(.din(n360), .dout(n361));
  jand g0313(.dina(n361), .dinb(n120), .dout(n362));
  jand g0314(.dina(n117), .dinb(n112), .dout(n363));
  jor  g0315(.dina(n363), .dinb(n302), .dout(n364));
  jnot g0316(.din(n364), .dout(n365));
  jor  g0317(.dina(n249), .dinb(n125), .dout(n366));
  jand g0318(.dina(n366), .dinb(n297), .dout(n367));
  jand g0319(.dina(n367), .dinb(n365), .dout(n368));
  jand g0320(.dina(n368), .dinb(n362), .dout(n369));
  jor  g0321(.dina(n135), .dinb(n99), .dout(n370));
  jand g0322(.dina(n215), .dinb(n206), .dout(n371));
  jand g0323(.dina(n371), .dinb(n370), .dout(n372));
  jor  g0324(.dina(n231), .dinb(n75), .dout(n373));
  jor  g0325(.dina(n373), .dinb(n100), .dout(n374));
  jand g0326(.dina(n374), .dinb(n207), .dout(n375));
  jand g0327(.dina(n375), .dinb(n372), .dout(n376));
  jor  g0328(.dina(n138), .dinb(n113), .dout(n377));
  jor  g0329(.dina(n165), .dinb(n78), .dout(n378));
  jand g0330(.dina(n378), .dinb(n377), .dout(n379));
  jand g0331(.dina(n236), .dinb(n162), .dout(n380));
  jand g0332(.dina(n380), .dinb(n379), .dout(n381));
  jor  g0333(.dina(n168), .dinb(n108), .dout(n382));
  jor  g0334(.dina(n165), .dinb(n336), .dout(n383));
  jor  g0335(.dina(n151), .dinb(n101), .dout(n384));
  jand g0336(.dina(n384), .dinb(n383), .dout(n385));
  jand g0337(.dina(n385), .dinb(n382), .dout(n386));
  jor  g0338(.dina(n268), .dinb(n101), .dout(n387));
  jand g0339(.dina(n387), .dinb(n310), .dout(n388));
  jor  g0340(.dina(n127), .dinb(n336), .dout(n389));
  jand g0341(.dina(n389), .dinb(n218), .dout(n390));
  jand g0342(.dina(n390), .dinb(n388), .dout(n391));
  jand g0343(.dina(n391), .dinb(n386), .dout(n392));
  jand g0344(.dina(n392), .dinb(n381), .dout(n393));
  jand g0345(.dina(n393), .dinb(n376), .dout(n394));
  jor  g0346(.dina(n217), .dinb(n93), .dout(n395));
  jand g0347(.dina(n395), .dinb(n321), .dout(n396));
  jand g0348(.dina(n396), .dinb(n255), .dout(n397));
  jand g0349(.dina(n397), .dinb(n309), .dout(n398));
  jand g0350(.dina(n311), .dinb(n118), .dout(n399));
  jand g0351(.dina(n263), .dinb(n174), .dout(n400));
  jor  g0352(.dina(n400), .dinb(n399), .dout(n401));
  jnot g0353(.din(n401), .dout(n402));
  jor  g0354(.dina(n141), .dinb(n75), .dout(n403));
  jor  g0355(.dina(n403), .dinb(n77), .dout(n404));
  jand g0356(.dina(n404), .dinb(n233), .dout(n405));
  jand g0357(.dina(n405), .dinb(n283), .dout(n406));
  jand g0358(.dina(n406), .dinb(n402), .dout(n407));
  jand g0359(.dina(n407), .dinb(n398), .dout(n408));
  jor  g0360(.dina(n165), .dinb(n125), .dout(n409));
  jand g0361(.dina(n171), .dinb(n118), .dout(n410));
  jnot g0362(.din(n410), .dout(n411));
  jand g0363(.dina(n411), .dinb(n409), .dout(n412));
  jand g0364(.dina(n230), .dinb(n223), .dout(n413));
  jand g0365(.dina(n413), .dinb(n100), .dout(n414));
  jnot g0366(.din(n414), .dout(n415));
  jand g0367(.dina(n415), .dinb(n286), .dout(n416));
  jand g0368(.dina(n416), .dinb(n412), .dout(n417));
  jor  g0369(.dina(n249), .dinb(n101), .dout(n418));
  jand g0370(.dina(n226), .dinb(n94), .dout(n419));
  jand g0371(.dina(n419), .dinb(n418), .dout(n420));
  jand g0372(.dina(n420), .dinb(n417), .dout(n421));
  jand g0373(.dina(n421), .dinb(n408), .dout(n422));
  jand g0374(.dina(n422), .dinb(n394), .dout(n423));
  jand g0375(.dina(n423), .dinb(n369), .dout(n424));
  jand g0376(.dina(n424), .dinb(n359), .dout(n425));
  jand g0377(.dina(n140), .dinb(n118), .dout(n426));
  jnot g0378(.din(n426), .dout(n427));
  jand g0379(.dina(n411), .dinb(n120), .dout(n428));
  jor  g0380(.dina(n127), .dinb(n78), .dout(n429));
  jand g0381(.dina(n429), .dinb(n278), .dout(n430));
  jand g0382(.dina(n430), .dinb(n428), .dout(n431));
  jand g0383(.dina(n431), .dinb(n352), .dout(n432));
  jand g0384(.dina(n311), .dinb(n174), .dout(n433));
  jnot g0385(.din(n433), .dout(n434));
  jor  g0386(.dina(n217), .dinb(n289), .dout(n435));
  jand g0387(.dina(n435), .dinb(n434), .dout(n436));
  jand g0388(.dina(n346), .dinb(n245), .dout(n437));
  jor  g0389(.dina(n217), .dinb(n99), .dout(n438));
  jor  g0390(.dina(n336), .dinb(n99), .dout(n439));
  jand g0391(.dina(n439), .dinb(n438), .dout(n440));
  jand g0392(.dina(n440), .dinb(n437), .dout(n441));
  jand g0393(.dina(n441), .dinb(n436), .dout(n442));
  jand g0394(.dina(n442), .dinb(n432), .dout(n443));
  jnot g0395(.din(n145), .dout(n444));
  jor  g0396(.dina(n217), .dinb(n444), .dout(n445));
  jnot g0397(.din(n399), .dout(n446));
  jand g0398(.dina(n174), .dinb(n140), .dout(n447));
  jnot g0399(.din(n447), .dout(n448));
  jand g0400(.dina(n448), .dinb(n446), .dout(n449));
  jand g0401(.dina(n449), .dinb(n445), .dout(n450));
  jand g0402(.dina(n450), .dinb(n275), .dout(n451));
  jand g0403(.dina(n451), .dinb(n443), .dout(n452));
  jand g0404(.dina(n452), .dinb(n427), .dout(n453));
  jnot g0405(.din(n453), .dout(n454));
  jand g0406(.dina(n344), .dinb(n327), .dout(n455));
  jand g0407(.dina(n455), .dinb(n310), .dout(n456));
  jnot g0408(.din(n301), .dout(n457));
  jand g0409(.dina(n457), .dinb(n124), .dout(n458));
  jand g0410(.dina(n458), .dinb(n456), .dout(n459));
  jor  g0411(.dina(n101), .dinb(n93), .dout(n460));
  jand g0412(.dina(n460), .dinb(n418), .dout(n461));
  jor  g0413(.dina(n249), .dinb(n78), .dout(n462));
  jand g0414(.dina(n462), .dinb(n374), .dout(n463));
  jand g0415(.dina(n463), .dinb(n461), .dout(n464));
  jand g0416(.dina(n464), .dinb(n459), .dout(n465));
  jnot g0417(.din(n465), .dout(n466));
  jor  g0418(.dina(n125), .dinb(n99), .dout(n467));
  jand g0419(.dina(n467), .dinb(n332), .dout(n468));
  jnot g0420(.din(n468), .dout(n469));
  jand g0421(.dina(n311), .dinb(n253), .dout(n470));
  jand g0422(.dina(n263), .dinb(n223), .dout(n471));
  jor  g0423(.dina(n471), .dinb(n470), .dout(n472));
  jor  g0424(.dina(n472), .dinb(n469), .dout(n473));
  jand g0425(.dina(n158), .dinb(n94), .dout(n474));
  jand g0426(.dina(n415), .dinb(n267), .dout(n475));
  jand g0427(.dina(n475), .dinb(n213), .dout(n476));
  jand g0428(.dina(n476), .dinb(n474), .dout(n477));
  jnot g0429(.din(n477), .dout(n478));
  jor  g0430(.dina(n478), .dinb(n473), .dout(n479));
  jor  g0431(.dina(n479), .dinb(n466), .dout(n480));
  jor  g0432(.dina(n193), .dinb(n217), .dout(n481));
  jand g0433(.dina(n481), .dinb(n218), .dout(n482));
  jand g0434(.dina(n482), .dinb(n383), .dout(n483));
  jnot g0435(.din(n483), .dout(n484));
  jor  g0436(.dina(n484), .dinb(n480), .dout(n485));
  jor  g0437(.dina(n485), .dinb(n454), .dout(n486));
  jand g0438(.dina(n167), .dinb(n253), .dout(n487));
  jnot g0439(.din(n487), .dout(n488));
  jor  g0440(.dina(n151), .dinb(n125), .dout(n489));
  jand g0441(.dina(n489), .dinb(n353), .dout(n490));
  jand g0442(.dina(n490), .dinb(n488), .dout(n491));
  jand g0443(.dina(n409), .dinb(n207), .dout(n492));
  jand g0444(.dina(n339), .dinb(n276), .dout(n493));
  jand g0445(.dina(n493), .dinb(n492), .dout(n494));
  jand g0446(.dina(n130), .dinb(n184), .dout(n495));
  jor  g0447(.dina(n495), .dinb(n254), .dout(n496));
  jnot g0448(.din(n496), .dout(n497));
  jand g0449(.dina(n497), .dinb(n382), .dout(n498));
  jand g0450(.dina(n498), .dinb(n494), .dout(n499));
  jand g0451(.dina(n499), .dinb(n491), .dout(n500));
  jand g0452(.dina(n430), .dinb(n351), .dout(n501));
  jand g0453(.dina(n501), .dinb(n500), .dout(n502));
  jnot g0454(.din(n502), .dout(n503));
  jor  g0455(.dina(n503), .dinb(n480), .dout(n504));
  jand g0456(.dina(n366), .dinb(n331), .dout(n505));
  jor  g0457(.dina(n231), .dinb(n125), .dout(n506));
  jand g0458(.dina(n506), .dinb(n333), .dout(n507));
  jand g0459(.dina(n507), .dinb(n114), .dout(n508));
  jand g0460(.dina(n508), .dinb(n505), .dout(n509));
  jor  g0461(.dina(n125), .dinb(n113), .dout(n510));
  jand g0462(.dina(n244), .dinb(n187), .dout(n511));
  jand g0463(.dina(n511), .dinb(n510), .dout(n512));
  jand g0464(.dina(n512), .dinb(n509), .dout(n513));
  jand g0465(.dina(n513), .dinb(n128), .dout(n514));
  jnot g0466(.din(n514), .dout(n515));
  jor  g0467(.dina(n515), .dinb(n504), .dout(n516));
  jxor g0468(.dina(n516), .dinb(n486), .dout(n517));
  jand g0469(.dina(n51), .dinb(n49), .dout(n518));
  jxor g0470(.dina(n518), .dinb(a3 ), .dout(n519));
  jand g0471(.dina(n519), .dinb(n517), .dout(n520));
  jnot g0472(.din(n520), .dout(n521));
  jand g0473(.dina(n388), .dinb(n250), .dout(n522));
  jand g0474(.dina(n253), .dinb(n116), .dout(n523));
  jor  g0475(.dina(n172), .dinb(n523), .dout(n524));
  jnot g0476(.din(n524), .dout(n525));
  jor  g0477(.dina(n151), .dinb(n216), .dout(n526));
  jor  g0478(.dina(n526), .dinb(n77), .dout(n527));
  jand g0479(.dina(n527), .dinb(n445), .dout(n528));
  jand g0480(.dina(n528), .dinb(n525), .dout(n529));
  jand g0481(.dina(n529), .dinb(n522), .dout(n530));
  jand g0482(.dina(n333), .dinb(n147), .dout(n531));
  jand g0483(.dina(n531), .dinb(n294), .dout(n532));
  jand g0484(.dina(n532), .dinb(n530), .dout(n533));
  jor  g0485(.dina(n99), .dinb(n78), .dout(n534));
  jor  g0486(.dina(n249), .dinb(n135), .dout(n535));
  jand g0487(.dina(n191), .dinb(n182), .dout(n536));
  jand g0488(.dina(n536), .dinb(n535), .dout(n537));
  jand g0489(.dina(n537), .dinb(n534), .dout(n538));
  jand g0490(.dina(n384), .dinb(n235), .dout(n539));
  jand g0491(.dina(n506), .dinb(n207), .dout(n540));
  jand g0492(.dina(n540), .dinb(n539), .dout(n541));
  jand g0493(.dina(n541), .dinb(n267), .dout(n542));
  jand g0494(.dina(n542), .dinb(n538), .dout(n543));
  jor  g0495(.dina(n495), .dinb(n312), .dout(n544));
  jnot g0496(.din(n544), .dout(n545));
  jand g0497(.dina(n382), .dinb(n204), .dout(n546));
  jand g0498(.dina(n546), .dinb(n133), .dout(n547));
  jand g0499(.dina(n547), .dinb(n545), .dout(n548));
  jand g0500(.dina(n548), .dinb(n407), .dout(n549));
  jand g0501(.dina(n549), .dinb(n543), .dout(n550));
  jand g0502(.dina(n550), .dinb(n533), .dout(n551));
  jand g0503(.dina(n331), .dinb(n114), .dout(n552));
  jand g0504(.dina(n112), .dinb(n262), .dout(n553));
  jor  g0505(.dina(n433), .dinb(n553), .dout(n554));
  jor  g0506(.dina(n554), .dinb(n296), .dout(n555));
  jnot g0507(.din(n555), .dout(n556));
  jand g0508(.dina(n269), .dinb(n252), .dout(n557));
  jand g0509(.dina(n395), .dinb(n160), .dout(n558));
  jand g0510(.dina(n558), .dinb(n557), .dout(n559));
  jand g0511(.dina(n559), .dinb(n556), .dout(n560));
  jor  g0512(.dina(n268), .dinb(n336), .dout(n561));
  jand g0513(.dina(n561), .dinb(n321), .dout(n562));
  jand g0514(.dina(n562), .dinb(n197), .dout(n563));
  jand g0515(.dina(n563), .dinb(n560), .dout(n564));
  jand g0516(.dina(n564), .dinb(n552), .dout(n565));
  jand g0517(.dina(n565), .dinb(n551), .dout(n566));
  jand g0518(.dina(n370), .dinb(n303), .dout(n567));
  jand g0519(.dina(n567), .dinb(n245), .dout(n568));
  jor  g0520(.dina(n135), .dinb(n113), .dout(n569));
  jor  g0521(.dina(n193), .dinb(n336), .dout(n570));
  jand g0522(.dina(n570), .dinb(n569), .dout(n571));
  jand g0523(.dina(n571), .dinb(n136), .dout(n572));
  jand g0524(.dina(n572), .dinb(n102), .dout(n573));
  jand g0525(.dina(n573), .dinb(n568), .dout(n574));
  jand g0526(.dina(n194), .dinb(n152), .dout(n575));
  jnot g0527(.din(n575), .dout(n576));
  jand g0528(.dina(n230), .dinb(n118), .dout(n577));
  jor  g0529(.dina(n577), .dinb(n205), .dout(n578));
  jand g0530(.dina(n118), .dinb(n98), .dout(n579));
  jor  g0531(.dina(n579), .dinb(n254), .dout(n580));
  jor  g0532(.dina(n580), .dinb(n578), .dout(n581));
  jor  g0533(.dina(n581), .dinb(n576), .dout(n582));
  jnot g0534(.din(n582), .dout(n583));
  jand g0535(.dina(n481), .dinb(n462), .dout(n584));
  jand g0536(.dina(n467), .dinb(n383), .dout(n585));
  jand g0537(.dina(n585), .dinb(n584), .dout(n586));
  jor  g0538(.dina(n151), .dinb(n78), .dout(n587));
  jand g0539(.dina(n587), .dinb(n166), .dout(n588));
  jand g0540(.dina(n232), .dinb(n128), .dout(n589));
  jand g0541(.dina(n589), .dinb(n588), .dout(n590));
  jand g0542(.dina(n590), .dinb(n586), .dout(n591));
  jand g0543(.dina(n438), .dinb(n244), .dout(n592));
  jand g0544(.dina(n592), .dinb(n248), .dout(n593));
  jand g0545(.dina(n409), .dinb(n290), .dout(n594));
  jand g0546(.dina(n594), .dinb(n378), .dout(n595));
  jand g0547(.dina(n595), .dinb(n593), .dout(n596));
  jand g0548(.dina(n596), .dinb(n591), .dout(n597));
  jand g0549(.dina(n597), .dinb(n583), .dout(n598));
  jand g0550(.dina(n185), .dinb(n118), .dout(n599));
  jnot g0551(.din(n599), .dout(n600));
  jand g0552(.dina(n600), .dinb(n418), .dout(n601));
  jand g0553(.dina(n309), .dinb(n236), .dout(n602));
  jand g0554(.dina(n602), .dinb(n305), .dout(n603));
  jand g0555(.dina(n603), .dinb(n601), .dout(n604));
  jand g0556(.dina(n604), .dinb(n598), .dout(n605));
  jand g0557(.dina(n605), .dinb(n574), .dout(n606));
  jand g0558(.dina(n606), .dinb(n566), .dout(n607));
  jnot g0559(.din(n417), .dout(n608));
  jand g0560(.dina(n192), .dinb(n154), .dout(n609));
  jand g0561(.dina(n154), .dinb(n98), .dout(n610));
  jor  g0562(.dina(n610), .dinb(n609), .dout(n611));
  jand g0563(.dina(n144), .dinb(n92), .dout(n612));
  jand g0564(.dina(n144), .dinb(n112), .dout(n613));
  jor  g0565(.dina(n613), .dinb(n612), .dout(n614));
  jor  g0566(.dina(n614), .dinb(n611), .dout(n615));
  jor  g0567(.dina(n615), .dinb(n360), .dout(n616));
  jand g0568(.dina(n144), .dinb(n98), .dout(n617));
  jand g0569(.dina(n116), .dinb(n184), .dout(n618));
  jand g0570(.dina(n126), .dinb(n253), .dout(n619));
  jor  g0571(.dina(n619), .dinb(n618), .dout(n620));
  jor  g0572(.dina(n266), .dinb(n620), .dout(n621));
  jor  g0573(.dina(n621), .dinb(n617), .dout(n622));
  jor  g0574(.dina(n622), .dinb(n616), .dout(n623));
  jand g0575(.dina(n116), .dinb(n223), .dout(n624));
  jand g0576(.dina(n624), .dinb(n100), .dout(n625));
  jand g0577(.dina(n263), .dinb(n224), .dout(n626));
  jor  g0578(.dina(n626), .dinb(n625), .dout(n627));
  jor  g0579(.dina(n627), .dinb(n599), .dout(n628));
  jor  g0580(.dina(n628), .dinb(n447), .dout(n629));
  jand g0581(.dina(n167), .dinb(n262), .dout(n630));
  jand g0582(.dina(n184), .dinb(n92), .dout(n631));
  jor  g0583(.dina(n631), .dinb(n630), .dout(n632));
  jor  g0584(.dina(n632), .dinb(n330), .dout(n633));
  jand g0585(.dina(n130), .dinb(n262), .dout(n634));
  jor  g0586(.dina(n634), .dinb(n633), .dout(n635));
  jor  g0587(.dina(n635), .dinb(n629), .dout(n636));
  jor  g0588(.dina(n636), .dinb(n623), .dout(n637));
  jor  g0589(.dina(n637), .dinb(n608), .dout(n638));
  jand g0590(.dina(n174), .dinb(n116), .dout(n639));
  jand g0591(.dina(n112), .dinb(n184), .dout(n640));
  jor  g0592(.dina(n295), .dinb(n640), .dout(n641));
  jor  g0593(.dina(n641), .dinb(n639), .dout(n642));
  jor  g0594(.dina(n642), .dinb(n301), .dout(n643));
  jor  g0595(.dina(n643), .dinb(n212), .dout(n644));
  jand g0596(.dina(n413), .dinb(n77), .dout(n645));
  jand g0597(.dina(n185), .dinb(n262), .dout(n646));
  jor  g0598(.dina(n646), .dinb(n645), .dout(n647));
  jand g0599(.dina(n185), .dinb(n253), .dout(n648));
  jor  g0600(.dina(n495), .dinb(n648), .dout(n649));
  jor  g0601(.dina(n649), .dinb(n647), .dout(n650));
  jand g0602(.dina(n311), .dinb(n262), .dout(n651));
  jand g0603(.dina(n263), .dinb(n154), .dout(n652));
  jor  g0604(.dina(n652), .dinb(n651), .dout(n653));
  jand g0605(.dina(n171), .dinb(n154), .dout(n654));
  jand g0606(.dina(n192), .dinb(n174), .dout(n655));
  jor  g0607(.dina(n655), .dinb(n654), .dout(n656));
  jor  g0608(.dina(n656), .dinb(n400), .dout(n657));
  jor  g0609(.dina(n657), .dinb(n653), .dout(n658));
  jor  g0610(.dina(n658), .dinb(n650), .dout(n659));
  jand g0611(.dina(n167), .dinb(n184), .dout(n660));
  jor  g0612(.dina(n660), .dinb(n470), .dout(n661));
  jand g0613(.dina(n174), .dinb(n126), .dout(n662));
  jand g0614(.dina(n185), .dinb(n224), .dout(n663));
  jor  g0615(.dina(n663), .dinb(n662), .dout(n664));
  jor  g0616(.dina(n664), .dinb(n661), .dout(n665));
  jand g0617(.dina(n311), .dinb(n143), .dout(n666));
  jand g0618(.dina(n666), .dinb(n100), .dout(n667));
  jor  g0619(.dina(n667), .dinb(n553), .dout(n668));
  jand g0620(.dina(n311), .dinb(n184), .dout(n669));
  jor  g0621(.dina(n669), .dinb(n668), .dout(n670));
  jor  g0622(.dina(n670), .dinb(n665), .dout(n671));
  jand g0623(.dina(n154), .dinb(n130), .dout(n672));
  jand g0624(.dina(n174), .dinb(n145), .dout(n673));
  jor  g0625(.dina(n673), .dinb(n672), .dout(n674));
  jand g0626(.dina(n192), .dinb(n184), .dout(n675));
  jand g0627(.dina(n112), .dinb(n224), .dout(n676));
  jand g0628(.dina(n155), .dinb(n262), .dout(n677));
  jor  g0629(.dina(n677), .dinb(n676), .dout(n678));
  jor  g0630(.dina(n678), .dinb(n675), .dout(n679));
  jor  g0631(.dina(n679), .dinb(n674), .dout(n680));
  jor  g0632(.dina(n680), .dinb(n671), .dout(n681));
  jor  g0633(.dina(n681), .dinb(n659), .dout(n682));
  jor  g0634(.dina(n682), .dinb(n644), .dout(n683));
  jand g0635(.dina(n131), .dinb(n100), .dout(n684));
  jand g0636(.dina(n185), .dinb(n154), .dout(n685));
  jand g0637(.dina(n154), .dinb(n112), .dout(n686));
  jor  g0638(.dina(n686), .dinb(n685), .dout(n687));
  jor  g0639(.dina(n687), .dinb(n684), .dout(n688));
  jand g0640(.dina(n155), .dinb(n224), .dout(n689));
  jand g0641(.dina(n263), .dinb(n118), .dout(n690));
  jor  g0642(.dina(n690), .dinb(n689), .dout(n691));
  jor  g0643(.dina(n691), .dinb(n314), .dout(n692));
  jor  g0644(.dina(n692), .dinb(n688), .dout(n693));
  jand g0645(.dina(n185), .dinb(n174), .dout(n694));
  jand g0646(.dina(n167), .dinb(n118), .dout(n695));
  jor  g0647(.dina(n695), .dinb(n694), .dout(n696));
  jand g0648(.dina(n143), .dinb(n126), .dout(n697));
  jor  g0649(.dina(n697), .dinb(n579), .dout(n698));
  jor  g0650(.dina(n698), .dinb(n696), .dout(n699));
  jand g0651(.dina(n174), .dinb(n155), .dout(n700));
  jand g0652(.dina(n118), .dinb(n112), .dout(n701));
  jor  g0653(.dina(n701), .dinb(n700), .dout(n702));
  jor  g0654(.dina(n702), .dinb(n699), .dout(n703));
  jor  g0655(.dina(n703), .dinb(n693), .dout(n704));
  jand g0656(.dina(n171), .dinb(n253), .dout(n705));
  jand g0657(.dina(n624), .dinb(n77), .dout(n706));
  jand g0658(.dina(n167), .dinb(n144), .dout(n707));
  jand g0659(.dina(n192), .dinb(n223), .dout(n708));
  jand g0660(.dina(n708), .dinb(n77), .dout(n709));
  jor  g0661(.dina(n709), .dinb(n707), .dout(n710));
  jor  g0662(.dina(n710), .dinb(n186), .dout(n711));
  jor  g0663(.dina(n711), .dinb(n706), .dout(n712));
  jor  g0664(.dina(n712), .dinb(n705), .dout(n713));
  jor  g0665(.dina(n713), .dinb(n704), .dout(n714));
  jor  g0666(.dina(n714), .dinb(n683), .dout(n715));
  jor  g0667(.dina(n715), .dinb(n638), .dout(n716));
  jor  g0668(.dina(n194), .dinb(n100), .dout(n717));
  jand g0669(.dina(n171), .dinb(n223), .dout(n718));
  jor  g0670(.dina(n718), .dinb(n673), .dout(n719));
  jnot g0671(.din(n719), .dout(n720));
  jand g0672(.dina(n720), .dinb(n717), .dout(n721));
  jand g0673(.dina(n240), .dinb(n197), .dout(n722));
  jand g0674(.dina(n722), .dinb(n721), .dout(n723));
  jnot g0675(.din(n723), .dout(n724));
  jor  g0676(.dina(n399), .dinb(n282), .dout(n725));
  jand g0677(.dina(n263), .dinb(n144), .dout(n726));
  jand g0678(.dina(n98), .dinb(n262), .dout(n727));
  jor  g0679(.dina(n727), .dinb(n726), .dout(n728));
  jand g0680(.dina(n174), .dinb(n92), .dout(n729));
  jor  g0681(.dina(n684), .dinb(n729), .dout(n730));
  jor  g0682(.dina(n730), .dinb(n728), .dout(n731));
  jor  g0683(.dina(n731), .dinb(n725), .dout(n732));
  jor  g0684(.dina(n630), .dinb(n652), .dout(n733));
  jor  g0685(.dina(n733), .dinb(n299), .dout(n734));
  jor  g0686(.dina(n734), .dinb(n677), .dout(n735));
  jor  g0687(.dina(n735), .dinb(n732), .dout(n736));
  jand g0688(.dina(n708), .dinb(n100), .dout(n737));
  jor  g0689(.dina(n737), .dinb(n706), .dout(n738));
  jor  g0690(.dina(n738), .dinb(n426), .dout(n739));
  jor  g0691(.dina(n739), .dinb(n400), .dout(n740));
  jand g0692(.dina(n126), .dinb(n224), .dout(n741));
  jor  g0693(.dina(n676), .dinb(n741), .dout(n742));
  jor  g0694(.dina(n690), .dinb(n742), .dout(n743));
  jor  g0695(.dina(n308), .dinb(n132), .dout(n744));
  jor  g0696(.dina(n744), .dinb(n743), .dout(n745));
  jor  g0697(.dina(n745), .dinb(n740), .dout(n746));
  jor  g0698(.dina(n746), .dinb(n736), .dout(n747));
  jor  g0699(.dina(n747), .dinb(n724), .dout(n748));
  jand g0700(.dina(n154), .dinb(n126), .dout(n749));
  jand g0701(.dina(n130), .dinb(n224), .dout(n750));
  jor  g0702(.dina(n750), .dinb(n749), .dout(n751));
  jand g0703(.dina(n144), .dinb(n116), .dout(n752));
  jand g0704(.dina(n126), .dinb(n118), .dout(n753));
  jor  g0705(.dina(n753), .dinb(n752), .dout(n754));
  jor  g0706(.dina(n754), .dinb(n617), .dout(n755));
  jor  g0707(.dina(n755), .dinb(n751), .dout(n756));
  jor  g0708(.dina(n756), .dinb(n264), .dout(n757));
  jand g0709(.dina(n154), .dinb(n116), .dout(n758));
  jand g0710(.dina(n192), .dinb(n118), .dout(n759));
  jor  g0711(.dina(n759), .dinb(n686), .dout(n760));
  jor  g0712(.dina(n760), .dinb(n758), .dout(n761));
  jand g0713(.dina(n140), .dinb(n144), .dout(n762));
  jand g0714(.dina(n155), .dinb(n184), .dout(n763));
  jor  g0715(.dina(n763), .dinb(n762), .dout(n764));
  jor  g0716(.dina(n764), .dinb(n761), .dout(n765));
  jand g0717(.dina(n230), .dinb(n253), .dout(n766));
  jand g0718(.dina(n174), .dinb(n171), .dout(n767));
  jand g0719(.dina(n144), .dinb(n130), .dout(n768));
  jor  g0720(.dina(n609), .dinb(n768), .dout(n769));
  jor  g0721(.dina(n769), .dinb(n767), .dout(n770));
  jor  g0722(.dina(n770), .dinb(n766), .dout(n771));
  jor  g0723(.dina(n771), .dinb(n765), .dout(n772));
  jor  g0724(.dina(n772), .dinb(n757), .dout(n773));
  jand g0725(.dina(n666), .dinb(n77), .dout(n774));
  jor  g0726(.dina(n689), .dinb(n774), .dout(n775));
  jor  g0727(.dina(n775), .dinb(n610), .dout(n776));
  jand g0728(.dina(n167), .dinb(n154), .dout(n777));
  jand g0729(.dina(n224), .dinb(n92), .dout(n778));
  jor  g0730(.dina(n778), .dinb(n663), .dout(n779));
  jor  g0731(.dina(n779), .dinb(n777), .dout(n780));
  jor  g0732(.dina(n780), .dinb(n702), .dout(n781));
  jor  g0733(.dina(n781), .dinb(n776), .dout(n782));
  jor  g0734(.dina(n782), .dinb(n644), .dout(n783));
  jor  g0735(.dina(n783), .dinb(n773), .dout(n784));
  jor  g0736(.dina(n410), .dinb(n266), .dout(n785));
  jor  g0737(.dina(n785), .dinb(n496), .dout(n786));
  jnot g0738(.din(n170), .dout(n787));
  jand g0739(.dina(n171), .dinb(n184), .dout(n788));
  jor  g0740(.dina(n669), .dinb(n788), .dout(n789));
  jor  g0741(.dina(n789), .dinb(n705), .dout(n790));
  jor  g0742(.dina(n790), .dinb(n787), .dout(n791));
  jor  g0743(.dina(n791), .dinb(n786), .dout(n792));
  jand g0744(.dina(n126), .dinb(n184), .dout(n793));
  jor  g0745(.dina(n645), .dinb(n793), .dout(n794));
  jand g0746(.dina(n130), .dinb(n253), .dout(n795));
  jand g0747(.dina(n253), .dinb(n112), .dout(n796));
  jor  g0748(.dina(n796), .dinb(n795), .dout(n797));
  jand g0749(.dina(n263), .dinb(n253), .dout(n798));
  jor  g0750(.dina(n648), .dinb(n798), .dout(n799));
  jor  g0751(.dina(n799), .dinb(n797), .dout(n800));
  jor  g0752(.dina(n800), .dinb(n794), .dout(n801));
  jand g0753(.dina(n230), .dinb(n154), .dout(n802));
  jor  g0754(.dina(n330), .dinb(n802), .dout(n803));
  jor  g0755(.dina(n803), .dinb(n801), .dout(n804));
  jor  g0756(.dina(n613), .dinb(n470), .dout(n805));
  jand g0757(.dina(n144), .dinb(n126), .dout(n806));
  jor  g0758(.dina(n806), .dinb(n523), .dout(n807));
  jor  g0759(.dina(n807), .dinb(n805), .dout(n808));
  jor  g0760(.dina(n808), .dinb(n146), .dout(n809));
  jor  g0761(.dina(n809), .dinb(n804), .dout(n810));
  jor  g0762(.dina(n810), .dinb(n792), .dout(n811));
  jor  g0763(.dina(n811), .dinb(n784), .dout(n812));
  jor  g0764(.dina(n812), .dinb(n748), .dout(n813));
  jand g0765(.dina(n813), .dinb(n716), .dout(n814));
  jor  g0766(.dina(n814), .dinb(n607), .dout(n815));
  jnot g0767(.din(n725), .dout(n816));
  jand g0768(.dina(n534), .dinb(n347), .dout(n817));
  jand g0769(.dina(n527), .dinb(n395), .dout(n818));
  jand g0770(.dina(n818), .dinb(n817), .dout(n819));
  jand g0771(.dina(n819), .dinb(n816), .dout(n820));
  jand g0772(.dina(n332), .dinb(n269), .dout(n821));
  jand g0773(.dina(n821), .dinb(n300), .dout(n822));
  jand g0774(.dina(n822), .dinb(n378), .dout(n823));
  jand g0775(.dina(n823), .dinb(n820), .dout(n824));
  jor  g0776(.dina(n268), .dinb(n217), .dout(n825));
  jand g0777(.dina(n195), .dinb(n160), .dout(n826));
  jand g0778(.dina(n826), .dinb(n427), .dout(n827));
  jand g0779(.dina(n827), .dinb(n825), .dout(n828));
  jand g0780(.dina(n561), .dinb(n351), .dout(n829));
  jnot g0781(.din(n744), .dout(n830));
  jand g0782(.dina(n830), .dinb(n829), .dout(n831));
  jand g0783(.dina(n831), .dinb(n828), .dout(n832));
  jand g0784(.dina(n832), .dinb(n824), .dout(n833));
  jand g0785(.dina(n833), .dinb(n723), .dout(n834));
  jand g0786(.dina(n389), .dinb(n191), .dout(n835));
  jand g0787(.dina(n835), .dinb(n294), .dout(n836));
  jand g0788(.dina(n836), .dinb(n539), .dout(n837));
  jand g0789(.dina(n837), .dinb(n265), .dout(n838));
  jand g0790(.dina(n276), .dinb(n142), .dout(n839));
  jand g0791(.dina(n839), .dinb(n572), .dout(n840));
  jand g0792(.dina(n221), .dinb(n162), .dout(n841));
  jand g0793(.dina(n841), .dinb(n435), .dout(n842));
  jand g0794(.dina(n842), .dinb(n506), .dout(n843));
  jand g0795(.dina(n843), .dinb(n840), .dout(n844));
  jand g0796(.dina(n844), .dinb(n838), .dout(n845));
  jand g0797(.dina(n403), .dinb(n114), .dout(n846));
  jand g0798(.dina(n846), .dinb(n245), .dout(n847));
  jand g0799(.dina(n847), .dinb(n457), .dout(n848));
  jand g0800(.dina(n848), .dinb(n213), .dout(n849));
  jand g0801(.dina(n321), .dinb(n286), .dout(n850));
  jand g0802(.dina(n850), .dinb(n370), .dout(n851));
  jor  g0803(.dina(n336), .dinb(n113), .dout(n852));
  jand g0804(.dina(n852), .dinb(n218), .dout(n853));
  jand g0805(.dina(n461), .dinb(n236), .dout(n854));
  jand g0806(.dina(n854), .dinb(n853), .dout(n855));
  jand g0807(.dina(n855), .dinb(n851), .dout(n856));
  jand g0808(.dina(n856), .dinb(n849), .dout(n857));
  jand g0809(.dina(n857), .dinb(n845), .dout(n858));
  jnot g0810(.din(n786), .dout(n859));
  jand g0811(.dina(n456), .dinb(n170), .dout(n860));
  jand g0812(.dina(n860), .dinb(n859), .dout(n861));
  jand g0813(.dina(n374), .dinb(n353), .dout(n862));
  jand g0814(.dina(n510), .dinb(n489), .dout(n863));
  jand g0815(.dina(n366), .dinb(n346), .dout(n864));
  jand g0816(.dina(n864), .dinb(n863), .dout(n865));
  jand g0817(.dina(n865), .dinb(n862), .dout(n866));
  jnot g0818(.din(n803), .dout(n867));
  jand g0819(.dina(n867), .dinb(n866), .dout(n868));
  jand g0820(.dina(n377), .dinb(n204), .dout(n869));
  jand g0821(.dina(n188), .dinb(n158), .dout(n870));
  jand g0822(.dina(n870), .dinb(n869), .dout(n871));
  jand g0823(.dina(n871), .dinb(n147), .dout(n872));
  jand g0824(.dina(n872), .dinb(n868), .dout(n873));
  jand g0825(.dina(n873), .dinb(n861), .dout(n874));
  jand g0826(.dina(n874), .dinb(n858), .dout(n875));
  jand g0827(.dina(n875), .dinb(n834), .dout(n876));
  jxor g0828(.dina(n876), .dinb(n716), .dout(n877));
  jand g0829(.dina(n877), .dinb(n815), .dout(n878));
  jand g0830(.dina(n57), .dinb(n49), .dout(n879));
  jxor g0831(.dina(n879), .dinb(a9 ), .dout(n880));
  jnot g0832(.din(n880), .dout(n881));
  jand g0833(.dina(n881), .dinb(n878), .dout(n882));
  jand g0834(.dina(n370), .dinb(n221), .dout(n883));
  jand g0835(.dina(n377), .dinb(n233), .dout(n884));
  jand g0836(.dina(n884), .dinb(n883), .dout(n885));
  jand g0837(.dina(n885), .dinb(n361), .dout(n886));
  jand g0838(.dina(n267), .dinb(n129), .dout(n887));
  jand g0839(.dina(n887), .dinb(n294), .dout(n888));
  jand g0840(.dina(n888), .dinb(n886), .dout(n889));
  jand g0841(.dina(n387), .dinb(n222), .dout(n890));
  jand g0842(.dina(n890), .dinb(n600), .dout(n891));
  jand g0843(.dina(n891), .dinb(n448), .dout(n892));
  jand g0844(.dina(n587), .dinb(n335), .dout(n893));
  jand g0845(.dina(n893), .dinb(n892), .dout(n894));
  jand g0846(.dina(n894), .dinb(n889), .dout(n895));
  jand g0847(.dina(n895), .dinb(n417), .dout(n896));
  jor  g0848(.dina(n151), .dinb(n108), .dout(n897));
  jand g0849(.dina(n897), .dinb(n366), .dout(n898));
  jand g0850(.dina(n898), .dinb(n463), .dout(n899));
  jand g0851(.dina(n481), .dinb(n290), .dout(n900));
  jand g0852(.dina(n900), .dinb(n825), .dout(n901));
  jand g0853(.dina(n901), .dinb(n557), .dout(n902));
  jand g0854(.dina(n902), .dinb(n899), .dout(n903));
  jand g0855(.dina(n418), .dinb(n261), .dout(n904));
  jand g0856(.dina(n904), .dinb(n546), .dout(n905));
  jand g0857(.dina(n344), .dinb(n281), .dout(n906));
  jand g0858(.dina(n906), .dinb(n905), .dout(n907));
  jand g0859(.dina(n445), .dinb(n152), .dout(n908));
  jand g0860(.dina(n378), .dinb(n305), .dout(n909));
  jand g0861(.dina(n909), .dinb(n339), .dout(n910));
  jand g0862(.dina(n910), .dinb(n908), .dout(n911));
  jand g0863(.dina(n911), .dinb(n907), .dout(n912));
  jand g0864(.dina(n912), .dinb(n903), .dout(n913));
  jand g0865(.dina(n913), .dinb(n849), .dout(n914));
  jand g0866(.dina(n569), .dinb(n535), .dout(n915));
  jand g0867(.dina(n915), .dinb(n527), .dout(n916));
  jand g0868(.dina(n562), .dinb(n315), .dout(n917));
  jand g0869(.dina(n917), .dinb(n916), .dout(n918));
  jnot g0870(.din(n697), .dout(n919));
  jand g0871(.dina(n919), .dinb(n439), .dout(n920));
  jand g0872(.dina(n920), .dinb(n338), .dout(n921));
  jand g0873(.dina(n853), .dinb(n921), .dout(n922));
  jand g0874(.dina(n922), .dinb(n918), .dout(n923));
  jand g0875(.dina(n717), .dinb(n169), .dout(n924));
  jand g0876(.dina(n924), .dinb(n187), .dout(n925));
  jand g0877(.dina(n925), .dinb(n160), .dout(n926));
  jand g0878(.dina(n926), .dinb(n310), .dout(n927));
  jand g0879(.dina(n927), .dinb(n923), .dout(n928));
  jand g0880(.dina(n928), .dinb(n914), .dout(n929));
  jand g0881(.dina(n929), .dinb(n896), .dout(n930));
  jand g0882(.dina(n876), .dinb(n930), .dout(n931));
  jnot g0883(.din(n522), .dout(n932));
  jnot g0884(.din(n528), .dout(n933));
  jor  g0885(.dina(n933), .dinb(n524), .dout(n934));
  jor  g0886(.dina(n934), .dinb(n932), .dout(n935));
  jnot g0887(.din(n532), .dout(n936));
  jor  g0888(.dina(n936), .dinb(n935), .dout(n937));
  jand g0889(.dina(n167), .dinb(n224), .dout(n938));
  jor  g0890(.dina(n752), .dinb(n938), .dout(n939));
  jor  g0891(.dina(n939), .dinb(n685), .dout(n940));
  jor  g0892(.dina(n940), .dinb(n727), .dout(n941));
  jand g0893(.dina(n192), .dinb(n253), .dout(n942));
  jor  g0894(.dina(n766), .dinb(n942), .dout(n943));
  jor  g0895(.dina(n943), .dinb(n751), .dout(n944));
  jor  g0896(.dina(n944), .dinb(n266), .dout(n945));
  jor  g0897(.dina(n945), .dinb(n941), .dout(n946));
  jand g0898(.dina(n295), .dinb(n100), .dout(n947));
  jor  g0899(.dina(n947), .dinb(n612), .dout(n948));
  jor  g0900(.dina(n948), .dinb(n282), .dout(n949));
  jor  g0901(.dina(n949), .dinb(n401), .dout(n950));
  jor  g0902(.dina(n661), .dinb(n132), .dout(n951));
  jor  g0903(.dina(n951), .dinb(n544), .dout(n952));
  jor  g0904(.dina(n952), .dinb(n950), .dout(n953));
  jor  g0905(.dina(n953), .dinb(n946), .dout(n954));
  jor  g0906(.dina(n954), .dinb(n937), .dout(n955));
  jnot g0907(.din(n552), .dout(n956));
  jnot g0908(.din(n559), .dout(n957));
  jor  g0909(.dina(n957), .dinb(n555), .dout(n958));
  jnot g0910(.din(n563), .dout(n959));
  jor  g0911(.dina(n959), .dinb(n958), .dout(n960));
  jor  g0912(.dina(n960), .dinb(n956), .dout(n961));
  jor  g0913(.dina(n961), .dinb(n955), .dout(n962));
  jnot g0914(.din(n574), .dout(n963));
  jor  g0915(.dina(n655), .dinb(n646), .dout(n964));
  jand g0916(.dina(n155), .dinb(n118), .dout(n965));
  jand g0917(.dina(n253), .dinb(n98), .dout(n966));
  jor  g0918(.dina(n966), .dinb(n965), .dout(n967));
  jor  g0919(.dina(n967), .dinb(n964), .dout(n968));
  jand g0920(.dina(n155), .dinb(n144), .dout(n969));
  jor  g0921(.dina(n634), .dinb(n969), .dout(n970));
  jor  g0922(.dina(n802), .dinb(n619), .dout(n971));
  jor  g0923(.dina(n971), .dinb(n970), .dout(n972));
  jor  g0924(.dina(n972), .dinb(n968), .dout(n973));
  jand g0925(.dina(n230), .dinb(n184), .dout(n974));
  jand g0926(.dina(n174), .dinb(n98), .dout(n975));
  jor  g0927(.dina(n975), .dinb(n974), .dout(n976));
  jor  g0928(.dina(n976), .dinb(n247), .dout(n977));
  jand g0929(.dina(n155), .dinb(n253), .dout(n978));
  jor  g0930(.dina(n978), .dinb(n654), .dout(n979));
  jor  g0931(.dina(n979), .dinb(n677), .dout(n980));
  jor  g0932(.dina(n980), .dinb(n977), .dout(n981));
  jor  g0933(.dina(n981), .dinb(n973), .dout(n982));
  jor  g0934(.dina(n982), .dinb(n582), .dout(n983));
  jnot g0935(.din(n604), .dout(n984));
  jor  g0936(.dina(n984), .dinb(n983), .dout(n985));
  jor  g0937(.dina(n985), .dinb(n963), .dout(n986));
  jor  g0938(.dina(n986), .dinb(n962), .dout(n987));
  jand g0939(.dina(n814), .dinb(n987), .dout(n988));
  jor  g0940(.dina(n988), .dinb(n931), .dout(n989));
  jand g0941(.dina(n989), .dinb(n880), .dout(n990));
  jor  g0942(.dina(n990), .dinb(n882), .dout(n991));
  jor  g0943(.dina(n931), .dinb(n815), .dout(n992));
  jand g0944(.dina(n58), .dinb(n49), .dout(n993));
  jxor g0945(.dina(n993), .dinb(a10 ), .dout(n994));
  jand g0946(.dina(n994), .dinb(n992), .dout(n995));
  jnot g0947(.din(n994), .dout(n996));
  jor  g0948(.dina(n877), .dinb(n987), .dout(n997));
  jand g0949(.dina(n997), .dinb(n996), .dout(n998));
  jor  g0950(.dina(n998), .dinb(n995), .dout(n999));
  jnot g0951(.din(n999), .dout(n1000));
  jor  g0952(.dina(n1000), .dinb(n991), .dout(n1001));
  jand g0953(.dina(n250), .dinb(n120), .dout(n1002));
  jand g0954(.dina(n488), .dinb(n409), .dout(n1003));
  jand g0955(.dina(n192), .dinb(n144), .dout(n1004));
  jnot g0956(.din(n1004), .dout(n1005));
  jand g0957(.dina(n1005), .dinb(n570), .dout(n1006));
  jand g0958(.dina(n333), .dinb(n245), .dout(n1007));
  jand g0959(.dina(n1007), .dinb(n1006), .dout(n1008));
  jand g0960(.dina(n1008), .dinb(n1003), .dout(n1009));
  jand g0961(.dina(n1009), .dinb(n352), .dout(n1010));
  jand g0962(.dina(n1010), .dinb(n1002), .dout(n1011));
  jand g0963(.dina(n344), .dinb(n187), .dout(n1012));
  jand g0964(.dina(n1012), .dinb(n897), .dout(n1013));
  jand g0965(.dina(n1013), .dinb(n398), .dout(n1014));
  jand g0966(.dina(n1014), .dinb(n166), .dout(n1015));
  jand g0967(.dina(n1015), .dinb(n1011), .dout(n1016));
  jnot g0968(.din(n785), .dout(n1017));
  jand g0969(.dina(n332), .dinb(n128), .dout(n1018));
  jand g0970(.dina(n404), .dinb(n252), .dout(n1019));
  jand g0971(.dina(n1019), .dinb(n841), .dout(n1020));
  jand g0972(.dina(n1020), .dinb(n1018), .dout(n1021));
  jand g0973(.dina(n1021), .dinb(n1017), .dout(n1022));
  jand g0974(.dina(n278), .dinb(n261), .dout(n1023));
  jand g0975(.dina(n1023), .dinb(n240), .dout(n1024));
  jand g0976(.dina(n195), .dinb(n158), .dout(n1025));
  jor  g0977(.dina(n965), .dinb(n314), .dout(n1026));
  jnot g0978(.din(n1026), .dout(n1027));
  jand g0979(.dina(n1027), .dinb(n1025), .dout(n1028));
  jand g0980(.dina(n1028), .dinb(n1024), .dout(n1029));
  jand g0981(.dina(n527), .dinb(n340), .dout(n1030));
  jand g0982(.dina(n1030), .dinb(n1029), .dout(n1031));
  jand g0983(.dina(n1031), .dinb(n1022), .dout(n1032));
  jand g0984(.dina(n275), .dinb(n152), .dout(n1033));
  jand g0985(.dina(n301), .dinb(n77), .dout(n1034));
  jnot g0986(.din(n1034), .dout(n1035));
  jand g0987(.dina(n1035), .dinb(n384), .dout(n1036));
  jand g0988(.dina(n506), .dinb(n438), .dout(n1037));
  jand g0989(.dina(n1037), .dinb(n1036), .dout(n1038));
  jand g0990(.dina(n1038), .dinb(n1033), .dout(n1039));
  jor  g0991(.dina(n796), .dinb(n426), .dout(n1040));
  jnot g0992(.din(n1040), .dout(n1041));
  jand g0993(.dina(n1041), .dinb(n234), .dout(n1042));
  jand g0994(.dina(n347), .dinb(n310), .dout(n1043));
  jand g0995(.dina(n1043), .dinb(n402), .dout(n1044));
  jand g0996(.dina(n1044), .dinb(n1042), .dout(n1045));
  jand g0997(.dina(n1045), .dinb(n159), .dout(n1046));
  jand g0998(.dina(n1046), .dinb(n1039), .dout(n1047));
  jand g0999(.dina(n1047), .dinb(n1032), .dout(n1048));
  jand g1000(.dina(n569), .dinb(n382), .dout(n1049));
  jand g1001(.dina(n1049), .dinb(n269), .dout(n1050));
  jand g1002(.dina(n1050), .dinb(n377), .dout(n1051));
  jand g1003(.dina(n420), .dinb(n248), .dout(n1052));
  jand g1004(.dina(n1052), .dinb(n1051), .dout(n1053));
  jand g1005(.dina(n1053), .dinb(n1048), .dout(n1054));
  jand g1006(.dina(n1054), .dinb(n1016), .dout(n1055));
  jand g1007(.dina(n915), .dinb(n133), .dout(n1056));
  jand g1008(.dina(n429), .dinb(n332), .dout(n1057));
  jand g1009(.dina(n1057), .dinb(n215), .dout(n1058));
  jand g1010(.dina(n1058), .dinb(n437), .dout(n1059));
  jand g1011(.dina(n1059), .dinb(n1056), .dout(n1060));
  jand g1012(.dina(n835), .dinb(n489), .dout(n1061));
  jand g1013(.dina(n497), .dinb(n238), .dout(n1062));
  jand g1014(.dina(n1062), .dinb(n1061), .dout(n1063));
  jand g1015(.dina(n300), .dinb(n136), .dout(n1064));
  jand g1016(.dina(n1064), .dinb(n148), .dout(n1065));
  jand g1017(.dina(n377), .dinb(n315), .dout(n1066));
  jand g1018(.dina(n1066), .dinb(n1065), .dout(n1067));
  jand g1019(.dina(n1067), .dinb(n1063), .dout(n1068));
  jand g1020(.dina(n1068), .dinb(n1060), .dout(n1069));
  jand g1021(.dina(n1069), .dinb(n570), .dout(n1070));
  jand g1022(.dina(n1070), .dinb(n370), .dout(n1071));
  jand g1023(.dina(n378), .dinb(n226), .dout(n1072));
  jnot g1024(.din(n577), .dout(n1073));
  jand g1025(.dina(n1073), .dinb(n460), .dout(n1074));
  jand g1026(.dina(n1074), .dinb(n197), .dout(n1075));
  jand g1027(.dina(n427), .dinb(n129), .dout(n1076));
  jand g1028(.dina(n1076), .dinb(n1075), .dout(n1077));
  jand g1029(.dina(n1077), .dinb(n904), .dout(n1078));
  jand g1030(.dina(n1078), .dinb(n1012), .dout(n1079));
  jand g1031(.dina(n445), .dinb(n395), .dout(n1080));
  jand g1032(.dina(n1080), .dinb(n850), .dout(n1081));
  jand g1033(.dina(n1081), .dinb(n1079), .dout(n1082));
  jand g1034(.dina(n1082), .dinb(n1072), .dout(n1083));
  jand g1035(.dina(n1083), .dinb(n1071), .dout(n1084));
  jand g1036(.dina(n310), .dinb(n222), .dout(n1085));
  jand g1037(.dina(n1085), .dinb(n435), .dout(n1086));
  jand g1038(.dina(n1086), .dinb(n248), .dout(n1087));
  jand g1039(.dina(n294), .dinb(n114), .dout(n1088));
  jand g1040(.dina(n1088), .dinb(n366), .dout(n1089));
  jand g1041(.dina(n1089), .dinb(n1087), .dout(n1090));
  jand g1042(.dina(n467), .dinb(n218), .dout(n1091));
  jand g1043(.dina(n313), .dinb(n276), .dout(n1092));
  jand g1044(.dina(n1092), .dinb(n1091), .dout(n1093));
  jand g1045(.dina(n185), .dinb(n144), .dout(n1094));
  jnot g1046(.din(n1094), .dout(n1095));
  jand g1047(.dina(n462), .dinb(n206), .dout(n1096));
  jand g1048(.dina(n1096), .dinb(n1095), .dout(n1097));
  jand g1049(.dina(n232), .dinb(n160), .dout(n1098));
  jand g1050(.dina(n1098), .dinb(n1097), .dout(n1099));
  jand g1051(.dina(n1099), .dinb(n1093), .dout(n1100));
  jand g1052(.dina(n290), .dinb(n204), .dout(n1101));
  jand g1053(.dina(n1101), .dinb(n446), .dout(n1102));
  jand g1054(.dina(n280), .dinb(n157), .dout(n1103));
  jand g1055(.dina(n1103), .dinb(n267), .dout(n1104));
  jand g1056(.dina(n506), .dinb(n404), .dout(n1105));
  jand g1057(.dina(n1105), .dinb(n362), .dout(n1106));
  jand g1058(.dina(n1106), .dinb(n1104), .dout(n1107));
  jand g1059(.dina(n1107), .dinb(n1102), .dout(n1108));
  jand g1060(.dina(n1108), .dinb(n1100), .dout(n1109));
  jand g1061(.dina(n717), .dinb(n173), .dout(n1110));
  jand g1062(.dina(n1110), .dinb(n288), .dout(n1111));
  jand g1063(.dina(n1111), .dinb(n1109), .dout(n1112));
  jand g1064(.dina(n1112), .dinb(n1090), .dout(n1113));
  jand g1065(.dina(n1113), .dinb(n1084), .dout(n1114));
  jxor g1066(.dina(n1114), .dinb(n1055), .dout(n1115));
  jor  g1067(.dina(n1114), .dinb(n1055), .dout(n1116));
  jand g1068(.dina(n1005), .dinb(n374), .dout(n1117));
  jand g1069(.dina(n446), .dinb(n267), .dout(n1118));
  jand g1070(.dina(n1118), .dinb(n1117), .dout(n1119));
  jand g1071(.dina(n1119), .dinb(n603), .dout(n1120));
  jand g1072(.dina(n467), .dinb(n339), .dout(n1121));
  jand g1073(.dina(n1121), .dinb(n346), .dout(n1122));
  jand g1074(.dina(n1088), .dinb(n492), .dout(n1123));
  jand g1075(.dina(n1123), .dinb(n448), .dout(n1124));
  jand g1076(.dina(n1124), .dinb(n1122), .dout(n1125));
  jand g1077(.dina(n1125), .dinb(n1120), .dout(n1126));
  jand g1078(.dina(n1073), .dinb(n313), .dout(n1127));
  jand g1079(.dina(n415), .dinb(n327), .dout(n1128));
  jand g1080(.dina(n429), .dinb(n252), .dout(n1129));
  jand g1081(.dina(n1129), .dinb(n1128), .dout(n1130));
  jand g1082(.dina(n1130), .dinb(n527), .dout(n1131));
  jand g1083(.dina(n570), .dinb(n297), .dout(n1132));
  jand g1084(.dina(n1132), .dinb(n222), .dout(n1133));
  jand g1085(.dina(n1133), .dinb(n255), .dout(n1134));
  jand g1086(.dina(n1134), .dinb(n238), .dout(n1135));
  jand g1087(.dina(n1135), .dinb(n1131), .dout(n1136));
  jand g1088(.dina(n1136), .dinb(n1127), .dout(n1137));
  jand g1089(.dina(n1137), .dinb(n1126), .dout(n1138));
  jand g1090(.dina(n510), .dinb(n221), .dout(n1139));
  jand g1091(.dina(n1139), .dinb(n180), .dout(n1140));
  jand g1092(.dina(n720), .dinb(n332), .dout(n1141));
  jand g1093(.dina(n1141), .dinb(n593), .dout(n1142));
  jand g1094(.dina(n1142), .dinb(n372), .dout(n1143));
  jand g1095(.dina(n1143), .dinb(n600), .dout(n1144));
  jand g1096(.dina(n921), .dinb(n191), .dout(n1145));
  jand g1097(.dina(n1145), .dinb(n293), .dout(n1146));
  jand g1098(.dina(n1146), .dinb(n1144), .dout(n1147));
  jand g1099(.dina(n1147), .dinb(n1140), .dout(n1148));
  jand g1100(.dina(n1148), .dinb(n1138), .dout(n1149));
  jnot g1101(.din(n1149), .dout(n1150));
  jand g1102(.dina(n1150), .dinb(n1116), .dout(n1151));
  jor  g1103(.dina(n1151), .dinb(n1115), .dout(n1152));
  jand g1104(.dina(n53), .dinb(n49), .dout(n1153));
  jxor g1105(.dina(n1153), .dinb(a5 ), .dout(n1154));
  jor  g1106(.dina(n1154), .dinb(n1152), .dout(n1155));
  jnot g1107(.din(n1154), .dout(n1156));
  jand g1108(.dina(n1114), .dinb(n1055), .dout(n1157));
  jnot g1109(.din(n1157), .dout(n1158));
  jand g1110(.dina(n1149), .dinb(n1158), .dout(n1159));
  jor  g1111(.dina(n1159), .dinb(n1115), .dout(n1160));
  jor  g1112(.dina(n1160), .dinb(n1156), .dout(n1161));
  jand g1113(.dina(n1161), .dinb(n1155), .dout(n1162));
  jand g1114(.dina(n1151), .dinb(n1158), .dout(n1163));
  jnot g1115(.din(n1163), .dout(n1164));
  jand g1116(.dina(n54), .dinb(n49), .dout(n1165));
  jxor g1117(.dina(n1165), .dinb(a6 ), .dout(n1166));
  jand g1118(.dina(n1166), .dinb(n1164), .dout(n1167));
  jnot g1119(.din(n1166), .dout(n1168));
  jnot g1120(.din(n1115), .dout(n1169));
  jor  g1121(.dina(n1150), .dinb(n1169), .dout(n1170));
  jand g1122(.dina(n1170), .dinb(n1168), .dout(n1171));
  jor  g1123(.dina(n1171), .dinb(n1167), .dout(n1172));
  jand g1124(.dina(n1172), .dinb(n1162), .dout(n1173));
  jnot g1125(.din(n1173), .dout(n1174));
  jor  g1126(.dina(n1174), .dinb(n1001), .dout(n1175));
  jand g1127(.dina(n827), .dinb(n506), .dout(n1176));
  jnot g1128(.din(n1176), .dout(n1177));
  jand g1129(.dina(n387), .dinb(n173), .dout(n1178));
  jnot g1130(.din(n1178), .dout(n1179));
  jor  g1131(.dina(n447), .dinb(n975), .dout(n1180));
  jor  g1132(.dina(n1180), .dinb(n634), .dout(n1181));
  jor  g1133(.dina(n1181), .dinb(n1179), .dout(n1182));
  jor  g1134(.dina(n1182), .dinb(n1177), .dout(n1183));
  jor  g1135(.dina(n1183), .dinb(n787), .dout(n1184));
  jor  g1136(.dina(n660), .dinb(n302), .dout(n1185));
  jor  g1137(.dina(n1185), .dinb(n282), .dout(n1186));
  jor  g1138(.dina(n1186), .dinb(n676), .dout(n1187));
  jor  g1139(.dina(n1187), .dinb(n274), .dout(n1188));
  jor  g1140(.dina(n1188), .dinb(n677), .dout(n1189));
  jor  g1141(.dina(n1189), .dinb(n1184), .dout(n1190));
  jand g1142(.dina(n374), .dinb(n276), .dout(n1191));
  jand g1143(.dina(n1191), .dinb(n1035), .dout(n1192));
  jand g1144(.dina(n1192), .dinb(n136), .dout(n1193));
  jand g1145(.dina(n863), .dinb(n244), .dout(n1194));
  jand g1146(.dina(n1194), .dinb(n1019), .dout(n1195));
  jand g1147(.dina(n1195), .dinb(n1193), .dout(n1196));
  jnot g1148(.din(n1196), .dout(n1197));
  jnot g1149(.din(n1056), .dout(n1198));
  jnot g1150(.din(n437), .dout(n1199));
  jand g1151(.dina(n126), .dinb(n262), .dout(n1200));
  jor  g1152(.dina(n1200), .dinb(n630), .dout(n1201));
  jor  g1153(.dina(n1201), .dinb(n214), .dout(n1202));
  jor  g1154(.dina(n1202), .dinb(n1199), .dout(n1203));
  jor  g1155(.dina(n1203), .dinb(n1198), .dout(n1204));
  jand g1156(.dina(n439), .dinb(n409), .dout(n1205));
  jnot g1157(.din(n1205), .dout(n1206));
  jor  g1158(.dina(n1206), .dinb(n1204), .dout(n1207));
  jor  g1159(.dina(n1207), .dinb(n1197), .dout(n1208));
  jor  g1160(.dina(n617), .dinb(n752), .dout(n1209));
  jor  g1161(.dina(n788), .dinb(n667), .dout(n1210));
  jor  g1162(.dina(n1210), .dinb(n1209), .dout(n1211));
  jor  g1163(.dina(n705), .dinb(n625), .dout(n1212));
  jor  g1164(.dina(n1212), .dinb(n654), .dout(n1213));
  jor  g1165(.dina(n1213), .dinb(n1211), .dout(n1214));
  jor  g1166(.dina(n287), .dinb(n777), .dout(n1215));
  jor  g1167(.dina(n1215), .dinb(n968), .dout(n1216));
  jor  g1168(.dina(n1216), .dinb(n1214), .dout(n1217));
  jand g1169(.dina(n92), .dinb(n262), .dout(n1218));
  jand g1170(.dina(n224), .dinb(n98), .dout(n1219));
  jor  g1171(.dina(n1219), .dinb(n1218), .dout(n1220));
  jor  g1172(.dina(n1094), .dinb(n1220), .dout(n1221));
  jor  g1173(.dina(n1221), .dinb(n700), .dout(n1222));
  jor  g1174(.dina(n1222), .dinb(n616), .dout(n1223));
  jor  g1175(.dina(n1223), .dinb(n1217), .dout(n1224));
  jand g1176(.dina(n1006), .dinb(n527), .dout(n1225));
  jand g1177(.dina(n1225), .dinb(n286), .dout(n1226));
  jnot g1178(.din(n1226), .dout(n1227));
  jor  g1179(.dina(n1227), .dinb(n1224), .dout(n1228));
  jor  g1180(.dina(n1228), .dinb(n1208), .dout(n1229));
  jor  g1181(.dina(n1229), .dinb(n1190), .dout(n1230));
  jand g1182(.dina(n1230), .dinb(n987), .dout(n1231));
  jor  g1183(.dina(n1231), .dinb(n1055), .dout(n1232));
  jnot g1184(.din(n1181), .dout(n1233));
  jand g1185(.dina(n1233), .dinb(n1178), .dout(n1234));
  jand g1186(.dina(n1234), .dinb(n1176), .dout(n1235));
  jand g1187(.dina(n1235), .dinb(n170), .dout(n1236));
  jnot g1188(.din(n1189), .dout(n1237));
  jand g1189(.dina(n1237), .dinb(n1236), .dout(n1238));
  jand g1190(.dina(n1205), .dinb(n1060), .dout(n1239));
  jand g1191(.dina(n1239), .dinb(n1196), .dout(n1240));
  jand g1192(.dina(n1085), .dinb(n290), .dout(n1241));
  jand g1193(.dina(n1241), .dinb(n329), .dout(n1242));
  jnot g1194(.din(n1215), .dout(n1243));
  jand g1195(.dina(n1243), .dinb(n586), .dout(n1244));
  jand g1196(.dina(n1244), .dinb(n1242), .dout(n1245));
  jand g1197(.dina(n1095), .dinb(n103), .dout(n1246));
  jand g1198(.dina(n1246), .dinb(n218), .dout(n1247));
  jand g1199(.dina(n1247), .dinb(n886), .dout(n1248));
  jand g1200(.dina(n1248), .dinb(n1245), .dout(n1249));
  jand g1201(.dina(n1226), .dinb(n1249), .dout(n1250));
  jand g1202(.dina(n1250), .dinb(n1240), .dout(n1251));
  jand g1203(.dina(n1251), .dinb(n1238), .dout(n1252));
  jand g1204(.dina(n1252), .dinb(n607), .dout(n1253));
  jor  g1205(.dina(n1253), .dinb(n1232), .dout(n1254));
  jnot g1206(.din(n1254), .dout(n1255));
  jand g1207(.dina(n56), .dinb(n49), .dout(n1256));
  jxor g1208(.dina(n1256), .dinb(a8 ), .dout(n1257));
  jand g1209(.dina(n1257), .dinb(n1255), .dout(n1258));
  jnot g1210(.din(n1257), .dout(n1259));
  jxor g1211(.dina(n1252), .dinb(n607), .dout(n1260));
  jand g1212(.dina(n1260), .dinb(n1055), .dout(n1261));
  jand g1213(.dina(n1261), .dinb(n1259), .dout(n1262));
  jor  g1214(.dina(n1262), .dinb(n1258), .dout(n1263));
  jnot g1215(.din(n1263), .dout(n1264));
  jand g1216(.dina(n55), .dinb(n49), .dout(n1265));
  jxor g1217(.dina(n1265), .dinb(a7 ), .dout(n1266));
  jnot g1218(.din(n1253), .dout(n1267));
  jor  g1219(.dina(n1252), .dinb(n607), .dout(n1268));
  jor  g1220(.dina(n1268), .dinb(n1055), .dout(n1269));
  jand g1221(.dina(n1269), .dinb(n1267), .dout(n1270));
  jand g1222(.dina(n1270), .dinb(n1266), .dout(n1271));
  jnot g1223(.din(n1266), .dout(n1272));
  jnot g1224(.din(n1016), .dout(n1273));
  jnot g1225(.din(n1022), .dout(n1274));
  jnot g1226(.din(n1024), .dout(n1275));
  jnot g1227(.din(n1025), .dout(n1276));
  jor  g1228(.dina(n1026), .dinb(n1276), .dout(n1277));
  jor  g1229(.dina(n1277), .dinb(n1275), .dout(n1278));
  jnot g1230(.din(n1030), .dout(n1279));
  jor  g1231(.dina(n1279), .dinb(n1278), .dout(n1280));
  jor  g1232(.dina(n1280), .dinb(n1274), .dout(n1281));
  jnot g1233(.din(n1039), .dout(n1282));
  jnot g1234(.din(n234), .dout(n1283));
  jor  g1235(.dina(n1040), .dinb(n1283), .dout(n1284));
  jnot g1236(.din(n1043), .dout(n1285));
  jor  g1237(.dina(n1285), .dinb(n401), .dout(n1286));
  jor  g1238(.dina(n1286), .dinb(n1284), .dout(n1287));
  jor  g1239(.dina(n1287), .dinb(n624), .dout(n1288));
  jor  g1240(.dina(n1288), .dinb(n1282), .dout(n1289));
  jor  g1241(.dina(n1289), .dinb(n1281), .dout(n1290));
  jnot g1242(.din(n1053), .dout(n1291));
  jor  g1243(.dina(n1291), .dinb(n1290), .dout(n1292));
  jor  g1244(.dina(n1292), .dinb(n1273), .dout(n1293));
  jand g1245(.dina(n1268), .dinb(n1293), .dout(n1294));
  jor  g1246(.dina(n1260), .dinb(n1294), .dout(n1295));
  jand g1247(.dina(n1295), .dinb(n1272), .dout(n1296));
  jor  g1248(.dina(n1296), .dinb(n1271), .dout(n1297));
  jand g1249(.dina(n1297), .dinb(n1264), .dout(n1298));
  jnot g1250(.din(n1298), .dout(n1299));
  jxor g1251(.dina(n1173), .dinb(n1001), .dout(n1300));
  jor  g1252(.dina(n1300), .dinb(n1299), .dout(n1301));
  jand g1253(.dina(n1301), .dinb(n1175), .dout(n1302));
  jor  g1254(.dina(n1302), .dinb(n521), .dout(n1303));
  jnot g1255(.din(n601), .dout(n1304));
  jor  g1256(.dina(n684), .dinb(n966), .dout(n1305));
  jor  g1257(.dina(n689), .dinb(n266), .dout(n1306));
  jor  g1258(.dina(n1306), .dinb(n1305), .dout(n1307));
  jnot g1259(.din(n1074), .dout(n1308));
  jor  g1260(.dina(n282), .dinb(n749), .dout(n1309));
  jor  g1261(.dina(n1309), .dinb(n1308), .dout(n1310));
  jor  g1262(.dina(n1310), .dinb(n1307), .dout(n1311));
  jor  g1263(.dina(n1311), .dinb(n1304), .dout(n1312));
  jand g1264(.dina(n353), .dinb(n197), .dout(n1313));
  jand g1265(.dina(n280), .dinb(n114), .dout(n1314));
  jand g1266(.dina(n1314), .dinb(n1313), .dout(n1315));
  jnot g1267(.din(n1315), .dout(n1316));
  jor  g1268(.dina(n1316), .dinb(n1312), .dout(n1317));
  jnot g1269(.din(n1105), .dout(n1318));
  jor  g1270(.dina(n1318), .dinb(n777), .dout(n1319));
  jor  g1271(.dina(n1319), .dinb(n974), .dout(n1320));
  jnot g1272(.din(n1320), .dout(n1321));
  jand g1273(.dina(n411), .dinb(n265), .dout(n1322));
  jand g1274(.dina(n1005), .dinb(n439), .dout(n1323));
  jand g1275(.dina(n1323), .dinb(n1322), .dout(n1324));
  jand g1276(.dina(n1064), .dinb(n826), .dout(n1325));
  jand g1277(.dina(n1325), .dinb(n1324), .dout(n1326));
  jor  g1278(.dina(n360), .dinb(n652), .dout(n1327));
  jnot g1279(.din(n1327), .dout(n1328));
  jand g1280(.dina(n1328), .dinb(n1130), .dout(n1329));
  jand g1281(.dina(n1329), .dinb(n1326), .dout(n1330));
  jand g1282(.dina(n1330), .dinb(n1321), .dout(n1331));
  jand g1283(.dina(n409), .dinb(n346), .dout(n1332));
  jand g1284(.dina(n374), .dinb(n288), .dout(n1333));
  jand g1285(.dina(n1333), .dinb(n1332), .dout(n1334));
  jand g1286(.dina(n1334), .dinb(n387), .dout(n1335));
  jand g1287(.dina(n434), .dinb(n255), .dout(n1336));
  jand g1288(.dina(n1336), .dinb(n133), .dout(n1337));
  jand g1289(.dina(n1337), .dinb(n561), .dout(n1338));
  jand g1290(.dina(n1338), .dinb(n1335), .dout(n1339));
  jand g1291(.dina(n232), .dinb(n206), .dout(n1340));
  jand g1292(.dina(n1340), .dinb(n226), .dout(n1341));
  jand g1293(.dina(n316), .dinb(n148), .dout(n1342));
  jand g1294(.dina(n1342), .dinb(n1341), .dout(n1343));
  jor  g1295(.dina(n239), .dinb(n119), .dout(n1344));
  jnot g1296(.din(n1344), .dout(n1345));
  jand g1297(.dina(n852), .dinb(n261), .dout(n1346));
  jand g1298(.dina(n1346), .dinb(n188), .dout(n1347));
  jand g1299(.dina(n1347), .dinb(n1345), .dout(n1348));
  jand g1300(.dina(n1348), .dinb(n1343), .dout(n1349));
  jand g1301(.dina(n1349), .dinb(n1339), .dout(n1350));
  jand g1302(.dina(n1350), .dinb(n1331), .dout(n1351));
  jnot g1303(.din(n1351), .dout(n1352));
  jor  g1304(.dina(n1352), .dinb(n1317), .dout(n1353));
  jnot g1305(.din(n1353), .dout(n1354));
  jand g1306(.dina(n59), .dinb(n49), .dout(n1355));
  jxor g1307(.dina(n1355), .dinb(a11 ), .dout(n1356));
  jand g1308(.dina(n1356), .dinb(n1354), .dout(n1357));
  jnot g1309(.din(n1357), .dout(n1358));
  jand g1310(.dina(n60), .dinb(n49), .dout(n1359));
  jxor g1311(.dina(n1359), .dinb(a12 ), .dout(n1360));
  jand g1312(.dina(n1360), .dinb(n1353), .dout(n1361));
  jxor g1313(.dina(n1361), .dinb(n716), .dout(n1362));
  jand g1314(.dina(n1362), .dinb(n1358), .dout(n1363));
  jand g1315(.dina(n1005), .dinb(n207), .dout(n1364));
  jand g1316(.dina(n1364), .dinb(n233), .dout(n1365));
  jand g1317(.dina(n434), .dinb(n415), .dout(n1366));
  jand g1318(.dina(n387), .dinb(n305), .dout(n1367));
  jand g1319(.dina(n1367), .dinb(n1366), .dout(n1368));
  jand g1320(.dina(n1368), .dinb(n1365), .dout(n1369));
  jand g1321(.dina(n1345), .dinb(n170), .dout(n1370));
  jand g1322(.dina(n1370), .dinb(n1243), .dout(n1371));
  jand g1323(.dina(n339), .dinb(n157), .dout(n1372));
  jand g1324(.dina(n1372), .dinb(n337), .dout(n1373));
  jand g1325(.dina(n1373), .dinb(n488), .dout(n1374));
  jand g1326(.dina(n1374), .dinb(n1371), .dout(n1375));
  jand g1327(.dina(n1375), .dinb(n1346), .dout(n1376));
  jand g1328(.dina(n345), .dinb(n152), .dout(n1377));
  jand g1329(.dina(n1377), .dinb(n276), .dout(n1378));
  jand g1330(.dina(n1378), .dinb(n1376), .dout(n1379));
  jand g1331(.dina(n1379), .dinb(n1369), .dout(n1380));
  jand g1332(.dina(n1380), .dinb(n1071), .dout(n1381));
  jand g1333(.dina(n177), .dinb(n103), .dout(n1382));
  jand g1334(.dina(n438), .dinb(n235), .dout(n1383));
  jand g1335(.dina(n1383), .dinb(n1382), .dout(n1384));
  jand g1336(.dina(n1384), .dinb(n1097), .dout(n1385));
  jand g1337(.dina(n1385), .dinb(n460), .dout(n1386));
  jand g1338(.dina(n1386), .dinb(n232), .dout(n1387));
  jand g1339(.dina(n817), .dinb(n382), .dout(n1388));
  jand g1340(.dina(n594), .dinb(n418), .dout(n1389));
  jand g1341(.dina(n294), .dinb(n286), .dout(n1390));
  jand g1342(.dina(n1390), .dinb(n1389), .dout(n1391));
  jand g1343(.dina(n1391), .dinb(n1388), .dout(n1392));
  jand g1344(.dina(n1392), .dinb(n281), .dout(n1393));
  jand g1345(.dina(n862), .dinb(n527), .dout(n1394));
  jand g1346(.dina(n1394), .dinb(n842), .dout(n1395));
  jand g1347(.dina(n1395), .dinb(n1322), .dout(n1396));
  jand g1348(.dina(n1396), .dinb(n439), .dout(n1397));
  jand g1349(.dina(n1397), .dinb(n1393), .dout(n1398));
  jand g1350(.dina(n1398), .dinb(n1387), .dout(n1399));
  jand g1351(.dina(n1399), .dinb(n1381), .dout(n1400));
  jor  g1352(.dina(n1400), .dinb(n1149), .dout(n1401));
  jand g1353(.dina(n1401), .dinb(n486), .dout(n1402));
  jxor g1354(.dina(n1400), .dinb(n1149), .dout(n1403));
  jand g1355(.dina(n1403), .dinb(n519), .dout(n1404));
  jnot g1356(.din(n1404), .dout(n1405));
  jand g1357(.dina(n1405), .dinb(n1402), .dout(n1406));
  jand g1358(.dina(n1406), .dinb(n1363), .dout(n1407));
  jand g1359(.dina(n1255), .dinb(n880), .dout(n1408));
  jand g1360(.dina(n1261), .dinb(n881), .dout(n1409));
  jor  g1361(.dina(n1409), .dinb(n1408), .dout(n1410));
  jnot g1362(.din(n1410), .dout(n1411));
  jand g1363(.dina(n1270), .dinb(n1257), .dout(n1412));
  jand g1364(.dina(n1295), .dinb(n1259), .dout(n1413));
  jor  g1365(.dina(n1413), .dinb(n1412), .dout(n1414));
  jand g1366(.dina(n1414), .dinb(n1411), .dout(n1415));
  jnot g1367(.din(n1152), .dout(n1416));
  jand g1368(.dina(n1168), .dinb(n1416), .dout(n1417));
  jnot g1369(.din(n1160), .dout(n1418));
  jand g1370(.dina(n1166), .dinb(n1418), .dout(n1419));
  jor  g1371(.dina(n1419), .dinb(n1417), .dout(n1420));
  jnot g1372(.din(n1420), .dout(n1421));
  jand g1373(.dina(n1266), .dinb(n1164), .dout(n1422));
  jand g1374(.dina(n1272), .dinb(n1170), .dout(n1423));
  jor  g1375(.dina(n1423), .dinb(n1422), .dout(n1424));
  jand g1376(.dina(n1424), .dinb(n1421), .dout(n1425));
  jxor g1377(.dina(n1425), .dinb(n1415), .dout(n1426));
  jxor g1378(.dina(n1426), .dinb(n1407), .dout(n1427));
  jnot g1379(.din(n1427), .dout(n1428));
  jxor g1380(.dina(n1302), .dinb(n521), .dout(n1429));
  jnot g1381(.din(n1429), .dout(n1430));
  jor  g1382(.dina(n1430), .dinb(n1428), .dout(n1431));
  jand g1383(.dina(n1431), .dinb(n1303), .dout(n1432));
  jand g1384(.dina(n61), .dinb(n49), .dout(n1433));
  jxor g1385(.dina(n1433), .dinb(a13 ), .dout(n1434));
  jand g1386(.dina(n1434), .dinb(n1354), .dout(n1435));
  jnot g1387(.din(n1435), .dout(n1436));
  jand g1388(.dina(n62), .dinb(n49), .dout(n1437));
  jxor g1389(.dina(n1437), .dinb(a14 ), .dout(n1438));
  jand g1390(.dina(n1438), .dinb(n1353), .dout(n1439));
  jxor g1391(.dina(n1439), .dinb(n716), .dout(n1440));
  jand g1392(.dina(n1440), .dinb(n1436), .dout(n1441));
  jand g1393(.dina(n516), .dinb(n486), .dout(n1442));
  jand g1394(.dina(n1343), .dinb(n361), .dout(n1443));
  jand g1395(.dina(n1443), .dinb(n252), .dout(n1444));
  jand g1396(.dina(n569), .dinb(n321), .dout(n1445));
  jand g1397(.dina(n1445), .dinb(n575), .dout(n1446));
  jand g1398(.dina(n1446), .dinb(n381), .dout(n1447));
  jand g1399(.dina(n347), .dinb(n102), .dout(n1448));
  jand g1400(.dina(n269), .dinb(n191), .dout(n1449));
  jand g1401(.dina(n1449), .dinb(n173), .dout(n1450));
  jand g1402(.dina(n1450), .dinb(n1448), .dout(n1451));
  jand g1403(.dina(n290), .dinb(n233), .dout(n1452));
  jand g1404(.dina(n1452), .dinb(n157), .dout(n1453));
  jand g1405(.dina(n1453), .dinb(n1451), .dout(n1454));
  jand g1406(.dina(n1454), .dinb(n1447), .dout(n1455));
  jand g1407(.dina(n1455), .dinb(n1444), .dout(n1456));
  jand g1408(.dina(n249), .dinb(n99), .dout(n1457));
  jor  g1409(.dina(n1457), .dinb(n134), .dout(n1458));
  jand g1410(.dina(n1005), .dinb(n283), .dout(n1459));
  jand g1411(.dina(n587), .dinb(n182), .dout(n1460));
  jand g1412(.dina(n309), .dinb(n403), .dout(n1461));
  jand g1413(.dina(n1461), .dinb(n1460), .dout(n1462));
  jand g1414(.dina(n1462), .dinb(n1459), .dout(n1463));
  jand g1415(.dina(n384), .dinb(n221), .dout(n1464));
  jand g1416(.dina(n1464), .dinb(n170), .dout(n1465));
  jand g1417(.dina(n1465), .dinb(n919), .dout(n1466));
  jand g1418(.dina(n1466), .dinb(n1463), .dout(n1467));
  jand g1419(.dina(n279), .dinb(n159), .dout(n1468));
  jand g1420(.dina(n1468), .dinb(n534), .dout(n1469));
  jand g1421(.dina(n1469), .dinb(n215), .dout(n1470));
  jand g1422(.dina(n1470), .dinb(n1064), .dout(n1471));
  jand g1423(.dina(n1471), .dinb(n1467), .dout(n1472));
  jand g1424(.dina(n1472), .dinb(n1458), .dout(n1473));
  jand g1425(.dina(n1473), .dinb(n1456), .dout(n1474));
  jxor g1426(.dina(n1494), .dinb(n1441), .dout(n1478));
  jnot g1427(.din(n1478), .dout(n1479));
  jnot g1428(.din(n1356), .dout(n1480));
  jand g1429(.dina(n1480), .dinb(n878), .dout(n1481));
  jand g1430(.dina(n1356), .dinb(n989), .dout(n1482));
  jor  g1431(.dina(n1482), .dinb(n1481), .dout(n1483));
  jand g1432(.dina(n1360), .dinb(n992), .dout(n1484));
  jnot g1433(.din(n1360), .dout(n1485));
  jand g1434(.dina(n1485), .dinb(n997), .dout(n1486));
  jor  g1435(.dina(n1486), .dinb(n1484), .dout(n1487));
  jnot g1436(.din(n1487), .dout(n1488));
  jor  g1437(.dina(n1488), .dinb(n1483), .dout(n1489));
  jnot g1438(.din(n517), .dout(n1490));
  jnot g1439(.din(n486), .dout(n1491));
  jnot g1440(.din(n516), .dout(n1492));
  jand g1441(.dina(n1492), .dinb(n1491), .dout(n1493));
  jnot g1442(.din(n1474), .dout(n1494));
  jand g1443(.dina(n1493), .dinb(n519), .dout(n1497));
  jand g1444(.dina(n52), .dinb(n49), .dout(n1498));
  jxor g1445(.dina(n1498), .dinb(a4 ), .dout(n1499));
  jnot g1446(.din(n1499), .dout(n1500));
  jxor g1447(.dina(n1500), .dinb(n1474), .dout(n1501));
  jor  g1448(.dina(n1501), .dinb(n1490), .dout(n1502));
  jnot g1449(.din(n1502), .dout(n1503));
  jnot g1450(.din(n519), .dout(n1504));
  jand g1451(.dina(n1474), .dinb(n1490), .dout(n1505));
  jand g1452(.dina(n1505), .dinb(n1504), .dout(n1506));
  jor  g1453(.dina(n1506), .dinb(n1503), .dout(n1507));
  jor  g1454(.dina(n1507), .dinb(n1497), .dout(n1508));
  jand g1455(.dina(n1508), .dinb(n1489), .dout(n1509));
  jnot g1456(.din(n1509), .dout(n1510));
  jor  g1457(.dina(n1508), .dinb(n1489), .dout(n1511));
  jand g1458(.dina(n1511), .dinb(n1478), .dout(n1512));
  jand g1459(.dina(n1512), .dinb(n1510), .dout(n1513));
  jor  g1460(.dina(n1513), .dinb(n1479), .dout(n1514));
  jnot g1461(.din(n1511), .dout(n1515));
  jor  g1462(.dina(n1513), .dinb(n1515), .dout(n1516));
  jor  g1463(.dina(n1516), .dinb(n1509), .dout(n1517));
  jand g1464(.dina(n1517), .dinb(n1514), .dout(n1518));
  jor  g1465(.dina(n1518), .dinb(n1432), .dout(n1519));
  jxor g1466(.dina(n1518), .dinb(n1432), .dout(n1520));
  jand g1467(.dina(n1425), .dinb(n1415), .dout(n1521));
  jand g1468(.dina(n1426), .dinb(n1407), .dout(n1522));
  jor  g1469(.dina(n1522), .dinb(n1521), .dout(n1523));
  jand g1470(.dina(n1360), .dinb(n1354), .dout(n1524));
  jnot g1471(.din(n1524), .dout(n1525));
  jand g1472(.dina(n1434), .dinb(n1353), .dout(n1526));
  jxor g1473(.dina(n1526), .dinb(n716), .dout(n1527));
  jand g1474(.dina(n1527), .dinb(n1525), .dout(n1528));
  jnot g1475(.din(n997), .dout(n1529));
  jand g1476(.dina(n1480), .dinb(n1529), .dout(n1530));
  jor  g1477(.dina(n876), .dinb(n930), .dout(n1531));
  jand g1478(.dina(n1531), .dinb(n987), .dout(n1532));
  jor  g1479(.dina(n813), .dinb(n716), .dout(n1533));
  jand g1480(.dina(n1533), .dinb(n1532), .dout(n1534));
  jand g1481(.dina(n1356), .dinb(n1534), .dout(n1535));
  jor  g1482(.dina(n1535), .dinb(n1530), .dout(n1536));
  jnot g1483(.din(n1536), .dout(n1537));
  jor  g1484(.dina(n1531), .dinb(n607), .dout(n1538));
  jand g1485(.dina(n1538), .dinb(n1533), .dout(n1539));
  jand g1486(.dina(n994), .dinb(n1539), .dout(n1540));
  jxor g1487(.dina(n876), .dinb(n930), .dout(n1541));
  jor  g1488(.dina(n1541), .dinb(n1532), .dout(n1542));
  jand g1489(.dina(n996), .dinb(n1542), .dout(n1543));
  jor  g1490(.dina(n1543), .dinb(n1540), .dout(n1544));
  jand g1491(.dina(n1544), .dinb(n1537), .dout(n1545));
  jand g1492(.dina(n1545), .dinb(n1528), .dout(n1546));
  jand g1493(.dina(n1400), .dinb(n1149), .dout(n1547));
  jnot g1494(.din(n1547), .dout(n1548));
  jand g1495(.dina(n1548), .dinb(n1402), .dout(n1549));
  jand g1496(.dina(n1549), .dinb(n1154), .dout(n1550));
  jand g1497(.dina(n1403), .dinb(n1491), .dout(n1551));
  jand g1498(.dina(n1551), .dinb(n1156), .dout(n1552));
  jor  g1499(.dina(n1552), .dinb(n1550), .dout(n1553));
  jnot g1500(.din(n1553), .dout(n1554));
  jnot g1501(.din(n1403), .dout(n1555));
  jor  g1502(.dina(n1547), .dinb(n486), .dout(n1556));
  jand g1503(.dina(n1556), .dinb(n1555), .dout(n1557));
  jnot g1504(.din(n1557), .dout(n1558));
  jand g1505(.dina(n1558), .dinb(n1499), .dout(n1559));
  jor  g1506(.dina(n1403), .dinb(n1402), .dout(n1560));
  jand g1507(.dina(n1560), .dinb(n1500), .dout(n1561));
  jor  g1508(.dina(n1561), .dinb(n1559), .dout(n1562));
  jand g1509(.dina(n1562), .dinb(n1554), .dout(n1563));
  jxor g1510(.dina(n1545), .dinb(n1528), .dout(n1564));
  jand g1511(.dina(n1564), .dinb(n1563), .dout(n1565));
  jor  g1512(.dina(n1565), .dinb(n1546), .dout(n1566));
  jxor g1513(.dina(n1566), .dinb(n1523), .dout(n1567));
  jand g1514(.dina(n1255), .dinb(n994), .dout(n1568));
  jand g1515(.dina(n1261), .dinb(n996), .dout(n1569));
  jor  g1516(.dina(n1569), .dinb(n1568), .dout(n1570));
  jnot g1517(.din(n1570), .dout(n1571));
  jand g1518(.dina(n1270), .dinb(n880), .dout(n1572));
  jand g1519(.dina(n1295), .dinb(n881), .dout(n1573));
  jor  g1520(.dina(n1573), .dinb(n1572), .dout(n1574));
  jand g1521(.dina(n1574), .dinb(n1571), .dout(n1575));
  jnot g1522(.din(n1170), .dout(n1576));
  jand g1523(.dina(n1259), .dinb(n1576), .dout(n1577));
  jand g1524(.dina(n1257), .dinb(n1163), .dout(n1578));
  jor  g1525(.dina(n1578), .dinb(n1577), .dout(n1579));
  jnot g1526(.din(n1579), .dout(n1580));
  jand g1527(.dina(n1266), .dinb(n1160), .dout(n1581));
  jand g1528(.dina(n1272), .dinb(n1152), .dout(n1582));
  jor  g1529(.dina(n1582), .dinb(n1581), .dout(n1583));
  jand g1530(.dina(n1583), .dinb(n1580), .dout(n1584));
  jand g1531(.dina(n1551), .dinb(n1168), .dout(n1585));
  jand g1532(.dina(n1549), .dinb(n1166), .dout(n1586));
  jor  g1533(.dina(n1586), .dinb(n1585), .dout(n1587));
  jnot g1534(.din(n1587), .dout(n1588));
  jand g1535(.dina(n1558), .dinb(n1154), .dout(n1589));
  jand g1536(.dina(n1560), .dinb(n1156), .dout(n1590));
  jor  g1537(.dina(n1590), .dinb(n1589), .dout(n1591));
  jand g1538(.dina(n1591), .dinb(n1588), .dout(n1592));
  jxor g1539(.dina(n1592), .dinb(n1584), .dout(n1593));
  jxor g1540(.dina(n1593), .dinb(n1575), .dout(n1594));
  jxor g1541(.dina(n1594), .dinb(n1567), .dout(n1595));
  jand g1542(.dina(n1595), .dinb(n1520), .dout(n1596));
  jnot g1543(.din(n1596), .dout(n1597));
  jand g1544(.dina(n1597), .dinb(n1519), .dout(n1598));
  jand g1545(.dina(n1566), .dinb(n1523), .dout(n1599));
  jand g1546(.dina(n1594), .dinb(n1567), .dout(n1600));
  jor  g1547(.dina(n1600), .dinb(n1599), .dout(n1601));
  jand g1548(.dina(n1592), .dinb(n1584), .dout(n1602));
  jand g1549(.dina(n1593), .dinb(n1575), .dout(n1603));
  jor  g1550(.dina(n1603), .dinb(n1602), .dout(n1604));
  jand g1551(.dina(n1494), .dinb(n1441), .dout(n1605));
  jand g1552(.dina(n1499), .dinb(n1493), .dout(n1606));
  jnot g1553(.din(n1606), .dout(n1607));
  jxor g1554(.dina(n1474), .dinb(n1156), .dout(n1608));
  jor  g1555(.dina(n1608), .dinb(n1490), .dout(n1609));
  jand g1556(.dina(n1505), .dinb(n1500), .dout(n1610));
  jnot g1557(.din(n1610), .dout(n1611));
  jand g1558(.dina(n1611), .dinb(n1609), .dout(n1612));
  jand g1559(.dina(n1612), .dinb(n1607), .dout(n1613));
  jxor g1560(.dina(n1613), .dinb(n1605), .dout(n1614));
  jxor g1561(.dina(n1614), .dinb(n1604), .dout(n1615));
  jxor g1562(.dina(n1615), .dinb(n1601), .dout(n1616));
  jand g1563(.dina(n1485), .dinb(n878), .dout(n1617));
  jand g1564(.dina(n1360), .dinb(n989), .dout(n1618));
  jor  g1565(.dina(n1618), .dinb(n1617), .dout(n1619));
  jnot g1566(.din(n1619), .dout(n1620));
  jand g1567(.dina(n1434), .dinb(n992), .dout(n1621));
  jnot g1568(.din(n1434), .dout(n1622));
  jand g1569(.dina(n1622), .dinb(n997), .dout(n1623));
  jor  g1570(.dina(n1623), .dinb(n1621), .dout(n1624));
  jand g1571(.dina(n1624), .dinb(n1620), .dout(n1625));
  jand g1572(.dina(n1494), .dinb(n519), .dout(n1626));
  jand g1573(.dina(n1438), .dinb(n1354), .dout(n1627));
  jor  g1574(.dina(n1627), .dinb(n930), .dout(n1628));
  jnot g1575(.din(n1628), .dout(n1629));
  jxor g1576(.dina(n1629), .dinb(n1626), .dout(n1630));
  jxor g1577(.dina(n1630), .dinb(n1625), .dout(n1631));
  jxor g1578(.dina(n1631), .dinb(n1516), .dout(n1632));
  jand g1579(.dina(n1551), .dinb(n1272), .dout(n1633));
  jand g1580(.dina(n1549), .dinb(n1266), .dout(n1634));
  jor  g1581(.dina(n1634), .dinb(n1633), .dout(n1635));
  jnot g1582(.din(n1635), .dout(n1636));
  jand g1583(.dina(n1558), .dinb(n1166), .dout(n1637));
  jand g1584(.dina(n1560), .dinb(n1168), .dout(n1638));
  jor  g1585(.dina(n1638), .dinb(n1637), .dout(n1639));
  jand g1586(.dina(n1639), .dinb(n1636), .dout(n1640));
  jand g1587(.dina(n1259), .dinb(n1416), .dout(n1641));
  jand g1588(.dina(n1257), .dinb(n1418), .dout(n1642));
  jor  g1589(.dina(n1642), .dinb(n1641), .dout(n1643));
  jnot g1590(.din(n1643), .dout(n1644));
  jand g1591(.dina(n1164), .dinb(n880), .dout(n1645));
  jand g1592(.dina(n1170), .dinb(n881), .dout(n1646));
  jor  g1593(.dina(n1646), .dinb(n1645), .dout(n1647));
  jand g1594(.dina(n1647), .dinb(n1644), .dout(n1648));
  jnot g1595(.din(n1295), .dout(n1649));
  jand g1596(.dina(n1649), .dinb(n996), .dout(n1650));
  jnot g1597(.din(n1270), .dout(n1651));
  jand g1598(.dina(n1651), .dinb(n994), .dout(n1652));
  jor  g1599(.dina(n1652), .dinb(n1650), .dout(n1653));
  jnot g1600(.din(n1653), .dout(n1654));
  jand g1601(.dina(n1356), .dinb(n1254), .dout(n1655));
  jnot g1602(.din(n1261), .dout(n1656));
  jand g1603(.dina(n1480), .dinb(n1656), .dout(n1657));
  jor  g1604(.dina(n1657), .dinb(n1655), .dout(n1658));
  jand g1605(.dina(n1658), .dinb(n1654), .dout(n1659));
  jxor g1606(.dina(n1659), .dinb(n1648), .dout(n1660));
  jxor g1607(.dina(n1660), .dinb(n1640), .dout(n1661));
  jxor g1608(.dina(n1661), .dinb(n1632), .dout(n1662));
  jxor g1609(.dina(n1662), .dinb(n1616), .dout(n1663));
  jxor g1610(.dina(n1663), .dinb(n1598), .dout(n1664));
  jand g1611(.dina(n1551), .dinb(n1500), .dout(n1665));
  jand g1612(.dina(n1549), .dinb(n1499), .dout(n1666));
  jor  g1613(.dina(n1666), .dinb(n1665), .dout(n1667));
  jnot g1614(.din(n1667), .dout(n1668));
  jor  g1615(.dina(n1557), .dinb(n1504), .dout(n1669));
  jnot g1616(.din(n1669), .dout(n1670));
  jand g1617(.dina(n1560), .dinb(n1504), .dout(n1671));
  jor  g1618(.dina(n1671), .dinb(n1670), .dout(n1672));
  jand g1619(.dina(n1672), .dinb(n1668), .dout(n1673));
  jxor g1620(.dina(n1406), .dinb(n1363), .dout(n1674));
  jand g1621(.dina(n1674), .dinb(n1673), .dout(n1675));
  jand g1622(.dina(n1354), .dinb(n994), .dout(n1676));
  jnot g1623(.din(n1676), .dout(n1677));
  jand g1624(.dina(n1356), .dinb(n1353), .dout(n1678));
  jxor g1625(.dina(n1678), .dinb(n716), .dout(n1679));
  jand g1626(.dina(n1679), .dinb(n1677), .dout(n1680));
  jor  g1627(.dina(n1257), .dinb(n1542), .dout(n1681));
  jor  g1628(.dina(n1259), .dinb(n1539), .dout(n1682));
  jand g1629(.dina(n1682), .dinb(n1681), .dout(n1683));
  jand g1630(.dina(n992), .dinb(n880), .dout(n1684));
  jand g1631(.dina(n997), .dinb(n881), .dout(n1685));
  jor  g1632(.dina(n1685), .dinb(n1684), .dout(n1686));
  jand g1633(.dina(n1686), .dinb(n1683), .dout(n1687));
  jand g1634(.dina(n1687), .dinb(n1680), .dout(n1688));
  jand g1635(.dina(n1266), .dinb(n1255), .dout(n1689));
  jand g1636(.dina(n1272), .dinb(n1261), .dout(n1690));
  jor  g1637(.dina(n1690), .dinb(n1689), .dout(n1691));
  jnot g1638(.din(n1691), .dout(n1692));
  jand g1639(.dina(n1270), .dinb(n1166), .dout(n1693));
  jand g1640(.dina(n1295), .dinb(n1168), .dout(n1694));
  jor  g1641(.dina(n1694), .dinb(n1693), .dout(n1695));
  jand g1642(.dina(n1695), .dinb(n1692), .dout(n1696));
  jxor g1643(.dina(n1687), .dinb(n1680), .dout(n1697));
  jand g1644(.dina(n1697), .dinb(n1696), .dout(n1698));
  jor  g1645(.dina(n1698), .dinb(n1688), .dout(n1699));
  jxor g1646(.dina(n1674), .dinb(n1673), .dout(n1700));
  jand g1647(.dina(n1700), .dinb(n1699), .dout(n1701));
  jor  g1648(.dina(n1701), .dinb(n1675), .dout(n1702));
  jxor g1649(.dina(n1564), .dinb(n1563), .dout(n1703));
  jand g1650(.dina(n1703), .dinb(n1702), .dout(n1704));
  jxor g1651(.dina(n1429), .dinb(n1427), .dout(n1705));
  jxor g1652(.dina(n1703), .dinb(n1702), .dout(n1706));
  jand g1653(.dina(n1706), .dinb(n1705), .dout(n1707));
  jor  g1654(.dina(n1707), .dinb(n1704), .dout(n1708));
  jxor g1655(.dina(n1595), .dinb(n1520), .dout(n1709));
  jand g1656(.dina(n1709), .dinb(n1708), .dout(n1710));
  jnot g1657(.din(n1710), .dout(n1711));
  jor  g1658(.dina(n1266), .dinb(n1542), .dout(n1712));
  jor  g1659(.dina(n1272), .dinb(n1539), .dout(n1713));
  jand g1660(.dina(n1713), .dinb(n1712), .dout(n1714));
  jand g1661(.dina(n1257), .dinb(n992), .dout(n1715));
  jand g1662(.dina(n1259), .dinb(n997), .dout(n1716));
  jor  g1663(.dina(n1716), .dinb(n1715), .dout(n1717));
  jand g1664(.dina(n1717), .dinb(n1714), .dout(n1718));
  jor  g1665(.dina(n1254), .dinb(n1168), .dout(n1719));
  jor  g1666(.dina(n1656), .dinb(n1166), .dout(n1720));
  jand g1667(.dina(n1720), .dinb(n1719), .dout(n1721));
  jand g1668(.dina(n1270), .dinb(n1154), .dout(n1722));
  jand g1669(.dina(n1295), .dinb(n1156), .dout(n1723));
  jor  g1670(.dina(n1723), .dinb(n1722), .dout(n1724));
  jand g1671(.dina(n1724), .dinb(n1721), .dout(n1725));
  jand g1672(.dina(n1725), .dinb(n1718), .dout(n1726));
  jor  g1673(.dina(n1499), .dinb(n1170), .dout(n1727));
  jor  g1674(.dina(n1500), .dinb(n1164), .dout(n1728));
  jand g1675(.dina(n1728), .dinb(n1727), .dout(n1729));
  jand g1676(.dina(n1160), .dinb(n519), .dout(n1730));
  jand g1677(.dina(n1152), .dinb(n1504), .dout(n1731));
  jor  g1678(.dina(n1731), .dinb(n1730), .dout(n1732));
  jand g1679(.dina(n1732), .dinb(n1729), .dout(n1733));
  jxor g1680(.dina(n1725), .dinb(n1718), .dout(n1734));
  jand g1681(.dina(n1734), .dinb(n1733), .dout(n1735));
  jor  g1682(.dina(n1735), .dinb(n1726), .dout(n1736));
  jxor g1683(.dina(n1697), .dinb(n1696), .dout(n1737));
  jand g1684(.dina(n1737), .dinb(n1736), .dout(n1738));
  jand g1685(.dina(n1354), .dinb(n880), .dout(n1739));
  jnot g1686(.din(n1739), .dout(n1740));
  jand g1687(.dina(n1353), .dinb(n994), .dout(n1741));
  jxor g1688(.dina(n1741), .dinb(n716), .dout(n1742));
  jand g1689(.dina(n1742), .dinb(n1740), .dout(n1743));
  jand g1690(.dina(n1115), .dinb(n519), .dout(n1744));
  jnot g1691(.din(n1744), .dout(n1745));
  jand g1692(.dina(n1745), .dinb(n1151), .dout(n1746));
  jand g1693(.dina(n1746), .dinb(n1743), .dout(n1747));
  jor  g1694(.dina(n1499), .dinb(n1152), .dout(n1748));
  jor  g1695(.dina(n1500), .dinb(n1160), .dout(n1749));
  jand g1696(.dina(n1749), .dinb(n1748), .dout(n1750));
  jand g1697(.dina(n1164), .dinb(n1154), .dout(n1751));
  jand g1698(.dina(n1170), .dinb(n1156), .dout(n1752));
  jor  g1699(.dina(n1752), .dinb(n1751), .dout(n1753));
  jand g1700(.dina(n1753), .dinb(n1750), .dout(n1754));
  jxor g1701(.dina(n1754), .dinb(n1747), .dout(n1755));
  jxor g1702(.dina(n1755), .dinb(n1404), .dout(n1756));
  jxor g1703(.dina(n1737), .dinb(n1736), .dout(n1757));
  jand g1704(.dina(n1757), .dinb(n1756), .dout(n1758));
  jor  g1705(.dina(n1758), .dinb(n1738), .dout(n1759));
  jnot g1706(.din(n1759), .dout(n1760));
  jand g1707(.dina(n1754), .dinb(n1747), .dout(n1761));
  jand g1708(.dina(n1755), .dinb(n1404), .dout(n1762));
  jor  g1709(.dina(n1762), .dinb(n1761), .dout(n1763));
  jxor g1710(.dina(n1300), .dinb(n1299), .dout(n1764));
  jxor g1711(.dina(n1764), .dinb(n1763), .dout(n1765));
  jxor g1712(.dina(n1700), .dinb(n1699), .dout(n1766));
  jxor g1713(.dina(n1766), .dinb(n1765), .dout(n1767));
  jnot g1714(.din(n1767), .dout(n1768));
  jxor g1715(.dina(n1746), .dinb(n1743), .dout(n1769));
  jnot g1716(.din(n1769), .dout(n1770));
  jand g1717(.dina(n1168), .dinb(n878), .dout(n1771));
  jand g1718(.dina(n1166), .dinb(n989), .dout(n1772));
  jor  g1719(.dina(n1772), .dinb(n1771), .dout(n1773));
  jand g1720(.dina(n1266), .dinb(n992), .dout(n1774));
  jand g1721(.dina(n1272), .dinb(n997), .dout(n1775));
  jor  g1722(.dina(n1775), .dinb(n1774), .dout(n1776));
  jnot g1723(.din(n1776), .dout(n1777));
  jor  g1724(.dina(n1777), .dinb(n1773), .dout(n1778));
  jand g1725(.dina(n1354), .dinb(n1257), .dout(n1779));
  jnot g1726(.din(n1779), .dout(n1780));
  jand g1727(.dina(n1353), .dinb(n880), .dout(n1781));
  jxor g1728(.dina(n1781), .dinb(n716), .dout(n1782));
  jand g1729(.dina(n1782), .dinb(n1780), .dout(n1783));
  jnot g1730(.din(n1783), .dout(n1784));
  jor  g1731(.dina(n1784), .dinb(n1778), .dout(n1785));
  jand g1732(.dina(n1255), .dinb(n1154), .dout(n1786));
  jand g1733(.dina(n1261), .dinb(n1156), .dout(n1787));
  jor  g1734(.dina(n1787), .dinb(n1786), .dout(n1788));
  jand g1735(.dina(n1499), .dinb(n1270), .dout(n1789));
  jand g1736(.dina(n1500), .dinb(n1295), .dout(n1790));
  jor  g1737(.dina(n1790), .dinb(n1789), .dout(n1791));
  jnot g1738(.din(n1791), .dout(n1792));
  jor  g1739(.dina(n1792), .dinb(n1788), .dout(n1793));
  jxor g1740(.dina(n1783), .dinb(n1778), .dout(n1794));
  jor  g1741(.dina(n1794), .dinb(n1793), .dout(n1795));
  jand g1742(.dina(n1795), .dinb(n1785), .dout(n1796));
  jor  g1743(.dina(n1796), .dinb(n1770), .dout(n1797));
  jnot g1744(.din(n1797), .dout(n1798));
  jxor g1745(.dina(n1796), .dinb(n1770), .dout(n1799));
  jxor g1746(.dina(n1734), .dinb(n1733), .dout(n1800));
  jand g1747(.dina(n1800), .dinb(n1799), .dout(n1801));
  jor  g1748(.dina(n1801), .dinb(n1798), .dout(n1802));
  jnot g1749(.din(n1802), .dout(n1803));
  jxor g1750(.dina(n1757), .dinb(n1756), .dout(n1804));
  jnot g1751(.din(n1804), .dout(n1805));
  jand g1752(.dina(n1805), .dinb(n1803), .dout(n1806));
  jand g1753(.dina(n1354), .dinb(n1266), .dout(n1807));
  jnot g1754(.din(n1807), .dout(n1808));
  jand g1755(.dina(n1353), .dinb(n1257), .dout(n1809));
  jxor g1756(.dina(n1809), .dinb(n716), .dout(n1810));
  jand g1757(.dina(n1810), .dinb(n1808), .dout(n1811));
  jnot g1758(.din(n1260), .dout(n1812));
  jor  g1759(.dina(n1812), .dinb(n1504), .dout(n1813));
  jand g1760(.dina(n1813), .dinb(n1294), .dout(n1814));
  jand g1761(.dina(n1814), .dinb(n1811), .dout(n1815));
  jand g1762(.dina(n1815), .dinb(n1744), .dout(n1816));
  jor  g1763(.dina(n1168), .dinb(n992), .dout(n1817));
  jor  g1764(.dina(n1166), .dinb(n997), .dout(n1818));
  jand g1765(.dina(n1818), .dinb(n1817), .dout(n1819));
  jand g1766(.dina(n1154), .dinb(n1539), .dout(n1820));
  jand g1767(.dina(n1156), .dinb(n1542), .dout(n1821));
  jor  g1768(.dina(n1821), .dinb(n1820), .dout(n1822));
  jand g1769(.dina(n1822), .dinb(n1819), .dout(n1823));
  jor  g1770(.dina(n1295), .dinb(n519), .dout(n1824));
  jor  g1771(.dina(n1270), .dinb(n1504), .dout(n1825));
  jand g1772(.dina(n1825), .dinb(n1824), .dout(n1826));
  jand g1773(.dina(n1499), .dinb(n1254), .dout(n1827));
  jand g1774(.dina(n1500), .dinb(n1656), .dout(n1828));
  jor  g1775(.dina(n1828), .dinb(n1827), .dout(n1829));
  jand g1776(.dina(n1829), .dinb(n1826), .dout(n1830));
  jand g1777(.dina(n1830), .dinb(n1823), .dout(n1831));
  jxor g1778(.dina(n1814), .dinb(n1811), .dout(n1832));
  jxor g1779(.dina(n1830), .dinb(n1823), .dout(n1833));
  jand g1780(.dina(n1833), .dinb(n1832), .dout(n1834));
  jor  g1781(.dina(n1834), .dinb(n1831), .dout(n1835));
  jxor g1782(.dina(n1815), .dinb(n1744), .dout(n1836));
  jand g1783(.dina(n1836), .dinb(n1835), .dout(n1837));
  jor  g1784(.dina(n1837), .dinb(n1816), .dout(n1838));
  jxor g1785(.dina(n1800), .dinb(n1799), .dout(n1839));
  jor  g1786(.dina(n1839), .dinb(n1838), .dout(n1840));
  jnot g1787(.din(n1840), .dout(n1841));
  jxor g1788(.dina(n1836), .dinb(n1835), .dout(n1842));
  jxor g1789(.dina(n1794), .dinb(n1793), .dout(n1843));
  jand g1790(.dina(n1843), .dinb(n1842), .dout(n1844));
  jnot g1791(.din(n1844), .dout(n1845));
  jor  g1792(.dina(n1843), .dinb(n1842), .dout(n1846));
  jnot g1793(.din(n1846), .dout(n1847));
  jand g1794(.dina(n877), .dinb(n519), .dout(n1848));
  jnot g1795(.din(n1848), .dout(n1849));
  jand g1796(.dina(n1541), .dinb(n519), .dout(n1850));
  jand g1797(.dina(n1850), .dinb(n1353), .dout(n1851));
  jand g1798(.dina(n1500), .dinb(n716), .dout(n1852));
  jor  g1799(.dina(n1852), .dinb(n1851), .dout(n1853));
  jand g1800(.dina(n1156), .dinb(n930), .dout(n1854));
  jand g1801(.dina(n1154), .dinb(n716), .dout(n1855));
  jand g1802(.dina(n1855), .dinb(n1353), .dout(n1856));
  jor  g1803(.dina(n1856), .dinb(n1854), .dout(n1857));
  jnot g1804(.din(n1857), .dout(n1858));
  jand g1805(.dina(n1858), .dinb(n1853), .dout(n1859));
  jand g1806(.dina(n1859), .dinb(n1849), .dout(n1860));
  jnot g1807(.din(n1860), .dout(n1861));
  jor  g1808(.dina(n1353), .dinb(n1156), .dout(n1862));
  jand g1809(.dina(n1353), .dinb(n1166), .dout(n1863));
  jxor g1810(.dina(n1863), .dinb(n716), .dout(n1864));
  jand g1811(.dina(n1864), .dinb(n1862), .dout(n1865));
  jor  g1812(.dina(n1850), .dinb(n815), .dout(n1866));
  jnot g1813(.din(n1866), .dout(n1867));
  jxor g1814(.dina(n1867), .dinb(n1865), .dout(n1868));
  jnot g1815(.din(n1868), .dout(n1869));
  jor  g1816(.dina(n878), .dinb(n519), .dout(n1870));
  jor  g1817(.dina(n989), .dinb(n1504), .dout(n1871));
  jand g1818(.dina(n1871), .dinb(n1870), .dout(n1872));
  jor  g1819(.dina(n1499), .dinb(n997), .dout(n1873));
  jnot g1820(.din(n1873), .dout(n1874));
  jand g1821(.dina(n1499), .dinb(n1534), .dout(n1875));
  jor  g1822(.dina(n1875), .dinb(n1874), .dout(n1876));
  jor  g1823(.dina(n1876), .dinb(n1872), .dout(n1877));
  jor  g1824(.dina(n1877), .dinb(n1869), .dout(n1878));
  jand g1825(.dina(n1878), .dinb(n1861), .dout(n1879));
  jand g1826(.dina(n1542), .dinb(n1504), .dout(n1880));
  jand g1827(.dina(n1539), .dinb(n519), .dout(n1881));
  jor  g1828(.dina(n1881), .dinb(n1880), .dout(n1882));
  jor  g1829(.dina(n1500), .dinb(n992), .dout(n1883));
  jand g1830(.dina(n1883), .dinb(n1873), .dout(n1884));
  jand g1831(.dina(n1884), .dinb(n1882), .dout(n1885));
  jor  g1832(.dina(n1885), .dinb(n1868), .dout(n1886));
  jnot g1833(.din(n1886), .dout(n1887));
  jor  g1834(.dina(n1887), .dinb(n1879), .dout(n1888));
  jor  g1835(.dina(n1888), .dinb(n1813), .dout(n1889));
  jand g1836(.dina(n1867), .dinb(n1865), .dout(n1890));
  jand g1837(.dina(n1354), .dinb(n1166), .dout(n1891));
  jnot g1838(.din(n1891), .dout(n1892));
  jand g1839(.dina(n1353), .dinb(n1266), .dout(n1893));
  jxor g1840(.dina(n1893), .dinb(n716), .dout(n1894));
  jand g1841(.dina(n1894), .dinb(n1892), .dout(n1895));
  jor  g1842(.dina(n1500), .dinb(n1539), .dout(n1896));
  jor  g1843(.dina(n1499), .dinb(n1542), .dout(n1897));
  jand g1844(.dina(n1897), .dinb(n1896), .dout(n1898));
  jand g1845(.dina(n1154), .dinb(n992), .dout(n1899));
  jand g1846(.dina(n1156), .dinb(n997), .dout(n1900));
  jor  g1847(.dina(n1900), .dinb(n1899), .dout(n1901));
  jand g1848(.dina(n1901), .dinb(n1898), .dout(n1902));
  jxor g1849(.dina(n1902), .dinb(n1895), .dout(n1903));
  jxor g1850(.dina(n1903), .dinb(n1890), .dout(n1904));
  jnot g1851(.din(n1904), .dout(n1905));
  jand g1852(.dina(n1905), .dinb(n1889), .dout(n1906));
  jand g1853(.dina(n1888), .dinb(n1813), .dout(n1907));
  jxor g1854(.dina(n1833), .dinb(n1832), .dout(n1908));
  jnot g1855(.din(n1908), .dout(n1909));
  jand g1856(.dina(n1902), .dinb(n1895), .dout(n1910));
  jnot g1857(.din(n1910), .dout(n1911));
  jnot g1858(.din(n1890), .dout(n1912));
  jnot g1859(.din(n1895), .dout(n1913));
  jxor g1860(.dina(n1902), .dinb(n1913), .dout(n1914));
  jor  g1861(.dina(n1914), .dinb(n1912), .dout(n1915));
  jand g1862(.dina(n1915), .dinb(n1911), .dout(n1916));
  jand g1863(.dina(n1916), .dinb(n1909), .dout(n1917));
  jor  g1864(.dina(n1917), .dinb(n1907), .dout(n1918));
  jor  g1865(.dina(n1918), .dinb(n1906), .dout(n1919));
  jand g1866(.dina(n1903), .dinb(n1890), .dout(n1920));
  jor  g1867(.dina(n1920), .dinb(n1910), .dout(n1921));
  jand g1868(.dina(n1921), .dinb(n1908), .dout(n1922));
  jnot g1869(.din(n1922), .dout(n1923));
  jand g1870(.dina(n1923), .dinb(n1919), .dout(n1924));
  jor  g1871(.dina(n1924), .dinb(n1847), .dout(n1925));
  jand g1872(.dina(n1925), .dinb(n1845), .dout(n1926));
  jor  g1873(.dina(n1926), .dinb(n1841), .dout(n1927));
  jand g1874(.dina(n1804), .dinb(n1802), .dout(n1928));
  jand g1875(.dina(n1839), .dinb(n1838), .dout(n1929));
  jor  g1876(.dina(n1929), .dinb(n1928), .dout(n1930));
  jnot g1877(.din(n1930), .dout(n1931));
  jand g1878(.dina(n1931), .dinb(n1927), .dout(n1932));
  jor  g1879(.dina(n1932), .dinb(n1806), .dout(n1933));
  jand g1880(.dina(n1933), .dinb(n1768), .dout(n1934));
  jor  g1881(.dina(n1934), .dinb(n1760), .dout(n1935));
  jand g1882(.dina(n1764), .dinb(n1763), .dout(n1936));
  jand g1883(.dina(n1766), .dinb(n1765), .dout(n1937));
  jor  g1884(.dina(n1937), .dinb(n1936), .dout(n1938));
  jxor g1885(.dina(n1706), .dinb(n1705), .dout(n1939));
  jand g1886(.dina(n1939), .dinb(n1938), .dout(n1940));
  jnot g1887(.din(n1940), .dout(n1941));
  jor  g1888(.dina(n1933), .dinb(n1768), .dout(n1942));
  jand g1889(.dina(n1942), .dinb(n1941), .dout(n1943));
  jand g1890(.dina(n1943), .dinb(n1935), .dout(n1944));
  jnot g1891(.din(n1938), .dout(n1945));
  jnot g1892(.din(n1939), .dout(n1946));
  jand g1893(.dina(n1946), .dinb(n1945), .dout(n1947));
  jnot g1894(.din(n1947), .dout(n1948));
  jor  g1895(.dina(n1709), .dinb(n1708), .dout(n1949));
  jand g1896(.dina(n1949), .dinb(n1948), .dout(n1950));
  jnot g1897(.din(n1950), .dout(n1951));
  jor  g1898(.dina(n1951), .dinb(n1944), .dout(n1952));
  jand g1899(.dina(n1952), .dinb(n1711), .dout(n1953));
  jxor g1900(.dina(n1953), .dinb(n1664), .dout(n1954));
  jxor g1901(.dina(n1954), .dinb(n425), .dout(n1955));
  jnot g1902(.din(n1955), .dout(n1956));
  jxor g1903(.dina(n1360), .dinb(n1480), .dout(n1957));
  jnot g1904(.din(n1957), .dout(n1958));
  jand g1905(.dina(n1958), .dinb(n1956), .dout(n1959));
  jand g1906(.dina(n1954), .dinb(n425), .dout(n1960));
  jand g1907(.dina(n445), .dinb(n327), .dout(n1961));
  jand g1908(.dina(n337), .dinb(n215), .dout(n1962));
  jand g1909(.dina(n467), .dinb(n147), .dout(n1963));
  jand g1910(.dina(n1963), .dinb(n1962), .dout(n1964));
  jand g1911(.dina(n1964), .dinb(n924), .dout(n1965));
  jand g1912(.dina(n1965), .dinb(n526), .dout(n1966));
  jand g1913(.dina(n534), .dinb(n290), .dout(n1967));
  jand g1914(.dina(n462), .dinb(n176), .dout(n1968));
  jand g1915(.dina(n1968), .dinb(n353), .dout(n1969));
  jand g1916(.dina(n1969), .dinb(n1967), .dout(n1970));
  jand g1917(.dina(n510), .dinb(n415), .dout(n1971));
  jand g1918(.dina(n1971), .dinb(n460), .dout(n1972));
  jand g1919(.dina(n1972), .dinb(n1970), .dout(n1973));
  jand g1920(.dina(n1973), .dinb(n1966), .dout(n1974));
  jand g1921(.dina(n1974), .dinb(n1961), .dout(n1975));
  jand g1922(.dina(n1087), .dinb(n297), .dout(n1976));
  jand g1923(.dina(n321), .dinb(n213), .dout(n1977));
  jand g1924(.dina(n1977), .dinb(n1005), .dout(n1978));
  jand g1925(.dina(n188), .dinb(n157), .dout(n1979));
  jand g1926(.dina(n1979), .dinb(n1978), .dout(n1980));
  jand g1927(.dina(n1980), .dinb(n1976), .dout(n1981));
  jand g1928(.dina(n1024), .dinb(n276), .dout(n1982));
  jand g1929(.dina(n546), .dinb(n207), .dout(n1983));
  jand g1930(.dina(n448), .dinb(n389), .dout(n1984));
  jand g1931(.dina(n1984), .dinb(n588), .dout(n1985));
  jand g1932(.dina(n1985), .dinb(n1983), .dout(n1986));
  jand g1933(.dina(n1986), .dinb(n1982), .dout(n1987));
  jand g1934(.dina(n437), .dinb(n103), .dout(n1988));
  jand g1935(.dina(n1988), .dinb(n383), .dout(n1989));
  jand g1936(.dina(n1989), .dinb(n1987), .dout(n1990));
  jand g1937(.dina(n1990), .dinb(n489), .dout(n1991));
  jand g1938(.dina(n1991), .dinb(n1981), .dout(n1992));
  jand g1939(.dina(n1992), .dinb(n1975), .dout(n1993));
  jnot g1940(.din(n1993), .dout(n1994));
  jnot g1941(.din(n1598), .dout(n1995));
  jand g1942(.dina(n1663), .dinb(n1995), .dout(n1996));
  jnot g1943(.din(n1664), .dout(n1997));
  jnot g1944(.din(n1806), .dout(n1998));
  jnot g1945(.din(n1813), .dout(n1999));
  jand g1946(.dina(n1885), .dinb(n1868), .dout(n2000));
  jor  g1947(.dina(n2000), .dinb(n1860), .dout(n2001));
  jand g1948(.dina(n1886), .dinb(n2001), .dout(n2002));
  jand g1949(.dina(n2002), .dinb(n1999), .dout(n2003));
  jor  g1950(.dina(n1904), .dinb(n2003), .dout(n2004));
  jor  g1951(.dina(n2002), .dinb(n1999), .dout(n2005));
  jor  g1952(.dina(n1921), .dinb(n1908), .dout(n2006));
  jand g1953(.dina(n2006), .dinb(n2005), .dout(n2007));
  jand g1954(.dina(n2007), .dinb(n2004), .dout(n2008));
  jor  g1955(.dina(n1922), .dinb(n2008), .dout(n2009));
  jand g1956(.dina(n2009), .dinb(n1846), .dout(n2010));
  jor  g1957(.dina(n2010), .dinb(n1844), .dout(n2011));
  jand g1958(.dina(n2011), .dinb(n1840), .dout(n2012));
  jor  g1959(.dina(n1930), .dinb(n2012), .dout(n2013));
  jand g1960(.dina(n2013), .dinb(n1998), .dout(n2014));
  jor  g1961(.dina(n2014), .dinb(n1767), .dout(n2015));
  jand g1962(.dina(n2015), .dinb(n1759), .dout(n2016));
  jand g1963(.dina(n2014), .dinb(n1767), .dout(n2017));
  jor  g1964(.dina(n2017), .dinb(n1940), .dout(n2018));
  jor  g1965(.dina(n2018), .dinb(n2016), .dout(n2019));
  jand g1966(.dina(n1950), .dinb(n2019), .dout(n2020));
  jor  g1967(.dina(n2020), .dinb(n1710), .dout(n2021));
  jand g1968(.dina(n2021), .dinb(n1997), .dout(n2022));
  jor  g1969(.dina(n2022), .dinb(n1996), .dout(n2023));
  jand g1970(.dina(n1615), .dinb(n1601), .dout(n2024));
  jand g1971(.dina(n1662), .dinb(n1616), .dout(n2025));
  jor  g1972(.dina(n2025), .dinb(n2024), .dout(n2026));
  jand g1973(.dina(n1631), .dinb(n1516), .dout(n2027));
  jand g1974(.dina(n1661), .dinb(n1632), .dout(n2028));
  jor  g1975(.dina(n2028), .dinb(n2027), .dout(n2029));
  jand g1976(.dina(n1493), .dinb(n1154), .dout(n2030));
  jnot g1977(.din(n2030), .dout(n2031));
  jxor g1978(.dina(n1474), .dinb(n1168), .dout(n2032));
  jor  g1979(.dina(n2032), .dinb(n1490), .dout(n2033));
  jand g1980(.dina(n1505), .dinb(n1156), .dout(n2034));
  jnot g1981(.din(n2034), .dout(n2035));
  jand g1982(.dina(n2035), .dinb(n2033), .dout(n2036));
  jand g1983(.dina(n2036), .dinb(n2031), .dout(n2037));
  jand g1984(.dina(n1629), .dinb(n1626), .dout(n2038));
  jand g1985(.dina(n1630), .dinb(n1625), .dout(n2039));
  jor  g1986(.dina(n2039), .dinb(n2038), .dout(n2040));
  jxor g1987(.dina(n2040), .dinb(n2037), .dout(n2041));
  jand g1988(.dina(n1659), .dinb(n1648), .dout(n2042));
  jand g1989(.dina(n1660), .dinb(n1640), .dout(n2043));
  jor  g1990(.dina(n2043), .dinb(n2042), .dout(n2044));
  jxor g1991(.dina(n2044), .dinb(n2041), .dout(n2045));
  jxor g1992(.dina(n2045), .dinb(n2029), .dout(n2046));
  jand g1993(.dina(n1613), .dinb(n1605), .dout(n2047));
  jand g1994(.dina(n1614), .dinb(n1604), .dout(n2048));
  jor  g1995(.dina(n2048), .dinb(n2047), .dout(n2049));
  jand g1996(.dina(n1438), .dinb(n1534), .dout(n2050));
  jnot g1997(.din(n1438), .dout(n2051));
  jand g1998(.dina(n2051), .dinb(n1529), .dout(n2052));
  jor  g1999(.dina(n2052), .dinb(n2050), .dout(n2053));
  jnot g2000(.din(n2053), .dout(n2054));
  jand g2001(.dina(n1434), .dinb(n1539), .dout(n2055));
  jand g2002(.dina(n1622), .dinb(n1542), .dout(n2056));
  jor  g2003(.dina(n2056), .dinb(n2055), .dout(n2057));
  jand g2004(.dina(n2057), .dinb(n2054), .dout(n2058));
  jand g2005(.dina(n1499), .dinb(n1494), .dout(n2059));
  jxor g2006(.dina(n2059), .dinb(n716), .dout(n2060));
  jxor g2007(.dina(n2060), .dinb(n2058), .dout(n2061));
  jxor g2008(.dina(n2061), .dinb(n2049), .dout(n2062));
  jand g2009(.dina(n1551), .dinb(n1259), .dout(n2063));
  jand g2010(.dina(n1549), .dinb(n1257), .dout(n2064));
  jor  g2011(.dina(n2064), .dinb(n2063), .dout(n2065));
  jnot g2012(.din(n2065), .dout(n2066));
  jand g2013(.dina(n1558), .dinb(n1266), .dout(n2067));
  jand g2014(.dina(n1560), .dinb(n1272), .dout(n2068));
  jor  g2015(.dina(n2068), .dinb(n2067), .dout(n2069));
  jand g2016(.dina(n2069), .dinb(n2066), .dout(n2070));
  jand g2017(.dina(n1416), .dinb(n881), .dout(n2071));
  jand g2018(.dina(n1418), .dinb(n880), .dout(n2072));
  jor  g2019(.dina(n2072), .dinb(n2071), .dout(n2073));
  jnot g2020(.din(n2073), .dout(n2074));
  jand g2021(.dina(n1164), .dinb(n994), .dout(n2075));
  jand g2022(.dina(n1170), .dinb(n996), .dout(n2076));
  jor  g2023(.dina(n2076), .dinb(n2075), .dout(n2077));
  jand g2024(.dina(n2077), .dinb(n2074), .dout(n2078));
  jand g2025(.dina(n1480), .dinb(n1649), .dout(n2079));
  jand g2026(.dina(n1356), .dinb(n1651), .dout(n2080));
  jor  g2027(.dina(n2080), .dinb(n2079), .dout(n2081));
  jnot g2028(.din(n2081), .dout(n2082));
  jand g2029(.dina(n1360), .dinb(n1254), .dout(n2083));
  jand g2030(.dina(n1485), .dinb(n1656), .dout(n2084));
  jor  g2031(.dina(n2084), .dinb(n2083), .dout(n2085));
  jand g2032(.dina(n2085), .dinb(n2082), .dout(n2086));
  jxor g2033(.dina(n2086), .dinb(n2078), .dout(n2087));
  jxor g2034(.dina(n2087), .dinb(n2070), .dout(n2088));
  jxor g2035(.dina(n2088), .dinb(n2062), .dout(n2089));
  jxor g2036(.dina(n2089), .dinb(n2046), .dout(n2090));
  jxor g2037(.dina(n2090), .dinb(n2026), .dout(n2091));
  jxor g2038(.dina(n2091), .dinb(n2023), .dout(n2092));
  jxor g2039(.dina(n2092), .dinb(n1994), .dout(n2093));
  jxor g2040(.dina(n2093), .dinb(n1960), .dout(n2094));
  jxor g2041(.dina(n2094), .dinb(n1955), .dout(n2095));
  jnot g2042(.din(n2095), .dout(n2096));
  jxor g2043(.dina(n1259), .dinb(n880), .dout(n2097));
  jnot g2044(.din(n2097), .dout(n2098));
  jxor g2045(.dina(n1356), .dinb(n996), .dout(n2099));
  jnot g2046(.din(n2099), .dout(n2100));
  jand g2047(.dina(n2100), .dinb(n2098), .dout(n2101));
  jand g2048(.dina(n2101), .dinb(n2096), .dout(n2102));
  jand g2049(.dina(n2099), .dinb(n2098), .dout(n2103));
  jand g2050(.dina(n2103), .dinb(n2094), .dout(n2104));
  jxor g2051(.dina(n994), .dinb(n881), .dout(n2105));
  jnot g2052(.din(n2105), .dout(n2106));
  jand g2053(.dina(n2106), .dinb(n2097), .dout(n2107));
  jand g2054(.dina(n2107), .dinb(n1956), .dout(n2108));
  jor  g2055(.dina(n2108), .dinb(n2104), .dout(n2109));
  jor  g2056(.dina(n2109), .dinb(n2102), .dout(n2110));
  jnot g2057(.din(n2110), .dout(n2111));
  jand g2058(.dina(n2098), .dinb(n1956), .dout(n2112));
  jnot g2059(.din(n2112), .dout(n2113));
  jand g2060(.dina(n2113), .dinb(n1356), .dout(n2114));
  jand g2061(.dina(n2114), .dinb(n2111), .dout(n2115));
  jnot g2062(.din(n2094), .dout(n2116));
  jor  g2063(.dina(n2116), .dinb(n1956), .dout(n2117));
  jnot g2064(.din(n1996), .dout(n2118));
  jor  g2065(.dina(n1953), .dinb(n1664), .dout(n2119));
  jand g2066(.dina(n2119), .dinb(n2118), .dout(n2120));
  jxor g2067(.dina(n2091), .dinb(n2120), .dout(n2121));
  jand g2068(.dina(n2121), .dinb(n1994), .dout(n2122));
  jnot g2069(.din(n1960), .dout(n2123));
  jxor g2070(.dina(n2092), .dinb(n1993), .dout(n2124));
  jand g2071(.dina(n2124), .dinb(n2123), .dout(n2125));
  jor  g2072(.dina(n2125), .dinb(n2122), .dout(n2126));
  jand g2073(.dina(n852), .dinb(n600), .dout(n2127));
  jand g2074(.dina(n331), .dinb(n204), .dout(n2128));
  jand g2075(.dina(n2128), .dinb(n435), .dout(n2129));
  jand g2076(.dina(n2129), .dinb(n2127), .dout(n2130));
  jand g2077(.dina(n2130), .dinb(n1961), .dout(n2131));
  jand g2078(.dina(n395), .dinb(n265), .dout(n2132));
  jand g2079(.dina(n2132), .dinb(n825), .dout(n2133));
  jand g2080(.dina(n2133), .dinb(n491), .dout(n2134));
  jnot g2081(.din(n1180), .dout(n2135));
  jand g2082(.dina(n1345), .dinb(n2135), .dout(n2136));
  jand g2083(.dina(n2136), .dinb(n2134), .dout(n2137));
  jand g2084(.dina(n2137), .dinb(n2131), .dout(n2138));
  jand g2085(.dina(n366), .dinb(n218), .dout(n2139));
  jand g2086(.dina(n2139), .dinb(n411), .dout(n2140));
  jand g2087(.dina(n1035), .dinb(n248), .dout(n2141));
  jand g2088(.dina(n2141), .dinb(n527), .dout(n2142));
  jand g2089(.dina(n2142), .dinb(n586), .dout(n2143));
  jand g2090(.dina(n2143), .dinb(n510), .dout(n2144));
  jand g2091(.dina(n2144), .dinb(n2140), .dout(n2145));
  jand g2092(.dina(n2145), .dinb(n2138), .dout(n2146));
  jand g2093(.dina(n562), .dinb(n543), .dout(n2147));
  jand g2094(.dina(n2147), .dinb(n2146), .dout(n2148));
  jand g2095(.dina(n114), .dinb(n102), .dout(n2149));
  jand g2096(.dina(n347), .dinb(n213), .dout(n2150));
  jand g2097(.dina(n2150), .dinb(n2149), .dout(n2151));
  jand g2098(.dina(n439), .dinb(n339), .dout(n2152));
  jand g2099(.dina(n2152), .dinb(n430), .dout(n2153));
  jand g2100(.dina(n2153), .dinb(n2151), .dout(n2154));
  jand g2101(.dina(n570), .dinb(n897), .dout(n2155));
  jand g2102(.dina(n374), .dinb(n250), .dout(n2156));
  jand g2103(.dina(n2156), .dinb(n2155), .dout(n2157));
  jand g2104(.dina(n1459), .dinb(n1072), .dout(n2158));
  jand g2105(.dina(n2158), .dinb(n2157), .dout(n2159));
  jand g2106(.dina(n2159), .dinb(n2154), .dout(n2160));
  jand g2107(.dina(n1095), .dinb(n886), .dout(n2161));
  jand g2108(.dina(n269), .dinb(n195), .dout(n2162));
  jand g2109(.dina(n2162), .dinb(n2161), .dout(n2163));
  jand g2110(.dina(n2163), .dinb(n2160), .dout(n2164));
  jand g2111(.dina(n2164), .dinb(n180), .dout(n2165));
  jand g2112(.dina(n2165), .dinb(n2148), .dout(n2166));
  jand g2113(.dina(n2090), .dinb(n2026), .dout(n2167));
  jand g2114(.dina(n2091), .dinb(n2023), .dout(n2168));
  jor  g2115(.dina(n2168), .dinb(n2167), .dout(n2169));
  jand g2116(.dina(n2045), .dinb(n2029), .dout(n2170));
  jand g2117(.dina(n2089), .dinb(n2046), .dout(n2171));
  jor  g2118(.dina(n2171), .dinb(n2170), .dout(n2172));
  jand g2119(.dina(n2061), .dinb(n2049), .dout(n2173));
  jand g2120(.dina(n2088), .dinb(n2062), .dout(n2174));
  jor  g2121(.dina(n2174), .dinb(n2173), .dout(n2175));
  jand g2122(.dina(n1505), .dinb(n1168), .dout(n2176));
  jnot g2123(.din(n2176), .dout(n2177));
  jxor g2124(.dina(n1474), .dinb(n1272), .dout(n2178));
  jor  g2125(.dina(n2178), .dinb(n1490), .dout(n2179));
  jand g2126(.dina(n1493), .dinb(n1166), .dout(n2180));
  jnot g2127(.din(n2180), .dout(n2181));
  jand g2128(.dina(n2181), .dinb(n2179), .dout(n2182));
  jand g2129(.dina(n2182), .dinb(n2177), .dout(n2183));
  jand g2130(.dina(n2059), .dinb(n716), .dout(n2184));
  jand g2131(.dina(n2060), .dinb(n2058), .dout(n2185));
  jor  g2132(.dina(n2185), .dinb(n2184), .dout(n2186));
  jxor g2133(.dina(n2186), .dinb(n2183), .dout(n2187));
  jand g2134(.dina(n2086), .dinb(n2078), .dout(n2188));
  jand g2135(.dina(n2087), .dinb(n2070), .dout(n2189));
  jor  g2136(.dina(n2189), .dinb(n2188), .dout(n2190));
  jxor g2137(.dina(n2190), .dinb(n2187), .dout(n2191));
  jxor g2138(.dina(n2191), .dinb(n2175), .dout(n2192));
  jand g2139(.dina(n2040), .dinb(n2037), .dout(n2193));
  jand g2140(.dina(n2044), .dinb(n2041), .dout(n2194));
  jor  g2141(.dina(n2194), .dinb(n2193), .dout(n2195));
  jand g2142(.dina(n1551), .dinb(n881), .dout(n2196));
  jand g2143(.dina(n1549), .dinb(n880), .dout(n2197));
  jor  g2144(.dina(n2197), .dinb(n2196), .dout(n2198));
  jnot g2145(.din(n2198), .dout(n2199));
  jand g2146(.dina(n1558), .dinb(n1257), .dout(n2200));
  jand g2147(.dina(n1560), .dinb(n1259), .dout(n2201));
  jor  g2148(.dina(n2201), .dinb(n2200), .dout(n2202));
  jand g2149(.dina(n2202), .dinb(n2199), .dout(n2203));
  jand g2150(.dina(n1434), .dinb(n1255), .dout(n2204));
  jand g2151(.dina(n1622), .dinb(n1261), .dout(n2205));
  jor  g2152(.dina(n2205), .dinb(n2204), .dout(n2206));
  jnot g2153(.din(n2206), .dout(n2207));
  jand g2154(.dina(n1360), .dinb(n1270), .dout(n2208));
  jand g2155(.dina(n1485), .dinb(n1295), .dout(n2209));
  jor  g2156(.dina(n2209), .dinb(n2208), .dout(n2210));
  jand g2157(.dina(n2210), .dinb(n2207), .dout(n2211));
  jand g2158(.dina(n1416), .dinb(n996), .dout(n2212));
  jand g2159(.dina(n1418), .dinb(n994), .dout(n2213));
  jor  g2160(.dina(n2213), .dinb(n2212), .dout(n2214));
  jnot g2161(.din(n2214), .dout(n2215));
  jand g2162(.dina(n1356), .dinb(n1164), .dout(n2216));
  jand g2163(.dina(n1480), .dinb(n1170), .dout(n2217));
  jor  g2164(.dina(n2217), .dinb(n2216), .dout(n2218));
  jand g2165(.dina(n2218), .dinb(n2215), .dout(n2219));
  jxor g2166(.dina(n2219), .dinb(n2211), .dout(n2220));
  jxor g2167(.dina(n2220), .dinb(n2203), .dout(n2221));
  jand g2168(.dina(n2051), .dinb(n815), .dout(n2222));
  jand g2169(.dina(n1438), .dinb(n989), .dout(n2223));
  jor  g2170(.dina(n2223), .dinb(n1529), .dout(n2224));
  jor  g2171(.dina(n2224), .dinb(n2222), .dout(n2225));
  jnot g2172(.din(n2225), .dout(n2226));
  jand g2173(.dina(n1494), .dinb(n1154), .dout(n2227));
  jxor g2174(.dina(n2227), .dinb(n716), .dout(n2228));
  jxor g2175(.dina(n2228), .dinb(n2226), .dout(n2229));
  jxor g2176(.dina(n2229), .dinb(n2221), .dout(n2230));
  jxor g2177(.dina(n2230), .dinb(n2195), .dout(n2231));
  jxor g2178(.dina(n2231), .dinb(n2192), .dout(n2232));
  jxor g2179(.dina(n2232), .dinb(n2172), .dout(n2233));
  jxor g2180(.dina(n2233), .dinb(n2169), .dout(n2234));
  jxor g2181(.dina(n2234), .dinb(n2166), .dout(n2235));
  jxor g2182(.dina(n2235), .dinb(n2126), .dout(n2236));
  jxor g2183(.dina(n2236), .dinb(n2117), .dout(n2237));
  jnot g2184(.din(n2237), .dout(n2238));
  jand g2185(.dina(n2238), .dinb(n2101), .dout(n2239));
  jand g2186(.dina(n2107), .dinb(n2094), .dout(n2240));
  jand g2187(.dina(n2236), .dinb(n2103), .dout(n2241));
  jor  g2188(.dina(n2241), .dinb(n2240), .dout(n2242));
  jand g2189(.dina(n2105), .dinb(n2097), .dout(n2243));
  jand g2190(.dina(n2243), .dinb(n2100), .dout(n2244));
  jand g2191(.dina(n2244), .dinb(n1956), .dout(n2245));
  jor  g2192(.dina(n2245), .dinb(n2242), .dout(n2246));
  jor  g2193(.dina(n2246), .dinb(n2239), .dout(n2247));
  jnot g2194(.din(n2247), .dout(n2248));
  jand g2195(.dina(n2248), .dinb(n2115), .dout(n2249));
  jand g2196(.dina(n2249), .dinb(n1959), .dout(n2250));
  jxor g2197(.dina(n2249), .dinb(n1959), .dout(n2251));
  jnot g2198(.din(n2101), .dout(n2252));
  jor  g2199(.dina(n2092), .dinb(n1993), .dout(n2253));
  jor  g2200(.dina(n2093), .dinb(n1960), .dout(n2254));
  jand g2201(.dina(n2254), .dinb(n2253), .dout(n2255));
  jxor g2202(.dina(n2235), .dinb(n2255), .dout(n2256));
  jand g2203(.dina(n2256), .dinb(n1955), .dout(n2257));
  jor  g2204(.dina(n2257), .dinb(n2116), .dout(n2258));
  jor  g2205(.dina(n2234), .dinb(n2166), .dout(n2259));
  jnot g2206(.din(n2166), .dout(n2260));
  jxor g2207(.dina(n2234), .dinb(n2260), .dout(n2261));
  jor  g2208(.dina(n2261), .dinb(n2255), .dout(n2262));
  jand g2209(.dina(n2262), .dinb(n2259), .dout(n2263));
  jand g2210(.dina(n1127), .dinb(n129), .dout(n2264));
  jand g2211(.dina(n2264), .dinb(n445), .dout(n2265));
  jand g2212(.dina(n2265), .dinb(n222), .dout(n2266));
  jand g2213(.dina(n2266), .dinb(n2154), .dout(n2267));
  jand g2214(.dina(n2267), .dinb(n1016), .dout(n2268));
  jand g2215(.dina(n434), .dinb(n221), .dout(n2269));
  jand g2216(.dina(n2269), .dinb(n244), .dout(n2270));
  jand g2217(.dina(n337), .dinb(n232), .dout(n2271));
  jand g2218(.dina(n717), .dinb(n197), .dout(n2272));
  jand g2219(.dina(n2272), .dinb(n2271), .dout(n2273));
  jand g2220(.dina(n2273), .dinb(n329), .dout(n2274));
  jand g2221(.dina(n2274), .dinb(n394), .dout(n2275));
  jand g2222(.dina(n2275), .dinb(n2270), .dout(n2276));
  jand g2223(.dina(n2276), .dinb(n2268), .dout(n2277));
  jand g2224(.dina(n2232), .dinb(n2172), .dout(n2278));
  jand g2225(.dina(n2233), .dinb(n2169), .dout(n2279));
  jor  g2226(.dina(n2279), .dinb(n2278), .dout(n2280));
  jand g2227(.dina(n2191), .dinb(n2175), .dout(n2281));
  jand g2228(.dina(n2231), .dinb(n2192), .dout(n2282));
  jor  g2229(.dina(n2282), .dinb(n2281), .dout(n2283));
  jand g2230(.dina(n2229), .dinb(n2221), .dout(n2284));
  jand g2231(.dina(n2230), .dinb(n2195), .dout(n2285));
  jor  g2232(.dina(n2285), .dinb(n2284), .dout(n2286));
  jand g2233(.dina(n2227), .dinb(n716), .dout(n2287));
  jand g2234(.dina(n2228), .dinb(n2226), .dout(n2288));
  jor  g2235(.dina(n2288), .dinb(n2287), .dout(n2289));
  jand g2236(.dina(n1485), .dinb(n1576), .dout(n2290));
  jand g2237(.dina(n1360), .dinb(n1163), .dout(n2291));
  jor  g2238(.dina(n2291), .dinb(n2290), .dout(n2292));
  jnot g2239(.din(n2292), .dout(n2293));
  jand g2240(.dina(n1356), .dinb(n1160), .dout(n2294));
  jand g2241(.dina(n1480), .dinb(n1152), .dout(n2295));
  jor  g2242(.dina(n2295), .dinb(n2294), .dout(n2296));
  jand g2243(.dina(n2296), .dinb(n2293), .dout(n2297));
  jand g2244(.dina(n1532), .dinb(n716), .dout(n2298));
  jnot g2245(.din(n2298), .dout(n2299));
  jand g2246(.dina(n930), .dinb(n607), .dout(n2300));
  jnot g2247(.din(n2300), .dout(n2301));
  jand g2248(.dina(n1494), .dinb(n1166), .dout(n2302));
  jand g2249(.dina(n2301), .dinb(n2302), .dout(n2303));
  jand g2250(.dina(n2303), .dinb(n2299), .dout(n2304));
  jnot g2251(.din(n2304), .dout(n2305));
  jand g2252(.dina(n2305), .dinb(n2301), .dout(n2306));
  jand g2253(.dina(n2306), .dinb(n2299), .dout(n2307));
  jand g2254(.dina(n2305), .dinb(n2302), .dout(n2308));
  jor  g2255(.dina(n2308), .dinb(n2307), .dout(n2309));
  jxor g2256(.dina(n2309), .dinb(n2297), .dout(n2310));
  jxor g2257(.dina(n2310), .dinb(n2289), .dout(n2311));
  jxor g2258(.dina(n2311), .dinb(n2286), .dout(n2312));
  jand g2259(.dina(n2186), .dinb(n2183), .dout(n2313));
  jand g2260(.dina(n2190), .dinb(n2187), .dout(n2314));
  jor  g2261(.dina(n2314), .dinb(n2313), .dout(n2315));
  jand g2262(.dina(n2219), .dinb(n2211), .dout(n2316));
  jand g2263(.dina(n2220), .dinb(n2203), .dout(n2317));
  jor  g2264(.dina(n2317), .dinb(n2316), .dout(n2318));
  jand g2265(.dina(n1622), .dinb(n1649), .dout(n2319));
  jand g2266(.dina(n1434), .dinb(n1651), .dout(n2320));
  jor  g2267(.dina(n2320), .dinb(n2319), .dout(n2321));
  jnot g2268(.din(n2321), .dout(n2322));
  jand g2269(.dina(n2051), .dinb(n1656), .dout(n2323));
  jand g2270(.dina(n1438), .dinb(n1254), .dout(n2324));
  jor  g2271(.dina(n2324), .dinb(n2323), .dout(n2325));
  jand g2272(.dina(n2325), .dinb(n2322), .dout(n2326));
  jand g2273(.dina(n1551), .dinb(n996), .dout(n2327));
  jand g2274(.dina(n1549), .dinb(n994), .dout(n2328));
  jor  g2275(.dina(n2328), .dinb(n2327), .dout(n2329));
  jnot g2276(.din(n2329), .dout(n2330));
  jand g2277(.dina(n1558), .dinb(n880), .dout(n2331));
  jand g2278(.dina(n1560), .dinb(n881), .dout(n2332));
  jor  g2279(.dina(n2332), .dinb(n2331), .dout(n2333));
  jand g2280(.dina(n2333), .dinb(n2330), .dout(n2334));
  jand g2281(.dina(n1505), .dinb(n1272), .dout(n2335));
  jnot g2282(.din(n2335), .dout(n2336));
  jxor g2283(.dina(n1474), .dinb(n1259), .dout(n2337));
  jor  g2284(.dina(n2337), .dinb(n1490), .dout(n2338));
  jand g2285(.dina(n1493), .dinb(n1266), .dout(n2339));
  jnot g2286(.din(n2339), .dout(n2340));
  jand g2287(.dina(n2340), .dinb(n2338), .dout(n2341));
  jand g2288(.dina(n2341), .dinb(n2336), .dout(n2342));
  jxor g2289(.dina(n2342), .dinb(n2334), .dout(n2343));
  jxor g2290(.dina(n2343), .dinb(n2326), .dout(n2344));
  jxor g2291(.dina(n2344), .dinb(n2318), .dout(n2345));
  jxor g2292(.dina(n2345), .dinb(n2315), .dout(n2346));
  jxor g2293(.dina(n2346), .dinb(n2312), .dout(n2347));
  jxor g2294(.dina(n2347), .dinb(n2283), .dout(n2348));
  jxor g2295(.dina(n2348), .dinb(n2280), .dout(n2349));
  jxor g2296(.dina(n2349), .dinb(n2277), .dout(n2350));
  jxor g2297(.dina(n2350), .dinb(n2263), .dout(n2351));
  jxor g2298(.dina(n2351), .dinb(n2256), .dout(n2352));
  jxor g2299(.dina(n2352), .dinb(n2258), .dout(n2353));
  jor  g2300(.dina(n2353), .dinb(n2252), .dout(n2354));
  jnot g2301(.din(n2103), .dout(n2355));
  jor  g2302(.dina(n2351), .dinb(n2355), .dout(n2356));
  jnot g2303(.din(n2244), .dout(n2357));
  jor  g2304(.dina(n2357), .dinb(n2116), .dout(n2358));
  jnot g2305(.din(n2107), .dout(n2359));
  jor  g2306(.dina(n2256), .dinb(n2359), .dout(n2360));
  jand g2307(.dina(n2360), .dinb(n2358), .dout(n2361));
  jand g2308(.dina(n2361), .dinb(n2356), .dout(n2362));
  jand g2309(.dina(n2362), .dinb(n2354), .dout(n2363));
  jxor g2310(.dina(n2363), .dinb(n1480), .dout(n2364));
  jand g2311(.dina(n2364), .dinb(n2251), .dout(n2365));
  jor  g2312(.dina(n2365), .dinb(n2250), .dout(n2366));
  jor  g2313(.dina(n2351), .dinb(n2256), .dout(n2367));
  jxor g2314(.dina(n2351), .dinb(n2236), .dout(n2368));
  jor  g2315(.dina(n2368), .dinb(n2258), .dout(n2369));
  jand g2316(.dina(n2369), .dinb(n2367), .dout(n2370));
  jor  g2317(.dina(n2349), .dinb(n2277), .dout(n2371));
  jnot g2318(.din(n2277), .dout(n2372));
  jxor g2319(.dina(n2349), .dinb(n2372), .dout(n2373));
  jor  g2320(.dina(n2373), .dinb(n2263), .dout(n2374));
  jand g2321(.dina(n2374), .dinb(n2371), .dout(n2375));
  jand g2322(.dina(n439), .dinb(n427), .dout(n2376));
  jand g2323(.dina(n2376), .dinb(n1096), .dout(n2377));
  jand g2324(.dina(n2377), .dinb(n283), .dout(n2378));
  jand g2325(.dina(n2378), .dinb(n866), .dout(n2379));
  jand g2326(.dina(n160), .dinb(n124), .dout(n2380));
  jand g2327(.dina(n2380), .dinb(n1345), .dout(n2381));
  jand g2328(.dina(n2381), .dinb(n218), .dout(n2382));
  jand g2329(.dina(n2382), .dinb(n1135), .dout(n2383));
  jand g2330(.dina(n2383), .dinb(n2379), .dout(n2384));
  jand g2331(.dina(n2384), .dinb(n137), .dout(n2385));
  jand g2332(.dina(n2385), .dinb(n404), .dout(n2386));
  jand g2333(.dina(n340), .dinb(n457), .dout(n2387));
  jand g2334(.dina(n2387), .dinb(n411), .dout(n2388));
  jand g2335(.dina(n467), .dinb(n235), .dout(n2389));
  jand g2336(.dina(n2389), .dinb(n309), .dout(n2390));
  jand g2337(.dina(n2390), .dinb(n294), .dout(n2391));
  jand g2338(.dina(n2391), .dinb(n2388), .dout(n2392));
  jand g2339(.dina(n337), .dinb(n102), .dout(n2393));
  jand g2340(.dina(n2393), .dinb(n327), .dout(n2394));
  jand g2341(.dina(n300), .dinb(n248), .dout(n2395));
  jand g2342(.dina(n2395), .dinb(n409), .dout(n2396));
  jand g2343(.dina(n2396), .dinb(n2394), .dout(n2397));
  jand g2344(.dina(n587), .dinb(n305), .dout(n2398));
  jand g2345(.dina(n2398), .dinb(n1057), .dout(n2399));
  jand g2346(.dina(n2399), .dinb(n315), .dout(n2400));
  jand g2347(.dina(n2400), .dinb(n530), .dout(n2401));
  jand g2348(.dina(n2401), .dinb(n2397), .dout(n2402));
  jand g2349(.dina(n2402), .dinb(n370), .dout(n2403));
  jand g2350(.dina(n534), .dinb(n245), .dout(n2404));
  jand g2351(.dina(n600), .dinb(n384), .dout(n2405));
  jand g2352(.dina(n2405), .dinb(n2404), .dout(n2406));
  jand g2353(.dina(n361), .dinb(n213), .dout(n2407));
  jand g2354(.dina(n2407), .dinb(n170), .dout(n2408));
  jand g2355(.dina(n2408), .dinb(n2406), .dout(n2409));
  jand g2356(.dina(n2409), .dinb(n2403), .dout(n2410));
  jand g2357(.dina(n2410), .dinb(n2392), .dout(n2411));
  jand g2358(.dina(n2411), .dinb(n2386), .dout(n2412));
  jand g2359(.dina(n2347), .dinb(n2283), .dout(n2413));
  jand g2360(.dina(n2348), .dinb(n2280), .dout(n2414));
  jor  g2361(.dina(n2414), .dinb(n2413), .dout(n2415));
  jand g2362(.dina(n2311), .dinb(n2286), .dout(n2416));
  jand g2363(.dina(n2346), .dinb(n2312), .dout(n2417));
  jor  g2364(.dina(n2417), .dinb(n2416), .dout(n2418));
  jand g2365(.dina(n2309), .dinb(n2297), .dout(n2419));
  jand g2366(.dina(n2310), .dinb(n2289), .dout(n2420));
  jor  g2367(.dina(n2420), .dinb(n2419), .dout(n2421));
  jand g2368(.dina(n2344), .dinb(n2318), .dout(n2422));
  jand g2369(.dina(n2345), .dinb(n2315), .dout(n2423));
  jor  g2370(.dina(n2423), .dinb(n2422), .dout(n2424));
  jxor g2371(.dina(n2424), .dinb(n2421), .dout(n2425));
  jnot g2372(.din(n2306), .dout(n2426));
  jand g2373(.dina(n1551), .dinb(n1480), .dout(n2427));
  jand g2374(.dina(n1549), .dinb(n1356), .dout(n2428));
  jor  g2375(.dina(n2428), .dinb(n2427), .dout(n2429));
  jnot g2376(.din(n2429), .dout(n2430));
  jand g2377(.dina(n1558), .dinb(n994), .dout(n2431));
  jand g2378(.dina(n1560), .dinb(n996), .dout(n2432));
  jor  g2379(.dina(n2432), .dinb(n2431), .dout(n2433));
  jand g2380(.dina(n2433), .dinb(n2430), .dout(n2434));
  jand g2381(.dina(n1493), .dinb(n1257), .dout(n2435));
  jnot g2382(.din(n2435), .dout(n2436));
  jxor g2383(.dina(n1474), .dinb(n881), .dout(n2437));
  jor  g2384(.dina(n2437), .dinb(n1490), .dout(n2438));
  jand g2385(.dina(n1505), .dinb(n1259), .dout(n2439));
  jnot g2386(.din(n2439), .dout(n2440));
  jand g2387(.dina(n2440), .dinb(n2438), .dout(n2441));
  jand g2388(.dina(n2441), .dinb(n2436), .dout(n2442));
  jxor g2389(.dina(n2442), .dinb(n2434), .dout(n2443));
  jxor g2390(.dina(n2443), .dinb(n2426), .dout(n2444));
  jand g2391(.dina(n2342), .dinb(n2334), .dout(n2445));
  jand g2392(.dina(n2343), .dinb(n2326), .dout(n2446));
  jor  g2393(.dina(n2446), .dinb(n2445), .dout(n2447));
  jand g2394(.dina(n1485), .dinb(n1416), .dout(n2448));
  jand g2395(.dina(n1360), .dinb(n1418), .dout(n2449));
  jor  g2396(.dina(n2449), .dinb(n2448), .dout(n2450));
  jnot g2397(.din(n2450), .dout(n2451));
  jand g2398(.dina(n1434), .dinb(n1164), .dout(n2452));
  jand g2399(.dina(n1622), .dinb(n1170), .dout(n2453));
  jor  g2400(.dina(n2453), .dinb(n2452), .dout(n2454));
  jand g2401(.dina(n2454), .dinb(n2451), .dout(n2455));
  jand g2402(.dina(n1494), .dinb(n1266), .dout(n2456));
  jnot g2403(.din(n2456), .dout(n2457));
  jand g2404(.dina(n1438), .dinb(n1651), .dout(n2458));
  jnot g2405(.din(n2458), .dout(n2459));
  jand g2406(.dina(n1438), .dinb(n1812), .dout(n2460));
  jor  g2407(.dina(n2460), .dinb(n1294), .dout(n2461));
  jand g2408(.dina(n2461), .dinb(n2459), .dout(n2462));
  jxor g2409(.dina(n2462), .dinb(n2457), .dout(n2463));
  jxor g2410(.dina(n2463), .dinb(n2455), .dout(n2464));
  jxor g2411(.dina(n2464), .dinb(n2447), .dout(n2465));
  jxor g2412(.dina(n2465), .dinb(n2444), .dout(n2466));
  jxor g2413(.dina(n2466), .dinb(n2425), .dout(n2467));
  jxor g2414(.dina(n2467), .dinb(n2418), .dout(n2468));
  jxor g2415(.dina(n2468), .dinb(n2415), .dout(n2469));
  jxor g2416(.dina(n2469), .dinb(n2412), .dout(n2470));
  jxor g2417(.dina(n2470), .dinb(n2375), .dout(n2471));
  jxor g2418(.dina(n2471), .dinb(n2351), .dout(n2472));
  jxor g2419(.dina(n2472), .dinb(n2370), .dout(n2473));
  jor  g2420(.dina(n2473), .dinb(n2252), .dout(n2474));
  jor  g2421(.dina(n2351), .dinb(n2359), .dout(n2475));
  jor  g2422(.dina(n2471), .dinb(n2355), .dout(n2476));
  jand g2423(.dina(n2476), .dinb(n2475), .dout(n2477));
  jor  g2424(.dina(n2357), .dinb(n2256), .dout(n2478));
  jand g2425(.dina(n2478), .dinb(n2477), .dout(n2479));
  jand g2426(.dina(n2479), .dinb(n2474), .dout(n2480));
  jxor g2427(.dina(n2480), .dinb(n1356), .dout(n2481));
  jnot g2428(.din(n2481), .dout(n2482));
  jxor g2429(.dina(n1438), .dinb(n1434), .dout(n2483));
  jand g2430(.dina(n2483), .dinb(n1958), .dout(n2484));
  jand g2431(.dina(n2484), .dinb(n2096), .dout(n2485));
  jxor g2432(.dina(n1434), .dinb(n1485), .dout(n2486));
  jnot g2433(.din(n2486), .dout(n2487));
  jand g2434(.dina(n2487), .dinb(n1957), .dout(n2488));
  jand g2435(.dina(n2488), .dinb(n1956), .dout(n2489));
  jnot g2436(.din(n2483), .dout(n2490));
  jand g2437(.dina(n2490), .dinb(n1958), .dout(n2491));
  jand g2438(.dina(n2491), .dinb(n2094), .dout(n2492));
  jor  g2439(.dina(n2492), .dinb(n2489), .dout(n2493));
  jor  g2440(.dina(n2493), .dinb(n2485), .dout(n2494));
  jand g2441(.dina(n1956), .dinb(n1438), .dout(n2495));
  jand g2442(.dina(n2495), .dinb(n1958), .dout(n2496));
  jxor g2443(.dina(n2496), .dinb(n2494), .dout(n2497));
  jxor g2444(.dina(n2497), .dinb(n2482), .dout(n2498));
  jxor g2445(.dina(n2498), .dinb(n2366), .dout(n2499));
  jnot g2446(.din(n2499), .dout(n2500));
  jxor g2447(.dina(n1166), .dinb(n1156), .dout(n2501));
  jnot g2448(.din(n2501), .dout(n2502));
  jxor g2449(.dina(n1272), .dinb(n1257), .dout(n2503));
  jnot g2450(.din(n2503), .dout(n2504));
  jand g2451(.dina(n2504), .dinb(n2502), .dout(n2505));
  jnot g2452(.din(n2505), .dout(n2506));
  jand g2453(.dina(n2134), .dinb(n583), .dout(n2507));
  jand g2454(.dina(n1366), .dinb(n238), .dout(n2508));
  jand g2455(.dina(n2508), .dinb(n2507), .dout(n2509));
  jand g2456(.dina(n1002), .dinb(n332), .dout(n2510));
  jand g2457(.dina(n2510), .dinb(n1987), .dout(n2511));
  jand g2458(.dina(n2511), .dinb(n2509), .dout(n2512));
  jand g2459(.dina(n162), .dinb(n124), .dout(n2513));
  jand g2460(.dina(n2513), .dinb(n1064), .dout(n2514));
  jand g2461(.dina(n847), .dinb(n539), .dout(n2515));
  jand g2462(.dina(n2515), .dinb(n2514), .dout(n2516));
  jand g2463(.dina(n2516), .dinb(n531), .dout(n2517));
  jand g2464(.dina(n2517), .dinb(n1249), .dout(n2518));
  jand g2465(.dina(n2518), .dinb(n2512), .dout(n2519));
  jnot g2466(.din(n2519), .dout(n2520));
  jand g2467(.dina(n2467), .dinb(n2418), .dout(n2521));
  jnot g2468(.din(n2521), .dout(n2522));
  jnot g2469(.din(n2413), .dout(n2523));
  jnot g2470(.din(n2278), .dout(n2524));
  jnot g2471(.din(n2167), .dout(n2525));
  jnot g2472(.din(n2091), .dout(n2526));
  jor  g2473(.dina(n2526), .dinb(n2120), .dout(n2527));
  jand g2474(.dina(n2527), .dinb(n2525), .dout(n2528));
  jnot g2475(.din(n2233), .dout(n2529));
  jor  g2476(.dina(n2529), .dinb(n2528), .dout(n2530));
  jand g2477(.dina(n2530), .dinb(n2524), .dout(n2531));
  jnot g2478(.din(n2348), .dout(n2532));
  jor  g2479(.dina(n2532), .dinb(n2531), .dout(n2533));
  jand g2480(.dina(n2533), .dinb(n2523), .dout(n2534));
  jnot g2481(.din(n2468), .dout(n2535));
  jor  g2482(.dina(n2535), .dinb(n2534), .dout(n2536));
  jand g2483(.dina(n2536), .dinb(n2522), .dout(n2537));
  jand g2484(.dina(n2424), .dinb(n2421), .dout(n2538));
  jand g2485(.dina(n2466), .dinb(n2425), .dout(n2539));
  jor  g2486(.dina(n2539), .dinb(n2538), .dout(n2540));
  jand g2487(.dina(n2464), .dinb(n2447), .dout(n2541));
  jand g2488(.dina(n2465), .dinb(n2444), .dout(n2542));
  jor  g2489(.dina(n2542), .dinb(n2541), .dout(n2543));
  jand g2490(.dina(n1505), .dinb(n881), .dout(n2544));
  jnot g2491(.din(n2544), .dout(n2545));
  jxor g2492(.dina(n1474), .dinb(n996), .dout(n2546));
  jor  g2493(.dina(n2546), .dinb(n1490), .dout(n2547));
  jand g2494(.dina(n1493), .dinb(n880), .dout(n2548));
  jnot g2495(.din(n2548), .dout(n2549));
  jand g2496(.dina(n2549), .dinb(n2547), .dout(n2550));
  jand g2497(.dina(n2550), .dinb(n2545), .dout(n2551));
  jand g2498(.dina(n1434), .dinb(n1418), .dout(n2552));
  jand g2499(.dina(n1622), .dinb(n1416), .dout(n2553));
  jor  g2500(.dina(n2553), .dinb(n2552), .dout(n2554));
  jnot g2501(.din(n2554), .dout(n2555));
  jand g2502(.dina(n2051), .dinb(n1170), .dout(n2556));
  jand g2503(.dina(n1438), .dinb(n1164), .dout(n2557));
  jor  g2504(.dina(n2557), .dinb(n2556), .dout(n2558));
  jand g2505(.dina(n2558), .dinb(n2555), .dout(n2559));
  jand g2506(.dina(n1551), .dinb(n1485), .dout(n2560));
  jand g2507(.dina(n1549), .dinb(n1360), .dout(n2561));
  jor  g2508(.dina(n2561), .dinb(n2560), .dout(n2562));
  jnot g2509(.din(n2562), .dout(n2563));
  jand g2510(.dina(n1558), .dinb(n1356), .dout(n2564));
  jand g2511(.dina(n1560), .dinb(n1480), .dout(n2565));
  jor  g2512(.dina(n2565), .dinb(n2564), .dout(n2566));
  jand g2513(.dina(n2566), .dinb(n2563), .dout(n2567));
  jxor g2514(.dina(n2567), .dinb(n2559), .dout(n2568));
  jxor g2515(.dina(n2568), .dinb(n2551), .dout(n2569));
  jxor g2516(.dina(n2569), .dinb(n2543), .dout(n2570));
  jand g2517(.dina(n2442), .dinb(n2434), .dout(n2571));
  jand g2518(.dina(n2443), .dinb(n2426), .dout(n2572));
  jor  g2519(.dina(n2572), .dinb(n2571), .dout(n2573));
  jand g2520(.dina(n2462), .dinb(n2457), .dout(n2574));
  jand g2521(.dina(n2463), .dinb(n2455), .dout(n2575));
  jor  g2522(.dina(n2575), .dinb(n2574), .dout(n2576));
  jxor g2523(.dina(n2576), .dinb(n2573), .dout(n2577));
  jand g2524(.dina(n1494), .dinb(n1257), .dout(n2578));
  jxor g2525(.dina(n2456), .dinb(n1232), .dout(n2579));
  jxor g2526(.dina(n2579), .dinb(n2578), .dout(n2580));
  jxor g2527(.dina(n2580), .dinb(n2577), .dout(n2581));
  jxor g2528(.dina(n2581), .dinb(n2570), .dout(n2582));
  jxor g2529(.dina(n2582), .dinb(n2540), .dout(n2583));
  jxor g2530(.dina(n2583), .dinb(n2537), .dout(n2584));
  jand g2531(.dina(n2584), .dinb(n2520), .dout(n2585));
  jnot g2532(.din(n2412), .dout(n2586));
  jxor g2533(.dina(n2468), .dinb(n2534), .dout(n2587));
  jand g2534(.dina(n2587), .dinb(n2586), .dout(n2588));
  jxor g2535(.dina(n2348), .dinb(n2531), .dout(n2589));
  jand g2536(.dina(n2589), .dinb(n2372), .dout(n2590));
  jxor g2537(.dina(n2233), .dinb(n2528), .dout(n2591));
  jand g2538(.dina(n2591), .dinb(n2260), .dout(n2592));
  jand g2539(.dina(n2235), .dinb(n2126), .dout(n2593));
  jor  g2540(.dina(n2593), .dinb(n2592), .dout(n2594));
  jand g2541(.dina(n2350), .dinb(n2594), .dout(n2595));
  jor  g2542(.dina(n2595), .dinb(n2590), .dout(n2596));
  jand g2543(.dina(n2470), .dinb(n2596), .dout(n2597));
  jor  g2544(.dina(n2597), .dinb(n2588), .dout(n2598));
  jand g2545(.dina(n2468), .dinb(n2415), .dout(n2599));
  jor  g2546(.dina(n2599), .dinb(n2521), .dout(n2600));
  jxor g2547(.dina(n2583), .dinb(n2600), .dout(n2601));
  jxor g2548(.dina(n2601), .dinb(n2519), .dout(n2602));
  jand g2549(.dina(n2602), .dinb(n2598), .dout(n2603));
  jor  g2550(.dina(n2603), .dinb(n2585), .dout(n2604));
  jand g2551(.dina(n389), .dinb(n120), .dout(n2605));
  jand g2552(.dina(n2605), .dinb(n551), .dout(n2606));
  jand g2553(.dina(n489), .dinb(n215), .dout(n2607));
  jand g2554(.dina(n244), .dinb(n162), .dout(n2608));
  jand g2555(.dina(n275), .dinb(n255), .dout(n2609));
  jand g2556(.dina(n2609), .dinb(n2608), .dout(n2610));
  jand g2557(.dina(n321), .dinb(n288), .dout(n2611));
  jand g2558(.dina(n2611), .dinb(n2610), .dout(n2612));
  jand g2559(.dina(n2612), .dinb(n2607), .dout(n2613));
  jand g2560(.dina(n448), .dinb(n238), .dout(n2614));
  jand g2561(.dina(n221), .dinb(n124), .dout(n2615));
  jand g2562(.dina(n2615), .dinb(n261), .dout(n2616));
  jand g2563(.dina(n2616), .dinb(n2614), .dout(n2617));
  jand g2564(.dina(n383), .dinb(n300), .dout(n2618));
  jand g2565(.dina(n2618), .dinb(n377), .dout(n2619));
  jand g2566(.dina(n2619), .dinb(n339), .dout(n2620));
  jand g2567(.dina(n2620), .dinb(n2617), .dout(n2621));
  jand g2568(.dina(n2621), .dinb(n2613), .dout(n2622));
  jand g2569(.dina(n427), .dinb(n206), .dout(n2623));
  jand g2570(.dina(n467), .dinb(n460), .dout(n2624));
  jand g2571(.dina(n2624), .dinb(n2623), .dout(n2625));
  jand g2572(.dina(n2625), .dinb(n853), .dout(n2626));
  jand g2573(.dina(n1322), .dinb(n170), .dout(n2627));
  jand g2574(.dina(n1035), .dinb(n1005), .dout(n2628));
  jand g2575(.dina(n2628), .dinb(n2627), .dout(n2629));
  jand g2576(.dina(n2629), .dinb(n2626), .dout(n2630));
  jand g2577(.dina(n2630), .dinb(n560), .dout(n2631));
  jand g2578(.dina(n2631), .dinb(n455), .dout(n2632));
  jand g2579(.dina(n1095), .dinb(n232), .dout(n2633));
  jand g2580(.dina(n2633), .dinb(n2632), .dout(n2634));
  jand g2581(.dina(n2634), .dinb(n2622), .dout(n2635));
  jand g2582(.dina(n2635), .dinb(n2606), .dout(n2636));
  jand g2583(.dina(n2582), .dinb(n2540), .dout(n2637));
  jand g2584(.dina(n2583), .dinb(n2600), .dout(n2638));
  jor  g2585(.dina(n2638), .dinb(n2637), .dout(n2639));
  jand g2586(.dina(n2569), .dinb(n2543), .dout(n2640));
  jand g2587(.dina(n2581), .dinb(n2570), .dout(n2641));
  jor  g2588(.dina(n2641), .dinb(n2640), .dout(n2642));
  jand g2589(.dina(n2576), .dinb(n2573), .dout(n2643));
  jand g2590(.dina(n2580), .dinb(n2577), .dout(n2644));
  jor  g2591(.dina(n2644), .dinb(n2643), .dout(n2645));
  jand g2592(.dina(n1551), .dinb(n1622), .dout(n2646));
  jand g2593(.dina(n1549), .dinb(n1434), .dout(n2647));
  jor  g2594(.dina(n2647), .dinb(n2646), .dout(n2648));
  jnot g2595(.din(n2648), .dout(n2649));
  jand g2596(.dina(n1558), .dinb(n1360), .dout(n2650));
  jand g2597(.dina(n1560), .dinb(n1485), .dout(n2651));
  jor  g2598(.dina(n2651), .dinb(n2650), .dout(n2652));
  jand g2599(.dina(n2652), .dinb(n2649), .dout(n2653));
  jand g2600(.dina(n1494), .dinb(n880), .dout(n2654));
  jnot g2601(.din(n1151), .dout(n2655));
  jand g2602(.dina(n2051), .dinb(n2655), .dout(n2656));
  jand g2603(.dina(n1438), .dinb(n1418), .dout(n2657));
  jor  g2604(.dina(n2657), .dinb(n1576), .dout(n2658));
  jor  g2605(.dina(n2658), .dinb(n2656), .dout(n2659));
  jxor g2606(.dina(n2659), .dinb(n2654), .dout(n2660));
  jxor g2607(.dina(n2660), .dinb(n2653), .dout(n2661));
  jxor g2608(.dina(n2661), .dinb(n2645), .dout(n2662));
  jand g2609(.dina(n2567), .dinb(n2559), .dout(n2663));
  jand g2610(.dina(n2568), .dinb(n2551), .dout(n2664));
  jor  g2611(.dina(n2664), .dinb(n2663), .dout(n2665));
  jand g2612(.dina(n1505), .dinb(n996), .dout(n2666));
  jnot g2613(.din(n2666), .dout(n2667));
  jxor g2614(.dina(n1474), .dinb(n1480), .dout(n2668));
  jor  g2615(.dina(n2668), .dinb(n1490), .dout(n2669));
  jand g2616(.dina(n1493), .dinb(n994), .dout(n2670));
  jnot g2617(.din(n2670), .dout(n2671));
  jand g2618(.dina(n2671), .dinb(n2669), .dout(n2672));
  jand g2619(.dina(n2672), .dinb(n2667), .dout(n2673));
  jand g2620(.dina(n2456), .dinb(n1232), .dout(n2674));
  jand g2621(.dina(n2579), .dinb(n2578), .dout(n2675));
  jor  g2622(.dina(n2675), .dinb(n2674), .dout(n2676));
  jxor g2623(.dina(n2676), .dinb(n2673), .dout(n2677));
  jxor g2624(.dina(n2677), .dinb(n2665), .dout(n2678));
  jxor g2625(.dina(n2678), .dinb(n2662), .dout(n2679));
  jxor g2626(.dina(n2679), .dinb(n2642), .dout(n2680));
  jxor g2627(.dina(n2680), .dinb(n2639), .dout(n2681));
  jxor g2628(.dina(n2681), .dinb(n2636), .dout(n2682));
  jxor g2629(.dina(n2682), .dinb(n2604), .dout(n2683));
  jxor g2630(.dina(n2602), .dinb(n2598), .dout(n2684));
  jand g2631(.dina(n2684), .dinb(n2683), .dout(n2685));
  jnot g2632(.din(n2685), .dout(n2686));
  jxor g2633(.dina(n2470), .dinb(n2596), .dout(n2687));
  jand g2634(.dina(n2684), .dinb(n2687), .dout(n2688));
  jnot g2635(.din(n2688), .dout(n2689));
  jxor g2636(.dina(n2350), .dinb(n2594), .dout(n2690));
  jand g2637(.dina(n2687), .dinb(n2690), .dout(n2691));
  jnot g2638(.din(n2691), .dout(n2692));
  jxor g2639(.dina(n2687), .dinb(n2351), .dout(n2693));
  jor  g2640(.dina(n2693), .dinb(n2370), .dout(n2694));
  jand g2641(.dina(n2694), .dinb(n2692), .dout(n2695));
  jxor g2642(.dina(n2684), .dinb(n2471), .dout(n2696));
  jor  g2643(.dina(n2696), .dinb(n2695), .dout(n2697));
  jand g2644(.dina(n2697), .dinb(n2689), .dout(n2698));
  jor  g2645(.dina(n2601), .dinb(n2519), .dout(n2699));
  jor  g2646(.dina(n2469), .dinb(n2412), .dout(n2700));
  jxor g2647(.dina(n2469), .dinb(n2586), .dout(n2701));
  jor  g2648(.dina(n2701), .dinb(n2375), .dout(n2702));
  jand g2649(.dina(n2702), .dinb(n2700), .dout(n2703));
  jxor g2650(.dina(n2601), .dinb(n2520), .dout(n2704));
  jor  g2651(.dina(n2704), .dinb(n2703), .dout(n2705));
  jand g2652(.dina(n2705), .dinb(n2699), .dout(n2706));
  jxor g2653(.dina(n2682), .dinb(n2706), .dout(n2707));
  jxor g2654(.dina(n2684), .dinb(n2707), .dout(n2708));
  jor  g2655(.dina(n2708), .dinb(n2698), .dout(n2709));
  jand g2656(.dina(n2709), .dinb(n2686), .dout(n2710));
  jor  g2657(.dina(n2681), .dinb(n2636), .dout(n2711));
  jnot g2658(.din(n2636), .dout(n2712));
  jxor g2659(.dina(n2681), .dinb(n2712), .dout(n2713));
  jor  g2660(.dina(n2713), .dinb(n2706), .dout(n2714));
  jand g2661(.dina(n2714), .dinb(n2711), .dout(n2715));
  jand g2662(.dina(n232), .dinb(n157), .dout(n2716));
  jand g2663(.dina(n2716), .dinb(n481), .dout(n2717));
  jand g2664(.dina(n246), .dinb(n235), .dout(n2718));
  jand g2665(.dina(n2718), .dinb(n2717), .dout(n2719));
  jand g2666(.dina(n817), .dinb(n904), .dout(n2720));
  jand g2667(.dina(n2720), .dinb(n2719), .dout(n2721));
  jand g2668(.dina(n370), .dinb(n355), .dout(n2722));
  jand g2669(.dina(n226), .dinb(n187), .dout(n2723));
  jand g2670(.dina(n1095), .dinb(n102), .dout(n2724));
  jand g2671(.dina(n2724), .dinb(n429), .dout(n2725));
  jand g2672(.dina(n2725), .dinb(n2723), .dout(n2726));
  jand g2673(.dina(n2726), .dinb(n2722), .dout(n2727));
  jand g2674(.dina(n2727), .dinb(n1135), .dout(n2728));
  jand g2675(.dina(n2728), .dinb(n2721), .dout(n2729));
  jand g2676(.dina(n445), .dinb(n147), .dout(n2730));
  jand g2677(.dina(n2730), .dinb(n240), .dout(n2731));
  jand g2678(.dina(n2731), .dinb(n2729), .dout(n2732));
  jand g2679(.dina(n460), .dinb(n169), .dout(n2733));
  jand g2680(.dina(n2733), .dinb(n600), .dout(n2734));
  jand g2681(.dina(n489), .dinb(n128), .dout(n2735));
  jand g2682(.dina(n2735), .dinb(n378), .dout(n2736));
  jand g2683(.dina(n2736), .dinb(n1093), .dout(n2737));
  jand g2684(.dina(n2737), .dinb(n2734), .dout(n2738));
  jand g2685(.dina(n2738), .dinb(n1105), .dout(n2739));
  jand g2686(.dina(n2739), .dinb(n384), .dout(n2740));
  jand g2687(.dina(n852), .dinb(n439), .dout(n2741));
  jand g2688(.dina(n488), .dinb(n438), .dout(n2742));
  jand g2689(.dina(n2742), .dinb(n280), .dout(n2743));
  jand g2690(.dina(n331), .dinb(n315), .dout(n2744));
  jand g2691(.dina(n510), .dinb(n166), .dout(n2745));
  jand g2692(.dina(n2745), .dinb(n2744), .dout(n2746));
  jand g2693(.dina(n2746), .dinb(n2743), .dout(n2747));
  jand g2694(.dina(n1459), .dinb(n191), .dout(n2748));
  jand g2695(.dina(n2748), .dinb(n456), .dout(n2749));
  jand g2696(.dina(n2749), .dinb(n2747), .dout(n2750));
  jand g2697(.dina(n2750), .dinb(n2741), .dout(n2751));
  jand g2698(.dina(n1452), .dinb(n373), .dout(n2752));
  jand g2699(.dina(n562), .dinb(n377), .dout(n2753));
  jand g2700(.dina(n2753), .dinb(n2752), .dout(n2754));
  jand g2701(.dina(n2142), .dinb(n602), .dout(n2755));
  jand g2702(.dina(n2755), .dinb(n2754), .dout(n2756));
  jand g2703(.dina(n2756), .dinb(n2751), .dout(n2757));
  jand g2704(.dina(n2757), .dinb(n2740), .dout(n2758));
  jand g2705(.dina(n2758), .dinb(n2732), .dout(n2759));
  jand g2706(.dina(n2679), .dinb(n2642), .dout(n2760));
  jand g2707(.dina(n2680), .dinb(n2639), .dout(n2761));
  jor  g2708(.dina(n2761), .dinb(n2760), .dout(n2762));
  jand g2709(.dina(n2661), .dinb(n2645), .dout(n2763));
  jand g2710(.dina(n2678), .dinb(n2662), .dout(n2764));
  jor  g2711(.dina(n2764), .dinb(n2763), .dout(n2765));
  jand g2712(.dina(n2676), .dinb(n2673), .dout(n2766));
  jand g2713(.dina(n2677), .dinb(n2665), .dout(n2767));
  jor  g2714(.dina(n2767), .dinb(n2766), .dout(n2768));
  jand g2715(.dina(n1494), .dinb(n994), .dout(n2769));
  jnot g2716(.din(n2654), .dout(n2770));
  jxor g2717(.dina(n2770), .dinb(n1151), .dout(n2771));
  jxor g2718(.dina(n2771), .dinb(n2769), .dout(n2772));
  jxor g2719(.dina(n2772), .dinb(n2768), .dout(n2773));
  jnot g2720(.din(n2659), .dout(n2774));
  jand g2721(.dina(n2774), .dinb(n2770), .dout(n2775));
  jand g2722(.dina(n2660), .dinb(n2653), .dout(n2776));
  jor  g2723(.dina(n2776), .dinb(n2775), .dout(n2777));
  jand g2724(.dina(n1549), .dinb(n1438), .dout(n2778));
  jand g2725(.dina(n1551), .dinb(n2051), .dout(n2779));
  jor  g2726(.dina(n2779), .dinb(n2778), .dout(n2780));
  jnot g2727(.din(n2780), .dout(n2781));
  jand g2728(.dina(n1558), .dinb(n1434), .dout(n2782));
  jand g2729(.dina(n1560), .dinb(n1622), .dout(n2783));
  jor  g2730(.dina(n2783), .dinb(n2782), .dout(n2784));
  jand g2731(.dina(n2784), .dinb(n2781), .dout(n2785));
  jand g2732(.dina(n1493), .dinb(n1356), .dout(n2786));
  jnot g2733(.din(n2786), .dout(n2787));
  jxor g2734(.dina(n1474), .dinb(n1485), .dout(n2788));
  jor  g2735(.dina(n2788), .dinb(n1490), .dout(n2789));
  jand g2736(.dina(n1505), .dinb(n1480), .dout(n2790));
  jnot g2737(.din(n2790), .dout(n2791));
  jand g2738(.dina(n2791), .dinb(n2789), .dout(n2792));
  jand g2739(.dina(n2792), .dinb(n2787), .dout(n2793));
  jxor g2740(.dina(n2793), .dinb(n2785), .dout(n2794));
  jxor g2741(.dina(n2794), .dinb(n2777), .dout(n2795));
  jxor g2742(.dina(n2795), .dinb(n2773), .dout(n2796));
  jxor g2743(.dina(n2796), .dinb(n2765), .dout(n2797));
  jxor g2744(.dina(n2797), .dinb(n2762), .dout(n2798));
  jxor g2745(.dina(n2798), .dinb(n2759), .dout(n2799));
  jxor g2746(.dina(n2799), .dinb(n2715), .dout(n2800));
  jxor g2747(.dina(n2800), .dinb(n2707), .dout(n2801));
  jxor g2748(.dina(n2801), .dinb(n2710), .dout(n2802));
  jor  g2749(.dina(n2802), .dinb(n2506), .dout(n2803));
  jxor g2750(.dina(n1266), .dinb(n1168), .dout(n2804));
  jnot g2751(.din(n2804), .dout(n2805));
  jand g2752(.dina(n2805), .dinb(n2501), .dout(n2806));
  jnot g2753(.din(n2806), .dout(n2807));
  jor  g2754(.dina(n2807), .dinb(n2707), .dout(n2808));
  jand g2755(.dina(n2503), .dinb(n2502), .dout(n2809));
  jnot g2756(.din(n2809), .dout(n2810));
  jor  g2757(.dina(n2810), .dinb(n2800), .dout(n2811));
  jand g2758(.dina(n2811), .dinb(n2808), .dout(n2812));
  jxor g2759(.dina(n2602), .dinb(n2703), .dout(n2813));
  jand g2760(.dina(n2804), .dinb(n2504), .dout(n2814));
  jand g2761(.dina(n2814), .dinb(n2501), .dout(n2815));
  jnot g2762(.din(n2815), .dout(n2816));
  jor  g2763(.dina(n2816), .dinb(n2813), .dout(n2817));
  jand g2764(.dina(n2817), .dinb(n2812), .dout(n2818));
  jand g2765(.dina(n2818), .dinb(n2803), .dout(n2819));
  jxor g2766(.dina(n2819), .dinb(n1257), .dout(n2820));
  jor  g2767(.dina(n2820), .dinb(n2500), .dout(n2821));
  jxor g2768(.dina(n2364), .dinb(n2251), .dout(n2822));
  jnot g2769(.din(n2822), .dout(n2823));
  jxor g2770(.dina(n2813), .dinb(n2707), .dout(n2824));
  jxor g2771(.dina(n2824), .dinb(n2698), .dout(n2825));
  jor  g2772(.dina(n2825), .dinb(n2506), .dout(n2826));
  jor  g2773(.dina(n2810), .dinb(n2707), .dout(n2827));
  jor  g2774(.dina(n2807), .dinb(n2813), .dout(n2828));
  jand g2775(.dina(n2828), .dinb(n2827), .dout(n2829));
  jor  g2776(.dina(n2816), .dinb(n2471), .dout(n2830));
  jand g2777(.dina(n2830), .dinb(n2829), .dout(n2831));
  jand g2778(.dina(n2831), .dinb(n2826), .dout(n2832));
  jxor g2779(.dina(n2832), .dinb(n1257), .dout(n2833));
  jor  g2780(.dina(n2833), .dinb(n2823), .dout(n2834));
  jxor g2781(.dina(n2813), .dinb(n2471), .dout(n2835));
  jxor g2782(.dina(n2835), .dinb(n2695), .dout(n2836));
  jor  g2783(.dina(n2836), .dinb(n2506), .dout(n2837));
  jor  g2784(.dina(n2807), .dinb(n2471), .dout(n2838));
  jor  g2785(.dina(n2810), .dinb(n2813), .dout(n2839));
  jand g2786(.dina(n2839), .dinb(n2838), .dout(n2840));
  jor  g2787(.dina(n2816), .dinb(n2351), .dout(n2841));
  jand g2788(.dina(n2841), .dinb(n2840), .dout(n2842));
  jand g2789(.dina(n2842), .dinb(n2837), .dout(n2843));
  jxor g2790(.dina(n2843), .dinb(n1257), .dout(n2844));
  jnot g2791(.din(n2844), .dout(n2845));
  jor  g2792(.dina(n2115), .dinb(n1480), .dout(n2846));
  jxor g2793(.dina(n2846), .dinb(n2248), .dout(n2847));
  jand g2794(.dina(n2847), .dinb(n2845), .dout(n2848));
  jor  g2795(.dina(n2506), .dinb(n2473), .dout(n2849));
  jor  g2796(.dina(n2807), .dinb(n2351), .dout(n2850));
  jor  g2797(.dina(n2810), .dinb(n2471), .dout(n2851));
  jand g2798(.dina(n2851), .dinb(n2850), .dout(n2852));
  jor  g2799(.dina(n2816), .dinb(n2256), .dout(n2853));
  jand g2800(.dina(n2853), .dinb(n2852), .dout(n2854));
  jand g2801(.dina(n2854), .dinb(n2849), .dout(n2855));
  jxor g2802(.dina(n2855), .dinb(n1257), .dout(n2856));
  jnot g2803(.din(n2856), .dout(n2857));
  jand g2804(.dina(n2112), .dinb(n1356), .dout(n2858));
  jxor g2805(.dina(n2858), .dinb(n2110), .dout(n2859));
  jand g2806(.dina(n2859), .dinb(n2857), .dout(n2860));
  jand g2807(.dina(n2505), .dinb(n2096), .dout(n2861));
  jand g2808(.dina(n2806), .dinb(n1956), .dout(n2862));
  jand g2809(.dina(n2809), .dinb(n2094), .dout(n2863));
  jor  g2810(.dina(n2863), .dinb(n2862), .dout(n2864));
  jor  g2811(.dina(n2864), .dinb(n2861), .dout(n2865));
  jnot g2812(.din(n2865), .dout(n2866));
  jand g2813(.dina(n2502), .dinb(n1956), .dout(n2867));
  jnot g2814(.din(n2867), .dout(n2868));
  jand g2815(.dina(n2868), .dinb(n1257), .dout(n2869));
  jand g2816(.dina(n2869), .dinb(n2866), .dout(n2870));
  jand g2817(.dina(n2505), .dinb(n2238), .dout(n2871));
  jand g2818(.dina(n2806), .dinb(n2094), .dout(n2872));
  jand g2819(.dina(n2809), .dinb(n2236), .dout(n2873));
  jor  g2820(.dina(n2873), .dinb(n2872), .dout(n2874));
  jand g2821(.dina(n2815), .dinb(n1956), .dout(n2875));
  jor  g2822(.dina(n2875), .dinb(n2874), .dout(n2876));
  jor  g2823(.dina(n2876), .dinb(n2871), .dout(n2877));
  jnot g2824(.din(n2877), .dout(n2878));
  jand g2825(.dina(n2878), .dinb(n2870), .dout(n2879));
  jand g2826(.dina(n2879), .dinb(n2112), .dout(n2880));
  jxor g2827(.dina(n2879), .dinb(n2112), .dout(n2881));
  jor  g2828(.dina(n2506), .dinb(n2353), .dout(n2882));
  jor  g2829(.dina(n2810), .dinb(n2351), .dout(n2883));
  jor  g2830(.dina(n2816), .dinb(n2116), .dout(n2884));
  jor  g2831(.dina(n2807), .dinb(n2256), .dout(n2885));
  jand g2832(.dina(n2885), .dinb(n2884), .dout(n2886));
  jand g2833(.dina(n2886), .dinb(n2883), .dout(n2887));
  jand g2834(.dina(n2887), .dinb(n2882), .dout(n2888));
  jxor g2835(.dina(n2888), .dinb(n1259), .dout(n2889));
  jand g2836(.dina(n2889), .dinb(n2881), .dout(n2890));
  jor  g2837(.dina(n2890), .dinb(n2880), .dout(n2891));
  jxor g2838(.dina(n2859), .dinb(n2857), .dout(n2892));
  jand g2839(.dina(n2892), .dinb(n2891), .dout(n2893));
  jor  g2840(.dina(n2893), .dinb(n2860), .dout(n2894));
  jxor g2841(.dina(n2847), .dinb(n2845), .dout(n2895));
  jand g2842(.dina(n2895), .dinb(n2894), .dout(n2896));
  jor  g2843(.dina(n2896), .dinb(n2848), .dout(n2897));
  jxor g2844(.dina(n2833), .dinb(n2823), .dout(n2898));
  jand g2845(.dina(n2898), .dinb(n2897), .dout(n2899));
  jnot g2846(.din(n2899), .dout(n2900));
  jand g2847(.dina(n2900), .dinb(n2834), .dout(n2901));
  jnot g2848(.din(n2901), .dout(n2902));
  jxor g2849(.dina(n2820), .dinb(n2500), .dout(n2903));
  jand g2850(.dina(n2903), .dinb(n2902), .dout(n2904));
  jnot g2851(.din(n2904), .dout(n2905));
  jand g2852(.dina(n2905), .dinb(n2821), .dout(n2906));
  jand g2853(.dina(n2497), .dinb(n2482), .dout(n2907));
  jand g2854(.dina(n2498), .dinb(n2366), .dout(n2908));
  jor  g2855(.dina(n2908), .dinb(n2907), .dout(n2909));
  jor  g2856(.dina(n2836), .dinb(n2252), .dout(n2910));
  jor  g2857(.dina(n2471), .dinb(n2359), .dout(n2911));
  jor  g2858(.dina(n2813), .dinb(n2355), .dout(n2912));
  jand g2859(.dina(n2912), .dinb(n2911), .dout(n2913));
  jor  g2860(.dina(n2351), .dinb(n2357), .dout(n2914));
  jand g2861(.dina(n2914), .dinb(n2913), .dout(n2915));
  jand g2862(.dina(n2915), .dinb(n2910), .dout(n2916));
  jxor g2863(.dina(n2916), .dinb(n1356), .dout(n2917));
  jnot g2864(.din(n2917), .dout(n2918));
  jand g2865(.dina(n2484), .dinb(n2238), .dout(n2919));
  jand g2866(.dina(n2491), .dinb(n2236), .dout(n2920));
  jand g2867(.dina(n2488), .dinb(n2094), .dout(n2921));
  jand g2868(.dina(n2483), .dinb(n1957), .dout(n2922));
  jand g2869(.dina(n2922), .dinb(n2486), .dout(n2923));
  jand g2870(.dina(n2923), .dinb(n1956), .dout(n2924));
  jor  g2871(.dina(n2924), .dinb(n2921), .dout(n2925));
  jor  g2872(.dina(n2925), .dinb(n2920), .dout(n2926));
  jor  g2873(.dina(n2926), .dinb(n2919), .dout(n2927));
  jor  g2874(.dina(n1959), .dinb(n2051), .dout(n2928));
  jor  g2875(.dina(n2928), .dinb(n2494), .dout(n2929));
  jand g2876(.dina(n2929), .dinb(n1438), .dout(n2930));
  jxor g2877(.dina(n2930), .dinb(n2927), .dout(n2931));
  jxor g2878(.dina(n2931), .dinb(n2918), .dout(n2932));
  jxor g2879(.dina(n2932), .dinb(n2909), .dout(n2933));
  jnot g2880(.din(n2933), .dout(n2934));
  jnot g2881(.din(n2637), .dout(n2935));
  jnot g2882(.din(n2583), .dout(n2936));
  jor  g2883(.dina(n2936), .dinb(n2537), .dout(n2937));
  jand g2884(.dina(n2937), .dinb(n2935), .dout(n2938));
  jxor g2885(.dina(n2680), .dinb(n2938), .dout(n2939));
  jand g2886(.dina(n2939), .dinb(n2712), .dout(n2940));
  jand g2887(.dina(n2682), .dinb(n2604), .dout(n2941));
  jor  g2888(.dina(n2941), .dinb(n2940), .dout(n2942));
  jxor g2889(.dina(n2799), .dinb(n2942), .dout(n2943));
  jand g2890(.dina(n2943), .dinb(n2683), .dout(n2944));
  jnot g2891(.din(n2944), .dout(n2945));
  jxor g2892(.dina(n2943), .dinb(n2707), .dout(n2946));
  jor  g2893(.dina(n2946), .dinb(n2710), .dout(n2947));
  jand g2894(.dina(n2947), .dinb(n2945), .dout(n2948));
  jor  g2895(.dina(n2798), .dinb(n2759), .dout(n2949));
  jnot g2896(.din(n2759), .dout(n2950));
  jxor g2897(.dina(n2798), .dinb(n2950), .dout(n2951));
  jor  g2898(.dina(n2951), .dinb(n2715), .dout(n2952));
  jand g2899(.dina(n2952), .dinb(n2949), .dout(n2953));
  jand g2900(.dina(n535), .dinb(n337), .dout(n2954));
  jand g2901(.dina(n2954), .dinb(n1120), .dout(n2955));
  jand g2902(.dina(n2955), .dinb(n2743), .dout(n2956));
  jand g2903(.dina(n2956), .dinb(n436), .dout(n2957));
  jand g2904(.dina(n1322), .dinb(n137), .dout(n2958));
  jand g2905(.dina(n717), .dinb(n386), .dout(n2959));
  jand g2906(.dina(n2959), .dinb(n2958), .dout(n2960));
  jand g2907(.dina(n2960), .dinb(n2957), .dout(n2961));
  jand g2908(.dina(n1124), .dinb(n396), .dout(n2962));
  jand g2909(.dina(n2962), .dinb(n215), .dout(n2963));
  jand g2910(.dina(n250), .dinb(n204), .dout(n2964));
  jand g2911(.dina(n2964), .dinb(n128), .dout(n2965));
  jand g2912(.dina(n1035), .dinb(n94), .dout(n2966));
  jand g2913(.dina(n2966), .dinb(n388), .dout(n2967));
  jand g2914(.dina(n2967), .dinb(n2965), .dout(n2968));
  jand g2915(.dina(n2968), .dinb(n361), .dout(n2969));
  jand g2916(.dina(n2969), .dinb(n1378), .dout(n2970));
  jand g2917(.dina(n2970), .dinb(n2963), .dout(n2971));
  jand g2918(.dina(n2971), .dinb(n2729), .dout(n2972));
  jand g2919(.dina(n2972), .dinb(n2961), .dout(n2973));
  jand g2920(.dina(n2796), .dinb(n2765), .dout(n2974));
  jand g2921(.dina(n2797), .dinb(n2762), .dout(n2975));
  jor  g2922(.dina(n2975), .dinb(n2974), .dout(n2976));
  jand g2923(.dina(n2772), .dinb(n2768), .dout(n2977));
  jand g2924(.dina(n2795), .dinb(n2773), .dout(n2978));
  jor  g2925(.dina(n2978), .dinb(n2977), .dout(n2979));
  jand g2926(.dina(n1505), .dinb(n1485), .dout(n2980));
  jnot g2927(.din(n2980), .dout(n2981));
  jxor g2928(.dina(n1474), .dinb(n1622), .dout(n2982));
  jor  g2929(.dina(n2982), .dinb(n1490), .dout(n2983));
  jand g2930(.dina(n1493), .dinb(n1360), .dout(n2984));
  jnot g2931(.din(n2984), .dout(n2985));
  jand g2932(.dina(n2985), .dinb(n2983), .dout(n2986));
  jand g2933(.dina(n2986), .dinb(n2981), .dout(n2987));
  jand g2934(.dina(n1494), .dinb(n1356), .dout(n2988));
  jand g2935(.dina(n1438), .dinb(n1555), .dout(n2989));
  jnot g2936(.din(n2989), .dout(n2990));
  jor  g2937(.dina(n2990), .dinb(n1556), .dout(n2991));
  jand g2938(.dina(n2990), .dinb(n1402), .dout(n2992));
  jnot g2939(.din(n2992), .dout(n2993));
  jand g2940(.dina(n2993), .dinb(n2991), .dout(n2994));
  jxor g2941(.dina(n2994), .dinb(n2988), .dout(n2995));
  jxor g2942(.dina(n2995), .dinb(n2987), .dout(n2996));
  jand g2943(.dina(n2654), .dinb(n2655), .dout(n2997));
  jand g2944(.dina(n2771), .dinb(n2769), .dout(n2998));
  jor  g2945(.dina(n2998), .dinb(n2997), .dout(n2999));
  jand g2946(.dina(n2793), .dinb(n2785), .dout(n3000));
  jand g2947(.dina(n2794), .dinb(n2777), .dout(n3001));
  jor  g2948(.dina(n3001), .dinb(n3000), .dout(n3002));
  jxor g2949(.dina(n3002), .dinb(n2999), .dout(n3003));
  jxor g2950(.dina(n3003), .dinb(n2996), .dout(n3004));
  jxor g2951(.dina(n3004), .dinb(n2979), .dout(n3005));
  jxor g2952(.dina(n3005), .dinb(n2976), .dout(n3006));
  jxor g2953(.dina(n3006), .dinb(n2973), .dout(n3007));
  jxor g2954(.dina(n3007), .dinb(n2953), .dout(n3008));
  jxor g2955(.dina(n3008), .dinb(n2800), .dout(n3009));
  jxor g2956(.dina(n3009), .dinb(n2948), .dout(n3010));
  jor  g2957(.dina(n3010), .dinb(n2506), .dout(n3011));
  jor  g2958(.dina(n3008), .dinb(n2810), .dout(n3012));
  jor  g2959(.dina(n2807), .dinb(n2800), .dout(n3013));
  jand g2960(.dina(n3013), .dinb(n3012), .dout(n3014));
  jor  g2961(.dina(n2816), .dinb(n2707), .dout(n3015));
  jand g2962(.dina(n3015), .dinb(n3014), .dout(n3016));
  jand g2963(.dina(n3016), .dinb(n3011), .dout(n3017));
  jxor g2964(.dina(n3017), .dinb(n1257), .dout(n3018));
  jxor g2965(.dina(n3018), .dinb(n2934), .dout(n3019));
  jxor g2966(.dina(n3019), .dinb(n2906), .dout(n3020));
  jnot g2967(.din(a2 ), .dout(n3021));
  jand g2968(.dina(n50), .dinb(n49), .dout(n3022));
  jxor g2969(.dina(n3022), .dinb(n3021), .dout(n3023));
  jxor g2970(.dina(n3023), .dinb(n519), .dout(n3024));
  jnot g2971(.din(n3024), .dout(n3025));
  jxor g2972(.dina(n1500), .dinb(n1154), .dout(n3026));
  jnot g2973(.din(n3026), .dout(n3027));
  jand g2974(.dina(n3027), .dinb(n3025), .dout(n3028));
  jnot g2975(.din(n3028), .dout(n3029));
  jand g2976(.dina(n1102), .dinb(n275), .dout(n3030));
  jand g2977(.dina(n3030), .dinb(n398), .dout(n3031));
  jand g2978(.dina(n3031), .dinb(n1375), .dout(n3032));
  jand g2979(.dina(n525), .dinb(n248), .dout(n3033));
  jand g2980(.dina(n3033), .dinb(n437), .dout(n3034));
  jand g2981(.dina(n817), .dinb(n366), .dout(n3035));
  jand g2982(.dina(n3035), .dinb(n460), .dout(n3036));
  jand g2983(.dina(n3036), .dinb(n3034), .dout(n3037));
  jand g2984(.dina(n3037), .dinb(n1196), .dout(n3038));
  jand g2985(.dina(n3038), .dinb(n3032), .dout(n3039));
  jand g2986(.dina(n537), .dinb(n344), .dout(n3040));
  jand g2987(.dina(n3040), .dinb(n3039), .dout(n3041));
  jand g2988(.dina(n3041), .dinb(n896), .dout(n3042));
  jnot g2989(.din(n3042), .dout(n3043));
  jand g2990(.dina(n3004), .dinb(n2979), .dout(n3044));
  jnot g2991(.din(n3044), .dout(n3045));
  jnot g2992(.din(n2974), .dout(n3046));
  jnot g2993(.din(n2760), .dout(n3047));
  jnot g2994(.din(n2680), .dout(n3048));
  jor  g2995(.dina(n3048), .dinb(n2938), .dout(n3049));
  jand g2996(.dina(n3049), .dinb(n3047), .dout(n3050));
  jnot g2997(.din(n2797), .dout(n3051));
  jor  g2998(.dina(n3051), .dinb(n3050), .dout(n3052));
  jand g2999(.dina(n3052), .dinb(n3046), .dout(n3053));
  jnot g3000(.din(n3005), .dout(n3054));
  jor  g3001(.dina(n3054), .dinb(n3053), .dout(n3055));
  jand g3002(.dina(n3055), .dinb(n3045), .dout(n3056));
  jand g3003(.dina(n3002), .dinb(n2999), .dout(n3057));
  jand g3004(.dina(n3003), .dinb(n2996), .dout(n3058));
  jor  g3005(.dina(n3058), .dinb(n3057), .dout(n3059));
  jand g3006(.dina(n1493), .dinb(n1434), .dout(n3060));
  jxor g3007(.dina(n1474), .dinb(n1438), .dout(n3061));
  jand g3008(.dina(n3061), .dinb(n517), .dout(n3062));
  jand g3009(.dina(n1505), .dinb(n1622), .dout(n3063));
  jor  g3010(.dina(n3063), .dinb(n3062), .dout(n3064));
  jor  g3011(.dina(n3064), .dinb(n3060), .dout(n3065));
  jor  g3012(.dina(n2994), .dinb(n2988), .dout(n3066));
  jand g3013(.dina(n2995), .dinb(n2987), .dout(n3067));
  jnot g3014(.din(n3067), .dout(n3068));
  jand g3015(.dina(n3068), .dinb(n3066), .dout(n3069));
  jxor g3016(.dina(n3069), .dinb(n3065), .dout(n3070));
  jand g3017(.dina(n1494), .dinb(n1360), .dout(n3071));
  jnot g3018(.din(n2988), .dout(n3072));
  jxor g3019(.dina(n3072), .dinb(n1402), .dout(n3073));
  jxor g3020(.dina(n3073), .dinb(n3071), .dout(n3074));
  jxor g3021(.dina(n3074), .dinb(n3070), .dout(n3075));
  jxor g3022(.dina(n3075), .dinb(n3059), .dout(n3076));
  jxor g3023(.dina(n3076), .dinb(n3056), .dout(n3077));
  jand g3024(.dina(n3077), .dinb(n3043), .dout(n3078));
  jnot g3025(.din(n2973), .dout(n3079));
  jxor g3026(.dina(n3005), .dinb(n3053), .dout(n3080));
  jand g3027(.dina(n3080), .dinb(n3079), .dout(n3081));
  jxor g3028(.dina(n2797), .dinb(n3050), .dout(n3082));
  jand g3029(.dina(n3082), .dinb(n2950), .dout(n3083));
  jand g3030(.dina(n2799), .dinb(n2942), .dout(n3084));
  jor  g3031(.dina(n3084), .dinb(n3083), .dout(n3085));
  jand g3032(.dina(n3007), .dinb(n3085), .dout(n3086));
  jor  g3033(.dina(n3086), .dinb(n3081), .dout(n3087));
  jand g3034(.dina(n3005), .dinb(n2976), .dout(n3088));
  jor  g3035(.dina(n3088), .dinb(n3044), .dout(n3089));
  jxor g3036(.dina(n3076), .dinb(n3089), .dout(n3090));
  jxor g3037(.dina(n3090), .dinb(n3042), .dout(n3091));
  jand g3038(.dina(n3091), .dinb(n3087), .dout(n3092));
  jor  g3039(.dina(n3092), .dinb(n3078), .dout(n3093));
  jand g3040(.dina(n1095), .dinb(n359), .dout(n3094));
  jand g3041(.dina(n429), .dinb(n94), .dout(n3095));
  jand g3042(.dina(n434), .dinb(n366), .dout(n3096));
  jand g3043(.dina(n3096), .dinb(n389), .dout(n3097));
  jand g3044(.dina(n3097), .dinb(n3095), .dout(n3098));
  jand g3045(.dina(n252), .dinb(n187), .dout(n3099));
  jand g3046(.dina(n3099), .dinb(n1017), .dout(n3100));
  jand g3047(.dina(n3100), .dinb(n3098), .dout(n3101));
  jand g3048(.dina(n309), .dinb(n303), .dout(n3102));
  jand g3049(.dina(n1073), .dinb(n395), .dout(n3103));
  jand g3050(.dina(n3103), .dinb(n222), .dout(n3104));
  jand g3051(.dina(n3104), .dinb(n3102), .dout(n3105));
  jand g3052(.dina(n3105), .dinb(n3101), .dout(n3106));
  jand g3053(.dina(n3106), .dinb(n897), .dout(n3107));
  jand g3054(.dina(n1110), .dinb(n221), .dout(n3108));
  jand g3055(.dina(n3108), .dinb(n2717), .dout(n3109));
  jand g3056(.dina(n3109), .dinb(n1039), .dout(n3110));
  jand g3057(.dina(n3110), .dinb(n240), .dout(n3111));
  jand g3058(.dina(n3111), .dinb(n3107), .dout(n3112));
  jand g3059(.dina(n1460), .dinb(n148), .dout(n3113));
  jand g3060(.dina(n3113), .dinb(n439), .dout(n3114));
  jand g3061(.dina(n3114), .dinb(n2738), .dout(n3115));
  jand g3062(.dina(n3115), .dinb(n278), .dout(n3116));
  jand g3063(.dina(n3116), .dinb(n3112), .dout(n3117));
  jand g3064(.dina(n3117), .dinb(n3094), .dout(n3118));
  jand g3065(.dina(n3075), .dinb(n3059), .dout(n3119));
  jand g3066(.dina(n3076), .dinb(n3089), .dout(n3120));
  jor  g3067(.dina(n3120), .dinb(n3119), .dout(n3121));
  jor  g3068(.dina(n3069), .dinb(n3065), .dout(n3122));
  jand g3069(.dina(n3074), .dinb(n3070), .dout(n3123));
  jnot g3070(.din(n3123), .dout(n3124));
  jand g3071(.dina(n3124), .dinb(n3122), .dout(n3125));
  jnot g3072(.din(n3125), .dout(n3126));
  jand g3073(.dina(n3073), .dinb(n3071), .dout(n3128));
  jnot g3074(.din(n3128), .dout(n3129));
  jand g3075(.dina(n3129), .dinb(n3072), .dout(n3130));
  jand g3076(.dina(n1494), .dinb(n1434), .dout(n3131));
  jand g3077(.dina(n1438), .dinb(n1490), .dout(n3132));
  jnot g3078(.din(n3132), .dout(n3133));
  jor  g3079(.dina(n3133), .dinb(n1493), .dout(n3134));
  jor  g3080(.dina(n3132), .dinb(n1474), .dout(n3135));
  jand g3081(.dina(n3135), .dinb(n3134), .dout(n3136));
  jxor g3082(.dina(n3136), .dinb(n3131), .dout(n3137));
  jnot g3083(.din(n3137), .dout(n3138));
  jxor g3084(.dina(n3138), .dinb(n3130), .dout(n3139));
  jxor g3085(.dina(n3139), .dinb(n3126), .dout(n3140));
  jxor g3086(.dina(n3140), .dinb(n3121), .dout(n3141));
  jxor g3087(.dina(n3141), .dinb(n3118), .dout(n3142));
  jxor g3088(.dina(n3142), .dinb(n3093), .dout(n3143));
  jxor g3089(.dina(n3091), .dinb(n3087), .dout(n3144));
  jand g3090(.dina(n3144), .dinb(n3143), .dout(n3145));
  jnot g3091(.din(n3145), .dout(n3146));
  jxor g3092(.dina(n3007), .dinb(n3085), .dout(n3147));
  jand g3093(.dina(n3144), .dinb(n3147), .dout(n3148));
  jnot g3094(.din(n3148), .dout(n3149));
  jand g3095(.dina(n3147), .dinb(n2943), .dout(n3150));
  jnot g3096(.din(n3150), .dout(n3151));
  jxor g3097(.dina(n3147), .dinb(n2800), .dout(n3152));
  jor  g3098(.dina(n3152), .dinb(n2948), .dout(n3153));
  jand g3099(.dina(n3153), .dinb(n3151), .dout(n3154));
  jxor g3100(.dina(n3144), .dinb(n3008), .dout(n3155));
  jor  g3101(.dina(n3155), .dinb(n3154), .dout(n3156));
  jand g3102(.dina(n3156), .dinb(n3149), .dout(n3157));
  jor  g3103(.dina(n3090), .dinb(n3042), .dout(n3158));
  jor  g3104(.dina(n3006), .dinb(n2973), .dout(n3159));
  jxor g3105(.dina(n3006), .dinb(n3079), .dout(n3160));
  jor  g3106(.dina(n3160), .dinb(n2953), .dout(n3161));
  jand g3107(.dina(n3161), .dinb(n3159), .dout(n3162));
  jxor g3108(.dina(n3090), .dinb(n3043), .dout(n3163));
  jor  g3109(.dina(n3163), .dinb(n3162), .dout(n3164));
  jand g3110(.dina(n3164), .dinb(n3158), .dout(n3165));
  jxor g3111(.dina(n3142), .dinb(n3165), .dout(n3166));
  jxor g3112(.dina(n3144), .dinb(n3166), .dout(n3167));
  jor  g3113(.dina(n3167), .dinb(n3157), .dout(n3168));
  jand g3114(.dina(n3168), .dinb(n3146), .dout(n3169));
  jor  g3115(.dina(n3141), .dinb(n3118), .dout(n3170));
  jnot g3116(.din(n3118), .dout(n3171));
  jxor g3117(.dina(n3141), .dinb(n3171), .dout(n3172));
  jor  g3118(.dina(n3172), .dinb(n3165), .dout(n3173));
  jand g3119(.dina(n3173), .dinb(n3170), .dout(n3174));
  jand g3120(.dina(n587), .dinb(n275), .dout(n3175));
  jand g3121(.dina(n3175), .dinb(n389), .dout(n3176));
  jand g3122(.dina(n3176), .dinb(n2725), .dout(n3177));
  jand g3123(.dina(n3177), .dinb(n198), .dout(n3178));
  jand g3124(.dina(n825), .dinb(n142), .dout(n3179));
  jand g3125(.dina(n3179), .dinb(n1979), .dout(n3180));
  jand g3126(.dina(n3180), .dinb(n3178), .dout(n3181));
  jand g3127(.dina(n3181), .dinb(n2147), .dout(n3182));
  jand g3128(.dina(n1005), .dinb(n717), .dout(n3183));
  jand g3129(.dina(n3183), .dinb(n2744), .dout(n3184));
  jand g3130(.dina(n3184), .dinb(n286), .dout(n3185));
  jand g3131(.dina(n3185), .dinb(n1366), .dout(n3186));
  jand g3132(.dina(n3186), .dinb(n912), .dout(n3187));
  jand g3133(.dina(n3187), .dinb(n468), .dout(n3188));
  jand g3134(.dina(n3188), .dinb(n3182), .dout(n3189));
  jand g3135(.dina(n3189), .dinb(n2386), .dout(n3190));
  jnot g3136(.din(n3190), .dout(n3191));
  jand g3137(.dina(n3139), .dinb(n3126), .dout(n3192));
  jand g3138(.dina(n3140), .dinb(n3121), .dout(n3193));
  jor  g3139(.dina(n3193), .dinb(n3192), .dout(n3194));
  jxor g3140(.dina(n2483), .dinb(n1442), .dout(n3195));
  jor  g3141(.dina(n3195), .dinb(n1474), .dout(n3196));
  jor  g3142(.dina(n3136), .dinb(n3131), .dout(n3197));
  jor  g3143(.dina(n3138), .dinb(n3130), .dout(n3198));
  jand g3144(.dina(n3198), .dinb(n3197), .dout(n3199));
  jxor g3145(.dina(n3199), .dinb(n3196), .dout(n3200));
  jxor g3146(.dina(n3200), .dinb(n3194), .dout(n3201));
  jxor g3147(.dina(n3201), .dinb(n3191), .dout(n3202));
  jxor g3148(.dina(n3202), .dinb(n3174), .dout(n3203));
  jxor g3149(.dina(n3203), .dinb(n3166), .dout(n3204));
  jxor g3150(.dina(n3204), .dinb(n3169), .dout(n3205));
  jor  g3151(.dina(n3205), .dinb(n3029), .dout(n3206));
  jxor g3152(.dina(n1499), .dinb(n1504), .dout(n3207));
  jnot g3153(.din(n3207), .dout(n3208));
  jand g3154(.dina(n3208), .dinb(n3024), .dout(n3209));
  jnot g3155(.din(n3209), .dout(n3210));
  jor  g3156(.dina(n3210), .dinb(n3166), .dout(n3211));
  jand g3157(.dina(n3026), .dinb(n3025), .dout(n3212));
  jnot g3158(.din(n3212), .dout(n3213));
  jor  g3159(.dina(n3213), .dinb(n3203), .dout(n3214));
  jand g3160(.dina(n3214), .dinb(n3211), .dout(n3215));
  jxor g3161(.dina(n3091), .dinb(n3162), .dout(n3216));
  jand g3162(.dina(n3207), .dinb(n3024), .dout(n3217));
  jand g3163(.dina(n3217), .dinb(n3027), .dout(n3218));
  jnot g3164(.din(n3218), .dout(n3219));
  jor  g3165(.dina(n3219), .dinb(n3216), .dout(n3220));
  jand g3166(.dina(n3220), .dinb(n3215), .dout(n3221));
  jand g3167(.dina(n3221), .dinb(n3206), .dout(n3222));
  jxor g3168(.dina(n3222), .dinb(n1154), .dout(n3223));
  jor  g3169(.dina(n3223), .dinb(n3020), .dout(n3224));
  jnot g3170(.din(n3224), .dout(n3225));
  jxor g3171(.dina(n2903), .dinb(n2902), .dout(n3226));
  jnot g3172(.din(n3226), .dout(n3227));
  jxor g3173(.dina(n3216), .dinb(n3166), .dout(n3228));
  jxor g3174(.dina(n3228), .dinb(n3157), .dout(n3229));
  jor  g3175(.dina(n3229), .dinb(n3029), .dout(n3230));
  jor  g3176(.dina(n3213), .dinb(n3166), .dout(n3231));
  jor  g3177(.dina(n3210), .dinb(n3216), .dout(n3232));
  jand g3178(.dina(n3232), .dinb(n3231), .dout(n3233));
  jor  g3179(.dina(n3219), .dinb(n3008), .dout(n3234));
  jand g3180(.dina(n3234), .dinb(n3233), .dout(n3235));
  jand g3181(.dina(n3235), .dinb(n3230), .dout(n3236));
  jxor g3182(.dina(n3236), .dinb(n1154), .dout(n3237));
  jor  g3183(.dina(n3237), .dinb(n3227), .dout(n3238));
  jnot g3184(.din(n3238), .dout(n3239));
  jxor g3185(.dina(n2898), .dinb(n2897), .dout(n3240));
  jxor g3186(.dina(n3216), .dinb(n3008), .dout(n3241));
  jxor g3187(.dina(n3241), .dinb(n3154), .dout(n3242));
  jor  g3188(.dina(n3242), .dinb(n3029), .dout(n3243));
  jor  g3189(.dina(n3213), .dinb(n3216), .dout(n3244));
  jor  g3190(.dina(n3210), .dinb(n3008), .dout(n3245));
  jor  g3191(.dina(n3219), .dinb(n2800), .dout(n3246));
  jand g3192(.dina(n3246), .dinb(n3245), .dout(n3247));
  jand g3193(.dina(n3247), .dinb(n3244), .dout(n3248));
  jand g3194(.dina(n3248), .dinb(n3243), .dout(n3249));
  jxor g3195(.dina(n3249), .dinb(n1156), .dout(n3250));
  jand g3196(.dina(n3250), .dinb(n3240), .dout(n3251));
  jxor g3197(.dina(n2895), .dinb(n2894), .dout(n3252));
  jor  g3198(.dina(n3029), .dinb(n3010), .dout(n3253));
  jor  g3199(.dina(n3210), .dinb(n2800), .dout(n3254));
  jor  g3200(.dina(n3213), .dinb(n3008), .dout(n3255));
  jor  g3201(.dina(n3219), .dinb(n2707), .dout(n3256));
  jand g3202(.dina(n3256), .dinb(n3255), .dout(n3257));
  jand g3203(.dina(n3257), .dinb(n3254), .dout(n3258));
  jand g3204(.dina(n3258), .dinb(n3253), .dout(n3259));
  jxor g3205(.dina(n3259), .dinb(n1156), .dout(n3260));
  jand g3206(.dina(n3260), .dinb(n3252), .dout(n3261));
  jxor g3207(.dina(n2892), .dinb(n2891), .dout(n3262));
  jor  g3208(.dina(n3029), .dinb(n2802), .dout(n3263));
  jor  g3209(.dina(n3213), .dinb(n2800), .dout(n3264));
  jor  g3210(.dina(n3210), .dinb(n2707), .dout(n3265));
  jor  g3211(.dina(n3219), .dinb(n2813), .dout(n3266));
  jand g3212(.dina(n3266), .dinb(n3265), .dout(n3267));
  jand g3213(.dina(n3267), .dinb(n3264), .dout(n3268));
  jand g3214(.dina(n3268), .dinb(n3263), .dout(n3269));
  jxor g3215(.dina(n3269), .dinb(n1156), .dout(n3270));
  jand g3216(.dina(n3270), .dinb(n3262), .dout(n3271));
  jxor g3217(.dina(n2889), .dinb(n2881), .dout(n3272));
  jor  g3218(.dina(n3029), .dinb(n2825), .dout(n3273));
  jor  g3219(.dina(n3210), .dinb(n2813), .dout(n3274));
  jor  g3220(.dina(n3213), .dinb(n2707), .dout(n3275));
  jor  g3221(.dina(n3219), .dinb(n2471), .dout(n3276));
  jand g3222(.dina(n3276), .dinb(n3275), .dout(n3277));
  jand g3223(.dina(n3277), .dinb(n3274), .dout(n3278));
  jand g3224(.dina(n3278), .dinb(n3273), .dout(n3279));
  jxor g3225(.dina(n3279), .dinb(n1156), .dout(n3280));
  jand g3226(.dina(n3280), .dinb(n3272), .dout(n3281));
  jor  g3227(.dina(n3029), .dinb(n2836), .dout(n3282));
  jor  g3228(.dina(n3210), .dinb(n2471), .dout(n3283));
  jor  g3229(.dina(n3213), .dinb(n2813), .dout(n3284));
  jand g3230(.dina(n3284), .dinb(n3283), .dout(n3285));
  jor  g3231(.dina(n3219), .dinb(n2351), .dout(n3286));
  jand g3232(.dina(n3286), .dinb(n3285), .dout(n3287));
  jand g3233(.dina(n3287), .dinb(n3282), .dout(n3288));
  jxor g3234(.dina(n3288), .dinb(n1154), .dout(n3289));
  jnot g3235(.din(n3289), .dout(n3290));
  jor  g3236(.dina(n2870), .dinb(n1259), .dout(n3291));
  jxor g3237(.dina(n3291), .dinb(n2878), .dout(n3292));
  jand g3238(.dina(n3292), .dinb(n3290), .dout(n3293));
  jor  g3239(.dina(n3029), .dinb(n2473), .dout(n3294));
  jor  g3240(.dina(n3210), .dinb(n2351), .dout(n3295));
  jor  g3241(.dina(n3213), .dinb(n2471), .dout(n3296));
  jand g3242(.dina(n3296), .dinb(n3295), .dout(n3297));
  jor  g3243(.dina(n3219), .dinb(n2256), .dout(n3298));
  jand g3244(.dina(n3298), .dinb(n3297), .dout(n3299));
  jand g3245(.dina(n3299), .dinb(n3294), .dout(n3300));
  jxor g3246(.dina(n3300), .dinb(n1154), .dout(n3301));
  jnot g3247(.din(n3301), .dout(n3302));
  jand g3248(.dina(n2867), .dinb(n1257), .dout(n3303));
  jxor g3249(.dina(n3303), .dinb(n2865), .dout(n3304));
  jand g3250(.dina(n3304), .dinb(n3302), .dout(n3305));
  jand g3251(.dina(n3028), .dinb(n2096), .dout(n3306));
  jand g3252(.dina(n3212), .dinb(n2094), .dout(n3307));
  jand g3253(.dina(n3209), .dinb(n1956), .dout(n3308));
  jor  g3254(.dina(n3308), .dinb(n3307), .dout(n3309));
  jor  g3255(.dina(n3309), .dinb(n3306), .dout(n3310));
  jnot g3256(.din(n3310), .dout(n3311));
  jand g3257(.dina(n3025), .dinb(n1956), .dout(n3312));
  jnot g3258(.din(n3312), .dout(n3313));
  jand g3259(.dina(n3313), .dinb(n1154), .dout(n3314));
  jand g3260(.dina(n3314), .dinb(n3311), .dout(n3315));
  jand g3261(.dina(n3028), .dinb(n2238), .dout(n3316));
  jand g3262(.dina(n3212), .dinb(n2236), .dout(n3317));
  jand g3263(.dina(n3209), .dinb(n2094), .dout(n3318));
  jand g3264(.dina(n3218), .dinb(n1956), .dout(n3319));
  jor  g3265(.dina(n3319), .dinb(n3318), .dout(n3320));
  jor  g3266(.dina(n3320), .dinb(n3317), .dout(n3321));
  jor  g3267(.dina(n3321), .dinb(n3316), .dout(n3322));
  jnot g3268(.din(n3322), .dout(n3323));
  jand g3269(.dina(n3323), .dinb(n3315), .dout(n3324));
  jand g3270(.dina(n3324), .dinb(n2867), .dout(n3325));
  jxor g3271(.dina(n3324), .dinb(n2867), .dout(n3326));
  jor  g3272(.dina(n3029), .dinb(n2353), .dout(n3327));
  jor  g3273(.dina(n3213), .dinb(n2351), .dout(n3328));
  jor  g3274(.dina(n3219), .dinb(n2116), .dout(n3329));
  jor  g3275(.dina(n3210), .dinb(n2256), .dout(n3330));
  jand g3276(.dina(n3330), .dinb(n3329), .dout(n3331));
  jand g3277(.dina(n3331), .dinb(n3328), .dout(n3332));
  jand g3278(.dina(n3332), .dinb(n3327), .dout(n3333));
  jxor g3279(.dina(n3333), .dinb(n1156), .dout(n3334));
  jand g3280(.dina(n3334), .dinb(n3326), .dout(n3335));
  jor  g3281(.dina(n3335), .dinb(n3325), .dout(n3336));
  jnot g3282(.din(n3336), .dout(n3337));
  jxor g3283(.dina(n3304), .dinb(n3301), .dout(n3338));
  jor  g3284(.dina(n3338), .dinb(n3337), .dout(n3339));
  jnot g3285(.din(n3339), .dout(n3340));
  jor  g3286(.dina(n3340), .dinb(n3305), .dout(n3341));
  jxor g3287(.dina(n3292), .dinb(n3289), .dout(n3342));
  jnot g3288(.din(n3342), .dout(n3343));
  jand g3289(.dina(n3343), .dinb(n3341), .dout(n3344));
  jor  g3290(.dina(n3344), .dinb(n3293), .dout(n3345));
  jxor g3291(.dina(n3280), .dinb(n3272), .dout(n3346));
  jand g3292(.dina(n3346), .dinb(n3345), .dout(n3347));
  jor  g3293(.dina(n3347), .dinb(n3281), .dout(n3348));
  jxor g3294(.dina(n3270), .dinb(n3262), .dout(n3349));
  jand g3295(.dina(n3349), .dinb(n3348), .dout(n3350));
  jor  g3296(.dina(n3350), .dinb(n3271), .dout(n3351));
  jxor g3297(.dina(n3260), .dinb(n3252), .dout(n3352));
  jand g3298(.dina(n3352), .dinb(n3351), .dout(n3353));
  jor  g3299(.dina(n3353), .dinb(n3261), .dout(n3354));
  jxor g3300(.dina(n3250), .dinb(n3240), .dout(n3355));
  jand g3301(.dina(n3355), .dinb(n3354), .dout(n3356));
  jor  g3302(.dina(n3356), .dinb(n3251), .dout(n3357));
  jxor g3303(.dina(n3237), .dinb(n3227), .dout(n3358));
  jand g3304(.dina(n3358), .dinb(n3357), .dout(n3359));
  jor  g3305(.dina(n3359), .dinb(n3239), .dout(n3360));
  jxor g3306(.dina(n3223), .dinb(n3020), .dout(n3361));
  jand g3307(.dina(n3361), .dinb(n3360), .dout(n3362));
  jor  g3308(.dina(n3362), .dinb(n3225), .dout(n3363));
  jor  g3309(.dina(n3018), .dinb(n2934), .dout(n3364));
  jnot g3310(.din(n3364), .dout(n3365));
  jnot g3311(.din(n2906), .dout(n3366));
  jand g3312(.dina(n3019), .dinb(n3366), .dout(n3367));
  jor  g3313(.dina(n3367), .dinb(n3365), .dout(n3368));
  jand g3314(.dina(n2931), .dinb(n2918), .dout(n3369));
  jand g3315(.dina(n2932), .dinb(n2909), .dout(n3370));
  jor  g3316(.dina(n3370), .dinb(n3369), .dout(n3371));
  jor  g3317(.dina(n2825), .dinb(n2252), .dout(n3372));
  jor  g3318(.dina(n2707), .dinb(n2355), .dout(n3373));
  jor  g3319(.dina(n2813), .dinb(n2359), .dout(n3374));
  jand g3320(.dina(n3374), .dinb(n3373), .dout(n3375));
  jor  g3321(.dina(n2471), .dinb(n2357), .dout(n3376));
  jand g3322(.dina(n3376), .dinb(n3375), .dout(n3377));
  jand g3323(.dina(n3377), .dinb(n3372), .dout(n3378));
  jxor g3324(.dina(n3378), .dinb(n1356), .dout(n3379));
  jnot g3325(.din(n3379), .dout(n3380));
  jnot g3326(.din(n2495), .dout(n3381));
  jor  g3327(.dina(n2929), .dinb(n2927), .dout(n3382));
  jxor g3328(.dina(n3382), .dinb(n3381), .dout(n3383));
  jnot g3329(.din(n2484), .dout(n3384));
  jor  g3330(.dina(n3384), .dinb(n2353), .dout(n3385));
  jnot g3331(.din(n2491), .dout(n3386));
  jor  g3332(.dina(n3386), .dinb(n2351), .dout(n3387));
  jnot g3333(.din(n2923), .dout(n3388));
  jor  g3334(.dina(n3388), .dinb(n2116), .dout(n3389));
  jnot g3335(.din(n2488), .dout(n3390));
  jor  g3336(.dina(n3390), .dinb(n2256), .dout(n3391));
  jand g3337(.dina(n3391), .dinb(n3389), .dout(n3392));
  jand g3338(.dina(n3392), .dinb(n3387), .dout(n3393));
  jand g3339(.dina(n3393), .dinb(n3385), .dout(n3394));
  jxor g3340(.dina(n3394), .dinb(n2051), .dout(n3395));
  jxor g3341(.dina(n3395), .dinb(n3383), .dout(n3396));
  jxor g3342(.dina(n3396), .dinb(n3380), .dout(n3397));
  jxor g3343(.dina(n3397), .dinb(n3371), .dout(n3398));
  jnot g3344(.din(n3398), .dout(n3399));
  jor  g3345(.dina(n3242), .dinb(n2506), .dout(n3400));
  jor  g3346(.dina(n3008), .dinb(n2807), .dout(n3401));
  jor  g3347(.dina(n3216), .dinb(n2810), .dout(n3402));
  jand g3348(.dina(n3402), .dinb(n3401), .dout(n3403));
  jor  g3349(.dina(n2816), .dinb(n2800), .dout(n3404));
  jand g3350(.dina(n3404), .dinb(n3403), .dout(n3405));
  jand g3351(.dina(n3405), .dinb(n3400), .dout(n3406));
  jxor g3352(.dina(n3406), .dinb(n1257), .dout(n3407));
  jxor g3353(.dina(n3407), .dinb(n3399), .dout(n3408));
  jxor g3354(.dina(n3408), .dinb(n3368), .dout(n3409));
  jnot g3355(.din(n3140), .dout(n3410));
  jxor g3356(.dina(n3410), .dinb(n3121), .dout(n3411));
  jand g3357(.dina(n3411), .dinb(n3171), .dout(n3412));
  jand g3358(.dina(n3142), .dinb(n3093), .dout(n3413));
  jor  g3359(.dina(n3413), .dinb(n3412), .dout(n3414));
  jxor g3360(.dina(n3202), .dinb(n3414), .dout(n3415));
  jand g3361(.dina(n3415), .dinb(n3143), .dout(n3416));
  jnot g3362(.din(n3416), .dout(n3417));
  jxor g3363(.dina(n3203), .dinb(n3143), .dout(n3418));
  jor  g3364(.dina(n3418), .dinb(n3169), .dout(n3419));
  jand g3365(.dina(n3419), .dinb(n3417), .dout(n3420));
  jand g3366(.dina(n1331), .dinb(n335), .dout(n3421));
  jand g3367(.dina(n436), .dinb(n218), .dout(n3422));
  jand g3368(.dina(n3422), .dinb(n1385), .dout(n3423));
  jand g3369(.dina(n3423), .dinb(n337), .dout(n3424));
  jand g3370(.dina(n3424), .dinb(n3421), .dout(n3425));
  jand g3371(.dina(n1066), .dinb(n427), .dout(n3426));
  jand g3372(.dina(n283), .dinb(n215), .dout(n3427));
  jand g3373(.dina(n3427), .dinb(n3426), .dout(n3428));
  jand g3374(.dina(n3428), .dinb(n1104), .dout(n3429));
  jand g3375(.dina(n567), .dinb(n527), .dout(n3430));
  jand g3376(.dina(n3430), .dinb(n378), .dout(n3431));
  jand g3377(.dina(n3431), .dinb(n1987), .dout(n3432));
  jand g3378(.dina(n3432), .dinb(n3429), .dout(n3433));
  jand g3379(.dina(n3433), .dinb(n129), .dout(n3434));
  jand g3380(.dina(n3434), .dinb(n3425), .dout(n3435));
  jnot g3381(.din(n3435), .dout(n3436));
  jor  g3382(.dina(n3201), .dinb(n3191), .dout(n3437));
  jand g3383(.dina(n3201), .dinb(n3191), .dout(n3438));
  jor  g3384(.dina(n3438), .dinb(n3414), .dout(n3439));
  jand g3385(.dina(n3439), .dinb(n3437), .dout(n3440));
  jxor g3386(.dina(n3440), .dinb(n3436), .dout(n3441));
  jxor g3387(.dina(n3441), .dinb(n3203), .dout(n3442));
  jxor g3388(.dina(n3442), .dinb(n3420), .dout(n3443));
  jor  g3389(.dina(n3443), .dinb(n3029), .dout(n3444));
  jor  g3390(.dina(n3210), .dinb(n3203), .dout(n3445));
  jor  g3391(.dina(n3441), .dinb(n3213), .dout(n3446));
  jor  g3392(.dina(n3219), .dinb(n3166), .dout(n3447));
  jand g3393(.dina(n3447), .dinb(n3446), .dout(n3448));
  jand g3394(.dina(n3448), .dinb(n3445), .dout(n3449));
  jand g3395(.dina(n3449), .dinb(n3444), .dout(n3450));
  jxor g3396(.dina(n3450), .dinb(n1156), .dout(n3451));
  jxor g3397(.dina(n3451), .dinb(n3409), .dout(n3452));
  jxor g3398(.dina(n3452), .dinb(n3363), .dout(n3453));
  jnot g3399(.din(n3453), .dout(n3454));
  jnot g3400(.din(n3023), .dout(n3455));
  jnot g3401(.din(a0 ), .dout(n3456));
  jor  g3402(.dina(a22 ), .dinb(n3456), .dout(n3457));
  jxor g3403(.dina(n3457), .dinb(a1 ), .dout(n3458));
  jxor g3404(.dina(n3458), .dinb(n3023), .dout(n3459));
  jand g3405(.dina(n3459), .dinb(a0 ), .dout(n3460));
  jnot g3406(.din(n3460), .dout(n3461));
  jnot g3407(.din(n3200), .dout(n3462));
  jxor g3408(.dina(n3462), .dinb(n3194), .dout(n3463));
  jand g3409(.dina(n3463), .dinb(n3190), .dout(n3464));
  jor  g3410(.dina(n3463), .dinb(n3190), .dout(n3465));
  jand g3411(.dina(n3465), .dinb(n3174), .dout(n3466));
  jor  g3412(.dina(n3466), .dinb(n3464), .dout(n3467));
  jand g3413(.dina(n3467), .dinb(n3435), .dout(n3468));
  jand g3414(.dina(n1110), .dinb(n389), .dout(n3469));
  jand g3415(.dina(n3469), .dinb(n418), .dout(n3470));
  jand g3416(.dina(n3470), .dinb(n1035), .dout(n3471));
  jand g3417(.dina(n2717), .dinb(n505), .dout(n3472));
  jand g3418(.dina(n3472), .dinb(n207), .dout(n3473));
  jand g3419(.dina(n3473), .dinb(n3471), .dout(n3474));
  jand g3420(.dina(n347), .dinb(n265), .dout(n3475));
  jand g3421(.dina(n3475), .dinb(n222), .dout(n3476));
  jand g3422(.dina(n462), .dinb(n434), .dout(n3477));
  jand g3423(.dina(n3477), .dinb(n120), .dout(n3478));
  jand g3424(.dina(n3478), .dinb(n307), .dout(n3479));
  jand g3425(.dina(n3479), .dinb(n3476), .dout(n3480));
  jand g3426(.dina(n3480), .dinb(n3474), .dout(n3481));
  jand g3427(.dina(n3481), .dinb(n1032), .dout(n3482));
  jand g3428(.dina(n2394), .dinb(n190), .dout(n3483));
  jand g3429(.dina(n3483), .dinb(n1009), .dout(n3484));
  jand g3430(.dina(n387), .dinb(n137), .dout(n3485));
  jand g3431(.dina(n3485), .dinb(n353), .dout(n3486));
  jand g3432(.dina(n3486), .dinb(n3484), .dout(n3487));
  jand g3433(.dina(n290), .dinb(n215), .dout(n3488));
  jand g3434(.dina(n313), .dinb(n142), .dout(n3489));
  jand g3435(.dina(n3489), .dinb(n236), .dout(n3490));
  jand g3436(.dina(n3490), .dinb(n3488), .dout(n3491));
  jand g3437(.dina(n3491), .dinb(n435), .dout(n3492));
  jand g3438(.dina(n3492), .dinb(n3487), .dout(n3493));
  jand g3439(.dina(n3493), .dinb(n3482), .dout(n3494));
  jxor g3440(.dina(n3494), .dinb(n3468), .dout(n3495));
  jand g3441(.dina(n3494), .dinb(n3468), .dout(n3496));
  jnot g3442(.din(n1185), .dout(n3497));
  jand g3443(.dina(n2127), .dinb(n3497), .dout(n3498));
  jand g3444(.dina(n561), .dinb(n344), .dout(n3499));
  jand g3445(.dina(n3499), .dinb(n1074), .dout(n3500));
  jand g3446(.dina(n3500), .dinb(n3498), .dout(n3501));
  jand g3447(.dina(n3501), .dinb(n2968), .dout(n3502));
  jand g3448(.dina(n897), .dinb(n197), .dout(n3503));
  jand g3449(.dina(n3503), .dinb(n267), .dout(n3504));
  jand g3450(.dina(n3504), .dinb(n248), .dout(n3505));
  jand g3451(.dina(n3505), .dinb(n2134), .dout(n3506));
  jand g3452(.dina(n3506), .dinb(n3502), .dout(n3507));
  jand g3453(.dina(n3507), .dinb(n443), .dout(n3508));
  jand g3454(.dina(n3508), .dinb(n1456), .dout(n3509));
  jxor g3455(.dina(n3509), .dinb(n3496), .dout(n3510));
  jor  g3456(.dina(n3510), .dinb(n3495), .dout(n3511));
  jor  g3457(.dina(n3495), .dinb(n3441), .dout(n3512));
  jxor g3458(.dina(n3440), .dinb(n3435), .dout(n3513));
  jand g3459(.dina(n3513), .dinb(n3415), .dout(n3514));
  jnot g3460(.din(n3514), .dout(n3515));
  jxor g3461(.dina(n3441), .dinb(n3415), .dout(n3516));
  jor  g3462(.dina(n3516), .dinb(n3420), .dout(n3517));
  jand g3463(.dina(n3517), .dinb(n3515), .dout(n3518));
  jnot g3464(.din(n3494), .dout(n3519));
  jxor g3465(.dina(n3519), .dinb(n3468), .dout(n3520));
  jand g3466(.dina(n3520), .dinb(n3513), .dout(n3521));
  jor  g3467(.dina(n3519), .dinb(n3513), .dout(n3522));
  jnot g3468(.din(n3522), .dout(n3523));
  jor  g3469(.dina(n3523), .dinb(n3521), .dout(n3524));
  jor  g3470(.dina(n3524), .dinb(n3518), .dout(n3525));
  jand g3471(.dina(n3525), .dinb(n3512), .dout(n3526));
  jand g3472(.dina(n3509), .dinb(n3495), .dout(n3527));
  jnot g3473(.din(n3527), .dout(n3528));
  jand g3474(.dina(n3528), .dinb(n3511), .dout(n3529));
  jnot g3475(.din(n3529), .dout(n3530));
  jor  g3476(.dina(n3530), .dinb(n3526), .dout(n3531));
  jand g3477(.dina(n3531), .dinb(n3511), .dout(n3532));
  jand g3478(.dina(n1470), .dinb(n513), .dout(n3533));
  jand g3479(.dina(n3533), .dinb(n459), .dout(n3534));
  jand g3480(.dina(n871), .dinb(n468), .dout(n3535));
  jand g3481(.dina(n1460), .dinb(n539), .dout(n3536));
  jand g3482(.dina(n569), .dinb(n157), .dout(n3537));
  jand g3483(.dina(n3537), .dinb(n169), .dout(n3538));
  jand g3484(.dina(n3538), .dinb(n3536), .dout(n3539));
  jand g3485(.dina(n3539), .dinb(n3535), .dout(n3540));
  jand g3486(.dina(n3540), .dinb(n443), .dout(n3541));
  jand g3487(.dina(n3541), .dinb(n1444), .dout(n3542));
  jand g3488(.dina(n3542), .dinb(n3534), .dout(n3543));
  jand g3489(.dina(n3543), .dinb(n3510), .dout(n3544));
  jnot g3490(.din(n3544), .dout(n3545));
  jand g3491(.dina(n3509), .dinb(n3496), .dout(n3546));
  jxor g3492(.dina(n3543), .dinb(n3546), .dout(n3547));
  jor  g3493(.dina(n3547), .dinb(n3510), .dout(n3548));
  jand g3494(.dina(n3548), .dinb(n3545), .dout(n3549));
  jxor g3495(.dina(n3549), .dinb(n3532), .dout(n3550));
  jor  g3496(.dina(n3550), .dinb(n3461), .dout(n3551));
  jor  g3497(.dina(n50), .dinb(n3021), .dout(n3552));
  jor  g3498(.dina(n3552), .dinb(n3495), .dout(n3553));
  jor  g3499(.dina(n3459), .dinb(n3456), .dout(n3554));
  jor  g3500(.dina(n3554), .dinb(n3547), .dout(n3555));
  jand g3501(.dina(n3555), .dinb(n3553), .dout(n3556));
  jand g3502(.dina(a1 ), .dinb(n3456), .dout(n3557));
  jnot g3503(.din(n3557), .dout(n3558));
  jor  g3504(.dina(n3558), .dinb(n3510), .dout(n3559));
  jand g3505(.dina(n3559), .dinb(n3556), .dout(n3560));
  jand g3506(.dina(n3560), .dinb(n3551), .dout(n3561));
  jxor g3507(.dina(n3561), .dinb(n3455), .dout(n3562));
  jor  g3508(.dina(n3562), .dinb(n3454), .dout(n3563));
  jnot g3509(.din(n3563), .dout(n3564));
  jxor g3510(.dina(n3361), .dinb(n3360), .dout(n3565));
  jxor g3511(.dina(n3529), .dinb(n3526), .dout(n3566));
  jor  g3512(.dina(n3566), .dinb(n3461), .dout(n3567));
  jor  g3513(.dina(n3554), .dinb(n3510), .dout(n3568));
  jor  g3514(.dina(n3558), .dinb(n3495), .dout(n3569));
  jor  g3515(.dina(n3552), .dinb(n3441), .dout(n3570));
  jand g3516(.dina(n3570), .dinb(n3569), .dout(n3571));
  jand g3517(.dina(n3571), .dinb(n3568), .dout(n3572));
  jand g3518(.dina(n3572), .dinb(n3567), .dout(n3573));
  jxor g3519(.dina(n3573), .dinb(n3023), .dout(n3574));
  jand g3520(.dina(n3574), .dinb(n3565), .dout(n3575));
  jxor g3521(.dina(n3574), .dinb(n3565), .dout(n3576));
  jxor g3522(.dina(n3358), .dinb(n3357), .dout(n3577));
  jand g3523(.dina(n3522), .dinb(n3512), .dout(n3578));
  jxor g3524(.dina(n3578), .dinb(n3518), .dout(n3579));
  jor  g3525(.dina(n3579), .dinb(n3461), .dout(n3580));
  jor  g3526(.dina(n3554), .dinb(n3495), .dout(n3581));
  jor  g3527(.dina(n3558), .dinb(n3441), .dout(n3582));
  jor  g3528(.dina(n3552), .dinb(n3203), .dout(n3583));
  jand g3529(.dina(n3583), .dinb(n3582), .dout(n3584));
  jand g3530(.dina(n3584), .dinb(n3581), .dout(n3585));
  jand g3531(.dina(n3585), .dinb(n3580), .dout(n3586));
  jxor g3532(.dina(n3586), .dinb(n3023), .dout(n3587));
  jand g3533(.dina(n3587), .dinb(n3577), .dout(n3588));
  jor  g3534(.dina(n3587), .dinb(n3577), .dout(n3589));
  jxor g3535(.dina(n3355), .dinb(n3354), .dout(n3590));
  jor  g3536(.dina(n3461), .dinb(n3443), .dout(n3591));
  jor  g3537(.dina(n3558), .dinb(n3203), .dout(n3592));
  jor  g3538(.dina(n3554), .dinb(n3441), .dout(n3593));
  jor  g3539(.dina(n3552), .dinb(n3166), .dout(n3594));
  jand g3540(.dina(n3594), .dinb(n3593), .dout(n3595));
  jand g3541(.dina(n3595), .dinb(n3592), .dout(n3596));
  jand g3542(.dina(n3596), .dinb(n3591), .dout(n3597));
  jxor g3543(.dina(n3597), .dinb(n3023), .dout(n3598));
  jor  g3544(.dina(n3598), .dinb(n3590), .dout(n3599));
  jand g3545(.dina(n3598), .dinb(n3590), .dout(n3600));
  jxor g3546(.dina(n3352), .dinb(n3351), .dout(n3601));
  jor  g3547(.dina(n3461), .dinb(n3205), .dout(n3602));
  jor  g3548(.dina(n3554), .dinb(n3203), .dout(n3603));
  jor  g3549(.dina(n3558), .dinb(n3166), .dout(n3604));
  jor  g3550(.dina(n3552), .dinb(n3216), .dout(n3605));
  jand g3551(.dina(n3605), .dinb(n3604), .dout(n3606));
  jand g3552(.dina(n3606), .dinb(n3603), .dout(n3607));
  jand g3553(.dina(n3607), .dinb(n3602), .dout(n3608));
  jxor g3554(.dina(n3608), .dinb(n3023), .dout(n3609));
  jor  g3555(.dina(n3609), .dinb(n3601), .dout(n3610));
  jand g3556(.dina(n3609), .dinb(n3601), .dout(n3611));
  jxor g3557(.dina(n3349), .dinb(n3348), .dout(n3612));
  jor  g3558(.dina(n3461), .dinb(n3229), .dout(n3613));
  jor  g3559(.dina(n3554), .dinb(n3166), .dout(n3614));
  jor  g3560(.dina(n3558), .dinb(n3216), .dout(n3615));
  jand g3561(.dina(n3615), .dinb(n3614), .dout(n3616));
  jor  g3562(.dina(n3552), .dinb(n3008), .dout(n3617));
  jand g3563(.dina(n3617), .dinb(n3616), .dout(n3618));
  jand g3564(.dina(n3618), .dinb(n3613), .dout(n3619));
  jxor g3565(.dina(n3619), .dinb(n3023), .dout(n3620));
  jor  g3566(.dina(n3620), .dinb(n3612), .dout(n3621));
  jand g3567(.dina(n3620), .dinb(n3612), .dout(n3622));
  jxor g3568(.dina(n3346), .dinb(n3345), .dout(n3623));
  jor  g3569(.dina(n3461), .dinb(n3242), .dout(n3624));
  jor  g3570(.dina(n3554), .dinb(n3216), .dout(n3625));
  jor  g3571(.dina(n3558), .dinb(n3008), .dout(n3626));
  jor  g3572(.dina(n3552), .dinb(n2800), .dout(n3627));
  jand g3573(.dina(n3627), .dinb(n3626), .dout(n3628));
  jand g3574(.dina(n3628), .dinb(n3625), .dout(n3629));
  jand g3575(.dina(n3629), .dinb(n3624), .dout(n3630));
  jxor g3576(.dina(n3630), .dinb(n3023), .dout(n3631));
  jor  g3577(.dina(n3631), .dinb(n3623), .dout(n3632));
  jand g3578(.dina(n3631), .dinb(n3623), .dout(n3633));
  jxor g3579(.dina(n3343), .dinb(n3341), .dout(n3634));
  jor  g3580(.dina(n3461), .dinb(n3010), .dout(n3635));
  jor  g3581(.dina(n3554), .dinb(n3008), .dout(n3636));
  jor  g3582(.dina(n3558), .dinb(n2800), .dout(n3637));
  jand g3583(.dina(n3637), .dinb(n3636), .dout(n3638));
  jor  g3584(.dina(n3552), .dinb(n2707), .dout(n3639));
  jand g3585(.dina(n3639), .dinb(n3638), .dout(n3640));
  jand g3586(.dina(n3640), .dinb(n3635), .dout(n3641));
  jxor g3587(.dina(n3641), .dinb(n3023), .dout(n3642));
  jor  g3588(.dina(n3642), .dinb(n3634), .dout(n3643));
  jand g3589(.dina(n3642), .dinb(n3634), .dout(n3644));
  jxor g3590(.dina(n3338), .dinb(n3337), .dout(n3645));
  jor  g3591(.dina(n3461), .dinb(n2802), .dout(n3646));
  jor  g3592(.dina(n3554), .dinb(n2800), .dout(n3647));
  jor  g3593(.dina(n3558), .dinb(n2707), .dout(n3648));
  jor  g3594(.dina(n3552), .dinb(n2813), .dout(n3649));
  jand g3595(.dina(n3649), .dinb(n3648), .dout(n3650));
  jand g3596(.dina(n3650), .dinb(n3647), .dout(n3651));
  jand g3597(.dina(n3651), .dinb(n3646), .dout(n3652));
  jxor g3598(.dina(n3652), .dinb(n3023), .dout(n3653));
  jor  g3599(.dina(n3653), .dinb(n3645), .dout(n3654));
  jand g3600(.dina(n3653), .dinb(n3645), .dout(n3655));
  jxor g3601(.dina(n3334), .dinb(n3326), .dout(n3656));
  jor  g3602(.dina(n3461), .dinb(n2825), .dout(n3657));
  jor  g3603(.dina(n3554), .dinb(n2707), .dout(n3658));
  jor  g3604(.dina(n3558), .dinb(n2813), .dout(n3659));
  jand g3605(.dina(n3659), .dinb(n3658), .dout(n3660));
  jor  g3606(.dina(n3552), .dinb(n2471), .dout(n3661));
  jand g3607(.dina(n3661), .dinb(n3660), .dout(n3662));
  jand g3608(.dina(n3662), .dinb(n3657), .dout(n3663));
  jxor g3609(.dina(n3663), .dinb(n3023), .dout(n3664));
  jor  g3610(.dina(n3664), .dinb(n3656), .dout(n3665));
  jand g3611(.dina(n3557), .dinb(n2094), .dout(n3666));
  jor  g3612(.dina(n3666), .dinb(n3023), .dout(n3667));
  jor  g3613(.dina(n3667), .dinb(n1956), .dout(n3668));
  jnot g3614(.din(n3668), .dout(n3669));
  jand g3615(.dina(n2256), .dinb(n2116), .dout(n3670));
  jor  g3616(.dina(n3670), .dinb(n3554), .dout(n3671));
  jand g3617(.dina(n2256), .dinb(n2095), .dout(n3672));
  jor  g3618(.dina(n3672), .dinb(n3461), .dout(n3673));
  jand g3619(.dina(n3673), .dinb(n3671), .dout(n3674));
  jand g3620(.dina(n3674), .dinb(n3669), .dout(n3675));
  jor  g3621(.dina(n3675), .dinb(n3312), .dout(n3676));
  jor  g3622(.dina(n2236), .dinb(n1956), .dout(n3677));
  jand g3623(.dina(n3677), .dinb(n2094), .dout(n3678));
  jxor g3624(.dina(n2352), .dinb(n3678), .dout(n3679));
  jand g3625(.dina(n3460), .dinb(n3679), .dout(n3680));
  jand g3626(.dina(n3557), .dinb(n2236), .dout(n3681));
  jnot g3627(.din(n3554), .dout(n3682));
  jand g3628(.dina(n3682), .dinb(n2690), .dout(n3683));
  jor  g3629(.dina(n3683), .dinb(n3681), .dout(n3684));
  jor  g3630(.dina(n3684), .dinb(n3680), .dout(n3685));
  jnot g3631(.din(n3552), .dout(n3686));
  jand g3632(.dina(n3686), .dinb(n2094), .dout(n3687));
  jor  g3633(.dina(n3687), .dinb(n3023), .dout(n3688));
  jnot g3634(.din(n3688), .dout(n3689));
  jor  g3635(.dina(n3689), .dinb(n3685), .dout(n3690));
  jor  g3636(.dina(n3461), .dinb(n2353), .dout(n3691));
  jnot g3637(.din(n3681), .dout(n3692));
  jor  g3638(.dina(n3554), .dinb(n2351), .dout(n3693));
  jand g3639(.dina(n3693), .dinb(n3692), .dout(n3694));
  jand g3640(.dina(n3694), .dinb(n3691), .dout(n3695));
  jor  g3641(.dina(n3695), .dinb(n3023), .dout(n3696));
  jand g3642(.dina(n3696), .dinb(n3690), .dout(n3697));
  jand g3643(.dina(n3697), .dinb(n3676), .dout(n3698));
  jand g3644(.dina(n3312), .dinb(n1154), .dout(n3699));
  jxor g3645(.dina(n3699), .dinb(n3311), .dout(n3700));
  jnot g3646(.din(n3700), .dout(n3701));
  jand g3647(.dina(n3701), .dinb(n3698), .dout(n3702));
  jor  g3648(.dina(n3701), .dinb(n3698), .dout(n3703));
  jor  g3649(.dina(n3461), .dinb(n2473), .dout(n3704));
  jand g3650(.dina(n3557), .dinb(n2690), .dout(n3705));
  jnot g3651(.din(n3705), .dout(n3706));
  jor  g3652(.dina(n3554), .dinb(n2471), .dout(n3707));
  jand g3653(.dina(n3707), .dinb(n3706), .dout(n3708));
  jand g3654(.dina(n3708), .dinb(n3704), .dout(n3709));
  jor  g3655(.dina(n3709), .dinb(n3023), .dout(n3710));
  jand g3656(.dina(n2690), .dinb(n2236), .dout(n3711));
  jand g3657(.dina(n2352), .dinb(n3678), .dout(n3712));
  jor  g3658(.dina(n3712), .dinb(n3711), .dout(n3713));
  jxor g3659(.dina(n2472), .dinb(n3713), .dout(n3714));
  jand g3660(.dina(n3460), .dinb(n3714), .dout(n3715));
  jand g3661(.dina(n3682), .dinb(n2687), .dout(n3716));
  jor  g3662(.dina(n3716), .dinb(n3705), .dout(n3717));
  jor  g3663(.dina(n3717), .dinb(n3715), .dout(n3718));
  jand g3664(.dina(n3686), .dinb(n2236), .dout(n3719));
  jor  g3665(.dina(n3719), .dinb(n3023), .dout(n3720));
  jnot g3666(.din(n3720), .dout(n3721));
  jor  g3667(.dina(n3721), .dinb(n3718), .dout(n3722));
  jand g3668(.dina(n3722), .dinb(n3710), .dout(n3723));
  jand g3669(.dina(n3723), .dinb(n3703), .dout(n3724));
  jor  g3670(.dina(n3724), .dinb(n3702), .dout(n3725));
  jor  g3671(.dina(n3461), .dinb(n2836), .dout(n3726));
  jor  g3672(.dina(n3554), .dinb(n2813), .dout(n3727));
  jor  g3673(.dina(n3558), .dinb(n2471), .dout(n3728));
  jor  g3674(.dina(n3552), .dinb(n2351), .dout(n3729));
  jand g3675(.dina(n3729), .dinb(n3728), .dout(n3730));
  jand g3676(.dina(n3730), .dinb(n3727), .dout(n3731));
  jand g3677(.dina(n3731), .dinb(n3726), .dout(n3732));
  jxor g3678(.dina(n3732), .dinb(n3023), .dout(n3733));
  jor  g3679(.dina(n3733), .dinb(n3725), .dout(n3734));
  jand g3680(.dina(n3733), .dinb(n3725), .dout(n3735));
  jnot g3681(.din(n3315), .dout(n3736));
  jand g3682(.dina(n3736), .dinb(n1154), .dout(n3737));
  jxor g3683(.dina(n3737), .dinb(n3323), .dout(n3738));
  jnot g3684(.din(n3738), .dout(n3739));
  jor  g3685(.dina(n3739), .dinb(n3735), .dout(n3740));
  jand g3686(.dina(n3740), .dinb(n3734), .dout(n3741));
  jand g3687(.dina(n3664), .dinb(n3656), .dout(n3742));
  jor  g3688(.dina(n3742), .dinb(n3741), .dout(n3743));
  jand g3689(.dina(n3743), .dinb(n3665), .dout(n3744));
  jor  g3690(.dina(n3744), .dinb(n3655), .dout(n3745));
  jand g3691(.dina(n3745), .dinb(n3654), .dout(n3746));
  jor  g3692(.dina(n3746), .dinb(n3644), .dout(n3747));
  jand g3693(.dina(n3747), .dinb(n3643), .dout(n3748));
  jor  g3694(.dina(n3748), .dinb(n3633), .dout(n3749));
  jand g3695(.dina(n3749), .dinb(n3632), .dout(n3750));
  jor  g3696(.dina(n3750), .dinb(n3622), .dout(n3751));
  jand g3697(.dina(n3751), .dinb(n3621), .dout(n3752));
  jor  g3698(.dina(n3752), .dinb(n3611), .dout(n3753));
  jand g3699(.dina(n3753), .dinb(n3610), .dout(n3754));
  jor  g3700(.dina(n3754), .dinb(n3600), .dout(n3755));
  jand g3701(.dina(n3755), .dinb(n3599), .dout(n3756));
  jand g3702(.dina(n3756), .dinb(n3589), .dout(n3757));
  jor  g3703(.dina(n3757), .dinb(n3588), .dout(n3758));
  jand g3704(.dina(n3758), .dinb(n3576), .dout(n3759));
  jor  g3705(.dina(n3759), .dinb(n3575), .dout(n3760));
  jxor g3706(.dina(n3562), .dinb(n3454), .dout(n3761));
  jand g3707(.dina(n3761), .dinb(n3760), .dout(n3762));
  jor  g3708(.dina(n3762), .dinb(n3564), .dout(n3763));
  jand g3709(.dina(n3451), .dinb(n3409), .dout(n3764));
  jand g3710(.dina(n3452), .dinb(n3363), .dout(n3765));
  jor  g3711(.dina(n3765), .dinb(n3764), .dout(n3766));
  jor  g3712(.dina(n3407), .dinb(n3399), .dout(n3767));
  jnot g3713(.din(n3767), .dout(n3768));
  jand g3714(.dina(n3408), .dinb(n3368), .dout(n3769));
  jor  g3715(.dina(n3769), .dinb(n3768), .dout(n3770));
  jand g3716(.dina(n3396), .dinb(n3380), .dout(n3771));
  jand g3717(.dina(n3397), .dinb(n3371), .dout(n3772));
  jor  g3718(.dina(n3772), .dinb(n3771), .dout(n3773));
  jand g3719(.dina(n3382), .dinb(n3381), .dout(n3774));
  jnot g3720(.din(n3774), .dout(n3775));
  jand g3721(.dina(n3395), .dinb(n3775), .dout(n3779));
  jnot g3722(.din(n3779), .dout(n3780));
  jand g3723(.dina(n2484), .dinb(n3714), .dout(n3781));
  jand g3724(.dina(n2491), .dinb(n2687), .dout(n3782));
  jand g3725(.dina(n2488), .dinb(n2690), .dout(n3783));
  jand g3726(.dina(n2923), .dinb(n2236), .dout(n3784));
  jor  g3727(.dina(n3784), .dinb(n3783), .dout(n3785));
  jor  g3728(.dina(n3785), .dinb(n3782), .dout(n3786));
  jor  g3729(.dina(n3786), .dinb(n3781), .dout(n3787));
  jor  g3730(.dina(n2094), .dinb(n2051), .dout(n3788));
  jxor g3731(.dina(n3788), .dinb(n3787), .dout(n3789));
  jxor g3732(.dina(n3789), .dinb(n3780), .dout(n3790));
  jor  g3733(.dina(n2802), .dinb(n2252), .dout(n3791));
  jor  g3734(.dina(n2800), .dinb(n2355), .dout(n3792));
  jor  g3735(.dina(n2707), .dinb(n2359), .dout(n3793));
  jor  g3736(.dina(n2813), .dinb(n2357), .dout(n3794));
  jand g3737(.dina(n3794), .dinb(n3793), .dout(n3795));
  jand g3738(.dina(n3795), .dinb(n3792), .dout(n3796));
  jand g3739(.dina(n3796), .dinb(n3791), .dout(n3797));
  jxor g3740(.dina(n3797), .dinb(n1480), .dout(n3798));
  jxor g3741(.dina(n3798), .dinb(n3790), .dout(n3799));
  jxor g3742(.dina(n3799), .dinb(n3773), .dout(n3800));
  jnot g3743(.din(n3800), .dout(n3801));
  jor  g3744(.dina(n3229), .dinb(n2506), .dout(n3802));
  jor  g3745(.dina(n3166), .dinb(n2810), .dout(n3803));
  jor  g3746(.dina(n3216), .dinb(n2807), .dout(n3804));
  jand g3747(.dina(n3804), .dinb(n3803), .dout(n3805));
  jor  g3748(.dina(n3008), .dinb(n2816), .dout(n3806));
  jand g3749(.dina(n3806), .dinb(n3805), .dout(n3807));
  jand g3750(.dina(n3807), .dinb(n3802), .dout(n3808));
  jxor g3751(.dina(n3808), .dinb(n1257), .dout(n3809));
  jxor g3752(.dina(n3809), .dinb(n3801), .dout(n3810));
  jxor g3753(.dina(n3810), .dinb(n3770), .dout(n3811));
  jor  g3754(.dina(n3579), .dinb(n3029), .dout(n3812));
  jor  g3755(.dina(n3495), .dinb(n3213), .dout(n3813));
  jor  g3756(.dina(n3441), .dinb(n3210), .dout(n3814));
  jor  g3757(.dina(n3219), .dinb(n3203), .dout(n3815));
  jand g3758(.dina(n3815), .dinb(n3814), .dout(n3816));
  jand g3759(.dina(n3816), .dinb(n3813), .dout(n3817));
  jand g3760(.dina(n3817), .dinb(n3812), .dout(n3818));
  jxor g3761(.dina(n3818), .dinb(n1156), .dout(n3819));
  jxor g3762(.dina(n3819), .dinb(n3811), .dout(n3820));
  jxor g3763(.dina(n3820), .dinb(n3766), .dout(n3821));
  jnot g3764(.din(n3549), .dout(n3822));
  jor  g3765(.dina(n3822), .dinb(n3532), .dout(n3823));
  jand g3766(.dina(n3823), .dinb(n3548), .dout(n3824));
  jnot g3767(.din(n3547), .dout(n3825));
  jand g3768(.dina(n514), .dinb(n332), .dout(n3826));
  jand g3769(.dina(n1467), .dinb(n443), .dout(n3827));
  jand g3770(.dina(n3827), .dinb(n3826), .dout(n3828));
  jand g3771(.dina(n232), .dinb(n213), .dout(n3829));
  jand g3772(.dina(n3829), .dinb(n315), .dout(n3830));
  jand g3773(.dina(n3830), .dinb(n500), .dout(n3831));
  jand g3774(.dina(n3831), .dinb(n1447), .dout(n3832));
  jand g3775(.dina(n3832), .dinb(n3828), .dout(n3833));
  jnot g3776(.din(n3833), .dout(n3834));
  jor  g3777(.dina(n3834), .dinb(n3825), .dout(n3835));
  jand g3778(.dina(n3543), .dinb(n3546), .dout(n3836));
  jxor g3779(.dina(n3833), .dinb(n3836), .dout(n3837));
  jnot g3780(.din(n3837), .dout(n3838));
  jand g3781(.dina(n3838), .dinb(n3825), .dout(n3839));
  jnot g3782(.din(n3839), .dout(n3840));
  jand g3783(.dina(n3840), .dinb(n3835), .dout(n3841));
  jxor g3784(.dina(n3841), .dinb(n3824), .dout(n3842));
  jor  g3785(.dina(n3842), .dinb(n3461), .dout(n3843));
  jor  g3786(.dina(n3837), .dinb(n3554), .dout(n3844));
  jor  g3787(.dina(n3558), .dinb(n3547), .dout(n3845));
  jor  g3788(.dina(n3552), .dinb(n3510), .dout(n3846));
  jand g3789(.dina(n3846), .dinb(n3845), .dout(n3847));
  jand g3790(.dina(n3847), .dinb(n3844), .dout(n3848));
  jand g3791(.dina(n3848), .dinb(n3843), .dout(n3849));
  jxor g3792(.dina(n3849), .dinb(n3023), .dout(n3850));
  jxor g3793(.dina(n3850), .dinb(n3821), .dout(n3851));
  jxor g3794(.dina(n3851), .dinb(n3763), .dout(n3852));
  jand g3795(.dina(n3852), .dinb(n325), .dout(n3853));
  jxor g3796(.dina(n3852), .dinb(n325), .dout(n3854));
  jand g3797(.dina(n344), .dinb(n152), .dout(n3855));
  jand g3798(.dina(n3855), .dinb(n884), .dout(n3856));
  jand g3799(.dina(n587), .dinb(n434), .dout(n3857));
  jand g3800(.dina(n3857), .dinb(n446), .dout(n3858));
  jand g3801(.dina(n3858), .dinb(n3856), .dout(n3859));
  jand g3802(.dina(n3859), .dinb(n1965), .dout(n3860));
  jand g3803(.dina(n383), .dinb(n333), .dout(n3861));
  jand g3804(.dina(n3861), .dinb(n241), .dout(n3862));
  jand g3805(.dina(n3862), .dinb(n497), .dout(n3863));
  jand g3806(.dina(n438), .dinb(n102), .dout(n3864));
  jand g3807(.dina(n3864), .dinb(n600), .dout(n3865));
  jand g3808(.dina(n3865), .dinb(n2377), .dout(n3866));
  jand g3809(.dina(n3866), .dinb(n3863), .dout(n3867));
  jand g3810(.dina(n3867), .dinb(n856), .dout(n3868));
  jand g3811(.dina(n1087), .dinb(n339), .dout(n3869));
  jand g3812(.dina(n3869), .dinb(n361), .dout(n3870));
  jand g3813(.dina(n3870), .dinb(n3868), .dout(n3871));
  jand g3814(.dina(n1072), .dinb(n166), .dout(n3872));
  jand g3815(.dina(n488), .dinb(n207), .dout(n3873));
  jand g3816(.dina(n3873), .dinb(n1080), .dout(n3874));
  jand g3817(.dina(n3874), .dinb(n133), .dout(n3875));
  jand g3818(.dina(n3875), .dinb(n3872), .dout(n3876));
  jand g3819(.dina(n510), .dinb(n384), .dout(n3877));
  jand g3820(.dina(n3877), .dinb(n161), .dout(n3878));
  jand g3821(.dina(n3878), .dinb(n120), .dout(n3879));
  jand g3822(.dina(n3879), .dinb(n3489), .dout(n3880));
  jand g3823(.dina(n3880), .dinb(n3876), .dout(n3881));
  jand g3824(.dina(n387), .dinb(n331), .dout(n3882));
  jand g3825(.dina(n3882), .dinb(n124), .dout(n3883));
  jand g3826(.dina(n3883), .dinb(n94), .dout(n3884));
  jand g3827(.dina(n3884), .dinb(n3881), .dout(n3885));
  jand g3828(.dina(n3885), .dinb(n3871), .dout(n3886));
  jand g3829(.dina(n3886), .dinb(n3860), .dout(n3887));
  jand g3830(.dina(n2613), .dinb(n1332), .dout(n3888));
  jand g3831(.dina(n1460), .dinb(n173), .dout(n3889));
  jand g3832(.dina(n3889), .dinb(n2142), .dout(n3890));
  jand g3833(.dina(n3890), .dinb(n435), .dout(n3891));
  jand g3834(.dina(n3891), .dinb(n3888), .dout(n3892));
  jand g3835(.dina(n152), .dinb(n136), .dout(n3893));
  jand g3836(.dina(n3893), .dinb(n3185), .dout(n3894));
  jand g3837(.dina(n3894), .dinb(n1078), .dout(n3895));
  jand g3838(.dina(n252), .dinb(n142), .dout(n3896));
  jand g3839(.dina(n535), .dinb(n283), .dout(n3897));
  jand g3840(.dina(n347), .dinb(n232), .dout(n3898));
  jand g3841(.dina(n3898), .dinb(n3897), .dout(n3899));
  jand g3842(.dina(n3899), .dinb(n3896), .dout(n3900));
  jand g3843(.dina(n463), .dinb(n382), .dout(n3901));
  jand g3844(.dina(n3901), .dinb(n1366), .dout(n3902));
  jand g3845(.dina(n3902), .dinb(n1961), .dout(n3903));
  jand g3846(.dina(n3903), .dinb(n2155), .dout(n3904));
  jand g3847(.dina(n3904), .dinb(n3900), .dout(n3905));
  jand g3848(.dina(n3905), .dinb(n3895), .dout(n3906));
  jand g3849(.dina(n3906), .dinb(n3892), .dout(n3907));
  jand g3850(.dina(n3907), .dinb(n2409), .dout(n3908));
  jnot g3851(.din(n3908), .dout(n3909));
  jnot g3852(.din(n3576), .dout(n3910));
  jnot g3853(.din(n3588), .dout(n3911));
  jnot g3854(.din(n3589), .dout(n3912));
  jnot g3855(.din(n3599), .dout(n3913));
  jnot g3856(.din(n3600), .dout(n3914));
  jnot g3857(.din(n3610), .dout(n3915));
  jnot g3858(.din(n3611), .dout(n3916));
  jnot g3859(.din(n3621), .dout(n3917));
  jnot g3860(.din(n3622), .dout(n3918));
  jnot g3861(.din(n3632), .dout(n3919));
  jnot g3862(.din(n3633), .dout(n3920));
  jnot g3863(.din(n3643), .dout(n3921));
  jnot g3864(.din(n3644), .dout(n3922));
  jnot g3865(.din(n3654), .dout(n3923));
  jnot g3866(.din(n3655), .dout(n3924));
  jnot g3867(.din(n3665), .dout(n3925));
  jnot g3868(.din(n3734), .dout(n3926));
  jnot g3869(.din(n3702), .dout(n3927));
  jnot g3870(.din(n3676), .dout(n3928));
  jand g3871(.dina(n3688), .dinb(n3695), .dout(n3929));
  jand g3872(.dina(n3685), .dinb(n3455), .dout(n3930));
  jor  g3873(.dina(n3930), .dinb(n3929), .dout(n3931));
  jor  g3874(.dina(n3931), .dinb(n3928), .dout(n3932));
  jand g3875(.dina(n3700), .dinb(n3932), .dout(n3933));
  jand g3876(.dina(n3718), .dinb(n3455), .dout(n3934));
  jand g3877(.dina(n3720), .dinb(n3709), .dout(n3935));
  jor  g3878(.dina(n3935), .dinb(n3934), .dout(n3936));
  jor  g3879(.dina(n3936), .dinb(n3933), .dout(n3937));
  jand g3880(.dina(n3937), .dinb(n3927), .dout(n3938));
  jnot g3881(.din(n3733), .dout(n3939));
  jor  g3882(.dina(n3939), .dinb(n3938), .dout(n3940));
  jand g3883(.dina(n3738), .dinb(n3940), .dout(n3941));
  jor  g3884(.dina(n3941), .dinb(n3926), .dout(n3942));
  jnot g3885(.din(n3742), .dout(n3943));
  jand g3886(.dina(n3943), .dinb(n3942), .dout(n3944));
  jor  g3887(.dina(n3944), .dinb(n3925), .dout(n3945));
  jand g3888(.dina(n3945), .dinb(n3924), .dout(n3946));
  jor  g3889(.dina(n3946), .dinb(n3923), .dout(n3947));
  jand g3890(.dina(n3947), .dinb(n3922), .dout(n3948));
  jor  g3891(.dina(n3948), .dinb(n3921), .dout(n3949));
  jand g3892(.dina(n3949), .dinb(n3920), .dout(n3950));
  jor  g3893(.dina(n3950), .dinb(n3919), .dout(n3951));
  jand g3894(.dina(n3951), .dinb(n3918), .dout(n3952));
  jor  g3895(.dina(n3952), .dinb(n3917), .dout(n3953));
  jand g3896(.dina(n3953), .dinb(n3916), .dout(n3954));
  jor  g3897(.dina(n3954), .dinb(n3915), .dout(n3955));
  jand g3898(.dina(n3955), .dinb(n3914), .dout(n3956));
  jor  g3899(.dina(n3956), .dinb(n3913), .dout(n3957));
  jor  g3900(.dina(n3957), .dinb(n3912), .dout(n3958));
  jand g3901(.dina(n3958), .dinb(n3911), .dout(n3959));
  jxor g3902(.dina(n3959), .dinb(n3910), .dout(n3960));
  jand g3903(.dina(n3960), .dinb(n3909), .dout(n3961));
  jnot g3904(.din(n3961), .dout(n3962));
  jand g3905(.dina(n3962), .dinb(n3887), .dout(n3963));
  jnot g3906(.din(n3963), .dout(n3964));
  jnot g3907(.din(n3887), .dout(n3965));
  jand g3908(.dina(n3961), .dinb(n3965), .dout(n3966));
  jxor g3909(.dina(n3761), .dinb(n3760), .dout(n3967));
  jor  g3910(.dina(n3967), .dinb(n3966), .dout(n3968));
  jand g3911(.dina(n3968), .dinb(n3964), .dout(n3969));
  jand g3912(.dina(n3969), .dinb(n3854), .dout(n3970));
  jor  g3913(.dina(n3970), .dinb(n3853), .dout(n3971));
  jand g3914(.dina(n3850), .dinb(n3821), .dout(n3972));
  jnot g3915(.din(n3972), .dout(n3973));
  jnot g3916(.din(n3575), .dout(n3974));
  jor  g3917(.dina(n3959), .dinb(n3910), .dout(n3975));
  jand g3918(.dina(n3975), .dinb(n3974), .dout(n3976));
  jnot g3919(.din(n3761), .dout(n3977));
  jor  g3920(.dina(n3977), .dinb(n3976), .dout(n3978));
  jand g3921(.dina(n3978), .dinb(n3563), .dout(n3979));
  jnot g3922(.din(n3851), .dout(n3980));
  jor  g3923(.dina(n3980), .dinb(n3979), .dout(n3981));
  jand g3924(.dina(n3981), .dinb(n3973), .dout(n3982));
  jand g3925(.dina(n3819), .dinb(n3811), .dout(n3983));
  jand g3926(.dina(n3820), .dinb(n3766), .dout(n3984));
  jor  g3927(.dina(n3984), .dinb(n3983), .dout(n3985));
  jor  g3928(.dina(n3809), .dinb(n3801), .dout(n3986));
  jnot g3929(.din(n3986), .dout(n3987));
  jand g3930(.dina(n3810), .dinb(n3770), .dout(n3988));
  jor  g3931(.dina(n3988), .dinb(n3987), .dout(n3989));
  jand g3932(.dina(n3798), .dinb(n3790), .dout(n3990));
  jand g3933(.dina(n3799), .dinb(n3773), .dout(n3991));
  jor  g3934(.dina(n3991), .dinb(n3990), .dout(n3992));
  jor  g3935(.dina(n3789), .dinb(n3780), .dout(n3993));
  jnot g3936(.din(n3787), .dout(n3994));
  jand g3937(.dina(n3994), .dinb(n1438), .dout(n3995));
  jand g3938(.dina(n3995), .dinb(n2094), .dout(n3996));
  jnot g3939(.din(n3996), .dout(n3997));
  jand g3940(.dina(n3997), .dinb(n3993), .dout(n3998));
  jor  g3941(.dina(n2836), .dinb(n3384), .dout(n3999));
  jand g3942(.dina(n2684), .dinb(n2491), .dout(n4000));
  jand g3943(.dina(n2488), .dinb(n2687), .dout(n4001));
  jand g3944(.dina(n2923), .dinb(n2690), .dout(n4002));
  jor  g3945(.dina(n4002), .dinb(n4001), .dout(n4003));
  jor  g3946(.dina(n4003), .dinb(n4000), .dout(n4004));
  jnot g3947(.din(n4004), .dout(n4005));
  jand g3948(.dina(n4005), .dinb(n3999), .dout(n4006));
  jand g3949(.dina(n2256), .dinb(n1438), .dout(n4007));
  jxor g3950(.dina(n4007), .dinb(n4006), .dout(n4008));
  jxor g3951(.dina(n4008), .dinb(n3998), .dout(n4009));
  jor  g3952(.dina(n3010), .dinb(n2252), .dout(n4010));
  jor  g3953(.dina(n2800), .dinb(n2359), .dout(n4011));
  jor  g3954(.dina(n3008), .dinb(n2355), .dout(n4012));
  jor  g3955(.dina(n2707), .dinb(n2357), .dout(n4013));
  jand g3956(.dina(n4013), .dinb(n4012), .dout(n4014));
  jand g3957(.dina(n4014), .dinb(n4011), .dout(n4015));
  jand g3958(.dina(n4015), .dinb(n4010), .dout(n4016));
  jxor g3959(.dina(n4016), .dinb(n1480), .dout(n4017));
  jxor g3960(.dina(n4017), .dinb(n4009), .dout(n4018));
  jxor g3961(.dina(n4018), .dinb(n3992), .dout(n4019));
  jnot g3962(.din(n4019), .dout(n4020));
  jor  g3963(.dina(n3205), .dinb(n2506), .dout(n4021));
  jor  g3964(.dina(n3166), .dinb(n2807), .dout(n4022));
  jor  g3965(.dina(n3203), .dinb(n2810), .dout(n4023));
  jand g3966(.dina(n4023), .dinb(n4022), .dout(n4024));
  jor  g3967(.dina(n3216), .dinb(n2816), .dout(n4025));
  jand g3968(.dina(n4025), .dinb(n4024), .dout(n4026));
  jand g3969(.dina(n4026), .dinb(n4021), .dout(n4027));
  jxor g3970(.dina(n4027), .dinb(n1257), .dout(n4028));
  jxor g3971(.dina(n4028), .dinb(n4020), .dout(n4029));
  jxor g3972(.dina(n4029), .dinb(n3989), .dout(n4030));
  jor  g3973(.dina(n3566), .dinb(n3029), .dout(n4031));
  jor  g3974(.dina(n3510), .dinb(n3213), .dout(n4032));
  jor  g3975(.dina(n3495), .dinb(n3210), .dout(n4033));
  jor  g3976(.dina(n3441), .dinb(n3219), .dout(n4034));
  jand g3977(.dina(n4034), .dinb(n4033), .dout(n4035));
  jand g3978(.dina(n4035), .dinb(n4032), .dout(n4036));
  jand g3979(.dina(n4036), .dinb(n4031), .dout(n4037));
  jxor g3980(.dina(n4037), .dinb(n1156), .dout(n4038));
  jxor g3981(.dina(n4038), .dinb(n4030), .dout(n4039));
  jxor g3982(.dina(n4039), .dinb(n3985), .dout(n4040));
  jnot g3983(.din(n3841), .dout(n4041));
  jor  g3984(.dina(n4041), .dinb(n3824), .dout(n4042));
  jand g3985(.dina(n4042), .dinb(n3840), .dout(n4043));
  jand g3986(.dina(n2954), .dinb(n1133), .dout(n4044));
  jand g3987(.dina(n4044), .dinb(n3177), .dout(n4045));
  jand g3988(.dina(n404), .dinb(n182), .dout(n4046));
  jand g3989(.dina(n4046), .dinb(n1127), .dout(n4047));
  jand g3990(.dina(n4047), .dinb(n448), .dout(n4048));
  jand g3991(.dina(n385), .dinb(n251), .dout(n4049));
  jand g3992(.dina(n4049), .dinb(n321), .dout(n4050));
  jand g3993(.dina(n4050), .dinb(n4048), .dout(n4051));
  jand g3994(.dina(n4051), .dinb(n4045), .dout(n4052));
  jand g3995(.dina(n2127), .dinb(n482), .dout(n4053));
  jand g3996(.dina(n4053), .dinb(n252), .dout(n4054));
  jand g3997(.dina(n4054), .dinb(n1023), .dout(n4055));
  jand g3998(.dina(n233), .dinb(n176), .dout(n4056));
  jand g3999(.dina(n4056), .dinb(n4055), .dout(n4057));
  jand g4000(.dina(n4057), .dinb(n4052), .dout(n4058));
  jand g4001(.dina(n4058), .dinb(n834), .dout(n4059));
  jand g4002(.dina(n4059), .dinb(n3837), .dout(n4060));
  jnot g4003(.din(n4060), .dout(n4061));
  jand g4004(.dina(n3833), .dinb(n3836), .dout(n4062));
  jxor g4005(.dina(n4059), .dinb(n4062), .dout(n4063));
  jor  g4006(.dina(n4063), .dinb(n3837), .dout(n4064));
  jand g4007(.dina(n4064), .dinb(n4061), .dout(n4065));
  jxor g4008(.dina(n4065), .dinb(n4043), .dout(n4066));
  jor  g4009(.dina(n4066), .dinb(n3461), .dout(n4067));
  jor  g4010(.dina(n3552), .dinb(n3547), .dout(n4068));
  jor  g4011(.dina(n3837), .dinb(n3558), .dout(n4069));
  jor  g4012(.dina(n4063), .dinb(n3554), .dout(n4070));
  jand g4013(.dina(n4070), .dinb(n4069), .dout(n4071));
  jand g4014(.dina(n4071), .dinb(n4068), .dout(n4072));
  jand g4015(.dina(n4072), .dinb(n4067), .dout(n4073));
  jxor g4016(.dina(n4073), .dinb(n3023), .dout(n4074));
  jxor g4017(.dina(n4074), .dinb(n4040), .dout(n4075));
  jxor g4018(.dina(n4075), .dinb(n3982), .dout(n4076));
  jnot g4019(.din(n190), .dout(n4077));
  jor  g4020(.dina(n1319), .dinb(n4077), .dout(n4078));
  jor  g4021(.dina(n4078), .dinb(n628), .dout(n4079));
  jnot g4022(.din(n4079), .dout(n4080));
  jand g4023(.dina(n4080), .dinb(n1392), .dout(n4081));
  jand g4024(.dina(n1072), .dinb(n251), .dout(n4082));
  jand g4025(.dina(n4082), .dinb(n128), .dout(n4083));
  jand g4026(.dina(n825), .dinb(n102), .dout(n4084));
  jand g4027(.dina(n4084), .dinb(n4083), .dout(n4085));
  jand g4028(.dina(n4085), .dinb(n4081), .dout(n4086));
  jand g4029(.dina(n2631), .dinb(n1069), .dout(n4087));
  jand g4030(.dina(n4087), .dinb(n4086), .dout(n4088));
  jxor g4031(.dina(n4088), .dinb(n4076), .dout(n4089));
  jxor g4032(.dina(n4089), .dinb(n3971), .dout(n4090));
  jxor g4033(.dina(n3969), .dinb(n3854), .dout(n4091));
  jxor g4034(.dina(n4091), .dinb(n4090), .dout(sin0 ));
  jxor g4035(.dina(a23 ), .dinb(a22 ), .dout(n4093));
  jand g4036(.dina(n4093), .dinb(sin0 ), .dout(n4094));
  jnot g4037(.din(n4094), .dout(n4095));
  jand g4038(.dina(n4091), .dinb(n4090), .dout(n4096));
  jor  g4039(.dina(n4088), .dinb(n4076), .dout(n4097));
  jnot g4040(.din(n4097), .dout(n4098));
  jand g4041(.dina(n4089), .dinb(n3971), .dout(n4099));
  jor  g4042(.dina(n4099), .dinb(n4098), .dout(n4100));
  jand g4043(.dina(n4074), .dinb(n4040), .dout(n4101));
  jnot g4044(.din(n4101), .dout(n4102));
  jnot g4045(.din(n4075), .dout(n4103));
  jor  g4046(.dina(n4103), .dinb(n3982), .dout(n4104));
  jand g4047(.dina(n4104), .dinb(n4102), .dout(n4105));
  jand g4048(.dina(n4038), .dinb(n4030), .dout(n4106));
  jand g4049(.dina(n4039), .dinb(n3985), .dout(n4107));
  jor  g4050(.dina(n4107), .dinb(n4106), .dout(n4108));
  jor  g4051(.dina(n4028), .dinb(n4020), .dout(n4109));
  jnot g4052(.din(n4109), .dout(n4110));
  jand g4053(.dina(n4029), .dinb(n3989), .dout(n4111));
  jor  g4054(.dina(n4111), .dinb(n4110), .dout(n4112));
  jand g4055(.dina(n4017), .dinb(n4009), .dout(n4113));
  jand g4056(.dina(n4018), .dinb(n3992), .dout(n4114));
  jor  g4057(.dina(n4114), .dinb(n4113), .dout(n4115));
  jor  g4058(.dina(n4008), .dinb(n3998), .dout(n4116));
  jand g4059(.dina(n4006), .dinb(n1438), .dout(n4117));
  jand g4060(.dina(n4117), .dinb(n2236), .dout(n4118));
  jnot g4061(.din(n4118), .dout(n4119));
  jand g4062(.dina(n4119), .dinb(n4116), .dout(n4120));
  jor  g4063(.dina(n2825), .dinb(n3384), .dout(n4121));
  jand g4064(.dina(n2684), .dinb(n2488), .dout(n4122));
  jand g4065(.dina(n2683), .dinb(n2491), .dout(n4123));
  jand g4066(.dina(n2923), .dinb(n2687), .dout(n4124));
  jor  g4067(.dina(n4124), .dinb(n4123), .dout(n4125));
  jor  g4068(.dina(n4125), .dinb(n4122), .dout(n4126));
  jnot g4069(.din(n4126), .dout(n4127));
  jand g4070(.dina(n4127), .dinb(n4121), .dout(n4128));
  jand g4071(.dina(n2351), .dinb(n1438), .dout(n4129));
  jxor g4072(.dina(n4129), .dinb(n4128), .dout(n4130));
  jxor g4073(.dina(n4130), .dinb(n4120), .dout(n4131));
  jnot g4074(.din(n4131), .dout(n4132));
  jor  g4075(.dina(n3242), .dinb(n2252), .dout(n4133));
  jor  g4076(.dina(n3008), .dinb(n2359), .dout(n4134));
  jor  g4077(.dina(n3216), .dinb(n2355), .dout(n4135));
  jand g4078(.dina(n4135), .dinb(n4134), .dout(n4136));
  jor  g4079(.dina(n2800), .dinb(n2357), .dout(n4137));
  jand g4080(.dina(n4137), .dinb(n4136), .dout(n4138));
  jand g4081(.dina(n4138), .dinb(n4133), .dout(n4139));
  jxor g4082(.dina(n4139), .dinb(n1356), .dout(n4140));
  jxor g4083(.dina(n4140), .dinb(n4132), .dout(n4141));
  jxor g4084(.dina(n4141), .dinb(n4115), .dout(n4142));
  jnot g4085(.din(n4142), .dout(n4143));
  jor  g4086(.dina(n3443), .dinb(n2506), .dout(n4144));
  jor  g4087(.dina(n3441), .dinb(n2810), .dout(n4145));
  jor  g4088(.dina(n3203), .dinb(n2807), .dout(n4146));
  jand g4089(.dina(n4146), .dinb(n4145), .dout(n4147));
  jor  g4090(.dina(n3166), .dinb(n2816), .dout(n4148));
  jand g4091(.dina(n4148), .dinb(n4147), .dout(n4149));
  jand g4092(.dina(n4149), .dinb(n4144), .dout(n4150));
  jxor g4093(.dina(n4150), .dinb(n1257), .dout(n4151));
  jxor g4094(.dina(n4151), .dinb(n4143), .dout(n4152));
  jxor g4095(.dina(n4152), .dinb(n4112), .dout(n4153));
  jor  g4096(.dina(n3550), .dinb(n3029), .dout(n4154));
  jor  g4097(.dina(n3547), .dinb(n3213), .dout(n4155));
  jor  g4098(.dina(n3510), .dinb(n3210), .dout(n4156));
  jor  g4099(.dina(n3495), .dinb(n3219), .dout(n4157));
  jand g4100(.dina(n4157), .dinb(n4156), .dout(n4158));
  jand g4101(.dina(n4158), .dinb(n4155), .dout(n4159));
  jand g4102(.dina(n4159), .dinb(n4154), .dout(n4160));
  jxor g4103(.dina(n4160), .dinb(n1156), .dout(n4161));
  jxor g4104(.dina(n4161), .dinb(n4153), .dout(n4162));
  jxor g4105(.dina(n4162), .dinb(n4108), .dout(n4163));
  jnot g4106(.din(n4064), .dout(n4164));
  jnot g4107(.din(n3548), .dout(n4165));
  jnot g4108(.din(n3511), .dout(n4166));
  jand g4109(.dina(n2472), .dinb(n3713), .dout(n4167));
  jor  g4110(.dina(n4167), .dinb(n2691), .dout(n4168));
  jand g4111(.dina(n2835), .dinb(n4168), .dout(n4169));
  jor  g4112(.dina(n4169), .dinb(n2688), .dout(n4170));
  jand g4113(.dina(n2824), .dinb(n4170), .dout(n4171));
  jor  g4114(.dina(n4171), .dinb(n2685), .dout(n4172));
  jand g4115(.dina(n2801), .dinb(n4172), .dout(n4173));
  jor  g4116(.dina(n4173), .dinb(n2944), .dout(n4174));
  jand g4117(.dina(n3009), .dinb(n4174), .dout(n4175));
  jor  g4118(.dina(n4175), .dinb(n3150), .dout(n4176));
  jand g4119(.dina(n3241), .dinb(n4176), .dout(n4177));
  jor  g4120(.dina(n4177), .dinb(n3148), .dout(n4178));
  jand g4121(.dina(n3228), .dinb(n4178), .dout(n4179));
  jor  g4122(.dina(n4179), .dinb(n3145), .dout(n4180));
  jand g4123(.dina(n3204), .dinb(n4180), .dout(n4181));
  jor  g4124(.dina(n4181), .dinb(n3416), .dout(n4182));
  jand g4125(.dina(n3442), .dinb(n4182), .dout(n4183));
  jor  g4126(.dina(n4183), .dinb(n3514), .dout(n4184));
  jand g4127(.dina(n3578), .dinb(n4184), .dout(n4185));
  jor  g4128(.dina(n4185), .dinb(n3521), .dout(n4186));
  jand g4129(.dina(n3529), .dinb(n4186), .dout(n4187));
  jor  g4130(.dina(n4187), .dinb(n4166), .dout(n4188));
  jand g4131(.dina(n3549), .dinb(n4188), .dout(n4189));
  jor  g4132(.dina(n4189), .dinb(n4165), .dout(n4190));
  jand g4133(.dina(n3841), .dinb(n4190), .dout(n4191));
  jor  g4134(.dina(n4191), .dinb(n3839), .dout(n4192));
  jand g4135(.dina(n4065), .dinb(n4192), .dout(n4193));
  jor  g4136(.dina(n4193), .dinb(n4164), .dout(n4194));
  jnot g4137(.din(n4062), .dout(n4195));
  jnot g4138(.din(n4059), .dout(n4196));
  jand g4139(.dina(n4196), .dinb(n4195), .dout(n4197));
  jand g4140(.dina(n2155), .dinb(n340), .dout(n4198));
  jand g4141(.dina(n310), .dinb(n114), .dout(n4199));
  jand g4142(.dina(n4199), .dinb(n277), .dout(n4200));
  jand g4143(.dina(n4200), .dinb(n246), .dout(n4201));
  jand g4144(.dina(n4201), .dinb(n477), .dout(n4202));
  jand g4145(.dina(n4202), .dinb(n4198), .dout(n4203));
  jand g4146(.dina(n4203), .dinb(n1079), .dout(n4204));
  jand g4147(.dina(n4204), .dinb(n1339), .dout(n4205));
  jand g4148(.dina(n3497), .dinb(n439), .dout(n4206));
  jand g4149(.dina(n4206), .dinb(n333), .dout(n4207));
  jand g4150(.dina(n389), .dinb(n338), .dout(n4208));
  jand g4151(.dina(n540), .dinb(n446), .dout(n4209));
  jand g4152(.dina(n4209), .dinb(n4208), .dout(n4210));
  jand g4153(.dina(n4210), .dinb(n4207), .dout(n4211));
  jand g4154(.dina(n4211), .dinb(n2146), .dout(n4212));
  jand g4155(.dina(n4212), .dinb(n4205), .dout(n4213));
  jxor g4156(.dina(n4213), .dinb(n4197), .dout(n4214));
  jxor g4157(.dina(n4214), .dinb(n4194), .dout(n4215));
  jor  g4158(.dina(n4215), .dinb(n3461), .dout(n4216));
  jor  g4159(.dina(n4213), .dinb(n3554), .dout(n4219));
  jor  g4160(.dina(n3837), .dinb(n3552), .dout(n4220));
  jand g4161(.dina(n4220), .dinb(n4219), .dout(n4221));
  jor  g4162(.dina(n4063), .dinb(n3558), .dout(n4222));
  jand g4163(.dina(n4222), .dinb(n4221), .dout(n4223));
  jand g4164(.dina(n4223), .dinb(n4216), .dout(n4224));
  jxor g4165(.dina(n4224), .dinb(n3023), .dout(n4225));
  jxor g4166(.dina(n4225), .dinb(n4163), .dout(n4226));
  jxor g4167(.dina(n4226), .dinb(n4105), .dout(n4227));
  jand g4168(.dina(n190), .dinb(n136), .dout(n4228));
  jand g4169(.dina(n4228), .dinb(n3470), .dout(n4229));
  jand g4170(.dina(n2513), .dinb(n340), .dout(n4230));
  jand g4171(.dina(n383), .dinb(n286), .dout(n4231));
  jand g4172(.dina(n4231), .dinb(n817), .dout(n4232));
  jand g4173(.dina(n4232), .dinb(n4230), .dout(n4233));
  jand g4174(.dina(n4233), .dinb(n305), .dout(n4234));
  jand g4175(.dina(n4234), .dinb(n4229), .dout(n4235));
  jand g4176(.dina(n1313), .dinb(n569), .dout(n4236));
  jand g4177(.dina(n4236), .dinb(n169), .dout(n4237));
  jand g4178(.dina(n4237), .dinb(n114), .dout(n4238));
  jand g4179(.dina(n4238), .dinb(n587), .dout(n4239));
  jand g4180(.dina(n4239), .dinb(n4235), .dout(n4240));
  jand g4181(.dina(n2751), .dinb(n260), .dout(n4241));
  jand g4182(.dina(n4241), .dinb(n4240), .dout(n4242));
  jxor g4183(.dina(n4242), .dinb(n4227), .dout(n4243));
  jxor g4184(.dina(n4243), .dinb(n4100), .dout(n4244));
  jxor g4185(.dina(n4244), .dinb(n4096), .dout(n4245));
  jand g4186(.dina(n4245), .dinb(n4095), .dout(n4246));
  jnot g4187(.din(n4244), .dout(n4247));
  jand g4188(.dina(n4247), .dinb(n4094), .dout(n4248));
  jor  g4189(.dina(n4248), .dinb(n4246), .dout(sin1 ));
  jand g4190(.dina(n4244), .dinb(n4096), .dout(n4250));
  jor  g4191(.dina(n4242), .dinb(n4227), .dout(n4251));
  jnot g4192(.din(n4251), .dout(n4252));
  jand g4193(.dina(n4243), .dinb(n4100), .dout(n4253));
  jor  g4194(.dina(n4253), .dinb(n4252), .dout(n4254));
  jand g4195(.dina(n897), .dinb(n460), .dout(n4255));
  jand g4196(.dina(n4255), .dinb(n389), .dout(n4256));
  jand g4197(.dina(n4256), .dinb(n488), .dout(n4257));
  jand g4198(.dina(n4257), .dinb(n1109), .dout(n4258));
  jand g4199(.dina(n384), .dinb(n339), .dout(n4259));
  jand g4200(.dina(n4259), .dinb(n1365), .dout(n4260));
  jand g4201(.dina(n4260), .dinb(n124), .dout(n4261));
  jand g4202(.dina(n3179), .dinb(n176), .dout(n4262));
  jand g4203(.dina(n377), .dinb(n191), .dout(n4263));
  jand g4204(.dina(n221), .dinb(n158), .dout(n4264));
  jand g4205(.dina(n4264), .dinb(n4263), .dout(n4265));
  jand g4206(.dina(n4265), .dinb(n4262), .dout(n4266));
  jand g4207(.dina(n4266), .dinb(n1448), .dout(n4267));
  jand g4208(.dina(n4267), .dinb(n4261), .dout(n4268));
  jand g4209(.dina(n4268), .dinb(n3892), .dout(n4269));
  jand g4210(.dina(n4269), .dinb(n4258), .dout(n4270));
  jnot g4211(.din(n4270), .dout(n4271));
  jand g4212(.dina(n4225), .dinb(n4163), .dout(n4272));
  jand g4213(.dina(n3851), .dinb(n3763), .dout(n4273));
  jor  g4214(.dina(n4273), .dinb(n3972), .dout(n4274));
  jand g4215(.dina(n4075), .dinb(n4274), .dout(n4275));
  jor  g4216(.dina(n4275), .dinb(n4101), .dout(n4276));
  jand g4217(.dina(n4226), .dinb(n4276), .dout(n4277));
  jor  g4218(.dina(n4277), .dinb(n4272), .dout(n4278));
  jand g4219(.dina(n4161), .dinb(n4153), .dout(n4279));
  jand g4220(.dina(n4162), .dinb(n4108), .dout(n4280));
  jor  g4221(.dina(n4280), .dinb(n4279), .dout(n4281));
  jor  g4222(.dina(n4151), .dinb(n4143), .dout(n4282));
  jnot g4223(.din(n4282), .dout(n4283));
  jand g4224(.dina(n4152), .dinb(n4112), .dout(n4284));
  jor  g4225(.dina(n4284), .dinb(n4283), .dout(n4285));
  jor  g4226(.dina(n4140), .dinb(n4132), .dout(n4286));
  jand g4227(.dina(n4141), .dinb(n4115), .dout(n4287));
  jnot g4228(.din(n4287), .dout(n4288));
  jand g4229(.dina(n4288), .dinb(n4286), .dout(n4289));
  jnot g4230(.din(n4289), .dout(n4290));
  jor  g4231(.dina(n4130), .dinb(n4120), .dout(n4291));
  jand g4232(.dina(n4128), .dinb(n1438), .dout(n4292));
  jand g4233(.dina(n4292), .dinb(n2690), .dout(n4293));
  jnot g4234(.din(n4293), .dout(n4294));
  jand g4235(.dina(n4294), .dinb(n4291), .dout(n4295));
  jor  g4236(.dina(n2802), .dinb(n3384), .dout(n4296));
  jand g4237(.dina(n2943), .dinb(n2491), .dout(n4297));
  jand g4238(.dina(n2683), .dinb(n2488), .dout(n4298));
  jand g4239(.dina(n2923), .dinb(n2684), .dout(n4299));
  jor  g4240(.dina(n4299), .dinb(n4298), .dout(n4300));
  jor  g4241(.dina(n4300), .dinb(n4297), .dout(n4301));
  jnot g4242(.din(n4301), .dout(n4302));
  jand g4243(.dina(n4302), .dinb(n4296), .dout(n4303));
  jand g4244(.dina(n2471), .dinb(n1438), .dout(n4304));
  jxor g4245(.dina(n4304), .dinb(n4303), .dout(n4305));
  jxor g4246(.dina(n4305), .dinb(n4295), .dout(n4306));
  jnot g4247(.din(n4306), .dout(n4307));
  jor  g4248(.dina(n3229), .dinb(n2252), .dout(n4308));
  jor  g4249(.dina(n3166), .dinb(n2355), .dout(n4309));
  jor  g4250(.dina(n3216), .dinb(n2359), .dout(n4310));
  jand g4251(.dina(n4310), .dinb(n4309), .dout(n4311));
  jor  g4252(.dina(n3008), .dinb(n2357), .dout(n4312));
  jand g4253(.dina(n4312), .dinb(n4311), .dout(n4313));
  jand g4254(.dina(n4313), .dinb(n4308), .dout(n4314));
  jxor g4255(.dina(n4314), .dinb(n1356), .dout(n4315));
  jxor g4256(.dina(n4315), .dinb(n4307), .dout(n4316));
  jxor g4257(.dina(n4316), .dinb(n4290), .dout(n4317));
  jor  g4258(.dina(n3579), .dinb(n2506), .dout(n4318));
  jor  g4259(.dina(n3495), .dinb(n2810), .dout(n4319));
  jor  g4260(.dina(n3203), .dinb(n2816), .dout(n4320));
  jor  g4261(.dina(n3441), .dinb(n2807), .dout(n4321));
  jand g4262(.dina(n4321), .dinb(n4320), .dout(n4322));
  jand g4263(.dina(n4322), .dinb(n4319), .dout(n4323));
  jand g4264(.dina(n4323), .dinb(n4318), .dout(n4324));
  jxor g4265(.dina(n4324), .dinb(n1259), .dout(n4325));
  jxor g4266(.dina(n4325), .dinb(n4317), .dout(n4326));
  jxor g4267(.dina(n4326), .dinb(n4285), .dout(n4327));
  jor  g4268(.dina(n3842), .dinb(n3029), .dout(n4328));
  jor  g4269(.dina(n3837), .dinb(n3213), .dout(n4329));
  jor  g4270(.dina(n3547), .dinb(n3210), .dout(n4330));
  jor  g4271(.dina(n3510), .dinb(n3219), .dout(n4331));
  jand g4272(.dina(n4331), .dinb(n4330), .dout(n4332));
  jand g4273(.dina(n4332), .dinb(n4329), .dout(n4333));
  jand g4274(.dina(n4333), .dinb(n4328), .dout(n4334));
  jxor g4275(.dina(n4334), .dinb(n1156), .dout(n4335));
  jxor g4276(.dina(n4335), .dinb(n4327), .dout(n4336));
  jxor g4277(.dina(n4336), .dinb(n4281), .dout(n4337));
  jnot g4278(.din(n4213), .dout(n4338));
  jnot g4279(.din(n4063), .dout(n4339));
  jnot g4280(.din(n4214), .dout(n4340));
  jand g4281(.dina(n4340), .dinb(n4194), .dout(n4341));
  jor  g4282(.dina(n4341), .dinb(n4339), .dout(n4342));
  jand g4283(.dina(n4342), .dinb(n4338), .dout(n4343));
  jnot g4284(.din(n4065), .dout(n4344));
  jor  g4285(.dina(n4344), .dinb(n4043), .dout(n4345));
  jand g4286(.dina(n4345), .dinb(n4064), .dout(n4346));
  jor  g4287(.dina(n4214), .dinb(n4346), .dout(n4347));
  jand g4288(.dina(n4213), .dinb(n4347), .dout(n4348));
  jor  g4289(.dina(n4348), .dinb(n4343), .dout(n4349));
  jor  g4290(.dina(n4349), .dinb(n3461), .dout(n4350));
  jor  g4291(.dina(n4063), .dinb(n3552), .dout(n4351));
  jor  g4292(.dina(n4213), .dinb(n3558), .dout(n4352));
  jand g4293(.dina(n4352), .dinb(n4351), .dout(n4353));
  jand g4294(.dina(n4353), .dinb(n4350), .dout(n4354));
  jxor g4295(.dina(n4354), .dinb(n3023), .dout(n4355));
  jxor g4296(.dina(n4355), .dinb(n4337), .dout(n4356));
  jxor g4297(.dina(n4356), .dinb(n4278), .dout(n4357));
  jxor g4298(.dina(n4357), .dinb(n4271), .dout(n4358));
  jxor g4299(.dina(n4358), .dinb(n4254), .dout(n4359));
  jxor g4300(.dina(n4359), .dinb(n4250), .dout(n4360));
  jor  g4301(.dina(n4245), .dinb(sin0 ), .dout(n4361));
  jand g4302(.dina(n4361), .dinb(n4093), .dout(n4362));
  jxor g4303(.dina(n4362), .dinb(n4360), .dout(sin2 ));
  jor  g4304(.dina(n4361), .dinb(n4360), .dout(n4364));
  jand g4305(.dina(n4364), .dinb(n4093), .dout(n4365));
  jand g4306(.dina(n4359), .dinb(n4250), .dout(n4366));
  jand g4307(.dina(n4357), .dinb(n4271), .dout(n4367));
  jand g4308(.dina(n4358), .dinb(n4254), .dout(n4368));
  jor  g4309(.dina(n4368), .dinb(n4367), .dout(n4369));
  jand g4310(.dina(n2964), .dinb(n535), .dout(n4370));
  jand g4311(.dina(n4370), .dinb(n2513), .dout(n4371));
  jand g4312(.dina(n4371), .dinb(n2738), .dout(n4372));
  jand g4313(.dina(n1460), .dinb(n462), .dout(n4373));
  jand g4314(.dina(n4373), .dinb(n1135), .dout(n4374));
  jand g4315(.dina(n4374), .dinb(n4372), .dout(n4375));
  jand g4316(.dina(n3875), .dinb(n197), .dout(n4376));
  jand g4317(.dina(n568), .dinb(n286), .dout(n4377));
  jand g4318(.dina(n4377), .dinb(n1045), .dout(n4378));
  jand g4319(.dina(n4378), .dinb(n4376), .dout(n4379));
  jand g4320(.dina(n4379), .dinb(n1331), .dout(n4380));
  jand g4321(.dina(n4380), .dinb(n4375), .dout(n4381));
  jnot g4322(.din(n4381), .dout(n4382));
  jand g4323(.dina(n4355), .dinb(n4337), .dout(n4383));
  jand g4324(.dina(n4356), .dinb(n4278), .dout(n4384));
  jor  g4325(.dina(n4384), .dinb(n4383), .dout(n4385));
  jand g4326(.dina(n4335), .dinb(n4327), .dout(n4386));
  jand g4327(.dina(n4336), .dinb(n4281), .dout(n4387));
  jor  g4328(.dina(n4387), .dinb(n4386), .dout(n4388));
  jand g4329(.dina(n4325), .dinb(n4317), .dout(n4389));
  jand g4330(.dina(n4326), .dinb(n4285), .dout(n4390));
  jor  g4331(.dina(n4390), .dinb(n4389), .dout(n4391));
  jor  g4332(.dina(n4315), .dinb(n4307), .dout(n4392));
  jand g4333(.dina(n4316), .dinb(n4290), .dout(n4393));
  jnot g4334(.din(n4393), .dout(n4394));
  jand g4335(.dina(n4394), .dinb(n4392), .dout(n4395));
  jnot g4336(.din(n4395), .dout(n4396));
  jor  g4337(.dina(n4305), .dinb(n4295), .dout(n4397));
  jand g4338(.dina(n4303), .dinb(n1438), .dout(n4398));
  jand g4339(.dina(n4398), .dinb(n2687), .dout(n4399));
  jnot g4340(.din(n4399), .dout(n4400));
  jand g4341(.dina(n4400), .dinb(n4397), .dout(n4401));
  jor  g4342(.dina(n3010), .dinb(n3384), .dout(n4402));
  jand g4343(.dina(n2943), .dinb(n2488), .dout(n4403));
  jand g4344(.dina(n3147), .dinb(n2491), .dout(n4404));
  jand g4345(.dina(n2923), .dinb(n2683), .dout(n4405));
  jor  g4346(.dina(n4405), .dinb(n4404), .dout(n4406));
  jor  g4347(.dina(n4406), .dinb(n4403), .dout(n4407));
  jnot g4348(.din(n4407), .dout(n4408));
  jand g4349(.dina(n4408), .dinb(n4402), .dout(n4409));
  jand g4350(.dina(n2813), .dinb(n1438), .dout(n4410));
  jxor g4351(.dina(n4410), .dinb(n4409), .dout(n4411));
  jxor g4352(.dina(n4411), .dinb(n4401), .dout(n4412));
  jnot g4353(.din(n4412), .dout(n4413));
  jor  g4354(.dina(n3205), .dinb(n2252), .dout(n4414));
  jor  g4355(.dina(n3166), .dinb(n2359), .dout(n4415));
  jor  g4356(.dina(n3203), .dinb(n2355), .dout(n4416));
  jand g4357(.dina(n4416), .dinb(n4415), .dout(n4417));
  jor  g4358(.dina(n3216), .dinb(n2357), .dout(n4418));
  jand g4359(.dina(n4418), .dinb(n4417), .dout(n4419));
  jand g4360(.dina(n4419), .dinb(n4414), .dout(n4420));
  jxor g4361(.dina(n4420), .dinb(n1356), .dout(n4421));
  jxor g4362(.dina(n4421), .dinb(n4413), .dout(n4422));
  jxor g4363(.dina(n4422), .dinb(n4396), .dout(n4423));
  jnot g4364(.din(n4423), .dout(n4424));
  jor  g4365(.dina(n3566), .dinb(n2506), .dout(n4425));
  jor  g4366(.dina(n3495), .dinb(n2807), .dout(n4426));
  jor  g4367(.dina(n3510), .dinb(n2810), .dout(n4427));
  jand g4368(.dina(n4427), .dinb(n4426), .dout(n4428));
  jor  g4369(.dina(n3441), .dinb(n2816), .dout(n4429));
  jand g4370(.dina(n4429), .dinb(n4428), .dout(n4430));
  jand g4371(.dina(n4430), .dinb(n4425), .dout(n4431));
  jxor g4372(.dina(n4431), .dinb(n1257), .dout(n4432));
  jxor g4373(.dina(n4432), .dinb(n4424), .dout(n4433));
  jxor g4374(.dina(n4433), .dinb(n4391), .dout(n4434));
  jor  g4375(.dina(n4066), .dinb(n3029), .dout(n4435));
  jor  g4376(.dina(n3837), .dinb(n3210), .dout(n4436));
  jor  g4377(.dina(n4063), .dinb(n3213), .dout(n4437));
  jand g4378(.dina(n4437), .dinb(n4436), .dout(n4438));
  jor  g4379(.dina(n3547), .dinb(n3219), .dout(n4439));
  jand g4380(.dina(n4439), .dinb(n4438), .dout(n4440));
  jand g4381(.dina(n4440), .dinb(n4435), .dout(n4441));
  jxor g4382(.dina(n4441), .dinb(n1154), .dout(n4442));
  jxor g4383(.dina(n4442), .dinb(n4434), .dout(n4443));
  jor  g4384(.dina(n4213), .dinb(n3552), .dout(n4444));
  jnot g4385(.din(n4343), .dout(n4445));
  jor  g4386(.dina(n4445), .dinb(n3461), .dout(n4446));
  jand g4387(.dina(n4446), .dinb(n4444), .dout(n4447));
  jxor g4388(.dina(n4447), .dinb(n3455), .dout(n4448));
  jxor g4389(.dina(n4448), .dinb(n4443), .dout(n4449));
  jxor g4390(.dina(n4449), .dinb(n4388), .dout(n4450));
  jxor g4391(.dina(n4450), .dinb(n4385), .dout(n4451));
  jxor g4392(.dina(n4451), .dinb(n4382), .dout(n4452));
  jxor g4393(.dina(n4452), .dinb(n4369), .dout(n4453));
  jxor g4394(.dina(n4453), .dinb(n4366), .dout(n4454));
  jxor g4395(.dina(n4454), .dinb(n4365), .dout(sin3 ));
  jand g4396(.dina(n4453), .dinb(n4366), .dout(n4456));
  jand g4397(.dina(n4451), .dinb(n4382), .dout(n4457));
  jand g4398(.dina(n4452), .dinb(n4369), .dout(n4458));
  jor  g4399(.dina(n4458), .dinb(n4457), .dout(n4459));
  jand g4400(.dina(n1073), .dinb(n280), .dout(n4460));
  jand g4401(.dina(n4460), .dinb(n1322), .dout(n4461));
  jand g4402(.dina(n4461), .dinb(n552), .dout(n4462));
  jand g4403(.dina(n4462), .dinb(n300), .dout(n4463));
  jand g4404(.dina(n2127), .dinb(n904), .dout(n4464));
  jand g4405(.dina(n4464), .dinb(n3179), .dout(n4465));
  jand g4406(.dina(n4465), .dinb(n1235), .dout(n4466));
  jand g4407(.dina(n4466), .dinb(n1974), .dout(n4467));
  jand g4408(.dina(n4467), .dinb(n1016), .dout(n4468));
  jand g4409(.dina(n4468), .dinb(n4463), .dout(n4469));
  jnot g4410(.din(n4469), .dout(n4470));
  jand g4411(.dina(n4449), .dinb(n4388), .dout(n4471));
  jand g4412(.dina(n4450), .dinb(n4385), .dout(n4472));
  jor  g4413(.dina(n4472), .dinb(n4471), .dout(n4473));
  jnot g4414(.din(n4434), .dout(n4474));
  jor  g4415(.dina(n4442), .dinb(n4474), .dout(n4475));
  jnot g4416(.din(n4475), .dout(n4476));
  jnot g4417(.din(n4443), .dout(n4477));
  jnot g4418(.din(n4448), .dout(n4478));
  jand g4419(.dina(n4478), .dinb(n4477), .dout(n4479));
  jor  g4420(.dina(n4479), .dinb(n4476), .dout(n4480));
  jor  g4421(.dina(n4432), .dinb(n4424), .dout(n4481));
  jand g4422(.dina(n4433), .dinb(n4391), .dout(n4482));
  jnot g4423(.din(n4482), .dout(n4483));
  jand g4424(.dina(n4483), .dinb(n4481), .dout(n4484));
  jor  g4425(.dina(n4421), .dinb(n4413), .dout(n4485));
  jand g4426(.dina(n4422), .dinb(n4396), .dout(n4486));
  jnot g4427(.din(n4486), .dout(n4487));
  jand g4428(.dina(n4487), .dinb(n4485), .dout(n4488));
  jnot g4429(.din(n4488), .dout(n4489));
  jor  g4430(.dina(n4411), .dinb(n4401), .dout(n4490));
  jand g4431(.dina(n4409), .dinb(n1438), .dout(n4491));
  jand g4432(.dina(n4491), .dinb(n2684), .dout(n4492));
  jnot g4433(.din(n4492), .dout(n4493));
  jand g4434(.dina(n4493), .dinb(n4490), .dout(n4494));
  jnot g4435(.din(n4494), .dout(n4495));
  jand g4436(.dina(n2683), .dinb(n1438), .dout(n4496));
  jxor g4437(.dina(n4496), .dinb(n3455), .dout(n4497));
  jor  g4438(.dina(n3242), .dinb(n3384), .dout(n4498));
  jor  g4439(.dina(n3008), .dinb(n3390), .dout(n4499));
  jor  g4440(.dina(n3216), .dinb(n3386), .dout(n4500));
  jand g4441(.dina(n4500), .dinb(n4499), .dout(n4501));
  jor  g4442(.dina(n3388), .dinb(n2800), .dout(n4502));
  jand g4443(.dina(n4502), .dinb(n4501), .dout(n4503));
  jand g4444(.dina(n4503), .dinb(n4498), .dout(n4504));
  jxor g4445(.dina(n4504), .dinb(n2051), .dout(n4505));
  jxor g4446(.dina(n4505), .dinb(n4497), .dout(n4506));
  jxor g4447(.dina(n4506), .dinb(n4495), .dout(n4507));
  jnot g4448(.din(n4507), .dout(n4508));
  jor  g4449(.dina(n3443), .dinb(n2252), .dout(n4509));
  jor  g4450(.dina(n3441), .dinb(n2355), .dout(n4510));
  jor  g4451(.dina(n3203), .dinb(n2359), .dout(n4511));
  jand g4452(.dina(n4511), .dinb(n4510), .dout(n4512));
  jor  g4453(.dina(n3166), .dinb(n2357), .dout(n4513));
  jand g4454(.dina(n4513), .dinb(n4512), .dout(n4514));
  jand g4455(.dina(n4514), .dinb(n4509), .dout(n4515));
  jxor g4456(.dina(n4515), .dinb(n1356), .dout(n4516));
  jxor g4457(.dina(n4516), .dinb(n4508), .dout(n4517));
  jxor g4458(.dina(n4517), .dinb(n4489), .dout(n4518));
  jor  g4459(.dina(n3550), .dinb(n2506), .dout(n4519));
  jor  g4460(.dina(n3547), .dinb(n2810), .dout(n4520));
  jor  g4461(.dina(n3510), .dinb(n2807), .dout(n4521));
  jor  g4462(.dina(n3495), .dinb(n2816), .dout(n4522));
  jand g4463(.dina(n4522), .dinb(n4521), .dout(n4523));
  jand g4464(.dina(n4523), .dinb(n4520), .dout(n4524));
  jand g4465(.dina(n4524), .dinb(n4519), .dout(n4525));
  jxor g4466(.dina(n4525), .dinb(n1259), .dout(n4526));
  jxor g4467(.dina(n4526), .dinb(n4518), .dout(n4527));
  jxor g4468(.dina(n4527), .dinb(n4484), .dout(n4528));
  jor  g4469(.dina(n4215), .dinb(n3029), .dout(n4529));
  jor  g4470(.dina(n4063), .dinb(n3210), .dout(n4530));
  jor  g4471(.dina(n3837), .dinb(n3219), .dout(n4531));
  jor  g4472(.dina(n4213), .dinb(n3213), .dout(n4532));
  jand g4473(.dina(n4532), .dinb(n4531), .dout(n4533));
  jand g4474(.dina(n4533), .dinb(n4530), .dout(n4534));
  jand g4475(.dina(n4534), .dinb(n4529), .dout(n4535));
  jxor g4476(.dina(n4535), .dinb(n1154), .dout(n4536));
  jxor g4477(.dina(n4536), .dinb(n4528), .dout(n4537));
  jxor g4478(.dina(n4537), .dinb(n4480), .dout(n4538));
  jxor g4479(.dina(n4538), .dinb(n4473), .dout(n4539));
  jxor g4480(.dina(n4539), .dinb(n4470), .dout(n4540));
  jxor g4481(.dina(n4540), .dinb(n4459), .dout(n4541));
  jxor g4482(.dina(n4541), .dinb(n4456), .dout(n4542));
  jor  g4483(.dina(n4454), .dinb(n4364), .dout(n4543));
  jand g4484(.dina(n4543), .dinb(n4093), .dout(n4544));
  jxor g4485(.dina(n4544), .dinb(n4542), .dout(sin4 ));
  jand g4486(.dina(n4541), .dinb(n4456), .dout(n4546));
  jand g4487(.dina(n4539), .dinb(n4470), .dout(n4547));
  jand g4488(.dina(n4540), .dinb(n4459), .dout(n4548));
  jor  g4489(.dina(n4548), .dinb(n4547), .dout(n4549));
  jand g4490(.dina(n361), .dinb(n280), .dout(n4550));
  jand g4491(.dina(n2617), .dinb(n850), .dout(n4551));
  jand g4492(.dina(n4551), .dinb(n4550), .dout(n4552));
  jand g4493(.dina(n4552), .dinb(n4203), .dout(n4553));
  jand g4494(.dina(n378), .dinb(n248), .dout(n4554));
  jand g4495(.dina(n4554), .dinb(n539), .dout(n4555));
  jand g4496(.dina(n2623), .dinb(n316), .dout(n4556));
  jand g4497(.dina(n510), .dinb(n411), .dout(n4557));
  jand g4498(.dina(n4557), .dinb(n535), .dout(n4558));
  jand g4499(.dina(n4558), .dinb(n4556), .dout(n4559));
  jand g4500(.dina(n4559), .dinb(n4555), .dout(n4560));
  jand g4501(.dina(n4560), .dinb(n4237), .dout(n4561));
  jand g4502(.dina(n4561), .dinb(n3481), .dout(n4562));
  jand g4503(.dina(n4562), .dinb(n4553), .dout(n4563));
  jnot g4504(.din(n4563), .dout(n4564));
  jand g4505(.dina(n4537), .dinb(n4480), .dout(n4565));
  jand g4506(.dina(n4538), .dinb(n4473), .dout(n4566));
  jor  g4507(.dina(n4566), .dinb(n4565), .dout(n4567));
  jnot g4508(.din(n4484), .dout(n4568));
  jand g4509(.dina(n4527), .dinb(n4568), .dout(n4569));
  jor  g4510(.dina(n4536), .dinb(n4528), .dout(n4570));
  jnot g4511(.din(n4570), .dout(n4571));
  jor  g4512(.dina(n4571), .dinb(n4569), .dout(n4572));
  jand g4513(.dina(n4517), .dinb(n4489), .dout(n4573));
  jand g4514(.dina(n4526), .dinb(n4518), .dout(n4574));
  jor  g4515(.dina(n4574), .dinb(n4573), .dout(n4575));
  jand g4516(.dina(n4506), .dinb(n4495), .dout(n4576));
  jnot g4517(.din(n4576), .dout(n4577));
  jor  g4518(.dina(n4516), .dinb(n4508), .dout(n4578));
  jand g4519(.dina(n4578), .dinb(n4577), .dout(n4579));
  jnot g4520(.din(n4579), .dout(n4580));
  jand g4521(.dina(n4496), .dinb(n3455), .dout(n4581));
  jand g4522(.dina(n4505), .dinb(n4497), .dout(n4582));
  jor  g4523(.dina(n4582), .dinb(n4581), .dout(n4583));
  jand g4524(.dina(n2943), .dinb(n1438), .dout(n4584));
  jxor g4525(.dina(n4584), .dinb(n3455), .dout(n4585));
  jxor g4526(.dina(n4585), .dinb(n4583), .dout(n4586));
  jor  g4527(.dina(n3229), .dinb(n3384), .dout(n4587));
  jor  g4528(.dina(n3166), .dinb(n3386), .dout(n4588));
  jor  g4529(.dina(n3216), .dinb(n3390), .dout(n4589));
  jand g4530(.dina(n4589), .dinb(n4588), .dout(n4590));
  jor  g4531(.dina(n3008), .dinb(n3388), .dout(n4591));
  jand g4532(.dina(n4591), .dinb(n4590), .dout(n4592));
  jand g4533(.dina(n4592), .dinb(n4587), .dout(n4593));
  jxor g4534(.dina(n4593), .dinb(n2051), .dout(n4594));
  jxor g4535(.dina(n4594), .dinb(n4586), .dout(n4595));
  jor  g4536(.dina(n3579), .dinb(n2252), .dout(n4596));
  jor  g4537(.dina(n3495), .dinb(n2355), .dout(n4597));
  jor  g4538(.dina(n3441), .dinb(n2359), .dout(n4598));
  jor  g4539(.dina(n3203), .dinb(n2357), .dout(n4599));
  jand g4540(.dina(n4599), .dinb(n4598), .dout(n4600));
  jand g4541(.dina(n4600), .dinb(n4597), .dout(n4601));
  jand g4542(.dina(n4601), .dinb(n4596), .dout(n4602));
  jxor g4543(.dina(n4602), .dinb(n1480), .dout(n4603));
  jxor g4544(.dina(n4603), .dinb(n4595), .dout(n4604));
  jxor g4545(.dina(n4604), .dinb(n4580), .dout(n4605));
  jnot g4546(.din(n4605), .dout(n4606));
  jor  g4547(.dina(n3842), .dinb(n2506), .dout(n4607));
  jor  g4548(.dina(n3547), .dinb(n2807), .dout(n4608));
  jor  g4549(.dina(n3837), .dinb(n2810), .dout(n4609));
  jand g4550(.dina(n4609), .dinb(n4608), .dout(n4610));
  jor  g4551(.dina(n3510), .dinb(n2816), .dout(n4611));
  jand g4552(.dina(n4611), .dinb(n4610), .dout(n4612));
  jand g4553(.dina(n4612), .dinb(n4607), .dout(n4613));
  jxor g4554(.dina(n4613), .dinb(n1257), .dout(n4614));
  jxor g4555(.dina(n4614), .dinb(n4606), .dout(n4615));
  jxor g4556(.dina(n4615), .dinb(n4575), .dout(n4616));
  jor  g4557(.dina(n4349), .dinb(n3029), .dout(n4617));
  jor  g4558(.dina(n4063), .dinb(n3219), .dout(n4618));
  jor  g4559(.dina(n4213), .dinb(n3210), .dout(n4619));
  jand g4560(.dina(n4619), .dinb(n4618), .dout(n4620));
  jand g4561(.dina(n4620), .dinb(n4617), .dout(n4621));
  jxor g4562(.dina(n4621), .dinb(n1156), .dout(n4622));
  jxor g4563(.dina(n4622), .dinb(n4616), .dout(n4623));
  jxor g4564(.dina(n4623), .dinb(n4572), .dout(n4624));
  jxor g4565(.dina(n4624), .dinb(n4567), .dout(n4625));
  jxor g4566(.dina(n4625), .dinb(n4564), .dout(n4626));
  jxor g4567(.dina(n4626), .dinb(n4549), .dout(n4627));
  jxor g4568(.dina(n4627), .dinb(n4546), .dout(n4628));
  jor  g4569(.dina(n4543), .dinb(n4542), .dout(n4629));
  jand g4570(.dina(n4629), .dinb(n4093), .dout(n4630));
  jxor g4571(.dina(n4630), .dinb(n4628), .dout(sin5 ));
  jand g4572(.dina(n4627), .dinb(n4546), .dout(n4632));
  jand g4573(.dina(n4625), .dinb(n4564), .dout(n4633));
  jand g4574(.dina(n4626), .dinb(n4549), .dout(n4634));
  jor  g4575(.dina(n4634), .dinb(n4633), .dout(n4635));
  jand g4576(.dina(n924), .dinb(n137), .dout(n4636));
  jand g4577(.dina(n4636), .dinb(n2623), .dout(n4637));
  jand g4578(.dina(n2513), .dinb(n540), .dout(n4638));
  jand g4579(.dina(n4638), .dinb(n4637), .dout(n4639));
  jand g4580(.dina(n3497), .dinb(n489), .dout(n4640));
  jand g4581(.dina(n4640), .dinb(n1122), .dout(n4641));
  jand g4582(.dina(n4641), .dinb(n2130), .dout(n4642));
  jand g4583(.dina(n4642), .dinb(n4639), .dout(n4643));
  jand g4584(.dina(n2628), .dinb(n276), .dout(n4644));
  jand g4585(.dina(n2135), .dinb(n128), .dout(n4645));
  jand g4586(.dina(n4645), .dinb(n4644), .dout(n4646));
  jand g4587(.dina(n4646), .dinb(n1970), .dout(n4647));
  jand g4588(.dina(n3537), .dinb(n142), .dout(n4648));
  jand g4589(.dina(n4648), .dinb(n288), .dout(n4649));
  jand g4590(.dina(n4649), .dinb(n4647), .dout(n4650));
  jand g4591(.dina(n4650), .dinb(n4643), .dout(n4651));
  jand g4592(.dina(n4651), .dinb(n273), .dout(n4652));
  jnot g4593(.din(n4652), .dout(n4653));
  jand g4594(.dina(n4623), .dinb(n4572), .dout(n4654));
  jand g4595(.dina(n4624), .dinb(n4567), .dout(n4655));
  jor  g4596(.dina(n4655), .dinb(n4654), .dout(n4656));
  jand g4597(.dina(n4615), .dinb(n4575), .dout(n4657));
  jand g4598(.dina(n4622), .dinb(n4616), .dout(n4658));
  jor  g4599(.dina(n4658), .dinb(n4657), .dout(n4659));
  jand g4600(.dina(n4604), .dinb(n4580), .dout(n4660));
  jnot g4601(.din(n4660), .dout(n4661));
  jor  g4602(.dina(n4614), .dinb(n4606), .dout(n4662));
  jand g4603(.dina(n4662), .dinb(n4661), .dout(n4663));
  jand g4604(.dina(n4338), .dinb(n3218), .dout(n4664));
  jand g4605(.dina(n4343), .dinb(n3028), .dout(n4665));
  jor  g4606(.dina(n4665), .dinb(n4664), .dout(n4666));
  jxor g4607(.dina(n4666), .dinb(n1156), .dout(n4667));
  jxor g4608(.dina(n4667), .dinb(n4663), .dout(n4668));
  jand g4609(.dina(n4594), .dinb(n4586), .dout(n4669));
  jand g4610(.dina(n4603), .dinb(n4595), .dout(n4670));
  jor  g4611(.dina(n4670), .dinb(n4669), .dout(n4671));
  jand g4612(.dina(n4584), .dinb(n3455), .dout(n4672));
  jand g4613(.dina(n4585), .dinb(n4583), .dout(n4673));
  jor  g4614(.dina(n4673), .dinb(n4672), .dout(n4674));
  jand g4615(.dina(n3147), .dinb(n1438), .dout(n4675));
  jxor g4616(.dina(n4675), .dinb(n3455), .dout(n4676));
  jxor g4617(.dina(n4676), .dinb(n4674), .dout(n4677));
  jor  g4618(.dina(n3205), .dinb(n3384), .dout(n4678));
  jor  g4619(.dina(n3166), .dinb(n3390), .dout(n4679));
  jor  g4620(.dina(n3203), .dinb(n3386), .dout(n4680));
  jand g4621(.dina(n4680), .dinb(n4679), .dout(n4681));
  jor  g4622(.dina(n3216), .dinb(n3388), .dout(n4682));
  jand g4623(.dina(n4682), .dinb(n4681), .dout(n4683));
  jand g4624(.dina(n4683), .dinb(n4678), .dout(n4684));
  jxor g4625(.dina(n4684), .dinb(n2051), .dout(n4685));
  jxor g4626(.dina(n4685), .dinb(n4677), .dout(n4686));
  jor  g4627(.dina(n3566), .dinb(n2252), .dout(n4687));
  jor  g4628(.dina(n3510), .dinb(n2355), .dout(n4688));
  jor  g4629(.dina(n3495), .dinb(n2359), .dout(n4689));
  jor  g4630(.dina(n3441), .dinb(n2357), .dout(n4690));
  jand g4631(.dina(n4690), .dinb(n4689), .dout(n4691));
  jand g4632(.dina(n4691), .dinb(n4688), .dout(n4692));
  jand g4633(.dina(n4692), .dinb(n4687), .dout(n4693));
  jxor g4634(.dina(n4693), .dinb(n1480), .dout(n4694));
  jxor g4635(.dina(n4694), .dinb(n4686), .dout(n4695));
  jxor g4636(.dina(n4695), .dinb(n4671), .dout(n4696));
  jnot g4637(.din(n4696), .dout(n4697));
  jor  g4638(.dina(n4066), .dinb(n2506), .dout(n4698));
  jor  g4639(.dina(n3837), .dinb(n2807), .dout(n4699));
  jor  g4640(.dina(n4063), .dinb(n2810), .dout(n4700));
  jand g4641(.dina(n4700), .dinb(n4699), .dout(n4701));
  jor  g4642(.dina(n3547), .dinb(n2816), .dout(n4702));
  jand g4643(.dina(n4702), .dinb(n4701), .dout(n4703));
  jand g4644(.dina(n4703), .dinb(n4698), .dout(n4704));
  jxor g4645(.dina(n4704), .dinb(n1257), .dout(n4705));
  jxor g4646(.dina(n4705), .dinb(n4697), .dout(n4706));
  jxor g4647(.dina(n4706), .dinb(n4668), .dout(n4707));
  jxor g4648(.dina(n4707), .dinb(n4659), .dout(n4708));
  jxor g4649(.dina(n4708), .dinb(n4656), .dout(n4709));
  jxor g4650(.dina(n4709), .dinb(n4653), .dout(n4710));
  jxor g4651(.dina(n4710), .dinb(n4635), .dout(n4711));
  jxor g4652(.dina(n4711), .dinb(n4632), .dout(n4712));
  jor  g4653(.dina(n4629), .dinb(n4628), .dout(n4713));
  jand g4654(.dina(n4713), .dinb(n4093), .dout(n4714));
  jxor g4655(.dina(n4714), .dinb(n4712), .dout(sin6 ));
  jand g4656(.dina(n4711), .dinb(n4632), .dout(n4716));
  jand g4657(.dina(n4709), .dinb(n4653), .dout(n4717));
  jand g4658(.dina(n4710), .dinb(n4635), .dout(n4718));
  jor  g4659(.dina(n4718), .dinb(n4717), .dout(n4719));
  jand g4660(.dina(n4707), .dinb(n4659), .dout(n4720));
  jand g4661(.dina(n4708), .dinb(n4656), .dout(n4721));
  jor  g4662(.dina(n4721), .dinb(n4720), .dout(n4722));
  jor  g4663(.dina(n4667), .dinb(n4663), .dout(n4723));
  jand g4664(.dina(n4706), .dinb(n4668), .dout(n4724));
  jnot g4665(.din(n4724), .dout(n4725));
  jand g4666(.dina(n4725), .dinb(n4723), .dout(n4726));
  jnot g4667(.din(n4726), .dout(n4727));
  jand g4668(.dina(n4695), .dinb(n4671), .dout(n4728));
  jnot g4669(.din(n4728), .dout(n4729));
  jor  g4670(.dina(n4705), .dinb(n4697), .dout(n4730));
  jand g4671(.dina(n4730), .dinb(n4729), .dout(n4731));
  jor  g4672(.dina(n4215), .dinb(n2506), .dout(n4732));
  jor  g4673(.dina(n4063), .dinb(n2807), .dout(n4733));
  jor  g4674(.dina(n3837), .dinb(n2816), .dout(n4734));
  jor  g4675(.dina(n4213), .dinb(n2810), .dout(n4735));
  jand g4676(.dina(n4735), .dinb(n4734), .dout(n4736));
  jand g4677(.dina(n4736), .dinb(n4733), .dout(n4737));
  jand g4678(.dina(n4737), .dinb(n4732), .dout(n4738));
  jxor g4679(.dina(n4738), .dinb(n1257), .dout(n4739));
  jxor g4680(.dina(n4739), .dinb(n4731), .dout(n4740));
  jand g4681(.dina(n4685), .dinb(n4677), .dout(n4741));
  jand g4682(.dina(n4694), .dinb(n4686), .dout(n4742));
  jor  g4683(.dina(n4742), .dinb(n4741), .dout(n4743));
  jand g4684(.dina(n4675), .dinb(n3455), .dout(n4744));
  jand g4685(.dina(n4676), .dinb(n4674), .dout(n4745));
  jor  g4686(.dina(n4745), .dinb(n4744), .dout(n4746));
  jand g4687(.dina(n3144), .dinb(n1438), .dout(n4747));
  jxor g4688(.dina(n3455), .dinb(n1154), .dout(n4748));
  jxor g4689(.dina(n4748), .dinb(n4747), .dout(n4749));
  jor  g4690(.dina(n3443), .dinb(n3384), .dout(n4750));
  jor  g4691(.dina(n3203), .dinb(n3390), .dout(n4751));
  jor  g4692(.dina(n3441), .dinb(n3386), .dout(n4752));
  jor  g4693(.dina(n3166), .dinb(n3388), .dout(n4753));
  jand g4694(.dina(n4753), .dinb(n4752), .dout(n4754));
  jand g4695(.dina(n4754), .dinb(n4751), .dout(n4755));
  jand g4696(.dina(n4755), .dinb(n4750), .dout(n4756));
  jxor g4697(.dina(n4756), .dinb(n2051), .dout(n4757));
  jxor g4698(.dina(n4757), .dinb(n4749), .dout(n4758));
  jxor g4699(.dina(n4758), .dinb(n4746), .dout(n4759));
  jor  g4700(.dina(n3550), .dinb(n2252), .dout(n4760));
  jor  g4701(.dina(n3547), .dinb(n2355), .dout(n4761));
  jor  g4702(.dina(n3510), .dinb(n2359), .dout(n4762));
  jor  g4703(.dina(n3495), .dinb(n2357), .dout(n4763));
  jand g4704(.dina(n4763), .dinb(n4762), .dout(n4764));
  jand g4705(.dina(n4764), .dinb(n4761), .dout(n4765));
  jand g4706(.dina(n4765), .dinb(n4760), .dout(n4766));
  jxor g4707(.dina(n4766), .dinb(n1480), .dout(n4767));
  jxor g4708(.dina(n4767), .dinb(n4759), .dout(n4768));
  jxor g4709(.dina(n4768), .dinb(n4743), .dout(n4769));
  jxor g4710(.dina(n4769), .dinb(n4740), .dout(n4770));
  jxor g4711(.dina(n4770), .dinb(n4727), .dout(n4771));
  jnot g4712(.din(n4771), .dout(n4772));
  jxor g4713(.dina(n4772), .dinb(n4722), .dout(n4773));
  jand g4714(.dina(n2618), .dinb(n588), .dout(n4774));
  jand g4715(.dina(n4774), .dinb(n4643), .dout(n4775));
  jand g4716(.dina(n1074), .dinb(n1033), .dout(n4776));
  jand g4717(.dina(n252), .dinb(n191), .dout(n4777));
  jand g4718(.dina(n4777), .dinb(n4776), .dout(n4778));
  jand g4719(.dina(n4778), .dinb(n4558), .dout(n4779));
  jand g4720(.dina(n4779), .dinb(n334), .dout(n4780));
  jand g4721(.dina(n4780), .dinb(n4775), .dout(n4781));
  jand g4722(.dina(n4781), .dinb(n2732), .dout(n4782));
  jxor g4723(.dina(n4782), .dinb(n4773), .dout(n4783));
  jxor g4724(.dina(n4783), .dinb(n4719), .dout(n4784));
  jxor g4725(.dina(n4784), .dinb(n4716), .dout(n4785));
  jor  g4726(.dina(n4713), .dinb(n4712), .dout(n4786));
  jand g4727(.dina(n4786), .dinb(n4093), .dout(n4787));
  jxor g4728(.dina(n4787), .dinb(n4785), .dout(sin7 ));
  jand g4729(.dina(n4784), .dinb(n4716), .dout(n4789));
  jor  g4730(.dina(n4782), .dinb(n4773), .dout(n4790));
  jnot g4731(.din(n4790), .dout(n4791));
  jand g4732(.dina(n4783), .dinb(n4719), .dout(n4792));
  jor  g4733(.dina(n4792), .dinb(n4791), .dout(n4793));
  jnot g4734(.din(n1188), .dout(n4794));
  jand g4735(.dina(n1984), .dinb(n1192), .dout(n4795));
  jand g4736(.dina(n4795), .dinb(n4794), .dout(n4796));
  jand g4737(.dina(n4796), .dinb(n195), .dout(n4797));
  jand g4738(.dina(n353), .dinb(n213), .dout(n4798));
  jand g4739(.dina(n4798), .dinb(n2510), .dout(n4799));
  jand g4740(.dina(n377), .dinb(n182), .dout(n4800));
  jand g4741(.dina(n4800), .dinb(n4799), .dout(n4801));
  jand g4742(.dina(n4801), .dinb(n4797), .dout(n4802));
  jand g4743(.dina(n387), .dinb(n235), .dout(n4803));
  jand g4744(.dina(n261), .dinb(n232), .dout(n4804));
  jand g4745(.dina(n4804), .dinb(n309), .dout(n4805));
  jand g4746(.dina(n4805), .dinb(n4803), .dout(n4806));
  jand g4747(.dina(n915), .dinb(n204), .dout(n4807));
  jand g4748(.dina(n4807), .dinb(n226), .dout(n4808));
  jand g4749(.dina(n4808), .dinb(n350), .dout(n4809));
  jand g4750(.dina(n4809), .dinb(n4806), .dout(n4810));
  jand g4751(.dina(n4810), .dinb(n180), .dout(n4811));
  jand g4752(.dina(n4811), .dinb(n3871), .dout(n4812));
  jand g4753(.dina(n4812), .dinb(n4802), .dout(n4813));
  jnot g4754(.din(n4813), .dout(n4814));
  jand g4755(.dina(n4770), .dinb(n4727), .dout(n4815));
  jand g4756(.dina(n4771), .dinb(n4722), .dout(n4816));
  jor  g4757(.dina(n4816), .dinb(n4815), .dout(n4817));
  jor  g4758(.dina(n4739), .dinb(n4731), .dout(n4818));
  jand g4759(.dina(n4769), .dinb(n4740), .dout(n4819));
  jnot g4760(.din(n4819), .dout(n4820));
  jand g4761(.dina(n4820), .dinb(n4818), .dout(n4821));
  jnot g4762(.din(n4821), .dout(n4822));
  jand g4763(.dina(n4767), .dinb(n4759), .dout(n4823));
  jand g4764(.dina(n4768), .dinb(n4743), .dout(n4824));
  jor  g4765(.dina(n4824), .dinb(n4823), .dout(n4825));
  jand g4766(.dina(n4757), .dinb(n4749), .dout(n4826));
  jand g4767(.dina(n4758), .dinb(n4746), .dout(n4827));
  jor  g4768(.dina(n4827), .dinb(n4826), .dout(n4828));
  jand g4769(.dina(n3143), .dinb(n1438), .dout(n4829));
  jnot g4770(.din(n4829), .dout(n4830));
  jand g4771(.dina(n3023), .dinb(n1156), .dout(n4831));
  jand g4772(.dina(n4748), .dinb(n4747), .dout(n4832));
  jor  g4773(.dina(n4832), .dinb(n4831), .dout(n4833));
  jxor g4774(.dina(n4833), .dinb(n4830), .dout(n4834));
  jor  g4775(.dina(n3579), .dinb(n3384), .dout(n4835));
  jor  g4776(.dina(n3495), .dinb(n3386), .dout(n4836));
  jor  g4777(.dina(n3203), .dinb(n3388), .dout(n4837));
  jor  g4778(.dina(n3441), .dinb(n3390), .dout(n4838));
  jand g4779(.dina(n4838), .dinb(n4837), .dout(n4839));
  jand g4780(.dina(n4839), .dinb(n4836), .dout(n4840));
  jand g4781(.dina(n4840), .dinb(n4835), .dout(n4841));
  jxor g4782(.dina(n4841), .dinb(n2051), .dout(n4842));
  jxor g4783(.dina(n4842), .dinb(n4834), .dout(n4843));
  jxor g4784(.dina(n4843), .dinb(n4828), .dout(n4844));
  jnot g4785(.din(n4844), .dout(n4845));
  jor  g4786(.dina(n3842), .dinb(n2252), .dout(n4846));
  jor  g4787(.dina(n3547), .dinb(n2359), .dout(n4847));
  jor  g4788(.dina(n3837), .dinb(n2355), .dout(n4848));
  jand g4789(.dina(n4848), .dinb(n4847), .dout(n4849));
  jor  g4790(.dina(n3510), .dinb(n2357), .dout(n4850));
  jand g4791(.dina(n4850), .dinb(n4849), .dout(n4851));
  jand g4792(.dina(n4851), .dinb(n4846), .dout(n4852));
  jxor g4793(.dina(n4852), .dinb(n1356), .dout(n4853));
  jxor g4794(.dina(n4853), .dinb(n4845), .dout(n4854));
  jxor g4795(.dina(n4854), .dinb(n4825), .dout(n4855));
  jor  g4796(.dina(n4349), .dinb(n2506), .dout(n4856));
  jor  g4797(.dina(n4063), .dinb(n2816), .dout(n4857));
  jor  g4798(.dina(n4213), .dinb(n2807), .dout(n4858));
  jand g4799(.dina(n4858), .dinb(n4857), .dout(n4859));
  jand g4800(.dina(n4859), .dinb(n4856), .dout(n4860));
  jxor g4801(.dina(n4860), .dinb(n1259), .dout(n4861));
  jxor g4802(.dina(n4861), .dinb(n4855), .dout(n4862));
  jxor g4803(.dina(n4862), .dinb(n4822), .dout(n4863));
  jxor g4804(.dina(n4863), .dinb(n4817), .dout(n4864));
  jxor g4805(.dina(n4864), .dinb(n4814), .dout(n4865));
  jxor g4806(.dina(n4865), .dinb(n4793), .dout(n4866));
  jxor g4807(.dina(n4866), .dinb(n4789), .dout(n4867));
  jor  g4808(.dina(n4786), .dinb(n4785), .dout(n4868));
  jand g4809(.dina(n4868), .dinb(n4093), .dout(n4869));
  jxor g4810(.dina(n4869), .dinb(n4867), .dout(sin8 ));
  jand g4811(.dina(n4866), .dinb(n4789), .dout(n4871));
  jand g4812(.dina(n4864), .dinb(n4814), .dout(n4872));
  jand g4813(.dina(n4865), .dinb(n4793), .dout(n4873));
  jor  g4814(.dina(n4873), .dinb(n4872), .dout(n4874));
  jand g4815(.dina(n3470), .dinb(n226), .dout(n4875));
  jand g4816(.dina(n1005), .dinb(n587), .dout(n4876));
  jand g4817(.dina(n346), .dinb(n160), .dout(n4877));
  jand g4818(.dina(n4877), .dinb(n4876), .dout(n4878));
  jand g4819(.dina(n3537), .dinb(n1074), .dout(n4879));
  jand g4820(.dina(n4879), .dinb(n4878), .dout(n4880));
  jand g4821(.dina(n255), .dinb(n244), .dout(n4881));
  jand g4822(.dina(n4881), .dinb(n1021), .dout(n4882));
  jand g4823(.dina(n4882), .dinb(n4880), .dout(n4883));
  jand g4824(.dina(n4883), .dinb(n4875), .dout(n4884));
  jand g4825(.dina(n4884), .dinb(n320), .dout(n4885));
  jand g4826(.dina(n4885), .dinb(n2146), .dout(n4886));
  jnot g4827(.din(n4886), .dout(n4887));
  jand g4828(.dina(n4862), .dinb(n4822), .dout(n4888));
  jand g4829(.dina(n4863), .dinb(n4817), .dout(n4889));
  jor  g4830(.dina(n4889), .dinb(n4888), .dout(n4890));
  jand g4831(.dina(n4854), .dinb(n4825), .dout(n4891));
  jand g4832(.dina(n4861), .dinb(n4855), .dout(n4892));
  jor  g4833(.dina(n4892), .dinb(n4891), .dout(n4893));
  jand g4834(.dina(n4843), .dinb(n4828), .dout(n4894));
  jnot g4835(.din(n4894), .dout(n4895));
  jor  g4836(.dina(n4853), .dinb(n4845), .dout(n4896));
  jand g4837(.dina(n4896), .dinb(n4895), .dout(n4897));
  jand g4838(.dina(n4338), .dinb(n2815), .dout(n4898));
  jand g4839(.dina(n4343), .dinb(n2505), .dout(n4899));
  jor  g4840(.dina(n4899), .dinb(n4898), .dout(n4900));
  jxor g4841(.dina(n4900), .dinb(n1259), .dout(n4901));
  jxor g4842(.dina(n4901), .dinb(n4897), .dout(n4902));
  jand g4843(.dina(n4833), .dinb(n4830), .dout(n4903));
  jand g4844(.dina(n4842), .dinb(n4834), .dout(n4904));
  jor  g4845(.dina(n4904), .dinb(n4903), .dout(n4905));
  jor  g4846(.dina(n3566), .dinb(n3384), .dout(n4906));
  jand g4847(.dina(n3520), .dinb(n2488), .dout(n4907));
  jnot g4848(.din(n3510), .dout(n4908));
  jand g4849(.dina(n4908), .dinb(n2491), .dout(n4909));
  jor  g4850(.dina(n4909), .dinb(n4907), .dout(n4910));
  jand g4851(.dina(n3513), .dinb(n2923), .dout(n4911));
  jor  g4852(.dina(n4911), .dinb(n4910), .dout(n4912));
  jnot g4853(.din(n4912), .dout(n4913));
  jand g4854(.dina(n4913), .dinb(n4906), .dout(n4914));
  jand g4855(.dina(n3418), .dinb(n1438), .dout(n4915));
  jxor g4856(.dina(n4915), .dinb(n4914), .dout(n4916));
  jxor g4857(.dina(n4916), .dinb(n4905), .dout(n4917));
  jnot g4858(.din(n4917), .dout(n4918));
  jor  g4859(.dina(n4066), .dinb(n2252), .dout(n4919));
  jor  g4860(.dina(n3837), .dinb(n2359), .dout(n4920));
  jor  g4861(.dina(n4063), .dinb(n2355), .dout(n4921));
  jand g4862(.dina(n4921), .dinb(n4920), .dout(n4922));
  jor  g4863(.dina(n3547), .dinb(n2357), .dout(n4923));
  jand g4864(.dina(n4923), .dinb(n4922), .dout(n4924));
  jand g4865(.dina(n4924), .dinb(n4919), .dout(n4925));
  jxor g4866(.dina(n4925), .dinb(n1356), .dout(n4926));
  jxor g4867(.dina(n4926), .dinb(n4918), .dout(n4927));
  jxor g4868(.dina(n4927), .dinb(n4902), .dout(n4928));
  jxor g4869(.dina(n4928), .dinb(n4893), .dout(n4929));
  jxor g4870(.dina(n4929), .dinb(n4890), .dout(n4930));
  jxor g4871(.dina(n4930), .dinb(n4887), .dout(n4931));
  jxor g4872(.dina(n4931), .dinb(n4874), .dout(n4932));
  jxor g4873(.dina(n4932), .dinb(n4871), .dout(n4933));
  jor  g4874(.dina(n4868), .dinb(n4867), .dout(n4934));
  jand g4875(.dina(n4934), .dinb(n4093), .dout(n4935));
  jxor g4876(.dina(n4935), .dinb(n4933), .dout(sin9 ));
  jand g4877(.dina(n4932), .dinb(n4871), .dout(n4937));
  jand g4878(.dina(n4930), .dinb(n4887), .dout(n4938));
  jand g4879(.dina(n4931), .dinb(n4874), .dout(n4939));
  jor  g4880(.dina(n4939), .dinb(n4938), .dout(n4940));
  jand g4881(.dina(n497), .dinb(n198), .dout(n4941));
  jand g4882(.dina(n3537), .dinb(n352), .dout(n4942));
  jand g4883(.dina(n4942), .dinb(n4941), .dout(n4943));
  jand g4884(.dina(n4943), .dinb(n1387), .dout(n4944));
  jand g4885(.dina(n534), .dinb(n190), .dout(n4945));
  jand g4886(.dina(n4945), .dinb(n297), .dout(n4946));
  jnot g4887(.din(n1186), .dout(n4947));
  jand g4888(.dina(n4947), .dinb(n506), .dout(n4948));
  jand g4889(.dina(n4948), .dinb(n4946), .dout(n4949));
  jand g4890(.dina(n4949), .dinb(n3881), .dout(n4950));
  jand g4891(.dina(n4950), .dinb(n896), .dout(n4951));
  jand g4892(.dina(n4951), .dinb(n4944), .dout(n4952));
  jnot g4893(.din(n4952), .dout(n4953));
  jand g4894(.dina(n4928), .dinb(n4893), .dout(n4954));
  jand g4895(.dina(n4929), .dinb(n4890), .dout(n4955));
  jor  g4896(.dina(n4955), .dinb(n4954), .dout(n4956));
  jor  g4897(.dina(n4901), .dinb(n4897), .dout(n4957));
  jand g4898(.dina(n4927), .dinb(n4902), .dout(n4958));
  jnot g4899(.din(n4958), .dout(n4959));
  jand g4900(.dina(n4959), .dinb(n4957), .dout(n4960));
  jnot g4901(.din(n4960), .dout(n4961));
  jor  g4902(.dina(n4914), .dinb(n1438), .dout(n4962));
  jand g4903(.dina(n4915), .dinb(n4914), .dout(n4963));
  jand g4904(.dina(n3415), .dinb(n1438), .dout(n4964));
  jand g4905(.dina(n4964), .dinb(n3166), .dout(n4965));
  jor  g4906(.dina(n4965), .dinb(n4963), .dout(n4966));
  jnot g4907(.din(n4966), .dout(n4967));
  jand g4908(.dina(n4967), .dinb(n4962), .dout(n4968));
  jnot g4909(.din(n4968), .dout(n4969));
  jand g4910(.dina(n3513), .dinb(n1438), .dout(n4970));
  jxor g4911(.dina(n4970), .dinb(n1259), .dout(n4971));
  jxor g4912(.dina(n4971), .dinb(n4829), .dout(n4972));
  jxor g4913(.dina(n4972), .dinb(n4969), .dout(n4973));
  jnot g4914(.din(n4973), .dout(n4974));
  jor  g4915(.dina(n3550), .dinb(n3384), .dout(n4975));
  jor  g4916(.dina(n3547), .dinb(n3386), .dout(n4976));
  jor  g4917(.dina(n3510), .dinb(n3390), .dout(n4977));
  jor  g4918(.dina(n3495), .dinb(n3388), .dout(n4978));
  jand g4919(.dina(n4978), .dinb(n4977), .dout(n4979));
  jand g4920(.dina(n4979), .dinb(n4976), .dout(n4980));
  jand g4921(.dina(n4980), .dinb(n4975), .dout(n4981));
  jxor g4922(.dina(n4981), .dinb(n1438), .dout(n4982));
  jxor g4923(.dina(n4982), .dinb(n4974), .dout(n4983));
  jand g4924(.dina(n4916), .dinb(n4905), .dout(n4984));
  jnot g4925(.din(n4984), .dout(n4985));
  jor  g4926(.dina(n4926), .dinb(n4918), .dout(n4986));
  jand g4927(.dina(n4986), .dinb(n4985), .dout(n4987));
  jnot g4928(.din(n4987), .dout(n4988));
  jor  g4929(.dina(n4215), .dinb(n2252), .dout(n4989));
  jor  g4930(.dina(n4213), .dinb(n2355), .dout(n4990));
  jor  g4931(.dina(n3837), .dinb(n2357), .dout(n4991));
  jand g4932(.dina(n4991), .dinb(n4990), .dout(n4992));
  jor  g4933(.dina(n4063), .dinb(n2359), .dout(n4993));
  jand g4934(.dina(n4993), .dinb(n4992), .dout(n4994));
  jand g4935(.dina(n4994), .dinb(n4989), .dout(n4995));
  jxor g4936(.dina(n4995), .dinb(n1480), .dout(n4996));
  jxor g4937(.dina(n4996), .dinb(n4988), .dout(n4997));
  jxor g4938(.dina(n4997), .dinb(n4983), .dout(n4998));
  jxor g4939(.dina(n4998), .dinb(n4961), .dout(n4999));
  jxor g4940(.dina(n4999), .dinb(n4956), .dout(n5000));
  jxor g4941(.dina(n5000), .dinb(n4953), .dout(n5001));
  jxor g4942(.dina(n5001), .dinb(n4940), .dout(n5002));
  jxor g4943(.dina(n5002), .dinb(n4937), .dout(n5003));
  jor  g4944(.dina(n4934), .dinb(n4933), .dout(n5004));
  jand g4945(.dina(n5004), .dinb(n4093), .dout(n5005));
  jxor g4946(.dina(n5005), .dinb(n5003), .dout(sin10 ));
  jand g4947(.dina(n5002), .dinb(n4937), .dout(n5007));
  jand g4948(.dina(n5000), .dinb(n4953), .dout(n5008));
  jand g4949(.dina(n5001), .dinb(n4940), .dout(n5009));
  jor  g4950(.dina(n5009), .dinb(n5008), .dout(n5010));
  jand g4951(.dina(n816), .dinb(n717), .dout(n5011));
  jand g4952(.dina(n5011), .dinb(n459), .dout(n5012));
  jand g4953(.dina(n5012), .dinb(n4051), .dout(n5013));
  jand g4954(.dina(n827), .dinb(n509), .dout(n5014));
  jand g4955(.dina(n5014), .dinb(n5013), .dout(n5015));
  jand g4956(.dina(n5015), .dinb(n1381), .dout(n5016));
  jnot g4957(.din(n5016), .dout(n5017));
  jand g4958(.dina(n4998), .dinb(n4961), .dout(n5018));
  jand g4959(.dina(n4999), .dinb(n4956), .dout(n5019));
  jor  g4960(.dina(n5019), .dinb(n5018), .dout(n5020));
  jand g4961(.dina(n4996), .dinb(n4988), .dout(n5021));
  jand g4962(.dina(n4997), .dinb(n4983), .dout(n5022));
  jor  g4963(.dina(n5022), .dinb(n5021), .dout(n5023));
  jand g4964(.dina(n4972), .dinb(n4969), .dout(n5024));
  jnot g4965(.din(n5024), .dout(n5025));
  jor  g4966(.dina(n4982), .dinb(n4974), .dout(n5026));
  jand g4967(.dina(n5026), .dinb(n5025), .dout(n5027));
  jnot g4968(.din(n5027), .dout(n5028));
  jand g4969(.dina(n3520), .dinb(n1438), .dout(n5029));
  jnot g4970(.din(n5029), .dout(n5030));
  jor  g4971(.dina(n4970), .dinb(n1259), .dout(n5031));
  jand g4972(.dina(n4970), .dinb(n1259), .dout(n5032));
  jor  g4973(.dina(n5032), .dinb(n4829), .dout(n5033));
  jand g4974(.dina(n5033), .dinb(n5031), .dout(n5034));
  jxor g4975(.dina(n5034), .dinb(n5030), .dout(n5035));
  jor  g4976(.dina(n3842), .dinb(n3384), .dout(n5036));
  jor  g4977(.dina(n3837), .dinb(n3386), .dout(n5037));
  jor  g4978(.dina(n3547), .dinb(n3390), .dout(n5038));
  jor  g4979(.dina(n3510), .dinb(n3388), .dout(n5039));
  jand g4980(.dina(n5039), .dinb(n5038), .dout(n5040));
  jand g4981(.dina(n5040), .dinb(n5037), .dout(n5041));
  jand g4982(.dina(n5041), .dinb(n5036), .dout(n5042));
  jxor g4983(.dina(n5042), .dinb(n2051), .dout(n5043));
  jxor g4984(.dina(n5043), .dinb(n5035), .dout(n5044));
  jxor g4985(.dina(n5044), .dinb(n5028), .dout(n5045));
  jor  g4986(.dina(n4349), .dinb(n2252), .dout(n5046));
  jor  g4987(.dina(n4063), .dinb(n2357), .dout(n5047));
  jor  g4988(.dina(n4213), .dinb(n2359), .dout(n5048));
  jand g4989(.dina(n5048), .dinb(n5047), .dout(n5049));
  jand g4990(.dina(n5049), .dinb(n5046), .dout(n5050));
  jxor g4991(.dina(n5050), .dinb(n1480), .dout(n5051));
  jxor g4992(.dina(n5051), .dinb(n5045), .dout(n5052));
  jxor g4993(.dina(n5052), .dinb(n5023), .dout(n5053));
  jxor g4994(.dina(n5053), .dinb(n5020), .dout(n5054));
  jxor g4995(.dina(n5054), .dinb(n5017), .dout(n5055));
  jxor g4996(.dina(n5055), .dinb(n5010), .dout(n5056));
  jxor g4997(.dina(n5056), .dinb(n5007), .dout(n5057));
  jor  g4998(.dina(n5004), .dinb(n5003), .dout(n5058));
  jand g4999(.dina(n5058), .dinb(n4093), .dout(n5059));
  jxor g5000(.dina(n5059), .dinb(n5057), .dout(sin11 ));
  jand g5001(.dina(n5056), .dinb(n5007), .dout(n5061));
  jand g5002(.dina(n5054), .dinb(n5017), .dout(n5062));
  jand g5003(.dina(n5055), .dinb(n5010), .dout(n5063));
  jor  g5004(.dina(n5063), .dinb(n5062), .dout(n5064));
  jand g5005(.dina(n2395), .dinb(n261), .dout(n5065));
  jand g5006(.dina(n5065), .dinb(n2971), .dout(n5066));
  jand g5007(.dina(n331), .dinb(n182), .dout(n5067));
  jand g5008(.dina(n313), .dinb(n278), .dout(n5068));
  jand g5009(.dina(n5068), .dinb(n244), .dout(n5069));
  jand g5010(.dina(n5069), .dinb(n5067), .dout(n5070));
  jand g5011(.dina(n5070), .dinb(n4266), .dout(n5071));
  jand g5012(.dina(n568), .dinb(n166), .dout(n5072));
  jand g5013(.dina(n5072), .dinb(n157), .dout(n5073));
  jand g5014(.dina(n5073), .dinb(n5071), .dout(n5074));
  jand g5015(.dina(n5074), .dinb(n2384), .dout(n5075));
  jand g5016(.dina(n5075), .dinb(n5066), .dout(n5076));
  jnot g5017(.din(n5076), .dout(n5077));
  jand g5018(.dina(n5052), .dinb(n5023), .dout(n5078));
  jand g5019(.dina(n5053), .dinb(n5020), .dout(n5079));
  jor  g5020(.dina(n5079), .dinb(n5078), .dout(n5080));
  jand g5021(.dina(n5044), .dinb(n5028), .dout(n5081));
  jand g5022(.dina(n5051), .dinb(n5045), .dout(n5082));
  jor  g5023(.dina(n5082), .dinb(n5081), .dout(n5083));
  jand g5024(.dina(n4338), .dinb(n2244), .dout(n5084));
  jand g5025(.dina(n4343), .dinb(n2101), .dout(n5085));
  jor  g5026(.dina(n5085), .dinb(n5084), .dout(n5086));
  jxor g5027(.dina(n5086), .dinb(n1356), .dout(n5087));
  jnot g5028(.din(n5087), .dout(n5088));
  jor  g5029(.dina(n4066), .dinb(n3384), .dout(n5089));
  jor  g5030(.dina(n3547), .dinb(n3388), .dout(n5090));
  jor  g5031(.dina(n3837), .dinb(n3390), .dout(n5091));
  jor  g5032(.dina(n4063), .dinb(n3386), .dout(n5092));
  jand g5033(.dina(n5092), .dinb(n5091), .dout(n5093));
  jand g5034(.dina(n5093), .dinb(n5090), .dout(n5094));
  jand g5035(.dina(n5094), .dinb(n5089), .dout(n5095));
  jxor g5036(.dina(n5095), .dinb(n1438), .dout(n5096));
  jxor g5037(.dina(n5096), .dinb(n5088), .dout(n5097));
  jand g5038(.dina(n5034), .dinb(n5030), .dout(n5098));
  jand g5039(.dina(n5043), .dinb(n5035), .dout(n5099));
  jor  g5040(.dina(n5099), .dinb(n5098), .dout(n5100));
  jand g5041(.dina(n5029), .dinb(n3510), .dout(n5101));
  jand g5042(.dina(n4908), .dinb(n1438), .dout(n5102));
  jand g5043(.dina(n5102), .dinb(n3495), .dout(n5103));
  jor  g5044(.dina(n5103), .dinb(n5101), .dout(n5104));
  jnot g5045(.din(n5104), .dout(n5105));
  jxor g5046(.dina(n5105), .dinb(n5100), .dout(n5106));
  jxor g5047(.dina(n5106), .dinb(n5097), .dout(n5107));
  jxor g5048(.dina(n5107), .dinb(n5083), .dout(n5108));
  jxor g5049(.dina(n5108), .dinb(n5080), .dout(n5109));
  jxor g5050(.dina(n5109), .dinb(n5077), .dout(n5110));
  jxor g5051(.dina(n5110), .dinb(n5064), .dout(n5111));
  jxor g5052(.dina(n5111), .dinb(n5061), .dout(n5112));
  jor  g5053(.dina(n5058), .dinb(n5057), .dout(n5113));
  jand g5054(.dina(n5113), .dinb(n4093), .dout(n5114));
  jxor g5055(.dina(n5114), .dinb(n5112), .dout(sin12 ));
  jand g5056(.dina(n5111), .dinb(n5061), .dout(n5116));
  jand g5057(.dina(n5109), .dinb(n5077), .dout(n5117));
  jand g5058(.dina(n5110), .dinb(n5064), .dout(n5118));
  jor  g5059(.dina(n5118), .dinb(n5117), .dout(n5119));
  jand g5060(.dina(n370), .dinb(n300), .dout(n5120));
  jand g5061(.dina(n2149), .dinb(n374), .dout(n5121));
  jand g5062(.dina(n5121), .dinb(n5120), .dout(n5122));
  jand g5063(.dina(n5122), .dinb(n4237), .dout(n5123));
  jand g5064(.dina(n5123), .dinb(n415), .dout(n5124));
  jand g5065(.dina(n5124), .dinb(n294), .dout(n5125));
  jand g5066(.dina(n5125), .dinb(n3892), .dout(n5126));
  jand g5067(.dina(n446), .dinb(n276), .dout(n5127));
  jand g5068(.dina(n5127), .dinb(n1025), .dout(n5128));
  jand g5069(.dina(n5128), .dinb(n884), .dout(n5129));
  jand g5070(.dina(n570), .dinb(n137), .dout(n5130));
  jand g5071(.dina(n5130), .dinb(n5129), .dout(n5131));
  jand g5072(.dina(n3106), .dinb(n912), .dout(n5132));
  jand g5073(.dina(n5132), .dinb(n5131), .dout(n5133));
  jand g5074(.dina(n5133), .dinb(n5126), .dout(n5134));
  jnot g5075(.din(n5134), .dout(n5135));
  jand g5076(.dina(n5107), .dinb(n5083), .dout(n5136));
  jand g5077(.dina(n5108), .dinb(n5080), .dout(n5137));
  jor  g5078(.dina(n5137), .dinb(n5136), .dout(n5138));
  jor  g5079(.dina(n5096), .dinb(n5088), .dout(n5139));
  jand g5080(.dina(n5106), .dinb(n5097), .dout(n5140));
  jnot g5081(.din(n5140), .dout(n5141));
  jand g5082(.dina(n5141), .dinb(n5139), .dout(n5142));
  jnot g5083(.din(n5142), .dout(n5143));
  jand g5084(.dina(n5105), .dinb(n5100), .dout(n5144));
  jor  g5085(.dina(n5144), .dinb(n5101), .dout(n5145));
  jxor g5086(.dina(n5102), .dinb(n1480), .dout(n5146));
  jand g5087(.dina(n3825), .dinb(n1438), .dout(n5147));
  jxor g5088(.dina(n5147), .dinb(n5146), .dout(n5148));
  jor  g5089(.dina(n4215), .dinb(n3384), .dout(n5149));
  jor  g5090(.dina(n4213), .dinb(n3386), .dout(n5150));
  jor  g5091(.dina(n3837), .dinb(n3388), .dout(n5151));
  jand g5092(.dina(n5151), .dinb(n5150), .dout(n5152));
  jor  g5093(.dina(n4063), .dinb(n3390), .dout(n5153));
  jand g5094(.dina(n5153), .dinb(n5152), .dout(n5154));
  jand g5095(.dina(n5154), .dinb(n5149), .dout(n5155));
  jxor g5096(.dina(n5155), .dinb(n2051), .dout(n5156));
  jxor g5097(.dina(n5156), .dinb(n5148), .dout(n5157));
  jxor g5098(.dina(n5157), .dinb(n5145), .dout(n5158));
  jxor g5099(.dina(n5158), .dinb(n5143), .dout(n5159));
  jxor g5100(.dina(n5159), .dinb(n5138), .dout(n5160));
  jxor g5101(.dina(n5160), .dinb(n5135), .dout(n5161));
  jxor g5102(.dina(n5161), .dinb(n5119), .dout(n5162));
  jxor g5103(.dina(n5162), .dinb(n5116), .dout(n5163));
  jor  g5104(.dina(n5113), .dinb(n5112), .dout(n5164));
  jand g5105(.dina(n5164), .dinb(n4093), .dout(n5165));
  jxor g5106(.dina(n5165), .dinb(n5163), .dout(sin13 ));
  jand g5107(.dina(n5162), .dinb(n5116), .dout(n5167));
  jand g5108(.dina(n5160), .dinb(n5135), .dout(n5168));
  jand g5109(.dina(n5161), .dinb(n5119), .dout(n5169));
  jor  g5110(.dina(n5169), .dinb(n5168), .dout(n5170));
  jand g5111(.dina(n2155), .dinb(n290), .dout(n5171));
  jand g5112(.dina(n5171), .dinb(n2395), .dout(n5172));
  jand g5113(.dina(n5172), .dinb(n886), .dout(n5173));
  jand g5114(.dina(n5173), .dinb(n1196), .dout(n5174));
  jand g5115(.dina(n1096), .dinb(n162), .dout(n5175));
  jand g5116(.dina(n5175), .dinb(n5174), .dout(n5176));
  jnot g5117(.din(n1312), .dout(n5177));
  jand g5118(.dina(n717), .dinb(n430), .dout(n5178));
  jand g5119(.dina(n5178), .dinb(n3537), .dout(n5179));
  jand g5120(.dina(n488), .dinb(n415), .dout(n5180));
  jand g5121(.dina(n5180), .dinb(n5179), .dout(n5181));
  jand g5122(.dina(n5181), .dinb(n5177), .dout(n5182));
  jand g5123(.dina(n5182), .dinb(n359), .dout(n5183));
  jand g5124(.dina(n5183), .dinb(n5176), .dout(n5184));
  jnot g5125(.din(n5184), .dout(n5185));
  jand g5126(.dina(n5158), .dinb(n5143), .dout(n5186));
  jand g5127(.dina(n5159), .dinb(n5138), .dout(n5187));
  jor  g5128(.dina(n5187), .dinb(n5186), .dout(n5188));
  jand g5129(.dina(n5156), .dinb(n5148), .dout(n5189));
  jand g5130(.dina(n5157), .dinb(n5145), .dout(n5190));
  jor  g5131(.dina(n5190), .dinb(n5189), .dout(n5191));
  jand g5132(.dina(n3838), .dinb(n1438), .dout(n5192));
  jnot g5133(.din(n5192), .dout(n5193));
  jand g5134(.dina(n5102), .dinb(n1480), .dout(n5194));
  jand g5135(.dina(n5147), .dinb(n5146), .dout(n5195));
  jor  g5136(.dina(n5195), .dinb(n5194), .dout(n5196));
  jxor g5137(.dina(n5196), .dinb(n5193), .dout(n5197));
  jor  g5138(.dina(n4349), .dinb(n3384), .dout(n5198));
  jor  g5139(.dina(n4063), .dinb(n3388), .dout(n5199));
  jor  g5140(.dina(n4213), .dinb(n3390), .dout(n5200));
  jand g5141(.dina(n5200), .dinb(n5199), .dout(n5201));
  jand g5142(.dina(n5201), .dinb(n5198), .dout(n5202));
  jxor g5143(.dina(n5202), .dinb(n2051), .dout(n5203));
  jxor g5144(.dina(n5203), .dinb(n5197), .dout(n5204));
  jxor g5145(.dina(n5204), .dinb(n5191), .dout(n5205));
  jxor g5146(.dina(n5205), .dinb(n5188), .dout(n5206));
  jxor g5147(.dina(n5206), .dinb(n5185), .dout(n5207));
  jxor g5148(.dina(n5207), .dinb(n5170), .dout(n5208));
  jxor g5149(.dina(n5208), .dinb(n5167), .dout(n5209));
  jor  g5150(.dina(n5164), .dinb(n5163), .dout(n5210));
  jand g5151(.dina(n5210), .dinb(n4093), .dout(n5211));
  jxor g5152(.dina(n5211), .dinb(n5209), .dout(sin14 ));
  jand g5153(.dina(n5208), .dinb(n5167), .dout(n5213));
  jand g5154(.dina(n5206), .dinb(n5185), .dout(n5214));
  jand g5155(.dina(n5207), .dinb(n5170), .dout(n5215));
  jor  g5156(.dina(n5215), .dinb(n5214), .dout(n5216));
  jand g5157(.dina(n1095), .dinb(n1005), .dout(n5217));
  jand g5158(.dina(n5217), .dinb(n94), .dout(n5218));
  jand g5159(.dina(n5218), .dinb(n858), .dout(n5219));
  jand g5160(.dina(n2402), .dinb(n206), .dout(n5220));
  jand g5161(.dina(n2135), .dinb(n395), .dout(n5221));
  jand g5162(.dina(n5221), .dinb(n2508), .dout(n5222));
  jand g5163(.dina(n346), .dinb(n222), .dout(n5223));
  jand g5164(.dina(n5223), .dinb(n5222), .dout(n5224));
  jand g5165(.dina(n5224), .dinb(n903), .dout(n5225));
  jand g5166(.dina(n5070), .dinb(n488), .dout(n5226));
  jand g5167(.dina(n5226), .dinb(n5225), .dout(n5227));
  jand g5168(.dina(n5227), .dinb(n5220), .dout(n5228));
  jand g5169(.dina(n5228), .dinb(n5219), .dout(n5229));
  jnot g5170(.din(n5229), .dout(n5230));
  jand g5171(.dina(n5196), .dinb(n5193), .dout(n5231));
  jand g5172(.dina(n5203), .dinb(n5197), .dout(n5232));
  jor  g5173(.dina(n5232), .dinb(n5231), .dout(n5233));
  jand g5174(.dina(n4338), .dinb(n2923), .dout(n5234));
  jand g5175(.dina(n4343), .dinb(n2484), .dout(n5235));
  jor  g5176(.dina(n5235), .dinb(n5234), .dout(n5236));
  jand g5177(.dina(n4344), .dinb(n1438), .dout(n5237));
  jnot g5178(.din(n5237), .dout(n5238));
  jxor g5179(.dina(n5238), .dinb(n5236), .dout(n5239));
  jxor g5180(.dina(n5239), .dinb(n5233), .dout(n5240));
  jand g5181(.dina(n5204), .dinb(n5191), .dout(n5241));
  jand g5182(.dina(n5205), .dinb(n5188), .dout(n5242));
  jor  g5183(.dina(n5242), .dinb(n5241), .dout(n5243));
  jxor g5184(.dina(n5243), .dinb(n5240), .dout(n5244));
  jxor g5185(.dina(n5244), .dinb(n5230), .dout(n5245));
  jxor g5186(.dina(n5245), .dinb(n5216), .dout(n5246));
  jxor g5187(.dina(n5246), .dinb(n5213), .dout(n5247));
  jor  g5188(.dina(n5210), .dinb(n5209), .dout(n5248));
  jand g5189(.dina(n5248), .dinb(n4093), .dout(n5249));
  jxor g5190(.dina(n5249), .dinb(n5247), .dout(sin15 ));
  jand g5191(.dina(n5246), .dinb(n5213), .dout(n5251));
  jnot g5192(.din(n5251), .dout(n5252));
  jand g5193(.dina(n5244), .dinb(n5230), .dout(n5253));
  jnot g5194(.din(n5253), .dout(n5254));
  jnot g5195(.din(n5214), .dout(n5255));
  jnot g5196(.din(n5168), .dout(n5256));
  jnot g5197(.din(n5117), .dout(n5257));
  jnot g5198(.din(n5062), .dout(n5258));
  jnot g5199(.din(n5008), .dout(n5259));
  jnot g5200(.din(n4938), .dout(n5260));
  jnot g5201(.din(n4872), .dout(n5261));
  jnot g5202(.din(n4717), .dout(n5262));
  jnot g5203(.din(n4633), .dout(n5263));
  jnot g5204(.din(n4547), .dout(n5264));
  jnot g5205(.din(n4457), .dout(n5265));
  jnot g5206(.din(n4367), .dout(n5266));
  jnot g5207(.din(n3853), .dout(n5267));
  jxor g5208(.dina(n3852), .dinb(n324), .dout(n5268));
  jnot g5209(.din(n3968), .dout(n5269));
  jor  g5210(.dina(n5269), .dinb(n3963), .dout(n5270));
  jor  g5211(.dina(n5270), .dinb(n5268), .dout(n5271));
  jand g5212(.dina(n5271), .dinb(n5267), .dout(n5272));
  jxor g5213(.dina(n4075), .dinb(n4274), .dout(n5273));
  jxor g5214(.dina(n4088), .dinb(n5273), .dout(n5274));
  jor  g5215(.dina(n5274), .dinb(n5272), .dout(n5275));
  jand g5216(.dina(n5275), .dinb(n4097), .dout(n5276));
  jxor g5217(.dina(n4226), .dinb(n4276), .dout(n5277));
  jxor g5218(.dina(n4242), .dinb(n5277), .dout(n5278));
  jor  g5219(.dina(n5278), .dinb(n5276), .dout(n5279));
  jand g5220(.dina(n5279), .dinb(n4251), .dout(n5280));
  jxor g5221(.dina(n4357), .dinb(n4270), .dout(n5281));
  jor  g5222(.dina(n5281), .dinb(n5280), .dout(n5282));
  jand g5223(.dina(n5282), .dinb(n5266), .dout(n5283));
  jxor g5224(.dina(n4451), .dinb(n4381), .dout(n5284));
  jor  g5225(.dina(n5284), .dinb(n5283), .dout(n5285));
  jand g5226(.dina(n5285), .dinb(n5265), .dout(n5286));
  jxor g5227(.dina(n4539), .dinb(n4469), .dout(n5287));
  jor  g5228(.dina(n5287), .dinb(n5286), .dout(n5288));
  jand g5229(.dina(n5288), .dinb(n5264), .dout(n5289));
  jxor g5230(.dina(n4625), .dinb(n4563), .dout(n5290));
  jor  g5231(.dina(n5290), .dinb(n5289), .dout(n5291));
  jand g5232(.dina(n5291), .dinb(n5263), .dout(n5292));
  jxor g5233(.dina(n4709), .dinb(n4652), .dout(n5293));
  jor  g5234(.dina(n5293), .dinb(n5292), .dout(n5294));
  jand g5235(.dina(n5294), .dinb(n5262), .dout(n5295));
  jxor g5236(.dina(n4771), .dinb(n4722), .dout(n5296));
  jxor g5237(.dina(n4782), .dinb(n5296), .dout(n5297));
  jor  g5238(.dina(n5297), .dinb(n5295), .dout(n5298));
  jand g5239(.dina(n5298), .dinb(n4790), .dout(n5299));
  jxor g5240(.dina(n4864), .dinb(n4813), .dout(n5300));
  jor  g5241(.dina(n5300), .dinb(n5299), .dout(n5301));
  jand g5242(.dina(n5301), .dinb(n5261), .dout(n5302));
  jxor g5243(.dina(n4930), .dinb(n4886), .dout(n5303));
  jor  g5244(.dina(n5303), .dinb(n5302), .dout(n5304));
  jand g5245(.dina(n5304), .dinb(n5260), .dout(n5305));
  jxor g5246(.dina(n5000), .dinb(n4952), .dout(n5306));
  jor  g5247(.dina(n5306), .dinb(n5305), .dout(n5307));
  jand g5248(.dina(n5307), .dinb(n5259), .dout(n5308));
  jxor g5249(.dina(n5054), .dinb(n5016), .dout(n5309));
  jor  g5250(.dina(n5309), .dinb(n5308), .dout(n5310));
  jand g5251(.dina(n5310), .dinb(n5258), .dout(n5311));
  jxor g5252(.dina(n5109), .dinb(n5076), .dout(n5312));
  jor  g5253(.dina(n5312), .dinb(n5311), .dout(n5313));
  jand g5254(.dina(n5313), .dinb(n5257), .dout(n5314));
  jxor g5255(.dina(n5160), .dinb(n5134), .dout(n5315));
  jor  g5256(.dina(n5315), .dinb(n5314), .dout(n5316));
  jand g5257(.dina(n5316), .dinb(n5256), .dout(n5317));
  jxor g5258(.dina(n5206), .dinb(n5184), .dout(n5318));
  jor  g5259(.dina(n5318), .dinb(n5317), .dout(n5319));
  jand g5260(.dina(n5319), .dinb(n5255), .dout(n5320));
  jxor g5261(.dina(n5244), .dinb(n5229), .dout(n5321));
  jor  g5262(.dina(n5321), .dinb(n5320), .dout(n5322));
  jand g5263(.dina(n5322), .dinb(n5254), .dout(n5323));
  jand g5264(.dina(n3895), .dinb(n1035), .dout(n5324));
  jand g5265(.dina(n594), .dinb(n351), .dout(n5325));
  jand g5266(.dina(n5325), .dinb(n2743), .dout(n5326));
  jand g5267(.dina(n5326), .dinb(n229), .dout(n5327));
  jand g5268(.dina(n5327), .dinb(n435), .dout(n5328));
  jand g5269(.dina(n5122), .dinb(n188), .dout(n5329));
  jand g5270(.dina(n5329), .dinb(n5328), .dout(n5330));
  jand g5271(.dina(n5330), .dinb(n5324), .dout(n5331));
  jand g5272(.dina(n5331), .dinb(n2606), .dout(n5332));
  jxor g5273(.dina(n4213), .dinb(n3838), .dout(n5333));
  jand g5274(.dina(n5333), .dinb(n1438), .dout(n5334));
  jnot g5275(.din(n5334), .dout(n5335));
  jand g5276(.dina(n5239), .dinb(n5233), .dout(n5336));
  jand g5277(.dina(n5243), .dinb(n5240), .dout(n5337));
  jor  g5278(.dina(n5337), .dinb(n5336), .dout(n5338));
  jor  g5279(.dina(n5238), .dinb(n5236), .dout(n5339));
  jnot g5280(.din(n5236), .dout(n5340));
  jor  g5281(.dina(n5340), .dinb(n1438), .dout(n5341));
  jand g5282(.dina(n5341), .dinb(n5339), .dout(n5342));
  jor  g5283(.dina(n4063), .dinb(n2051), .dout(n5343));
  jor  g5284(.dina(n5343), .dinb(n3838), .dout(n5344));
  jand g5285(.dina(n5344), .dinb(n5342), .dout(n5345));
  jxor g5286(.dina(n5345), .dinb(n5338), .dout(n5346));
  jxor g5287(.dina(n5346), .dinb(n5335), .dout(n5347));
  jxor g5288(.dina(n5347), .dinb(n5332), .dout(n5348));
  jxor g5289(.dina(n5348), .dinb(n5323), .dout(n5349));
  jxor g5290(.dina(n5349), .dinb(n5252), .dout(n5350));
  jor  g5291(.dina(n5248), .dinb(n5247), .dout(n5351));
  jand g5292(.dina(n5351), .dinb(n4093), .dout(n5352));
  jxor g5293(.dina(n5352), .dinb(n5350), .dout(sin16 ));
  jor  g5294(.dina(n5351), .dinb(n5350), .dout(n5354));
  jand g5295(.dina(n5354), .dinb(n4093), .dout(n5355));
  jor  g5296(.dina(n5349), .dinb(n5252), .dout(n5356));
  jnot g5297(.din(n5356), .dout(n5357));
  jand g5298(.dina(n198), .dinb(n166), .dout(n5358));
  jand g5299(.dina(n5358), .dinb(n1050), .dout(n5359));
  jand g5300(.dina(n5359), .dinb(n3481), .dout(n5360));
  jand g5301(.dina(n427), .dinb(n240), .dout(n5361));
  jand g5302(.dina(n5361), .dinb(n388), .dout(n5362));
  jand g5303(.dina(n344), .dinb(n182), .dout(n5363));
  jand g5304(.dina(n5363), .dinb(n5362), .dout(n5364));
  jand g5305(.dina(n5364), .dinb(n150), .dout(n5365));
  jand g5306(.dina(n5365), .dinb(n884), .dout(n5366));
  jand g5307(.dina(n5366), .dinb(n1147), .dout(n5367));
  jand g5308(.dina(n5367), .dinb(n5360), .dout(n5368));
  jnot g5309(.din(n5368), .dout(n5369));
  jnot g5310(.din(n5332), .dout(n5370));
  jxor g5311(.dina(n5346), .dinb(n5334), .dout(n5371));
  jor  g5312(.dina(n5371), .dinb(n5370), .dout(n5372));
  jand g5313(.dina(n5245), .dinb(n5216), .dout(n5373));
  jor  g5314(.dina(n5373), .dinb(n5253), .dout(n5374));
  jand g5315(.dina(n5371), .dinb(n5370), .dout(n5375));
  jor  g5316(.dina(n5375), .dinb(n5374), .dout(n5376));
  jand g5317(.dina(n5376), .dinb(n5372), .dout(n5377));
  jxor g5318(.dina(n5377), .dinb(n5369), .dout(n5378));
  jxor g5319(.dina(n5378), .dinb(n5357), .dout(n5379));
  jxor g5320(.dina(n5379), .dinb(n5355), .dout(sin17 ));
  jand g5321(.dina(n489), .dinb(n250), .dout(n5381));
  jand g5322(.dina(n5381), .dinb(n3488), .dout(n5382));
  jand g5323(.dina(n5382), .dinb(n1365), .dout(n5383));
  jand g5324(.dina(n5383), .dinb(n849), .dout(n5384));
  jand g5325(.dina(n5384), .dinb(n1140), .dout(n5385));
  jand g5326(.dina(n329), .dinb(n182), .dout(n5386));
  jand g5327(.dina(n5386), .dinb(n3098), .dout(n5387));
  jand g5328(.dina(n3868), .dinb(n824), .dout(n5388));
  jand g5329(.dina(n5388), .dinb(n5387), .dout(n5389));
  jand g5330(.dina(n5389), .dinb(n5385), .dout(n5390));
  jand g5331(.dina(n5347), .dinb(n5332), .dout(n5391));
  jor  g5332(.dina(n5347), .dinb(n5332), .dout(n5392));
  jand g5333(.dina(n5392), .dinb(n5323), .dout(n5393));
  jor  g5334(.dina(n5393), .dinb(n5391), .dout(n5394));
  jor  g5335(.dina(n5394), .dinb(n5368), .dout(n5395));
  jxor g5336(.dina(n5377), .dinb(n5368), .dout(n5396));
  jor  g5337(.dina(n5396), .dinb(n5356), .dout(n5397));
  jand g5338(.dina(n5397), .dinb(n5395), .dout(n5398));
  jxor g5339(.dina(n5398), .dinb(n5390), .dout(n5399));
  jor  g5340(.dina(n5379), .dinb(n5354), .dout(n5400));
  jand g5341(.dina(n5400), .dinb(n4093), .dout(n5401));
  jxor g5342(.dina(n5401), .dinb(n5399), .dout(sin18 ));
  jand g5343(.dina(n5378), .dinb(n5357), .dout(n5403));
  jnot g5344(.din(n5390), .dout(n5404));
  jand g5345(.dina(n5404), .dinb(n5403), .dout(n5405));
  jor  g5346(.dina(n5390), .dinb(n5395), .dout(n5406));
  jand g5347(.dina(n5219), .dinb(n189), .dout(n5407));
  jand g5348(.dina(n4558), .dinb(n1345), .dout(n5408));
  jand g5349(.dina(n5408), .dinb(n339), .dout(n5409));
  jand g5350(.dina(n5409), .dinb(n3429), .dout(n5410));
  jand g5351(.dina(n5410), .dinb(n598), .dout(n5411));
  jand g5352(.dina(n1178), .dinb(n169), .dout(n5412));
  jand g5353(.dina(n5412), .dinb(n147), .dout(n5413));
  jand g5354(.dina(n5413), .dinb(n5411), .dout(n5414));
  jand g5355(.dina(n5414), .dinb(n5407), .dout(n5415));
  jxor g5356(.dina(n5415), .dinb(n5406), .dout(n5416));
  jxor g5357(.dina(n5416), .dinb(n5405), .dout(n5417));
  jor  g5358(.dina(n5400), .dinb(n5399), .dout(n5418));
  jand g5359(.dina(n5418), .dinb(n4093), .dout(n5419));
  jxor g5360(.dina(n5419), .dinb(n5417), .dout(sin19 ));
  jor  g5361(.dina(n5415), .dinb(n5406), .dout(n5421));
  jand g5362(.dina(n4556), .dinb(n300), .dout(n5422));
  jand g5363(.dina(n5422), .dinb(n252), .dout(n5423));
  jand g5364(.dina(n1962), .dinb(n513), .dout(n5424));
  jand g5365(.dina(n534), .dinb(n267), .dout(n5425));
  jand g5366(.dina(n5425), .dinb(n461), .dout(n5426));
  jand g5367(.dina(n5426), .dinb(n265), .dout(n5427));
  jand g5368(.dina(n5427), .dinb(n5424), .dout(n5428));
  jand g5369(.dina(n5428), .dinb(n5423), .dout(n5429));
  jand g5370(.dina(n4811), .dinb(n1250), .dout(n5430));
  jand g5371(.dina(n5430), .dinb(n5429), .dout(n5431));
  jor  g5372(.dina(n5431), .dinb(n5421), .dout(n5432));
  jor  g5373(.dina(n5390), .dinb(n5397), .dout(n5433));
  jand g5374(.dina(n5377), .dinb(n5369), .dout(n5434));
  jand g5375(.dina(n5404), .dinb(n5434), .dout(n5435));
  jxor g5376(.dina(n5415), .dinb(n5435), .dout(n5436));
  jor  g5377(.dina(n5436), .dinb(n5433), .dout(n5437));
  jand g5378(.dina(n5431), .dinb(n5421), .dout(n5438));
  jxor g5379(.dina(n5438), .dinb(n5437), .dout(n5439));
  jand g5380(.dina(n5439), .dinb(n5432), .dout(n5440));
  jor  g5381(.dina(n5418), .dinb(n5417), .dout(n5441));
  jand g5382(.dina(n5441), .dinb(n4093), .dout(n5442));
  jxor g5383(.dina(n5442), .dinb(n5440), .dout(sin20 ));
  jand g5384(.dina(n5416), .dinb(n5405), .dout(n5444));
  jnot g5385(.din(n5415), .dout(n5445));
  jand g5386(.dina(n5445), .dinb(n5435), .dout(n5446));
  jnot g5387(.din(n5431), .dout(n5447));
  jor  g5388(.dina(n5447), .dinb(n5446), .dout(n5448));
  jand g5389(.dina(n5448), .dinb(n5444), .dout(n5449));
  jand g5390(.dina(n452), .dinb(n373), .dout(n5450));
  jand g5391(.dina(n5450), .dinb(n3826), .dout(n5451));
  jand g5392(.dina(n5451), .dinb(n1474), .dout(n5452));
  jxor g5393(.dina(n5452), .dinb(n5432), .dout(n5453));
  jxor g5394(.dina(n5453), .dinb(n5449), .dout(n5454));
  jor  g5395(.dina(n5441), .dinb(n5440), .dout(n5455));
  jand g5396(.dina(n5455), .dinb(n4093), .dout(n5456));
  jxor g5397(.dina(n5456), .dinb(n5454), .dout(sin21 ));
  jand g5398(.dina(n5453), .dinb(n5449), .dout(n5458));
  jand g5399(.dina(n5447), .dinb(n5446), .dout(n5459));
  jnot g5400(.din(n5452), .dout(n5460));
  jand g5401(.dina(n5460), .dinb(n5459), .dout(n5461));
  jor  g5402(.dina(n1494), .dinb(n504), .dout(n5462));
  jor  g5403(.dina(n5462), .dinb(n5461), .dout(n5463));
  jor  g5404(.dina(n5463), .dinb(n5458), .dout(n5464));
  jor  g5405(.dina(n5452), .dinb(n5432), .dout(n5465));
  jnot g5406(.din(n5462), .dout(n5466));
  jand g5407(.dina(n5466), .dinb(n5465), .dout(n5467));
  jor  g5408(.dina(n5438), .dinb(n5437), .dout(n5468));
  jxor g5409(.dina(n5452), .dinb(n5459), .dout(n5469));
  jor  g5410(.dina(n5469), .dinb(n5468), .dout(n5470));
  jor  g5411(.dina(n5466), .dinb(n5465), .dout(n5471));
  jand g5412(.dina(n5471), .dinb(n5470), .dout(n5472));
  jor  g5413(.dina(n5472), .dinb(n5467), .dout(n5473));
  jand g5414(.dina(n5473), .dinb(n5464), .dout(n5474));
  jor  g5415(.dina(n5455), .dinb(n5454), .dout(n5475));
  jand g5416(.dina(n5475), .dinb(n4093), .dout(n5476));
  jxor g5417(.dina(n5476), .dinb(n5474), .dout(sin22 ));
  jnot g5418(.din(n72), .dout(n5478));
  jand g5419(.dina(n5478), .dinb(n49), .dout(n5479));
  jand g5420(.dina(n5479), .dinb(n71), .dout(n5480));
  jand g5421(.dina(n5462), .dinb(n5461), .dout(n5481));
  jor  g5422(.dina(n5481), .dinb(n5458), .dout(n5482));
  jand g5423(.dina(n5482), .dinb(n5463), .dout(n5483));
  jor  g5424(.dina(n5471), .dinb(n5470), .dout(n5484));
  jand g5425(.dina(n5484), .dinb(n5483), .dout(n5485));
  jand g5426(.dina(n5474), .dinb(n4093), .dout(n5486));
  jor  g5427(.dina(n5486), .dinb(n5476), .dout(n5487));
  jxor g5428(.dina(n5487), .dinb(n5485), .dout(n5488));
  jor  g5429(.dina(n5488), .dinb(n5480), .dout(sin23 ));
  jand g5430(.dina(n5487), .dinb(n5484), .dout(n5490));
  jnot g5431(.din(n5454), .dout(n5491));
  jxor g5432(.dina(n5438), .dinb(n5444), .dout(n5492));
  jor  g5433(.dina(n5492), .dinb(n5459), .dout(n5493));
  jnot g5434(.din(n5417), .dout(n5494));
  jxor g5435(.dina(n5398), .dinb(n5404), .dout(n5495));
  jnot g5436(.din(n5400), .dout(n5496));
  jand g5437(.dina(n5496), .dinb(n5495), .dout(n5497));
  jand g5438(.dina(n5497), .dinb(n5494), .dout(n5498));
  jand g5439(.dina(n5498), .dinb(n5493), .dout(n5499));
  jand g5440(.dina(n5499), .dinb(n5491), .dout(n5500));
  jand g5441(.dina(n5500), .dinb(n5483), .dout(n5501));
  jor  g5442(.dina(n5501), .dinb(n5480), .dout(n5502));
  jand g5443(.dina(n5502), .dinb(n4093), .dout(n5503));
  jor  g5444(.dina(n5503), .dinb(n5490), .dout(sin24 ));
endmodule


