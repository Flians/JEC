/*

top:
	jspl: 1960
	jspl3: 418
	jnot: 1214
	jdff: 214
	jand: 1896
	jor: 1282

Summary:
	jspl: 1960
	jspl3: 418
	jnot: 1214
	jdff: 214
	jand: 1896
	jor: 1282

The maximum logic level gap of any gate:
	top: 209
*/

module gf_max(gclk, in00, in01, in02, in03, in04, in05, in06, in07, in08, in09, in010, in011, in012, in013, in014, in015, in016, in017, in018, in019, in020, in021, in022, in023, in024, in025, in026, in027, in028, in029, in030, in031, in032, in033, in034, in035, in036, in037, in038, in039, in040, in041, in042, in043, in044, in045, in046, in047, in048, in049, in050, in051, in052, in053, in054, in055, in056, in057, in058, in059, in060, in061, in062, in063, in064, in065, in066, in067, in068, in069, in070, in071, in072, in073, in074, in075, in076, in077, in078, in079, in080, in081, in082, in083, in084, in085, in086, in087, in088, in089, in090, in091, in092, in093, in094, in095, in096, in097, in098, in099, in0100, in0101, in0102, in0103, in0104, in0105, in0106, in0107, in0108, in0109, in0110, in0111, in0112, in0113, in0114, in0115, in0116, in0117, in0118, in0119, in0120, in0121, in0122, in0123, in0124, in0125, in0126, in0127, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in1100, in1101, in1102, in1103, in1104, in1105, in1106, in1107, in1108, in1109, in1110, in1111, in1112, in1113, in1114, in1115, in1116, in1117, in1118, in1119, in1120, in1121, in1122, in1123, in1124, in1125, in1126, in1127, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, in256, in257, in258, in259, in260, in261, in262, in263, in264, in265, in266, in267, in268, in269, in270, in271, in272, in273, in274, in275, in276, in277, in278, in279, in280, in281, in282, in283, in284, in285, in286, in287, in288, in289, in290, in291, in292, in293, in294, in295, in296, in297, in298, in299, in2100, in2101, in2102, in2103, in2104, in2105, in2106, in2107, in2108, in2109, in2110, in2111, in2112, in2113, in2114, in2115, in2116, in2117, in2118, in2119, in2120, in2121, in2122, in2123, in2124, in2125, in2126, in2127, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in310, in311, in312, in313, in314, in315, in316, in317, in318, in319, in320, in321, in322, in323, in324, in325, in326, in327, in328, in329, in330, in331, in332, in333, in334, in335, in336, in337, in338, in339, in340, in341, in342, in343, in344, in345, in346, in347, in348, in349, in350, in351, in352, in353, in354, in355, in356, in357, in358, in359, in360, in361, in362, in363, in364, in365, in366, in367, in368, in369, in370, in371, in372, in373, in374, in375, in376, in377, in378, in379, in380, in381, in382, in383, in384, in385, in386, in387, in388, in389, in390, in391, in392, in393, in394, in395, in396, in397, in398, in399, in3100, in3101, in3102, in3103, in3104, in3105, in3106, in3107, in3108, in3109, in3110, in3111, in3112, in3113, in3114, in3115, in3116, in3117, in3118, in3119, in3120, in3121, in3122, in3123, in3124, in3125, in3126, in3127, result0, result1, result2, result3, result4, result5, result6, result7, result8, result9, result10, result11, result12, result13, result14, result15, result16, result17, result18, result19, result20, result21, result22, result23, result24, result25, result26, result27, result28, result29, result30, result31, result32, result33, result34, result35, result36, result37, result38, result39, result40, result41, result42, result43, result44, result45, result46, result47, result48, result49, result50, result51, result52, result53, result54, result55, result56, result57, result58, result59, result60, result61, result62, result63, result64, result65, result66, result67, result68, result69, result70, result71, result72, result73, result74, result75, result76, result77, result78, result79, result80, result81, result82, result83, result84, result85, result86, result87, result88, result89, result90, result91, result92, result93, result94, result95, result96, result97, result98, result99, result100, result101, result102, result103, result104, result105, result106, result107, result108, result109, result110, result111, result112, result113, result114, result115, result116, result117, result118, result119, result120, result121, result122, result123, result124, result125, result126, result127, address0, address1);
	input gclk;
	input in00;
	input in01;
	input in02;
	input in03;
	input in04;
	input in05;
	input in06;
	input in07;
	input in08;
	input in09;
	input in010;
	input in011;
	input in012;
	input in013;
	input in014;
	input in015;
	input in016;
	input in017;
	input in018;
	input in019;
	input in020;
	input in021;
	input in022;
	input in023;
	input in024;
	input in025;
	input in026;
	input in027;
	input in028;
	input in029;
	input in030;
	input in031;
	input in032;
	input in033;
	input in034;
	input in035;
	input in036;
	input in037;
	input in038;
	input in039;
	input in040;
	input in041;
	input in042;
	input in043;
	input in044;
	input in045;
	input in046;
	input in047;
	input in048;
	input in049;
	input in050;
	input in051;
	input in052;
	input in053;
	input in054;
	input in055;
	input in056;
	input in057;
	input in058;
	input in059;
	input in060;
	input in061;
	input in062;
	input in063;
	input in064;
	input in065;
	input in066;
	input in067;
	input in068;
	input in069;
	input in070;
	input in071;
	input in072;
	input in073;
	input in074;
	input in075;
	input in076;
	input in077;
	input in078;
	input in079;
	input in080;
	input in081;
	input in082;
	input in083;
	input in084;
	input in085;
	input in086;
	input in087;
	input in088;
	input in089;
	input in090;
	input in091;
	input in092;
	input in093;
	input in094;
	input in095;
	input in096;
	input in097;
	input in098;
	input in099;
	input in0100;
	input in0101;
	input in0102;
	input in0103;
	input in0104;
	input in0105;
	input in0106;
	input in0107;
	input in0108;
	input in0109;
	input in0110;
	input in0111;
	input in0112;
	input in0113;
	input in0114;
	input in0115;
	input in0116;
	input in0117;
	input in0118;
	input in0119;
	input in0120;
	input in0121;
	input in0122;
	input in0123;
	input in0124;
	input in0125;
	input in0126;
	input in0127;
	input in10;
	input in11;
	input in12;
	input in13;
	input in14;
	input in15;
	input in16;
	input in17;
	input in18;
	input in19;
	input in110;
	input in111;
	input in112;
	input in113;
	input in114;
	input in115;
	input in116;
	input in117;
	input in118;
	input in119;
	input in120;
	input in121;
	input in122;
	input in123;
	input in124;
	input in125;
	input in126;
	input in127;
	input in128;
	input in129;
	input in130;
	input in131;
	input in132;
	input in133;
	input in134;
	input in135;
	input in136;
	input in137;
	input in138;
	input in139;
	input in140;
	input in141;
	input in142;
	input in143;
	input in144;
	input in145;
	input in146;
	input in147;
	input in148;
	input in149;
	input in150;
	input in151;
	input in152;
	input in153;
	input in154;
	input in155;
	input in156;
	input in157;
	input in158;
	input in159;
	input in160;
	input in161;
	input in162;
	input in163;
	input in164;
	input in165;
	input in166;
	input in167;
	input in168;
	input in169;
	input in170;
	input in171;
	input in172;
	input in173;
	input in174;
	input in175;
	input in176;
	input in177;
	input in178;
	input in179;
	input in180;
	input in181;
	input in182;
	input in183;
	input in184;
	input in185;
	input in186;
	input in187;
	input in188;
	input in189;
	input in190;
	input in191;
	input in192;
	input in193;
	input in194;
	input in195;
	input in196;
	input in197;
	input in198;
	input in199;
	input in1100;
	input in1101;
	input in1102;
	input in1103;
	input in1104;
	input in1105;
	input in1106;
	input in1107;
	input in1108;
	input in1109;
	input in1110;
	input in1111;
	input in1112;
	input in1113;
	input in1114;
	input in1115;
	input in1116;
	input in1117;
	input in1118;
	input in1119;
	input in1120;
	input in1121;
	input in1122;
	input in1123;
	input in1124;
	input in1125;
	input in1126;
	input in1127;
	input in20;
	input in21;
	input in22;
	input in23;
	input in24;
	input in25;
	input in26;
	input in27;
	input in28;
	input in29;
	input in210;
	input in211;
	input in212;
	input in213;
	input in214;
	input in215;
	input in216;
	input in217;
	input in218;
	input in219;
	input in220;
	input in221;
	input in222;
	input in223;
	input in224;
	input in225;
	input in226;
	input in227;
	input in228;
	input in229;
	input in230;
	input in231;
	input in232;
	input in233;
	input in234;
	input in235;
	input in236;
	input in237;
	input in238;
	input in239;
	input in240;
	input in241;
	input in242;
	input in243;
	input in244;
	input in245;
	input in246;
	input in247;
	input in248;
	input in249;
	input in250;
	input in251;
	input in252;
	input in253;
	input in254;
	input in255;
	input in256;
	input in257;
	input in258;
	input in259;
	input in260;
	input in261;
	input in262;
	input in263;
	input in264;
	input in265;
	input in266;
	input in267;
	input in268;
	input in269;
	input in270;
	input in271;
	input in272;
	input in273;
	input in274;
	input in275;
	input in276;
	input in277;
	input in278;
	input in279;
	input in280;
	input in281;
	input in282;
	input in283;
	input in284;
	input in285;
	input in286;
	input in287;
	input in288;
	input in289;
	input in290;
	input in291;
	input in292;
	input in293;
	input in294;
	input in295;
	input in296;
	input in297;
	input in298;
	input in299;
	input in2100;
	input in2101;
	input in2102;
	input in2103;
	input in2104;
	input in2105;
	input in2106;
	input in2107;
	input in2108;
	input in2109;
	input in2110;
	input in2111;
	input in2112;
	input in2113;
	input in2114;
	input in2115;
	input in2116;
	input in2117;
	input in2118;
	input in2119;
	input in2120;
	input in2121;
	input in2122;
	input in2123;
	input in2124;
	input in2125;
	input in2126;
	input in2127;
	input in30;
	input in31;
	input in32;
	input in33;
	input in34;
	input in35;
	input in36;
	input in37;
	input in38;
	input in39;
	input in310;
	input in311;
	input in312;
	input in313;
	input in314;
	input in315;
	input in316;
	input in317;
	input in318;
	input in319;
	input in320;
	input in321;
	input in322;
	input in323;
	input in324;
	input in325;
	input in326;
	input in327;
	input in328;
	input in329;
	input in330;
	input in331;
	input in332;
	input in333;
	input in334;
	input in335;
	input in336;
	input in337;
	input in338;
	input in339;
	input in340;
	input in341;
	input in342;
	input in343;
	input in344;
	input in345;
	input in346;
	input in347;
	input in348;
	input in349;
	input in350;
	input in351;
	input in352;
	input in353;
	input in354;
	input in355;
	input in356;
	input in357;
	input in358;
	input in359;
	input in360;
	input in361;
	input in362;
	input in363;
	input in364;
	input in365;
	input in366;
	input in367;
	input in368;
	input in369;
	input in370;
	input in371;
	input in372;
	input in373;
	input in374;
	input in375;
	input in376;
	input in377;
	input in378;
	input in379;
	input in380;
	input in381;
	input in382;
	input in383;
	input in384;
	input in385;
	input in386;
	input in387;
	input in388;
	input in389;
	input in390;
	input in391;
	input in392;
	input in393;
	input in394;
	input in395;
	input in396;
	input in397;
	input in398;
	input in399;
	input in3100;
	input in3101;
	input in3102;
	input in3103;
	input in3104;
	input in3105;
	input in3106;
	input in3107;
	input in3108;
	input in3109;
	input in3110;
	input in3111;
	input in3112;
	input in3113;
	input in3114;
	input in3115;
	input in3116;
	input in3117;
	input in3118;
	input in3119;
	input in3120;
	input in3121;
	input in3122;
	input in3123;
	input in3124;
	input in3125;
	input in3126;
	input in3127;
	output result0;
	output result1;
	output result2;
	output result3;
	output result4;
	output result5;
	output result6;
	output result7;
	output result8;
	output result9;
	output result10;
	output result11;
	output result12;
	output result13;
	output result14;
	output result15;
	output result16;
	output result17;
	output result18;
	output result19;
	output result20;
	output result21;
	output result22;
	output result23;
	output result24;
	output result25;
	output result26;
	output result27;
	output result28;
	output result29;
	output result30;
	output result31;
	output result32;
	output result33;
	output result34;
	output result35;
	output result36;
	output result37;
	output result38;
	output result39;
	output result40;
	output result41;
	output result42;
	output result43;
	output result44;
	output result45;
	output result46;
	output result47;
	output result48;
	output result49;
	output result50;
	output result51;
	output result52;
	output result53;
	output result54;
	output result55;
	output result56;
	output result57;
	output result58;
	output result59;
	output result60;
	output result61;
	output result62;
	output result63;
	output result64;
	output result65;
	output result66;
	output result67;
	output result68;
	output result69;
	output result70;
	output result71;
	output result72;
	output result73;
	output result74;
	output result75;
	output result76;
	output result77;
	output result78;
	output result79;
	output result80;
	output result81;
	output result82;
	output result83;
	output result84;
	output result85;
	output result86;
	output result87;
	output result88;
	output result89;
	output result90;
	output result91;
	output result92;
	output result93;
	output result94;
	output result95;
	output result96;
	output result97;
	output result98;
	output result99;
	output result100;
	output result101;
	output result102;
	output result103;
	output result104;
	output result105;
	output result106;
	output result107;
	output result108;
	output result109;
	output result110;
	output result111;
	output result112;
	output result113;
	output result114;
	output result115;
	output result116;
	output result117;
	output result118;
	output result119;
	output result120;
	output result121;
	output result122;
	output result123;
	output result124;
	output result125;
	output result126;
	output result127;
	output address0;
	output address1;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1903;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1921;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1976;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1994;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2006;
	wire n2007;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2011;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2049;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2067;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2102;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2122;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2140;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2195;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2204;
	wire n2205;
	wire n2206;
	wire n2207;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2213;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2230;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2237;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2247;
	wire n2248;
	wire n2249;
	wire n2250;
	wire n2251;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2264;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2268;
	wire n2269;
	wire n2270;
	wire n2271;
	wire n2272;
	wire n2273;
	wire n2274;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2281;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2298;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2315;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2332;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2341;
	wire n2342;
	wire n2343;
	wire n2344;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2349;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2366;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2383;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2400;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2414;
	wire n2415;
	wire n2416;
	wire n2417;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2421;
	wire n2422;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2426;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2431;
	wire n2432;
	wire n2433;
	wire n2434;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2448;
	wire n2449;
	wire n2450;
	wire n2451;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2465;
	wire n2466;
	wire n2467;
	wire n2468;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2482;
	wire n2483;
	wire n2484;
	wire n2485;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2499;
	wire n2500;
	wire n2501;
	wire n2502;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2516;
	wire n2517;
	wire n2518;
	wire n2519;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2533;
	wire n2534;
	wire n2535;
	wire n2536;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2550;
	wire n2551;
	wire n2552;
	wire n2553;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2562;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2567;
	wire n2568;
	wire n2569;
	wire n2570;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2584;
	wire n2585;
	wire n2586;
	wire n2587;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2601;
	wire n2602;
	wire n2603;
	wire n2604;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2618;
	wire n2619;
	wire n2620;
	wire n2621;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2631;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2635;
	wire n2636;
	wire n2637;
	wire n2638;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2652;
	wire n2653;
	wire n2654;
	wire n2655;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2669;
	wire n2670;
	wire n2671;
	wire n2672;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2686;
	wire n2687;
	wire n2688;
	wire n2689;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2703;
	wire n2704;
	wire n2705;
	wire n2706;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2718;
	wire n2719;
	wire n2720;
	wire n2721;
	wire n2722;
	wire n2723;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2731;
	wire n2732;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2737;
	wire n2738;
	wire n2739;
	wire n2740;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2745;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2754;
	wire n2755;
	wire n2756;
	wire n2757;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2771;
	wire n2772;
	wire n2773;
	wire n2774;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2788;
	wire n2789;
	wire n2790;
	wire n2791;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2805;
	wire n2806;
	wire n2807;
	wire n2808;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2822;
	wire n2823;
	wire n2824;
	wire n2825;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2832;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2839;
	wire n2840;
	wire n2841;
	wire n2842;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2856;
	wire n2857;
	wire n2858;
	wire n2859;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2871;
	wire n2872;
	wire n2873;
	wire n2874;
	wire n2875;
	wire n2876;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2890;
	wire n2891;
	wire n2892;
	wire n2893;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2907;
	wire n2908;
	wire n2909;
	wire n2910;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2924;
	wire n2925;
	wire n2926;
	wire n2927;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2941;
	wire n2942;
	wire n2943;
	wire n2944;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2958;
	wire n2959;
	wire n2960;
	wire n2961;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2975;
	wire n2976;
	wire n2977;
	wire n2978;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2992;
	wire n2993;
	wire n2994;
	wire n2995;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3009;
	wire n3010;
	wire n3011;
	wire n3012;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3026;
	wire n3027;
	wire n3028;
	wire n3029;
	wire n3030;
	wire n3031;
	wire n3032;
	wire n3033;
	wire n3034;
	wire n3035;
	wire n3036;
	wire n3037;
	wire n3038;
	wire n3039;
	wire n3040;
	wire n3041;
	wire n3042;
	wire n3043;
	wire n3044;
	wire n3045;
	wire n3046;
	wire n3047;
	wire n3048;
	wire n3049;
	wire n3050;
	wire n3051;
	wire n3052;
	wire n3053;
	wire n3054;
	wire n3055;
	wire n3056;
	wire n3057;
	wire n3058;
	wire n3059;
	wire n3060;
	wire n3061;
	wire n3062;
	wire n3063;
	wire n3064;
	wire n3065;
	wire n3066;
	wire n3067;
	wire n3068;
	wire n3069;
	wire n3070;
	wire n3071;
	wire n3072;
	wire n3073;
	wire n3074;
	wire n3075;
	wire n3076;
	wire n3077;
	wire n3078;
	wire n3079;
	wire n3080;
	wire n3081;
	wire n3082;
	wire n3083;
	wire n3084;
	wire n3085;
	wire n3086;
	wire n3087;
	wire n3088;
	wire n3089;
	wire n3090;
	wire n3091;
	wire n3092;
	wire n3093;
	wire n3094;
	wire n3095;
	wire n3096;
	wire n3097;
	wire n3098;
	wire n3099;
	wire n3100;
	wire n3101;
	wire n3102;
	wire n3103;
	wire n3104;
	wire n3105;
	wire n3106;
	wire n3107;
	wire n3108;
	wire n3109;
	wire n3110;
	wire n3111;
	wire n3112;
	wire n3113;
	wire n3114;
	wire n3115;
	wire n3116;
	wire n3117;
	wire n3118;
	wire n3119;
	wire n3120;
	wire n3121;
	wire n3122;
	wire n3123;
	wire n3124;
	wire n3125;
	wire n3126;
	wire n3127;
	wire n3128;
	wire n3129;
	wire n3130;
	wire n3131;
	wire n3132;
	wire n3133;
	wire n3134;
	wire n3135;
	wire n3136;
	wire n3137;
	wire n3138;
	wire n3139;
	wire n3140;
	wire n3141;
	wire n3142;
	wire n3143;
	wire n3144;
	wire n3145;
	wire n3146;
	wire n3147;
	wire n3148;
	wire n3149;
	wire n3150;
	wire n3151;
	wire n3152;
	wire n3153;
	wire n3154;
	wire n3155;
	wire n3156;
	wire n3157;
	wire n3158;
	wire n3159;
	wire n3160;
	wire n3161;
	wire n3162;
	wire n3163;
	wire n3164;
	wire n3165;
	wire n3166;
	wire n3167;
	wire n3168;
	wire n3169;
	wire n3170;
	wire n3171;
	wire n3172;
	wire n3173;
	wire n3174;
	wire n3175;
	wire n3176;
	wire n3177;
	wire n3178;
	wire n3179;
	wire n3180;
	wire n3181;
	wire n3182;
	wire n3183;
	wire n3184;
	wire n3185;
	wire n3186;
	wire n3187;
	wire n3188;
	wire n3189;
	wire n3190;
	wire n3191;
	wire n3192;
	wire n3193;
	wire n3194;
	wire n3195;
	wire n3196;
	wire n3197;
	wire n3198;
	wire n3199;
	wire n3200;
	wire n3201;
	wire n3202;
	wire n3203;
	wire n3204;
	wire n3205;
	wire n3206;
	wire n3207;
	wire n3208;
	wire n3209;
	wire n3210;
	wire n3211;
	wire n3212;
	wire n3213;
	wire n3214;
	wire n3215;
	wire n3216;
	wire n3217;
	wire n3218;
	wire n3219;
	wire n3220;
	wire n3221;
	wire n3222;
	wire n3223;
	wire n3224;
	wire n3225;
	wire n3226;
	wire n3227;
	wire n3228;
	wire n3229;
	wire n3230;
	wire n3231;
	wire n3232;
	wire n3233;
	wire n3234;
	wire n3235;
	wire n3236;
	wire n3237;
	wire n3238;
	wire n3239;
	wire n3240;
	wire n3241;
	wire n3242;
	wire n3243;
	wire n3244;
	wire n3245;
	wire n3246;
	wire n3247;
	wire n3248;
	wire n3249;
	wire n3250;
	wire n3251;
	wire n3252;
	wire n3253;
	wire n3254;
	wire n3255;
	wire n3256;
	wire n3257;
	wire n3258;
	wire n3259;
	wire n3260;
	wire n3261;
	wire n3262;
	wire n3263;
	wire n3264;
	wire n3265;
	wire n3266;
	wire n3267;
	wire n3268;
	wire n3269;
	wire n3270;
	wire n3271;
	wire n3272;
	wire n3273;
	wire n3274;
	wire n3275;
	wire n3276;
	wire n3277;
	wire n3278;
	wire n3279;
	wire n3280;
	wire n3281;
	wire n3282;
	wire n3283;
	wire n3284;
	wire n3285;
	wire n3286;
	wire n3287;
	wire n3288;
	wire n3289;
	wire n3290;
	wire n3291;
	wire n3292;
	wire n3293;
	wire n3294;
	wire n3295;
	wire n3296;
	wire n3297;
	wire n3298;
	wire n3299;
	wire n3300;
	wire n3301;
	wire n3302;
	wire n3303;
	wire n3304;
	wire n3305;
	wire n3306;
	wire n3307;
	wire n3308;
	wire n3309;
	wire n3310;
	wire n3311;
	wire n3312;
	wire n3313;
	wire n3314;
	wire n3315;
	wire n3316;
	wire n3317;
	wire n3318;
	wire n3319;
	wire n3320;
	wire n3321;
	wire n3322;
	wire n3323;
	wire n3324;
	wire n3325;
	wire n3326;
	wire n3327;
	wire n3328;
	wire n3329;
	wire n3330;
	wire n3331;
	wire n3332;
	wire n3333;
	wire n3334;
	wire n3335;
	wire n3336;
	wire n3337;
	wire n3338;
	wire n3339;
	wire n3340;
	wire n3341;
	wire n3342;
	wire n3343;
	wire n3344;
	wire n3345;
	wire n3346;
	wire n3347;
	wire n3348;
	wire n3349;
	wire n3350;
	wire n3351;
	wire n3352;
	wire n3353;
	wire n3354;
	wire n3355;
	wire n3356;
	wire n3357;
	wire n3358;
	wire n3359;
	wire n3360;
	wire n3361;
	wire n3362;
	wire n3363;
	wire n3364;
	wire n3365;
	wire n3366;
	wire n3367;
	wire n3368;
	wire n3369;
	wire n3370;
	wire n3371;
	wire n3372;
	wire n3373;
	wire n3374;
	wire n3375;
	wire n3376;
	wire n3377;
	wire n3378;
	wire n3379;
	wire n3380;
	wire n3381;
	wire n3382;
	wire n3383;
	wire n3384;
	wire n3385;
	wire n3386;
	wire n3387;
	wire n3388;
	wire n3389;
	wire n3390;
	wire n3391;
	wire n3392;
	wire n3393;
	wire n3394;
	wire n3395;
	wire n3396;
	wire n3397;
	wire n3398;
	wire n3399;
	wire n3400;
	wire n3401;
	wire n3402;
	wire n3403;
	wire n3404;
	wire n3405;
	wire n3406;
	wire n3407;
	wire n3408;
	wire n3409;
	wire n3410;
	wire n3411;
	wire n3412;
	wire n3413;
	wire n3414;
	wire n3415;
	wire n3416;
	wire n3417;
	wire n3418;
	wire n3419;
	wire n3420;
	wire n3421;
	wire n3422;
	wire n3423;
	wire n3424;
	wire n3425;
	wire n3426;
	wire n3427;
	wire n3428;
	wire n3429;
	wire n3430;
	wire n3431;
	wire n3432;
	wire n3433;
	wire n3434;
	wire n3435;
	wire n3436;
	wire n3437;
	wire n3438;
	wire n3439;
	wire n3440;
	wire n3441;
	wire n3442;
	wire n3443;
	wire n3444;
	wire n3445;
	wire n3446;
	wire n3447;
	wire n3448;
	wire n3449;
	wire n3450;
	wire n3451;
	wire n3452;
	wire n3453;
	wire n3454;
	wire n3455;
	wire n3456;
	wire n3457;
	wire n3458;
	wire n3459;
	wire n3460;
	wire n3461;
	wire n3462;
	wire n3463;
	wire n3464;
	wire n3465;
	wire n3466;
	wire n3467;
	wire n3468;
	wire n3469;
	wire n3470;
	wire n3471;
	wire n3472;
	wire n3473;
	wire n3474;
	wire n3475;
	wire n3476;
	wire n3477;
	wire n3478;
	wire n3479;
	wire n3480;
	wire n3481;
	wire n3482;
	wire n3483;
	wire n3484;
	wire n3485;
	wire n3486;
	wire n3487;
	wire n3488;
	wire n3489;
	wire n3490;
	wire n3491;
	wire n3492;
	wire n3493;
	wire n3494;
	wire n3495;
	wire n3496;
	wire n3497;
	wire n3498;
	wire n3499;
	wire n3500;
	wire n3501;
	wire n3502;
	wire n3503;
	wire n3504;
	wire n3505;
	wire n3506;
	wire n3507;
	wire n3508;
	wire n3509;
	wire n3510;
	wire n3511;
	wire n3512;
	wire n3513;
	wire n3514;
	wire n3515;
	wire n3516;
	wire n3517;
	wire n3518;
	wire n3519;
	wire n3520;
	wire n3521;
	wire n3522;
	wire n3523;
	wire n3524;
	wire n3525;
	wire n3526;
	wire n3527;
	wire n3528;
	wire n3529;
	wire n3530;
	wire n3531;
	wire n3532;
	wire n3533;
	wire n3534;
	wire n3535;
	wire n3536;
	wire n3537;
	wire n3538;
	wire n3539;
	wire n3540;
	wire n3541;
	wire n3542;
	wire n3543;
	wire n3544;
	wire n3545;
	wire n3546;
	wire n3547;
	wire n3548;
	wire n3549;
	wire n3550;
	wire n3551;
	wire n3552;
	wire n3553;
	wire n3554;
	wire n3555;
	wire n3556;
	wire n3557;
	wire n3558;
	wire n3559;
	wire n3560;
	wire n3561;
	wire n3562;
	wire n3563;
	wire n3564;
	wire n3565;
	wire n3566;
	wire n3567;
	wire n3568;
	wire n3569;
	wire n3570;
	wire n3571;
	wire n3572;
	wire n3573;
	wire n3574;
	wire n3575;
	wire n3576;
	wire n3577;
	wire n3578;
	wire n3579;
	wire n3580;
	wire n3581;
	wire n3582;
	wire n3583;
	wire n3584;
	wire n3585;
	wire n3586;
	wire n3587;
	wire n3588;
	wire n3589;
	wire n3590;
	wire n3591;
	wire n3592;
	wire n3593;
	wire n3594;
	wire n3595;
	wire n3596;
	wire n3597;
	wire n3598;
	wire n3599;
	wire n3600;
	wire n3601;
	wire n3602;
	wire n3603;
	wire n3604;
	wire n3605;
	wire n3606;
	wire n3607;
	wire n3608;
	wire n3609;
	wire n3610;
	wire n3611;
	wire n3612;
	wire n3613;
	wire n3614;
	wire n3615;
	wire n3616;
	wire n3617;
	wire n3618;
	wire n3619;
	wire n3620;
	wire n3621;
	wire n3622;
	wire n3623;
	wire n3624;
	wire n3625;
	wire n3626;
	wire n3627;
	wire n3628;
	wire n3629;
	wire n3630;
	wire n3631;
	wire n3632;
	wire n3633;
	wire n3634;
	wire n3635;
	wire n3636;
	wire n3637;
	wire n3638;
	wire n3639;
	wire n3640;
	wire n3641;
	wire n3642;
	wire n3643;
	wire n3644;
	wire n3645;
	wire n3646;
	wire n3647;
	wire n3648;
	wire n3649;
	wire n3650;
	wire n3651;
	wire n3652;
	wire n3653;
	wire n3654;
	wire n3655;
	wire n3656;
	wire n3657;
	wire n3658;
	wire n3659;
	wire n3660;
	wire n3661;
	wire n3662;
	wire n3663;
	wire n3664;
	wire n3665;
	wire n3666;
	wire n3667;
	wire n3668;
	wire n3669;
	wire n3670;
	wire n3671;
	wire n3672;
	wire n3673;
	wire n3674;
	wire n3675;
	wire n3676;
	wire n3677;
	wire n3678;
	wire n3679;
	wire n3680;
	wire n3681;
	wire n3682;
	wire n3683;
	wire n3684;
	wire n3685;
	wire n3686;
	wire n3687;
	wire n3688;
	wire n3689;
	wire n3690;
	wire n3691;
	wire n3692;
	wire n3693;
	wire n3694;
	wire n3695;
	wire n3696;
	wire n3697;
	wire n3698;
	wire n3699;
	wire n3700;
	wire n3701;
	wire n3702;
	wire n3703;
	wire n3704;
	wire n3705;
	wire n3706;
	wire n3707;
	wire n3708;
	wire n3709;
	wire n3710;
	wire n3711;
	wire n3712;
	wire n3713;
	wire n3714;
	wire n3715;
	wire n3716;
	wire n3717;
	wire n3718;
	wire n3719;
	wire n3720;
	wire n3721;
	wire n3722;
	wire n3723;
	wire n3724;
	wire n3725;
	wire n3726;
	wire n3727;
	wire n3728;
	wire n3729;
	wire n3730;
	wire n3731;
	wire n3732;
	wire n3733;
	wire n3734;
	wire n3735;
	wire n3736;
	wire n3737;
	wire n3738;
	wire n3739;
	wire n3740;
	wire n3741;
	wire n3742;
	wire n3743;
	wire n3744;
	wire n3745;
	wire n3746;
	wire n3747;
	wire n3748;
	wire n3749;
	wire n3750;
	wire n3751;
	wire n3752;
	wire n3753;
	wire n3754;
	wire n3755;
	wire n3756;
	wire n3757;
	wire n3758;
	wire n3759;
	wire n3760;
	wire n3761;
	wire n3762;
	wire n3763;
	wire n3764;
	wire n3765;
	wire n3766;
	wire n3767;
	wire n3768;
	wire n3769;
	wire n3770;
	wire n3771;
	wire n3772;
	wire n3773;
	wire n3774;
	wire n3775;
	wire n3776;
	wire n3777;
	wire n3778;
	wire n3779;
	wire n3780;
	wire n3781;
	wire n3782;
	wire n3783;
	wire n3784;
	wire n3785;
	wire n3786;
	wire n3787;
	wire n3788;
	wire n3789;
	wire n3790;
	wire n3791;
	wire n3792;
	wire n3793;
	wire n3794;
	wire n3795;
	wire n3796;
	wire n3797;
	wire n3798;
	wire n3799;
	wire n3800;
	wire n3801;
	wire n3802;
	wire n3803;
	wire n3804;
	wire n3805;
	wire n3806;
	wire n3807;
	wire n3808;
	wire n3809;
	wire n3810;
	wire n3811;
	wire n3812;
	wire n3813;
	wire n3814;
	wire n3815;
	wire n3816;
	wire n3817;
	wire n3818;
	wire n3819;
	wire n3820;
	wire n3821;
	wire n3822;
	wire n3823;
	wire n3824;
	wire n3825;
	wire n3826;
	wire n3827;
	wire n3828;
	wire n3829;
	wire n3830;
	wire n3831;
	wire n3832;
	wire n3833;
	wire n3834;
	wire n3835;
	wire n3836;
	wire n3837;
	wire n3838;
	wire n3839;
	wire n3840;
	wire n3841;
	wire n3842;
	wire n3843;
	wire n3844;
	wire n3845;
	wire n3846;
	wire n3847;
	wire n3848;
	wire n3849;
	wire n3850;
	wire n3851;
	wire n3852;
	wire n3853;
	wire n3854;
	wire n3855;
	wire n3856;
	wire n3857;
	wire n3858;
	wire n3859;
	wire n3860;
	wire n3861;
	wire n3862;
	wire n3863;
	wire n3864;
	wire n3865;
	wire n3866;
	wire n3867;
	wire n3868;
	wire n3869;
	wire n3870;
	wire n3871;
	wire n3872;
	wire n3873;
	wire n3874;
	wire n3875;
	wire n3876;
	wire n3877;
	wire n3878;
	wire n3879;
	wire n3880;
	wire n3881;
	wire n3882;
	wire n3883;
	wire n3884;
	wire n3885;
	wire n3886;
	wire n3887;
	wire n3888;
	wire n3889;
	wire n3890;
	wire n3891;
	wire n3892;
	wire n3893;
	wire n3894;
	wire n3895;
	wire n3896;
	wire n3897;
	wire n3898;
	wire n3899;
	wire n3900;
	wire n3901;
	wire n3902;
	wire n3903;
	wire n3904;
	wire n3905;
	wire n3906;
	wire n3907;
	wire n3908;
	wire n3909;
	wire n3910;
	wire n3911;
	wire n3912;
	wire n3913;
	wire n3914;
	wire n3915;
	wire n3916;
	wire n3917;
	wire n3918;
	wire n3919;
	wire n3920;
	wire n3921;
	wire n3922;
	wire n3923;
	wire n3924;
	wire n3925;
	wire n3926;
	wire n3927;
	wire n3928;
	wire n3929;
	wire n3930;
	wire n3931;
	wire n3932;
	wire n3933;
	wire n3934;
	wire n3935;
	wire n3936;
	wire n3937;
	wire n3938;
	wire n3939;
	wire n3940;
	wire n3941;
	wire n3942;
	wire n3943;
	wire n3944;
	wire n3945;
	wire n3946;
	wire n3947;
	wire n3948;
	wire n3949;
	wire n3950;
	wire n3951;
	wire n3952;
	wire n3953;
	wire n3954;
	wire n3955;
	wire n3956;
	wire n3957;
	wire n3958;
	wire n3959;
	wire n3960;
	wire n3961;
	wire n3962;
	wire n3963;
	wire n3964;
	wire n3965;
	wire n3966;
	wire n3967;
	wire n3968;
	wire n3969;
	wire n3970;
	wire n3971;
	wire n3972;
	wire n3973;
	wire n3974;
	wire n3975;
	wire n3976;
	wire n3977;
	wire n3978;
	wire n3979;
	wire n3980;
	wire n3981;
	wire n3982;
	wire n3983;
	wire n3984;
	wire n3985;
	wire n3986;
	wire n3987;
	wire n3988;
	wire n3989;
	wire n3990;
	wire n3991;
	wire n3992;
	wire n3993;
	wire n3994;
	wire n3995;
	wire n3996;
	wire n3997;
	wire n3998;
	wire n3999;
	wire n4000;
	wire n4001;
	wire n4002;
	wire n4003;
	wire n4004;
	wire n4005;
	wire n4006;
	wire n4007;
	wire n4008;
	wire n4009;
	wire n4010;
	wire n4011;
	wire n4012;
	wire n4013;
	wire n4014;
	wire n4015;
	wire n4016;
	wire n4017;
	wire n4018;
	wire n4019;
	wire n4020;
	wire n4021;
	wire n4022;
	wire n4023;
	wire n4024;
	wire n4025;
	wire n4026;
	wire n4027;
	wire n4028;
	wire n4029;
	wire n4030;
	wire n4031;
	wire n4032;
	wire n4033;
	wire n4034;
	wire n4035;
	wire n4036;
	wire n4037;
	wire n4038;
	wire n4039;
	wire n4040;
	wire n4041;
	wire n4042;
	wire n4043;
	wire n4044;
	wire n4045;
	wire n4046;
	wire n4047;
	wire n4048;
	wire n4049;
	wire n4050;
	wire n4051;
	wire n4052;
	wire n4053;
	wire n4054;
	wire n4055;
	wire n4056;
	wire n4057;
	wire n4058;
	wire n4059;
	wire n4060;
	wire n4061;
	wire n4062;
	wire n4063;
	wire n4064;
	wire n4065;
	wire n4066;
	wire n4067;
	wire n4068;
	wire n4069;
	wire n4070;
	wire n4071;
	wire n4072;
	wire n4073;
	wire n4074;
	wire n4075;
	wire n4076;
	wire n4077;
	wire n4078;
	wire n4079;
	wire n4080;
	wire n4081;
	wire n4082;
	wire n4083;
	wire n4084;
	wire n4085;
	wire n4086;
	wire n4087;
	wire n4088;
	wire n4089;
	wire n4090;
	wire n4091;
	wire n4092;
	wire n4093;
	wire n4094;
	wire n4095;
	wire n4096;
	wire n4097;
	wire n4098;
	wire n4099;
	wire n4100;
	wire n4101;
	wire n4102;
	wire n4103;
	wire n4104;
	wire n4105;
	wire n4106;
	wire n4107;
	wire n4108;
	wire n4109;
	wire n4110;
	wire n4111;
	wire n4112;
	wire n4113;
	wire n4114;
	wire n4115;
	wire n4116;
	wire n4117;
	wire n4118;
	wire n4119;
	wire n4120;
	wire n4121;
	wire n4122;
	wire n4123;
	wire n4124;
	wire n4125;
	wire n4126;
	wire n4127;
	wire n4128;
	wire n4129;
	wire n4130;
	wire n4131;
	wire n4132;
	wire n4133;
	wire n4134;
	wire n4135;
	wire n4136;
	wire n4137;
	wire n4138;
	wire n4139;
	wire n4140;
	wire n4141;
	wire n4142;
	wire n4143;
	wire n4144;
	wire n4145;
	wire n4146;
	wire n4147;
	wire n4148;
	wire n4149;
	wire n4150;
	wire n4151;
	wire n4152;
	wire n4153;
	wire n4154;
	wire n4155;
	wire n4156;
	wire n4157;
	wire n4158;
	wire n4159;
	wire n4160;
	wire n4161;
	wire n4162;
	wire n4163;
	wire n4164;
	wire n4165;
	wire n4166;
	wire n4167;
	wire n4168;
	wire n4169;
	wire n4170;
	wire n4171;
	wire n4172;
	wire n4173;
	wire n4174;
	wire n4175;
	wire n4176;
	wire n4177;
	wire n4178;
	wire n4179;
	wire n4180;
	wire n4181;
	wire n4182;
	wire n4183;
	wire n4184;
	wire n4185;
	wire n4186;
	wire n4187;
	wire n4188;
	wire n4189;
	wire n4190;
	wire n4191;
	wire n4192;
	wire n4193;
	wire n4194;
	wire n4195;
	wire n4196;
	wire n4197;
	wire n4198;
	wire n4199;
	wire n4200;
	wire n4201;
	wire n4202;
	wire n4203;
	wire n4204;
	wire n4205;
	wire n4206;
	wire n4207;
	wire n4208;
	wire n4209;
	wire n4210;
	wire n4211;
	wire n4212;
	wire n4213;
	wire n4214;
	wire n4215;
	wire n4216;
	wire n4217;
	wire n4218;
	wire n4219;
	wire n4220;
	wire n4221;
	wire n4222;
	wire n4223;
	wire n4224;
	wire n4225;
	wire n4226;
	wire n4227;
	wire n4228;
	wire n4229;
	wire n4230;
	wire n4231;
	wire n4232;
	wire n4233;
	wire n4234;
	wire n4235;
	wire n4236;
	wire n4237;
	wire n4238;
	wire n4239;
	wire n4240;
	wire n4241;
	wire n4242;
	wire n4243;
	wire n4244;
	wire n4245;
	wire n4246;
	wire n4247;
	wire n4248;
	wire n4249;
	wire n4250;
	wire n4251;
	wire n4252;
	wire n4253;
	wire n4254;
	wire n4255;
	wire n4256;
	wire n4257;
	wire n4258;
	wire n4259;
	wire n4260;
	wire n4261;
	wire n4262;
	wire n4263;
	wire n4264;
	wire n4265;
	wire n4266;
	wire n4267;
	wire n4268;
	wire n4269;
	wire n4270;
	wire n4271;
	wire n4272;
	wire n4273;
	wire n4274;
	wire n4275;
	wire n4276;
	wire n4277;
	wire n4278;
	wire n4279;
	wire n4280;
	wire n4281;
	wire n4282;
	wire n4283;
	wire n4284;
	wire n4285;
	wire n4286;
	wire n4287;
	wire n4288;
	wire n4289;
	wire n4290;
	wire n4291;
	wire n4292;
	wire n4293;
	wire n4294;
	wire n4295;
	wire n4296;
	wire n4297;
	wire n4298;
	wire n4299;
	wire n4300;
	wire n4301;
	wire n4302;
	wire n4303;
	wire n4304;
	wire n4305;
	wire n4306;
	wire n4307;
	wire n4308;
	wire n4309;
	wire n4310;
	wire n4311;
	wire n4312;
	wire n4313;
	wire n4314;
	wire n4315;
	wire n4316;
	wire n4317;
	wire n4318;
	wire n4319;
	wire n4320;
	wire n4321;
	wire n4322;
	wire n4323;
	wire n4324;
	wire n4325;
	wire n4326;
	wire n4327;
	wire n4328;
	wire n4329;
	wire n4330;
	wire n4331;
	wire n4332;
	wire n4333;
	wire n4334;
	wire n4335;
	wire n4336;
	wire n4337;
	wire n4338;
	wire n4339;
	wire n4340;
	wire n4341;
	wire n4342;
	wire n4343;
	wire n4344;
	wire n4345;
	wire n4346;
	wire n4347;
	wire n4348;
	wire n4349;
	wire n4350;
	wire n4351;
	wire n4352;
	wire n4353;
	wire n4354;
	wire n4355;
	wire n4356;
	wire n4357;
	wire n4358;
	wire n4359;
	wire n4360;
	wire n4361;
	wire n4362;
	wire n4363;
	wire n4364;
	wire n4365;
	wire n4366;
	wire n4367;
	wire n4368;
	wire n4369;
	wire n4370;
	wire n4371;
	wire n4372;
	wire n4373;
	wire n4374;
	wire n4375;
	wire n4376;
	wire n4377;
	wire n4378;
	wire n4379;
	wire n4380;
	wire n4381;
	wire n4382;
	wire n4383;
	wire n4384;
	wire n4385;
	wire n4386;
	wire n4387;
	wire n4388;
	wire n4389;
	wire n4390;
	wire n4391;
	wire n4392;
	wire n4393;
	wire n4394;
	wire n4395;
	wire n4396;
	wire n4397;
	wire n4398;
	wire n4399;
	wire n4400;
	wire n4401;
	wire n4402;
	wire n4403;
	wire n4404;
	wire n4405;
	wire n4406;
	wire n4407;
	wire n4408;
	wire n4409;
	wire n4410;
	wire n4411;
	wire n4412;
	wire n4413;
	wire n4414;
	wire n4415;
	wire n4416;
	wire n4417;
	wire n4418;
	wire n4419;
	wire n4420;
	wire n4421;
	wire n4422;
	wire n4423;
	wire n4424;
	wire n4425;
	wire n4426;
	wire n4427;
	wire n4428;
	wire n4429;
	wire n4430;
	wire n4431;
	wire n4432;
	wire n4433;
	wire n4434;
	wire n4435;
	wire n4436;
	wire n4437;
	wire n4438;
	wire n4439;
	wire n4440;
	wire n4441;
	wire n4442;
	wire n4443;
	wire n4444;
	wire n4445;
	wire n4446;
	wire n4447;
	wire n4448;
	wire n4449;
	wire n4450;
	wire n4451;
	wire n4452;
	wire n4453;
	wire n4454;
	wire n4455;
	wire n4456;
	wire n4457;
	wire n4458;
	wire n4459;
	wire n4460;
	wire n4461;
	wire n4462;
	wire n4463;
	wire n4464;
	wire n4465;
	wire n4466;
	wire n4467;
	wire n4468;
	wire n4469;
	wire n4470;
	wire n4471;
	wire n4472;
	wire n4473;
	wire n4474;
	wire n4475;
	wire n4477;
	wire n4478;
	wire n4479;
	wire n4480;
	wire n4481;
	wire n4482;
	wire n4483;
	wire n4484;
	wire n4485;
	wire n4486;
	wire n4487;
	wire n4488;
	wire n4489;
	wire n4490;
	wire n4491;
	wire n4492;
	wire n4493;
	wire n4494;
	wire n4495;
	wire n4496;
	wire n4497;
	wire n4498;
	wire n4499;
	wire n4500;
	wire n4501;
	wire n4502;
	wire n4503;
	wire n4504;
	wire n4505;
	wire n4506;
	wire n4507;
	wire n4508;
	wire n4509;
	wire n4510;
	wire n4511;
	wire n4512;
	wire n4513;
	wire n4514;
	wire n4515;
	wire n4516;
	wire n4517;
	wire n4518;
	wire n4519;
	wire n4520;
	wire n4521;
	wire n4522;
	wire n4523;
	wire n4524;
	wire n4525;
	wire n4526;
	wire n4527;
	wire n4528;
	wire n4529;
	wire n4530;
	wire n4531;
	wire n4532;
	wire n4533;
	wire n4534;
	wire n4535;
	wire n4536;
	wire n4537;
	wire n4538;
	wire n4539;
	wire n4540;
	wire n4541;
	wire n4542;
	wire n4543;
	wire n4544;
	wire n4545;
	wire n4546;
	wire n4547;
	wire n4548;
	wire n4549;
	wire n4550;
	wire n4551;
	wire n4552;
	wire n4553;
	wire n4554;
	wire n4555;
	wire n4556;
	wire n4557;
	wire n4558;
	wire n4559;
	wire n4560;
	wire n4561;
	wire n4562;
	wire n4563;
	wire n4564;
	wire n4565;
	wire n4566;
	wire n4567;
	wire n4568;
	wire n4569;
	wire n4570;
	wire n4571;
	wire n4572;
	wire n4573;
	wire n4574;
	wire n4575;
	wire n4576;
	wire n4577;
	wire n4578;
	wire n4579;
	wire n4580;
	wire n4581;
	wire n4582;
	wire n4583;
	wire n4584;
	wire n4585;
	wire n4586;
	wire n4587;
	wire n4588;
	wire n4589;
	wire n4590;
	wire n4591;
	wire n4592;
	wire n4593;
	wire n4594;
	wire n4595;
	wire n4596;
	wire n4597;
	wire n4598;
	wire n4599;
	wire n4600;
	wire n4601;
	wire n4602;
	wire n4603;
	wire n4604;
	wire n4605;
	wire n4606;
	wire n4607;
	wire n4608;
	wire n4609;
	wire n4610;
	wire n4611;
	wire n4612;
	wire n4613;
	wire n4614;
	wire n4615;
	wire n4616;
	wire n4617;
	wire n4618;
	wire n4619;
	wire n4620;
	wire n4621;
	wire n4622;
	wire n4623;
	wire n4624;
	wire n4625;
	wire n4626;
	wire n4627;
	wire n4628;
	wire n4629;
	wire n4630;
	wire n4631;
	wire n4632;
	wire n4633;
	wire n4634;
	wire n4635;
	wire n4636;
	wire n4637;
	wire n4638;
	wire n4639;
	wire n4640;
	wire n4641;
	wire n4642;
	wire n4643;
	wire n4644;
	wire n4645;
	wire n4646;
	wire n4647;
	wire n4648;
	wire n4649;
	wire n4651;
	wire n4652;
	wire n4654;
	wire n4655;
	wire n4657;
	wire n4658;
	wire n4660;
	wire n4661;
	wire n4663;
	wire n4664;
	wire n4666;
	wire n4667;
	wire n4669;
	wire n4670;
	wire n4672;
	wire n4673;
	wire n4675;
	wire n4676;
	wire n4678;
	wire n4679;
	wire n4681;
	wire n4682;
	wire n4684;
	wire n4685;
	wire n4687;
	wire n4688;
	wire n4690;
	wire n4691;
	wire n4693;
	wire n4694;
	wire n4696;
	wire n4697;
	wire n4699;
	wire n4700;
	wire n4702;
	wire n4703;
	wire n4705;
	wire n4706;
	wire n4708;
	wire n4709;
	wire n4711;
	wire n4712;
	wire n4714;
	wire n4715;
	wire n4717;
	wire n4718;
	wire n4720;
	wire n4721;
	wire n4723;
	wire n4724;
	wire n4726;
	wire n4727;
	wire n4729;
	wire n4730;
	wire n4732;
	wire n4733;
	wire n4735;
	wire n4736;
	wire n4738;
	wire n4739;
	wire n4741;
	wire n4742;
	wire n4744;
	wire n4745;
	wire n4747;
	wire n4748;
	wire n4750;
	wire n4751;
	wire n4753;
	wire n4754;
	wire n4756;
	wire n4757;
	wire n4759;
	wire n4760;
	wire n4762;
	wire n4763;
	wire n4765;
	wire n4766;
	wire n4768;
	wire n4769;
	wire n4771;
	wire n4772;
	wire n4774;
	wire n4775;
	wire n4777;
	wire n4778;
	wire n4779;
	wire n4781;
	wire n4782;
	wire n4784;
	wire n4785;
	wire n4787;
	wire n4788;
	wire n4790;
	wire n4791;
	wire n4793;
	wire n4794;
	wire n4796;
	wire n4797;
	wire n4799;
	wire n4800;
	wire n4802;
	wire n4803;
	wire n4805;
	wire n4806;
	wire n4808;
	wire n4809;
	wire n4811;
	wire n4812;
	wire n4814;
	wire n4815;
	wire n4817;
	wire n4818;
	wire n4820;
	wire n4821;
	wire n4823;
	wire n4824;
	wire n4826;
	wire n4827;
	wire n4829;
	wire n4830;
	wire n4832;
	wire n4833;
	wire n4835;
	wire n4836;
	wire n4838;
	wire n4839;
	wire n4841;
	wire n4842;
	wire n4844;
	wire n4845;
	wire n4847;
	wire n4848;
	wire n4850;
	wire n4851;
	wire n4853;
	wire n4854;
	wire n4856;
	wire n4857;
	wire n4859;
	wire n4860;
	wire n4862;
	wire n4863;
	wire n4865;
	wire n4866;
	wire n4868;
	wire n4869;
	wire n4871;
	wire n4872;
	wire n4874;
	wire n4875;
	wire n4877;
	wire n4878;
	wire n4880;
	wire n4881;
	wire n4883;
	wire n4884;
	wire n4886;
	wire n4887;
	wire n4889;
	wire n4890;
	wire n4892;
	wire n4893;
	wire n4895;
	wire n4896;
	wire n4898;
	wire n4899;
	wire n4901;
	wire n4902;
	wire n4904;
	wire n4905;
	wire n4907;
	wire n4908;
	wire n4910;
	wire n4911;
	wire n4913;
	wire n4914;
	wire n4916;
	wire n4917;
	wire n4919;
	wire n4920;
	wire n4922;
	wire n4923;
	wire n4925;
	wire n4926;
	wire n4928;
	wire n4929;
	wire n4931;
	wire n4932;
	wire n4934;
	wire n4935;
	wire n4937;
	wire n4938;
	wire n4940;
	wire n4941;
	wire n4943;
	wire n4944;
	wire n4946;
	wire n4947;
	wire n4949;
	wire n4950;
	wire n4952;
	wire n4953;
	wire n4955;
	wire n4956;
	wire n4958;
	wire n4959;
	wire n4961;
	wire n4962;
	wire n4964;
	wire n4965;
	wire n4967;
	wire n4968;
	wire n4970;
	wire n4971;
	wire n4973;
	wire n4974;
	wire n4976;
	wire n4977;
	wire n4979;
	wire n4980;
	wire n4982;
	wire n4983;
	wire n4985;
	wire n4986;
	wire n4988;
	wire n4989;
	wire n4991;
	wire n4992;
	wire n4994;
	wire n4995;
	wire n4997;
	wire n4998;
	wire n5000;
	wire n5001;
	wire n5003;
	wire n5004;
	wire n5006;
	wire n5007;
	wire n5009;
	wire n5010;
	wire n5012;
	wire n5013;
	wire n5015;
	wire n5016;
	wire n5018;
	wire n5019;
	wire n5021;
	wire n5022;
	wire n5024;
	wire n5025;
	wire n5027;
	wire n5028;
	wire n5031;
	wire n5032;
	wire[2:0] w_in00_0;
	wire[2:0] w_in01_0;
	wire[1:0] w_in01_1;
	wire[2:0] w_in02_0;
	wire[1:0] w_in02_1;
	wire[2:0] w_in03_0;
	wire[1:0] w_in04_0;
	wire[1:0] w_in05_0;
	wire[1:0] w_in06_0;
	wire[1:0] w_in07_0;
	wire[1:0] w_in08_0;
	wire[1:0] w_in09_0;
	wire[1:0] w_in010_0;
	wire[1:0] w_in011_0;
	wire[1:0] w_in012_0;
	wire[1:0] w_in013_0;
	wire[1:0] w_in014_0;
	wire[1:0] w_in015_0;
	wire[1:0] w_in016_0;
	wire[1:0] w_in017_0;
	wire[1:0] w_in018_0;
	wire[1:0] w_in019_0;
	wire[1:0] w_in020_0;
	wire[1:0] w_in021_0;
	wire[1:0] w_in022_0;
	wire[1:0] w_in023_0;
	wire[1:0] w_in024_0;
	wire[1:0] w_in025_0;
	wire[1:0] w_in026_0;
	wire[1:0] w_in027_0;
	wire[1:0] w_in028_0;
	wire[1:0] w_in029_0;
	wire[1:0] w_in030_0;
	wire[1:0] w_in031_0;
	wire[1:0] w_in032_0;
	wire[1:0] w_in033_0;
	wire[1:0] w_in034_0;
	wire[1:0] w_in035_0;
	wire[1:0] w_in036_0;
	wire[1:0] w_in037_0;
	wire[1:0] w_in038_0;
	wire[1:0] w_in039_0;
	wire[1:0] w_in040_0;
	wire[1:0] w_in041_0;
	wire[1:0] w_in042_0;
	wire[1:0] w_in044_0;
	wire[1:0] w_in045_0;
	wire[1:0] w_in046_0;
	wire[1:0] w_in047_0;
	wire[1:0] w_in048_0;
	wire[1:0] w_in049_0;
	wire[1:0] w_in050_0;
	wire[1:0] w_in051_0;
	wire[1:0] w_in052_0;
	wire[1:0] w_in053_0;
	wire[1:0] w_in054_0;
	wire[1:0] w_in055_0;
	wire[1:0] w_in056_0;
	wire[1:0] w_in057_0;
	wire[1:0] w_in058_0;
	wire[1:0] w_in059_0;
	wire[1:0] w_in060_0;
	wire[1:0] w_in061_0;
	wire[1:0] w_in062_0;
	wire[1:0] w_in063_0;
	wire[1:0] w_in064_0;
	wire[1:0] w_in065_0;
	wire[1:0] w_in066_0;
	wire[1:0] w_in067_0;
	wire[1:0] w_in068_0;
	wire[1:0] w_in069_0;
	wire[1:0] w_in070_0;
	wire[1:0] w_in071_0;
	wire[1:0] w_in072_0;
	wire[1:0] w_in073_0;
	wire[1:0] w_in074_0;
	wire[1:0] w_in075_0;
	wire[1:0] w_in076_0;
	wire[1:0] w_in077_0;
	wire[1:0] w_in078_0;
	wire[1:0] w_in079_0;
	wire[1:0] w_in080_0;
	wire[1:0] w_in081_0;
	wire[1:0] w_in082_0;
	wire[1:0] w_in083_0;
	wire[1:0] w_in084_0;
	wire[1:0] w_in085_0;
	wire[1:0] w_in086_0;
	wire[1:0] w_in087_0;
	wire[1:0] w_in088_0;
	wire[1:0] w_in089_0;
	wire[1:0] w_in090_0;
	wire[1:0] w_in091_0;
	wire[1:0] w_in092_0;
	wire[1:0] w_in093_0;
	wire[1:0] w_in094_0;
	wire[1:0] w_in095_0;
	wire[1:0] w_in096_0;
	wire[1:0] w_in097_0;
	wire[1:0] w_in098_0;
	wire[1:0] w_in099_0;
	wire[1:0] w_in0100_0;
	wire[1:0] w_in0101_0;
	wire[1:0] w_in0102_0;
	wire[1:0] w_in0103_0;
	wire[1:0] w_in0104_0;
	wire[1:0] w_in0105_0;
	wire[1:0] w_in0106_0;
	wire[1:0] w_in0107_0;
	wire[1:0] w_in0108_0;
	wire[1:0] w_in0109_0;
	wire[1:0] w_in0110_0;
	wire[1:0] w_in0111_0;
	wire[1:0] w_in0112_0;
	wire[1:0] w_in0113_0;
	wire[1:0] w_in0114_0;
	wire[1:0] w_in0115_0;
	wire[1:0] w_in0116_0;
	wire[1:0] w_in0117_0;
	wire[1:0] w_in0118_0;
	wire[1:0] w_in0119_0;
	wire[1:0] w_in0120_0;
	wire[1:0] w_in0121_0;
	wire[1:0] w_in0122_0;
	wire[1:0] w_in0123_0;
	wire[1:0] w_in0124_0;
	wire[1:0] w_in0125_0;
	wire[1:0] w_in0126_0;
	wire[2:0] w_in0127_0;
	wire[2:0] w_in10_0;
	wire[2:0] w_in11_0;
	wire[1:0] w_in11_1;
	wire[2:0] w_in12_0;
	wire[2:0] w_in13_0;
	wire[1:0] w_in14_0;
	wire[1:0] w_in15_0;
	wire[1:0] w_in16_0;
	wire[1:0] w_in17_0;
	wire[1:0] w_in18_0;
	wire[1:0] w_in19_0;
	wire[1:0] w_in110_0;
	wire[1:0] w_in111_0;
	wire[1:0] w_in112_0;
	wire[1:0] w_in113_0;
	wire[1:0] w_in114_0;
	wire[1:0] w_in115_0;
	wire[1:0] w_in116_0;
	wire[1:0] w_in117_0;
	wire[1:0] w_in118_0;
	wire[1:0] w_in119_0;
	wire[1:0] w_in120_0;
	wire[1:0] w_in121_0;
	wire[1:0] w_in122_0;
	wire[1:0] w_in123_0;
	wire[1:0] w_in124_0;
	wire[1:0] w_in125_0;
	wire[1:0] w_in126_0;
	wire[1:0] w_in127_0;
	wire[1:0] w_in128_0;
	wire[1:0] w_in129_0;
	wire[1:0] w_in130_0;
	wire[1:0] w_in131_0;
	wire[1:0] w_in132_0;
	wire[1:0] w_in133_0;
	wire[1:0] w_in134_0;
	wire[1:0] w_in135_0;
	wire[1:0] w_in136_0;
	wire[1:0] w_in137_0;
	wire[1:0] w_in138_0;
	wire[1:0] w_in139_0;
	wire[1:0] w_in140_0;
	wire[1:0] w_in141_0;
	wire[1:0] w_in142_0;
	wire[2:0] w_in143_0;
	wire[1:0] w_in144_0;
	wire[1:0] w_in145_0;
	wire[1:0] w_in146_0;
	wire[1:0] w_in147_0;
	wire[1:0] w_in148_0;
	wire[1:0] w_in149_0;
	wire[1:0] w_in150_0;
	wire[1:0] w_in151_0;
	wire[1:0] w_in152_0;
	wire[1:0] w_in153_0;
	wire[1:0] w_in154_0;
	wire[1:0] w_in155_0;
	wire[1:0] w_in156_0;
	wire[1:0] w_in157_0;
	wire[1:0] w_in158_0;
	wire[1:0] w_in159_0;
	wire[1:0] w_in160_0;
	wire[1:0] w_in161_0;
	wire[1:0] w_in162_0;
	wire[1:0] w_in163_0;
	wire[1:0] w_in164_0;
	wire[1:0] w_in165_0;
	wire[1:0] w_in166_0;
	wire[1:0] w_in167_0;
	wire[1:0] w_in168_0;
	wire[1:0] w_in169_0;
	wire[1:0] w_in170_0;
	wire[1:0] w_in171_0;
	wire[1:0] w_in172_0;
	wire[1:0] w_in173_0;
	wire[1:0] w_in174_0;
	wire[1:0] w_in175_0;
	wire[1:0] w_in176_0;
	wire[1:0] w_in177_0;
	wire[1:0] w_in178_0;
	wire[1:0] w_in179_0;
	wire[1:0] w_in180_0;
	wire[1:0] w_in181_0;
	wire[1:0] w_in182_0;
	wire[1:0] w_in183_0;
	wire[1:0] w_in184_0;
	wire[1:0] w_in185_0;
	wire[1:0] w_in186_0;
	wire[1:0] w_in187_0;
	wire[1:0] w_in188_0;
	wire[1:0] w_in189_0;
	wire[1:0] w_in190_0;
	wire[1:0] w_in191_0;
	wire[1:0] w_in192_0;
	wire[1:0] w_in193_0;
	wire[1:0] w_in194_0;
	wire[1:0] w_in195_0;
	wire[1:0] w_in196_0;
	wire[1:0] w_in197_0;
	wire[1:0] w_in198_0;
	wire[1:0] w_in199_0;
	wire[1:0] w_in1100_0;
	wire[1:0] w_in1101_0;
	wire[1:0] w_in1102_0;
	wire[1:0] w_in1103_0;
	wire[1:0] w_in1104_0;
	wire[1:0] w_in1105_0;
	wire[1:0] w_in1106_0;
	wire[1:0] w_in1107_0;
	wire[1:0] w_in1108_0;
	wire[1:0] w_in1109_0;
	wire[1:0] w_in1110_0;
	wire[1:0] w_in1111_0;
	wire[1:0] w_in1112_0;
	wire[1:0] w_in1113_0;
	wire[1:0] w_in1114_0;
	wire[1:0] w_in1115_0;
	wire[1:0] w_in1116_0;
	wire[1:0] w_in1117_0;
	wire[1:0] w_in1118_0;
	wire[1:0] w_in1119_0;
	wire[1:0] w_in1120_0;
	wire[1:0] w_in1121_0;
	wire[1:0] w_in1122_0;
	wire[1:0] w_in1123_0;
	wire[1:0] w_in1124_0;
	wire[1:0] w_in1125_0;
	wire[1:0] w_in1126_0;
	wire[2:0] w_in1127_0;
	wire[2:0] w_in20_0;
	wire[2:0] w_in21_0;
	wire[1:0] w_in21_1;
	wire[2:0] w_in22_0;
	wire[1:0] w_in23_0;
	wire[1:0] w_in24_0;
	wire[1:0] w_in25_0;
	wire[1:0] w_in26_0;
	wire[1:0] w_in27_0;
	wire[1:0] w_in28_0;
	wire[1:0] w_in29_0;
	wire[1:0] w_in210_0;
	wire[1:0] w_in211_0;
	wire[1:0] w_in212_0;
	wire[1:0] w_in213_0;
	wire[1:0] w_in214_0;
	wire[1:0] w_in215_0;
	wire[1:0] w_in216_0;
	wire[1:0] w_in217_0;
	wire[1:0] w_in218_0;
	wire[1:0] w_in219_0;
	wire[1:0] w_in220_0;
	wire[1:0] w_in221_0;
	wire[1:0] w_in222_0;
	wire[1:0] w_in223_0;
	wire[1:0] w_in224_0;
	wire[1:0] w_in225_0;
	wire[1:0] w_in226_0;
	wire[1:0] w_in227_0;
	wire[1:0] w_in228_0;
	wire[1:0] w_in229_0;
	wire[1:0] w_in230_0;
	wire[1:0] w_in231_0;
	wire[1:0] w_in232_0;
	wire[1:0] w_in233_0;
	wire[1:0] w_in234_0;
	wire[1:0] w_in235_0;
	wire[1:0] w_in236_0;
	wire[1:0] w_in237_0;
	wire[1:0] w_in238_0;
	wire[1:0] w_in239_0;
	wire[1:0] w_in240_0;
	wire[1:0] w_in241_0;
	wire[1:0] w_in242_0;
	wire[1:0] w_in243_0;
	wire[1:0] w_in244_0;
	wire[1:0] w_in245_0;
	wire[1:0] w_in246_0;
	wire[1:0] w_in247_0;
	wire[1:0] w_in248_0;
	wire[1:0] w_in249_0;
	wire[1:0] w_in250_0;
	wire[1:0] w_in251_0;
	wire[1:0] w_in252_0;
	wire[1:0] w_in253_0;
	wire[1:0] w_in254_0;
	wire[1:0] w_in255_0;
	wire[1:0] w_in256_0;
	wire[1:0] w_in257_0;
	wire[1:0] w_in258_0;
	wire[1:0] w_in259_0;
	wire[1:0] w_in260_0;
	wire[1:0] w_in261_0;
	wire[1:0] w_in262_0;
	wire[1:0] w_in263_0;
	wire[1:0] w_in264_0;
	wire[1:0] w_in265_0;
	wire[1:0] w_in266_0;
	wire[1:0] w_in267_0;
	wire[1:0] w_in268_0;
	wire[1:0] w_in269_0;
	wire[1:0] w_in270_0;
	wire[1:0] w_in271_0;
	wire[1:0] w_in272_0;
	wire[1:0] w_in273_0;
	wire[1:0] w_in274_0;
	wire[1:0] w_in275_0;
	wire[1:0] w_in276_0;
	wire[1:0] w_in277_0;
	wire[1:0] w_in278_0;
	wire[1:0] w_in279_0;
	wire[1:0] w_in280_0;
	wire[1:0] w_in281_0;
	wire[1:0] w_in282_0;
	wire[1:0] w_in283_0;
	wire[1:0] w_in284_0;
	wire[1:0] w_in285_0;
	wire[1:0] w_in286_0;
	wire[1:0] w_in287_0;
	wire[1:0] w_in288_0;
	wire[1:0] w_in289_0;
	wire[1:0] w_in290_0;
	wire[1:0] w_in291_0;
	wire[1:0] w_in292_0;
	wire[1:0] w_in293_0;
	wire[1:0] w_in294_0;
	wire[1:0] w_in295_0;
	wire[1:0] w_in296_0;
	wire[1:0] w_in297_0;
	wire[1:0] w_in298_0;
	wire[1:0] w_in299_0;
	wire[1:0] w_in2100_0;
	wire[1:0] w_in2101_0;
	wire[1:0] w_in2102_0;
	wire[1:0] w_in2103_0;
	wire[1:0] w_in2104_0;
	wire[1:0] w_in2105_0;
	wire[1:0] w_in2106_0;
	wire[1:0] w_in2107_0;
	wire[1:0] w_in2108_0;
	wire[1:0] w_in2109_0;
	wire[1:0] w_in2110_0;
	wire[1:0] w_in2111_0;
	wire[1:0] w_in2112_0;
	wire[1:0] w_in2113_0;
	wire[1:0] w_in2114_0;
	wire[1:0] w_in2115_0;
	wire[1:0] w_in2116_0;
	wire[1:0] w_in2117_0;
	wire[1:0] w_in2118_0;
	wire[1:0] w_in2119_0;
	wire[1:0] w_in2120_0;
	wire[1:0] w_in2121_0;
	wire[1:0] w_in2122_0;
	wire[1:0] w_in2123_0;
	wire[1:0] w_in2124_0;
	wire[1:0] w_in2125_0;
	wire[1:0] w_in2126_0;
	wire[2:0] w_in2127_0;
	wire[2:0] w_in30_0;
	wire[2:0] w_in31_0;
	wire[2:0] w_in32_0;
	wire[1:0] w_in33_0;
	wire[1:0] w_in34_0;
	wire[1:0] w_in35_0;
	wire[1:0] w_in36_0;
	wire[1:0] w_in37_0;
	wire[1:0] w_in38_0;
	wire[1:0] w_in39_0;
	wire[1:0] w_in310_0;
	wire[1:0] w_in311_0;
	wire[1:0] w_in312_0;
	wire[1:0] w_in313_0;
	wire[1:0] w_in314_0;
	wire[1:0] w_in315_0;
	wire[1:0] w_in316_0;
	wire[1:0] w_in317_0;
	wire[1:0] w_in318_0;
	wire[1:0] w_in319_0;
	wire[1:0] w_in320_0;
	wire[1:0] w_in321_0;
	wire[1:0] w_in322_0;
	wire[1:0] w_in323_0;
	wire[1:0] w_in324_0;
	wire[1:0] w_in325_0;
	wire[1:0] w_in326_0;
	wire[1:0] w_in327_0;
	wire[1:0] w_in328_0;
	wire[1:0] w_in329_0;
	wire[1:0] w_in330_0;
	wire[1:0] w_in331_0;
	wire[1:0] w_in332_0;
	wire[1:0] w_in333_0;
	wire[1:0] w_in334_0;
	wire[1:0] w_in335_0;
	wire[1:0] w_in336_0;
	wire[1:0] w_in337_0;
	wire[1:0] w_in338_0;
	wire[1:0] w_in339_0;
	wire[1:0] w_in340_0;
	wire[1:0] w_in341_0;
	wire[1:0] w_in342_0;
	wire[1:0] w_in343_0;
	wire[1:0] w_in344_0;
	wire[1:0] w_in345_0;
	wire[1:0] w_in346_0;
	wire[1:0] w_in347_0;
	wire[1:0] w_in348_0;
	wire[1:0] w_in349_0;
	wire[1:0] w_in350_0;
	wire[1:0] w_in351_0;
	wire[1:0] w_in352_0;
	wire[1:0] w_in353_0;
	wire[1:0] w_in354_0;
	wire[1:0] w_in355_0;
	wire[1:0] w_in356_0;
	wire[1:0] w_in357_0;
	wire[1:0] w_in358_0;
	wire[1:0] w_in359_0;
	wire[1:0] w_in360_0;
	wire[1:0] w_in361_0;
	wire[1:0] w_in362_0;
	wire[1:0] w_in363_0;
	wire[1:0] w_in364_0;
	wire[1:0] w_in365_0;
	wire[1:0] w_in366_0;
	wire[1:0] w_in367_0;
	wire[1:0] w_in368_0;
	wire[1:0] w_in369_0;
	wire[1:0] w_in370_0;
	wire[1:0] w_in371_0;
	wire[1:0] w_in372_0;
	wire[1:0] w_in373_0;
	wire[1:0] w_in374_0;
	wire[1:0] w_in375_0;
	wire[1:0] w_in376_0;
	wire[1:0] w_in377_0;
	wire[1:0] w_in378_0;
	wire[1:0] w_in379_0;
	wire[1:0] w_in380_0;
	wire[1:0] w_in381_0;
	wire[1:0] w_in382_0;
	wire[1:0] w_in383_0;
	wire[1:0] w_in384_0;
	wire[1:0] w_in385_0;
	wire[1:0] w_in386_0;
	wire[1:0] w_in387_0;
	wire[1:0] w_in388_0;
	wire[1:0] w_in389_0;
	wire[1:0] w_in390_0;
	wire[1:0] w_in391_0;
	wire[1:0] w_in392_0;
	wire[1:0] w_in393_0;
	wire[1:0] w_in394_0;
	wire[1:0] w_in395_0;
	wire[1:0] w_in396_0;
	wire[1:0] w_in397_0;
	wire[1:0] w_in398_0;
	wire[1:0] w_in399_0;
	wire[1:0] w_in3100_0;
	wire[1:0] w_in3101_0;
	wire[1:0] w_in3102_0;
	wire[1:0] w_in3103_0;
	wire[1:0] w_in3104_0;
	wire[1:0] w_in3105_0;
	wire[1:0] w_in3106_0;
	wire[1:0] w_in3107_0;
	wire[1:0] w_in3108_0;
	wire[1:0] w_in3109_0;
	wire[1:0] w_in3110_0;
	wire[1:0] w_in3111_0;
	wire[1:0] w_in3112_0;
	wire[1:0] w_in3113_0;
	wire[1:0] w_in3114_0;
	wire[1:0] w_in3115_0;
	wire[1:0] w_in3116_0;
	wire[1:0] w_in3117_0;
	wire[1:0] w_in3118_0;
	wire[1:0] w_in3119_0;
	wire[1:0] w_in3120_0;
	wire[1:0] w_in3121_0;
	wire[1:0] w_in3122_0;
	wire[1:0] w_in3123_0;
	wire[1:0] w_in3124_0;
	wire[1:0] w_in3125_0;
	wire[1:0] w_in3126_0;
	wire[1:0] w_in3127_0;
	wire[2:0] w_address1_0;
	wire[2:0] w_address1_1;
	wire[2:0] w_address1_2;
	wire[2:0] w_address1_3;
	wire[2:0] w_address1_4;
	wire[2:0] w_address1_5;
	wire[2:0] w_address1_6;
	wire[2:0] w_address1_7;
	wire[2:0] w_address1_8;
	wire[2:0] w_address1_9;
	wire[2:0] w_address1_10;
	wire[2:0] w_address1_11;
	wire[2:0] w_address1_12;
	wire[2:0] w_address1_13;
	wire[2:0] w_address1_14;
	wire[2:0] w_address1_15;
	wire[2:0] w_address1_16;
	wire[2:0] w_address1_17;
	wire[2:0] w_address1_18;
	wire[2:0] w_address1_19;
	wire[2:0] w_address1_20;
	wire[2:0] w_address1_21;
	wire[2:0] w_address1_22;
	wire[2:0] w_address1_23;
	wire[2:0] w_address1_24;
	wire[2:0] w_address1_25;
	wire[2:0] w_address1_26;
	wire[2:0] w_address1_27;
	wire[2:0] w_address1_28;
	wire[2:0] w_address1_29;
	wire[2:0] w_address1_30;
	wire[2:0] w_address1_31;
	wire[2:0] w_address1_32;
	wire[2:0] w_address1_33;
	wire[2:0] w_address1_34;
	wire[2:0] w_address1_35;
	wire[2:0] w_address1_36;
	wire[2:0] w_address1_37;
	wire[2:0] w_address1_38;
	wire[2:0] w_address1_39;
	wire[2:0] w_address1_40;
	wire[2:0] w_address1_41;
	wire[2:0] w_address1_42;
	wire[2:0] w_address1_43;
	wire[2:0] w_address1_44;
	wire[2:0] w_address1_45;
	wire[2:0] w_address1_46;
	wire[2:0] w_address1_47;
	wire[2:0] w_address1_48;
	wire[2:0] w_address1_49;
	wire[2:0] w_address1_50;
	wire[2:0] w_address1_51;
	wire[2:0] w_address1_52;
	wire[2:0] w_address1_53;
	wire[2:0] w_address1_54;
	wire[2:0] w_address1_55;
	wire[2:0] w_address1_56;
	wire[2:0] w_address1_57;
	wire[2:0] w_address1_58;
	wire[2:0] w_address1_59;
	wire[2:0] w_address1_60;
	wire[2:0] w_address1_61;
	wire[2:0] w_address1_62;
	wire[1:0] w_address1_63;
	wire address1_fa_;
	wire[1:0] w_n642_0;
	wire[1:0] w_n643_0;
	wire[1:0] w_n645_0;
	wire[1:0] w_n647_0;
	wire[1:0] w_n648_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n653_0;
	wire[1:0] w_n654_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n659_0;
	wire[1:0] w_n661_0;
	wire[1:0] w_n666_0;
	wire[1:0] w_n668_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n674_0;
	wire[1:0] w_n675_0;
	wire[1:0] w_n677_0;
	wire[1:0] w_n678_0;
	wire[1:0] w_n679_0;
	wire[1:0] w_n681_0;
	wire[1:0] w_n682_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n691_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n698_0;
	wire[1:0] w_n700_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n707_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[1:0] w_n713_0;
	wire[1:0] w_n714_0;
	wire[1:0] w_n716_0;
	wire[1:0] w_n717_0;
	wire[1:0] w_n718_0;
	wire[1:0] w_n721_0;
	wire[1:0] w_n723_0;
	wire[1:0] w_n725_0;
	wire[1:0] w_n730_0;
	wire[1:0] w_n732_0;
	wire[1:0] w_n736_0;
	wire[1:0] w_n738_0;
	wire[1:0] w_n739_0;
	wire[1:0] w_n741_0;
	wire[1:0] w_n742_0;
	wire[1:0] w_n743_0;
	wire[1:0] w_n745_0;
	wire[1:0] w_n746_0;
	wire[1:0] w_n748_0;
	wire[1:0] w_n749_0;
	wire[1:0] w_n750_0;
	wire[1:0] w_n753_0;
	wire[1:0] w_n755_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n762_0;
	wire[1:0] w_n764_0;
	wire[1:0] w_n768_0;
	wire[1:0] w_n770_0;
	wire[1:0] w_n771_0;
	wire[1:0] w_n773_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n776_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n780_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n784_0;
	wire[1:0] w_n789_0;
	wire[1:0] w_n791_0;
	wire[1:0] w_n795_0;
	wire[1:0] w_n797_0;
	wire[1:0] w_n798_0;
	wire[1:0] w_n800_0;
	wire[1:0] w_n801_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n804_0;
	wire[1:0] w_n805_0;
	wire[1:0] w_n807_0;
	wire[1:0] w_n808_0;
	wire[1:0] w_n809_0;
	wire[1:0] w_n812_0;
	wire[1:0] w_n814_0;
	wire[1:0] w_n816_0;
	wire[1:0] w_n821_0;
	wire[1:0] w_n823_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n829_0;
	wire[1:0] w_n830_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n834_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n836_0;
	wire[1:0] w_n837_0;
	wire[1:0] w_n839_0;
	wire[1:0] w_n840_0;
	wire[1:0] w_n841_0;
	wire[1:0] w_n844_0;
	wire[1:0] w_n846_0;
	wire[1:0] w_n848_0;
	wire[1:0] w_n853_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n861_0;
	wire[1:0] w_n862_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n865_0;
	wire[1:0] w_n867_0;
	wire[1:0] w_n870_0;
	wire[1:0] w_n872_0;
	wire[1:0] w_n875_0;
	wire[1:0] w_n877_0;
	wire[1:0] w_n878_0;
	wire[1:0] w_n880_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n882_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n887_0;
	wire[1:0] w_n888_0;
	wire[1:0] w_n891_0;
	wire[1:0] w_n893_0;
	wire[1:0] w_n894_0;
	wire[1:0] w_n895_0;
	wire[1:0] w_n896_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n900_0;
	wire[1:0] w_n901_0;
	wire[1:0] w_n904_0;
	wire[1:0] w_n907_0;
	wire[1:0] w_n909_0;
	wire[1:0] w_n911_0;
	wire[1:0] w_n912_0;
	wire[1:0] w_n913_0;
	wire[1:0] w_n915_0;
	wire[1:0] w_n918_0;
	wire[1:0] w_n919_0;
	wire[1:0] w_n920_0;
	wire[2:0] w_n922_0;
	wire[1:0] w_n925_0;
	wire[1:0] w_n927_0;
	wire[1:0] w_n929_0;
	wire[1:0] w_n931_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n934_0;
	wire[1:0] w_n939_0;
	wire[1:0] w_n941_0;
	wire[1:0] w_n943_0;
	wire[1:0] w_n946_0;
	wire[1:0] w_n947_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n953_0;
	wire[1:0] w_n955_0;
	wire[1:0] w_n958_0;
	wire[1:0] w_n960_0;
	wire[1:0] w_n962_0;
	wire[1:0] w_n963_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n967_0;
	wire[1:0] w_n968_0;
	wire[1:0] w_n969_0;
	wire[1:0] w_n971_0;
	wire[1:0] w_n973_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n975_0;
	wire[1:0] w_n976_0;
	wire[1:0] w_n978_0;
	wire[1:0] w_n979_0;
	wire[1:0] w_n980_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n983_0;
	wire[1:0] w_n984_0;
	wire[1:0] w_n985_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n988_0;
	wire[1:0] w_n989_0;
	wire[1:0] w_n990_0;
	wire[1:0] w_n991_0;
	wire[1:0] w_n993_0;
	wire[1:0] w_n994_0;
	wire[1:0] w_n995_0;
	wire[1:0] w_n996_0;
	wire[1:0] w_n997_0;
	wire[1:0] w_n998_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1002_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1005_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1010_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1012_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1015_0;
	wire[1:0] w_n1016_0;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1019_0;
	wire[1:0] w_n1020_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[1:0] w_n1024_0;
	wire[1:0] w_n1025_0;
	wire[1:0] w_n1027_0;
	wire[1:0] w_n1028_0;
	wire[1:0] w_n1029_0;
	wire[1:0] w_n1030_0;
	wire[1:0] w_n1032_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1034_0;
	wire[1:0] w_n1035_0;
	wire[1:0] w_n1037_0;
	wire[1:0] w_n1038_0;
	wire[1:0] w_n1039_0;
	wire[1:0] w_n1040_0;
	wire[2:0] w_n1041_0;
	wire[1:0] w_n1042_0;
	wire[2:0] w_n1044_0;
	wire[1:0] w_n1046_0;
	wire[1:0] w_n1049_0;
	wire[1:0] w_n1054_0;
	wire[1:0] w_n1055_0;
	wire[1:0] w_n1059_0;
	wire[1:0] w_n1060_0;
	wire[1:0] w_n1063_0;
	wire[1:0] w_n1065_0;
	wire[1:0] w_n1067_0;
	wire[1:0] w_n1070_0;
	wire[1:0] w_n1072_0;
	wire[1:0] w_n1074_0;
	wire[1:0] w_n1076_0;
	wire[1:0] w_n1078_0;
	wire[1:0] w_n1080_0;
	wire[1:0] w_n1083_0;
	wire[1:0] w_n1084_0;
	wire[1:0] w_n1087_0;
	wire[1:0] w_n1089_0;
	wire[1:0] w_n1091_0;
	wire[1:0] w_n1094_0;
	wire[1:0] w_n1096_0;
	wire[1:0] w_n1098_0;
	wire[1:0] w_n1108_0;
	wire[1:0] w_n1110_0;
	wire[1:0] w_n1112_0;
	wire[1:0] w_n1115_0;
	wire[1:0] w_n1116_0;
	wire[1:0] w_n1119_0;
	wire[1:0] w_n1121_0;
	wire[1:0] w_n1123_0;
	wire[1:0] w_n1126_0;
	wire[1:0] w_n1128_0;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1140_0;
	wire[1:0] w_n1142_0;
	wire[1:0] w_n1144_0;
	wire[1:0] w_n1147_0;
	wire[1:0] w_n1148_0;
	wire[1:0] w_n1151_0;
	wire[1:0] w_n1153_0;
	wire[1:0] w_n1155_0;
	wire[1:0] w_n1158_0;
	wire[1:0] w_n1160_0;
	wire[1:0] w_n1162_0;
	wire[1:0] w_n1172_0;
	wire[1:0] w_n1174_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1179_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1185_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1190_0;
	wire[1:0] w_n1195_0;
	wire[1:0] w_n1198_0;
	wire[1:0] w_n1201_0;
	wire[1:0] w_n1206_0;
	wire[1:0] w_n1210_0;
	wire[1:0] w_n1213_0;
	wire[1:0] w_n1216_0;
	wire[1:0] w_n1218_0;
	wire[1:0] w_n1223_0;
	wire[1:0] w_n1225_0;
	wire[1:0] w_n1233_0;
	wire[1:0] w_n1236_0;
	wire[1:0] w_n1239_0;
	wire[1:0] w_n1241_0;
	wire[1:0] w_n1242_0;
	wire[1:0] w_n1244_0;
	wire[1:0] w_n1248_0;
	wire[1:0] w_n1250_0;
	wire[1:0] w_n1253_0;
	wire[1:0] w_n1255_0;
	wire[1:0] w_n1258_0;
	wire[1:0] w_n1263_0;
	wire[1:0] w_n1267_0;
	wire[1:0] w_n1270_0;
	wire[1:0] w_n1272_0;
	wire[1:0] w_n1278_0;
	wire[1:0] w_n1282_0;
	wire[1:0] w_n1285_0;
	wire[1:0] w_n1287_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1290_0;
	wire[1:0] w_n1294_0;
	wire[1:0] w_n1296_0;
	wire[1:0] w_n1299_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1304_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1319_0;
	wire[1:0] w_n1324_0;
	wire[1:0] w_n1328_0;
	wire[1:0] w_n1330_0;
	wire[1:0] w_n1333_0;
	wire[1:0] w_n1335_0;
	wire[1:0] w_n1337_0;
	wire[1:0] w_n1340_0;
	wire[1:0] w_n1342_0;
	wire[1:0] w_n1345_0;
	wire[1:0] w_n1347_0;
	wire[1:0] w_n1349_0;
	wire[1:0] w_n1352_0;
	wire[1:0] w_n1353_0;
	wire[1:0] w_n1355_0;
	wire[1:0] w_n1359_0;
	wire[1:0] w_n1363_0;
	wire[1:0] w_n1367_0;
	wire[1:0] w_n1369_0;
	wire[1:0] w_n1372_0;
	wire[1:0] w_n1374_0;
	wire[1:0] w_n1376_0;
	wire[1:0] w_n1379_0;
	wire[1:0] w_n1380_0;
	wire[1:0] w_n1382_0;
	wire[1:0] w_n1386_0;
	wire[1:0] w_n1390_0;
	wire[1:0] w_n1394_0;
	wire[1:0] w_n1396_0;
	wire[1:0] w_n1399_0;
	wire[1:0] w_n1401_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1404_0;
	wire[1:0] w_n1406_0;
	wire[1:0] w_n1407_0;
	wire[1:0] w_n1409_0;
	wire[1:0] w_n1412_0;
	wire[1:0] w_n1414_0;
	wire[1:0] w_n1418_0;
	wire[1:0] w_n1422_0;
	wire[1:0] w_n1426_0;
	wire[1:0] w_n1428_0;
	wire[1:0] w_n1431_0;
	wire[1:0] w_n1433_0;
	wire[1:0] w_n1435_0;
	wire[1:0] w_n1438_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1449_0;
	wire[1:0] w_n1453_0;
	wire[1:0] w_n1455_0;
	wire[1:0] w_n1458_0;
	wire[1:0] w_n1460_0;
	wire[1:0] w_n1462_0;
	wire[1:0] w_n1465_0;
	wire[1:0] w_n1466_0;
	wire[1:0] w_n1468_0;
	wire[1:0] w_n1472_0;
	wire[1:0] w_n1476_0;
	wire[1:0] w_n1480_0;
	wire[1:0] w_n1482_0;
	wire[1:0] w_n1485_0;
	wire[1:0] w_n1487_0;
	wire[1:0] w_n1489_0;
	wire[1:0] w_n1492_0;
	wire[1:0] w_n1493_0;
	wire[1:0] w_n1495_0;
	wire[1:0] w_n1499_0;
	wire[1:0] w_n1503_0;
	wire[1:0] w_n1507_0;
	wire[1:0] w_n1509_0;
	wire[1:0] w_n1512_0;
	wire[1:0] w_n1514_0;
	wire[1:0] w_n1516_0;
	wire[1:0] w_n1519_0;
	wire[1:0] w_n1520_0;
	wire[1:0] w_n1522_0;
	wire[1:0] w_n1526_0;
	wire[1:0] w_n1530_0;
	wire[1:0] w_n1534_0;
	wire[1:0] w_n1536_0;
	wire[1:0] w_n1538_0;
	wire[1:0] w_n1539_0;
	wire[1:0] w_n1542_0;
	wire[1:0] w_n1544_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1554_0;
	wire[1:0] w_n1560_0;
	wire[2:0] w_n1562_0;
	wire[2:0] w_n1562_1;
	wire[2:0] w_n1562_2;
	wire[2:0] w_n1562_3;
	wire[2:0] w_n1562_4;
	wire[2:0] w_n1562_5;
	wire[2:0] w_n1562_6;
	wire[2:0] w_n1562_7;
	wire[2:0] w_n1562_8;
	wire[2:0] w_n1562_9;
	wire[2:0] w_n1562_10;
	wire[2:0] w_n1562_11;
	wire[2:0] w_n1562_12;
	wire[2:0] w_n1562_13;
	wire[2:0] w_n1562_14;
	wire[2:0] w_n1562_15;
	wire[2:0] w_n1562_16;
	wire[2:0] w_n1562_17;
	wire[2:0] w_n1562_18;
	wire[2:0] w_n1562_19;
	wire[2:0] w_n1562_20;
	wire[2:0] w_n1562_21;
	wire[2:0] w_n1562_22;
	wire[2:0] w_n1562_23;
	wire[2:0] w_n1562_24;
	wire[2:0] w_n1562_25;
	wire[2:0] w_n1562_26;
	wire[2:0] w_n1562_27;
	wire[2:0] w_n1562_28;
	wire[2:0] w_n1562_29;
	wire[2:0] w_n1562_30;
	wire[2:0] w_n1562_31;
	wire[2:0] w_n1562_32;
	wire[2:0] w_n1562_33;
	wire[2:0] w_n1562_34;
	wire[2:0] w_n1562_35;
	wire[2:0] w_n1562_36;
	wire[2:0] w_n1562_37;
	wire[2:0] w_n1562_38;
	wire[2:0] w_n1562_39;
	wire[2:0] w_n1562_40;
	wire[2:0] w_n1562_41;
	wire[2:0] w_n1562_42;
	wire[2:0] w_n1562_43;
	wire[2:0] w_n1562_44;
	wire[2:0] w_n1562_45;
	wire[2:0] w_n1562_46;
	wire[2:0] w_n1562_47;
	wire[2:0] w_n1562_48;
	wire[2:0] w_n1562_49;
	wire[2:0] w_n1562_50;
	wire[2:0] w_n1562_51;
	wire[2:0] w_n1562_52;
	wire[2:0] w_n1562_53;
	wire[2:0] w_n1562_54;
	wire[2:0] w_n1562_55;
	wire[2:0] w_n1562_56;
	wire[2:0] w_n1562_57;
	wire[2:0] w_n1562_58;
	wire[2:0] w_n1562_59;
	wire[2:0] w_n1562_60;
	wire[2:0] w_n1562_61;
	wire[2:0] w_n1562_62;
	wire[2:0] w_n1562_63;
	wire[2:0] w_n1562_64;
	wire[2:0] w_n1586_0;
	wire[1:0] w_n1588_0;
	wire[2:0] w_n1721_0;
	wire[2:0] w_n1721_1;
	wire[2:0] w_n1721_2;
	wire[2:0] w_n1721_3;
	wire[2:0] w_n1721_4;
	wire[2:0] w_n1721_5;
	wire[2:0] w_n1721_6;
	wire[2:0] w_n1721_7;
	wire[2:0] w_n1721_8;
	wire[2:0] w_n1721_9;
	wire[2:0] w_n1721_10;
	wire[2:0] w_n1721_11;
	wire[2:0] w_n1721_12;
	wire[2:0] w_n1721_13;
	wire[2:0] w_n1721_14;
	wire[2:0] w_n1721_15;
	wire[2:0] w_n1721_16;
	wire[2:0] w_n1721_17;
	wire[2:0] w_n1721_18;
	wire[2:0] w_n1721_19;
	wire[2:0] w_n1721_20;
	wire[2:0] w_n1721_21;
	wire[2:0] w_n1721_22;
	wire[2:0] w_n1721_23;
	wire[2:0] w_n1721_24;
	wire[2:0] w_n1721_25;
	wire[2:0] w_n1721_26;
	wire[2:0] w_n1721_27;
	wire[2:0] w_n1721_28;
	wire[2:0] w_n1721_29;
	wire[2:0] w_n1721_30;
	wire[2:0] w_n1721_31;
	wire[2:0] w_n1721_32;
	wire[2:0] w_n1721_33;
	wire[2:0] w_n1721_34;
	wire[2:0] w_n1721_35;
	wire[2:0] w_n1721_36;
	wire[2:0] w_n1721_37;
	wire[2:0] w_n1721_38;
	wire[2:0] w_n1721_39;
	wire[2:0] w_n1721_40;
	wire[2:0] w_n1721_41;
	wire[2:0] w_n1721_42;
	wire[2:0] w_n1721_43;
	wire[2:0] w_n1721_44;
	wire[2:0] w_n1721_45;
	wire[2:0] w_n1721_46;
	wire[2:0] w_n1721_47;
	wire[2:0] w_n1721_48;
	wire[2:0] w_n1721_49;
	wire[2:0] w_n1721_50;
	wire[2:0] w_n1721_51;
	wire[2:0] w_n1721_52;
	wire[2:0] w_n1721_53;
	wire[2:0] w_n1721_54;
	wire[2:0] w_n1721_55;
	wire[2:0] w_n1721_56;
	wire[2:0] w_n1721_57;
	wire[2:0] w_n1721_58;
	wire[2:0] w_n1721_59;
	wire[2:0] w_n1721_60;
	wire[2:0] w_n1721_61;
	wire[2:0] w_n1721_62;
	wire[2:0] w_n1721_63;
	wire[2:0] w_n1721_64;
	wire[1:0] w_n1721_65;
	wire[1:0] w_n1723_0;
	wire[1:0] w_n1724_0;
	wire[1:0] w_n1726_0;
	wire[1:0] w_n1728_0;
	wire[1:0] w_n1730_0;
	wire[1:0] w_n1732_0;
	wire[1:0] w_n1736_0;
	wire[1:0] w_n1738_0;
	wire[1:0] w_n1740_0;
	wire[1:0] w_n1741_0;
	wire[1:0] w_n1743_0;
	wire[1:0] w_n1745_0;
	wire[1:0] w_n1746_0;
	wire[1:0] w_n1747_0;
	wire[1:0] w_n1750_0;
	wire[1:0] w_n1752_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1759_0;
	wire[1:0] w_n1761_0;
	wire[1:0] w_n1765_0;
	wire[1:0] w_n1767_0;
	wire[1:0] w_n1768_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1771_0;
	wire[1:0] w_n1772_0;
	wire[1:0] w_n1774_0;
	wire[1:0] w_n1775_0;
	wire[1:0] w_n1777_0;
	wire[1:0] w_n1778_0;
	wire[1:0] w_n1779_0;
	wire[1:0] w_n1782_0;
	wire[1:0] w_n1784_0;
	wire[1:0] w_n1786_0;
	wire[1:0] w_n1791_0;
	wire[1:0] w_n1793_0;
	wire[1:0] w_n1797_0;
	wire[1:0] w_n1799_0;
	wire[1:0] w_n1800_0;
	wire[1:0] w_n1802_0;
	wire[1:0] w_n1804_0;
	wire[1:0] w_n1805_0;
	wire[1:0] w_n1806_0;
	wire[1:0] w_n1809_0;
	wire[1:0] w_n1811_0;
	wire[1:0] w_n1813_0;
	wire[1:0] w_n1818_0;
	wire[1:0] w_n1820_0;
	wire[1:0] w_n1824_0;
	wire[1:0] w_n1826_0;
	wire[1:0] w_n1827_0;
	wire[1:0] w_n1829_0;
	wire[1:0] w_n1830_0;
	wire[1:0] w_n1831_0;
	wire[1:0] w_n1833_0;
	wire[1:0] w_n1834_0;
	wire[1:0] w_n1836_0;
	wire[1:0] w_n1837_0;
	wire[1:0] w_n1838_0;
	wire[1:0] w_n1841_0;
	wire[1:0] w_n1843_0;
	wire[1:0] w_n1845_0;
	wire[1:0] w_n1850_0;
	wire[1:0] w_n1852_0;
	wire[1:0] w_n1856_0;
	wire[1:0] w_n1858_0;
	wire[1:0] w_n1859_0;
	wire[1:0] w_n1861_0;
	wire[1:0] w_n1863_0;
	wire[1:0] w_n1864_0;
	wire[1:0] w_n1865_0;
	wire[1:0] w_n1868_0;
	wire[1:0] w_n1870_0;
	wire[1:0] w_n1872_0;
	wire[1:0] w_n1877_0;
	wire[1:0] w_n1879_0;
	wire[1:0] w_n1883_0;
	wire[1:0] w_n1885_0;
	wire[1:0] w_n1886_0;
	wire[1:0] w_n1888_0;
	wire[1:0] w_n1889_0;
	wire[1:0] w_n1890_0;
	wire[1:0] w_n1892_0;
	wire[1:0] w_n1893_0;
	wire[1:0] w_n1895_0;
	wire[1:0] w_n1896_0;
	wire[1:0] w_n1897_0;
	wire[1:0] w_n1900_0;
	wire[1:0] w_n1902_0;
	wire[1:0] w_n1904_0;
	wire[1:0] w_n1909_0;
	wire[1:0] w_n1911_0;
	wire[1:0] w_n1915_0;
	wire[1:0] w_n1917_0;
	wire[1:0] w_n1918_0;
	wire[1:0] w_n1920_0;
	wire[1:0] w_n1922_0;
	wire[1:0] w_n1923_0;
	wire[1:0] w_n1924_0;
	wire[1:0] w_n1927_0;
	wire[1:0] w_n1929_0;
	wire[1:0] w_n1931_0;
	wire[1:0] w_n1936_0;
	wire[1:0] w_n1938_0;
	wire[1:0] w_n1942_0;
	wire[1:0] w_n1944_0;
	wire[1:0] w_n1945_0;
	wire[1:0] w_n1947_0;
	wire[1:0] w_n1948_0;
	wire[1:0] w_n1950_0;
	wire[1:0] w_n1953_0;
	wire[1:0] w_n1955_0;
	wire[1:0] w_n1958_0;
	wire[1:0] w_n1960_0;
	wire[1:0] w_n1961_0;
	wire[1:0] w_n1963_0;
	wire[1:0] w_n1964_0;
	wire[1:0] w_n1965_0;
	wire[1:0] w_n1967_0;
	wire[1:0] w_n1970_0;
	wire[1:0] w_n1971_0;
	wire[1:0] w_n1974_0;
	wire[1:0] w_n1976_0;
	wire[1:0] w_n1977_0;
	wire[1:0] w_n1978_0;
	wire[1:0] w_n1979_0;
	wire[1:0] w_n1981_0;
	wire[1:0] w_n1983_0;
	wire[1:0] w_n1984_0;
	wire[1:0] w_n1987_0;
	wire[1:0] w_n1990_0;
	wire[1:0] w_n1992_0;
	wire[1:0] w_n1993_0;
	wire[1:0] w_n1995_0;
	wire[1:0] w_n1996_0;
	wire[1:0] w_n1997_0;
	wire[1:0] w_n1999_0;
	wire[1:0] w_n2002_0;
	wire[1:0] w_n2003_0;
	wire[1:0] w_n2006_0;
	wire[1:0] w_n2008_0;
	wire[1:0] w_n2010_0;
	wire[1:0] w_n2013_0;
	wire[1:0] w_n2014_0;
	wire[1:0] w_n2016_0;
	wire[1:0] w_n2020_0;
	wire[1:0] w_n2022_0;
	wire[1:0] w_n2025_0;
	wire[1:0] w_n2027_0;
	wire[1:0] w_n2029_0;
	wire[1:0] w_n2030_0;
	wire[1:0] w_n2031_0;
	wire[1:0] w_n2034_0;
	wire[1:0] w_n2035_0;
	wire[1:0] w_n2036_0;
	wire[1:0] w_n2038_0;
	wire[1:0] w_n2040_0;
	wire[1:0] w_n2041_0;
	wire[1:0] w_n2042_0;
	wire[1:0] w_n2043_0;
	wire[1:0] w_n2045_0;
	wire[1:0] w_n2046_0;
	wire[1:0] w_n2047_0;
	wire[1:0] w_n2048_0;
	wire[1:0] w_n2050_0;
	wire[1:0] w_n2051_0;
	wire[1:0] w_n2052_0;
	wire[1:0] w_n2053_0;
	wire[1:0] w_n2055_0;
	wire[1:0] w_n2056_0;
	wire[1:0] w_n2057_0;
	wire[1:0] w_n2058_0;
	wire[1:0] w_n2060_0;
	wire[1:0] w_n2061_0;
	wire[1:0] w_n2062_0;
	wire[1:0] w_n2063_0;
	wire[1:0] w_n2064_0;
	wire[1:0] w_n2065_0;
	wire[1:0] w_n2067_0;
	wire[1:0] w_n2068_0;
	wire[1:0] w_n2069_0;
	wire[1:0] w_n2070_0;
	wire[1:0] w_n2072_0;
	wire[1:0] w_n2073_0;
	wire[1:0] w_n2074_0;
	wire[1:0] w_n2075_0;
	wire[1:0] w_n2077_0;
	wire[1:0] w_n2078_0;
	wire[1:0] w_n2079_0;
	wire[1:0] w_n2080_0;
	wire[1:0] w_n2082_0;
	wire[1:0] w_n2083_0;
	wire[1:0] w_n2084_0;
	wire[1:0] w_n2085_0;
	wire[1:0] w_n2086_0;
	wire[1:0] w_n2087_0;
	wire[1:0] w_n2089_0;
	wire[1:0] w_n2090_0;
	wire[1:0] w_n2091_0;
	wire[1:0] w_n2092_0;
	wire[1:0] w_n2094_0;
	wire[1:0] w_n2095_0;
	wire[1:0] w_n2096_0;
	wire[1:0] w_n2097_0;
	wire[1:0] w_n2099_0;
	wire[1:0] w_n2100_0;
	wire[1:0] w_n2101_0;
	wire[1:0] w_n2102_0;
	wire[1:0] w_n2104_0;
	wire[1:0] w_n2105_0;
	wire[1:0] w_n2106_0;
	wire[1:0] w_n2107_0;
	wire[1:0] w_n2108_0;
	wire[1:0] w_n2109_0;
	wire[2:0] w_n2110_0;
	wire[1:0] w_n2111_0;
	wire[1:0] w_n2113_0;
	wire[1:0] w_n2115_0;
	wire[1:0] w_n2120_0;
	wire[1:0] w_n2122_0;
	wire[1:0] w_n2124_0;
	wire[1:0] w_n2127_0;
	wire[1:0] w_n2128_0;
	wire[1:0] w_n2131_0;
	wire[1:0] w_n2133_0;
	wire[1:0] w_n2135_0;
	wire[1:0] w_n2138_0;
	wire[1:0] w_n2140_0;
	wire[1:0] w_n2142_0;
	wire[1:0] w_n2144_0;
	wire[1:0] w_n2146_0;
	wire[1:0] w_n2148_0;
	wire[1:0] w_n2151_0;
	wire[1:0] w_n2152_0;
	wire[1:0] w_n2155_0;
	wire[1:0] w_n2157_0;
	wire[1:0] w_n2159_0;
	wire[1:0] w_n2162_0;
	wire[1:0] w_n2164_0;
	wire[1:0] w_n2166_0;
	wire[1:0] w_n2176_0;
	wire[1:0] w_n2178_0;
	wire[1:0] w_n2180_0;
	wire[1:0] w_n2183_0;
	wire[1:0] w_n2184_0;
	wire[1:0] w_n2187_0;
	wire[1:0] w_n2189_0;
	wire[1:0] w_n2191_0;
	wire[1:0] w_n2194_0;
	wire[1:0] w_n2196_0;
	wire[1:0] w_n2198_0;
	wire[1:0] w_n2208_0;
	wire[1:0] w_n2210_0;
	wire[1:0] w_n2212_0;
	wire[1:0] w_n2215_0;
	wire[1:0] w_n2216_0;
	wire[1:0] w_n2219_0;
	wire[1:0] w_n2221_0;
	wire[1:0] w_n2223_0;
	wire[1:0] w_n2226_0;
	wire[1:0] w_n2228_0;
	wire[1:0] w_n2230_0;
	wire[1:0] w_n2240_0;
	wire[1:0] w_n2242_0;
	wire[1:0] w_n2244_0;
	wire[1:0] w_n2247_0;
	wire[1:0] w_n2249_0;
	wire[1:0] w_n2253_0;
	wire[1:0] w_n2256_0;
	wire[1:0] w_n2258_0;
	wire[1:0] w_n2263_0;
	wire[1:0] w_n2266_0;
	wire[1:0] w_n2269_0;
	wire[1:0] w_n2274_0;
	wire[1:0] w_n2278_0;
	wire[1:0] w_n2281_0;
	wire[1:0] w_n2283_0;
	wire[1:0] w_n2284_0;
	wire[1:0] w_n2286_0;
	wire[1:0] w_n2290_0;
	wire[1:0] w_n2292_0;
	wire[1:0] w_n2295_0;
	wire[1:0] w_n2297_0;
	wire[1:0] w_n2300_0;
	wire[1:0] w_n2306_0;
	wire[1:0] w_n2308_0;
	wire[1:0] w_n2313_0;
	wire[1:0] w_n2315_0;
	wire[1:0] w_n2320_0;
	wire[1:0] w_n2324_0;
	wire[1:0] w_n2327_0;
	wire[1:0] w_n2329_0;
	wire[1:0] w_n2330_0;
	wire[1:0] w_n2332_0;
	wire[1:0] w_n2336_0;
	wire[1:0] w_n2338_0;
	wire[1:0] w_n2341_0;
	wire[1:0] w_n2343_0;
	wire[1:0] w_n2346_0;
	wire[1:0] w_n2351_0;
	wire[1:0] w_n2355_0;
	wire[1:0] w_n2358_0;
	wire[1:0] w_n2360_0;
	wire[1:0] w_n2366_0;
	wire[1:0] w_n2370_0;
	wire[1:0] w_n2373_0;
	wire[1:0] w_n2375_0;
	wire[1:0] w_n2376_0;
	wire[1:0] w_n2378_0;
	wire[1:0] w_n2382_0;
	wire[1:0] w_n2384_0;
	wire[1:0] w_n2387_0;
	wire[1:0] w_n2389_0;
	wire[1:0] w_n2392_0;
	wire[1:0] w_n2398_0;
	wire[1:0] w_n2400_0;
	wire[1:0] w_n2405_0;
	wire[1:0] w_n2407_0;
	wire[1:0] w_n2412_0;
	wire[1:0] w_n2416_0;
	wire[1:0] w_n2418_0;
	wire[1:0] w_n2421_0;
	wire[1:0] w_n2423_0;
	wire[1:0] w_n2425_0;
	wire[1:0] w_n2428_0;
	wire[1:0] w_n2430_0;
	wire[1:0] w_n2433_0;
	wire[1:0] w_n2435_0;
	wire[1:0] w_n2437_0;
	wire[1:0] w_n2438_0;
	wire[1:0] w_n2440_0;
	wire[1:0] w_n2441_0;
	wire[1:0] w_n2443_0;
	wire[1:0] w_n2446_0;
	wire[1:0] w_n2448_0;
	wire[1:0] w_n2452_0;
	wire[1:0] w_n2456_0;
	wire[1:0] w_n2460_0;
	wire[1:0] w_n2462_0;
	wire[1:0] w_n2465_0;
	wire[1:0] w_n2467_0;
	wire[1:0] w_n2469_0;
	wire[1:0] w_n2472_0;
	wire[1:0] w_n2473_0;
	wire[1:0] w_n2475_0;
	wire[1:0] w_n2479_0;
	wire[1:0] w_n2483_0;
	wire[1:0] w_n2487_0;
	wire[1:0] w_n2489_0;
	wire[1:0] w_n2492_0;
	wire[1:0] w_n2494_0;
	wire[1:0] w_n2496_0;
	wire[1:0] w_n2497_0;
	wire[1:0] w_n2499_0;
	wire[1:0] w_n2500_0;
	wire[1:0] w_n2502_0;
	wire[1:0] w_n2505_0;
	wire[1:0] w_n2507_0;
	wire[1:0] w_n2511_0;
	wire[1:0] w_n2515_0;
	wire[1:0] w_n2519_0;
	wire[1:0] w_n2521_0;
	wire[1:0] w_n2524_0;
	wire[1:0] w_n2526_0;
	wire[1:0] w_n2528_0;
	wire[1:0] w_n2531_0;
	wire[1:0] w_n2532_0;
	wire[1:0] w_n2534_0;
	wire[1:0] w_n2538_0;
	wire[1:0] w_n2542_0;
	wire[1:0] w_n2546_0;
	wire[1:0] w_n2548_0;
	wire[1:0] w_n2551_0;
	wire[1:0] w_n2553_0;
	wire[1:0] w_n2555_0;
	wire[1:0] w_n2556_0;
	wire[1:0] w_n2558_0;
	wire[1:0] w_n2559_0;
	wire[1:0] w_n2561_0;
	wire[1:0] w_n2564_0;
	wire[1:0] w_n2566_0;
	wire[1:0] w_n2570_0;
	wire[1:0] w_n2574_0;
	wire[1:0] w_n2578_0;
	wire[1:0] w_n2580_0;
	wire[1:0] w_n2583_0;
	wire[1:0] w_n2585_0;
	wire[1:0] w_n2587_0;
	wire[1:0] w_n2590_0;
	wire[1:0] w_n2591_0;
	wire[1:0] w_n2593_0;
	wire[1:0] w_n2597_0;
	wire[1:0] w_n2601_0;
	wire[1:0] w_n2605_0;
	wire[1:0] w_n2607_0;
	wire[1:0] w_n2610_0;
	wire[1:0] w_n2612_0;
	wire[1:0] w_n2614_0;
	wire[1:0] w_n2615_0;
	wire[1:0] w_n2617_0;
	wire[1:0] w_n2618_0;
	wire[1:0] w_n2620_0;
	wire[1:0] w_n2623_0;
	wire[1:0] w_n2625_0;
	wire[1:0] w_n2629_0;
	wire[1:0] w_n2633_0;
	wire[1:0] w_n2637_0;
	wire[1:0] w_n2639_0;
	wire[2:0] w_n2641_0;
	wire[1:0] w_n2642_0;
	wire[2:0] w_n2643_0;
	wire[1:0] w_n2643_1;
	wire[1:0] w_n2644_0;
	wire[1:0] w_n2647_0;
	wire[1:0] w_n2648_0;
	wire[1:0] w_n2649_0;
	wire[1:0] w_n2672_0;
	wire[1:0] w_n2801_0;
	wire[2:0] w_n2803_0;
	wire[2:0] w_n2803_1;
	wire[2:0] w_n2803_2;
	wire[2:0] w_n2803_3;
	wire[2:0] w_n2803_4;
	wire[2:0] w_n2803_5;
	wire[2:0] w_n2803_6;
	wire[2:0] w_n2803_7;
	wire[2:0] w_n2803_8;
	wire[2:0] w_n2803_9;
	wire[2:0] w_n2803_10;
	wire[2:0] w_n2803_11;
	wire[2:0] w_n2803_12;
	wire[2:0] w_n2803_13;
	wire[2:0] w_n2803_14;
	wire[2:0] w_n2803_15;
	wire[2:0] w_n2803_16;
	wire[2:0] w_n2803_17;
	wire[2:0] w_n2803_18;
	wire[2:0] w_n2803_19;
	wire[2:0] w_n2803_20;
	wire[2:0] w_n2803_21;
	wire[2:0] w_n2803_22;
	wire[2:0] w_n2803_23;
	wire[2:0] w_n2803_24;
	wire[2:0] w_n2803_25;
	wire[2:0] w_n2803_26;
	wire[2:0] w_n2803_27;
	wire[2:0] w_n2803_28;
	wire[2:0] w_n2803_29;
	wire[2:0] w_n2803_30;
	wire[2:0] w_n2803_31;
	wire[2:0] w_n2803_32;
	wire[2:0] w_n2803_33;
	wire[2:0] w_n2803_34;
	wire[2:0] w_n2803_35;
	wire[2:0] w_n2803_36;
	wire[2:0] w_n2803_37;
	wire[2:0] w_n2803_38;
	wire[2:0] w_n2803_39;
	wire[2:0] w_n2803_40;
	wire[2:0] w_n2803_41;
	wire[2:0] w_n2803_42;
	wire[2:0] w_n2803_43;
	wire[2:0] w_n2803_44;
	wire[2:0] w_n2803_45;
	wire[2:0] w_n2803_46;
	wire[2:0] w_n2803_47;
	wire[2:0] w_n2803_48;
	wire[2:0] w_n2803_49;
	wire[2:0] w_n2803_50;
	wire[2:0] w_n2803_51;
	wire[2:0] w_n2803_52;
	wire[2:0] w_n2803_53;
	wire[2:0] w_n2803_54;
	wire[2:0] w_n2803_55;
	wire[2:0] w_n2803_56;
	wire[2:0] w_n2803_57;
	wire[2:0] w_n2803_58;
	wire[2:0] w_n2803_59;
	wire[2:0] w_n2803_60;
	wire[2:0] w_n2803_61;
	wire[2:0] w_n2803_62;
	wire[2:0] w_n2803_63;
	wire[1:0] w_n2803_64;
	wire[2:0] w_n2808_0;
	wire[2:0] w_n2808_1;
	wire[2:0] w_n2808_2;
	wire[2:0] w_n2808_3;
	wire[2:0] w_n2808_4;
	wire[2:0] w_n2808_5;
	wire[2:0] w_n2808_6;
	wire[2:0] w_n2808_7;
	wire[2:0] w_n2808_8;
	wire[2:0] w_n2808_9;
	wire[2:0] w_n2808_10;
	wire[2:0] w_n2808_11;
	wire[2:0] w_n2808_12;
	wire[2:0] w_n2808_13;
	wire[2:0] w_n2808_14;
	wire[2:0] w_n2808_15;
	wire[2:0] w_n2808_16;
	wire[2:0] w_n2808_17;
	wire[2:0] w_n2808_18;
	wire[2:0] w_n2808_19;
	wire[2:0] w_n2808_20;
	wire[2:0] w_n2808_21;
	wire[2:0] w_n2808_22;
	wire[2:0] w_n2808_23;
	wire[2:0] w_n2808_24;
	wire[2:0] w_n2808_25;
	wire[2:0] w_n2808_26;
	wire[2:0] w_n2808_27;
	wire[2:0] w_n2808_28;
	wire[2:0] w_n2808_29;
	wire[2:0] w_n2808_30;
	wire[2:0] w_n2808_31;
	wire[2:0] w_n2808_32;
	wire[2:0] w_n2808_33;
	wire[2:0] w_n2808_34;
	wire[2:0] w_n2808_35;
	wire[2:0] w_n2808_36;
	wire[2:0] w_n2808_37;
	wire[2:0] w_n2808_38;
	wire[2:0] w_n2808_39;
	wire[2:0] w_n2808_40;
	wire[2:0] w_n2808_41;
	wire[2:0] w_n2808_42;
	wire[2:0] w_n2808_43;
	wire[2:0] w_n2808_44;
	wire[2:0] w_n2808_45;
	wire[2:0] w_n2808_46;
	wire[2:0] w_n2808_47;
	wire[2:0] w_n2808_48;
	wire[2:0] w_n2808_49;
	wire[2:0] w_n2808_50;
	wire[2:0] w_n2808_51;
	wire[2:0] w_n2808_52;
	wire[2:0] w_n2808_53;
	wire[2:0] w_n2808_54;
	wire[2:0] w_n2808_55;
	wire[2:0] w_n2808_56;
	wire[2:0] w_n2808_57;
	wire[2:0] w_n2808_58;
	wire[2:0] w_n2808_59;
	wire[2:0] w_n2808_60;
	wire[2:0] w_n2808_61;
	wire[2:0] w_n2808_62;
	wire[2:0] w_n2808_63;
	wire[2:0] w_n2808_64;
	wire[1:0] w_n2810_0;
	wire[1:0] w_n2811_0;
	wire[1:0] w_n2815_0;
	wire[1:0] w_n2818_0;
	wire[1:0] w_n2819_0;
	wire[1:0] w_n2821_0;
	wire[1:0] w_n2825_0;
	wire[1:0] w_n2826_0;
	wire[1:0] w_n2829_0;
	wire[1:0] w_n2831_0;
	wire[1:0] w_n2835_0;
	wire[1:0] w_n2837_0;
	wire[1:0] w_n2839_0;
	wire[1:0] w_n2841_0;
	wire[1:0] w_n2844_0;
	wire[1:0] w_n2845_0;
	wire[1:0] w_n2848_0;
	wire[1:0] w_n2852_0;
	wire[1:0] w_n2855_0;
	wire[1:0] w_n2856_0;
	wire[1:0] w_n2857_0;
	wire[1:0] w_n2860_0;
	wire[1:0] w_n2863_0;
	wire[1:0] w_n2864_0;
	wire[1:0] w_n2867_0;
	wire[1:0] w_n2869_0;
	wire[1:0] w_n2873_0;
	wire[1:0] w_n2874_0;
	wire[1:0] w_n2877_0;
	wire[1:0] w_n2882_0;
	wire[1:0] w_n2884_0;
	wire[1:0] w_n2888_0;
	wire[1:0] w_n2892_0;
	wire[1:0] w_n2893_0;
	wire[1:0] w_n2896_0;
	wire[1:0] w_n2897_0;
	wire[1:0] w_n2901_0;
	wire[1:0] w_n2902_0;
	wire[1:0] w_n2905_0;
	wire[1:0] w_n2909_0;
	wire[1:0] w_n2912_0;
	wire[1:0] w_n2913_0;
	wire[1:0] w_n2914_0;
	wire[1:0] w_n2917_0;
	wire[1:0] w_n2920_0;
	wire[1:0] w_n2921_0;
	wire[1:0] w_n2924_0;
	wire[1:0] w_n2926_0;
	wire[1:0] w_n2930_0;
	wire[1:0] w_n2931_0;
	wire[1:0] w_n2934_0;
	wire[1:0] w_n2937_0;
	wire[1:0] w_n2939_0;
	wire[1:0] w_n2941_0;
	wire[1:0] w_n2944_0;
	wire[1:0] w_n2947_0;
	wire[1:0] w_n2948_0;
	wire[1:0] w_n2952_0;
	wire[1:0] w_n2953_0;
	wire[1:0] w_n2956_0;
	wire[1:0] w_n2958_0;
	wire[1:0] w_n2961_0;
	wire[1:0] w_n2964_0;
	wire[1:0] w_n2965_0;
	wire[1:0] w_n2966_0;
	wire[1:0] w_n2969_0;
	wire[1:0] w_n2970_0;
	wire[1:0] w_n2973_0;
	wire[1:0] w_n2976_0;
	wire[1:0] w_n2979_0;
	wire[1:0] w_n2982_0;
	wire[1:0] w_n2983_0;
	wire[1:0] w_n2987_0;
	wire[1:0] w_n2988_0;
	wire[1:0] w_n2991_0;
	wire[1:0] w_n2995_0;
	wire[1:0] w_n2998_0;
	wire[1:0] w_n2999_0;
	wire[1:0] w_n3000_0;
	wire[1:0] w_n3003_0;
	wire[1:0] w_n3006_0;
	wire[1:0] w_n3007_0;
	wire[1:0] w_n3010_0;
	wire[1:0] w_n3011_0;
	wire[1:0] w_n3014_0;
	wire[1:0] w_n3017_0;
	wire[1:0] w_n3018_0;
	wire[1:0] w_n3022_0;
	wire[1:0] w_n3023_0;
	wire[1:0] w_n3026_0;
	wire[1:0] w_n3028_0;
	wire[1:0] w_n3031_0;
	wire[1:0] w_n3034_0;
	wire[1:0] w_n3035_0;
	wire[1:0] w_n3036_0;
	wire[1:0] w_n3039_0;
	wire[1:0] w_n3040_0;
	wire[1:0] w_n3043_0;
	wire[1:0] w_n3046_0;
	wire[1:0] w_n3049_0;
	wire[1:0] w_n3052_0;
	wire[1:0] w_n3053_0;
	wire[1:0] w_n3057_0;
	wire[1:0] w_n3058_0;
	wire[1:0] w_n3061_0;
	wire[1:0] w_n3065_0;
	wire[1:0] w_n3068_0;
	wire[1:0] w_n3069_0;
	wire[1:0] w_n3070_0;
	wire[1:0] w_n3073_0;
	wire[1:0] w_n3076_0;
	wire[1:0] w_n3077_0;
	wire[1:0] w_n3080_0;
	wire[1:0] w_n3081_0;
	wire[1:0] w_n3084_0;
	wire[1:0] w_n3087_0;
	wire[1:0] w_n3088_0;
	wire[1:0] w_n3092_0;
	wire[1:0] w_n3093_0;
	wire[1:0] w_n3096_0;
	wire[1:0] w_n3098_0;
	wire[1:0] w_n3101_0;
	wire[1:0] w_n3104_0;
	wire[1:0] w_n3105_0;
	wire[1:0] w_n3106_0;
	wire[1:0] w_n3109_0;
	wire[1:0] w_n3110_0;
	wire[1:0] w_n3113_0;
	wire[1:0] w_n3116_0;
	wire[1:0] w_n3119_0;
	wire[1:0] w_n3120_0;
	wire[1:0] w_n3123_0;
	wire[1:0] w_n3127_0;
	wire[1:0] w_n3130_0;
	wire[1:0] w_n3131_0;
	wire[1:0] w_n3132_0;
	wire[1:0] w_n3135_0;
	wire[1:0] w_n3138_0;
	wire[1:0] w_n3139_0;
	wire[1:0] w_n3142_0;
	wire[1:0] w_n3144_0;
	wire[1:0] w_n3148_0;
	wire[1:0] w_n3149_0;
	wire[1:0] w_n3152_0;
	wire[1:0] w_n3155_0;
	wire[1:0] w_n3158_0;
	wire[1:0] w_n3160_0;
	wire[1:0] w_n3163_0;
	wire[1:0] w_n3167_0;
	wire[1:0] w_n3168_0;
	wire[1:0] w_n3171_0;
	wire[1:0] w_n3172_0;
	wire[1:0] w_n3174_0;
	wire[1:0] w_n3178_0;
	wire[1:0] w_n3179_0;
	wire[1:0] w_n3182_0;
	wire[1:0] w_n3184_0;
	wire[1:0] w_n3187_0;
	wire[1:0] w_n3190_0;
	wire[1:0] w_n3191_0;
	wire[1:0] w_n3192_0;
	wire[1:0] w_n3195_0;
	wire[1:0] w_n3196_0;
	wire[1:0] w_n3199_0;
	wire[1:0] w_n3202_0;
	wire[1:0] w_n3205_0;
	wire[1:0] w_n3208_0;
	wire[1:0] w_n3209_0;
	wire[1:0] w_n3213_0;
	wire[1:0] w_n3214_0;
	wire[1:0] w_n3217_0;
	wire[1:0] w_n3221_0;
	wire[1:0] w_n3224_0;
	wire[1:0] w_n3225_0;
	wire[1:0] w_n3226_0;
	wire[1:0] w_n3229_0;
	wire[1:0] w_n3232_0;
	wire[1:0] w_n3233_0;
	wire[1:0] w_n3236_0;
	wire[1:0] w_n3237_0;
	wire[1:0] w_n3240_0;
	wire[1:0] w_n3241_0;
	wire[1:0] w_n3244_0;
	wire[1:0] w_n3248_0;
	wire[1:0] w_n3251_0;
	wire[1:0] w_n3252_0;
	wire[1:0] w_n3253_0;
	wire[1:0] w_n3256_0;
	wire[1:0] w_n3259_0;
	wire[1:0] w_n3260_0;
	wire[1:0] w_n3263_0;
	wire[1:0] w_n3265_0;
	wire[1:0] w_n3269_0;
	wire[1:0] w_n3270_0;
	wire[1:0] w_n3273_0;
	wire[1:0] w_n3278_0;
	wire[1:0] w_n3280_0;
	wire[1:0] w_n3284_0;
	wire[1:0] w_n3288_0;
	wire[1:0] w_n3289_0;
	wire[1:0] w_n3292_0;
	wire[1:0] w_n3293_0;
	wire[1:0] w_n3297_0;
	wire[1:0] w_n3300_0;
	wire[1:0] w_n3301_0;
	wire[1:0] w_n3305_0;
	wire[1:0] w_n3306_0;
	wire[1:0] w_n3309_0;
	wire[1:0] w_n3311_0;
	wire[1:0] w_n3312_0;
	wire[1:0] w_n3316_0;
	wire[1:0] w_n3319_0;
	wire[1:0] w_n3320_0;
	wire[1:0] w_n3324_0;
	wire[1:0] w_n3328_0;
	wire[1:0] w_n3331_0;
	wire[1:0] w_n3332_0;
	wire[1:0] w_n3336_0;
	wire[1:0] w_n3337_0;
	wire[1:0] w_n3340_0;
	wire[1:0] w_n3344_0;
	wire[1:0] w_n3347_0;
	wire[1:0] w_n3348_0;
	wire[1:0] w_n3349_0;
	wire[1:0] w_n3352_0;
	wire[1:0] w_n3355_0;
	wire[1:0] w_n3356_0;
	wire[1:0] w_n3359_0;
	wire[1:0] w_n3360_0;
	wire[1:0] w_n3364_0;
	wire[1:0] w_n3365_0;
	wire[1:0] w_n3368_0;
	wire[1:0] w_n3370_0;
	wire[1:0] w_n3374_0;
	wire[1:0] w_n3377_0;
	wire[1:0] w_n3378_0;
	wire[1:0] w_n3380_0;
	wire[1:0] w_n3382_0;
	wire[1:0] w_n3386_0;
	wire[1:0] w_n3389_0;
	wire[1:0] w_n3390_0;
	wire[1:0] w_n3391_0;
	wire[1:0] w_n3395_0;
	wire[1:0] w_n3396_0;
	wire[1:0] w_n3399_0;
	wire[1:0] w_n3402_0;
	wire[1:0] w_n3408_0;
	wire[1:0] w_n3412_0;
	wire[1:0] w_n3413_0;
	wire[1:0] w_n3416_0;
	wire[1:0] w_n3417_0;
	wire[2:0] w_n3421_0;
	wire[1:0] w_n3424_0;
	wire[1:0] w_n3427_0;
	wire[1:0] w_n3428_0;
	wire[1:0] w_n3433_0;
	wire[1:0] w_n3436_0;
	wire[1:0] w_n3437_0;
	wire[1:0] w_n3438_0;
	wire[1:0] w_n3441_0;
	wire[1:0] w_n3442_0;
	wire[1:0] w_n3445_0;
	wire[1:0] w_n3448_0;
	wire[1:0] w_n3451_0;
	wire[1:0] w_n3454_0;
	wire[1:0] w_n3455_0;
	wire[1:0] w_n3457_0;
	wire[1:0] w_n3459_0;
	wire[2:0] w_n3463_0;
	wire[1:0] w_n3465_0;
	wire[1:0] w_n3469_0;
	wire[1:0] w_n3472_0;
	wire[1:0] w_n3473_0;
	wire[1:0] w_n3475_0;
	wire[1:0] w_n3478_0;
	wire[1:0] w_n3479_0;
	wire[1:0] w_n3482_0;
	wire[1:0] w_n3486_0;
	wire[1:0] w_n3489_0;
	wire[1:0] w_n3490_0;
	wire[1:0] w_n3493_0;
	wire[1:0] w_n3494_0;
	wire[1:0] w_n3498_0;
	wire[1:0] w_n3499_0;
	wire[1:0] w_n3502_0;
	wire[1:0] w_n3505_0;
	wire[1:0] w_n3507_0;
	wire[1:0] w_n3510_0;
	wire[1:0] w_n3513_0;
	wire[1:0] w_n3514_0;
	wire[1:0] w_n3515_0;
	wire[1:0] w_n3519_0;
	wire[1:0] w_n3522_0;
	wire[1:0] w_n3523_0;
	wire[1:0] w_n3527_0;
	wire[1:0] w_n3528_0;
	wire[1:0] w_n3531_0;
	wire[1:0] w_n3533_0;
	wire[1:0] w_n3534_0;
	wire[1:0] w_n3537_0;
	wire[1:0] w_n3540_0;
	wire[1:0] w_n3541_0;
	wire[1:0] w_n3543_0;
	wire[1:0] w_n3547_0;
	wire[1:0] w_n3549_0;
	wire[1:0] w_n3557_0;
	wire[1:0] w_n3559_0;
	wire[1:0] w_n3563_0;
	wire[1:0] w_n3567_0;
	wire[1:0] w_n3568_0;
	wire[1:0] w_n3571_0;
	wire[1:0] w_n3572_0;
	wire[1:0] w_n3576_0;
	wire[1:0] w_n3579_0;
	wire[1:0] w_n3580_0;
	wire[1:0] w_n3581_0;
	wire[1:0] w_n3584_0;
	wire[1:0] w_n3585_0;
	wire[1:0] w_n3588_0;
	wire[1:0] w_n3589_0;
	wire[1:0] w_n3593_0;
	wire[1:0] w_n3596_0;
	wire[1:0] w_n3597_0;
	wire[1:0] w_n3598_0;
	wire[1:0] w_n3601_0;
	wire[1:0] w_n3604_0;
	wire[1:0] w_n3605_0;
	wire[1:0] w_n3609_0;
	wire[1:0] w_n3612_0;
	wire[1:0] w_n3613_0;
	wire[1:0] w_n3615_0;
	wire[1:0] w_n3619_0;
	wire[1:0] w_n3620_0;
	wire[1:0] w_n3623_0;
	wire[1:0] w_n3624_0;
	wire[1:0] w_n3628_0;
	wire[1:0] w_n3631_0;
	wire[1:0] w_n3632_0;
	wire[1:0] w_n3633_0;
	wire[1:0] w_n3636_0;
	wire[1:0] w_n3639_0;
	wire[1:0] w_n3640_0;
	wire[1:0] w_n3641_0;
	wire[1:0] w_n3642_0;
	wire[1:0] w_n3643_0;
	wire[1:0] w_n3647_0;
	wire[1:0] w_n3650_0;
	wire[1:0] w_n3651_0;
	wire[1:0] w_n3652_0;
	wire[1:0] w_n3655_0;
	wire[1:0] w_n3658_0;
	wire[1:0] w_n3659_0;
	wire[1:0] w_n3660_0;
	wire[1:0] w_n3663_0;
	wire[1:0] w_n3666_0;
	wire[1:0] w_n3667_0;
	wire[1:0] w_n3668_0;
	wire[1:0] w_n3672_0;
	wire[1:0] w_n3675_0;
	wire[1:0] w_n3676_0;
	wire[1:0] w_n3677_0;
	wire[1:0] w_n3680_0;
	wire[1:0] w_n3683_0;
	wire[1:0] w_n3684_0;
	wire[1:0] w_n3685_0;
	wire[1:0] w_n3688_0;
	wire[1:0] w_n3689_0;
	wire[1:0] w_n3692_0;
	wire[1:0] w_n3693_0;
	wire[1:0] w_n3695_0;
	wire[1:0] w_n3696_0;
	wire[1:0] w_n3699_0;
	wire[1:0] w_n3700_0;
	wire[1:0] w_n3703_0;
	wire[1:0] w_n3704_0;
	wire[1:0] w_n3708_0;
	wire[1:0] w_n3711_0;
	wire[1:0] w_n3712_0;
	wire[1:0] w_n3713_0;
	wire[1:0] w_n3716_0;
	wire[1:0] w_n3719_0;
	wire[1:0] w_n3720_0;
	wire[1:0] w_n3721_0;
	wire[1:0] w_n3725_0;
	wire[1:0] w_n3728_0;
	wire[1:0] w_n3729_0;
	wire[1:0] w_n3730_0;
	wire[1:0] w_n3733_0;
	wire[1:0] w_n3734_0;
	wire[1:0] w_n3737_0;
	wire[1:0] w_n3738_0;
	wire[1:0] w_n3741_0;
	wire[1:0] w_n3744_0;
	wire[1:0] w_n3745_0;
	wire[1:0] w_n3746_0;
	wire[1:0] w_n3748_0;
	wire[1:0] w_n3749_0;
	wire[1:0] w_n3752_0;
	wire[1:0] w_n3755_0;
	wire[1:0] w_n3756_0;
	wire[1:0] w_n3757_0;
	wire[2:0] w_n3761_0;
	wire[1:0] w_n3764_0;
	wire[1:0] w_n3771_0;
	wire[1:0] w_n3776_0;
	wire[2:0] w_n3779_0;
	wire[1:0] w_n3787_0;
	wire[1:0] w_n3790_0;
	wire[2:0] w_n3791_0;
	wire[1:0] w_n3795_0;
	wire[1:0] w_n3798_0;
	wire[1:0] w_n3804_0;
	wire[1:0] w_n3806_0;
	wire[1:0] w_n3808_0;
	wire[1:0] w_n3811_0;
	wire[1:0] w_n3812_0;
	wire[1:0] w_n3817_0;
	wire[1:0] w_n3820_0;
	wire[1:0] w_n3821_0;
	wire[1:0] w_n3822_0;
	wire[1:0] w_n3826_0;
	wire[1:0] w_n3827_0;
	wire[1:0] w_n3830_0;
	wire[1:0] w_n3834_0;
	wire[1:0] w_n3835_0;
	wire[1:0] w_n3838_0;
	wire[1:0] w_n3840_0;
	wire[1:0] w_n3843_0;
	wire[1:0] w_n3845_0;
	wire[1:0] w_n3847_0;
	wire[1:0] w_n3853_0;
	wire[1:0] w_n3855_0;
	wire[1:0] w_n3857_0;
	wire[1:0] w_n3860_0;
	wire[1:0] w_n3861_0;
	wire[1:0] w_n3866_0;
	wire[1:0] w_n3869_0;
	wire[1:0] w_n3870_0;
	wire[1:0] w_n3871_0;
	wire[1:0] w_n3875_0;
	wire[1:0] w_n3876_0;
	wire[1:0] w_n3879_0;
	wire[1:0] w_n3881_0;
	wire[1:0] w_n3883_0;
	wire[1:0] w_n3890_0;
	wire[1:0] w_n3893_0;
	wire[1:0] w_n3894_0;
	wire[1:0] w_n3895_0;
	wire[1:0] w_n3898_0;
	wire[1:0] w_n3900_0;
	wire[1:0] w_n3902_0;
	wire[1:0] w_n3907_0;
	wire[1:0] w_n3909_0;
	wire[1:0] w_n3911_0;
	wire[1:0] w_n3914_0;
	wire[1:0] w_n3915_0;
	wire[1:0] w_n3918_0;
	wire[1:0] w_n3922_0;
	wire[1:0] w_n3923_0;
	wire[1:0] w_n3926_0;
	wire[1:0] w_n3928_0;
	wire[1:0] w_n3931_0;
	wire[1:0] w_n3933_0;
	wire[1:0] w_n3935_0;
	wire[1:0] w_n3941_0;
	wire[1:0] w_n3942_0;
	wire[1:0] w_n3945_0;
	wire[1:0] w_n3947_0;
	wire[1:0] w_n3949_0;
	wire[1:0] w_n3952_0;
	wire[1:0] w_n3954_0;
	wire[1:0] w_n3956_0;
	wire[1:0] w_n3960_0;
	wire[1:0] w_n3965_0;
	wire[1:0] w_n3972_0;
	wire[1:0] w_n3975_0;
	wire[1:0] w_n3976_0;
	wire[1:0] w_n3977_0;
	wire[1:0] w_n3980_0;
	wire[1:0] w_n3983_0;
	wire[1:0] w_n3984_0;
	wire[1:0] w_n3988_0;
	wire[1:0] w_n3991_0;
	wire[1:0] w_n3992_0;
	wire[1:0] w_n3997_0;
	wire[1:0] w_n4000_0;
	wire[1:0] w_n4002_0;
	wire[1:0] w_n4005_0;
	wire[1:0] w_n4008_0;
	wire[1:0] w_n4013_0;
	wire[1:0] w_n4015_0;
	wire[1:0] w_n4021_0;
	wire[1:0] w_n4023_0;
	wire[1:0] w_n4028_0;
	wire[1:0] w_n4034_0;
	wire[1:0] w_n4037_0;
	wire[1:0] w_n4038_0;
	wire[1:0] w_n4042_0;
	wire[1:0] w_n4043_0;
	wire[1:0] w_n4046_0;
	wire[1:0] w_n4048_0;
	wire[1:0] w_n4051_0;
	wire[1:0] w_n4052_0;
	wire[1:0] w_n4055_0;
	wire[1:0] w_n4059_0;
	wire[1:0] w_n4062_0;
	wire[1:0] w_n4063_0;
	wire[1:0] w_n4065_0;
	wire[1:0] w_n4066_0;
	wire[1:0] w_n4070_0;
	wire[1:0] w_n4071_0;
	wire[1:0] w_n4074_0;
	wire[1:0] w_n4076_0;
	wire[1:0] w_n4079_0;
	wire[1:0] w_n4080_0;
	wire[1:0] w_n4083_0;
	wire[1:0] w_n4087_0;
	wire[1:0] w_n4090_0;
	wire[1:0] w_n4091_0;
	wire[1:0] w_n4092_0;
	wire[1:0] w_n4096_0;
	wire[1:0] w_n4099_0;
	wire[1:0] w_n4101_0;
	wire[1:0] w_n4104_0;
	wire[1:0] w_n4108_0;
	wire[1:0] w_n4110_0;
	wire[1:0] w_n4114_0;
	wire[1:0] w_n4116_0;
	wire[1:0] w_n4125_0;
	wire[1:0] w_n4129_0;
	wire[1:0] w_n4133_0;
	wire[1:0] w_n4136_0;
	wire[1:0] w_n4138_0;
	wire[1:0] w_n4143_0;
	wire[1:0] w_n4145_0;
	wire[1:0] w_n4149_0;
	wire[1:0] w_n4153_0;
	wire[1:0] w_n4155_0;
	wire[1:0] w_n4158_0;
	wire[1:0] w_n4160_0;
	wire[1:0] w_n4162_0;
	wire[1:0] w_n4165_0;
	wire[1:0] w_n4167_0;
	wire[1:0] w_n4172_0;
	wire[1:0] w_n4173_0;
	wire[1:0] w_n4176_0;
	wire[1:0] w_n4181_0;
	wire[1:0] w_n4184_0;
	wire[1:0] w_n4185_0;
	wire[1:0] w_n4189_0;
	wire[1:0] w_n4190_0;
	wire[1:0] w_n4193_0;
	wire[1:0] w_n4196_0;
	wire[1:0] w_n4199_0;
	wire[1:0] w_n4202_0;
	wire[1:0] w_n4203_0;
	wire[1:0] w_n4205_0;
	wire[1:0] w_n4207_0;
	wire[1:0] w_n4210_0;
	wire[1:0] w_n4212_0;
	wire[1:0] w_n4214_0;
	wire[1:0] w_n4217_0;
	wire[1:0] w_n4222_0;
	wire[1:0] w_n4227_0;
	wire[1:0] w_n4229_0;
	wire[1:0] w_n4234_0;
	wire[1:0] w_n4236_0;
	wire[1:0] w_n4240_0;
	wire[1:0] w_n4245_0;
	wire[1:0] w_n4248_0;
	wire[1:0] w_n4251_0;
	wire[1:0] w_n4255_0;
	wire[1:0] w_n4259_0;
	wire[1:0] w_n4261_0;
	wire[1:0] w_n4266_0;
	wire[1:0] w_n4269_0;
	wire[1:0] w_n4272_0;
	wire[1:0] w_n4275_0;
	wire[1:0] w_n4280_0;
	wire[1:0] w_n4285_0;
	wire[1:0] w_n4287_0;
	wire[1:0] w_n4292_0;
	wire[1:0] w_n4294_0;
	wire[1:0] w_n4298_0;
	wire[1:0] w_n4302_0;
	wire[1:0] w_n4305_0;
	wire[1:0] w_n4308_0;
	wire[1:0] w_n4311_0;
	wire[1:0] w_n4316_0;
	wire[1:0] w_n4321_0;
	wire[1:0] w_n4323_0;
	wire[1:0] w_n4328_0;
	wire[1:0] w_n4330_0;
	wire[1:0] w_n4334_0;
	wire[1:0] w_n4338_0;
	wire[1:0] w_n4341_0;
	wire[1:0] w_n4344_0;
	wire[1:0] w_n4347_0;
	wire[1:0] w_n4352_0;
	wire[1:0] w_n4357_0;
	wire[1:0] w_n4359_0;
	wire[1:0] w_n4362_0;
	wire[1:0] w_n4368_0;
	wire[1:0] w_n4371_0;
	wire[1:0] w_n4372_0;
	wire[1:0] w_n4373_0;
	wire[1:0] w_n4374_0;
	wire[1:0] w_n4378_0;
	wire[1:0] w_n4379_0;
	wire[1:0] w_n4382_0;
	wire[1:0] w_n4384_0;
	wire[1:0] w_n4387_0;
	wire[1:0] w_n4388_0;
	wire[1:0] w_n4391_0;
	wire[1:0] w_n4394_0;
	wire[1:0] w_n4397_0;
	wire[1:0] w_n4400_0;
	wire[1:0] w_n4403_0;
	wire[1:0] w_n4407_0;
	wire[1:0] w_n4411_0;
	wire[1:0] w_n4413_0;
	wire[1:0] w_n4418_0;
	wire[1:0] w_n4419_0;
	wire[1:0] w_n4422_0;
	wire[1:0] w_n4427_0;
	wire[1:0] w_n4430_0;
	wire[1:0] w_n4431_0;
	wire[1:0] w_n4435_0;
	wire[1:0] w_n4436_0;
	wire[1:0] w_n4439_0;
	wire[1:0] w_n4442_0;
	wire[1:0] w_n4445_0;
	wire[1:0] w_n4448_0;
	wire[1:0] w_n4449_0;
	wire[1:0] w_n4451_0;
	wire[1:0] w_n4453_0;
	wire[1:0] w_n4456_0;
	wire[1:0] w_n4458_0;
	wire[1:0] w_n4460_0;
	wire[1:0] w_n4463_0;
	wire[1:0] w_n4468_0;
	wire[1:0] w_n4473_0;
	wire[1:0] w_n4503_0;
	wire[2:0] w_n4506_0;
	wire[2:0] w_n4515_0;
	wire[1:0] w_n4518_0;
	wire[1:0] w_n4526_0;
	wire[1:0] w_n4644_0;
	wire[2:0] w_n4648_0;
	wire[2:0] w_n4648_1;
	wire[2:0] w_n4648_2;
	wire[2:0] w_n4648_3;
	wire[2:0] w_n4648_4;
	wire[2:0] w_n4648_5;
	wire[2:0] w_n4648_6;
	wire[2:0] w_n4648_7;
	wire[2:0] w_n4648_8;
	wire[2:0] w_n4648_9;
	wire[2:0] w_n4648_10;
	wire[2:0] w_n4648_11;
	wire[2:0] w_n4648_12;
	wire[2:0] w_n4648_13;
	wire[2:0] w_n4648_14;
	wire[2:0] w_n4648_15;
	wire[2:0] w_n4648_16;
	wire[2:0] w_n4648_17;
	wire[2:0] w_n4648_18;
	wire[2:0] w_n4648_19;
	wire[2:0] w_n4648_20;
	wire[2:0] w_n4648_21;
	wire[2:0] w_n4648_22;
	wire[2:0] w_n4648_23;
	wire[2:0] w_n4648_24;
	wire[2:0] w_n4648_25;
	wire[2:0] w_n4648_26;
	wire[2:0] w_n4648_27;
	wire[2:0] w_n4648_28;
	wire[2:0] w_n4648_29;
	wire[2:0] w_n4648_30;
	wire[2:0] w_n4648_31;
	wire[2:0] w_n4648_32;
	wire[2:0] w_n4648_33;
	wire[2:0] w_n4648_34;
	wire[2:0] w_n4648_35;
	wire[2:0] w_n4648_36;
	wire[2:0] w_n4648_37;
	wire[2:0] w_n4648_38;
	wire[2:0] w_n4648_39;
	wire[2:0] w_n4648_40;
	wire[2:0] w_n4648_41;
	wire[2:0] w_n4648_42;
	wire[2:0] w_n4648_43;
	wire[2:0] w_n4648_44;
	wire[2:0] w_n4648_45;
	wire[2:0] w_n4648_46;
	wire[2:0] w_n4648_47;
	wire[2:0] w_n4648_48;
	wire[2:0] w_n4648_49;
	wire[2:0] w_n4648_50;
	wire[2:0] w_n4648_51;
	wire[2:0] w_n4648_52;
	wire[2:0] w_n4648_53;
	wire[2:0] w_n4648_54;
	wire[2:0] w_n4648_55;
	wire[2:0] w_n4648_56;
	wire[2:0] w_n4648_57;
	wire[2:0] w_n4648_58;
	wire[2:0] w_n4648_59;
	wire[2:0] w_n4648_60;
	wire[2:0] w_n4648_61;
	wire[2:0] w_n4648_62;
	wire[1:0] w_n4648_63;
	wire w_dff_A_4jf92R4g9_2;
	wire w_dff_A_WvrfUvCs4_0;
	wire w_dff_A_w2HmUyZ48_0;
	wire w_dff_A_cEcZOE7F6_0;
	wire w_dff_A_vRk2r0SD6_0;
	wire w_dff_A_qewfvzh80_0;
	wire w_dff_A_LulQbJwz3_0;
	wire w_dff_A_cYvKdfOF7_0;
	wire w_dff_A_9kGlvLfv2_0;
	wire w_dff_A_KiKbdZ2f2_0;
	wire w_dff_A_Bb0zsgpd0_0;
	wire w_dff_A_NyxQ7mA05_0;
	wire w_dff_A_X6eyEOAP9_0;
	wire w_dff_A_k0ryneHL6_0;
	wire w_dff_A_AHlgEB6R8_0;
	wire w_dff_A_nDuQPgox8_0;
	wire w_dff_A_RkK6Y4jk9_0;
	wire w_dff_A_Mva2ZKpy1_0;
	wire w_dff_A_NM8nigdI3_0;
	wire w_dff_A_LSf5wbfi1_0;
	wire w_dff_A_MlsONPWJ1_0;
	wire w_dff_A_7llmVHmU1_0;
	wire w_dff_A_2EwzNxVk7_0;
	wire w_dff_A_uyTbEu456_0;
	wire w_dff_A_73IGuFAb6_0;
	wire w_dff_A_164mSSGv9_0;
	wire w_dff_A_r8wBZGB90_0;
	wire w_dff_A_zxTqd09L3_0;
	wire w_dff_A_ZfBg7EOm3_0;
	wire w_dff_A_eAoBdlQn5_0;
	wire w_dff_A_UxAkDqS77_0;
	wire w_dff_A_GUFhpf3f0_0;
	wire w_dff_A_C2haGvds5_0;
	wire w_dff_A_iFd7aNBs5_0;
	wire w_dff_A_NUwyw1zB8_0;
	wire w_dff_A_oW4Z1SBK2_0;
	wire w_dff_A_GkCBajpz2_0;
	wire w_dff_A_24eK7md31_0;
	wire w_dff_A_MQhPxitl4_0;
	wire w_dff_A_WemNEdjD0_0;
	wire w_dff_A_BjmyDr9S7_0;
	wire w_dff_A_79a9Un1M3_0;
	wire w_dff_A_ZgAAD1X23_0;
	wire w_dff_A_W0hJcJng0_0;
	wire w_dff_A_15VK5Byw3_0;
	wire w_dff_A_YXQp2haH1_0;
	wire w_dff_A_R013b8kh1_0;
	wire w_dff_A_LcCBDxSe1_0;
	wire w_dff_A_5wIbKRAj5_0;
	wire w_dff_A_0QxsLgfB0_0;
	wire w_dff_A_3jFrOwCd1_0;
	wire w_dff_A_y9jp4VX77_0;
	wire w_dff_A_4Qlnpg9M5_0;
	wire w_dff_A_uYaPzqZA3_0;
	wire w_dff_A_kq1RummO1_0;
	wire w_dff_A_GfhJdHXK4_0;
	wire w_dff_A_vEYKv4WB4_0;
	wire w_dff_A_CDjyd4pp2_0;
	wire w_dff_A_jmRc3lFI4_0;
	wire w_dff_A_vw8shElw8_0;
	wire w_dff_A_y3Lzx6BD0_0;
	wire w_dff_A_SP5SySG57_0;
	wire w_dff_A_2moUPmxi5_0;
	wire w_dff_A_X19Xa4qX4_0;
	wire w_dff_A_DiDjfcNx9_0;
	wire w_dff_A_gJQ7MzSx4_0;
	wire w_dff_A_frWp3oTl2_0;
	wire w_dff_A_zHUiaLRr5_0;
	wire w_dff_A_EUKunzJq7_0;
	wire w_dff_A_oQwMs0mW5_0;
	wire w_dff_A_LSKIU1R72_0;
	wire w_dff_A_YUFMEqV59_0;
	wire w_dff_A_T9pDQtWE9_0;
	wire w_dff_A_t1ixKgFx5_0;
	wire w_dff_A_AGuJGsML4_0;
	wire w_dff_A_Q2yISQDn5_0;
	wire w_dff_A_6ukHgAXp8_0;
	wire w_dff_A_zxbKaZ869_0;
	wire w_dff_A_24sfdZXr3_0;
	wire w_dff_A_GhuuM4nu2_0;
	wire w_dff_A_vKtwxVRJ5_0;
	wire w_dff_A_JXDjRnst9_0;
	wire w_dff_A_4TbC2bHw6_0;
	wire w_dff_A_uYSMAWWk0_0;
	wire w_dff_A_SJgKgLkE7_0;
	wire w_dff_A_VTeFanvL9_0;
	wire w_dff_A_sMHiCaPq4_0;
	wire w_dff_A_6janH4c82_0;
	wire w_dff_A_7jRGideT8_0;
	wire w_dff_A_dO38tszJ1_0;
	wire w_dff_A_ruoAbtlZ9_0;
	wire w_dff_A_4fiXhAXU2_0;
	wire w_dff_A_egevUpLL9_0;
	wire w_dff_A_Nhdw7Kox2_0;
	wire w_dff_A_rhyNALCV1_0;
	wire w_dff_A_E9BTpH219_0;
	wire w_dff_A_vKsq5QJb0_0;
	wire w_dff_A_AgztGxiK8_0;
	wire w_dff_A_t4IJCiJa6_0;
	wire w_dff_A_N2ne8qw09_0;
	wire w_dff_A_G7kqdhof8_0;
	wire w_dff_A_FBvnzSKB4_0;
	wire w_dff_A_L0pTsOk01_0;
	wire w_dff_A_i7MpsIXU1_0;
	wire w_dff_A_Nx3X5url6_0;
	wire w_dff_A_fUFtcc7W4_0;
	wire w_dff_A_fKGTRAXk4_0;
	wire w_dff_A_TrFMigrB8_0;
	wire w_dff_A_oY4d4AN77_0;
	wire w_dff_A_4rHXoMaq5_0;
	wire w_dff_A_ne5OJtTS8_0;
	wire w_dff_A_TybogAPB0_0;
	wire w_dff_A_7an3FYwm6_0;
	wire w_dff_A_KVbc8xCN0_0;
	wire w_dff_A_LfXOHS0O4_0;
	wire w_dff_A_4NFpnNuN3_0;
	wire w_dff_A_y4WunLpr2_0;
	wire w_dff_A_rkjJcYFu4_0;
	wire w_dff_A_btioAenC8_0;
	wire w_dff_A_zMWFq7u72_0;
	wire w_dff_A_5J0aoye44_0;
	wire w_dff_A_JnTC9t918_0;
	wire w_dff_A_fuigrAIF3_0;
	wire w_dff_A_k0vpDHaf5_0;
	wire w_dff_A_n2Og61yG7_0;
	wire w_dff_A_BwaUDQlb7_0;
	wire w_dff_A_jvIRd8RD9_0;
	wire w_dff_A_t6DmL0hs4_0;
	wire w_dff_A_vKttdw0P8_0;
	wire w_dff_A_zil5QNhd3_0;
	wire w_dff_A_eChi8Hp90_0;
	wire w_dff_A_h8NfFE6T9_0;
	wire w_dff_A_WxOwicXM7_0;
	wire w_dff_A_53ozTV0t8_0;
	wire w_dff_A_sHAhLXI65_0;
	wire w_dff_A_p6cK4d8e3_0;
	wire w_dff_A_cNAUyyp40_0;
	wire w_dff_A_B0ajDMg55_0;
	wire w_dff_A_bDDsIjFK5_0;
	wire w_dff_A_zWmd4dhB0_0;
	wire w_dff_A_dFzYkT2w9_0;
	wire w_dff_A_WwnrpaUb3_0;
	wire w_dff_A_jCq1zhJR6_0;
	wire w_dff_A_3DB2Aomd0_0;
	wire w_dff_A_0MeMQ0W84_0;
	wire w_dff_A_rMxVGIVT7_0;
	wire w_dff_A_xWgZWwKi6_0;
	wire w_dff_A_OxDGxcuy0_0;
	wire w_dff_A_BAHS0BlU4_0;
	wire w_dff_A_1ur5BZkO0_0;
	wire w_dff_A_zU2Az30p3_0;
	wire w_dff_A_pxdk0SaI5_0;
	wire w_dff_A_IufjhC9z3_0;
	wire w_dff_A_bUxsefr51_0;
	wire w_dff_A_Nfv1pWz89_0;
	wire w_dff_A_Mi6vWPQd2_0;
	wire w_dff_A_iZRgV53k8_0;
	wire w_dff_A_y9cqJ74O8_0;
	wire w_dff_A_Yb7ypwXw3_0;
	wire w_dff_A_ObOVeJRp9_0;
	wire w_dff_A_KrQIAAHE3_0;
	wire w_dff_A_aoGDhvui2_0;
	wire w_dff_A_KM4GCFim7_0;
	wire w_dff_A_kGuuD0dn6_0;
	wire w_dff_A_TpFMWBtX0_0;
	wire w_dff_A_8ByzbrMU2_0;
	wire w_dff_A_AabcLQEi4_0;
	wire w_dff_A_rTZdbN3s7_0;
	wire w_dff_A_ck0PEhff7_0;
	wire w_dff_A_cpY2kb4V7_0;
	wire w_dff_A_p1PukFDF4_0;
	wire w_dff_A_mVDadcX61_0;
	wire w_dff_A_dy2I0UeI4_0;
	wire w_dff_A_cLy6gKfo5_0;
	wire w_dff_A_PRxsZe801_0;
	wire w_dff_A_sicOs0hc7_0;
	wire w_dff_A_dSVYS6Sb0_0;
	wire w_dff_A_Y9MPNg2g7_0;
	wire w_dff_A_ENC5HKRE6_0;
	wire w_dff_A_rTDKpKiJ5_0;
	wire w_dff_A_n1KDeIFP5_0;
	wire w_dff_A_QrykYaRi5_0;
	wire w_dff_A_tX8FSWOw9_0;
	wire w_dff_A_unj9VdsQ4_0;
	wire w_dff_A_y7AeHnxY2_0;
	wire w_dff_A_suiUbgLz3_0;
	wire w_dff_A_Nt1BUMao2_0;
	wire w_dff_A_E1qwy4311_0;
	wire w_dff_A_FEoc5rfZ4_0;
	wire w_dff_A_zAIw19Ld1_0;
	wire w_dff_A_gbW1I6Xw7_0;
	wire w_dff_A_fjV7yB6Y1_0;
	wire w_dff_A_u9eCVOjx8_0;
	wire w_dff_A_vxbIwSN15_0;
	wire w_dff_A_habLXnNM8_0;
	wire w_dff_A_HpcRdr2p2_0;
	wire w_dff_A_JpdZBD5e9_0;
	wire w_dff_A_CxWhO9FU8_0;
	wire w_dff_A_uZPd6kIb3_0;
	wire w_dff_A_mypM8eLS6_0;
	wire w_dff_A_426B4d8m3_0;
	wire w_dff_A_hYPFUOh12_0;
	wire w_dff_A_jPWtj9QZ3_0;
	wire w_dff_A_pHcPiXMP2_0;
	wire w_dff_A_0brnFmns3_0;
	wire w_dff_A_i4dkcnEv4_0;
	wire w_dff_A_1ZsJQvPo9_0;
	wire w_dff_A_CfvqN9Yh0_0;
	wire w_dff_A_gVxwUDTJ2_0;
	wire w_dff_A_VSKG0pS21_0;
	wire w_dff_A_m6FTD2XC1_0;
	wire w_dff_A_IUnjpRHq6_0;
	wire w_dff_A_J7blzP2R6_2;
	wire w_dff_A_PyOOYhAQ5_0;
	jnot g0000(.din(w_in1123_0[1]),.dout(n642),.clk(gclk));
	jand g0001(.dina(w_n642_0[1]),.dinb(w_in0123_0[1]),.dout(n643),.clk(gclk));
	jnot g0002(.din(w_n643_0[1]),.dout(n644),.clk(gclk));
	jnot g0003(.din(w_in0120_0[1]),.dout(n645),.clk(gclk));
	jand g0004(.dina(w_in1120_0[1]),.dinb(w_n645_0[1]),.dout(n646),.clk(gclk));
	jnot g0005(.din(w_in0121_0[1]),.dout(n647),.clk(gclk));
	jand g0006(.dina(w_in1121_0[1]),.dinb(w_n647_0[1]),.dout(n648),.clk(gclk));
	jor g0007(.dina(w_n648_0[1]),.dinb(n646),.dout(n649),.clk(gclk));
	jnot g0008(.din(w_in0118_0[1]),.dout(n650),.clk(gclk));
	jand g0009(.dina(w_in1118_0[1]),.dinb(w_n650_0[1]),.dout(n651),.clk(gclk));
	jnot g0010(.din(w_in0119_0[1]),.dout(n652),.clk(gclk));
	jand g0011(.dina(w_in1119_0[1]),.dinb(w_n652_0[1]),.dout(n653),.clk(gclk));
	jnot g0012(.din(w_in0117_0[1]),.dout(n654),.clk(gclk));
	jand g0013(.dina(w_in1117_0[1]),.dinb(w_n654_0[1]),.dout(n655),.clk(gclk));
	jor g0014(.dina(n655),.dinb(w_n653_0[1]),.dout(n656),.clk(gclk));
	jor g0015(.dina(n656),.dinb(n651),.dout(n657),.clk(gclk));
	jnot g0016(.din(w_n657_0[1]),.dout(n658),.clk(gclk));
	jnot g0017(.din(w_in1117_0[0]),.dout(n659),.clk(gclk));
	jand g0018(.dina(w_n659_0[1]),.dinb(w_in0117_0[0]),.dout(n660),.clk(gclk));
	jnot g0019(.din(w_in1116_0[1]),.dout(n661),.clk(gclk));
	jand g0020(.dina(w_n661_0[1]),.dinb(w_in0116_0[1]),.dout(n662),.clk(gclk));
	jor g0021(.dina(n662),.dinb(n660),.dout(n663),.clk(gclk));
	jand g0022(.dina(n663),.dinb(n658),.dout(n664),.clk(gclk));
	jnot g0023(.din(w_n653_0[0]),.dout(n665),.clk(gclk));
	jnot g0024(.din(w_in1119_0[0]),.dout(n666),.clk(gclk));
	jand g0025(.dina(w_n666_0[1]),.dinb(w_in0119_0[0]),.dout(n667),.clk(gclk));
	jnot g0026(.din(w_in1118_0[0]),.dout(n668),.clk(gclk));
	jand g0027(.dina(w_n668_0[1]),.dinb(w_in0118_0[0]),.dout(n669),.clk(gclk));
	jor g0028(.dina(n669),.dinb(n667),.dout(n670),.clk(gclk));
	jand g0029(.dina(n670),.dinb(n665),.dout(n671),.clk(gclk));
	jor g0030(.dina(n671),.dinb(n664),.dout(n672),.clk(gclk));
	jnot g0031(.din(w_n672_0[1]),.dout(n673),.clk(gclk));
	jnot g0032(.din(w_in1115_0[1]),.dout(n674),.clk(gclk));
	jand g0033(.dina(w_n674_0[1]),.dinb(w_in0115_0[1]),.dout(n675),.clk(gclk));
	jnot g0034(.din(w_n675_0[1]),.dout(n676),.clk(gclk));
	jnot g0035(.din(w_in0113_0[1]),.dout(n677),.clk(gclk));
	jand g0036(.dina(w_in1113_0[1]),.dinb(w_n677_0[1]),.dout(n678),.clk(gclk));
	jnot g0037(.din(w_in0112_0[1]),.dout(n679),.clk(gclk));
	jand g0038(.dina(w_in1112_0[1]),.dinb(w_n679_0[1]),.dout(n680),.clk(gclk));
	jor g0039(.dina(n680),.dinb(w_n678_0[1]),.dout(n681),.clk(gclk));
	jnot g0040(.din(w_in0110_0[1]),.dout(n682),.clk(gclk));
	jand g0041(.dina(w_in1110_0[1]),.dinb(w_n682_0[1]),.dout(n683),.clk(gclk));
	jnot g0042(.din(w_in0111_0[1]),.dout(n684),.clk(gclk));
	jand g0043(.dina(w_in1111_0[1]),.dinb(w_n684_0[1]),.dout(n685),.clk(gclk));
	jnot g0044(.din(w_in0109_0[1]),.dout(n686),.clk(gclk));
	jand g0045(.dina(w_in1109_0[1]),.dinb(w_n686_0[1]),.dout(n687),.clk(gclk));
	jor g0046(.dina(n687),.dinb(w_n685_0[1]),.dout(n688),.clk(gclk));
	jor g0047(.dina(n688),.dinb(n683),.dout(n689),.clk(gclk));
	jnot g0048(.din(w_n689_0[1]),.dout(n690),.clk(gclk));
	jnot g0049(.din(w_in1109_0[0]),.dout(n691),.clk(gclk));
	jand g0050(.dina(w_n691_0[1]),.dinb(w_in0109_0[0]),.dout(n692),.clk(gclk));
	jnot g0051(.din(w_in1108_0[1]),.dout(n693),.clk(gclk));
	jand g0052(.dina(w_n693_0[1]),.dinb(w_in0108_0[1]),.dout(n694),.clk(gclk));
	jor g0053(.dina(n694),.dinb(n692),.dout(n695),.clk(gclk));
	jand g0054(.dina(n695),.dinb(n690),.dout(n696),.clk(gclk));
	jnot g0055(.din(w_n685_0[0]),.dout(n697),.clk(gclk));
	jnot g0056(.din(w_in1111_0[0]),.dout(n698),.clk(gclk));
	jand g0057(.dina(w_n698_0[1]),.dinb(w_in0111_0[0]),.dout(n699),.clk(gclk));
	jnot g0058(.din(w_in1110_0[0]),.dout(n700),.clk(gclk));
	jand g0059(.dina(w_n700_0[1]),.dinb(w_in0110_0[0]),.dout(n701),.clk(gclk));
	jor g0060(.dina(n701),.dinb(n699),.dout(n702),.clk(gclk));
	jand g0061(.dina(n702),.dinb(n697),.dout(n703),.clk(gclk));
	jor g0062(.dina(n703),.dinb(n696),.dout(n704),.clk(gclk));
	jnot g0063(.din(w_n704_0[1]),.dout(n705),.clk(gclk));
	jnot g0064(.din(w_in1107_0[1]),.dout(n706),.clk(gclk));
	jand g0065(.dina(w_n706_0[1]),.dinb(w_in0107_0[1]),.dout(n707),.clk(gclk));
	jnot g0066(.din(w_n707_0[1]),.dout(n708),.clk(gclk));
	jnot g0067(.din(w_in0104_0[1]),.dout(n709),.clk(gclk));
	jand g0068(.dina(w_in1104_0[1]),.dinb(w_n709_0[1]),.dout(n710),.clk(gclk));
	jnot g0069(.din(w_in0105_0[1]),.dout(n711),.clk(gclk));
	jand g0070(.dina(w_in1105_0[1]),.dinb(w_n711_0[1]),.dout(n712),.clk(gclk));
	jor g0071(.dina(w_n712_0[1]),.dinb(n710),.dout(n713),.clk(gclk));
	jnot g0072(.din(w_in0102_0[1]),.dout(n714),.clk(gclk));
	jand g0073(.dina(w_in1102_0[1]),.dinb(w_n714_0[1]),.dout(n715),.clk(gclk));
	jnot g0074(.din(w_in0103_0[1]),.dout(n716),.clk(gclk));
	jand g0075(.dina(w_in1103_0[1]),.dinb(w_n716_0[1]),.dout(n717),.clk(gclk));
	jnot g0076(.din(w_in0101_0[1]),.dout(n718),.clk(gclk));
	jand g0077(.dina(w_in1101_0[1]),.dinb(w_n718_0[1]),.dout(n719),.clk(gclk));
	jor g0078(.dina(n719),.dinb(w_n717_0[1]),.dout(n720),.clk(gclk));
	jor g0079(.dina(n720),.dinb(n715),.dout(n721),.clk(gclk));
	jnot g0080(.din(w_n721_0[1]),.dout(n722),.clk(gclk));
	jnot g0081(.din(w_in1101_0[0]),.dout(n723),.clk(gclk));
	jand g0082(.dina(w_n723_0[1]),.dinb(w_in0101_0[0]),.dout(n724),.clk(gclk));
	jnot g0083(.din(w_in1100_0[1]),.dout(n725),.clk(gclk));
	jand g0084(.dina(w_n725_0[1]),.dinb(w_in0100_0[1]),.dout(n726),.clk(gclk));
	jor g0085(.dina(n726),.dinb(n724),.dout(n727),.clk(gclk));
	jand g0086(.dina(n727),.dinb(n722),.dout(n728),.clk(gclk));
	jnot g0087(.din(w_n717_0[0]),.dout(n729),.clk(gclk));
	jnot g0088(.din(w_in1103_0[0]),.dout(n730),.clk(gclk));
	jand g0089(.dina(w_n730_0[1]),.dinb(w_in0103_0[0]),.dout(n731),.clk(gclk));
	jnot g0090(.din(w_in1102_0[0]),.dout(n732),.clk(gclk));
	jand g0091(.dina(w_n732_0[1]),.dinb(w_in0102_0[0]),.dout(n733),.clk(gclk));
	jor g0092(.dina(n733),.dinb(n731),.dout(n734),.clk(gclk));
	jand g0093(.dina(n734),.dinb(n729),.dout(n735),.clk(gclk));
	jor g0094(.dina(n735),.dinb(n728),.dout(n736),.clk(gclk));
	jnot g0095(.din(w_n736_0[1]),.dout(n737),.clk(gclk));
	jnot g0096(.din(w_in199_0[1]),.dout(n738),.clk(gclk));
	jand g0097(.dina(w_n738_0[1]),.dinb(w_in099_0[1]),.dout(n739),.clk(gclk));
	jnot g0098(.din(w_n739_0[1]),.dout(n740),.clk(gclk));
	jnot g0099(.din(w_in097_0[1]),.dout(n741),.clk(gclk));
	jand g0100(.dina(w_in197_0[1]),.dinb(w_n741_0[1]),.dout(n742),.clk(gclk));
	jnot g0101(.din(w_in096_0[1]),.dout(n743),.clk(gclk));
	jand g0102(.dina(w_in196_0[1]),.dinb(w_n743_0[1]),.dout(n744),.clk(gclk));
	jor g0103(.dina(n744),.dinb(w_n742_0[1]),.dout(n745),.clk(gclk));
	jnot g0104(.din(w_in094_0[1]),.dout(n746),.clk(gclk));
	jand g0105(.dina(w_in194_0[1]),.dinb(w_n746_0[1]),.dout(n747),.clk(gclk));
	jnot g0106(.din(w_in095_0[1]),.dout(n748),.clk(gclk));
	jand g0107(.dina(w_in195_0[1]),.dinb(w_n748_0[1]),.dout(n749),.clk(gclk));
	jnot g0108(.din(w_in093_0[1]),.dout(n750),.clk(gclk));
	jand g0109(.dina(w_in193_0[1]),.dinb(w_n750_0[1]),.dout(n751),.clk(gclk));
	jor g0110(.dina(n751),.dinb(w_n749_0[1]),.dout(n752),.clk(gclk));
	jor g0111(.dina(n752),.dinb(n747),.dout(n753),.clk(gclk));
	jnot g0112(.din(w_n753_0[1]),.dout(n754),.clk(gclk));
	jnot g0113(.din(w_in193_0[0]),.dout(n755),.clk(gclk));
	jand g0114(.dina(w_n755_0[1]),.dinb(w_in093_0[0]),.dout(n756),.clk(gclk));
	jnot g0115(.din(w_in192_0[1]),.dout(n757),.clk(gclk));
	jand g0116(.dina(w_n757_0[1]),.dinb(w_in092_0[1]),.dout(n758),.clk(gclk));
	jor g0117(.dina(n758),.dinb(n756),.dout(n759),.clk(gclk));
	jand g0118(.dina(n759),.dinb(n754),.dout(n760),.clk(gclk));
	jnot g0119(.din(w_n749_0[0]),.dout(n761),.clk(gclk));
	jnot g0120(.din(w_in195_0[0]),.dout(n762),.clk(gclk));
	jand g0121(.dina(w_n762_0[1]),.dinb(w_in095_0[0]),.dout(n763),.clk(gclk));
	jnot g0122(.din(w_in194_0[0]),.dout(n764),.clk(gclk));
	jand g0123(.dina(w_n764_0[1]),.dinb(w_in094_0[0]),.dout(n765),.clk(gclk));
	jor g0124(.dina(n765),.dinb(n763),.dout(n766),.clk(gclk));
	jand g0125(.dina(n766),.dinb(n761),.dout(n767),.clk(gclk));
	jor g0126(.dina(n767),.dinb(n760),.dout(n768),.clk(gclk));
	jnot g0127(.din(w_n768_0[1]),.dout(n769),.clk(gclk));
	jnot g0128(.din(w_in191_0[1]),.dout(n770),.clk(gclk));
	jand g0129(.dina(w_n770_0[1]),.dinb(w_in091_0[1]),.dout(n771),.clk(gclk));
	jnot g0130(.din(w_n771_0[1]),.dout(n772),.clk(gclk));
	jnot g0131(.din(w_in086_0[1]),.dout(n773),.clk(gclk));
	jand g0132(.dina(w_in186_0[1]),.dinb(w_n773_0[1]),.dout(n774),.clk(gclk));
	jnot g0133(.din(w_in087_0[1]),.dout(n775),.clk(gclk));
	jand g0134(.dina(w_in187_0[1]),.dinb(w_n775_0[1]),.dout(n776),.clk(gclk));
	jnot g0135(.din(w_in085_0[1]),.dout(n777),.clk(gclk));
	jand g0136(.dina(w_in185_0[1]),.dinb(w_n777_0[1]),.dout(n778),.clk(gclk));
	jor g0137(.dina(n778),.dinb(w_n776_0[1]),.dout(n779),.clk(gclk));
	jor g0138(.dina(n779),.dinb(n774),.dout(n780),.clk(gclk));
	jnot g0139(.din(w_n780_0[1]),.dout(n781),.clk(gclk));
	jnot g0140(.din(w_in185_0[0]),.dout(n782),.clk(gclk));
	jand g0141(.dina(w_n782_0[1]),.dinb(w_in085_0[0]),.dout(n783),.clk(gclk));
	jnot g0142(.din(w_in184_0[1]),.dout(n784),.clk(gclk));
	jand g0143(.dina(w_n784_0[1]),.dinb(w_in084_0[1]),.dout(n785),.clk(gclk));
	jor g0144(.dina(n785),.dinb(n783),.dout(n786),.clk(gclk));
	jand g0145(.dina(n786),.dinb(n781),.dout(n787),.clk(gclk));
	jnot g0146(.din(w_n776_0[0]),.dout(n788),.clk(gclk));
	jnot g0147(.din(w_in187_0[0]),.dout(n789),.clk(gclk));
	jand g0148(.dina(w_n789_0[1]),.dinb(w_in087_0[0]),.dout(n790),.clk(gclk));
	jnot g0149(.din(w_in186_0[0]),.dout(n791),.clk(gclk));
	jand g0150(.dina(w_n791_0[1]),.dinb(w_in086_0[0]),.dout(n792),.clk(gclk));
	jor g0151(.dina(n792),.dinb(n790),.dout(n793),.clk(gclk));
	jand g0152(.dina(n793),.dinb(n788),.dout(n794),.clk(gclk));
	jor g0153(.dina(n794),.dinb(n787),.dout(n795),.clk(gclk));
	jnot g0154(.din(w_n795_0[1]),.dout(n796),.clk(gclk));
	jnot g0155(.din(w_in183_0[1]),.dout(n797),.clk(gclk));
	jand g0156(.dina(w_n797_0[1]),.dinb(w_in083_0[1]),.dout(n798),.clk(gclk));
	jnot g0157(.din(w_n798_0[1]),.dout(n799),.clk(gclk));
	jnot g0158(.din(w_in081_0[1]),.dout(n800),.clk(gclk));
	jand g0159(.dina(w_in181_0[1]),.dinb(w_n800_0[1]),.dout(n801),.clk(gclk));
	jnot g0160(.din(w_in080_0[1]),.dout(n802),.clk(gclk));
	jand g0161(.dina(w_in180_0[1]),.dinb(w_n802_0[1]),.dout(n803),.clk(gclk));
	jor g0162(.dina(n803),.dinb(w_n801_0[1]),.dout(n804),.clk(gclk));
	jnot g0163(.din(w_in078_0[1]),.dout(n805),.clk(gclk));
	jand g0164(.dina(w_in178_0[1]),.dinb(w_n805_0[1]),.dout(n806),.clk(gclk));
	jnot g0165(.din(w_in079_0[1]),.dout(n807),.clk(gclk));
	jand g0166(.dina(w_in179_0[1]),.dinb(w_n807_0[1]),.dout(n808),.clk(gclk));
	jnot g0167(.din(w_in077_0[1]),.dout(n809),.clk(gclk));
	jand g0168(.dina(w_in177_0[1]),.dinb(w_n809_0[1]),.dout(n810),.clk(gclk));
	jor g0169(.dina(n810),.dinb(w_n808_0[1]),.dout(n811),.clk(gclk));
	jor g0170(.dina(n811),.dinb(n806),.dout(n812),.clk(gclk));
	jnot g0171(.din(w_n812_0[1]),.dout(n813),.clk(gclk));
	jnot g0172(.din(w_in177_0[0]),.dout(n814),.clk(gclk));
	jand g0173(.dina(w_n814_0[1]),.dinb(w_in077_0[0]),.dout(n815),.clk(gclk));
	jnot g0174(.din(w_in176_0[1]),.dout(n816),.clk(gclk));
	jand g0175(.dina(w_n816_0[1]),.dinb(w_in076_0[1]),.dout(n817),.clk(gclk));
	jor g0176(.dina(n817),.dinb(n815),.dout(n818),.clk(gclk));
	jand g0177(.dina(n818),.dinb(n813),.dout(n819),.clk(gclk));
	jnot g0178(.din(w_n808_0[0]),.dout(n820),.clk(gclk));
	jnot g0179(.din(w_in179_0[0]),.dout(n821),.clk(gclk));
	jand g0180(.dina(w_n821_0[1]),.dinb(w_in079_0[0]),.dout(n822),.clk(gclk));
	jnot g0181(.din(w_in178_0[0]),.dout(n823),.clk(gclk));
	jand g0182(.dina(w_n823_0[1]),.dinb(w_in078_0[0]),.dout(n824),.clk(gclk));
	jor g0183(.dina(n824),.dinb(n822),.dout(n825),.clk(gclk));
	jand g0184(.dina(n825),.dinb(n820),.dout(n826),.clk(gclk));
	jor g0185(.dina(n826),.dinb(n819),.dout(n827),.clk(gclk));
	jnot g0186(.din(w_n827_0[1]),.dout(n828),.clk(gclk));
	jnot g0187(.din(w_in175_0[1]),.dout(n829),.clk(gclk));
	jand g0188(.dina(w_n829_0[1]),.dinb(w_in075_0[1]),.dout(n830),.clk(gclk));
	jnot g0189(.din(w_n830_0[1]),.dout(n831),.clk(gclk));
	jnot g0190(.din(w_in072_0[1]),.dout(n832),.clk(gclk));
	jand g0191(.dina(w_in172_0[1]),.dinb(w_n832_0[1]),.dout(n833),.clk(gclk));
	jnot g0192(.din(w_in073_0[1]),.dout(n834),.clk(gclk));
	jand g0193(.dina(w_in173_0[1]),.dinb(w_n834_0[1]),.dout(n835),.clk(gclk));
	jor g0194(.dina(w_n835_0[1]),.dinb(n833),.dout(n836),.clk(gclk));
	jnot g0195(.din(w_in070_0[1]),.dout(n837),.clk(gclk));
	jand g0196(.dina(w_in170_0[1]),.dinb(w_n837_0[1]),.dout(n838),.clk(gclk));
	jnot g0197(.din(w_in071_0[1]),.dout(n839),.clk(gclk));
	jand g0198(.dina(w_in171_0[1]),.dinb(w_n839_0[1]),.dout(n840),.clk(gclk));
	jnot g0199(.din(w_in069_0[1]),.dout(n841),.clk(gclk));
	jand g0200(.dina(w_in169_0[1]),.dinb(w_n841_0[1]),.dout(n842),.clk(gclk));
	jor g0201(.dina(n842),.dinb(w_n840_0[1]),.dout(n843),.clk(gclk));
	jor g0202(.dina(n843),.dinb(n838),.dout(n844),.clk(gclk));
	jnot g0203(.din(w_n844_0[1]),.dout(n845),.clk(gclk));
	jnot g0204(.din(w_in169_0[0]),.dout(n846),.clk(gclk));
	jand g0205(.dina(w_n846_0[1]),.dinb(w_in069_0[0]),.dout(n847),.clk(gclk));
	jnot g0206(.din(w_in168_0[1]),.dout(n848),.clk(gclk));
	jand g0207(.dina(w_n848_0[1]),.dinb(w_in068_0[1]),.dout(n849),.clk(gclk));
	jor g0208(.dina(n849),.dinb(n847),.dout(n850),.clk(gclk));
	jand g0209(.dina(n850),.dinb(n845),.dout(n851),.clk(gclk));
	jnot g0210(.din(w_n840_0[0]),.dout(n852),.clk(gclk));
	jnot g0211(.din(w_in171_0[0]),.dout(n853),.clk(gclk));
	jand g0212(.dina(w_n853_0[1]),.dinb(w_in071_0[0]),.dout(n854),.clk(gclk));
	jnot g0213(.din(w_in170_0[0]),.dout(n855),.clk(gclk));
	jand g0214(.dina(w_n855_0[1]),.dinb(w_in070_0[0]),.dout(n856),.clk(gclk));
	jor g0215(.dina(n856),.dinb(n854),.dout(n857),.clk(gclk));
	jand g0216(.dina(n857),.dinb(n852),.dout(n858),.clk(gclk));
	jor g0217(.dina(n858),.dinb(n851),.dout(n859),.clk(gclk));
	jnot g0218(.din(w_n859_0[1]),.dout(n860),.clk(gclk));
	jnot g0219(.din(w_in167_0[1]),.dout(n861),.clk(gclk));
	jand g0220(.dina(w_n861_0[1]),.dinb(w_in067_0[1]),.dout(n862),.clk(gclk));
	jnot g0221(.din(w_n862_0[1]),.dout(n863),.clk(gclk));
	jnot g0222(.din(w_in065_0[1]),.dout(n864),.clk(gclk));
	jand g0223(.dina(w_in165_0[1]),.dinb(w_n864_0[1]),.dout(n865),.clk(gclk));
	jnot g0224(.din(w_n865_0[1]),.dout(n866),.clk(gclk));
	jnot g0225(.din(w_in164_0[1]),.dout(n867),.clk(gclk));
	jand g0226(.dina(w_n867_0[1]),.dinb(w_in064_0[1]),.dout(n868),.clk(gclk));
	jand g0227(.dina(n868),.dinb(n866),.dout(n869),.clk(gclk));
	jnot g0228(.din(w_in166_0[1]),.dout(n870),.clk(gclk));
	jand g0229(.dina(w_n870_0[1]),.dinb(w_in066_0[1]),.dout(n871),.clk(gclk));
	jnot g0230(.din(w_in165_0[0]),.dout(n872),.clk(gclk));
	jand g0231(.dina(w_n872_0[1]),.dinb(w_in065_0[0]),.dout(n873),.clk(gclk));
	jor g0232(.dina(n873),.dinb(n871),.dout(n874),.clk(gclk));
	jor g0233(.dina(n874),.dinb(n869),.dout(n875),.clk(gclk));
	jnot g0234(.din(w_n875_0[1]),.dout(n876),.clk(gclk));
	jnot g0235(.din(w_in159_0[1]),.dout(n877),.clk(gclk));
	jnot g0236(.din(w_in060_0[1]),.dout(n878),.clk(gclk));
	jand g0237(.dina(w_in160_0[1]),.dinb(w_n878_0[1]),.dout(n879),.clk(gclk));
	jnot g0238(.din(w_in063_0[1]),.dout(n880),.clk(gclk));
	jand g0239(.dina(w_in163_0[1]),.dinb(w_n880_0[1]),.dout(n881),.clk(gclk));
	jnot g0240(.din(w_in061_0[1]),.dout(n882),.clk(gclk));
	jand g0241(.dina(w_in161_0[1]),.dinb(w_n882_0[1]),.dout(n883),.clk(gclk));
	jnot g0242(.din(w_in062_0[1]),.dout(n884),.clk(gclk));
	jand g0243(.dina(w_in162_0[1]),.dinb(w_n884_0[1]),.dout(n885),.clk(gclk));
	jor g0244(.dina(n885),.dinb(n883),.dout(n886),.clk(gclk));
	jor g0245(.dina(n886),.dinb(w_n881_0[1]),.dout(n887),.clk(gclk));
	jor g0246(.dina(w_n887_0[1]),.dinb(n879),.dout(n888),.clk(gclk));
	jnot g0247(.din(w_n888_0[1]),.dout(n889),.clk(gclk));
	jand g0248(.dina(n889),.dinb(w_in059_0[1]),.dout(n890),.clk(gclk));
	jand g0249(.dina(n890),.dinb(w_n877_0[1]),.dout(n891),.clk(gclk));
	jnot g0250(.din(w_n891_0[1]),.dout(n892),.clk(gclk));
	jnot g0251(.din(w_in151_0[1]),.dout(n893),.clk(gclk));
	jnot g0252(.din(w_in053_0[1]),.dout(n894),.clk(gclk));
	jand g0253(.dina(w_in153_0[1]),.dinb(w_n894_0[1]),.dout(n895),.clk(gclk));
	jnot g0254(.din(w_in055_0[1]),.dout(n896),.clk(gclk));
	jand g0255(.dina(w_in155_0[1]),.dinb(w_n896_0[1]),.dout(n897),.clk(gclk));
	jnot g0256(.din(w_in054_0[1]),.dout(n898),.clk(gclk));
	jand g0257(.dina(w_in154_0[1]),.dinb(w_n898_0[1]),.dout(n899),.clk(gclk));
	jor g0258(.dina(n899),.dinb(n897),.dout(n900),.clk(gclk));
	jnot g0259(.din(w_in052_0[1]),.dout(n901),.clk(gclk));
	jand g0260(.dina(w_in152_0[1]),.dinb(w_n901_0[1]),.dout(n902),.clk(gclk));
	jor g0261(.dina(n902),.dinb(w_n900_0[1]),.dout(n903),.clk(gclk));
	jor g0262(.dina(n903),.dinb(w_n895_0[1]),.dout(n904),.clk(gclk));
	jnot g0263(.din(w_n904_0[1]),.dout(n905),.clk(gclk));
	jand g0264(.dina(n905),.dinb(w_in051_0[1]),.dout(n906),.clk(gclk));
	jand g0265(.dina(n906),.dinb(w_n893_0[1]),.dout(n907),.clk(gclk));
	jnot g0266(.din(w_n907_0[1]),.dout(n908),.clk(gclk));
	jnot g0267(.din(w_in044_0[1]),.dout(n909),.clk(gclk));
	jand g0268(.dina(w_in144_0[1]),.dinb(w_n909_0[1]),.dout(n910),.clk(gclk));
	jnot g0269(.din(w_in047_0[1]),.dout(n911),.clk(gclk));
	jand g0270(.dina(w_in147_0[1]),.dinb(w_n911_0[1]),.dout(n912),.clk(gclk));
	jnot g0271(.din(w_in045_0[1]),.dout(n913),.clk(gclk));
	jand g0272(.dina(w_in145_0[1]),.dinb(w_n913_0[1]),.dout(n914),.clk(gclk));
	jnot g0273(.din(w_in046_0[1]),.dout(n915),.clk(gclk));
	jand g0274(.dina(w_in146_0[1]),.dinb(w_n915_0[1]),.dout(n916),.clk(gclk));
	jor g0275(.dina(n916),.dinb(n914),.dout(n917),.clk(gclk));
	jor g0276(.dina(n917),.dinb(w_n912_0[1]),.dout(n918),.clk(gclk));
	jor g0277(.dina(w_n918_0[1]),.dinb(n910),.dout(n919),.clk(gclk));
	jnot g0278(.din(w_in042_0[1]),.dout(n920),.clk(gclk));
	jand g0279(.dina(w_in142_0[1]),.dinb(w_n920_0[1]),.dout(n921),.clk(gclk));
	jnot g0280(.din(in043),.dout(n922),.clk(gclk));
	jand g0281(.dina(w_in143_0[2]),.dinb(w_n922_0[2]),.dout(n923),.clk(gclk));
	jor g0282(.dina(n923),.dinb(n921),.dout(n924),.clk(gclk));
	jor g0283(.dina(n924),.dinb(w_n919_0[1]),.dout(n925),.clk(gclk));
	jnot g0284(.din(w_n925_0[1]),.dout(n926),.clk(gclk));
	jnot g0285(.din(w_in142_0[0]),.dout(n927),.clk(gclk));
	jand g0286(.dina(w_n927_0[1]),.dinb(w_in042_0[0]),.dout(n928),.clk(gclk));
	jnot g0287(.din(w_in141_0[1]),.dout(n929),.clk(gclk));
	jand g0288(.dina(w_n929_0[1]),.dinb(w_in041_0[1]),.dout(n930),.clk(gclk));
	jnot g0289(.din(w_in041_0[0]),.dout(n931),.clk(gclk));
	jand g0290(.dina(w_in141_0[0]),.dinb(w_n931_0[1]),.dout(n932),.clk(gclk));
	jnot g0291(.din(w_n932_0[1]),.dout(n933),.clk(gclk));
	jnot g0292(.din(w_in140_0[1]),.dout(n934),.clk(gclk));
	jand g0293(.dina(w_n934_0[1]),.dinb(w_in040_0[1]),.dout(n935),.clk(gclk));
	jand g0294(.dina(n935),.dinb(n933),.dout(n936),.clk(gclk));
	jor g0295(.dina(n936),.dinb(n930),.dout(n937),.clk(gclk));
	jor g0296(.dina(n937),.dinb(n928),.dout(n938),.clk(gclk));
	jand g0297(.dina(n938),.dinb(n926),.dout(n939),.clk(gclk));
	jnot g0298(.din(w_n939_0[1]),.dout(n940),.clk(gclk));
	jnot g0299(.din(w_in133_0[1]),.dout(n941),.clk(gclk));
	jand g0300(.dina(w_n941_0[1]),.dinb(w_in033_0[1]),.dout(n942),.clk(gclk));
	jnot g0301(.din(w_in134_0[1]),.dout(n943),.clk(gclk));
	jand g0302(.dina(w_n943_0[1]),.dinb(w_in034_0[1]),.dout(n944),.clk(gclk));
	jor g0303(.dina(n944),.dinb(n942),.dout(n945),.clk(gclk));
	jnot g0304(.din(w_in033_0[0]),.dout(n946),.clk(gclk));
	jand g0305(.dina(w_in133_0[0]),.dinb(w_n946_0[1]),.dout(n947),.clk(gclk));
	jnot g0306(.din(w_n947_0[1]),.dout(n948),.clk(gclk));
	jnot g0307(.din(w_in132_0[1]),.dout(n949),.clk(gclk));
	jand g0308(.dina(w_n949_0[1]),.dinb(w_in032_0[1]),.dout(n950),.clk(gclk));
	jand g0309(.dina(n950),.dinb(n948),.dout(n951),.clk(gclk));
	jor g0310(.dina(n951),.dinb(n945),.dout(n952),.clk(gclk));
	jnot g0311(.din(w_in035_0[1]),.dout(n953),.clk(gclk));
	jand g0312(.dina(w_in135_0[1]),.dinb(w_n953_0[1]),.dout(n954),.clk(gclk));
	jnot g0313(.din(w_in034_0[0]),.dout(n955),.clk(gclk));
	jand g0314(.dina(w_in134_0[0]),.dinb(w_n955_0[1]),.dout(n956),.clk(gclk));
	jor g0315(.dina(n956),.dinb(n954),.dout(n957),.clk(gclk));
	jnot g0316(.din(w_in036_0[1]),.dout(n958),.clk(gclk));
	jand g0317(.dina(w_in136_0[1]),.dinb(w_n958_0[1]),.dout(n959),.clk(gclk));
	jnot g0318(.din(w_in038_0[1]),.dout(n960),.clk(gclk));
	jand g0319(.dina(w_in138_0[1]),.dinb(w_n960_0[1]),.dout(n961),.clk(gclk));
	jnot g0320(.din(w_in039_0[1]),.dout(n962),.clk(gclk));
	jand g0321(.dina(w_in139_0[1]),.dinb(w_n962_0[1]),.dout(n963),.clk(gclk));
	jnot g0322(.din(w_in037_0[1]),.dout(n964),.clk(gclk));
	jand g0323(.dina(w_in137_0[1]),.dinb(w_n964_0[1]),.dout(n965),.clk(gclk));
	jor g0324(.dina(n965),.dinb(w_n963_0[1]),.dout(n966),.clk(gclk));
	jor g0325(.dina(n966),.dinb(n961),.dout(n967),.clk(gclk));
	jor g0326(.dina(w_n967_0[1]),.dinb(n959),.dout(n968),.clk(gclk));
	jor g0327(.dina(w_n968_0[1]),.dinb(n957),.dout(n969),.clk(gclk));
	jnot g0328(.din(w_n969_0[1]),.dout(n970),.clk(gclk));
	jand g0329(.dina(n970),.dinb(n952),.dout(n971),.clk(gclk));
	jnot g0330(.din(w_n971_0[1]),.dout(n972),.clk(gclk));
	jnot g0331(.din(w_in030_0[1]),.dout(n973),.clk(gclk));
	jand g0332(.dina(w_in130_0[1]),.dinb(w_n973_0[1]),.dout(n974),.clk(gclk));
	jnot g0333(.din(w_in129_0[1]),.dout(n975),.clk(gclk));
	jand g0334(.dina(w_n975_0[1]),.dinb(w_in029_0[1]),.dout(n976),.clk(gclk));
	jnot g0335(.din(w_n976_0[1]),.dout(n977),.clk(gclk));
	jnot g0336(.din(w_in029_0[0]),.dout(n978),.clk(gclk));
	jand g0337(.dina(w_in129_0[0]),.dinb(w_n978_0[1]),.dout(n979),.clk(gclk));
	jnot g0338(.din(w_in128_0[1]),.dout(n980),.clk(gclk));
	jand g0339(.dina(w_n980_0[1]),.dinb(w_in028_0[1]),.dout(n981),.clk(gclk));
	jnot g0340(.din(w_n981_0[1]),.dout(n982),.clk(gclk));
	jnot g0341(.din(w_in028_0[0]),.dout(n983),.clk(gclk));
	jand g0342(.dina(w_in128_0[0]),.dinb(w_n983_0[1]),.dout(n984),.clk(gclk));
	jnot g0343(.din(w_in127_0[1]),.dout(n985),.clk(gclk));
	jand g0344(.dina(w_n985_0[1]),.dinb(w_in027_0[1]),.dout(n986),.clk(gclk));
	jnot g0345(.din(w_n986_0[1]),.dout(n987),.clk(gclk));
	jnot g0346(.din(w_in027_0[0]),.dout(n988),.clk(gclk));
	jand g0347(.dina(w_in127_0[0]),.dinb(w_n988_0[1]),.dout(n989),.clk(gclk));
	jnot g0348(.din(w_in126_0[1]),.dout(n990),.clk(gclk));
	jand g0349(.dina(w_n990_0[1]),.dinb(w_in026_0[1]),.dout(n991),.clk(gclk));
	jnot g0350(.din(w_n991_0[1]),.dout(n992),.clk(gclk));
	jnot g0351(.din(w_in023_0[1]),.dout(n993),.clk(gclk));
	jand g0352(.dina(w_in123_0[1]),.dinb(w_n993_0[1]),.dout(n994),.clk(gclk));
	jnot g0353(.din(w_in022_0[1]),.dout(n995),.clk(gclk));
	jand g0354(.dina(w_in122_0[1]),.dinb(w_n995_0[1]),.dout(n996),.clk(gclk));
	jnot g0355(.din(w_in121_0[1]),.dout(n997),.clk(gclk));
	jand g0356(.dina(w_n997_0[1]),.dinb(w_in021_0[1]),.dout(n998),.clk(gclk));
	jnot g0357(.din(w_n998_0[1]),.dout(n999),.clk(gclk));
	jnot g0358(.din(w_in021_0[0]),.dout(n1000),.clk(gclk));
	jand g0359(.dina(w_in121_0[0]),.dinb(w_n1000_0[1]),.dout(n1001),.clk(gclk));
	jnot g0360(.din(w_in120_0[1]),.dout(n1002),.clk(gclk));
	jand g0361(.dina(w_n1002_0[1]),.dinb(w_in020_0[1]),.dout(n1003),.clk(gclk));
	jnot g0362(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jnot g0363(.din(w_in020_0[0]),.dout(n1005),.clk(gclk));
	jand g0364(.dina(w_in120_0[0]),.dinb(w_n1005_0[1]),.dout(n1006),.clk(gclk));
	jnot g0365(.din(w_in119_0[1]),.dout(n1007),.clk(gclk));
	jand g0366(.dina(w_n1007_0[1]),.dinb(w_in019_0[1]),.dout(n1008),.clk(gclk));
	jnot g0367(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jnot g0368(.din(w_in019_0[0]),.dout(n1010),.clk(gclk));
	jand g0369(.dina(w_in119_0[0]),.dinb(w_n1010_0[1]),.dout(n1011),.clk(gclk));
	jnot g0370(.din(w_in118_0[1]),.dout(n1012),.clk(gclk));
	jand g0371(.dina(w_n1012_0[1]),.dinb(w_in018_0[1]),.dout(n1013),.clk(gclk));
	jnot g0372(.din(w_n1013_0[1]),.dout(n1014),.clk(gclk));
	jnot g0373(.din(w_in015_0[1]),.dout(n1015),.clk(gclk));
	jand g0374(.dina(w_in115_0[1]),.dinb(w_n1015_0[1]),.dout(n1016),.clk(gclk));
	jnot g0375(.din(w_in014_0[1]),.dout(n1017),.clk(gclk));
	jand g0376(.dina(w_in114_0[1]),.dinb(w_n1017_0[1]),.dout(n1018),.clk(gclk));
	jnot g0377(.din(w_in113_0[1]),.dout(n1019),.clk(gclk));
	jand g0378(.dina(w_n1019_0[1]),.dinb(w_in013_0[1]),.dout(n1020),.clk(gclk));
	jnot g0379(.din(w_n1020_0[1]),.dout(n1021),.clk(gclk));
	jnot g0380(.din(w_in013_0[0]),.dout(n1022),.clk(gclk));
	jand g0381(.dina(w_in113_0[0]),.dinb(w_n1022_0[1]),.dout(n1023),.clk(gclk));
	jnot g0382(.din(w_in112_0[1]),.dout(n1024),.clk(gclk));
	jand g0383(.dina(w_n1024_0[1]),.dinb(w_in012_0[1]),.dout(n1025),.clk(gclk));
	jnot g0384(.din(w_n1025_0[1]),.dout(n1026),.clk(gclk));
	jnot g0385(.din(w_in012_0[0]),.dout(n1027),.clk(gclk));
	jand g0386(.dina(w_in112_0[0]),.dinb(w_n1027_0[1]),.dout(n1028),.clk(gclk));
	jnot g0387(.din(w_in111_0[1]),.dout(n1029),.clk(gclk));
	jand g0388(.dina(w_n1029_0[1]),.dinb(w_in011_0[1]),.dout(n1030),.clk(gclk));
	jnot g0389(.din(w_n1030_0[1]),.dout(n1031),.clk(gclk));
	jnot g0390(.din(w_in011_0[0]),.dout(n1032),.clk(gclk));
	jand g0391(.dina(w_in111_0[0]),.dinb(w_n1032_0[1]),.dout(n1033),.clk(gclk));
	jnot g0392(.din(w_in110_0[1]),.dout(n1034),.clk(gclk));
	jand g0393(.dina(w_n1034_0[1]),.dinb(w_in010_0[1]),.dout(n1035),.clk(gclk));
	jnot g0394(.din(w_n1035_0[1]),.dout(n1036),.clk(gclk));
	jnot g0395(.din(w_in07_0[1]),.dout(n1037),.clk(gclk));
	jand g0396(.dina(w_in17_0[1]),.dinb(w_n1037_0[1]),.dout(n1038),.clk(gclk));
	jnot g0397(.din(w_in03_0[2]),.dout(n1039),.clk(gclk));
	jand g0398(.dina(w_in13_0[2]),.dinb(w_n1039_0[1]),.dout(n1040),.clk(gclk));
	jnot g0399(.din(w_in12_0[2]),.dout(n1041),.clk(gclk));
	jand g0400(.dina(w_n1041_0[2]),.dinb(w_in02_1[1]),.dout(n1042),.clk(gclk));
	jnot g0401(.din(w_n1042_0[1]),.dout(n1043),.clk(gclk));
	jnot g0402(.din(w_in01_1[1]),.dout(n1044),.clk(gclk));
	jor g0403(.dina(w_in11_1[1]),.dinb(w_n1044_0[2]),.dout(n1045),.clk(gclk));
	jnot g0404(.din(w_in00_0[2]),.dout(n1046),.clk(gclk));
	jor g0405(.dina(w_in10_0[2]),.dinb(w_n1046_0[1]),.dout(n1047),.clk(gclk));
	jand g0406(.dina(n1047),.dinb(n1045),.dout(n1048),.clk(gclk));
	jnot g0407(.din(w_in02_1[0]),.dout(n1049),.clk(gclk));
	jand g0408(.dina(w_in12_0[1]),.dinb(w_n1049_0[1]),.dout(n1050),.clk(gclk));
	jand g0409(.dina(w_in11_1[0]),.dinb(w_n1044_0[1]),.dout(n1051),.clk(gclk));
	jor g0410(.dina(n1051),.dinb(n1050),.dout(n1052),.clk(gclk));
	jor g0411(.dina(n1052),.dinb(n1048),.dout(n1053),.clk(gclk));
	jnot g0412(.din(w_in13_0[1]),.dout(n1054),.clk(gclk));
	jand g0413(.dina(w_n1054_0[1]),.dinb(w_in03_0[1]),.dout(n1055),.clk(gclk));
	jnot g0414(.din(w_n1055_0[1]),.dout(n1056),.clk(gclk));
	jand g0415(.dina(n1056),.dinb(n1053),.dout(n1057),.clk(gclk));
	jand g0416(.dina(n1057),.dinb(n1043),.dout(n1058),.clk(gclk));
	jnot g0417(.din(w_in04_0[1]),.dout(n1059),.clk(gclk));
	jand g0418(.dina(w_in14_0[1]),.dinb(w_n1059_0[1]),.dout(n1060),.clk(gclk));
	jor g0419(.dina(w_n1060_0[1]),.dinb(n1058),.dout(n1061),.clk(gclk));
	jor g0420(.dina(n1061),.dinb(w_n1040_0[1]),.dout(n1062),.clk(gclk));
	jnot g0421(.din(w_in14_0[0]),.dout(n1063),.clk(gclk));
	jand g0422(.dina(w_n1063_0[1]),.dinb(w_in04_0[0]),.dout(n1064),.clk(gclk));
	jnot g0423(.din(w_in15_0[1]),.dout(n1065),.clk(gclk));
	jand g0424(.dina(w_n1065_0[1]),.dinb(w_in05_0[1]),.dout(n1066),.clk(gclk));
	jor g0425(.dina(n1066),.dinb(n1064),.dout(n1067),.clk(gclk));
	jnot g0426(.din(w_n1067_0[1]),.dout(n1068),.clk(gclk));
	jand g0427(.dina(n1068),.dinb(n1062),.dout(n1069),.clk(gclk));
	jnot g0428(.din(w_in06_0[1]),.dout(n1070),.clk(gclk));
	jand g0429(.dina(w_in16_0[1]),.dinb(w_n1070_0[1]),.dout(n1071),.clk(gclk));
	jnot g0430(.din(w_in05_0[0]),.dout(n1072),.clk(gclk));
	jand g0431(.dina(w_in15_0[0]),.dinb(w_n1072_0[1]),.dout(n1073),.clk(gclk));
	jor g0432(.dina(n1073),.dinb(n1071),.dout(n1074),.clk(gclk));
	jor g0433(.dina(w_n1074_0[1]),.dinb(n1069),.dout(n1075),.clk(gclk));
	jnot g0434(.din(w_in17_0[0]),.dout(n1076),.clk(gclk));
	jand g0435(.dina(w_n1076_0[1]),.dinb(w_in07_0[0]),.dout(n1077),.clk(gclk));
	jnot g0436(.din(w_in16_0[0]),.dout(n1078),.clk(gclk));
	jand g0437(.dina(w_n1078_0[1]),.dinb(w_in06_0[0]),.dout(n1079),.clk(gclk));
	jor g0438(.dina(n1079),.dinb(n1077),.dout(n1080),.clk(gclk));
	jnot g0439(.din(w_n1080_0[1]),.dout(n1081),.clk(gclk));
	jand g0440(.dina(n1081),.dinb(n1075),.dout(n1082),.clk(gclk));
	jnot g0441(.din(w_in08_0[1]),.dout(n1083),.clk(gclk));
	jand g0442(.dina(w_in18_0[1]),.dinb(w_n1083_0[1]),.dout(n1084),.clk(gclk));
	jor g0443(.dina(w_n1084_0[1]),.dinb(n1082),.dout(n1085),.clk(gclk));
	jor g0444(.dina(n1085),.dinb(w_n1038_0[1]),.dout(n1086),.clk(gclk));
	jnot g0445(.din(w_in18_0[0]),.dout(n1087),.clk(gclk));
	jand g0446(.dina(w_n1087_0[1]),.dinb(w_in08_0[0]),.dout(n1088),.clk(gclk));
	jnot g0447(.din(w_in19_0[1]),.dout(n1089),.clk(gclk));
	jand g0448(.dina(w_n1089_0[1]),.dinb(w_in09_0[1]),.dout(n1090),.clk(gclk));
	jor g0449(.dina(n1090),.dinb(n1088),.dout(n1091),.clk(gclk));
	jnot g0450(.din(w_n1091_0[1]),.dout(n1092),.clk(gclk));
	jand g0451(.dina(n1092),.dinb(n1086),.dout(n1093),.clk(gclk));
	jnot g0452(.din(w_in010_0[0]),.dout(n1094),.clk(gclk));
	jand g0453(.dina(w_in110_0[0]),.dinb(w_n1094_0[1]),.dout(n1095),.clk(gclk));
	jnot g0454(.din(w_in09_0[0]),.dout(n1096),.clk(gclk));
	jand g0455(.dina(w_in19_0[0]),.dinb(w_n1096_0[1]),.dout(n1097),.clk(gclk));
	jor g0456(.dina(n1097),.dinb(n1095),.dout(n1098),.clk(gclk));
	jor g0457(.dina(w_n1098_0[1]),.dinb(n1093),.dout(n1099),.clk(gclk));
	jand g0458(.dina(n1099),.dinb(n1036),.dout(n1100),.clk(gclk));
	jor g0459(.dina(n1100),.dinb(w_n1033_0[1]),.dout(n1101),.clk(gclk));
	jand g0460(.dina(n1101),.dinb(n1031),.dout(n1102),.clk(gclk));
	jor g0461(.dina(n1102),.dinb(w_n1028_0[1]),.dout(n1103),.clk(gclk));
	jand g0462(.dina(n1103),.dinb(n1026),.dout(n1104),.clk(gclk));
	jor g0463(.dina(n1104),.dinb(w_n1023_0[1]),.dout(n1105),.clk(gclk));
	jand g0464(.dina(n1105),.dinb(n1021),.dout(n1106),.clk(gclk));
	jor g0465(.dina(n1106),.dinb(w_n1018_0[1]),.dout(n1107),.clk(gclk));
	jnot g0466(.din(w_in115_0[0]),.dout(n1108),.clk(gclk));
	jand g0467(.dina(w_n1108_0[1]),.dinb(w_in015_0[0]),.dout(n1109),.clk(gclk));
	jnot g0468(.din(w_in114_0[0]),.dout(n1110),.clk(gclk));
	jand g0469(.dina(w_n1110_0[1]),.dinb(w_in014_0[0]),.dout(n1111),.clk(gclk));
	jor g0470(.dina(n1111),.dinb(n1109),.dout(n1112),.clk(gclk));
	jnot g0471(.din(w_n1112_0[1]),.dout(n1113),.clk(gclk));
	jand g0472(.dina(n1113),.dinb(n1107),.dout(n1114),.clk(gclk));
	jnot g0473(.din(w_in016_0[1]),.dout(n1115),.clk(gclk));
	jand g0474(.dina(w_in116_0[1]),.dinb(w_n1115_0[1]),.dout(n1116),.clk(gclk));
	jor g0475(.dina(w_n1116_0[1]),.dinb(n1114),.dout(n1117),.clk(gclk));
	jor g0476(.dina(n1117),.dinb(w_n1016_0[1]),.dout(n1118),.clk(gclk));
	jnot g0477(.din(w_in116_0[0]),.dout(n1119),.clk(gclk));
	jand g0478(.dina(w_n1119_0[1]),.dinb(w_in016_0[0]),.dout(n1120),.clk(gclk));
	jnot g0479(.din(w_in117_0[1]),.dout(n1121),.clk(gclk));
	jand g0480(.dina(w_n1121_0[1]),.dinb(w_in017_0[1]),.dout(n1122),.clk(gclk));
	jor g0481(.dina(n1122),.dinb(n1120),.dout(n1123),.clk(gclk));
	jnot g0482(.din(w_n1123_0[1]),.dout(n1124),.clk(gclk));
	jand g0483(.dina(n1124),.dinb(n1118),.dout(n1125),.clk(gclk));
	jnot g0484(.din(w_in018_0[0]),.dout(n1126),.clk(gclk));
	jand g0485(.dina(w_in118_0[0]),.dinb(w_n1126_0[1]),.dout(n1127),.clk(gclk));
	jnot g0486(.din(w_in017_0[0]),.dout(n1128),.clk(gclk));
	jand g0487(.dina(w_in117_0[0]),.dinb(w_n1128_0[1]),.dout(n1129),.clk(gclk));
	jor g0488(.dina(n1129),.dinb(n1127),.dout(n1130),.clk(gclk));
	jor g0489(.dina(w_n1130_0[1]),.dinb(n1125),.dout(n1131),.clk(gclk));
	jand g0490(.dina(n1131),.dinb(n1014),.dout(n1132),.clk(gclk));
	jor g0491(.dina(n1132),.dinb(w_n1011_0[1]),.dout(n1133),.clk(gclk));
	jand g0492(.dina(n1133),.dinb(n1009),.dout(n1134),.clk(gclk));
	jor g0493(.dina(n1134),.dinb(w_n1006_0[1]),.dout(n1135),.clk(gclk));
	jand g0494(.dina(n1135),.dinb(n1004),.dout(n1136),.clk(gclk));
	jor g0495(.dina(n1136),.dinb(w_n1001_0[1]),.dout(n1137),.clk(gclk));
	jand g0496(.dina(n1137),.dinb(n999),.dout(n1138),.clk(gclk));
	jor g0497(.dina(n1138),.dinb(w_n996_0[1]),.dout(n1139),.clk(gclk));
	jnot g0498(.din(w_in123_0[0]),.dout(n1140),.clk(gclk));
	jand g0499(.dina(w_n1140_0[1]),.dinb(w_in023_0[0]),.dout(n1141),.clk(gclk));
	jnot g0500(.din(w_in122_0[0]),.dout(n1142),.clk(gclk));
	jand g0501(.dina(w_n1142_0[1]),.dinb(w_in022_0[0]),.dout(n1143),.clk(gclk));
	jor g0502(.dina(n1143),.dinb(n1141),.dout(n1144),.clk(gclk));
	jnot g0503(.din(w_n1144_0[1]),.dout(n1145),.clk(gclk));
	jand g0504(.dina(n1145),.dinb(n1139),.dout(n1146),.clk(gclk));
	jnot g0505(.din(w_in024_0[1]),.dout(n1147),.clk(gclk));
	jand g0506(.dina(w_in124_0[1]),.dinb(w_n1147_0[1]),.dout(n1148),.clk(gclk));
	jor g0507(.dina(w_n1148_0[1]),.dinb(n1146),.dout(n1149),.clk(gclk));
	jor g0508(.dina(n1149),.dinb(w_n994_0[1]),.dout(n1150),.clk(gclk));
	jnot g0509(.din(w_in124_0[0]),.dout(n1151),.clk(gclk));
	jand g0510(.dina(w_n1151_0[1]),.dinb(w_in024_0[0]),.dout(n1152),.clk(gclk));
	jnot g0511(.din(w_in125_0[1]),.dout(n1153),.clk(gclk));
	jand g0512(.dina(w_n1153_0[1]),.dinb(w_in025_0[1]),.dout(n1154),.clk(gclk));
	jor g0513(.dina(n1154),.dinb(n1152),.dout(n1155),.clk(gclk));
	jnot g0514(.din(w_n1155_0[1]),.dout(n1156),.clk(gclk));
	jand g0515(.dina(n1156),.dinb(n1150),.dout(n1157),.clk(gclk));
	jnot g0516(.din(w_in026_0[0]),.dout(n1158),.clk(gclk));
	jand g0517(.dina(w_in126_0[0]),.dinb(w_n1158_0[1]),.dout(n1159),.clk(gclk));
	jnot g0518(.din(w_in025_0[0]),.dout(n1160),.clk(gclk));
	jand g0519(.dina(w_in125_0[0]),.dinb(w_n1160_0[1]),.dout(n1161),.clk(gclk));
	jor g0520(.dina(n1161),.dinb(n1159),.dout(n1162),.clk(gclk));
	jor g0521(.dina(w_n1162_0[1]),.dinb(n1157),.dout(n1163),.clk(gclk));
	jand g0522(.dina(n1163),.dinb(n992),.dout(n1164),.clk(gclk));
	jor g0523(.dina(n1164),.dinb(w_n989_0[1]),.dout(n1165),.clk(gclk));
	jand g0524(.dina(n1165),.dinb(n987),.dout(n1166),.clk(gclk));
	jor g0525(.dina(n1166),.dinb(w_n984_0[1]),.dout(n1167),.clk(gclk));
	jand g0526(.dina(n1167),.dinb(n982),.dout(n1168),.clk(gclk));
	jor g0527(.dina(n1168),.dinb(w_n979_0[1]),.dout(n1169),.clk(gclk));
	jand g0528(.dina(n1169),.dinb(n977),.dout(n1170),.clk(gclk));
	jor g0529(.dina(n1170),.dinb(w_n974_0[1]),.dout(n1171),.clk(gclk));
	jnot g0530(.din(w_in131_0[1]),.dout(n1172),.clk(gclk));
	jand g0531(.dina(w_n1172_0[1]),.dinb(w_in031_0[1]),.dout(n1173),.clk(gclk));
	jnot g0532(.din(w_in130_0[0]),.dout(n1174),.clk(gclk));
	jand g0533(.dina(w_n1174_0[1]),.dinb(w_in030_0[0]),.dout(n1175),.clk(gclk));
	jor g0534(.dina(n1175),.dinb(n1173),.dout(n1176),.clk(gclk));
	jnot g0535(.din(w_n1176_0[1]),.dout(n1177),.clk(gclk));
	jand g0536(.dina(n1177),.dinb(n1171),.dout(n1178),.clk(gclk));
	jnot g0537(.din(w_in031_0[0]),.dout(n1179),.clk(gclk));
	jand g0538(.dina(w_in131_0[0]),.dinb(w_n1179_0[1]),.dout(n1180),.clk(gclk));
	jnot g0539(.din(w_in032_0[0]),.dout(n1181),.clk(gclk));
	jand g0540(.dina(w_in132_0[0]),.dinb(w_n1181_0[1]),.dout(n1182),.clk(gclk));
	jor g0541(.dina(n1182),.dinb(n1180),.dout(n1183),.clk(gclk));
	jor g0542(.dina(n1183),.dinb(w_n947_0[0]),.dout(n1184),.clk(gclk));
	jor g0543(.dina(n1184),.dinb(w_n969_0[0]),.dout(n1185),.clk(gclk));
	jor g0544(.dina(w_n1185_0[1]),.dinb(n1178),.dout(n1186),.clk(gclk));
	jnot g0545(.din(w_n967_0[0]),.dout(n1187),.clk(gclk));
	jnot g0546(.din(w_in137_0[0]),.dout(n1188),.clk(gclk));
	jand g0547(.dina(w_n1188_0[1]),.dinb(w_in037_0[0]),.dout(n1189),.clk(gclk));
	jnot g0548(.din(w_in136_0[0]),.dout(n1190),.clk(gclk));
	jand g0549(.dina(w_n1190_0[1]),.dinb(w_in036_0[0]),.dout(n1191),.clk(gclk));
	jor g0550(.dina(n1191),.dinb(n1189),.dout(n1192),.clk(gclk));
	jand g0551(.dina(n1192),.dinb(n1187),.dout(n1193),.clk(gclk));
	jnot g0552(.din(w_n968_0[0]),.dout(n1194),.clk(gclk));
	jnot g0553(.din(w_in135_0[0]),.dout(n1195),.clk(gclk));
	jand g0554(.dina(w_n1195_0[1]),.dinb(w_in035_0[0]),.dout(n1196),.clk(gclk));
	jand g0555(.dina(n1196),.dinb(n1194),.dout(n1197),.clk(gclk));
	jnot g0556(.din(w_in139_0[0]),.dout(n1198),.clk(gclk));
	jand g0557(.dina(w_n1198_0[1]),.dinb(w_in039_0[0]),.dout(n1199),.clk(gclk));
	jnot g0558(.din(w_n963_0[0]),.dout(n1200),.clk(gclk));
	jnot g0559(.din(w_in138_0[0]),.dout(n1201),.clk(gclk));
	jand g0560(.dina(w_n1201_0[1]),.dinb(w_in038_0[0]),.dout(n1202),.clk(gclk));
	jand g0561(.dina(n1202),.dinb(n1200),.dout(n1203),.clk(gclk));
	jor g0562(.dina(n1203),.dinb(n1199),.dout(n1204),.clk(gclk));
	jor g0563(.dina(n1204),.dinb(n1197),.dout(n1205),.clk(gclk));
	jor g0564(.dina(n1205),.dinb(n1193),.dout(n1206),.clk(gclk));
	jnot g0565(.din(w_n1206_0[1]),.dout(n1207),.clk(gclk));
	jand g0566(.dina(n1207),.dinb(n1186),.dout(n1208),.clk(gclk));
	jand g0567(.dina(n1208),.dinb(n972),.dout(n1209),.clk(gclk));
	jnot g0568(.din(w_in040_0[0]),.dout(n1210),.clk(gclk));
	jand g0569(.dina(w_in140_0[0]),.dinb(w_n1210_0[1]),.dout(n1211),.clk(gclk));
	jor g0570(.dina(n1211),.dinb(w_n925_0[0]),.dout(n1212),.clk(gclk));
	jor g0571(.dina(n1212),.dinb(w_n932_0[0]),.dout(n1213),.clk(gclk));
	jor g0572(.dina(w_n1213_0[1]),.dinb(n1209),.dout(n1214),.clk(gclk));
	jnot g0573(.din(w_n918_0[0]),.dout(n1215),.clk(gclk));
	jnot g0574(.din(w_in145_0[0]),.dout(n1216),.clk(gclk));
	jand g0575(.dina(w_n1216_0[1]),.dinb(w_in045_0[0]),.dout(n1217),.clk(gclk));
	jnot g0576(.din(w_in144_0[0]),.dout(n1218),.clk(gclk));
	jand g0577(.dina(w_n1218_0[1]),.dinb(w_in044_0[0]),.dout(n1219),.clk(gclk));
	jor g0578(.dina(n1219),.dinb(n1217),.dout(n1220),.clk(gclk));
	jand g0579(.dina(n1220),.dinb(n1215),.dout(n1221),.clk(gclk));
	jnot g0580(.din(w_n912_0[0]),.dout(n1222),.clk(gclk));
	jnot g0581(.din(w_in147_0[0]),.dout(n1223),.clk(gclk));
	jand g0582(.dina(w_n1223_0[1]),.dinb(w_in047_0[0]),.dout(n1224),.clk(gclk));
	jnot g0583(.din(w_in146_0[0]),.dout(n1225),.clk(gclk));
	jand g0584(.dina(w_n1225_0[1]),.dinb(w_in046_0[0]),.dout(n1226),.clk(gclk));
	jor g0585(.dina(n1226),.dinb(n1224),.dout(n1227),.clk(gclk));
	jand g0586(.dina(n1227),.dinb(n1222),.dout(n1228),.clk(gclk));
	jor g0587(.dina(n1228),.dinb(n1221),.dout(n1229),.clk(gclk));
	jnot g0588(.din(n1229),.dout(n1230),.clk(gclk));
	jor g0589(.dina(w_n919_0[0]),.dinb(w_in143_0[1]),.dout(n1231),.clk(gclk));
	jor g0590(.dina(n1231),.dinb(w_n922_0[1]),.dout(n1232),.clk(gclk));
	jand g0591(.dina(n1232),.dinb(n1230),.dout(n1233),.clk(gclk));
	jand g0592(.dina(w_n1233_0[1]),.dinb(n1214),.dout(n1234),.clk(gclk));
	jand g0593(.dina(n1234),.dinb(n940),.dout(n1235),.clk(gclk));
	jnot g0594(.din(w_in048_0[1]),.dout(n1236),.clk(gclk));
	jand g0595(.dina(w_in148_0[1]),.dinb(w_n1236_0[1]),.dout(n1237),.clk(gclk));
	jnot g0596(.din(n1237),.dout(n1238),.clk(gclk));
	jnot g0597(.din(w_in049_0[1]),.dout(n1239),.clk(gclk));
	jand g0598(.dina(w_in149_0[1]),.dinb(w_n1239_0[1]),.dout(n1240),.clk(gclk));
	jnot g0599(.din(n1240),.dout(n1241),.clk(gclk));
	jnot g0600(.din(w_in050_0[1]),.dout(n1242),.clk(gclk));
	jand g0601(.dina(w_in150_0[1]),.dinb(w_n1242_0[1]),.dout(n1243),.clk(gclk));
	jnot g0602(.din(w_in051_0[0]),.dout(n1244),.clk(gclk));
	jand g0603(.dina(w_in151_0[0]),.dinb(w_n1244_0[1]),.dout(n1245),.clk(gclk));
	jor g0604(.dina(n1245),.dinb(n1243),.dout(n1246),.clk(gclk));
	jor g0605(.dina(n1246),.dinb(w_n904_0[0]),.dout(n1247),.clk(gclk));
	jnot g0606(.din(n1247),.dout(n1248),.clk(gclk));
	jand g0607(.dina(w_n1248_0[1]),.dinb(w_n1241_0[1]),.dout(n1249),.clk(gclk));
	jand g0608(.dina(n1249),.dinb(n1238),.dout(n1250),.clk(gclk));
	jnot g0609(.din(w_n1250_0[1]),.dout(n1251),.clk(gclk));
	jor g0610(.dina(n1251),.dinb(n1235),.dout(n1252),.clk(gclk));
	jnot g0611(.din(w_in149_0[0]),.dout(n1253),.clk(gclk));
	jand g0612(.dina(w_n1253_0[1]),.dinb(w_in049_0[0]),.dout(n1254),.clk(gclk));
	jnot g0613(.din(w_in150_0[0]),.dout(n1255),.clk(gclk));
	jand g0614(.dina(w_n1255_0[1]),.dinb(w_in050_0[0]),.dout(n1256),.clk(gclk));
	jor g0615(.dina(n1256),.dinb(n1254),.dout(n1257),.clk(gclk));
	jnot g0616(.din(w_in148_0[0]),.dout(n1258),.clk(gclk));
	jand g0617(.dina(w_n1258_0[1]),.dinb(w_in048_0[0]),.dout(n1259),.clk(gclk));
	jand g0618(.dina(n1259),.dinb(w_n1241_0[0]),.dout(n1260),.clk(gclk));
	jor g0619(.dina(n1260),.dinb(n1257),.dout(n1261),.clk(gclk));
	jand g0620(.dina(n1261),.dinb(w_n1248_0[0]),.dout(n1262),.clk(gclk));
	jnot g0621(.din(w_in155_0[0]),.dout(n1263),.clk(gclk));
	jand g0622(.dina(w_n1263_0[1]),.dinb(w_in055_0[0]),.dout(n1264),.clk(gclk));
	jnot g0623(.din(w_n900_0[0]),.dout(n1265),.clk(gclk));
	jnot g0624(.din(w_n895_0[0]),.dout(n1266),.clk(gclk));
	jnot g0625(.din(w_in152_0[0]),.dout(n1267),.clk(gclk));
	jand g0626(.dina(w_n1267_0[1]),.dinb(w_in052_0[0]),.dout(n1268),.clk(gclk));
	jand g0627(.dina(n1268),.dinb(n1266),.dout(n1269),.clk(gclk));
	jnot g0628(.din(w_in154_0[0]),.dout(n1270),.clk(gclk));
	jand g0629(.dina(w_n1270_0[1]),.dinb(w_in054_0[0]),.dout(n1271),.clk(gclk));
	jnot g0630(.din(w_in153_0[0]),.dout(n1272),.clk(gclk));
	jand g0631(.dina(w_n1272_0[1]),.dinb(w_in053_0[0]),.dout(n1273),.clk(gclk));
	jor g0632(.dina(n1273),.dinb(n1271),.dout(n1274),.clk(gclk));
	jor g0633(.dina(n1274),.dinb(n1269),.dout(n1275),.clk(gclk));
	jand g0634(.dina(n1275),.dinb(n1265),.dout(n1276),.clk(gclk));
	jor g0635(.dina(n1276),.dinb(n1264),.dout(n1277),.clk(gclk));
	jor g0636(.dina(n1277),.dinb(n1262),.dout(n1278),.clk(gclk));
	jnot g0637(.din(w_n1278_0[1]),.dout(n1279),.clk(gclk));
	jand g0638(.dina(n1279),.dinb(n1252),.dout(n1280),.clk(gclk));
	jand g0639(.dina(n1280),.dinb(n908),.dout(n1281),.clk(gclk));
	jnot g0640(.din(w_in056_0[1]),.dout(n1282),.clk(gclk));
	jand g0641(.dina(w_in156_0[1]),.dinb(w_n1282_0[1]),.dout(n1283),.clk(gclk));
	jnot g0642(.din(n1283),.dout(n1284),.clk(gclk));
	jnot g0643(.din(w_in057_0[1]),.dout(n1285),.clk(gclk));
	jand g0644(.dina(w_in157_0[1]),.dinb(w_n1285_0[1]),.dout(n1286),.clk(gclk));
	jnot g0645(.din(n1286),.dout(n1287),.clk(gclk));
	jnot g0646(.din(w_in058_0[1]),.dout(n1288),.clk(gclk));
	jand g0647(.dina(w_in158_0[1]),.dinb(w_n1288_0[1]),.dout(n1289),.clk(gclk));
	jnot g0648(.din(w_in059_0[0]),.dout(n1290),.clk(gclk));
	jand g0649(.dina(w_in159_0[0]),.dinb(w_n1290_0[1]),.dout(n1291),.clk(gclk));
	jor g0650(.dina(n1291),.dinb(n1289),.dout(n1292),.clk(gclk));
	jor g0651(.dina(n1292),.dinb(w_n888_0[0]),.dout(n1293),.clk(gclk));
	jnot g0652(.din(n1293),.dout(n1294),.clk(gclk));
	jand g0653(.dina(w_n1294_0[1]),.dinb(w_n1287_0[1]),.dout(n1295),.clk(gclk));
	jand g0654(.dina(n1295),.dinb(n1284),.dout(n1296),.clk(gclk));
	jnot g0655(.din(w_n1296_0[1]),.dout(n1297),.clk(gclk));
	jor g0656(.dina(n1297),.dinb(n1281),.dout(n1298),.clk(gclk));
	jnot g0657(.din(w_in157_0[0]),.dout(n1299),.clk(gclk));
	jand g0658(.dina(w_n1299_0[1]),.dinb(w_in057_0[0]),.dout(n1300),.clk(gclk));
	jnot g0659(.din(w_in158_0[0]),.dout(n1301),.clk(gclk));
	jand g0660(.dina(w_n1301_0[1]),.dinb(w_in058_0[0]),.dout(n1302),.clk(gclk));
	jor g0661(.dina(n1302),.dinb(n1300),.dout(n1303),.clk(gclk));
	jnot g0662(.din(w_in156_0[0]),.dout(n1304),.clk(gclk));
	jand g0663(.dina(w_n1304_0[1]),.dinb(w_in056_0[0]),.dout(n1305),.clk(gclk));
	jand g0664(.dina(n1305),.dinb(w_n1287_0[0]),.dout(n1306),.clk(gclk));
	jor g0665(.dina(n1306),.dinb(n1303),.dout(n1307),.clk(gclk));
	jand g0666(.dina(n1307),.dinb(w_n1294_0[0]),.dout(n1308),.clk(gclk));
	jnot g0667(.din(w_n887_0[0]),.dout(n1309),.clk(gclk));
	jnot g0668(.din(w_in161_0[0]),.dout(n1310),.clk(gclk));
	jand g0669(.dina(w_n1310_0[1]),.dinb(w_in061_0[0]),.dout(n1311),.clk(gclk));
	jnot g0670(.din(w_in160_0[0]),.dout(n1312),.clk(gclk));
	jand g0671(.dina(w_n1312_0[1]),.dinb(w_in060_0[0]),.dout(n1313),.clk(gclk));
	jor g0672(.dina(n1313),.dinb(n1311),.dout(n1314),.clk(gclk));
	jand g0673(.dina(n1314),.dinb(n1309),.dout(n1315),.clk(gclk));
	jnot g0674(.din(w_n881_0[0]),.dout(n1316),.clk(gclk));
	jnot g0675(.din(w_in163_0[0]),.dout(n1317),.clk(gclk));
	jand g0676(.dina(w_n1317_0[1]),.dinb(w_in063_0[0]),.dout(n1318),.clk(gclk));
	jnot g0677(.din(w_in162_0[0]),.dout(n1319),.clk(gclk));
	jand g0678(.dina(w_n1319_0[1]),.dinb(w_in062_0[0]),.dout(n1320),.clk(gclk));
	jor g0679(.dina(n1320),.dinb(n1318),.dout(n1321),.clk(gclk));
	jand g0680(.dina(n1321),.dinb(n1316),.dout(n1322),.clk(gclk));
	jor g0681(.dina(n1322),.dinb(n1315),.dout(n1323),.clk(gclk));
	jor g0682(.dina(n1323),.dinb(n1308),.dout(n1324),.clk(gclk));
	jnot g0683(.din(w_n1324_0[1]),.dout(n1325),.clk(gclk));
	jand g0684(.dina(n1325),.dinb(n1298),.dout(n1326),.clk(gclk));
	jand g0685(.dina(n1326),.dinb(n892),.dout(n1327),.clk(gclk));
	jnot g0686(.din(w_in064_0[0]),.dout(n1328),.clk(gclk));
	jand g0687(.dina(w_in164_0[0]),.dinb(w_n1328_0[1]),.dout(n1329),.clk(gclk));
	jor g0688(.dina(n1329),.dinb(w_n865_0[0]),.dout(n1330),.clk(gclk));
	jor g0689(.dina(w_n1330_0[1]),.dinb(n1327),.dout(n1331),.clk(gclk));
	jand g0690(.dina(n1331),.dinb(n876),.dout(n1332),.clk(gclk));
	jnot g0691(.din(w_in067_0[0]),.dout(n1333),.clk(gclk));
	jand g0692(.dina(w_in167_0[0]),.dinb(w_n1333_0[1]),.dout(n1334),.clk(gclk));
	jnot g0693(.din(w_in066_0[0]),.dout(n1335),.clk(gclk));
	jand g0694(.dina(w_in166_0[0]),.dinb(w_n1335_0[1]),.dout(n1336),.clk(gclk));
	jor g0695(.dina(n1336),.dinb(n1334),.dout(n1337),.clk(gclk));
	jor g0696(.dina(w_n1337_0[1]),.dinb(n1332),.dout(n1338),.clk(gclk));
	jand g0697(.dina(n1338),.dinb(n863),.dout(n1339),.clk(gclk));
	jnot g0698(.din(w_in068_0[0]),.dout(n1340),.clk(gclk));
	jand g0699(.dina(w_in168_0[0]),.dinb(w_n1340_0[1]),.dout(n1341),.clk(gclk));
	jor g0700(.dina(n1341),.dinb(w_n844_0[0]),.dout(n1342),.clk(gclk));
	jor g0701(.dina(w_n1342_0[1]),.dinb(n1339),.dout(n1343),.clk(gclk));
	jand g0702(.dina(n1343),.dinb(n860),.dout(n1344),.clk(gclk));
	jnot g0703(.din(w_in075_0[0]),.dout(n1345),.clk(gclk));
	jand g0704(.dina(w_in175_0[0]),.dinb(w_n1345_0[1]),.dout(n1346),.clk(gclk));
	jnot g0705(.din(w_in074_0[1]),.dout(n1347),.clk(gclk));
	jand g0706(.dina(w_in174_0[1]),.dinb(w_n1347_0[1]),.dout(n1348),.clk(gclk));
	jor g0707(.dina(n1348),.dinb(n1346),.dout(n1349),.clk(gclk));
	jor g0708(.dina(w_n1349_0[1]),.dinb(n1344),.dout(n1350),.clk(gclk));
	jor g0709(.dina(n1350),.dinb(w_n836_0[1]),.dout(n1351),.clk(gclk));
	jnot g0710(.din(w_n1349_0[0]),.dout(n1352),.clk(gclk));
	jnot g0711(.din(w_in173_0[0]),.dout(n1353),.clk(gclk));
	jand g0712(.dina(w_n1353_0[1]),.dinb(w_in073_0[0]),.dout(n1354),.clk(gclk));
	jnot g0713(.din(w_in174_0[0]),.dout(n1355),.clk(gclk));
	jand g0714(.dina(w_n1355_0[1]),.dinb(w_in074_0[0]),.dout(n1356),.clk(gclk));
	jor g0715(.dina(n1356),.dinb(n1354),.dout(n1357),.clk(gclk));
	jnot g0716(.din(w_n835_0[0]),.dout(n1358),.clk(gclk));
	jnot g0717(.din(w_in172_0[0]),.dout(n1359),.clk(gclk));
	jand g0718(.dina(w_n1359_0[1]),.dinb(w_in072_0[0]),.dout(n1360),.clk(gclk));
	jand g0719(.dina(n1360),.dinb(n1358),.dout(n1361),.clk(gclk));
	jor g0720(.dina(n1361),.dinb(n1357),.dout(n1362),.clk(gclk));
	jand g0721(.dina(n1362),.dinb(w_n1352_0[1]),.dout(n1363),.clk(gclk));
	jnot g0722(.din(w_n1363_0[1]),.dout(n1364),.clk(gclk));
	jand g0723(.dina(n1364),.dinb(n1351),.dout(n1365),.clk(gclk));
	jand g0724(.dina(n1365),.dinb(n831),.dout(n1366),.clk(gclk));
	jnot g0725(.din(w_in076_0[0]),.dout(n1367),.clk(gclk));
	jand g0726(.dina(w_in176_0[0]),.dinb(w_n1367_0[1]),.dout(n1368),.clk(gclk));
	jor g0727(.dina(n1368),.dinb(w_n812_0[0]),.dout(n1369),.clk(gclk));
	jor g0728(.dina(w_n1369_0[1]),.dinb(n1366),.dout(n1370),.clk(gclk));
	jand g0729(.dina(n1370),.dinb(n828),.dout(n1371),.clk(gclk));
	jnot g0730(.din(w_in083_0[0]),.dout(n1372),.clk(gclk));
	jand g0731(.dina(w_in183_0[0]),.dinb(w_n1372_0[1]),.dout(n1373),.clk(gclk));
	jnot g0732(.din(w_in082_0[1]),.dout(n1374),.clk(gclk));
	jand g0733(.dina(w_in182_0[1]),.dinb(w_n1374_0[1]),.dout(n1375),.clk(gclk));
	jor g0734(.dina(n1375),.dinb(n1373),.dout(n1376),.clk(gclk));
	jor g0735(.dina(w_n1376_0[1]),.dinb(n1371),.dout(n1377),.clk(gclk));
	jor g0736(.dina(n1377),.dinb(w_n804_0[1]),.dout(n1378),.clk(gclk));
	jnot g0737(.din(w_n1376_0[0]),.dout(n1379),.clk(gclk));
	jnot g0738(.din(w_in181_0[0]),.dout(n1380),.clk(gclk));
	jand g0739(.dina(w_n1380_0[1]),.dinb(w_in081_0[0]),.dout(n1381),.clk(gclk));
	jnot g0740(.din(w_in182_0[0]),.dout(n1382),.clk(gclk));
	jand g0741(.dina(w_n1382_0[1]),.dinb(w_in082_0[0]),.dout(n1383),.clk(gclk));
	jor g0742(.dina(n1383),.dinb(n1381),.dout(n1384),.clk(gclk));
	jnot g0743(.din(w_n801_0[0]),.dout(n1385),.clk(gclk));
	jnot g0744(.din(w_in180_0[0]),.dout(n1386),.clk(gclk));
	jand g0745(.dina(w_n1386_0[1]),.dinb(w_in080_0[0]),.dout(n1387),.clk(gclk));
	jand g0746(.dina(n1387),.dinb(n1385),.dout(n1388),.clk(gclk));
	jor g0747(.dina(n1388),.dinb(n1384),.dout(n1389),.clk(gclk));
	jand g0748(.dina(n1389),.dinb(w_n1379_0[1]),.dout(n1390),.clk(gclk));
	jnot g0749(.din(w_n1390_0[1]),.dout(n1391),.clk(gclk));
	jand g0750(.dina(n1391),.dinb(n1378),.dout(n1392),.clk(gclk));
	jand g0751(.dina(n1392),.dinb(n799),.dout(n1393),.clk(gclk));
	jnot g0752(.din(w_in084_0[0]),.dout(n1394),.clk(gclk));
	jand g0753(.dina(w_in184_0[0]),.dinb(w_n1394_0[1]),.dout(n1395),.clk(gclk));
	jor g0754(.dina(n1395),.dinb(w_n780_0[0]),.dout(n1396),.clk(gclk));
	jor g0755(.dina(w_n1396_0[1]),.dinb(n1393),.dout(n1397),.clk(gclk));
	jand g0756(.dina(n1397),.dinb(n796),.dout(n1398),.clk(gclk));
	jnot g0757(.din(w_in091_0[0]),.dout(n1399),.clk(gclk));
	jand g0758(.dina(w_in191_0[0]),.dinb(w_n1399_0[1]),.dout(n1400),.clk(gclk));
	jnot g0759(.din(w_in090_0[1]),.dout(n1401),.clk(gclk));
	jand g0760(.dina(w_in190_0[1]),.dinb(w_n1401_0[1]),.dout(n1402),.clk(gclk));
	jor g0761(.dina(n1402),.dinb(n1400),.dout(n1403),.clk(gclk));
	jnot g0762(.din(w_in088_0[1]),.dout(n1404),.clk(gclk));
	jand g0763(.dina(w_in188_0[1]),.dinb(w_n1404_0[1]),.dout(n1405),.clk(gclk));
	jnot g0764(.din(w_in089_0[1]),.dout(n1406),.clk(gclk));
	jand g0765(.dina(w_in189_0[1]),.dinb(w_n1406_0[1]),.dout(n1407),.clk(gclk));
	jor g0766(.dina(w_n1407_0[1]),.dinb(n1405),.dout(n1408),.clk(gclk));
	jor g0767(.dina(n1408),.dinb(w_n1403_0[1]),.dout(n1409),.clk(gclk));
	jor g0768(.dina(w_n1409_0[1]),.dinb(n1398),.dout(n1410),.clk(gclk));
	jnot g0769(.din(w_n1403_0[0]),.dout(n1411),.clk(gclk));
	jnot g0770(.din(w_in189_0[0]),.dout(n1412),.clk(gclk));
	jand g0771(.dina(w_n1412_0[1]),.dinb(w_in089_0[0]),.dout(n1413),.clk(gclk));
	jnot g0772(.din(w_in190_0[0]),.dout(n1414),.clk(gclk));
	jand g0773(.dina(w_n1414_0[1]),.dinb(w_in090_0[0]),.dout(n1415),.clk(gclk));
	jor g0774(.dina(n1415),.dinb(n1413),.dout(n1416),.clk(gclk));
	jnot g0775(.din(w_n1407_0[0]),.dout(n1417),.clk(gclk));
	jnot g0776(.din(w_in188_0[0]),.dout(n1418),.clk(gclk));
	jand g0777(.dina(w_n1418_0[1]),.dinb(w_in088_0[0]),.dout(n1419),.clk(gclk));
	jand g0778(.dina(n1419),.dinb(n1417),.dout(n1420),.clk(gclk));
	jor g0779(.dina(n1420),.dinb(n1416),.dout(n1421),.clk(gclk));
	jand g0780(.dina(n1421),.dinb(n1411),.dout(n1422),.clk(gclk));
	jnot g0781(.din(w_n1422_0[1]),.dout(n1423),.clk(gclk));
	jand g0782(.dina(n1423),.dinb(n1410),.dout(n1424),.clk(gclk));
	jand g0783(.dina(n1424),.dinb(n772),.dout(n1425),.clk(gclk));
	jnot g0784(.din(w_in092_0[0]),.dout(n1426),.clk(gclk));
	jand g0785(.dina(w_in192_0[0]),.dinb(w_n1426_0[1]),.dout(n1427),.clk(gclk));
	jor g0786(.dina(n1427),.dinb(w_n753_0[0]),.dout(n1428),.clk(gclk));
	jor g0787(.dina(w_n1428_0[1]),.dinb(n1425),.dout(n1429),.clk(gclk));
	jand g0788(.dina(n1429),.dinb(n769),.dout(n1430),.clk(gclk));
	jnot g0789(.din(w_in099_0[0]),.dout(n1431),.clk(gclk));
	jand g0790(.dina(w_in199_0[0]),.dinb(w_n1431_0[1]),.dout(n1432),.clk(gclk));
	jnot g0791(.din(w_in098_0[1]),.dout(n1433),.clk(gclk));
	jand g0792(.dina(w_in198_0[1]),.dinb(w_n1433_0[1]),.dout(n1434),.clk(gclk));
	jor g0793(.dina(n1434),.dinb(n1432),.dout(n1435),.clk(gclk));
	jor g0794(.dina(w_n1435_0[1]),.dinb(n1430),.dout(n1436),.clk(gclk));
	jor g0795(.dina(n1436),.dinb(w_n745_0[1]),.dout(n1437),.clk(gclk));
	jnot g0796(.din(w_n1435_0[0]),.dout(n1438),.clk(gclk));
	jnot g0797(.din(w_in197_0[0]),.dout(n1439),.clk(gclk));
	jand g0798(.dina(w_n1439_0[1]),.dinb(w_in097_0[0]),.dout(n1440),.clk(gclk));
	jnot g0799(.din(w_in198_0[0]),.dout(n1441),.clk(gclk));
	jand g0800(.dina(w_n1441_0[1]),.dinb(w_in098_0[0]),.dout(n1442),.clk(gclk));
	jor g0801(.dina(n1442),.dinb(n1440),.dout(n1443),.clk(gclk));
	jnot g0802(.din(w_n742_0[0]),.dout(n1444),.clk(gclk));
	jnot g0803(.din(w_in196_0[0]),.dout(n1445),.clk(gclk));
	jand g0804(.dina(w_n1445_0[1]),.dinb(w_in096_0[0]),.dout(n1446),.clk(gclk));
	jand g0805(.dina(n1446),.dinb(n1444),.dout(n1447),.clk(gclk));
	jor g0806(.dina(n1447),.dinb(n1443),.dout(n1448),.clk(gclk));
	jand g0807(.dina(n1448),.dinb(w_n1438_0[1]),.dout(n1449),.clk(gclk));
	jnot g0808(.din(w_n1449_0[1]),.dout(n1450),.clk(gclk));
	jand g0809(.dina(n1450),.dinb(n1437),.dout(n1451),.clk(gclk));
	jand g0810(.dina(n1451),.dinb(n740),.dout(n1452),.clk(gclk));
	jnot g0811(.din(w_in0100_0[0]),.dout(n1453),.clk(gclk));
	jand g0812(.dina(w_in1100_0[0]),.dinb(w_n1453_0[1]),.dout(n1454),.clk(gclk));
	jor g0813(.dina(n1454),.dinb(w_n721_0[0]),.dout(n1455),.clk(gclk));
	jor g0814(.dina(w_n1455_0[1]),.dinb(n1452),.dout(n1456),.clk(gclk));
	jand g0815(.dina(n1456),.dinb(n737),.dout(n1457),.clk(gclk));
	jnot g0816(.din(w_in0107_0[0]),.dout(n1458),.clk(gclk));
	jand g0817(.dina(w_in1107_0[0]),.dinb(w_n1458_0[1]),.dout(n1459),.clk(gclk));
	jnot g0818(.din(w_in0106_0[1]),.dout(n1460),.clk(gclk));
	jand g0819(.dina(w_in1106_0[1]),.dinb(w_n1460_0[1]),.dout(n1461),.clk(gclk));
	jor g0820(.dina(n1461),.dinb(n1459),.dout(n1462),.clk(gclk));
	jor g0821(.dina(w_n1462_0[1]),.dinb(n1457),.dout(n1463),.clk(gclk));
	jor g0822(.dina(n1463),.dinb(w_n713_0[1]),.dout(n1464),.clk(gclk));
	jnot g0823(.din(w_n1462_0[0]),.dout(n1465),.clk(gclk));
	jnot g0824(.din(w_in1105_0[0]),.dout(n1466),.clk(gclk));
	jand g0825(.dina(w_n1466_0[1]),.dinb(w_in0105_0[0]),.dout(n1467),.clk(gclk));
	jnot g0826(.din(w_in1106_0[0]),.dout(n1468),.clk(gclk));
	jand g0827(.dina(w_n1468_0[1]),.dinb(w_in0106_0[0]),.dout(n1469),.clk(gclk));
	jor g0828(.dina(n1469),.dinb(n1467),.dout(n1470),.clk(gclk));
	jnot g0829(.din(w_n712_0[0]),.dout(n1471),.clk(gclk));
	jnot g0830(.din(w_in1104_0[0]),.dout(n1472),.clk(gclk));
	jand g0831(.dina(w_n1472_0[1]),.dinb(w_in0104_0[0]),.dout(n1473),.clk(gclk));
	jand g0832(.dina(n1473),.dinb(n1471),.dout(n1474),.clk(gclk));
	jor g0833(.dina(n1474),.dinb(n1470),.dout(n1475),.clk(gclk));
	jand g0834(.dina(n1475),.dinb(w_n1465_0[1]),.dout(n1476),.clk(gclk));
	jnot g0835(.din(w_n1476_0[1]),.dout(n1477),.clk(gclk));
	jand g0836(.dina(n1477),.dinb(n1464),.dout(n1478),.clk(gclk));
	jand g0837(.dina(n1478),.dinb(n708),.dout(n1479),.clk(gclk));
	jnot g0838(.din(w_in0108_0[0]),.dout(n1480),.clk(gclk));
	jand g0839(.dina(w_in1108_0[0]),.dinb(w_n1480_0[1]),.dout(n1481),.clk(gclk));
	jor g0840(.dina(n1481),.dinb(w_n689_0[0]),.dout(n1482),.clk(gclk));
	jor g0841(.dina(w_n1482_0[1]),.dinb(n1479),.dout(n1483),.clk(gclk));
	jand g0842(.dina(n1483),.dinb(n705),.dout(n1484),.clk(gclk));
	jnot g0843(.din(w_in0115_0[0]),.dout(n1485),.clk(gclk));
	jand g0844(.dina(w_in1115_0[0]),.dinb(w_n1485_0[1]),.dout(n1486),.clk(gclk));
	jnot g0845(.din(w_in0114_0[1]),.dout(n1487),.clk(gclk));
	jand g0846(.dina(w_in1114_0[1]),.dinb(w_n1487_0[1]),.dout(n1488),.clk(gclk));
	jor g0847(.dina(n1488),.dinb(n1486),.dout(n1489),.clk(gclk));
	jor g0848(.dina(w_n1489_0[1]),.dinb(n1484),.dout(n1490),.clk(gclk));
	jor g0849(.dina(n1490),.dinb(w_n681_0[1]),.dout(n1491),.clk(gclk));
	jnot g0850(.din(w_n1489_0[0]),.dout(n1492),.clk(gclk));
	jnot g0851(.din(w_in1113_0[0]),.dout(n1493),.clk(gclk));
	jand g0852(.dina(w_n1493_0[1]),.dinb(w_in0113_0[0]),.dout(n1494),.clk(gclk));
	jnot g0853(.din(w_in1114_0[0]),.dout(n1495),.clk(gclk));
	jand g0854(.dina(w_n1495_0[1]),.dinb(w_in0114_0[0]),.dout(n1496),.clk(gclk));
	jor g0855(.dina(n1496),.dinb(n1494),.dout(n1497),.clk(gclk));
	jnot g0856(.din(w_n678_0[0]),.dout(n1498),.clk(gclk));
	jnot g0857(.din(w_in1112_0[0]),.dout(n1499),.clk(gclk));
	jand g0858(.dina(w_n1499_0[1]),.dinb(w_in0112_0[0]),.dout(n1500),.clk(gclk));
	jand g0859(.dina(n1500),.dinb(n1498),.dout(n1501),.clk(gclk));
	jor g0860(.dina(n1501),.dinb(n1497),.dout(n1502),.clk(gclk));
	jand g0861(.dina(n1502),.dinb(w_n1492_0[1]),.dout(n1503),.clk(gclk));
	jnot g0862(.din(w_n1503_0[1]),.dout(n1504),.clk(gclk));
	jand g0863(.dina(n1504),.dinb(n1491),.dout(n1505),.clk(gclk));
	jand g0864(.dina(n1505),.dinb(n676),.dout(n1506),.clk(gclk));
	jnot g0865(.din(w_in0116_0[0]),.dout(n1507),.clk(gclk));
	jand g0866(.dina(w_in1116_0[0]),.dinb(w_n1507_0[1]),.dout(n1508),.clk(gclk));
	jor g0867(.dina(n1508),.dinb(w_n657_0[0]),.dout(n1509),.clk(gclk));
	jor g0868(.dina(w_n1509_0[1]),.dinb(n1506),.dout(n1510),.clk(gclk));
	jand g0869(.dina(n1510),.dinb(n673),.dout(n1511),.clk(gclk));
	jnot g0870(.din(w_in0123_0[0]),.dout(n1512),.clk(gclk));
	jand g0871(.dina(w_in1123_0[0]),.dinb(w_n1512_0[1]),.dout(n1513),.clk(gclk));
	jnot g0872(.din(w_in0122_0[1]),.dout(n1514),.clk(gclk));
	jand g0873(.dina(w_in1122_0[1]),.dinb(w_n1514_0[1]),.dout(n1515),.clk(gclk));
	jor g0874(.dina(n1515),.dinb(n1513),.dout(n1516),.clk(gclk));
	jor g0875(.dina(w_n1516_0[1]),.dinb(n1511),.dout(n1517),.clk(gclk));
	jor g0876(.dina(n1517),.dinb(w_n649_0[1]),.dout(n1518),.clk(gclk));
	jnot g0877(.din(w_n1516_0[0]),.dout(n1519),.clk(gclk));
	jnot g0878(.din(w_in1121_0[0]),.dout(n1520),.clk(gclk));
	jand g0879(.dina(w_n1520_0[1]),.dinb(w_in0121_0[0]),.dout(n1521),.clk(gclk));
	jnot g0880(.din(w_in1122_0[0]),.dout(n1522),.clk(gclk));
	jand g0881(.dina(w_n1522_0[1]),.dinb(w_in0122_0[0]),.dout(n1523),.clk(gclk));
	jor g0882(.dina(n1523),.dinb(n1521),.dout(n1524),.clk(gclk));
	jnot g0883(.din(w_n648_0[0]),.dout(n1525),.clk(gclk));
	jnot g0884(.din(w_in1120_0[0]),.dout(n1526),.clk(gclk));
	jand g0885(.dina(w_n1526_0[1]),.dinb(w_in0120_0[0]),.dout(n1527),.clk(gclk));
	jand g0886(.dina(n1527),.dinb(n1525),.dout(n1528),.clk(gclk));
	jor g0887(.dina(n1528),.dinb(n1524),.dout(n1529),.clk(gclk));
	jand g0888(.dina(n1529),.dinb(w_n1519_0[1]),.dout(n1530),.clk(gclk));
	jnot g0889(.din(w_n1530_0[1]),.dout(n1531),.clk(gclk));
	jand g0890(.dina(n1531),.dinb(n1518),.dout(n1532),.clk(gclk));
	jand g0891(.dina(n1532),.dinb(n644),.dout(n1533),.clk(gclk));
	jnot g0892(.din(w_in0126_0[1]),.dout(n1534),.clk(gclk));
	jand g0893(.dina(w_in1126_0[1]),.dinb(w_n1534_0[1]),.dout(n1535),.clk(gclk));
	jnot g0894(.din(w_in0125_0[1]),.dout(n1536),.clk(gclk));
	jand g0895(.dina(w_in1125_0[1]),.dinb(w_n1536_0[1]),.dout(n1537),.clk(gclk));
	jor g0896(.dina(n1537),.dinb(n1535),.dout(n1538),.clk(gclk));
	jnot g0897(.din(w_in0124_0[1]),.dout(n1539),.clk(gclk));
	jand g0898(.dina(w_in1124_0[1]),.dinb(w_n1539_0[1]),.dout(n1540),.clk(gclk));
	jnot g0899(.din(w_in1127_0[2]),.dout(n1541),.clk(gclk));
	jand g0900(.dina(n1541),.dinb(w_in0127_0[2]),.dout(n1542),.clk(gclk));
	jor g0901(.dina(w_n1542_0[1]),.dinb(n1540),.dout(n1543),.clk(gclk));
	jor g0902(.dina(n1543),.dinb(w_n1538_0[1]),.dout(n1544),.clk(gclk));
	jor g0903(.dina(w_n1544_0[1]),.dinb(n1533),.dout(n1545),.clk(gclk));
	jnot g0904(.din(w_n1542_0[0]),.dout(n1546),.clk(gclk));
	jnot g0905(.din(w_n1538_0[0]),.dout(n1547),.clk(gclk));
	jnot g0906(.din(w_in1124_0[0]),.dout(n1548),.clk(gclk));
	jand g0907(.dina(w_n1548_0[1]),.dinb(w_in0124_0[0]),.dout(n1549),.clk(gclk));
	jnot g0908(.din(w_in1125_0[0]),.dout(n1550),.clk(gclk));
	jand g0909(.dina(w_n1550_0[1]),.dinb(w_in0125_0[0]),.dout(n1551),.clk(gclk));
	jor g0910(.dina(n1551),.dinb(n1549),.dout(n1552),.clk(gclk));
	jand g0911(.dina(n1552),.dinb(n1547),.dout(n1553),.clk(gclk));
	jnot g0912(.din(w_in1126_0[0]),.dout(n1554),.clk(gclk));
	jand g0913(.dina(w_n1554_0[1]),.dinb(w_in0126_0[0]),.dout(n1555),.clk(gclk));
	jnot g0914(.din(w_in0127_0[1]),.dout(n1556),.clk(gclk));
	jand g0915(.dina(w_in1127_0[1]),.dinb(n1556),.dout(n1557),.clk(gclk));
	jor g0916(.dina(n1557),.dinb(n1555),.dout(n1558),.clk(gclk));
	jor g0917(.dina(n1558),.dinb(n1553),.dout(n1559),.clk(gclk));
	jand g0918(.dina(n1559),.dinb(n1546),.dout(n1560),.clk(gclk));
	jnot g0919(.din(w_n1560_0[1]),.dout(n1561),.clk(gclk));
	jand g0920(.dina(n1561),.dinb(n1545),.dout(n1562),.clk(gclk));
	jor g0921(.dina(w_n1562_64[2]),.dinb(w_in00_0[1]),.dout(n1563),.clk(gclk));
	jnot g0922(.din(w_n649_0[0]),.dout(n1564),.clk(gclk));
	jnot g0923(.din(w_n681_0[0]),.dout(n1565),.clk(gclk));
	jnot g0924(.din(w_n713_0[0]),.dout(n1566),.clk(gclk));
	jnot g0925(.din(w_n745_0[0]),.dout(n1567),.clk(gclk));
	jnot g0926(.din(w_n804_0[0]),.dout(n1568),.clk(gclk));
	jnot g0927(.din(w_n836_0[0]),.dout(n1569),.clk(gclk));
	jnot g0928(.din(w_n974_0[0]),.dout(n1570),.clk(gclk));
	jnot g0929(.din(w_n979_0[0]),.dout(n1571),.clk(gclk));
	jnot g0930(.din(w_n984_0[0]),.dout(n1572),.clk(gclk));
	jnot g0931(.din(w_n989_0[0]),.dout(n1573),.clk(gclk));
	jnot g0932(.din(w_n994_0[0]),.dout(n1574),.clk(gclk));
	jnot g0933(.din(w_n996_0[0]),.dout(n1575),.clk(gclk));
	jnot g0934(.din(w_n1001_0[0]),.dout(n1576),.clk(gclk));
	jnot g0935(.din(w_n1006_0[0]),.dout(n1577),.clk(gclk));
	jnot g0936(.din(w_n1011_0[0]),.dout(n1578),.clk(gclk));
	jnot g0937(.din(w_n1016_0[0]),.dout(n1579),.clk(gclk));
	jnot g0938(.din(w_n1018_0[0]),.dout(n1580),.clk(gclk));
	jnot g0939(.din(w_n1023_0[0]),.dout(n1581),.clk(gclk));
	jnot g0940(.din(w_n1028_0[0]),.dout(n1582),.clk(gclk));
	jnot g0941(.din(w_n1033_0[0]),.dout(n1583),.clk(gclk));
	jnot g0942(.din(w_n1038_0[0]),.dout(n1584),.clk(gclk));
	jnot g0943(.din(w_n1040_0[0]),.dout(n1585),.clk(gclk));
	jnot g0944(.din(w_in11_0[2]),.dout(n1586),.clk(gclk));
	jand g0945(.dina(w_n1586_0[2]),.dinb(w_in01_1[0]),.dout(n1587),.clk(gclk));
	jnot g0946(.din(w_in10_0[1]),.dout(n1588),.clk(gclk));
	jand g0947(.dina(w_n1588_0[1]),.dinb(w_in00_0[0]),.dout(n1589),.clk(gclk));
	jor g0948(.dina(n1589),.dinb(n1587),.dout(n1590),.clk(gclk));
	jor g0949(.dina(w_n1041_0[1]),.dinb(w_in02_0[2]),.dout(n1591),.clk(gclk));
	jor g0950(.dina(w_n1586_0[1]),.dinb(w_in01_0[2]),.dout(n1592),.clk(gclk));
	jand g0951(.dina(n1592),.dinb(n1591),.dout(n1593),.clk(gclk));
	jand g0952(.dina(n1593),.dinb(n1590),.dout(n1594),.clk(gclk));
	jor g0953(.dina(w_n1055_0[0]),.dinb(n1594),.dout(n1595),.clk(gclk));
	jor g0954(.dina(n1595),.dinb(w_n1042_0[0]),.dout(n1596),.clk(gclk));
	jnot g0955(.din(w_n1060_0[0]),.dout(n1597),.clk(gclk));
	jand g0956(.dina(n1597),.dinb(n1596),.dout(n1598),.clk(gclk));
	jand g0957(.dina(n1598),.dinb(n1585),.dout(n1599),.clk(gclk));
	jor g0958(.dina(w_n1067_0[0]),.dinb(n1599),.dout(n1600),.clk(gclk));
	jnot g0959(.din(w_n1074_0[0]),.dout(n1601),.clk(gclk));
	jand g0960(.dina(n1601),.dinb(n1600),.dout(n1602),.clk(gclk));
	jor g0961(.dina(w_n1080_0[0]),.dinb(n1602),.dout(n1603),.clk(gclk));
	jnot g0962(.din(w_n1084_0[0]),.dout(n1604),.clk(gclk));
	jand g0963(.dina(n1604),.dinb(n1603),.dout(n1605),.clk(gclk));
	jand g0964(.dina(n1605),.dinb(n1584),.dout(n1606),.clk(gclk));
	jor g0965(.dina(w_n1091_0[0]),.dinb(n1606),.dout(n1607),.clk(gclk));
	jnot g0966(.din(w_n1098_0[0]),.dout(n1608),.clk(gclk));
	jand g0967(.dina(n1608),.dinb(n1607),.dout(n1609),.clk(gclk));
	jor g0968(.dina(n1609),.dinb(w_n1035_0[0]),.dout(n1610),.clk(gclk));
	jand g0969(.dina(n1610),.dinb(n1583),.dout(n1611),.clk(gclk));
	jor g0970(.dina(n1611),.dinb(w_n1030_0[0]),.dout(n1612),.clk(gclk));
	jand g0971(.dina(n1612),.dinb(n1582),.dout(n1613),.clk(gclk));
	jor g0972(.dina(n1613),.dinb(w_n1025_0[0]),.dout(n1614),.clk(gclk));
	jand g0973(.dina(n1614),.dinb(n1581),.dout(n1615),.clk(gclk));
	jor g0974(.dina(n1615),.dinb(w_n1020_0[0]),.dout(n1616),.clk(gclk));
	jand g0975(.dina(n1616),.dinb(n1580),.dout(n1617),.clk(gclk));
	jor g0976(.dina(w_n1112_0[0]),.dinb(n1617),.dout(n1618),.clk(gclk));
	jnot g0977(.din(w_n1116_0[0]),.dout(n1619),.clk(gclk));
	jand g0978(.dina(n1619),.dinb(n1618),.dout(n1620),.clk(gclk));
	jand g0979(.dina(n1620),.dinb(n1579),.dout(n1621),.clk(gclk));
	jor g0980(.dina(w_n1123_0[0]),.dinb(n1621),.dout(n1622),.clk(gclk));
	jnot g0981(.din(w_n1130_0[0]),.dout(n1623),.clk(gclk));
	jand g0982(.dina(n1623),.dinb(n1622),.dout(n1624),.clk(gclk));
	jor g0983(.dina(n1624),.dinb(w_n1013_0[0]),.dout(n1625),.clk(gclk));
	jand g0984(.dina(n1625),.dinb(n1578),.dout(n1626),.clk(gclk));
	jor g0985(.dina(n1626),.dinb(w_n1008_0[0]),.dout(n1627),.clk(gclk));
	jand g0986(.dina(n1627),.dinb(n1577),.dout(n1628),.clk(gclk));
	jor g0987(.dina(n1628),.dinb(w_n1003_0[0]),.dout(n1629),.clk(gclk));
	jand g0988(.dina(n1629),.dinb(n1576),.dout(n1630),.clk(gclk));
	jor g0989(.dina(n1630),.dinb(w_n998_0[0]),.dout(n1631),.clk(gclk));
	jand g0990(.dina(n1631),.dinb(n1575),.dout(n1632),.clk(gclk));
	jor g0991(.dina(w_n1144_0[0]),.dinb(n1632),.dout(n1633),.clk(gclk));
	jnot g0992(.din(w_n1148_0[0]),.dout(n1634),.clk(gclk));
	jand g0993(.dina(n1634),.dinb(n1633),.dout(n1635),.clk(gclk));
	jand g0994(.dina(n1635),.dinb(n1574),.dout(n1636),.clk(gclk));
	jor g0995(.dina(w_n1155_0[0]),.dinb(n1636),.dout(n1637),.clk(gclk));
	jnot g0996(.din(w_n1162_0[0]),.dout(n1638),.clk(gclk));
	jand g0997(.dina(n1638),.dinb(n1637),.dout(n1639),.clk(gclk));
	jor g0998(.dina(n1639),.dinb(w_n991_0[0]),.dout(n1640),.clk(gclk));
	jand g0999(.dina(n1640),.dinb(n1573),.dout(n1641),.clk(gclk));
	jor g1000(.dina(n1641),.dinb(w_n986_0[0]),.dout(n1642),.clk(gclk));
	jand g1001(.dina(n1642),.dinb(n1572),.dout(n1643),.clk(gclk));
	jor g1002(.dina(n1643),.dinb(w_n981_0[0]),.dout(n1644),.clk(gclk));
	jand g1003(.dina(n1644),.dinb(n1571),.dout(n1645),.clk(gclk));
	jor g1004(.dina(n1645),.dinb(w_n976_0[0]),.dout(n1646),.clk(gclk));
	jand g1005(.dina(n1646),.dinb(n1570),.dout(n1647),.clk(gclk));
	jor g1006(.dina(w_n1176_0[0]),.dinb(n1647),.dout(n1648),.clk(gclk));
	jnot g1007(.din(w_n1185_0[0]),.dout(n1649),.clk(gclk));
	jand g1008(.dina(n1649),.dinb(n1648),.dout(n1650),.clk(gclk));
	jor g1009(.dina(w_n1206_0[0]),.dinb(n1650),.dout(n1651),.clk(gclk));
	jor g1010(.dina(n1651),.dinb(w_n971_0[0]),.dout(n1652),.clk(gclk));
	jnot g1011(.din(w_n1213_0[0]),.dout(n1653),.clk(gclk));
	jand g1012(.dina(n1653),.dinb(n1652),.dout(n1654),.clk(gclk));
	jnot g1013(.din(w_n1233_0[0]),.dout(n1655),.clk(gclk));
	jor g1014(.dina(n1655),.dinb(n1654),.dout(n1656),.clk(gclk));
	jor g1015(.dina(n1656),.dinb(w_n939_0[0]),.dout(n1657),.clk(gclk));
	jand g1016(.dina(w_n1250_0[0]),.dinb(n1657),.dout(n1658),.clk(gclk));
	jor g1017(.dina(w_n1278_0[0]),.dinb(n1658),.dout(n1659),.clk(gclk));
	jor g1018(.dina(n1659),.dinb(w_n907_0[0]),.dout(n1660),.clk(gclk));
	jand g1019(.dina(w_n1296_0[0]),.dinb(n1660),.dout(n1661),.clk(gclk));
	jor g1020(.dina(w_n1324_0[0]),.dinb(n1661),.dout(n1662),.clk(gclk));
	jor g1021(.dina(n1662),.dinb(w_n891_0[0]),.dout(n1663),.clk(gclk));
	jnot g1022(.din(w_n1330_0[0]),.dout(n1664),.clk(gclk));
	jand g1023(.dina(n1664),.dinb(n1663),.dout(n1665),.clk(gclk));
	jor g1024(.dina(n1665),.dinb(w_n875_0[0]),.dout(n1666),.clk(gclk));
	jnot g1025(.din(w_n1337_0[0]),.dout(n1667),.clk(gclk));
	jand g1026(.dina(n1667),.dinb(n1666),.dout(n1668),.clk(gclk));
	jor g1027(.dina(n1668),.dinb(w_n862_0[0]),.dout(n1669),.clk(gclk));
	jnot g1028(.din(w_n1342_0[0]),.dout(n1670),.clk(gclk));
	jand g1029(.dina(n1670),.dinb(n1669),.dout(n1671),.clk(gclk));
	jor g1030(.dina(n1671),.dinb(w_n859_0[0]),.dout(n1672),.clk(gclk));
	jand g1031(.dina(w_n1352_0[0]),.dinb(n1672),.dout(n1673),.clk(gclk));
	jand g1032(.dina(n1673),.dinb(n1569),.dout(n1674),.clk(gclk));
	jor g1033(.dina(w_n1363_0[0]),.dinb(n1674),.dout(n1675),.clk(gclk));
	jor g1034(.dina(n1675),.dinb(w_n830_0[0]),.dout(n1676),.clk(gclk));
	jnot g1035(.din(w_n1369_0[0]),.dout(n1677),.clk(gclk));
	jand g1036(.dina(n1677),.dinb(n1676),.dout(n1678),.clk(gclk));
	jor g1037(.dina(n1678),.dinb(w_n827_0[0]),.dout(n1679),.clk(gclk));
	jand g1038(.dina(w_n1379_0[0]),.dinb(n1679),.dout(n1680),.clk(gclk));
	jand g1039(.dina(n1680),.dinb(n1568),.dout(n1681),.clk(gclk));
	jor g1040(.dina(w_n1390_0[0]),.dinb(n1681),.dout(n1682),.clk(gclk));
	jor g1041(.dina(n1682),.dinb(w_n798_0[0]),.dout(n1683),.clk(gclk));
	jnot g1042(.din(w_n1396_0[0]),.dout(n1684),.clk(gclk));
	jand g1043(.dina(n1684),.dinb(n1683),.dout(n1685),.clk(gclk));
	jor g1044(.dina(n1685),.dinb(w_n795_0[0]),.dout(n1686),.clk(gclk));
	jnot g1045(.din(w_n1409_0[0]),.dout(n1687),.clk(gclk));
	jand g1046(.dina(n1687),.dinb(n1686),.dout(n1688),.clk(gclk));
	jor g1047(.dina(w_n1422_0[0]),.dinb(n1688),.dout(n1689),.clk(gclk));
	jor g1048(.dina(n1689),.dinb(w_n771_0[0]),.dout(n1690),.clk(gclk));
	jnot g1049(.din(w_n1428_0[0]),.dout(n1691),.clk(gclk));
	jand g1050(.dina(n1691),.dinb(n1690),.dout(n1692),.clk(gclk));
	jor g1051(.dina(n1692),.dinb(w_n768_0[0]),.dout(n1693),.clk(gclk));
	jand g1052(.dina(w_n1438_0[0]),.dinb(n1693),.dout(n1694),.clk(gclk));
	jand g1053(.dina(n1694),.dinb(n1567),.dout(n1695),.clk(gclk));
	jor g1054(.dina(w_n1449_0[0]),.dinb(n1695),.dout(n1696),.clk(gclk));
	jor g1055(.dina(n1696),.dinb(w_n739_0[0]),.dout(n1697),.clk(gclk));
	jnot g1056(.din(w_n1455_0[0]),.dout(n1698),.clk(gclk));
	jand g1057(.dina(n1698),.dinb(n1697),.dout(n1699),.clk(gclk));
	jor g1058(.dina(n1699),.dinb(w_n736_0[0]),.dout(n1700),.clk(gclk));
	jand g1059(.dina(w_n1465_0[0]),.dinb(n1700),.dout(n1701),.clk(gclk));
	jand g1060(.dina(n1701),.dinb(n1566),.dout(n1702),.clk(gclk));
	jor g1061(.dina(w_n1476_0[0]),.dinb(n1702),.dout(n1703),.clk(gclk));
	jor g1062(.dina(n1703),.dinb(w_n707_0[0]),.dout(n1704),.clk(gclk));
	jnot g1063(.din(w_n1482_0[0]),.dout(n1705),.clk(gclk));
	jand g1064(.dina(n1705),.dinb(n1704),.dout(n1706),.clk(gclk));
	jor g1065(.dina(n1706),.dinb(w_n704_0[0]),.dout(n1707),.clk(gclk));
	jand g1066(.dina(w_n1492_0[0]),.dinb(n1707),.dout(n1708),.clk(gclk));
	jand g1067(.dina(n1708),.dinb(n1565),.dout(n1709),.clk(gclk));
	jor g1068(.dina(w_n1503_0[0]),.dinb(n1709),.dout(n1710),.clk(gclk));
	jor g1069(.dina(n1710),.dinb(w_n675_0[0]),.dout(n1711),.clk(gclk));
	jnot g1070(.din(w_n1509_0[0]),.dout(n1712),.clk(gclk));
	jand g1071(.dina(n1712),.dinb(n1711),.dout(n1713),.clk(gclk));
	jor g1072(.dina(n1713),.dinb(w_n672_0[0]),.dout(n1714),.clk(gclk));
	jand g1073(.dina(w_n1519_0[0]),.dinb(n1714),.dout(n1715),.clk(gclk));
	jand g1074(.dina(n1715),.dinb(n1564),.dout(n1716),.clk(gclk));
	jor g1075(.dina(w_n1530_0[0]),.dinb(n1716),.dout(n1717),.clk(gclk));
	jor g1076(.dina(n1717),.dinb(w_n643_0[0]),.dout(n1718),.clk(gclk));
	jnot g1077(.din(w_n1544_0[0]),.dout(n1719),.clk(gclk));
	jand g1078(.dina(n1719),.dinb(n1718),.dout(n1720),.clk(gclk));
	jor g1079(.dina(w_n1560_0[0]),.dinb(n1720),.dout(n1721),.clk(gclk));
	jor g1080(.dina(w_n1721_65[1]),.dinb(w_in10_0[0]),.dout(n1722),.clk(gclk));
	jand g1081(.dina(n1722),.dinb(n1563),.dout(n1723),.clk(gclk));
	jnot g1082(.din(w_in2126_0[1]),.dout(n1724),.clk(gclk));
	jand g1083(.dina(w_in3126_0[1]),.dinb(w_n1724_0[1]),.dout(n1725),.clk(gclk));
	jnot g1084(.din(w_in2125_0[1]),.dout(n1726),.clk(gclk));
	jand g1085(.dina(w_in3125_0[1]),.dinb(w_n1726_0[1]),.dout(n1727),.clk(gclk));
	jor g1086(.dina(n1727),.dinb(n1725),.dout(n1728),.clk(gclk));
	jnot g1087(.din(w_n1728_0[1]),.dout(n1729),.clk(gclk));
	jnot g1088(.din(w_in3124_0[1]),.dout(n1730),.clk(gclk));
	jand g1089(.dina(w_n1730_0[1]),.dinb(w_in2124_0[1]),.dout(n1731),.clk(gclk));
	jnot g1090(.din(w_in3125_0[0]),.dout(n1732),.clk(gclk));
	jand g1091(.dina(w_n1732_0[1]),.dinb(w_in2125_0[0]),.dout(n1733),.clk(gclk));
	jor g1092(.dina(n1733),.dinb(n1731),.dout(n1734),.clk(gclk));
	jand g1093(.dina(n1734),.dinb(n1729),.dout(n1735),.clk(gclk));
	jnot g1094(.din(w_in3126_0[0]),.dout(n1736),.clk(gclk));
	jand g1095(.dina(w_n1736_0[1]),.dinb(w_in2126_0[0]),.dout(n1737),.clk(gclk));
	jor g1096(.dina(n1737),.dinb(n1735),.dout(n1738),.clk(gclk));
	jnot g1097(.din(w_n1738_0[1]),.dout(n1739),.clk(gclk));
	jnot g1098(.din(w_in3123_0[1]),.dout(n1740),.clk(gclk));
	jand g1099(.dina(w_n1740_0[1]),.dinb(w_in2123_0[1]),.dout(n1741),.clk(gclk));
	jnot g1100(.din(w_n1741_0[1]),.dout(n1742),.clk(gclk));
	jnot g1101(.din(w_in2118_0[1]),.dout(n1743),.clk(gclk));
	jand g1102(.dina(w_in3118_0[1]),.dinb(w_n1743_0[1]),.dout(n1744),.clk(gclk));
	jnot g1103(.din(w_in2119_0[1]),.dout(n1745),.clk(gclk));
	jand g1104(.dina(w_in3119_0[1]),.dinb(w_n1745_0[1]),.dout(n1746),.clk(gclk));
	jnot g1105(.din(w_in2117_0[1]),.dout(n1747),.clk(gclk));
	jand g1106(.dina(w_in3117_0[1]),.dinb(w_n1747_0[1]),.dout(n1748),.clk(gclk));
	jor g1107(.dina(n1748),.dinb(w_n1746_0[1]),.dout(n1749),.clk(gclk));
	jor g1108(.dina(n1749),.dinb(n1744),.dout(n1750),.clk(gclk));
	jnot g1109(.din(w_n1750_0[1]),.dout(n1751),.clk(gclk));
	jnot g1110(.din(w_in3117_0[0]),.dout(n1752),.clk(gclk));
	jand g1111(.dina(w_n1752_0[1]),.dinb(w_in2117_0[0]),.dout(n1753),.clk(gclk));
	jnot g1112(.din(w_in3116_0[1]),.dout(n1754),.clk(gclk));
	jand g1113(.dina(w_n1754_0[1]),.dinb(w_in2116_0[1]),.dout(n1755),.clk(gclk));
	jor g1114(.dina(n1755),.dinb(n1753),.dout(n1756),.clk(gclk));
	jand g1115(.dina(n1756),.dinb(n1751),.dout(n1757),.clk(gclk));
	jnot g1116(.din(w_n1746_0[0]),.dout(n1758),.clk(gclk));
	jnot g1117(.din(w_in3119_0[0]),.dout(n1759),.clk(gclk));
	jand g1118(.dina(w_n1759_0[1]),.dinb(w_in2119_0[0]),.dout(n1760),.clk(gclk));
	jnot g1119(.din(w_in3118_0[0]),.dout(n1761),.clk(gclk));
	jand g1120(.dina(w_n1761_0[1]),.dinb(w_in2118_0[0]),.dout(n1762),.clk(gclk));
	jor g1121(.dina(n1762),.dinb(n1760),.dout(n1763),.clk(gclk));
	jand g1122(.dina(n1763),.dinb(n1758),.dout(n1764),.clk(gclk));
	jor g1123(.dina(n1764),.dinb(n1757),.dout(n1765),.clk(gclk));
	jnot g1124(.din(w_n1765_0[1]),.dout(n1766),.clk(gclk));
	jnot g1125(.din(w_in3115_0[1]),.dout(n1767),.clk(gclk));
	jand g1126(.dina(w_n1767_0[1]),.dinb(w_in2115_0[1]),.dout(n1768),.clk(gclk));
	jnot g1127(.din(w_n1768_0[1]),.dout(n1769),.clk(gclk));
	jnot g1128(.din(w_in2113_0[1]),.dout(n1770),.clk(gclk));
	jand g1129(.dina(w_in3113_0[1]),.dinb(w_n1770_0[1]),.dout(n1771),.clk(gclk));
	jnot g1130(.din(w_in2112_0[1]),.dout(n1772),.clk(gclk));
	jand g1131(.dina(w_in3112_0[1]),.dinb(w_n1772_0[1]),.dout(n1773),.clk(gclk));
	jor g1132(.dina(n1773),.dinb(w_n1771_0[1]),.dout(n1774),.clk(gclk));
	jnot g1133(.din(w_in2110_0[1]),.dout(n1775),.clk(gclk));
	jand g1134(.dina(w_in3110_0[1]),.dinb(w_n1775_0[1]),.dout(n1776),.clk(gclk));
	jnot g1135(.din(w_in2111_0[1]),.dout(n1777),.clk(gclk));
	jand g1136(.dina(w_in3111_0[1]),.dinb(w_n1777_0[1]),.dout(n1778),.clk(gclk));
	jnot g1137(.din(w_in2109_0[1]),.dout(n1779),.clk(gclk));
	jand g1138(.dina(w_in3109_0[1]),.dinb(w_n1779_0[1]),.dout(n1780),.clk(gclk));
	jor g1139(.dina(n1780),.dinb(w_n1778_0[1]),.dout(n1781),.clk(gclk));
	jor g1140(.dina(n1781),.dinb(n1776),.dout(n1782),.clk(gclk));
	jnot g1141(.din(w_n1782_0[1]),.dout(n1783),.clk(gclk));
	jnot g1142(.din(w_in3109_0[0]),.dout(n1784),.clk(gclk));
	jand g1143(.dina(w_n1784_0[1]),.dinb(w_in2109_0[0]),.dout(n1785),.clk(gclk));
	jnot g1144(.din(w_in3108_0[1]),.dout(n1786),.clk(gclk));
	jand g1145(.dina(w_n1786_0[1]),.dinb(w_in2108_0[1]),.dout(n1787),.clk(gclk));
	jor g1146(.dina(n1787),.dinb(n1785),.dout(n1788),.clk(gclk));
	jand g1147(.dina(n1788),.dinb(n1783),.dout(n1789),.clk(gclk));
	jnot g1148(.din(w_n1778_0[0]),.dout(n1790),.clk(gclk));
	jnot g1149(.din(w_in3111_0[0]),.dout(n1791),.clk(gclk));
	jand g1150(.dina(w_n1791_0[1]),.dinb(w_in2111_0[0]),.dout(n1792),.clk(gclk));
	jnot g1151(.din(w_in3110_0[0]),.dout(n1793),.clk(gclk));
	jand g1152(.dina(w_n1793_0[1]),.dinb(w_in2110_0[0]),.dout(n1794),.clk(gclk));
	jor g1153(.dina(n1794),.dinb(n1792),.dout(n1795),.clk(gclk));
	jand g1154(.dina(n1795),.dinb(n1790),.dout(n1796),.clk(gclk));
	jor g1155(.dina(n1796),.dinb(n1789),.dout(n1797),.clk(gclk));
	jnot g1156(.din(w_n1797_0[1]),.dout(n1798),.clk(gclk));
	jnot g1157(.din(w_in3107_0[1]),.dout(n1799),.clk(gclk));
	jand g1158(.dina(w_n1799_0[1]),.dinb(w_in2107_0[1]),.dout(n1800),.clk(gclk));
	jnot g1159(.din(w_n1800_0[1]),.dout(n1801),.clk(gclk));
	jnot g1160(.din(w_in2102_0[1]),.dout(n1802),.clk(gclk));
	jand g1161(.dina(w_in3102_0[1]),.dinb(w_n1802_0[1]),.dout(n1803),.clk(gclk));
	jnot g1162(.din(w_in2103_0[1]),.dout(n1804),.clk(gclk));
	jand g1163(.dina(w_in3103_0[1]),.dinb(w_n1804_0[1]),.dout(n1805),.clk(gclk));
	jnot g1164(.din(w_in2101_0[1]),.dout(n1806),.clk(gclk));
	jand g1165(.dina(w_in3101_0[1]),.dinb(w_n1806_0[1]),.dout(n1807),.clk(gclk));
	jor g1166(.dina(n1807),.dinb(w_n1805_0[1]),.dout(n1808),.clk(gclk));
	jor g1167(.dina(n1808),.dinb(n1803),.dout(n1809),.clk(gclk));
	jnot g1168(.din(w_n1809_0[1]),.dout(n1810),.clk(gclk));
	jnot g1169(.din(w_in3101_0[0]),.dout(n1811),.clk(gclk));
	jand g1170(.dina(w_n1811_0[1]),.dinb(w_in2101_0[0]),.dout(n1812),.clk(gclk));
	jnot g1171(.din(w_in3100_0[1]),.dout(n1813),.clk(gclk));
	jand g1172(.dina(w_n1813_0[1]),.dinb(w_in2100_0[1]),.dout(n1814),.clk(gclk));
	jor g1173(.dina(n1814),.dinb(n1812),.dout(n1815),.clk(gclk));
	jand g1174(.dina(n1815),.dinb(n1810),.dout(n1816),.clk(gclk));
	jnot g1175(.din(w_n1805_0[0]),.dout(n1817),.clk(gclk));
	jnot g1176(.din(w_in3103_0[0]),.dout(n1818),.clk(gclk));
	jand g1177(.dina(w_n1818_0[1]),.dinb(w_in2103_0[0]),.dout(n1819),.clk(gclk));
	jnot g1178(.din(w_in3102_0[0]),.dout(n1820),.clk(gclk));
	jand g1179(.dina(w_n1820_0[1]),.dinb(w_in2102_0[0]),.dout(n1821),.clk(gclk));
	jor g1180(.dina(n1821),.dinb(n1819),.dout(n1822),.clk(gclk));
	jand g1181(.dina(n1822),.dinb(n1817),.dout(n1823),.clk(gclk));
	jor g1182(.dina(n1823),.dinb(n1816),.dout(n1824),.clk(gclk));
	jnot g1183(.din(w_n1824_0[1]),.dout(n1825),.clk(gclk));
	jnot g1184(.din(w_in399_0[1]),.dout(n1826),.clk(gclk));
	jand g1185(.dina(w_n1826_0[1]),.dinb(w_in299_0[1]),.dout(n1827),.clk(gclk));
	jnot g1186(.din(w_n1827_0[1]),.dout(n1828),.clk(gclk));
	jnot g1187(.din(w_in297_0[1]),.dout(n1829),.clk(gclk));
	jand g1188(.dina(w_in397_0[1]),.dinb(w_n1829_0[1]),.dout(n1830),.clk(gclk));
	jnot g1189(.din(w_in296_0[1]),.dout(n1831),.clk(gclk));
	jand g1190(.dina(w_in396_0[1]),.dinb(w_n1831_0[1]),.dout(n1832),.clk(gclk));
	jor g1191(.dina(n1832),.dinb(w_n1830_0[1]),.dout(n1833),.clk(gclk));
	jnot g1192(.din(w_in294_0[1]),.dout(n1834),.clk(gclk));
	jand g1193(.dina(w_in394_0[1]),.dinb(w_n1834_0[1]),.dout(n1835),.clk(gclk));
	jnot g1194(.din(w_in295_0[1]),.dout(n1836),.clk(gclk));
	jand g1195(.dina(w_in395_0[1]),.dinb(w_n1836_0[1]),.dout(n1837),.clk(gclk));
	jnot g1196(.din(w_in293_0[1]),.dout(n1838),.clk(gclk));
	jand g1197(.dina(w_in393_0[1]),.dinb(w_n1838_0[1]),.dout(n1839),.clk(gclk));
	jor g1198(.dina(n1839),.dinb(w_n1837_0[1]),.dout(n1840),.clk(gclk));
	jor g1199(.dina(n1840),.dinb(n1835),.dout(n1841),.clk(gclk));
	jnot g1200(.din(w_n1841_0[1]),.dout(n1842),.clk(gclk));
	jnot g1201(.din(w_in393_0[0]),.dout(n1843),.clk(gclk));
	jand g1202(.dina(w_n1843_0[1]),.dinb(w_in293_0[0]),.dout(n1844),.clk(gclk));
	jnot g1203(.din(w_in392_0[1]),.dout(n1845),.clk(gclk));
	jand g1204(.dina(w_n1845_0[1]),.dinb(w_in292_0[1]),.dout(n1846),.clk(gclk));
	jor g1205(.dina(n1846),.dinb(n1844),.dout(n1847),.clk(gclk));
	jand g1206(.dina(n1847),.dinb(n1842),.dout(n1848),.clk(gclk));
	jnot g1207(.din(w_n1837_0[0]),.dout(n1849),.clk(gclk));
	jnot g1208(.din(w_in395_0[0]),.dout(n1850),.clk(gclk));
	jand g1209(.dina(w_n1850_0[1]),.dinb(w_in295_0[0]),.dout(n1851),.clk(gclk));
	jnot g1210(.din(w_in394_0[0]),.dout(n1852),.clk(gclk));
	jand g1211(.dina(w_n1852_0[1]),.dinb(w_in294_0[0]),.dout(n1853),.clk(gclk));
	jor g1212(.dina(n1853),.dinb(n1851),.dout(n1854),.clk(gclk));
	jand g1213(.dina(n1854),.dinb(n1849),.dout(n1855),.clk(gclk));
	jor g1214(.dina(n1855),.dinb(n1848),.dout(n1856),.clk(gclk));
	jnot g1215(.din(w_n1856_0[1]),.dout(n1857),.clk(gclk));
	jnot g1216(.din(w_in391_0[1]),.dout(n1858),.clk(gclk));
	jand g1217(.dina(w_n1858_0[1]),.dinb(w_in291_0[1]),.dout(n1859),.clk(gclk));
	jnot g1218(.din(w_n1859_0[1]),.dout(n1860),.clk(gclk));
	jnot g1219(.din(w_in286_0[1]),.dout(n1861),.clk(gclk));
	jand g1220(.dina(w_in386_0[1]),.dinb(w_n1861_0[1]),.dout(n1862),.clk(gclk));
	jnot g1221(.din(w_in287_0[1]),.dout(n1863),.clk(gclk));
	jand g1222(.dina(w_in387_0[1]),.dinb(w_n1863_0[1]),.dout(n1864),.clk(gclk));
	jnot g1223(.din(w_in285_0[1]),.dout(n1865),.clk(gclk));
	jand g1224(.dina(w_in385_0[1]),.dinb(w_n1865_0[1]),.dout(n1866),.clk(gclk));
	jor g1225(.dina(n1866),.dinb(w_n1864_0[1]),.dout(n1867),.clk(gclk));
	jor g1226(.dina(n1867),.dinb(n1862),.dout(n1868),.clk(gclk));
	jnot g1227(.din(w_n1868_0[1]),.dout(n1869),.clk(gclk));
	jnot g1228(.din(w_in385_0[0]),.dout(n1870),.clk(gclk));
	jand g1229(.dina(w_n1870_0[1]),.dinb(w_in285_0[0]),.dout(n1871),.clk(gclk));
	jnot g1230(.din(w_in384_0[1]),.dout(n1872),.clk(gclk));
	jand g1231(.dina(w_n1872_0[1]),.dinb(w_in284_0[1]),.dout(n1873),.clk(gclk));
	jor g1232(.dina(n1873),.dinb(n1871),.dout(n1874),.clk(gclk));
	jand g1233(.dina(n1874),.dinb(n1869),.dout(n1875),.clk(gclk));
	jnot g1234(.din(w_n1864_0[0]),.dout(n1876),.clk(gclk));
	jnot g1235(.din(w_in387_0[0]),.dout(n1877),.clk(gclk));
	jand g1236(.dina(w_n1877_0[1]),.dinb(w_in287_0[0]),.dout(n1878),.clk(gclk));
	jnot g1237(.din(w_in386_0[0]),.dout(n1879),.clk(gclk));
	jand g1238(.dina(w_n1879_0[1]),.dinb(w_in286_0[0]),.dout(n1880),.clk(gclk));
	jor g1239(.dina(n1880),.dinb(n1878),.dout(n1881),.clk(gclk));
	jand g1240(.dina(n1881),.dinb(n1876),.dout(n1882),.clk(gclk));
	jor g1241(.dina(n1882),.dinb(n1875),.dout(n1883),.clk(gclk));
	jnot g1242(.din(w_n1883_0[1]),.dout(n1884),.clk(gclk));
	jnot g1243(.din(w_in383_0[1]),.dout(n1885),.clk(gclk));
	jand g1244(.dina(w_n1885_0[1]),.dinb(w_in283_0[1]),.dout(n1886),.clk(gclk));
	jnot g1245(.din(w_n1886_0[1]),.dout(n1887),.clk(gclk));
	jnot g1246(.din(w_in281_0[1]),.dout(n1888),.clk(gclk));
	jand g1247(.dina(w_in381_0[1]),.dinb(w_n1888_0[1]),.dout(n1889),.clk(gclk));
	jnot g1248(.din(w_in280_0[1]),.dout(n1890),.clk(gclk));
	jand g1249(.dina(w_in380_0[1]),.dinb(w_n1890_0[1]),.dout(n1891),.clk(gclk));
	jor g1250(.dina(n1891),.dinb(w_n1889_0[1]),.dout(n1892),.clk(gclk));
	jnot g1251(.din(w_in278_0[1]),.dout(n1893),.clk(gclk));
	jand g1252(.dina(w_in378_0[1]),.dinb(w_n1893_0[1]),.dout(n1894),.clk(gclk));
	jnot g1253(.din(w_in279_0[1]),.dout(n1895),.clk(gclk));
	jand g1254(.dina(w_in379_0[1]),.dinb(w_n1895_0[1]),.dout(n1896),.clk(gclk));
	jnot g1255(.din(w_in277_0[1]),.dout(n1897),.clk(gclk));
	jand g1256(.dina(w_in377_0[1]),.dinb(w_n1897_0[1]),.dout(n1898),.clk(gclk));
	jor g1257(.dina(n1898),.dinb(w_n1896_0[1]),.dout(n1899),.clk(gclk));
	jor g1258(.dina(n1899),.dinb(n1894),.dout(n1900),.clk(gclk));
	jnot g1259(.din(w_n1900_0[1]),.dout(n1901),.clk(gclk));
	jnot g1260(.din(w_in377_0[0]),.dout(n1902),.clk(gclk));
	jand g1261(.dina(w_n1902_0[1]),.dinb(w_in277_0[0]),.dout(n1903),.clk(gclk));
	jnot g1262(.din(w_in376_0[1]),.dout(n1904),.clk(gclk));
	jand g1263(.dina(w_n1904_0[1]),.dinb(w_in276_0[1]),.dout(n1905),.clk(gclk));
	jor g1264(.dina(n1905),.dinb(n1903),.dout(n1906),.clk(gclk));
	jand g1265(.dina(n1906),.dinb(n1901),.dout(n1907),.clk(gclk));
	jnot g1266(.din(w_n1896_0[0]),.dout(n1908),.clk(gclk));
	jnot g1267(.din(w_in379_0[0]),.dout(n1909),.clk(gclk));
	jand g1268(.dina(w_n1909_0[1]),.dinb(w_in279_0[0]),.dout(n1910),.clk(gclk));
	jnot g1269(.din(w_in378_0[0]),.dout(n1911),.clk(gclk));
	jand g1270(.dina(w_n1911_0[1]),.dinb(w_in278_0[0]),.dout(n1912),.clk(gclk));
	jor g1271(.dina(n1912),.dinb(n1910),.dout(n1913),.clk(gclk));
	jand g1272(.dina(n1913),.dinb(n1908),.dout(n1914),.clk(gclk));
	jor g1273(.dina(n1914),.dinb(n1907),.dout(n1915),.clk(gclk));
	jnot g1274(.din(w_n1915_0[1]),.dout(n1916),.clk(gclk));
	jnot g1275(.din(w_in375_0[1]),.dout(n1917),.clk(gclk));
	jand g1276(.dina(w_n1917_0[1]),.dinb(w_in275_0[1]),.dout(n1918),.clk(gclk));
	jnot g1277(.din(w_n1918_0[1]),.dout(n1919),.clk(gclk));
	jnot g1278(.din(w_in270_0[1]),.dout(n1920),.clk(gclk));
	jand g1279(.dina(w_in370_0[1]),.dinb(w_n1920_0[1]),.dout(n1921),.clk(gclk));
	jnot g1280(.din(w_in271_0[1]),.dout(n1922),.clk(gclk));
	jand g1281(.dina(w_in371_0[1]),.dinb(w_n1922_0[1]),.dout(n1923),.clk(gclk));
	jnot g1282(.din(w_in269_0[1]),.dout(n1924),.clk(gclk));
	jand g1283(.dina(w_in369_0[1]),.dinb(w_n1924_0[1]),.dout(n1925),.clk(gclk));
	jor g1284(.dina(n1925),.dinb(w_n1923_0[1]),.dout(n1926),.clk(gclk));
	jor g1285(.dina(n1926),.dinb(n1921),.dout(n1927),.clk(gclk));
	jnot g1286(.din(w_n1927_0[1]),.dout(n1928),.clk(gclk));
	jnot g1287(.din(w_in369_0[0]),.dout(n1929),.clk(gclk));
	jand g1288(.dina(w_n1929_0[1]),.dinb(w_in269_0[0]),.dout(n1930),.clk(gclk));
	jnot g1289(.din(w_in368_0[1]),.dout(n1931),.clk(gclk));
	jand g1290(.dina(w_n1931_0[1]),.dinb(w_in268_0[1]),.dout(n1932),.clk(gclk));
	jor g1291(.dina(n1932),.dinb(n1930),.dout(n1933),.clk(gclk));
	jand g1292(.dina(n1933),.dinb(n1928),.dout(n1934),.clk(gclk));
	jnot g1293(.din(w_n1923_0[0]),.dout(n1935),.clk(gclk));
	jnot g1294(.din(w_in371_0[0]),.dout(n1936),.clk(gclk));
	jand g1295(.dina(w_n1936_0[1]),.dinb(w_in271_0[0]),.dout(n1937),.clk(gclk));
	jnot g1296(.din(w_in370_0[0]),.dout(n1938),.clk(gclk));
	jand g1297(.dina(w_n1938_0[1]),.dinb(w_in270_0[0]),.dout(n1939),.clk(gclk));
	jor g1298(.dina(n1939),.dinb(n1937),.dout(n1940),.clk(gclk));
	jand g1299(.dina(n1940),.dinb(n1935),.dout(n1941),.clk(gclk));
	jor g1300(.dina(n1941),.dinb(n1934),.dout(n1942),.clk(gclk));
	jnot g1301(.din(w_n1942_0[1]),.dout(n1943),.clk(gclk));
	jnot g1302(.din(w_in367_0[1]),.dout(n1944),.clk(gclk));
	jand g1303(.dina(w_n1944_0[1]),.dinb(w_in267_0[1]),.dout(n1945),.clk(gclk));
	jnot g1304(.din(w_n1945_0[1]),.dout(n1946),.clk(gclk));
	jnot g1305(.din(w_in265_0[1]),.dout(n1947),.clk(gclk));
	jand g1306(.dina(w_in365_0[1]),.dinb(w_n1947_0[1]),.dout(n1948),.clk(gclk));
	jnot g1307(.din(w_n1948_0[1]),.dout(n1949),.clk(gclk));
	jnot g1308(.din(w_in364_0[1]),.dout(n1950),.clk(gclk));
	jand g1309(.dina(w_n1950_0[1]),.dinb(w_in264_0[1]),.dout(n1951),.clk(gclk));
	jand g1310(.dina(n1951),.dinb(n1949),.dout(n1952),.clk(gclk));
	jnot g1311(.din(w_in366_0[1]),.dout(n1953),.clk(gclk));
	jand g1312(.dina(w_n1953_0[1]),.dinb(w_in266_0[1]),.dout(n1954),.clk(gclk));
	jnot g1313(.din(w_in365_0[0]),.dout(n1955),.clk(gclk));
	jand g1314(.dina(w_n1955_0[1]),.dinb(w_in265_0[0]),.dout(n1956),.clk(gclk));
	jor g1315(.dina(n1956),.dinb(n1954),.dout(n1957),.clk(gclk));
	jor g1316(.dina(n1957),.dinb(n1952),.dout(n1958),.clk(gclk));
	jnot g1317(.din(w_n1958_0[1]),.dout(n1959),.clk(gclk));
	jnot g1318(.din(w_in359_0[1]),.dout(n1960),.clk(gclk));
	jnot g1319(.din(w_in260_0[1]),.dout(n1961),.clk(gclk));
	jand g1320(.dina(w_in360_0[1]),.dinb(w_n1961_0[1]),.dout(n1962),.clk(gclk));
	jnot g1321(.din(w_in263_0[1]),.dout(n1963),.clk(gclk));
	jand g1322(.dina(w_in363_0[1]),.dinb(w_n1963_0[1]),.dout(n1964),.clk(gclk));
	jnot g1323(.din(w_in261_0[1]),.dout(n1965),.clk(gclk));
	jand g1324(.dina(w_in361_0[1]),.dinb(w_n1965_0[1]),.dout(n1966),.clk(gclk));
	jnot g1325(.din(w_in262_0[1]),.dout(n1967),.clk(gclk));
	jand g1326(.dina(w_in362_0[1]),.dinb(w_n1967_0[1]),.dout(n1968),.clk(gclk));
	jor g1327(.dina(n1968),.dinb(n1966),.dout(n1969),.clk(gclk));
	jor g1328(.dina(n1969),.dinb(w_n1964_0[1]),.dout(n1970),.clk(gclk));
	jor g1329(.dina(w_n1970_0[1]),.dinb(n1962),.dout(n1971),.clk(gclk));
	jnot g1330(.din(w_n1971_0[1]),.dout(n1972),.clk(gclk));
	jand g1331(.dina(n1972),.dinb(w_in259_0[1]),.dout(n1973),.clk(gclk));
	jand g1332(.dina(n1973),.dinb(w_n1960_0[1]),.dout(n1974),.clk(gclk));
	jnot g1333(.din(w_n1974_0[1]),.dout(n1975),.clk(gclk));
	jnot g1334(.din(w_in351_0[1]),.dout(n1976),.clk(gclk));
	jnot g1335(.din(w_in253_0[1]),.dout(n1977),.clk(gclk));
	jand g1336(.dina(w_in353_0[1]),.dinb(w_n1977_0[1]),.dout(n1978),.clk(gclk));
	jnot g1337(.din(w_in255_0[1]),.dout(n1979),.clk(gclk));
	jand g1338(.dina(w_in355_0[1]),.dinb(w_n1979_0[1]),.dout(n1980),.clk(gclk));
	jnot g1339(.din(w_in254_0[1]),.dout(n1981),.clk(gclk));
	jand g1340(.dina(w_in354_0[1]),.dinb(w_n1981_0[1]),.dout(n1982),.clk(gclk));
	jor g1341(.dina(n1982),.dinb(n1980),.dout(n1983),.clk(gclk));
	jnot g1342(.din(w_in252_0[1]),.dout(n1984),.clk(gclk));
	jand g1343(.dina(w_in352_0[1]),.dinb(w_n1984_0[1]),.dout(n1985),.clk(gclk));
	jor g1344(.dina(n1985),.dinb(w_n1983_0[1]),.dout(n1986),.clk(gclk));
	jor g1345(.dina(n1986),.dinb(w_n1978_0[1]),.dout(n1987),.clk(gclk));
	jnot g1346(.din(w_n1987_0[1]),.dout(n1988),.clk(gclk));
	jand g1347(.dina(n1988),.dinb(w_in251_0[1]),.dout(n1989),.clk(gclk));
	jand g1348(.dina(n1989),.dinb(w_n1976_0[1]),.dout(n1990),.clk(gclk));
	jnot g1349(.din(w_n1990_0[1]),.dout(n1991),.clk(gclk));
	jnot g1350(.din(w_in343_0[1]),.dout(n1992),.clk(gclk));
	jnot g1351(.din(w_in244_0[1]),.dout(n1993),.clk(gclk));
	jand g1352(.dina(w_in344_0[1]),.dinb(w_n1993_0[1]),.dout(n1994),.clk(gclk));
	jnot g1353(.din(w_in247_0[1]),.dout(n1995),.clk(gclk));
	jand g1354(.dina(w_in347_0[1]),.dinb(w_n1995_0[1]),.dout(n1996),.clk(gclk));
	jnot g1355(.din(w_in245_0[1]),.dout(n1997),.clk(gclk));
	jand g1356(.dina(w_in345_0[1]),.dinb(w_n1997_0[1]),.dout(n1998),.clk(gclk));
	jnot g1357(.din(w_in246_0[1]),.dout(n1999),.clk(gclk));
	jand g1358(.dina(w_in346_0[1]),.dinb(w_n1999_0[1]),.dout(n2000),.clk(gclk));
	jor g1359(.dina(n2000),.dinb(n1998),.dout(n2001),.clk(gclk));
	jor g1360(.dina(n2001),.dinb(w_n1996_0[1]),.dout(n2002),.clk(gclk));
	jor g1361(.dina(w_n2002_0[1]),.dinb(n1994),.dout(n2003),.clk(gclk));
	jnot g1362(.din(w_n2003_0[1]),.dout(n2004),.clk(gclk));
	jand g1363(.dina(n2004),.dinb(w_in243_0[1]),.dout(n2005),.clk(gclk));
	jand g1364(.dina(n2005),.dinb(w_n1992_0[1]),.dout(n2006),.clk(gclk));
	jnot g1365(.din(w_n2006_0[1]),.dout(n2007),.clk(gclk));
	jnot g1366(.din(w_in333_0[1]),.dout(n2008),.clk(gclk));
	jand g1367(.dina(w_n2008_0[1]),.dinb(w_in233_0[1]),.dout(n2009),.clk(gclk));
	jnot g1368(.din(w_in334_0[1]),.dout(n2010),.clk(gclk));
	jand g1369(.dina(w_n2010_0[1]),.dinb(w_in234_0[1]),.dout(n2011),.clk(gclk));
	jor g1370(.dina(n2011),.dinb(n2009),.dout(n2012),.clk(gclk));
	jnot g1371(.din(w_in233_0[0]),.dout(n2013),.clk(gclk));
	jand g1372(.dina(w_in333_0[0]),.dinb(w_n2013_0[1]),.dout(n2014),.clk(gclk));
	jnot g1373(.din(w_n2014_0[1]),.dout(n2015),.clk(gclk));
	jnot g1374(.din(w_in332_0[1]),.dout(n2016),.clk(gclk));
	jand g1375(.dina(w_n2016_0[1]),.dinb(w_in232_0[1]),.dout(n2017),.clk(gclk));
	jand g1376(.dina(n2017),.dinb(n2015),.dout(n2018),.clk(gclk));
	jor g1377(.dina(n2018),.dinb(n2012),.dout(n2019),.clk(gclk));
	jnot g1378(.din(w_in235_0[1]),.dout(n2020),.clk(gclk));
	jand g1379(.dina(w_in335_0[1]),.dinb(w_n2020_0[1]),.dout(n2021),.clk(gclk));
	jnot g1380(.din(w_in234_0[0]),.dout(n2022),.clk(gclk));
	jand g1381(.dina(w_in334_0[0]),.dinb(w_n2022_0[1]),.dout(n2023),.clk(gclk));
	jor g1382(.dina(n2023),.dinb(n2021),.dout(n2024),.clk(gclk));
	jnot g1383(.din(w_in236_0[1]),.dout(n2025),.clk(gclk));
	jand g1384(.dina(w_in336_0[1]),.dinb(w_n2025_0[1]),.dout(n2026),.clk(gclk));
	jnot g1385(.din(w_in238_0[1]),.dout(n2027),.clk(gclk));
	jand g1386(.dina(w_in338_0[1]),.dinb(w_n2027_0[1]),.dout(n2028),.clk(gclk));
	jnot g1387(.din(w_in239_0[1]),.dout(n2029),.clk(gclk));
	jand g1388(.dina(w_in339_0[1]),.dinb(w_n2029_0[1]),.dout(n2030),.clk(gclk));
	jnot g1389(.din(w_in237_0[1]),.dout(n2031),.clk(gclk));
	jand g1390(.dina(w_in337_0[1]),.dinb(w_n2031_0[1]),.dout(n2032),.clk(gclk));
	jor g1391(.dina(n2032),.dinb(w_n2030_0[1]),.dout(n2033),.clk(gclk));
	jor g1392(.dina(n2033),.dinb(n2028),.dout(n2034),.clk(gclk));
	jor g1393(.dina(w_n2034_0[1]),.dinb(n2026),.dout(n2035),.clk(gclk));
	jor g1394(.dina(w_n2035_0[1]),.dinb(n2024),.dout(n2036),.clk(gclk));
	jnot g1395(.din(w_n2036_0[1]),.dout(n2037),.clk(gclk));
	jand g1396(.dina(n2037),.dinb(n2019),.dout(n2038),.clk(gclk));
	jnot g1397(.din(w_n2038_0[1]),.dout(n2039),.clk(gclk));
	jnot g1398(.din(w_in230_0[1]),.dout(n2040),.clk(gclk));
	jand g1399(.dina(w_in330_0[1]),.dinb(w_n2040_0[1]),.dout(n2041),.clk(gclk));
	jnot g1400(.din(w_in329_0[1]),.dout(n2042),.clk(gclk));
	jand g1401(.dina(w_n2042_0[1]),.dinb(w_in229_0[1]),.dout(n2043),.clk(gclk));
	jnot g1402(.din(w_n2043_0[1]),.dout(n2044),.clk(gclk));
	jnot g1403(.din(w_in229_0[0]),.dout(n2045),.clk(gclk));
	jand g1404(.dina(w_in329_0[0]),.dinb(w_n2045_0[1]),.dout(n2046),.clk(gclk));
	jnot g1405(.din(w_in328_0[1]),.dout(n2047),.clk(gclk));
	jand g1406(.dina(w_n2047_0[1]),.dinb(w_in228_0[1]),.dout(n2048),.clk(gclk));
	jnot g1407(.din(w_n2048_0[1]),.dout(n2049),.clk(gclk));
	jnot g1408(.din(w_in228_0[0]),.dout(n2050),.clk(gclk));
	jand g1409(.dina(w_in328_0[0]),.dinb(w_n2050_0[1]),.dout(n2051),.clk(gclk));
	jnot g1410(.din(w_in327_0[1]),.dout(n2052),.clk(gclk));
	jand g1411(.dina(w_n2052_0[1]),.dinb(w_in227_0[1]),.dout(n2053),.clk(gclk));
	jnot g1412(.din(w_n2053_0[1]),.dout(n2054),.clk(gclk));
	jnot g1413(.din(w_in227_0[0]),.dout(n2055),.clk(gclk));
	jand g1414(.dina(w_in327_0[0]),.dinb(w_n2055_0[1]),.dout(n2056),.clk(gclk));
	jnot g1415(.din(w_in326_0[1]),.dout(n2057),.clk(gclk));
	jand g1416(.dina(w_n2057_0[1]),.dinb(w_in226_0[1]),.dout(n2058),.clk(gclk));
	jnot g1417(.din(w_n2058_0[1]),.dout(n2059),.clk(gclk));
	jnot g1418(.din(w_in223_0[1]),.dout(n2060),.clk(gclk));
	jand g1419(.dina(w_in323_0[1]),.dinb(w_n2060_0[1]),.dout(n2061),.clk(gclk));
	jnot g1420(.din(w_in222_0[1]),.dout(n2062),.clk(gclk));
	jand g1421(.dina(w_in322_0[1]),.dinb(w_n2062_0[1]),.dout(n2063),.clk(gclk));
	jnot g1422(.din(w_in321_0[1]),.dout(n2064),.clk(gclk));
	jand g1423(.dina(w_n2064_0[1]),.dinb(w_in221_0[1]),.dout(n2065),.clk(gclk));
	jnot g1424(.din(w_n2065_0[1]),.dout(n2066),.clk(gclk));
	jnot g1425(.din(w_in221_0[0]),.dout(n2067),.clk(gclk));
	jand g1426(.dina(w_in321_0[0]),.dinb(w_n2067_0[1]),.dout(n2068),.clk(gclk));
	jnot g1427(.din(w_in320_0[1]),.dout(n2069),.clk(gclk));
	jand g1428(.dina(w_n2069_0[1]),.dinb(w_in220_0[1]),.dout(n2070),.clk(gclk));
	jnot g1429(.din(w_n2070_0[1]),.dout(n2071),.clk(gclk));
	jnot g1430(.din(w_in220_0[0]),.dout(n2072),.clk(gclk));
	jand g1431(.dina(w_in320_0[0]),.dinb(w_n2072_0[1]),.dout(n2073),.clk(gclk));
	jnot g1432(.din(w_in319_0[1]),.dout(n2074),.clk(gclk));
	jand g1433(.dina(w_n2074_0[1]),.dinb(w_in219_0[1]),.dout(n2075),.clk(gclk));
	jnot g1434(.din(w_n2075_0[1]),.dout(n2076),.clk(gclk));
	jnot g1435(.din(w_in219_0[0]),.dout(n2077),.clk(gclk));
	jand g1436(.dina(w_in319_0[0]),.dinb(w_n2077_0[1]),.dout(n2078),.clk(gclk));
	jnot g1437(.din(w_in318_0[1]),.dout(n2079),.clk(gclk));
	jand g1438(.dina(w_n2079_0[1]),.dinb(w_in218_0[1]),.dout(n2080),.clk(gclk));
	jnot g1439(.din(w_n2080_0[1]),.dout(n2081),.clk(gclk));
	jnot g1440(.din(w_in215_0[1]),.dout(n2082),.clk(gclk));
	jand g1441(.dina(w_in315_0[1]),.dinb(w_n2082_0[1]),.dout(n2083),.clk(gclk));
	jnot g1442(.din(w_in214_0[1]),.dout(n2084),.clk(gclk));
	jand g1443(.dina(w_in314_0[1]),.dinb(w_n2084_0[1]),.dout(n2085),.clk(gclk));
	jnot g1444(.din(w_in313_0[1]),.dout(n2086),.clk(gclk));
	jand g1445(.dina(w_n2086_0[1]),.dinb(w_in213_0[1]),.dout(n2087),.clk(gclk));
	jnot g1446(.din(w_n2087_0[1]),.dout(n2088),.clk(gclk));
	jnot g1447(.din(w_in213_0[0]),.dout(n2089),.clk(gclk));
	jand g1448(.dina(w_in313_0[0]),.dinb(w_n2089_0[1]),.dout(n2090),.clk(gclk));
	jnot g1449(.din(w_in312_0[1]),.dout(n2091),.clk(gclk));
	jand g1450(.dina(w_n2091_0[1]),.dinb(w_in212_0[1]),.dout(n2092),.clk(gclk));
	jnot g1451(.din(w_n2092_0[1]),.dout(n2093),.clk(gclk));
	jnot g1452(.din(w_in212_0[0]),.dout(n2094),.clk(gclk));
	jand g1453(.dina(w_in312_0[0]),.dinb(w_n2094_0[1]),.dout(n2095),.clk(gclk));
	jnot g1454(.din(w_in311_0[1]),.dout(n2096),.clk(gclk));
	jand g1455(.dina(w_n2096_0[1]),.dinb(w_in211_0[1]),.dout(n2097),.clk(gclk));
	jnot g1456(.din(w_n2097_0[1]),.dout(n2098),.clk(gclk));
	jnot g1457(.din(w_in211_0[0]),.dout(n2099),.clk(gclk));
	jand g1458(.dina(w_in311_0[0]),.dinb(w_n2099_0[1]),.dout(n2100),.clk(gclk));
	jnot g1459(.din(w_in310_0[1]),.dout(n2101),.clk(gclk));
	jand g1460(.dina(w_n2101_0[1]),.dinb(w_in210_0[1]),.dout(n2102),.clk(gclk));
	jnot g1461(.din(w_n2102_0[1]),.dout(n2103),.clk(gclk));
	jnot g1462(.din(w_in27_0[1]),.dout(n2104),.clk(gclk));
	jand g1463(.dina(w_in37_0[1]),.dinb(w_n2104_0[1]),.dout(n2105),.clk(gclk));
	jnot g1464(.din(w_in23_0[1]),.dout(n2106),.clk(gclk));
	jand g1465(.dina(w_in33_0[1]),.dinb(w_n2106_0[1]),.dout(n2107),.clk(gclk));
	jnot g1466(.din(w_in22_0[2]),.dout(n2108),.clk(gclk));
	jand g1467(.dina(w_in32_0[2]),.dinb(w_n2108_0[1]),.dout(n2109),.clk(gclk));
	jnot g1468(.din(w_in31_0[2]),.dout(n2110),.clk(gclk));
	jand g1469(.dina(w_n2110_0[2]),.dinb(w_in21_1[1]),.dout(n2111),.clk(gclk));
	jnot g1470(.din(w_n2111_0[1]),.dout(n2112),.clk(gclk));
	jnot g1471(.din(w_in21_1[0]),.dout(n2113),.clk(gclk));
	jand g1472(.dina(w_in31_0[1]),.dinb(w_n2113_0[1]),.dout(n2114),.clk(gclk));
	jnot g1473(.din(w_in20_0[2]),.dout(n2115),.clk(gclk));
	jor g1474(.dina(w_in30_0[2]),.dinb(w_n2115_0[1]),.dout(n2116),.clk(gclk));
	jor g1475(.dina(n2116),.dinb(n2114),.dout(n2117),.clk(gclk));
	jand g1476(.dina(n2117),.dinb(n2112),.dout(n2118),.clk(gclk));
	jor g1477(.dina(n2118),.dinb(w_n2109_0[1]),.dout(n2119),.clk(gclk));
	jnot g1478(.din(w_in33_0[0]),.dout(n2120),.clk(gclk));
	jand g1479(.dina(w_n2120_0[1]),.dinb(w_in23_0[0]),.dout(n2121),.clk(gclk));
	jnot g1480(.din(w_in32_0[1]),.dout(n2122),.clk(gclk));
	jand g1481(.dina(w_n2122_0[1]),.dinb(w_in22_0[1]),.dout(n2123),.clk(gclk));
	jor g1482(.dina(n2123),.dinb(n2121),.dout(n2124),.clk(gclk));
	jnot g1483(.din(w_n2124_0[1]),.dout(n2125),.clk(gclk));
	jand g1484(.dina(n2125),.dinb(n2119),.dout(n2126),.clk(gclk));
	jnot g1485(.din(w_in24_0[1]),.dout(n2127),.clk(gclk));
	jand g1486(.dina(w_in34_0[1]),.dinb(w_n2127_0[1]),.dout(n2128),.clk(gclk));
	jor g1487(.dina(w_n2128_0[1]),.dinb(n2126),.dout(n2129),.clk(gclk));
	jor g1488(.dina(n2129),.dinb(w_n2107_0[1]),.dout(n2130),.clk(gclk));
	jnot g1489(.din(w_in34_0[0]),.dout(n2131),.clk(gclk));
	jand g1490(.dina(w_n2131_0[1]),.dinb(w_in24_0[0]),.dout(n2132),.clk(gclk));
	jnot g1491(.din(w_in35_0[1]),.dout(n2133),.clk(gclk));
	jand g1492(.dina(w_n2133_0[1]),.dinb(w_in25_0[1]),.dout(n2134),.clk(gclk));
	jor g1493(.dina(n2134),.dinb(n2132),.dout(n2135),.clk(gclk));
	jnot g1494(.din(w_n2135_0[1]),.dout(n2136),.clk(gclk));
	jand g1495(.dina(n2136),.dinb(n2130),.dout(n2137),.clk(gclk));
	jnot g1496(.din(w_in26_0[1]),.dout(n2138),.clk(gclk));
	jand g1497(.dina(w_in36_0[1]),.dinb(w_n2138_0[1]),.dout(n2139),.clk(gclk));
	jnot g1498(.din(w_in25_0[0]),.dout(n2140),.clk(gclk));
	jand g1499(.dina(w_in35_0[0]),.dinb(w_n2140_0[1]),.dout(n2141),.clk(gclk));
	jor g1500(.dina(n2141),.dinb(n2139),.dout(n2142),.clk(gclk));
	jor g1501(.dina(w_n2142_0[1]),.dinb(n2137),.dout(n2143),.clk(gclk));
	jnot g1502(.din(w_in37_0[0]),.dout(n2144),.clk(gclk));
	jand g1503(.dina(w_n2144_0[1]),.dinb(w_in27_0[0]),.dout(n2145),.clk(gclk));
	jnot g1504(.din(w_in36_0[0]),.dout(n2146),.clk(gclk));
	jand g1505(.dina(w_n2146_0[1]),.dinb(w_in26_0[0]),.dout(n2147),.clk(gclk));
	jor g1506(.dina(n2147),.dinb(n2145),.dout(n2148),.clk(gclk));
	jnot g1507(.din(w_n2148_0[1]),.dout(n2149),.clk(gclk));
	jand g1508(.dina(n2149),.dinb(n2143),.dout(n2150),.clk(gclk));
	jnot g1509(.din(w_in28_0[1]),.dout(n2151),.clk(gclk));
	jand g1510(.dina(w_in38_0[1]),.dinb(w_n2151_0[1]),.dout(n2152),.clk(gclk));
	jor g1511(.dina(w_n2152_0[1]),.dinb(n2150),.dout(n2153),.clk(gclk));
	jor g1512(.dina(n2153),.dinb(w_n2105_0[1]),.dout(n2154),.clk(gclk));
	jnot g1513(.din(w_in38_0[0]),.dout(n2155),.clk(gclk));
	jand g1514(.dina(w_n2155_0[1]),.dinb(w_in28_0[0]),.dout(n2156),.clk(gclk));
	jnot g1515(.din(w_in39_0[1]),.dout(n2157),.clk(gclk));
	jand g1516(.dina(w_n2157_0[1]),.dinb(w_in29_0[1]),.dout(n2158),.clk(gclk));
	jor g1517(.dina(n2158),.dinb(n2156),.dout(n2159),.clk(gclk));
	jnot g1518(.din(w_n2159_0[1]),.dout(n2160),.clk(gclk));
	jand g1519(.dina(n2160),.dinb(n2154),.dout(n2161),.clk(gclk));
	jnot g1520(.din(w_in210_0[0]),.dout(n2162),.clk(gclk));
	jand g1521(.dina(w_in310_0[0]),.dinb(w_n2162_0[1]),.dout(n2163),.clk(gclk));
	jnot g1522(.din(w_in29_0[0]),.dout(n2164),.clk(gclk));
	jand g1523(.dina(w_in39_0[0]),.dinb(w_n2164_0[1]),.dout(n2165),.clk(gclk));
	jor g1524(.dina(n2165),.dinb(n2163),.dout(n2166),.clk(gclk));
	jor g1525(.dina(w_n2166_0[1]),.dinb(n2161),.dout(n2167),.clk(gclk));
	jand g1526(.dina(n2167),.dinb(n2103),.dout(n2168),.clk(gclk));
	jor g1527(.dina(n2168),.dinb(w_n2100_0[1]),.dout(n2169),.clk(gclk));
	jand g1528(.dina(n2169),.dinb(n2098),.dout(n2170),.clk(gclk));
	jor g1529(.dina(n2170),.dinb(w_n2095_0[1]),.dout(n2171),.clk(gclk));
	jand g1530(.dina(n2171),.dinb(n2093),.dout(n2172),.clk(gclk));
	jor g1531(.dina(n2172),.dinb(w_n2090_0[1]),.dout(n2173),.clk(gclk));
	jand g1532(.dina(n2173),.dinb(n2088),.dout(n2174),.clk(gclk));
	jor g1533(.dina(n2174),.dinb(w_n2085_0[1]),.dout(n2175),.clk(gclk));
	jnot g1534(.din(w_in315_0[0]),.dout(n2176),.clk(gclk));
	jand g1535(.dina(w_n2176_0[1]),.dinb(w_in215_0[0]),.dout(n2177),.clk(gclk));
	jnot g1536(.din(w_in314_0[0]),.dout(n2178),.clk(gclk));
	jand g1537(.dina(w_n2178_0[1]),.dinb(w_in214_0[0]),.dout(n2179),.clk(gclk));
	jor g1538(.dina(n2179),.dinb(n2177),.dout(n2180),.clk(gclk));
	jnot g1539(.din(w_n2180_0[1]),.dout(n2181),.clk(gclk));
	jand g1540(.dina(n2181),.dinb(n2175),.dout(n2182),.clk(gclk));
	jnot g1541(.din(w_in216_0[1]),.dout(n2183),.clk(gclk));
	jand g1542(.dina(w_in316_0[1]),.dinb(w_n2183_0[1]),.dout(n2184),.clk(gclk));
	jor g1543(.dina(w_n2184_0[1]),.dinb(n2182),.dout(n2185),.clk(gclk));
	jor g1544(.dina(n2185),.dinb(w_n2083_0[1]),.dout(n2186),.clk(gclk));
	jnot g1545(.din(w_in316_0[0]),.dout(n2187),.clk(gclk));
	jand g1546(.dina(w_n2187_0[1]),.dinb(w_in216_0[0]),.dout(n2188),.clk(gclk));
	jnot g1547(.din(w_in317_0[1]),.dout(n2189),.clk(gclk));
	jand g1548(.dina(w_n2189_0[1]),.dinb(w_in217_0[1]),.dout(n2190),.clk(gclk));
	jor g1549(.dina(n2190),.dinb(n2188),.dout(n2191),.clk(gclk));
	jnot g1550(.din(w_n2191_0[1]),.dout(n2192),.clk(gclk));
	jand g1551(.dina(n2192),.dinb(n2186),.dout(n2193),.clk(gclk));
	jnot g1552(.din(w_in218_0[0]),.dout(n2194),.clk(gclk));
	jand g1553(.dina(w_in318_0[0]),.dinb(w_n2194_0[1]),.dout(n2195),.clk(gclk));
	jnot g1554(.din(w_in217_0[0]),.dout(n2196),.clk(gclk));
	jand g1555(.dina(w_in317_0[0]),.dinb(w_n2196_0[1]),.dout(n2197),.clk(gclk));
	jor g1556(.dina(n2197),.dinb(n2195),.dout(n2198),.clk(gclk));
	jor g1557(.dina(w_n2198_0[1]),.dinb(n2193),.dout(n2199),.clk(gclk));
	jand g1558(.dina(n2199),.dinb(n2081),.dout(n2200),.clk(gclk));
	jor g1559(.dina(n2200),.dinb(w_n2078_0[1]),.dout(n2201),.clk(gclk));
	jand g1560(.dina(n2201),.dinb(n2076),.dout(n2202),.clk(gclk));
	jor g1561(.dina(n2202),.dinb(w_n2073_0[1]),.dout(n2203),.clk(gclk));
	jand g1562(.dina(n2203),.dinb(n2071),.dout(n2204),.clk(gclk));
	jor g1563(.dina(n2204),.dinb(w_n2068_0[1]),.dout(n2205),.clk(gclk));
	jand g1564(.dina(n2205),.dinb(n2066),.dout(n2206),.clk(gclk));
	jor g1565(.dina(n2206),.dinb(w_n2063_0[1]),.dout(n2207),.clk(gclk));
	jnot g1566(.din(w_in323_0[0]),.dout(n2208),.clk(gclk));
	jand g1567(.dina(w_n2208_0[1]),.dinb(w_in223_0[0]),.dout(n2209),.clk(gclk));
	jnot g1568(.din(w_in322_0[0]),.dout(n2210),.clk(gclk));
	jand g1569(.dina(w_n2210_0[1]),.dinb(w_in222_0[0]),.dout(n2211),.clk(gclk));
	jor g1570(.dina(n2211),.dinb(n2209),.dout(n2212),.clk(gclk));
	jnot g1571(.din(w_n2212_0[1]),.dout(n2213),.clk(gclk));
	jand g1572(.dina(n2213),.dinb(n2207),.dout(n2214),.clk(gclk));
	jnot g1573(.din(w_in224_0[1]),.dout(n2215),.clk(gclk));
	jand g1574(.dina(w_in324_0[1]),.dinb(w_n2215_0[1]),.dout(n2216),.clk(gclk));
	jor g1575(.dina(w_n2216_0[1]),.dinb(n2214),.dout(n2217),.clk(gclk));
	jor g1576(.dina(n2217),.dinb(w_n2061_0[1]),.dout(n2218),.clk(gclk));
	jnot g1577(.din(w_in324_0[0]),.dout(n2219),.clk(gclk));
	jand g1578(.dina(w_n2219_0[1]),.dinb(w_in224_0[0]),.dout(n2220),.clk(gclk));
	jnot g1579(.din(w_in325_0[1]),.dout(n2221),.clk(gclk));
	jand g1580(.dina(w_n2221_0[1]),.dinb(w_in225_0[1]),.dout(n2222),.clk(gclk));
	jor g1581(.dina(n2222),.dinb(n2220),.dout(n2223),.clk(gclk));
	jnot g1582(.din(w_n2223_0[1]),.dout(n2224),.clk(gclk));
	jand g1583(.dina(n2224),.dinb(n2218),.dout(n2225),.clk(gclk));
	jnot g1584(.din(w_in226_0[0]),.dout(n2226),.clk(gclk));
	jand g1585(.dina(w_in326_0[0]),.dinb(w_n2226_0[1]),.dout(n2227),.clk(gclk));
	jnot g1586(.din(w_in225_0[0]),.dout(n2228),.clk(gclk));
	jand g1587(.dina(w_in325_0[0]),.dinb(w_n2228_0[1]),.dout(n2229),.clk(gclk));
	jor g1588(.dina(n2229),.dinb(n2227),.dout(n2230),.clk(gclk));
	jor g1589(.dina(w_n2230_0[1]),.dinb(n2225),.dout(n2231),.clk(gclk));
	jand g1590(.dina(n2231),.dinb(n2059),.dout(n2232),.clk(gclk));
	jor g1591(.dina(n2232),.dinb(w_n2056_0[1]),.dout(n2233),.clk(gclk));
	jand g1592(.dina(n2233),.dinb(n2054),.dout(n2234),.clk(gclk));
	jor g1593(.dina(n2234),.dinb(w_n2051_0[1]),.dout(n2235),.clk(gclk));
	jand g1594(.dina(n2235),.dinb(n2049),.dout(n2236),.clk(gclk));
	jor g1595(.dina(n2236),.dinb(w_n2046_0[1]),.dout(n2237),.clk(gclk));
	jand g1596(.dina(n2237),.dinb(n2044),.dout(n2238),.clk(gclk));
	jor g1597(.dina(n2238),.dinb(w_n2041_0[1]),.dout(n2239),.clk(gclk));
	jnot g1598(.din(w_in331_0[1]),.dout(n2240),.clk(gclk));
	jand g1599(.dina(w_n2240_0[1]),.dinb(w_in231_0[1]),.dout(n2241),.clk(gclk));
	jnot g1600(.din(w_in330_0[0]),.dout(n2242),.clk(gclk));
	jand g1601(.dina(w_n2242_0[1]),.dinb(w_in230_0[0]),.dout(n2243),.clk(gclk));
	jor g1602(.dina(n2243),.dinb(n2241),.dout(n2244),.clk(gclk));
	jnot g1603(.din(w_n2244_0[1]),.dout(n2245),.clk(gclk));
	jand g1604(.dina(n2245),.dinb(n2239),.dout(n2246),.clk(gclk));
	jnot g1605(.din(w_in231_0[0]),.dout(n2247),.clk(gclk));
	jand g1606(.dina(w_in331_0[0]),.dinb(w_n2247_0[1]),.dout(n2248),.clk(gclk));
	jnot g1607(.din(w_in232_0[0]),.dout(n2249),.clk(gclk));
	jand g1608(.dina(w_in332_0[0]),.dinb(w_n2249_0[1]),.dout(n2250),.clk(gclk));
	jor g1609(.dina(n2250),.dinb(n2248),.dout(n2251),.clk(gclk));
	jor g1610(.dina(n2251),.dinb(w_n2014_0[0]),.dout(n2252),.clk(gclk));
	jor g1611(.dina(n2252),.dinb(w_n2036_0[0]),.dout(n2253),.clk(gclk));
	jor g1612(.dina(w_n2253_0[1]),.dinb(n2246),.dout(n2254),.clk(gclk));
	jnot g1613(.din(w_n2034_0[0]),.dout(n2255),.clk(gclk));
	jnot g1614(.din(w_in337_0[0]),.dout(n2256),.clk(gclk));
	jand g1615(.dina(w_n2256_0[1]),.dinb(w_in237_0[0]),.dout(n2257),.clk(gclk));
	jnot g1616(.din(w_in336_0[0]),.dout(n2258),.clk(gclk));
	jand g1617(.dina(w_n2258_0[1]),.dinb(w_in236_0[0]),.dout(n2259),.clk(gclk));
	jor g1618(.dina(n2259),.dinb(n2257),.dout(n2260),.clk(gclk));
	jand g1619(.dina(n2260),.dinb(n2255),.dout(n2261),.clk(gclk));
	jnot g1620(.din(w_n2035_0[0]),.dout(n2262),.clk(gclk));
	jnot g1621(.din(w_in335_0[0]),.dout(n2263),.clk(gclk));
	jand g1622(.dina(w_n2263_0[1]),.dinb(w_in235_0[0]),.dout(n2264),.clk(gclk));
	jand g1623(.dina(n2264),.dinb(n2262),.dout(n2265),.clk(gclk));
	jnot g1624(.din(w_in339_0[0]),.dout(n2266),.clk(gclk));
	jand g1625(.dina(w_n2266_0[1]),.dinb(w_in239_0[0]),.dout(n2267),.clk(gclk));
	jnot g1626(.din(w_n2030_0[0]),.dout(n2268),.clk(gclk));
	jnot g1627(.din(w_in338_0[0]),.dout(n2269),.clk(gclk));
	jand g1628(.dina(w_n2269_0[1]),.dinb(w_in238_0[0]),.dout(n2270),.clk(gclk));
	jand g1629(.dina(n2270),.dinb(n2268),.dout(n2271),.clk(gclk));
	jor g1630(.dina(n2271),.dinb(n2267),.dout(n2272),.clk(gclk));
	jor g1631(.dina(n2272),.dinb(n2265),.dout(n2273),.clk(gclk));
	jor g1632(.dina(n2273),.dinb(n2261),.dout(n2274),.clk(gclk));
	jnot g1633(.din(w_n2274_0[1]),.dout(n2275),.clk(gclk));
	jand g1634(.dina(n2275),.dinb(n2254),.dout(n2276),.clk(gclk));
	jand g1635(.dina(n2276),.dinb(n2039),.dout(n2277),.clk(gclk));
	jnot g1636(.din(w_in240_0[1]),.dout(n2278),.clk(gclk));
	jand g1637(.dina(w_in340_0[1]),.dinb(w_n2278_0[1]),.dout(n2279),.clk(gclk));
	jnot g1638(.din(n2279),.dout(n2280),.clk(gclk));
	jnot g1639(.din(w_in241_0[1]),.dout(n2281),.clk(gclk));
	jand g1640(.dina(w_in341_0[1]),.dinb(w_n2281_0[1]),.dout(n2282),.clk(gclk));
	jnot g1641(.din(n2282),.dout(n2283),.clk(gclk));
	jnot g1642(.din(w_in242_0[1]),.dout(n2284),.clk(gclk));
	jand g1643(.dina(w_in342_0[1]),.dinb(w_n2284_0[1]),.dout(n2285),.clk(gclk));
	jnot g1644(.din(w_in243_0[0]),.dout(n2286),.clk(gclk));
	jand g1645(.dina(w_in343_0[0]),.dinb(w_n2286_0[1]),.dout(n2287),.clk(gclk));
	jor g1646(.dina(n2287),.dinb(n2285),.dout(n2288),.clk(gclk));
	jor g1647(.dina(n2288),.dinb(w_n2003_0[0]),.dout(n2289),.clk(gclk));
	jnot g1648(.din(n2289),.dout(n2290),.clk(gclk));
	jand g1649(.dina(w_n2290_0[1]),.dinb(w_n2283_0[1]),.dout(n2291),.clk(gclk));
	jand g1650(.dina(n2291),.dinb(n2280),.dout(n2292),.clk(gclk));
	jnot g1651(.din(w_n2292_0[1]),.dout(n2293),.clk(gclk));
	jor g1652(.dina(n2293),.dinb(n2277),.dout(n2294),.clk(gclk));
	jnot g1653(.din(w_in341_0[0]),.dout(n2295),.clk(gclk));
	jand g1654(.dina(w_n2295_0[1]),.dinb(w_in241_0[0]),.dout(n2296),.clk(gclk));
	jnot g1655(.din(w_in342_0[0]),.dout(n2297),.clk(gclk));
	jand g1656(.dina(w_n2297_0[1]),.dinb(w_in242_0[0]),.dout(n2298),.clk(gclk));
	jor g1657(.dina(n2298),.dinb(n2296),.dout(n2299),.clk(gclk));
	jnot g1658(.din(w_in340_0[0]),.dout(n2300),.clk(gclk));
	jand g1659(.dina(w_n2300_0[1]),.dinb(w_in240_0[0]),.dout(n2301),.clk(gclk));
	jand g1660(.dina(n2301),.dinb(w_n2283_0[0]),.dout(n2302),.clk(gclk));
	jor g1661(.dina(n2302),.dinb(n2299),.dout(n2303),.clk(gclk));
	jand g1662(.dina(n2303),.dinb(w_n2290_0[0]),.dout(n2304),.clk(gclk));
	jnot g1663(.din(w_n2002_0[0]),.dout(n2305),.clk(gclk));
	jnot g1664(.din(w_in345_0[0]),.dout(n2306),.clk(gclk));
	jand g1665(.dina(w_n2306_0[1]),.dinb(w_in245_0[0]),.dout(n2307),.clk(gclk));
	jnot g1666(.din(w_in344_0[0]),.dout(n2308),.clk(gclk));
	jand g1667(.dina(w_n2308_0[1]),.dinb(w_in244_0[0]),.dout(n2309),.clk(gclk));
	jor g1668(.dina(n2309),.dinb(n2307),.dout(n2310),.clk(gclk));
	jand g1669(.dina(n2310),.dinb(n2305),.dout(n2311),.clk(gclk));
	jnot g1670(.din(w_n1996_0[0]),.dout(n2312),.clk(gclk));
	jnot g1671(.din(w_in347_0[0]),.dout(n2313),.clk(gclk));
	jand g1672(.dina(w_n2313_0[1]),.dinb(w_in247_0[0]),.dout(n2314),.clk(gclk));
	jnot g1673(.din(w_in346_0[0]),.dout(n2315),.clk(gclk));
	jand g1674(.dina(w_n2315_0[1]),.dinb(w_in246_0[0]),.dout(n2316),.clk(gclk));
	jor g1675(.dina(n2316),.dinb(n2314),.dout(n2317),.clk(gclk));
	jand g1676(.dina(n2317),.dinb(n2312),.dout(n2318),.clk(gclk));
	jor g1677(.dina(n2318),.dinb(n2311),.dout(n2319),.clk(gclk));
	jor g1678(.dina(n2319),.dinb(n2304),.dout(n2320),.clk(gclk));
	jnot g1679(.din(w_n2320_0[1]),.dout(n2321),.clk(gclk));
	jand g1680(.dina(n2321),.dinb(n2294),.dout(n2322),.clk(gclk));
	jand g1681(.dina(n2322),.dinb(n2007),.dout(n2323),.clk(gclk));
	jnot g1682(.din(w_in248_0[1]),.dout(n2324),.clk(gclk));
	jand g1683(.dina(w_in348_0[1]),.dinb(w_n2324_0[1]),.dout(n2325),.clk(gclk));
	jnot g1684(.din(n2325),.dout(n2326),.clk(gclk));
	jnot g1685(.din(w_in249_0[1]),.dout(n2327),.clk(gclk));
	jand g1686(.dina(w_in349_0[1]),.dinb(w_n2327_0[1]),.dout(n2328),.clk(gclk));
	jnot g1687(.din(n2328),.dout(n2329),.clk(gclk));
	jnot g1688(.din(w_in250_0[1]),.dout(n2330),.clk(gclk));
	jand g1689(.dina(w_in350_0[1]),.dinb(w_n2330_0[1]),.dout(n2331),.clk(gclk));
	jnot g1690(.din(w_in251_0[0]),.dout(n2332),.clk(gclk));
	jand g1691(.dina(w_in351_0[0]),.dinb(w_n2332_0[1]),.dout(n2333),.clk(gclk));
	jor g1692(.dina(n2333),.dinb(n2331),.dout(n2334),.clk(gclk));
	jor g1693(.dina(n2334),.dinb(w_n1987_0[0]),.dout(n2335),.clk(gclk));
	jnot g1694(.din(n2335),.dout(n2336),.clk(gclk));
	jand g1695(.dina(w_n2336_0[1]),.dinb(w_n2329_0[1]),.dout(n2337),.clk(gclk));
	jand g1696(.dina(n2337),.dinb(n2326),.dout(n2338),.clk(gclk));
	jnot g1697(.din(w_n2338_0[1]),.dout(n2339),.clk(gclk));
	jor g1698(.dina(n2339),.dinb(n2323),.dout(n2340),.clk(gclk));
	jnot g1699(.din(w_in349_0[0]),.dout(n2341),.clk(gclk));
	jand g1700(.dina(w_n2341_0[1]),.dinb(w_in249_0[0]),.dout(n2342),.clk(gclk));
	jnot g1701(.din(w_in350_0[0]),.dout(n2343),.clk(gclk));
	jand g1702(.dina(w_n2343_0[1]),.dinb(w_in250_0[0]),.dout(n2344),.clk(gclk));
	jor g1703(.dina(n2344),.dinb(n2342),.dout(n2345),.clk(gclk));
	jnot g1704(.din(w_in348_0[0]),.dout(n2346),.clk(gclk));
	jand g1705(.dina(w_n2346_0[1]),.dinb(w_in248_0[0]),.dout(n2347),.clk(gclk));
	jand g1706(.dina(n2347),.dinb(w_n2329_0[0]),.dout(n2348),.clk(gclk));
	jor g1707(.dina(n2348),.dinb(n2345),.dout(n2349),.clk(gclk));
	jand g1708(.dina(n2349),.dinb(w_n2336_0[0]),.dout(n2350),.clk(gclk));
	jnot g1709(.din(w_in355_0[0]),.dout(n2351),.clk(gclk));
	jand g1710(.dina(w_n2351_0[1]),.dinb(w_in255_0[0]),.dout(n2352),.clk(gclk));
	jnot g1711(.din(w_n1983_0[0]),.dout(n2353),.clk(gclk));
	jnot g1712(.din(w_n1978_0[0]),.dout(n2354),.clk(gclk));
	jnot g1713(.din(w_in352_0[0]),.dout(n2355),.clk(gclk));
	jand g1714(.dina(w_n2355_0[1]),.dinb(w_in252_0[0]),.dout(n2356),.clk(gclk));
	jand g1715(.dina(n2356),.dinb(n2354),.dout(n2357),.clk(gclk));
	jnot g1716(.din(w_in354_0[0]),.dout(n2358),.clk(gclk));
	jand g1717(.dina(w_n2358_0[1]),.dinb(w_in254_0[0]),.dout(n2359),.clk(gclk));
	jnot g1718(.din(w_in353_0[0]),.dout(n2360),.clk(gclk));
	jand g1719(.dina(w_n2360_0[1]),.dinb(w_in253_0[0]),.dout(n2361),.clk(gclk));
	jor g1720(.dina(n2361),.dinb(n2359),.dout(n2362),.clk(gclk));
	jor g1721(.dina(n2362),.dinb(n2357),.dout(n2363),.clk(gclk));
	jand g1722(.dina(n2363),.dinb(n2353),.dout(n2364),.clk(gclk));
	jor g1723(.dina(n2364),.dinb(n2352),.dout(n2365),.clk(gclk));
	jor g1724(.dina(n2365),.dinb(n2350),.dout(n2366),.clk(gclk));
	jnot g1725(.din(w_n2366_0[1]),.dout(n2367),.clk(gclk));
	jand g1726(.dina(n2367),.dinb(n2340),.dout(n2368),.clk(gclk));
	jand g1727(.dina(n2368),.dinb(n1991),.dout(n2369),.clk(gclk));
	jnot g1728(.din(w_in256_0[1]),.dout(n2370),.clk(gclk));
	jand g1729(.dina(w_in356_0[1]),.dinb(w_n2370_0[1]),.dout(n2371),.clk(gclk));
	jnot g1730(.din(n2371),.dout(n2372),.clk(gclk));
	jnot g1731(.din(w_in257_0[1]),.dout(n2373),.clk(gclk));
	jand g1732(.dina(w_in357_0[1]),.dinb(w_n2373_0[1]),.dout(n2374),.clk(gclk));
	jnot g1733(.din(n2374),.dout(n2375),.clk(gclk));
	jnot g1734(.din(w_in258_0[1]),.dout(n2376),.clk(gclk));
	jand g1735(.dina(w_in358_0[1]),.dinb(w_n2376_0[1]),.dout(n2377),.clk(gclk));
	jnot g1736(.din(w_in259_0[0]),.dout(n2378),.clk(gclk));
	jand g1737(.dina(w_in359_0[0]),.dinb(w_n2378_0[1]),.dout(n2379),.clk(gclk));
	jor g1738(.dina(n2379),.dinb(n2377),.dout(n2380),.clk(gclk));
	jor g1739(.dina(n2380),.dinb(w_n1971_0[0]),.dout(n2381),.clk(gclk));
	jnot g1740(.din(n2381),.dout(n2382),.clk(gclk));
	jand g1741(.dina(w_n2382_0[1]),.dinb(w_n2375_0[1]),.dout(n2383),.clk(gclk));
	jand g1742(.dina(n2383),.dinb(n2372),.dout(n2384),.clk(gclk));
	jnot g1743(.din(w_n2384_0[1]),.dout(n2385),.clk(gclk));
	jor g1744(.dina(n2385),.dinb(n2369),.dout(n2386),.clk(gclk));
	jnot g1745(.din(w_in357_0[0]),.dout(n2387),.clk(gclk));
	jand g1746(.dina(w_n2387_0[1]),.dinb(w_in257_0[0]),.dout(n2388),.clk(gclk));
	jnot g1747(.din(w_in358_0[0]),.dout(n2389),.clk(gclk));
	jand g1748(.dina(w_n2389_0[1]),.dinb(w_in258_0[0]),.dout(n2390),.clk(gclk));
	jor g1749(.dina(n2390),.dinb(n2388),.dout(n2391),.clk(gclk));
	jnot g1750(.din(w_in356_0[0]),.dout(n2392),.clk(gclk));
	jand g1751(.dina(w_n2392_0[1]),.dinb(w_in256_0[0]),.dout(n2393),.clk(gclk));
	jand g1752(.dina(n2393),.dinb(w_n2375_0[0]),.dout(n2394),.clk(gclk));
	jor g1753(.dina(n2394),.dinb(n2391),.dout(n2395),.clk(gclk));
	jand g1754(.dina(n2395),.dinb(w_n2382_0[0]),.dout(n2396),.clk(gclk));
	jnot g1755(.din(w_n1970_0[0]),.dout(n2397),.clk(gclk));
	jnot g1756(.din(w_in361_0[0]),.dout(n2398),.clk(gclk));
	jand g1757(.dina(w_n2398_0[1]),.dinb(w_in261_0[0]),.dout(n2399),.clk(gclk));
	jnot g1758(.din(w_in360_0[0]),.dout(n2400),.clk(gclk));
	jand g1759(.dina(w_n2400_0[1]),.dinb(w_in260_0[0]),.dout(n2401),.clk(gclk));
	jor g1760(.dina(n2401),.dinb(n2399),.dout(n2402),.clk(gclk));
	jand g1761(.dina(n2402),.dinb(n2397),.dout(n2403),.clk(gclk));
	jnot g1762(.din(w_n1964_0[0]),.dout(n2404),.clk(gclk));
	jnot g1763(.din(w_in363_0[0]),.dout(n2405),.clk(gclk));
	jand g1764(.dina(w_n2405_0[1]),.dinb(w_in263_0[0]),.dout(n2406),.clk(gclk));
	jnot g1765(.din(w_in362_0[0]),.dout(n2407),.clk(gclk));
	jand g1766(.dina(w_n2407_0[1]),.dinb(w_in262_0[0]),.dout(n2408),.clk(gclk));
	jor g1767(.dina(n2408),.dinb(n2406),.dout(n2409),.clk(gclk));
	jand g1768(.dina(n2409),.dinb(n2404),.dout(n2410),.clk(gclk));
	jor g1769(.dina(n2410),.dinb(n2403),.dout(n2411),.clk(gclk));
	jor g1770(.dina(n2411),.dinb(n2396),.dout(n2412),.clk(gclk));
	jnot g1771(.din(w_n2412_0[1]),.dout(n2413),.clk(gclk));
	jand g1772(.dina(n2413),.dinb(n2386),.dout(n2414),.clk(gclk));
	jand g1773(.dina(n2414),.dinb(n1975),.dout(n2415),.clk(gclk));
	jnot g1774(.din(w_in264_0[0]),.dout(n2416),.clk(gclk));
	jand g1775(.dina(w_in364_0[0]),.dinb(w_n2416_0[1]),.dout(n2417),.clk(gclk));
	jor g1776(.dina(n2417),.dinb(w_n1948_0[0]),.dout(n2418),.clk(gclk));
	jor g1777(.dina(w_n2418_0[1]),.dinb(n2415),.dout(n2419),.clk(gclk));
	jand g1778(.dina(n2419),.dinb(n1959),.dout(n2420),.clk(gclk));
	jnot g1779(.din(w_in267_0[0]),.dout(n2421),.clk(gclk));
	jand g1780(.dina(w_in367_0[0]),.dinb(w_n2421_0[1]),.dout(n2422),.clk(gclk));
	jnot g1781(.din(w_in266_0[0]),.dout(n2423),.clk(gclk));
	jand g1782(.dina(w_in366_0[0]),.dinb(w_n2423_0[1]),.dout(n2424),.clk(gclk));
	jor g1783(.dina(n2424),.dinb(n2422),.dout(n2425),.clk(gclk));
	jor g1784(.dina(w_n2425_0[1]),.dinb(n2420),.dout(n2426),.clk(gclk));
	jand g1785(.dina(n2426),.dinb(n1946),.dout(n2427),.clk(gclk));
	jnot g1786(.din(w_in268_0[0]),.dout(n2428),.clk(gclk));
	jand g1787(.dina(w_in368_0[0]),.dinb(w_n2428_0[1]),.dout(n2429),.clk(gclk));
	jor g1788(.dina(n2429),.dinb(w_n1927_0[0]),.dout(n2430),.clk(gclk));
	jor g1789(.dina(w_n2430_0[1]),.dinb(n2427),.dout(n2431),.clk(gclk));
	jand g1790(.dina(n2431),.dinb(n1943),.dout(n2432),.clk(gclk));
	jnot g1791(.din(w_in275_0[0]),.dout(n2433),.clk(gclk));
	jand g1792(.dina(w_in375_0[0]),.dinb(w_n2433_0[1]),.dout(n2434),.clk(gclk));
	jnot g1793(.din(w_in274_0[1]),.dout(n2435),.clk(gclk));
	jand g1794(.dina(w_in374_0[1]),.dinb(w_n2435_0[1]),.dout(n2436),.clk(gclk));
	jor g1795(.dina(n2436),.dinb(n2434),.dout(n2437),.clk(gclk));
	jnot g1796(.din(w_in272_0[1]),.dout(n2438),.clk(gclk));
	jand g1797(.dina(w_in372_0[1]),.dinb(w_n2438_0[1]),.dout(n2439),.clk(gclk));
	jnot g1798(.din(w_in273_0[1]),.dout(n2440),.clk(gclk));
	jand g1799(.dina(w_in373_0[1]),.dinb(w_n2440_0[1]),.dout(n2441),.clk(gclk));
	jor g1800(.dina(w_n2441_0[1]),.dinb(n2439),.dout(n2442),.clk(gclk));
	jor g1801(.dina(n2442),.dinb(w_n2437_0[1]),.dout(n2443),.clk(gclk));
	jor g1802(.dina(w_n2443_0[1]),.dinb(n2432),.dout(n2444),.clk(gclk));
	jnot g1803(.din(w_n2437_0[0]),.dout(n2445),.clk(gclk));
	jnot g1804(.din(w_in373_0[0]),.dout(n2446),.clk(gclk));
	jand g1805(.dina(w_n2446_0[1]),.dinb(w_in273_0[0]),.dout(n2447),.clk(gclk));
	jnot g1806(.din(w_in374_0[0]),.dout(n2448),.clk(gclk));
	jand g1807(.dina(w_n2448_0[1]),.dinb(w_in274_0[0]),.dout(n2449),.clk(gclk));
	jor g1808(.dina(n2449),.dinb(n2447),.dout(n2450),.clk(gclk));
	jnot g1809(.din(w_n2441_0[0]),.dout(n2451),.clk(gclk));
	jnot g1810(.din(w_in372_0[0]),.dout(n2452),.clk(gclk));
	jand g1811(.dina(w_n2452_0[1]),.dinb(w_in272_0[0]),.dout(n2453),.clk(gclk));
	jand g1812(.dina(n2453),.dinb(n2451),.dout(n2454),.clk(gclk));
	jor g1813(.dina(n2454),.dinb(n2450),.dout(n2455),.clk(gclk));
	jand g1814(.dina(n2455),.dinb(n2445),.dout(n2456),.clk(gclk));
	jnot g1815(.din(w_n2456_0[1]),.dout(n2457),.clk(gclk));
	jand g1816(.dina(n2457),.dinb(n2444),.dout(n2458),.clk(gclk));
	jand g1817(.dina(n2458),.dinb(n1919),.dout(n2459),.clk(gclk));
	jnot g1818(.din(w_in276_0[0]),.dout(n2460),.clk(gclk));
	jand g1819(.dina(w_in376_0[0]),.dinb(w_n2460_0[1]),.dout(n2461),.clk(gclk));
	jor g1820(.dina(n2461),.dinb(w_n1900_0[0]),.dout(n2462),.clk(gclk));
	jor g1821(.dina(w_n2462_0[1]),.dinb(n2459),.dout(n2463),.clk(gclk));
	jand g1822(.dina(n2463),.dinb(n1916),.dout(n2464),.clk(gclk));
	jnot g1823(.din(w_in283_0[0]),.dout(n2465),.clk(gclk));
	jand g1824(.dina(w_in383_0[0]),.dinb(w_n2465_0[1]),.dout(n2466),.clk(gclk));
	jnot g1825(.din(w_in282_0[1]),.dout(n2467),.clk(gclk));
	jand g1826(.dina(w_in382_0[1]),.dinb(w_n2467_0[1]),.dout(n2468),.clk(gclk));
	jor g1827(.dina(n2468),.dinb(n2466),.dout(n2469),.clk(gclk));
	jor g1828(.dina(w_n2469_0[1]),.dinb(n2464),.dout(n2470),.clk(gclk));
	jor g1829(.dina(n2470),.dinb(w_n1892_0[1]),.dout(n2471),.clk(gclk));
	jnot g1830(.din(w_n2469_0[0]),.dout(n2472),.clk(gclk));
	jnot g1831(.din(w_in381_0[0]),.dout(n2473),.clk(gclk));
	jand g1832(.dina(w_n2473_0[1]),.dinb(w_in281_0[0]),.dout(n2474),.clk(gclk));
	jnot g1833(.din(w_in382_0[0]),.dout(n2475),.clk(gclk));
	jand g1834(.dina(w_n2475_0[1]),.dinb(w_in282_0[0]),.dout(n2476),.clk(gclk));
	jor g1835(.dina(n2476),.dinb(n2474),.dout(n2477),.clk(gclk));
	jnot g1836(.din(w_n1889_0[0]),.dout(n2478),.clk(gclk));
	jnot g1837(.din(w_in380_0[0]),.dout(n2479),.clk(gclk));
	jand g1838(.dina(w_n2479_0[1]),.dinb(w_in280_0[0]),.dout(n2480),.clk(gclk));
	jand g1839(.dina(n2480),.dinb(n2478),.dout(n2481),.clk(gclk));
	jor g1840(.dina(n2481),.dinb(n2477),.dout(n2482),.clk(gclk));
	jand g1841(.dina(n2482),.dinb(w_n2472_0[1]),.dout(n2483),.clk(gclk));
	jnot g1842(.din(w_n2483_0[1]),.dout(n2484),.clk(gclk));
	jand g1843(.dina(n2484),.dinb(n2471),.dout(n2485),.clk(gclk));
	jand g1844(.dina(n2485),.dinb(n1887),.dout(n2486),.clk(gclk));
	jnot g1845(.din(w_in284_0[0]),.dout(n2487),.clk(gclk));
	jand g1846(.dina(w_in384_0[0]),.dinb(w_n2487_0[1]),.dout(n2488),.clk(gclk));
	jor g1847(.dina(n2488),.dinb(w_n1868_0[0]),.dout(n2489),.clk(gclk));
	jor g1848(.dina(w_n2489_0[1]),.dinb(n2486),.dout(n2490),.clk(gclk));
	jand g1849(.dina(n2490),.dinb(n1884),.dout(n2491),.clk(gclk));
	jnot g1850(.din(w_in291_0[0]),.dout(n2492),.clk(gclk));
	jand g1851(.dina(w_in391_0[0]),.dinb(w_n2492_0[1]),.dout(n2493),.clk(gclk));
	jnot g1852(.din(w_in290_0[1]),.dout(n2494),.clk(gclk));
	jand g1853(.dina(w_in390_0[1]),.dinb(w_n2494_0[1]),.dout(n2495),.clk(gclk));
	jor g1854(.dina(n2495),.dinb(n2493),.dout(n2496),.clk(gclk));
	jnot g1855(.din(w_in288_0[1]),.dout(n2497),.clk(gclk));
	jand g1856(.dina(w_in388_0[1]),.dinb(w_n2497_0[1]),.dout(n2498),.clk(gclk));
	jnot g1857(.din(w_in289_0[1]),.dout(n2499),.clk(gclk));
	jand g1858(.dina(w_in389_0[1]),.dinb(w_n2499_0[1]),.dout(n2500),.clk(gclk));
	jor g1859(.dina(w_n2500_0[1]),.dinb(n2498),.dout(n2501),.clk(gclk));
	jor g1860(.dina(n2501),.dinb(w_n2496_0[1]),.dout(n2502),.clk(gclk));
	jor g1861(.dina(w_n2502_0[1]),.dinb(n2491),.dout(n2503),.clk(gclk));
	jnot g1862(.din(w_n2496_0[0]),.dout(n2504),.clk(gclk));
	jnot g1863(.din(w_in389_0[0]),.dout(n2505),.clk(gclk));
	jand g1864(.dina(w_n2505_0[1]),.dinb(w_in289_0[0]),.dout(n2506),.clk(gclk));
	jnot g1865(.din(w_in390_0[0]),.dout(n2507),.clk(gclk));
	jand g1866(.dina(w_n2507_0[1]),.dinb(w_in290_0[0]),.dout(n2508),.clk(gclk));
	jor g1867(.dina(n2508),.dinb(n2506),.dout(n2509),.clk(gclk));
	jnot g1868(.din(w_n2500_0[0]),.dout(n2510),.clk(gclk));
	jnot g1869(.din(w_in388_0[0]),.dout(n2511),.clk(gclk));
	jand g1870(.dina(w_n2511_0[1]),.dinb(w_in288_0[0]),.dout(n2512),.clk(gclk));
	jand g1871(.dina(n2512),.dinb(n2510),.dout(n2513),.clk(gclk));
	jor g1872(.dina(n2513),.dinb(n2509),.dout(n2514),.clk(gclk));
	jand g1873(.dina(n2514),.dinb(n2504),.dout(n2515),.clk(gclk));
	jnot g1874(.din(w_n2515_0[1]),.dout(n2516),.clk(gclk));
	jand g1875(.dina(n2516),.dinb(n2503),.dout(n2517),.clk(gclk));
	jand g1876(.dina(n2517),.dinb(n1860),.dout(n2518),.clk(gclk));
	jnot g1877(.din(w_in292_0[0]),.dout(n2519),.clk(gclk));
	jand g1878(.dina(w_in392_0[0]),.dinb(w_n2519_0[1]),.dout(n2520),.clk(gclk));
	jor g1879(.dina(n2520),.dinb(w_n1841_0[0]),.dout(n2521),.clk(gclk));
	jor g1880(.dina(w_n2521_0[1]),.dinb(n2518),.dout(n2522),.clk(gclk));
	jand g1881(.dina(n2522),.dinb(n1857),.dout(n2523),.clk(gclk));
	jnot g1882(.din(w_in299_0[0]),.dout(n2524),.clk(gclk));
	jand g1883(.dina(w_in399_0[0]),.dinb(w_n2524_0[1]),.dout(n2525),.clk(gclk));
	jnot g1884(.din(w_in298_0[1]),.dout(n2526),.clk(gclk));
	jand g1885(.dina(w_in398_0[1]),.dinb(w_n2526_0[1]),.dout(n2527),.clk(gclk));
	jor g1886(.dina(n2527),.dinb(n2525),.dout(n2528),.clk(gclk));
	jor g1887(.dina(w_n2528_0[1]),.dinb(n2523),.dout(n2529),.clk(gclk));
	jor g1888(.dina(n2529),.dinb(w_n1833_0[1]),.dout(n2530),.clk(gclk));
	jnot g1889(.din(w_n2528_0[0]),.dout(n2531),.clk(gclk));
	jnot g1890(.din(w_in397_0[0]),.dout(n2532),.clk(gclk));
	jand g1891(.dina(w_n2532_0[1]),.dinb(w_in297_0[0]),.dout(n2533),.clk(gclk));
	jnot g1892(.din(w_in398_0[0]),.dout(n2534),.clk(gclk));
	jand g1893(.dina(w_n2534_0[1]),.dinb(w_in298_0[0]),.dout(n2535),.clk(gclk));
	jor g1894(.dina(n2535),.dinb(n2533),.dout(n2536),.clk(gclk));
	jnot g1895(.din(w_n1830_0[0]),.dout(n2537),.clk(gclk));
	jnot g1896(.din(w_in396_0[0]),.dout(n2538),.clk(gclk));
	jand g1897(.dina(w_n2538_0[1]),.dinb(w_in296_0[0]),.dout(n2539),.clk(gclk));
	jand g1898(.dina(n2539),.dinb(n2537),.dout(n2540),.clk(gclk));
	jor g1899(.dina(n2540),.dinb(n2536),.dout(n2541),.clk(gclk));
	jand g1900(.dina(n2541),.dinb(w_n2531_0[1]),.dout(n2542),.clk(gclk));
	jnot g1901(.din(w_n2542_0[1]),.dout(n2543),.clk(gclk));
	jand g1902(.dina(n2543),.dinb(n2530),.dout(n2544),.clk(gclk));
	jand g1903(.dina(n2544),.dinb(n1828),.dout(n2545),.clk(gclk));
	jnot g1904(.din(w_in2100_0[0]),.dout(n2546),.clk(gclk));
	jand g1905(.dina(w_in3100_0[0]),.dinb(w_n2546_0[1]),.dout(n2547),.clk(gclk));
	jor g1906(.dina(n2547),.dinb(w_n1809_0[0]),.dout(n2548),.clk(gclk));
	jor g1907(.dina(w_n2548_0[1]),.dinb(n2545),.dout(n2549),.clk(gclk));
	jand g1908(.dina(n2549),.dinb(n1825),.dout(n2550),.clk(gclk));
	jnot g1909(.din(w_in2107_0[0]),.dout(n2551),.clk(gclk));
	jand g1910(.dina(w_in3107_0[0]),.dinb(w_n2551_0[1]),.dout(n2552),.clk(gclk));
	jnot g1911(.din(w_in2106_0[1]),.dout(n2553),.clk(gclk));
	jand g1912(.dina(w_in3106_0[1]),.dinb(w_n2553_0[1]),.dout(n2554),.clk(gclk));
	jor g1913(.dina(n2554),.dinb(n2552),.dout(n2555),.clk(gclk));
	jnot g1914(.din(w_in2104_0[1]),.dout(n2556),.clk(gclk));
	jand g1915(.dina(w_in3104_0[1]),.dinb(w_n2556_0[1]),.dout(n2557),.clk(gclk));
	jnot g1916(.din(w_in2105_0[1]),.dout(n2558),.clk(gclk));
	jand g1917(.dina(w_in3105_0[1]),.dinb(w_n2558_0[1]),.dout(n2559),.clk(gclk));
	jor g1918(.dina(w_n2559_0[1]),.dinb(n2557),.dout(n2560),.clk(gclk));
	jor g1919(.dina(n2560),.dinb(w_n2555_0[1]),.dout(n2561),.clk(gclk));
	jor g1920(.dina(w_n2561_0[1]),.dinb(n2550),.dout(n2562),.clk(gclk));
	jnot g1921(.din(w_n2555_0[0]),.dout(n2563),.clk(gclk));
	jnot g1922(.din(w_in3105_0[0]),.dout(n2564),.clk(gclk));
	jand g1923(.dina(w_n2564_0[1]),.dinb(w_in2105_0[0]),.dout(n2565),.clk(gclk));
	jnot g1924(.din(w_in3106_0[0]),.dout(n2566),.clk(gclk));
	jand g1925(.dina(w_n2566_0[1]),.dinb(w_in2106_0[0]),.dout(n2567),.clk(gclk));
	jor g1926(.dina(n2567),.dinb(n2565),.dout(n2568),.clk(gclk));
	jnot g1927(.din(w_n2559_0[0]),.dout(n2569),.clk(gclk));
	jnot g1928(.din(w_in3104_0[0]),.dout(n2570),.clk(gclk));
	jand g1929(.dina(w_n2570_0[1]),.dinb(w_in2104_0[0]),.dout(n2571),.clk(gclk));
	jand g1930(.dina(n2571),.dinb(n2569),.dout(n2572),.clk(gclk));
	jor g1931(.dina(n2572),.dinb(n2568),.dout(n2573),.clk(gclk));
	jand g1932(.dina(n2573),.dinb(n2563),.dout(n2574),.clk(gclk));
	jnot g1933(.din(w_n2574_0[1]),.dout(n2575),.clk(gclk));
	jand g1934(.dina(n2575),.dinb(n2562),.dout(n2576),.clk(gclk));
	jand g1935(.dina(n2576),.dinb(n1801),.dout(n2577),.clk(gclk));
	jnot g1936(.din(w_in2108_0[0]),.dout(n2578),.clk(gclk));
	jand g1937(.dina(w_in3108_0[0]),.dinb(w_n2578_0[1]),.dout(n2579),.clk(gclk));
	jor g1938(.dina(n2579),.dinb(w_n1782_0[0]),.dout(n2580),.clk(gclk));
	jor g1939(.dina(w_n2580_0[1]),.dinb(n2577),.dout(n2581),.clk(gclk));
	jand g1940(.dina(n2581),.dinb(n1798),.dout(n2582),.clk(gclk));
	jnot g1941(.din(w_in2115_0[0]),.dout(n2583),.clk(gclk));
	jand g1942(.dina(w_in3115_0[0]),.dinb(w_n2583_0[1]),.dout(n2584),.clk(gclk));
	jnot g1943(.din(w_in2114_0[1]),.dout(n2585),.clk(gclk));
	jand g1944(.dina(w_in3114_0[1]),.dinb(w_n2585_0[1]),.dout(n2586),.clk(gclk));
	jor g1945(.dina(n2586),.dinb(n2584),.dout(n2587),.clk(gclk));
	jor g1946(.dina(w_n2587_0[1]),.dinb(n2582),.dout(n2588),.clk(gclk));
	jor g1947(.dina(n2588),.dinb(w_n1774_0[1]),.dout(n2589),.clk(gclk));
	jnot g1948(.din(w_n2587_0[0]),.dout(n2590),.clk(gclk));
	jnot g1949(.din(w_in3113_0[0]),.dout(n2591),.clk(gclk));
	jand g1950(.dina(w_n2591_0[1]),.dinb(w_in2113_0[0]),.dout(n2592),.clk(gclk));
	jnot g1951(.din(w_in3114_0[0]),.dout(n2593),.clk(gclk));
	jand g1952(.dina(w_n2593_0[1]),.dinb(w_in2114_0[0]),.dout(n2594),.clk(gclk));
	jor g1953(.dina(n2594),.dinb(n2592),.dout(n2595),.clk(gclk));
	jnot g1954(.din(w_n1771_0[0]),.dout(n2596),.clk(gclk));
	jnot g1955(.din(w_in3112_0[0]),.dout(n2597),.clk(gclk));
	jand g1956(.dina(w_n2597_0[1]),.dinb(w_in2112_0[0]),.dout(n2598),.clk(gclk));
	jand g1957(.dina(n2598),.dinb(n2596),.dout(n2599),.clk(gclk));
	jor g1958(.dina(n2599),.dinb(n2595),.dout(n2600),.clk(gclk));
	jand g1959(.dina(n2600),.dinb(w_n2590_0[1]),.dout(n2601),.clk(gclk));
	jnot g1960(.din(w_n2601_0[1]),.dout(n2602),.clk(gclk));
	jand g1961(.dina(n2602),.dinb(n2589),.dout(n2603),.clk(gclk));
	jand g1962(.dina(n2603),.dinb(n1769),.dout(n2604),.clk(gclk));
	jnot g1963(.din(w_in2116_0[0]),.dout(n2605),.clk(gclk));
	jand g1964(.dina(w_in3116_0[0]),.dinb(w_n2605_0[1]),.dout(n2606),.clk(gclk));
	jor g1965(.dina(n2606),.dinb(w_n1750_0[0]),.dout(n2607),.clk(gclk));
	jor g1966(.dina(w_n2607_0[1]),.dinb(n2604),.dout(n2608),.clk(gclk));
	jand g1967(.dina(n2608),.dinb(n1766),.dout(n2609),.clk(gclk));
	jnot g1968(.din(w_in2123_0[0]),.dout(n2610),.clk(gclk));
	jand g1969(.dina(w_in3123_0[0]),.dinb(w_n2610_0[1]),.dout(n2611),.clk(gclk));
	jnot g1970(.din(w_in2122_0[1]),.dout(n2612),.clk(gclk));
	jand g1971(.dina(w_in3122_0[1]),.dinb(w_n2612_0[1]),.dout(n2613),.clk(gclk));
	jor g1972(.dina(n2613),.dinb(n2611),.dout(n2614),.clk(gclk));
	jnot g1973(.din(w_in2120_0[1]),.dout(n2615),.clk(gclk));
	jand g1974(.dina(w_in3120_0[1]),.dinb(w_n2615_0[1]),.dout(n2616),.clk(gclk));
	jnot g1975(.din(w_in2121_0[1]),.dout(n2617),.clk(gclk));
	jand g1976(.dina(w_in3121_0[1]),.dinb(w_n2617_0[1]),.dout(n2618),.clk(gclk));
	jor g1977(.dina(w_n2618_0[1]),.dinb(n2616),.dout(n2619),.clk(gclk));
	jor g1978(.dina(n2619),.dinb(w_n2614_0[1]),.dout(n2620),.clk(gclk));
	jor g1979(.dina(w_n2620_0[1]),.dinb(n2609),.dout(n2621),.clk(gclk));
	jnot g1980(.din(w_n2614_0[0]),.dout(n2622),.clk(gclk));
	jnot g1981(.din(w_in3121_0[0]),.dout(n2623),.clk(gclk));
	jand g1982(.dina(w_n2623_0[1]),.dinb(w_in2121_0[0]),.dout(n2624),.clk(gclk));
	jnot g1983(.din(w_in3122_0[0]),.dout(n2625),.clk(gclk));
	jand g1984(.dina(w_n2625_0[1]),.dinb(w_in2122_0[0]),.dout(n2626),.clk(gclk));
	jor g1985(.dina(n2626),.dinb(n2624),.dout(n2627),.clk(gclk));
	jnot g1986(.din(w_n2618_0[0]),.dout(n2628),.clk(gclk));
	jnot g1987(.din(w_in3120_0[0]),.dout(n2629),.clk(gclk));
	jand g1988(.dina(w_n2629_0[1]),.dinb(w_in2120_0[0]),.dout(n2630),.clk(gclk));
	jand g1989(.dina(n2630),.dinb(n2628),.dout(n2631),.clk(gclk));
	jor g1990(.dina(n2631),.dinb(n2627),.dout(n2632),.clk(gclk));
	jand g1991(.dina(n2632),.dinb(n2622),.dout(n2633),.clk(gclk));
	jnot g1992(.din(w_n2633_0[1]),.dout(n2634),.clk(gclk));
	jand g1993(.dina(n2634),.dinb(n2621),.dout(n2635),.clk(gclk));
	jand g1994(.dina(n2635),.dinb(n1742),.dout(n2636),.clk(gclk));
	jnot g1995(.din(w_in2124_0[0]),.dout(n2637),.clk(gclk));
	jand g1996(.dina(w_in3124_0[0]),.dinb(w_n2637_0[1]),.dout(n2638),.clk(gclk));
	jor g1997(.dina(n2638),.dinb(w_n1728_0[0]),.dout(n2639),.clk(gclk));
	jnot g1998(.din(w_n2639_0[1]),.dout(n2640),.clk(gclk));
	jand g1999(.dina(w_in3127_0[1]),.dinb(w_in2127_0[2]),.dout(n2641),.clk(gclk));
	jnot g2000(.din(w_n2641_0[2]),.dout(n2642),.clk(gclk));
	jand g2001(.dina(w_in1127_0[0]),.dinb(w_in0127_0[0]),.dout(n2643),.clk(gclk));
	jand g2002(.dina(w_n2643_1[1]),.dinb(w_n2642_0[1]),.dout(n2644),.clk(gclk));
	jand g2003(.dina(w_n1721_65[0]),.dinb(w_n1534_0[0]),.dout(n2645),.clk(gclk));
	jand g2004(.dina(w_n1562_64[1]),.dinb(w_n1554_0[0]),.dout(n2646),.clk(gclk));
	jor g2005(.dina(n2646),.dinb(n2645),.dout(n2647),.clk(gclk));
	jnot g2006(.din(w_in3127_0[0]),.dout(n2648),.clk(gclk));
	jand g2007(.dina(w_n2648_0[1]),.dinb(w_in2127_0[1]),.dout(n2649),.clk(gclk));
	jnot g2008(.din(w_n2649_0[1]),.dout(n2650),.clk(gclk));
	jnot g2009(.din(w_n1774_0[0]),.dout(n2651),.clk(gclk));
	jnot g2010(.din(w_n1833_0[0]),.dout(n2652),.clk(gclk));
	jnot g2011(.din(w_n1892_0[0]),.dout(n2653),.clk(gclk));
	jnot g2012(.din(w_n2041_0[0]),.dout(n2654),.clk(gclk));
	jnot g2013(.din(w_n2046_0[0]),.dout(n2655),.clk(gclk));
	jnot g2014(.din(w_n2051_0[0]),.dout(n2656),.clk(gclk));
	jnot g2015(.din(w_n2056_0[0]),.dout(n2657),.clk(gclk));
	jnot g2016(.din(w_n2061_0[0]),.dout(n2658),.clk(gclk));
	jnot g2017(.din(w_n2063_0[0]),.dout(n2659),.clk(gclk));
	jnot g2018(.din(w_n2068_0[0]),.dout(n2660),.clk(gclk));
	jnot g2019(.din(w_n2073_0[0]),.dout(n2661),.clk(gclk));
	jnot g2020(.din(w_n2078_0[0]),.dout(n2662),.clk(gclk));
	jnot g2021(.din(w_n2083_0[0]),.dout(n2663),.clk(gclk));
	jnot g2022(.din(w_n2085_0[0]),.dout(n2664),.clk(gclk));
	jnot g2023(.din(w_n2090_0[0]),.dout(n2665),.clk(gclk));
	jnot g2024(.din(w_n2095_0[0]),.dout(n2666),.clk(gclk));
	jnot g2025(.din(w_n2100_0[0]),.dout(n2667),.clk(gclk));
	jnot g2026(.din(w_n2105_0[0]),.dout(n2668),.clk(gclk));
	jnot g2027(.din(w_n2107_0[0]),.dout(n2669),.clk(gclk));
	jnot g2028(.din(w_n2109_0[0]),.dout(n2670),.clk(gclk));
	jor g2029(.dina(w_n2110_0[1]),.dinb(w_in21_0[2]),.dout(n2671),.clk(gclk));
	jnot g2030(.din(w_in30_0[1]),.dout(n2672),.clk(gclk));
	jand g2031(.dina(w_n2672_0[1]),.dinb(w_in20_0[1]),.dout(n2673),.clk(gclk));
	jand g2032(.dina(n2673),.dinb(n2671),.dout(n2674),.clk(gclk));
	jor g2033(.dina(n2674),.dinb(w_n2111_0[0]),.dout(n2675),.clk(gclk));
	jand g2034(.dina(n2675),.dinb(n2670),.dout(n2676),.clk(gclk));
	jor g2035(.dina(w_n2124_0[0]),.dinb(n2676),.dout(n2677),.clk(gclk));
	jnot g2036(.din(w_n2128_0[0]),.dout(n2678),.clk(gclk));
	jand g2037(.dina(n2678),.dinb(n2677),.dout(n2679),.clk(gclk));
	jand g2038(.dina(n2679),.dinb(n2669),.dout(n2680),.clk(gclk));
	jor g2039(.dina(w_n2135_0[0]),.dinb(n2680),.dout(n2681),.clk(gclk));
	jnot g2040(.din(w_n2142_0[0]),.dout(n2682),.clk(gclk));
	jand g2041(.dina(n2682),.dinb(n2681),.dout(n2683),.clk(gclk));
	jor g2042(.dina(w_n2148_0[0]),.dinb(n2683),.dout(n2684),.clk(gclk));
	jnot g2043(.din(w_n2152_0[0]),.dout(n2685),.clk(gclk));
	jand g2044(.dina(n2685),.dinb(n2684),.dout(n2686),.clk(gclk));
	jand g2045(.dina(n2686),.dinb(n2668),.dout(n2687),.clk(gclk));
	jor g2046(.dina(w_n2159_0[0]),.dinb(n2687),.dout(n2688),.clk(gclk));
	jnot g2047(.din(w_n2166_0[0]),.dout(n2689),.clk(gclk));
	jand g2048(.dina(n2689),.dinb(n2688),.dout(n2690),.clk(gclk));
	jor g2049(.dina(n2690),.dinb(w_n2102_0[0]),.dout(n2691),.clk(gclk));
	jand g2050(.dina(n2691),.dinb(n2667),.dout(n2692),.clk(gclk));
	jor g2051(.dina(n2692),.dinb(w_n2097_0[0]),.dout(n2693),.clk(gclk));
	jand g2052(.dina(n2693),.dinb(n2666),.dout(n2694),.clk(gclk));
	jor g2053(.dina(n2694),.dinb(w_n2092_0[0]),.dout(n2695),.clk(gclk));
	jand g2054(.dina(n2695),.dinb(n2665),.dout(n2696),.clk(gclk));
	jor g2055(.dina(n2696),.dinb(w_n2087_0[0]),.dout(n2697),.clk(gclk));
	jand g2056(.dina(n2697),.dinb(n2664),.dout(n2698),.clk(gclk));
	jor g2057(.dina(w_n2180_0[0]),.dinb(n2698),.dout(n2699),.clk(gclk));
	jnot g2058(.din(w_n2184_0[0]),.dout(n2700),.clk(gclk));
	jand g2059(.dina(n2700),.dinb(n2699),.dout(n2701),.clk(gclk));
	jand g2060(.dina(n2701),.dinb(n2663),.dout(n2702),.clk(gclk));
	jor g2061(.dina(w_n2191_0[0]),.dinb(n2702),.dout(n2703),.clk(gclk));
	jnot g2062(.din(w_n2198_0[0]),.dout(n2704),.clk(gclk));
	jand g2063(.dina(n2704),.dinb(n2703),.dout(n2705),.clk(gclk));
	jor g2064(.dina(n2705),.dinb(w_n2080_0[0]),.dout(n2706),.clk(gclk));
	jand g2065(.dina(n2706),.dinb(n2662),.dout(n2707),.clk(gclk));
	jor g2066(.dina(n2707),.dinb(w_n2075_0[0]),.dout(n2708),.clk(gclk));
	jand g2067(.dina(n2708),.dinb(n2661),.dout(n2709),.clk(gclk));
	jor g2068(.dina(n2709),.dinb(w_n2070_0[0]),.dout(n2710),.clk(gclk));
	jand g2069(.dina(n2710),.dinb(n2660),.dout(n2711),.clk(gclk));
	jor g2070(.dina(n2711),.dinb(w_n2065_0[0]),.dout(n2712),.clk(gclk));
	jand g2071(.dina(n2712),.dinb(n2659),.dout(n2713),.clk(gclk));
	jor g2072(.dina(w_n2212_0[0]),.dinb(n2713),.dout(n2714),.clk(gclk));
	jnot g2073(.din(w_n2216_0[0]),.dout(n2715),.clk(gclk));
	jand g2074(.dina(n2715),.dinb(n2714),.dout(n2716),.clk(gclk));
	jand g2075(.dina(n2716),.dinb(n2658),.dout(n2717),.clk(gclk));
	jor g2076(.dina(w_n2223_0[0]),.dinb(n2717),.dout(n2718),.clk(gclk));
	jnot g2077(.din(w_n2230_0[0]),.dout(n2719),.clk(gclk));
	jand g2078(.dina(n2719),.dinb(n2718),.dout(n2720),.clk(gclk));
	jor g2079(.dina(n2720),.dinb(w_n2058_0[0]),.dout(n2721),.clk(gclk));
	jand g2080(.dina(n2721),.dinb(n2657),.dout(n2722),.clk(gclk));
	jor g2081(.dina(n2722),.dinb(w_n2053_0[0]),.dout(n2723),.clk(gclk));
	jand g2082(.dina(n2723),.dinb(n2656),.dout(n2724),.clk(gclk));
	jor g2083(.dina(n2724),.dinb(w_n2048_0[0]),.dout(n2725),.clk(gclk));
	jand g2084(.dina(n2725),.dinb(n2655),.dout(n2726),.clk(gclk));
	jor g2085(.dina(n2726),.dinb(w_n2043_0[0]),.dout(n2727),.clk(gclk));
	jand g2086(.dina(n2727),.dinb(n2654),.dout(n2728),.clk(gclk));
	jor g2087(.dina(w_n2244_0[0]),.dinb(n2728),.dout(n2729),.clk(gclk));
	jnot g2088(.din(w_n2253_0[0]),.dout(n2730),.clk(gclk));
	jand g2089(.dina(n2730),.dinb(n2729),.dout(n2731),.clk(gclk));
	jor g2090(.dina(w_n2274_0[0]),.dinb(n2731),.dout(n2732),.clk(gclk));
	jor g2091(.dina(n2732),.dinb(w_n2038_0[0]),.dout(n2733),.clk(gclk));
	jand g2092(.dina(w_n2292_0[0]),.dinb(n2733),.dout(n2734),.clk(gclk));
	jor g2093(.dina(w_n2320_0[0]),.dinb(n2734),.dout(n2735),.clk(gclk));
	jor g2094(.dina(n2735),.dinb(w_n2006_0[0]),.dout(n2736),.clk(gclk));
	jand g2095(.dina(w_n2338_0[0]),.dinb(n2736),.dout(n2737),.clk(gclk));
	jor g2096(.dina(w_n2366_0[0]),.dinb(n2737),.dout(n2738),.clk(gclk));
	jor g2097(.dina(n2738),.dinb(w_n1990_0[0]),.dout(n2739),.clk(gclk));
	jand g2098(.dina(w_n2384_0[0]),.dinb(n2739),.dout(n2740),.clk(gclk));
	jor g2099(.dina(w_n2412_0[0]),.dinb(n2740),.dout(n2741),.clk(gclk));
	jor g2100(.dina(n2741),.dinb(w_n1974_0[0]),.dout(n2742),.clk(gclk));
	jnot g2101(.din(w_n2418_0[0]),.dout(n2743),.clk(gclk));
	jand g2102(.dina(n2743),.dinb(n2742),.dout(n2744),.clk(gclk));
	jor g2103(.dina(n2744),.dinb(w_n1958_0[0]),.dout(n2745),.clk(gclk));
	jnot g2104(.din(w_n2425_0[0]),.dout(n2746),.clk(gclk));
	jand g2105(.dina(n2746),.dinb(n2745),.dout(n2747),.clk(gclk));
	jor g2106(.dina(n2747),.dinb(w_n1945_0[0]),.dout(n2748),.clk(gclk));
	jnot g2107(.din(w_n2430_0[0]),.dout(n2749),.clk(gclk));
	jand g2108(.dina(n2749),.dinb(n2748),.dout(n2750),.clk(gclk));
	jor g2109(.dina(n2750),.dinb(w_n1942_0[0]),.dout(n2751),.clk(gclk));
	jnot g2110(.din(w_n2443_0[0]),.dout(n2752),.clk(gclk));
	jand g2111(.dina(n2752),.dinb(n2751),.dout(n2753),.clk(gclk));
	jor g2112(.dina(w_n2456_0[0]),.dinb(n2753),.dout(n2754),.clk(gclk));
	jor g2113(.dina(n2754),.dinb(w_n1918_0[0]),.dout(n2755),.clk(gclk));
	jnot g2114(.din(w_n2462_0[0]),.dout(n2756),.clk(gclk));
	jand g2115(.dina(n2756),.dinb(n2755),.dout(n2757),.clk(gclk));
	jor g2116(.dina(n2757),.dinb(w_n1915_0[0]),.dout(n2758),.clk(gclk));
	jand g2117(.dina(w_n2472_0[0]),.dinb(n2758),.dout(n2759),.clk(gclk));
	jand g2118(.dina(n2759),.dinb(n2653),.dout(n2760),.clk(gclk));
	jor g2119(.dina(w_n2483_0[0]),.dinb(n2760),.dout(n2761),.clk(gclk));
	jor g2120(.dina(n2761),.dinb(w_n1886_0[0]),.dout(n2762),.clk(gclk));
	jnot g2121(.din(w_n2489_0[0]),.dout(n2763),.clk(gclk));
	jand g2122(.dina(n2763),.dinb(n2762),.dout(n2764),.clk(gclk));
	jor g2123(.dina(n2764),.dinb(w_n1883_0[0]),.dout(n2765),.clk(gclk));
	jnot g2124(.din(w_n2502_0[0]),.dout(n2766),.clk(gclk));
	jand g2125(.dina(n2766),.dinb(n2765),.dout(n2767),.clk(gclk));
	jor g2126(.dina(w_n2515_0[0]),.dinb(n2767),.dout(n2768),.clk(gclk));
	jor g2127(.dina(n2768),.dinb(w_n1859_0[0]),.dout(n2769),.clk(gclk));
	jnot g2128(.din(w_n2521_0[0]),.dout(n2770),.clk(gclk));
	jand g2129(.dina(n2770),.dinb(n2769),.dout(n2771),.clk(gclk));
	jor g2130(.dina(n2771),.dinb(w_n1856_0[0]),.dout(n2772),.clk(gclk));
	jand g2131(.dina(w_n2531_0[0]),.dinb(n2772),.dout(n2773),.clk(gclk));
	jand g2132(.dina(n2773),.dinb(n2652),.dout(n2774),.clk(gclk));
	jor g2133(.dina(w_n2542_0[0]),.dinb(n2774),.dout(n2775),.clk(gclk));
	jor g2134(.dina(n2775),.dinb(w_n1827_0[0]),.dout(n2776),.clk(gclk));
	jnot g2135(.din(w_n2548_0[0]),.dout(n2777),.clk(gclk));
	jand g2136(.dina(n2777),.dinb(n2776),.dout(n2778),.clk(gclk));
	jor g2137(.dina(n2778),.dinb(w_n1824_0[0]),.dout(n2779),.clk(gclk));
	jnot g2138(.din(w_n2561_0[0]),.dout(n2780),.clk(gclk));
	jand g2139(.dina(n2780),.dinb(n2779),.dout(n2781),.clk(gclk));
	jor g2140(.dina(w_n2574_0[0]),.dinb(n2781),.dout(n2782),.clk(gclk));
	jor g2141(.dina(n2782),.dinb(w_n1800_0[0]),.dout(n2783),.clk(gclk));
	jnot g2142(.din(w_n2580_0[0]),.dout(n2784),.clk(gclk));
	jand g2143(.dina(n2784),.dinb(n2783),.dout(n2785),.clk(gclk));
	jor g2144(.dina(n2785),.dinb(w_n1797_0[0]),.dout(n2786),.clk(gclk));
	jand g2145(.dina(w_n2590_0[0]),.dinb(n2786),.dout(n2787),.clk(gclk));
	jand g2146(.dina(n2787),.dinb(n2651),.dout(n2788),.clk(gclk));
	jor g2147(.dina(w_n2601_0[0]),.dinb(n2788),.dout(n2789),.clk(gclk));
	jor g2148(.dina(n2789),.dinb(w_n1768_0[0]),.dout(n2790),.clk(gclk));
	jnot g2149(.din(w_n2607_0[0]),.dout(n2791),.clk(gclk));
	jand g2150(.dina(n2791),.dinb(n2790),.dout(n2792),.clk(gclk));
	jor g2151(.dina(n2792),.dinb(w_n1765_0[0]),.dout(n2793),.clk(gclk));
	jnot g2152(.din(w_n2620_0[0]),.dout(n2794),.clk(gclk));
	jand g2153(.dina(n2794),.dinb(n2793),.dout(n2795),.clk(gclk));
	jor g2154(.dina(w_n2633_0[0]),.dinb(n2795),.dout(n2796),.clk(gclk));
	jor g2155(.dina(n2796),.dinb(w_n1741_0[0]),.dout(n2797),.clk(gclk));
	jand g2156(.dina(n2640),.dinb(n2797),.dout(n2798),.clk(gclk));
	jor g2157(.dina(n2798),.dinb(w_n1738_0[0]),.dout(n2799),.clk(gclk));
	jand g2158(.dina(n2799),.dinb(n2650),.dout(n2800),.clk(gclk));
	jor g2159(.dina(w_n2648_0[0]),.dinb(w_in2127_0[0]),.dout(n2801),.clk(gclk));
	jnot g2160(.din(w_n2801_0[1]),.dout(n2802),.clk(gclk));
	jor g2161(.dina(n2802),.dinb(n2800),.dout(n2803),.clk(gclk));
	jand g2162(.dina(w_n2803_64[1]),.dinb(w_n1724_0[0]),.dout(n2804),.clk(gclk));
	jor g2163(.dina(w_n2639_0[0]),.dinb(n2636),.dout(n2805),.clk(gclk));
	jand g2164(.dina(n2805),.dinb(n1739),.dout(n2806),.clk(gclk));
	jor g2165(.dina(n2806),.dinb(w_n2649_0[0]),.dout(n2807),.clk(gclk));
	jand g2166(.dina(w_n2801_0[0]),.dinb(n2807),.dout(n2808),.clk(gclk));
	jand g2167(.dina(w_n2808_64[2]),.dinb(w_n1736_0[0]),.dout(n2809),.clk(gclk));
	jor g2168(.dina(n2809),.dinb(n2804),.dout(n2810),.clk(gclk));
	jnot g2169(.din(w_n2810_0[1]),.dout(n2811),.clk(gclk));
	jand g2170(.dina(w_n2811_0[1]),.dinb(w_n2647_0[1]),.dout(n2812),.clk(gclk));
	jand g2171(.dina(w_n1721_64[2]),.dinb(w_n1536_0[0]),.dout(n2813),.clk(gclk));
	jand g2172(.dina(w_n1562_64[0]),.dinb(w_n1550_0[0]),.dout(n2814),.clk(gclk));
	jor g2173(.dina(n2814),.dinb(n2813),.dout(n2815),.clk(gclk));
	jand g2174(.dina(w_n2803_64[0]),.dinb(w_n1726_0[0]),.dout(n2816),.clk(gclk));
	jand g2175(.dina(w_n2808_64[1]),.dinb(w_n1732_0[0]),.dout(n2817),.clk(gclk));
	jor g2176(.dina(n2817),.dinb(n2816),.dout(n2818),.clk(gclk));
	jnot g2177(.din(w_n2818_0[1]),.dout(n2819),.clk(gclk));
	jand g2178(.dina(w_n2819_0[1]),.dinb(w_n2815_0[1]),.dout(n2820),.clk(gclk));
	jor g2179(.dina(n2820),.dinb(n2812),.dout(n2821),.clk(gclk));
	jnot g2180(.din(w_n2821_0[1]),.dout(n2822),.clk(gclk));
	jand g2181(.dina(w_n1721_64[1]),.dinb(w_n1539_0[0]),.dout(n2823),.clk(gclk));
	jand g2182(.dina(w_n1562_63[2]),.dinb(w_n1548_0[0]),.dout(n2824),.clk(gclk));
	jor g2183(.dina(n2824),.dinb(n2823),.dout(n2825),.clk(gclk));
	jnot g2184(.din(w_n2825_0[1]),.dout(n2826),.clk(gclk));
	jand g2185(.dina(w_n2803_63[2]),.dinb(w_n2637_0[0]),.dout(n2827),.clk(gclk));
	jand g2186(.dina(w_n2808_64[0]),.dinb(w_n1730_0[0]),.dout(n2828),.clk(gclk));
	jor g2187(.dina(n2828),.dinb(n2827),.dout(n2829),.clk(gclk));
	jand g2188(.dina(w_n2829_0[1]),.dinb(w_n2826_0[1]),.dout(n2830),.clk(gclk));
	jnot g2189(.din(w_n2815_0[0]),.dout(n2831),.clk(gclk));
	jand g2190(.dina(w_n2818_0[0]),.dinb(w_n2831_0[1]),.dout(n2832),.clk(gclk));
	jor g2191(.dina(n2832),.dinb(n2830),.dout(n2833),.clk(gclk));
	jand g2192(.dina(n2833),.dinb(n2822),.dout(n2834),.clk(gclk));
	jnot g2193(.din(w_n2647_0[0]),.dout(n2835),.clk(gclk));
	jand g2194(.dina(w_n2810_0[0]),.dinb(w_n2835_0[1]),.dout(n2836),.clk(gclk));
	jor g2195(.dina(n2836),.dinb(n2834),.dout(n2837),.clk(gclk));
	jnot g2196(.din(w_n2837_0[1]),.dout(n2838),.clk(gclk));
	jnot g2197(.din(w_n2829_0[0]),.dout(n2839),.clk(gclk));
	jand g2198(.dina(w_n2839_0[1]),.dinb(w_n2825_0[0]),.dout(n2840),.clk(gclk));
	jor g2199(.dina(n2840),.dinb(w_n2821_0[0]),.dout(n2841),.clk(gclk));
	jand g2200(.dina(w_n2803_63[1]),.dinb(w_n1743_0[0]),.dout(n2842),.clk(gclk));
	jand g2201(.dina(w_n2808_63[2]),.dinb(w_n1761_0[0]),.dout(n2843),.clk(gclk));
	jor g2202(.dina(n2843),.dinb(n2842),.dout(n2844),.clk(gclk));
	jnot g2203(.din(w_n2844_0[1]),.dout(n2845),.clk(gclk));
	jand g2204(.dina(w_n1721_64[0]),.dinb(w_n650_0[0]),.dout(n2846),.clk(gclk));
	jand g2205(.dina(w_n1562_63[1]),.dinb(w_n668_0[0]),.dout(n2847),.clk(gclk));
	jor g2206(.dina(n2847),.dinb(n2846),.dout(n2848),.clk(gclk));
	jand g2207(.dina(w_n2848_0[1]),.dinb(w_n2845_0[1]),.dout(n2849),.clk(gclk));
	jand g2208(.dina(w_n1721_63[2]),.dinb(w_n652_0[0]),.dout(n2850),.clk(gclk));
	jand g2209(.dina(w_n1562_63[0]),.dinb(w_n666_0[0]),.dout(n2851),.clk(gclk));
	jor g2210(.dina(n2851),.dinb(n2850),.dout(n2852),.clk(gclk));
	jand g2211(.dina(w_n2803_63[0]),.dinb(w_n1745_0[0]),.dout(n2853),.clk(gclk));
	jand g2212(.dina(w_n2808_63[1]),.dinb(w_n1759_0[0]),.dout(n2854),.clk(gclk));
	jor g2213(.dina(n2854),.dinb(n2853),.dout(n2855),.clk(gclk));
	jnot g2214(.din(w_n2855_0[1]),.dout(n2856),.clk(gclk));
	jand g2215(.dina(w_n2856_0[1]),.dinb(w_n2852_0[1]),.dout(n2857),.clk(gclk));
	jand g2216(.dina(w_n1721_63[1]),.dinb(w_n654_0[0]),.dout(n2858),.clk(gclk));
	jand g2217(.dina(w_n1562_62[2]),.dinb(w_n659_0[0]),.dout(n2859),.clk(gclk));
	jor g2218(.dina(n2859),.dinb(n2858),.dout(n2860),.clk(gclk));
	jand g2219(.dina(w_n2803_62[2]),.dinb(w_n1747_0[0]),.dout(n2861),.clk(gclk));
	jand g2220(.dina(w_n2808_63[0]),.dinb(w_n1752_0[0]),.dout(n2862),.clk(gclk));
	jor g2221(.dina(n2862),.dinb(n2861),.dout(n2863),.clk(gclk));
	jnot g2222(.din(w_n2863_0[1]),.dout(n2864),.clk(gclk));
	jand g2223(.dina(w_n2864_0[1]),.dinb(w_n2860_0[1]),.dout(n2865),.clk(gclk));
	jor g2224(.dina(n2865),.dinb(w_n2857_0[1]),.dout(n2866),.clk(gclk));
	jor g2225(.dina(n2866),.dinb(n2849),.dout(n2867),.clk(gclk));
	jnot g2226(.din(w_n2867_0[1]),.dout(n2868),.clk(gclk));
	jnot g2227(.din(w_n2860_0[0]),.dout(n2869),.clk(gclk));
	jand g2228(.dina(w_n2863_0[0]),.dinb(w_n2869_0[1]),.dout(n2870),.clk(gclk));
	jand g2229(.dina(w_n1721_63[0]),.dinb(w_n1507_0[0]),.dout(n2871),.clk(gclk));
	jand g2230(.dina(w_n1562_62[1]),.dinb(w_n661_0[0]),.dout(n2872),.clk(gclk));
	jor g2231(.dina(n2872),.dinb(n2871),.dout(n2873),.clk(gclk));
	jnot g2232(.din(w_n2873_0[1]),.dout(n2874),.clk(gclk));
	jand g2233(.dina(w_n2803_62[1]),.dinb(w_n2605_0[0]),.dout(n2875),.clk(gclk));
	jand g2234(.dina(w_n2808_62[2]),.dinb(w_n1754_0[0]),.dout(n2876),.clk(gclk));
	jor g2235(.dina(n2876),.dinb(n2875),.dout(n2877),.clk(gclk));
	jand g2236(.dina(w_n2877_0[1]),.dinb(w_n2874_0[1]),.dout(n2878),.clk(gclk));
	jor g2237(.dina(n2878),.dinb(n2870),.dout(n2879),.clk(gclk));
	jand g2238(.dina(n2879),.dinb(n2868),.dout(n2880),.clk(gclk));
	jnot g2239(.din(w_n2857_0[0]),.dout(n2881),.clk(gclk));
	jnot g2240(.din(w_n2852_0[0]),.dout(n2882),.clk(gclk));
	jand g2241(.dina(w_n2855_0[0]),.dinb(w_n2882_0[1]),.dout(n2883),.clk(gclk));
	jnot g2242(.din(w_n2848_0[0]),.dout(n2884),.clk(gclk));
	jand g2243(.dina(w_n2884_0[1]),.dinb(w_n2844_0[0]),.dout(n2885),.clk(gclk));
	jor g2244(.dina(n2885),.dinb(n2883),.dout(n2886),.clk(gclk));
	jand g2245(.dina(n2886),.dinb(n2881),.dout(n2887),.clk(gclk));
	jor g2246(.dina(n2887),.dinb(n2880),.dout(n2888),.clk(gclk));
	jnot g2247(.din(w_n2888_0[1]),.dout(n2889),.clk(gclk));
	jand g2248(.dina(w_n1721_62[2]),.dinb(w_n1485_0[0]),.dout(n2890),.clk(gclk));
	jand g2249(.dina(w_n1562_62[0]),.dinb(w_n674_0[0]),.dout(n2891),.clk(gclk));
	jor g2250(.dina(n2891),.dinb(n2890),.dout(n2892),.clk(gclk));
	jnot g2251(.din(w_n2892_0[1]),.dout(n2893),.clk(gclk));
	jand g2252(.dina(w_n2803_62[0]),.dinb(w_n2583_0[0]),.dout(n2894),.clk(gclk));
	jand g2253(.dina(w_n2808_62[1]),.dinb(w_n1767_0[0]),.dout(n2895),.clk(gclk));
	jor g2254(.dina(n2895),.dinb(n2894),.dout(n2896),.clk(gclk));
	jand g2255(.dina(w_n2896_0[1]),.dinb(w_n2893_0[1]),.dout(n2897),.clk(gclk));
	jnot g2256(.din(w_n2897_0[1]),.dout(n2898),.clk(gclk));
	jand g2257(.dina(w_n2803_61[2]),.dinb(w_n1775_0[0]),.dout(n2899),.clk(gclk));
	jand g2258(.dina(w_n2808_62[0]),.dinb(w_n1793_0[0]),.dout(n2900),.clk(gclk));
	jor g2259(.dina(n2900),.dinb(n2899),.dout(n2901),.clk(gclk));
	jnot g2260(.din(w_n2901_0[1]),.dout(n2902),.clk(gclk));
	jand g2261(.dina(w_n1721_62[1]),.dinb(w_n682_0[0]),.dout(n2903),.clk(gclk));
	jand g2262(.dina(w_n1562_61[2]),.dinb(w_n700_0[0]),.dout(n2904),.clk(gclk));
	jor g2263(.dina(n2904),.dinb(n2903),.dout(n2905),.clk(gclk));
	jand g2264(.dina(w_n2905_0[1]),.dinb(w_n2902_0[1]),.dout(n2906),.clk(gclk));
	jand g2265(.dina(w_n1721_62[0]),.dinb(w_n684_0[0]),.dout(n2907),.clk(gclk));
	jand g2266(.dina(w_n1562_61[1]),.dinb(w_n698_0[0]),.dout(n2908),.clk(gclk));
	jor g2267(.dina(n2908),.dinb(n2907),.dout(n2909),.clk(gclk));
	jand g2268(.dina(w_n2803_61[1]),.dinb(w_n1777_0[0]),.dout(n2910),.clk(gclk));
	jand g2269(.dina(w_n2808_61[2]),.dinb(w_n1791_0[0]),.dout(n2911),.clk(gclk));
	jor g2270(.dina(n2911),.dinb(n2910),.dout(n2912),.clk(gclk));
	jnot g2271(.din(w_n2912_0[1]),.dout(n2913),.clk(gclk));
	jand g2272(.dina(w_n2913_0[1]),.dinb(w_n2909_0[1]),.dout(n2914),.clk(gclk));
	jand g2273(.dina(w_n1721_61[2]),.dinb(w_n686_0[0]),.dout(n2915),.clk(gclk));
	jand g2274(.dina(w_n1562_61[0]),.dinb(w_n691_0[0]),.dout(n2916),.clk(gclk));
	jor g2275(.dina(n2916),.dinb(n2915),.dout(n2917),.clk(gclk));
	jand g2276(.dina(w_n2803_61[0]),.dinb(w_n1779_0[0]),.dout(n2918),.clk(gclk));
	jand g2277(.dina(w_n2808_61[1]),.dinb(w_n1784_0[0]),.dout(n2919),.clk(gclk));
	jor g2278(.dina(n2919),.dinb(n2918),.dout(n2920),.clk(gclk));
	jnot g2279(.din(w_n2920_0[1]),.dout(n2921),.clk(gclk));
	jand g2280(.dina(w_n2921_0[1]),.dinb(w_n2917_0[1]),.dout(n2922),.clk(gclk));
	jor g2281(.dina(n2922),.dinb(w_n2914_0[1]),.dout(n2923),.clk(gclk));
	jor g2282(.dina(n2923),.dinb(n2906),.dout(n2924),.clk(gclk));
	jnot g2283(.din(w_n2924_0[1]),.dout(n2925),.clk(gclk));
	jnot g2284(.din(w_n2917_0[0]),.dout(n2926),.clk(gclk));
	jand g2285(.dina(w_n2920_0[0]),.dinb(w_n2926_0[1]),.dout(n2927),.clk(gclk));
	jand g2286(.dina(w_n1721_61[1]),.dinb(w_n1480_0[0]),.dout(n2928),.clk(gclk));
	jand g2287(.dina(w_n1562_60[2]),.dinb(w_n693_0[0]),.dout(n2929),.clk(gclk));
	jor g2288(.dina(n2929),.dinb(n2928),.dout(n2930),.clk(gclk));
	jnot g2289(.din(w_n2930_0[1]),.dout(n2931),.clk(gclk));
	jand g2290(.dina(w_n2803_60[2]),.dinb(w_n2578_0[0]),.dout(n2932),.clk(gclk));
	jand g2291(.dina(w_n2808_61[0]),.dinb(w_n1786_0[0]),.dout(n2933),.clk(gclk));
	jor g2292(.dina(n2933),.dinb(n2932),.dout(n2934),.clk(gclk));
	jand g2293(.dina(w_n2934_0[1]),.dinb(w_n2931_0[1]),.dout(n2935),.clk(gclk));
	jor g2294(.dina(n2935),.dinb(n2927),.dout(n2936),.clk(gclk));
	jand g2295(.dina(n2936),.dinb(n2925),.dout(n2937),.clk(gclk));
	jnot g2296(.din(w_n2937_0[1]),.dout(n2938),.clk(gclk));
	jnot g2297(.din(w_n2934_0[0]),.dout(n2939),.clk(gclk));
	jand g2298(.dina(w_n2939_0[1]),.dinb(w_n2930_0[0]),.dout(n2940),.clk(gclk));
	jor g2299(.dina(n2940),.dinb(w_n2924_0[0]),.dout(n2941),.clk(gclk));
	jand g2300(.dina(w_n1721_61[0]),.dinb(w_n1458_0[0]),.dout(n2942),.clk(gclk));
	jand g2301(.dina(w_n1562_60[1]),.dinb(w_n706_0[0]),.dout(n2943),.clk(gclk));
	jor g2302(.dina(n2943),.dinb(n2942),.dout(n2944),.clk(gclk));
	jand g2303(.dina(w_n2803_60[1]),.dinb(w_n2551_0[0]),.dout(n2945),.clk(gclk));
	jand g2304(.dina(w_n2808_60[2]),.dinb(w_n1799_0[0]),.dout(n2946),.clk(gclk));
	jor g2305(.dina(n2946),.dinb(n2945),.dout(n2947),.clk(gclk));
	jnot g2306(.din(w_n2947_0[1]),.dout(n2948),.clk(gclk));
	jand g2307(.dina(w_n2948_0[1]),.dinb(w_n2944_0[1]),.dout(n2949),.clk(gclk));
	jand g2308(.dina(w_n2803_60[0]),.dinb(w_n2553_0[0]),.dout(n2950),.clk(gclk));
	jand g2309(.dina(w_n2808_60[1]),.dinb(w_n2566_0[0]),.dout(n2951),.clk(gclk));
	jor g2310(.dina(n2951),.dinb(n2950),.dout(n2952),.clk(gclk));
	jnot g2311(.din(w_n2952_0[1]),.dout(n2953),.clk(gclk));
	jand g2312(.dina(w_n1721_60[2]),.dinb(w_n1460_0[0]),.dout(n2954),.clk(gclk));
	jand g2313(.dina(w_n1562_60[0]),.dinb(w_n1468_0[0]),.dout(n2955),.clk(gclk));
	jor g2314(.dina(n2955),.dinb(n2954),.dout(n2956),.clk(gclk));
	jand g2315(.dina(w_n2956_0[1]),.dinb(w_n2953_0[1]),.dout(n2957),.clk(gclk));
	jor g2316(.dina(n2957),.dinb(n2949),.dout(n2958),.clk(gclk));
	jand g2317(.dina(w_n1721_60[1]),.dinb(w_n711_0[0]),.dout(n2959),.clk(gclk));
	jand g2318(.dina(w_n1562_59[2]),.dinb(w_n1466_0[0]),.dout(n2960),.clk(gclk));
	jor g2319(.dina(n2960),.dinb(n2959),.dout(n2961),.clk(gclk));
	jand g2320(.dina(w_n2803_59[2]),.dinb(w_n2558_0[0]),.dout(n2962),.clk(gclk));
	jand g2321(.dina(w_n2808_60[0]),.dinb(w_n2564_0[0]),.dout(n2963),.clk(gclk));
	jor g2322(.dina(n2963),.dinb(n2962),.dout(n2964),.clk(gclk));
	jnot g2323(.din(w_n2964_0[1]),.dout(n2965),.clk(gclk));
	jand g2324(.dina(w_n2965_0[1]),.dinb(w_n2961_0[1]),.dout(n2966),.clk(gclk));
	jand g2325(.dina(w_n2803_59[1]),.dinb(w_n2556_0[0]),.dout(n2967),.clk(gclk));
	jand g2326(.dina(w_n2808_59[2]),.dinb(w_n2570_0[0]),.dout(n2968),.clk(gclk));
	jor g2327(.dina(n2968),.dinb(n2967),.dout(n2969),.clk(gclk));
	jnot g2328(.din(w_n2969_0[1]),.dout(n2970),.clk(gclk));
	jand g2329(.dina(w_n1721_60[0]),.dinb(w_n709_0[0]),.dout(n2971),.clk(gclk));
	jand g2330(.dina(w_n1562_59[1]),.dinb(w_n1472_0[0]),.dout(n2972),.clk(gclk));
	jor g2331(.dina(n2972),.dinb(n2971),.dout(n2973),.clk(gclk));
	jand g2332(.dina(w_n2973_0[1]),.dinb(w_n2970_0[1]),.dout(n2974),.clk(gclk));
	jor g2333(.dina(n2974),.dinb(w_n2966_0[1]),.dout(n2975),.clk(gclk));
	jor g2334(.dina(n2975),.dinb(w_n2958_0[1]),.dout(n2976),.clk(gclk));
	jand g2335(.dina(w_n1721_59[2]),.dinb(w_n1453_0[0]),.dout(n2977),.clk(gclk));
	jand g2336(.dina(w_n1562_59[0]),.dinb(w_n725_0[0]),.dout(n2978),.clk(gclk));
	jor g2337(.dina(n2978),.dinb(n2977),.dout(n2979),.clk(gclk));
	jand g2338(.dina(w_n2803_59[0]),.dinb(w_n2546_0[0]),.dout(n2980),.clk(gclk));
	jand g2339(.dina(w_n2808_59[1]),.dinb(w_n1813_0[0]),.dout(n2981),.clk(gclk));
	jor g2340(.dina(n2981),.dinb(n2980),.dout(n2982),.clk(gclk));
	jnot g2341(.din(w_n2982_0[1]),.dout(n2983),.clk(gclk));
	jand g2342(.dina(w_n2983_0[1]),.dinb(w_n2979_0[1]),.dout(n2984),.clk(gclk));
	jand g2343(.dina(w_n2803_58[2]),.dinb(w_n1802_0[0]),.dout(n2985),.clk(gclk));
	jand g2344(.dina(w_n2808_59[0]),.dinb(w_n1820_0[0]),.dout(n2986),.clk(gclk));
	jor g2345(.dina(n2986),.dinb(n2985),.dout(n2987),.clk(gclk));
	jnot g2346(.din(w_n2987_0[1]),.dout(n2988),.clk(gclk));
	jand g2347(.dina(w_n1721_59[1]),.dinb(w_n714_0[0]),.dout(n2989),.clk(gclk));
	jand g2348(.dina(w_n1562_58[2]),.dinb(w_n732_0[0]),.dout(n2990),.clk(gclk));
	jor g2349(.dina(n2990),.dinb(n2989),.dout(n2991),.clk(gclk));
	jand g2350(.dina(w_n2991_0[1]),.dinb(w_n2988_0[1]),.dout(n2992),.clk(gclk));
	jand g2351(.dina(w_n1721_59[0]),.dinb(w_n716_0[0]),.dout(n2993),.clk(gclk));
	jand g2352(.dina(w_n1562_58[1]),.dinb(w_n730_0[0]),.dout(n2994),.clk(gclk));
	jor g2353(.dina(n2994),.dinb(n2993),.dout(n2995),.clk(gclk));
	jand g2354(.dina(w_n2803_58[1]),.dinb(w_n1804_0[0]),.dout(n2996),.clk(gclk));
	jand g2355(.dina(w_n2808_58[2]),.dinb(w_n1818_0[0]),.dout(n2997),.clk(gclk));
	jor g2356(.dina(n2997),.dinb(n2996),.dout(n2998),.clk(gclk));
	jnot g2357(.din(w_n2998_0[1]),.dout(n2999),.clk(gclk));
	jand g2358(.dina(w_n2999_0[1]),.dinb(w_n2995_0[1]),.dout(n3000),.clk(gclk));
	jand g2359(.dina(w_n1721_58[2]),.dinb(w_n718_0[0]),.dout(n3001),.clk(gclk));
	jand g2360(.dina(w_n1562_58[0]),.dinb(w_n723_0[0]),.dout(n3002),.clk(gclk));
	jor g2361(.dina(n3002),.dinb(n3001),.dout(n3003),.clk(gclk));
	jand g2362(.dina(w_n2803_58[0]),.dinb(w_n1806_0[0]),.dout(n3004),.clk(gclk));
	jand g2363(.dina(w_n2808_58[1]),.dinb(w_n1811_0[0]),.dout(n3005),.clk(gclk));
	jor g2364(.dina(n3005),.dinb(n3004),.dout(n3006),.clk(gclk));
	jnot g2365(.din(w_n3006_0[1]),.dout(n3007),.clk(gclk));
	jand g2366(.dina(w_n3007_0[1]),.dinb(w_n3003_0[1]),.dout(n3008),.clk(gclk));
	jor g2367(.dina(n3008),.dinb(w_n3000_0[1]),.dout(n3009),.clk(gclk));
	jor g2368(.dina(n3009),.dinb(n2992),.dout(n3010),.clk(gclk));
	jor g2369(.dina(w_n3010_0[1]),.dinb(n2984),.dout(n3011),.clk(gclk));
	jand g2370(.dina(w_n1721_58[1]),.dinb(w_n1431_0[0]),.dout(n3012),.clk(gclk));
	jand g2371(.dina(w_n1562_57[2]),.dinb(w_n738_0[0]),.dout(n3013),.clk(gclk));
	jor g2372(.dina(n3013),.dinb(n3012),.dout(n3014),.clk(gclk));
	jand g2373(.dina(w_n2803_57[2]),.dinb(w_n2524_0[0]),.dout(n3015),.clk(gclk));
	jand g2374(.dina(w_n2808_58[0]),.dinb(w_n1826_0[0]),.dout(n3016),.clk(gclk));
	jor g2375(.dina(n3016),.dinb(n3015),.dout(n3017),.clk(gclk));
	jnot g2376(.din(w_n3017_0[1]),.dout(n3018),.clk(gclk));
	jand g2377(.dina(w_n3018_0[1]),.dinb(w_n3014_0[1]),.dout(n3019),.clk(gclk));
	jand g2378(.dina(w_n2803_57[1]),.dinb(w_n2526_0[0]),.dout(n3020),.clk(gclk));
	jand g2379(.dina(w_n2808_57[2]),.dinb(w_n2534_0[0]),.dout(n3021),.clk(gclk));
	jor g2380(.dina(n3021),.dinb(n3020),.dout(n3022),.clk(gclk));
	jnot g2381(.din(w_n3022_0[1]),.dout(n3023),.clk(gclk));
	jand g2382(.dina(w_n1721_58[0]),.dinb(w_n1433_0[0]),.dout(n3024),.clk(gclk));
	jand g2383(.dina(w_n1562_57[1]),.dinb(w_n1441_0[0]),.dout(n3025),.clk(gclk));
	jor g2384(.dina(n3025),.dinb(n3024),.dout(n3026),.clk(gclk));
	jand g2385(.dina(w_n3026_0[1]),.dinb(w_n3023_0[1]),.dout(n3027),.clk(gclk));
	jor g2386(.dina(n3027),.dinb(n3019),.dout(n3028),.clk(gclk));
	jand g2387(.dina(w_n1721_57[2]),.dinb(w_n741_0[0]),.dout(n3029),.clk(gclk));
	jand g2388(.dina(w_n1562_57[0]),.dinb(w_n1439_0[0]),.dout(n3030),.clk(gclk));
	jor g2389(.dina(n3030),.dinb(n3029),.dout(n3031),.clk(gclk));
	jand g2390(.dina(w_n2803_57[0]),.dinb(w_n1829_0[0]),.dout(n3032),.clk(gclk));
	jand g2391(.dina(w_n2808_57[1]),.dinb(w_n2532_0[0]),.dout(n3033),.clk(gclk));
	jor g2392(.dina(n3033),.dinb(n3032),.dout(n3034),.clk(gclk));
	jnot g2393(.din(w_n3034_0[1]),.dout(n3035),.clk(gclk));
	jand g2394(.dina(w_n3035_0[1]),.dinb(w_n3031_0[1]),.dout(n3036),.clk(gclk));
	jand g2395(.dina(w_n2803_56[2]),.dinb(w_n1831_0[0]),.dout(n3037),.clk(gclk));
	jand g2396(.dina(w_n2808_57[0]),.dinb(w_n2538_0[0]),.dout(n3038),.clk(gclk));
	jor g2397(.dina(n3038),.dinb(n3037),.dout(n3039),.clk(gclk));
	jnot g2398(.din(w_n3039_0[1]),.dout(n3040),.clk(gclk));
	jand g2399(.dina(w_n1721_57[1]),.dinb(w_n743_0[0]),.dout(n3041),.clk(gclk));
	jand g2400(.dina(w_n1562_56[2]),.dinb(w_n1445_0[0]),.dout(n3042),.clk(gclk));
	jor g2401(.dina(n3042),.dinb(n3041),.dout(n3043),.clk(gclk));
	jand g2402(.dina(w_n3043_0[1]),.dinb(w_n3040_0[1]),.dout(n3044),.clk(gclk));
	jor g2403(.dina(n3044),.dinb(w_n3036_0[1]),.dout(n3045),.clk(gclk));
	jor g2404(.dina(n3045),.dinb(w_n3028_0[1]),.dout(n3046),.clk(gclk));
	jand g2405(.dina(w_n1721_57[0]),.dinb(w_n1426_0[0]),.dout(n3047),.clk(gclk));
	jand g2406(.dina(w_n1562_56[1]),.dinb(w_n757_0[0]),.dout(n3048),.clk(gclk));
	jor g2407(.dina(n3048),.dinb(n3047),.dout(n3049),.clk(gclk));
	jand g2408(.dina(w_n2803_56[1]),.dinb(w_n2519_0[0]),.dout(n3050),.clk(gclk));
	jand g2409(.dina(w_n2808_56[2]),.dinb(w_n1845_0[0]),.dout(n3051),.clk(gclk));
	jor g2410(.dina(n3051),.dinb(n3050),.dout(n3052),.clk(gclk));
	jnot g2411(.din(w_n3052_0[1]),.dout(n3053),.clk(gclk));
	jand g2412(.dina(w_n3053_0[1]),.dinb(w_n3049_0[1]),.dout(n3054),.clk(gclk));
	jand g2413(.dina(w_n2803_56[0]),.dinb(w_n1834_0[0]),.dout(n3055),.clk(gclk));
	jand g2414(.dina(w_n2808_56[1]),.dinb(w_n1852_0[0]),.dout(n3056),.clk(gclk));
	jor g2415(.dina(n3056),.dinb(n3055),.dout(n3057),.clk(gclk));
	jnot g2416(.din(w_n3057_0[1]),.dout(n3058),.clk(gclk));
	jand g2417(.dina(w_n1721_56[2]),.dinb(w_n746_0[0]),.dout(n3059),.clk(gclk));
	jand g2418(.dina(w_n1562_56[0]),.dinb(w_n764_0[0]),.dout(n3060),.clk(gclk));
	jor g2419(.dina(n3060),.dinb(n3059),.dout(n3061),.clk(gclk));
	jand g2420(.dina(w_n3061_0[1]),.dinb(w_n3058_0[1]),.dout(n3062),.clk(gclk));
	jand g2421(.dina(w_n1721_56[1]),.dinb(w_n748_0[0]),.dout(n3063),.clk(gclk));
	jand g2422(.dina(w_n1562_55[2]),.dinb(w_n762_0[0]),.dout(n3064),.clk(gclk));
	jor g2423(.dina(n3064),.dinb(n3063),.dout(n3065),.clk(gclk));
	jand g2424(.dina(w_n2803_55[2]),.dinb(w_n1836_0[0]),.dout(n3066),.clk(gclk));
	jand g2425(.dina(w_n2808_56[0]),.dinb(w_n1850_0[0]),.dout(n3067),.clk(gclk));
	jor g2426(.dina(n3067),.dinb(n3066),.dout(n3068),.clk(gclk));
	jnot g2427(.din(w_n3068_0[1]),.dout(n3069),.clk(gclk));
	jand g2428(.dina(w_n3069_0[1]),.dinb(w_n3065_0[1]),.dout(n3070),.clk(gclk));
	jand g2429(.dina(w_n1721_56[0]),.dinb(w_n750_0[0]),.dout(n3071),.clk(gclk));
	jand g2430(.dina(w_n1562_55[1]),.dinb(w_n755_0[0]),.dout(n3072),.clk(gclk));
	jor g2431(.dina(n3072),.dinb(n3071),.dout(n3073),.clk(gclk));
	jand g2432(.dina(w_n2803_55[1]),.dinb(w_n1838_0[0]),.dout(n3074),.clk(gclk));
	jand g2433(.dina(w_n2808_55[2]),.dinb(w_n1843_0[0]),.dout(n3075),.clk(gclk));
	jor g2434(.dina(n3075),.dinb(n3074),.dout(n3076),.clk(gclk));
	jnot g2435(.din(w_n3076_0[1]),.dout(n3077),.clk(gclk));
	jand g2436(.dina(w_n3077_0[1]),.dinb(w_n3073_0[1]),.dout(n3078),.clk(gclk));
	jor g2437(.dina(n3078),.dinb(w_n3070_0[1]),.dout(n3079),.clk(gclk));
	jor g2438(.dina(n3079),.dinb(n3062),.dout(n3080),.clk(gclk));
	jor g2439(.dina(w_n3080_0[1]),.dinb(n3054),.dout(n3081),.clk(gclk));
	jand g2440(.dina(w_n1721_55[2]),.dinb(w_n1399_0[0]),.dout(n3082),.clk(gclk));
	jand g2441(.dina(w_n1562_55[0]),.dinb(w_n770_0[0]),.dout(n3083),.clk(gclk));
	jor g2442(.dina(n3083),.dinb(n3082),.dout(n3084),.clk(gclk));
	jand g2443(.dina(w_n2803_55[0]),.dinb(w_n2492_0[0]),.dout(n3085),.clk(gclk));
	jand g2444(.dina(w_n2808_55[1]),.dinb(w_n1858_0[0]),.dout(n3086),.clk(gclk));
	jor g2445(.dina(n3086),.dinb(n3085),.dout(n3087),.clk(gclk));
	jnot g2446(.din(w_n3087_0[1]),.dout(n3088),.clk(gclk));
	jand g2447(.dina(w_n3088_0[1]),.dinb(w_n3084_0[1]),.dout(n3089),.clk(gclk));
	jand g2448(.dina(w_n2803_54[2]),.dinb(w_n2494_0[0]),.dout(n3090),.clk(gclk));
	jand g2449(.dina(w_n2808_55[0]),.dinb(w_n2507_0[0]),.dout(n3091),.clk(gclk));
	jor g2450(.dina(n3091),.dinb(n3090),.dout(n3092),.clk(gclk));
	jnot g2451(.din(w_n3092_0[1]),.dout(n3093),.clk(gclk));
	jand g2452(.dina(w_n1721_55[1]),.dinb(w_n1401_0[0]),.dout(n3094),.clk(gclk));
	jand g2453(.dina(w_n1562_54[2]),.dinb(w_n1414_0[0]),.dout(n3095),.clk(gclk));
	jor g2454(.dina(n3095),.dinb(n3094),.dout(n3096),.clk(gclk));
	jand g2455(.dina(w_n3096_0[1]),.dinb(w_n3093_0[1]),.dout(n3097),.clk(gclk));
	jor g2456(.dina(n3097),.dinb(n3089),.dout(n3098),.clk(gclk));
	jand g2457(.dina(w_n1721_55[0]),.dinb(w_n1406_0[0]),.dout(n3099),.clk(gclk));
	jand g2458(.dina(w_n1562_54[1]),.dinb(w_n1412_0[0]),.dout(n3100),.clk(gclk));
	jor g2459(.dina(n3100),.dinb(n3099),.dout(n3101),.clk(gclk));
	jand g2460(.dina(w_n2803_54[1]),.dinb(w_n2499_0[0]),.dout(n3102),.clk(gclk));
	jand g2461(.dina(w_n2808_54[2]),.dinb(w_n2505_0[0]),.dout(n3103),.clk(gclk));
	jor g2462(.dina(n3103),.dinb(n3102),.dout(n3104),.clk(gclk));
	jnot g2463(.din(w_n3104_0[1]),.dout(n3105),.clk(gclk));
	jand g2464(.dina(w_n3105_0[1]),.dinb(w_n3101_0[1]),.dout(n3106),.clk(gclk));
	jand g2465(.dina(w_n2803_54[0]),.dinb(w_n2497_0[0]),.dout(n3107),.clk(gclk));
	jand g2466(.dina(w_n2808_54[1]),.dinb(w_n2511_0[0]),.dout(n3108),.clk(gclk));
	jor g2467(.dina(n3108),.dinb(n3107),.dout(n3109),.clk(gclk));
	jnot g2468(.din(w_n3109_0[1]),.dout(n3110),.clk(gclk));
	jand g2469(.dina(w_n1721_54[2]),.dinb(w_n1404_0[0]),.dout(n3111),.clk(gclk));
	jand g2470(.dina(w_n1562_54[0]),.dinb(w_n1418_0[0]),.dout(n3112),.clk(gclk));
	jor g2471(.dina(n3112),.dinb(n3111),.dout(n3113),.clk(gclk));
	jand g2472(.dina(w_n3113_0[1]),.dinb(w_n3110_0[1]),.dout(n3114),.clk(gclk));
	jor g2473(.dina(n3114),.dinb(w_n3106_0[1]),.dout(n3115),.clk(gclk));
	jor g2474(.dina(n3115),.dinb(w_n3098_0[1]),.dout(n3116),.clk(gclk));
	jand g2475(.dina(w_n2803_53[2]),.dinb(w_n1861_0[0]),.dout(n3117),.clk(gclk));
	jand g2476(.dina(w_n2808_54[0]),.dinb(w_n1879_0[0]),.dout(n3118),.clk(gclk));
	jor g2477(.dina(n3118),.dinb(n3117),.dout(n3119),.clk(gclk));
	jnot g2478(.din(w_n3119_0[1]),.dout(n3120),.clk(gclk));
	jand g2479(.dina(w_n1721_54[1]),.dinb(w_n773_0[0]),.dout(n3121),.clk(gclk));
	jand g2480(.dina(w_n1562_53[2]),.dinb(w_n791_0[0]),.dout(n3122),.clk(gclk));
	jor g2481(.dina(n3122),.dinb(n3121),.dout(n3123),.clk(gclk));
	jand g2482(.dina(w_n3123_0[1]),.dinb(w_n3120_0[1]),.dout(n3124),.clk(gclk));
	jand g2483(.dina(w_n1721_54[0]),.dinb(w_n775_0[0]),.dout(n3125),.clk(gclk));
	jand g2484(.dina(w_n1562_53[1]),.dinb(w_n789_0[0]),.dout(n3126),.clk(gclk));
	jor g2485(.dina(n3126),.dinb(n3125),.dout(n3127),.clk(gclk));
	jand g2486(.dina(w_n2803_53[1]),.dinb(w_n1863_0[0]),.dout(n3128),.clk(gclk));
	jand g2487(.dina(w_n2808_53[2]),.dinb(w_n1877_0[0]),.dout(n3129),.clk(gclk));
	jor g2488(.dina(n3129),.dinb(n3128),.dout(n3130),.clk(gclk));
	jnot g2489(.din(w_n3130_0[1]),.dout(n3131),.clk(gclk));
	jand g2490(.dina(w_n3131_0[1]),.dinb(w_n3127_0[1]),.dout(n3132),.clk(gclk));
	jand g2491(.dina(w_n1721_53[2]),.dinb(w_n777_0[0]),.dout(n3133),.clk(gclk));
	jand g2492(.dina(w_n1562_53[0]),.dinb(w_n782_0[0]),.dout(n3134),.clk(gclk));
	jor g2493(.dina(n3134),.dinb(n3133),.dout(n3135),.clk(gclk));
	jand g2494(.dina(w_n2803_53[0]),.dinb(w_n1865_0[0]),.dout(n3136),.clk(gclk));
	jand g2495(.dina(w_n2808_53[1]),.dinb(w_n1870_0[0]),.dout(n3137),.clk(gclk));
	jor g2496(.dina(n3137),.dinb(n3136),.dout(n3138),.clk(gclk));
	jnot g2497(.din(w_n3138_0[1]),.dout(n3139),.clk(gclk));
	jand g2498(.dina(w_n3139_0[1]),.dinb(w_n3135_0[1]),.dout(n3140),.clk(gclk));
	jor g2499(.dina(n3140),.dinb(w_n3132_0[1]),.dout(n3141),.clk(gclk));
	jor g2500(.dina(n3141),.dinb(n3124),.dout(n3142),.clk(gclk));
	jnot g2501(.din(w_n3142_0[1]),.dout(n3143),.clk(gclk));
	jnot g2502(.din(w_n3135_0[0]),.dout(n3144),.clk(gclk));
	jand g2503(.dina(w_n3138_0[0]),.dinb(w_n3144_0[1]),.dout(n3145),.clk(gclk));
	jand g2504(.dina(w_n1721_53[1]),.dinb(w_n1394_0[0]),.dout(n3146),.clk(gclk));
	jand g2505(.dina(w_n1562_52[2]),.dinb(w_n784_0[0]),.dout(n3147),.clk(gclk));
	jor g2506(.dina(n3147),.dinb(n3146),.dout(n3148),.clk(gclk));
	jnot g2507(.din(w_n3148_0[1]),.dout(n3149),.clk(gclk));
	jand g2508(.dina(w_n2803_52[2]),.dinb(w_n2487_0[0]),.dout(n3150),.clk(gclk));
	jand g2509(.dina(w_n2808_53[0]),.dinb(w_n1872_0[0]),.dout(n3151),.clk(gclk));
	jor g2510(.dina(n3151),.dinb(n3150),.dout(n3152),.clk(gclk));
	jand g2511(.dina(w_n3152_0[1]),.dinb(w_n3149_0[1]),.dout(n3153),.clk(gclk));
	jor g2512(.dina(n3153),.dinb(n3145),.dout(n3154),.clk(gclk));
	jand g2513(.dina(n3154),.dinb(n3143),.dout(n3155),.clk(gclk));
	jnot g2514(.din(w_n3155_0[1]),.dout(n3156),.clk(gclk));
	jnot g2515(.din(w_n3132_0[0]),.dout(n3157),.clk(gclk));
	jnot g2516(.din(w_n3127_0[0]),.dout(n3158),.clk(gclk));
	jand g2517(.dina(w_n3130_0[0]),.dinb(w_n3158_0[1]),.dout(n3159),.clk(gclk));
	jnot g2518(.din(w_n3123_0[0]),.dout(n3160),.clk(gclk));
	jand g2519(.dina(w_n3160_0[1]),.dinb(w_n3119_0[0]),.dout(n3161),.clk(gclk));
	jor g2520(.dina(n3161),.dinb(n3159),.dout(n3162),.clk(gclk));
	jand g2521(.dina(n3162),.dinb(n3157),.dout(n3163),.clk(gclk));
	jnot g2522(.din(w_n3163_0[1]),.dout(n3164),.clk(gclk));
	jand g2523(.dina(w_n1721_53[0]),.dinb(w_n1372_0[0]),.dout(n3165),.clk(gclk));
	jand g2524(.dina(w_n1562_52[1]),.dinb(w_n797_0[0]),.dout(n3166),.clk(gclk));
	jor g2525(.dina(n3166),.dinb(n3165),.dout(n3167),.clk(gclk));
	jnot g2526(.din(w_n3167_0[1]),.dout(n3168),.clk(gclk));
	jand g2527(.dina(w_n2803_52[1]),.dinb(w_n2465_0[0]),.dout(n3169),.clk(gclk));
	jand g2528(.dina(w_n2808_52[2]),.dinb(w_n1885_0[0]),.dout(n3170),.clk(gclk));
	jor g2529(.dina(n3170),.dinb(n3169),.dout(n3171),.clk(gclk));
	jand g2530(.dina(w_n3171_0[1]),.dinb(w_n3168_0[1]),.dout(n3172),.clk(gclk));
	jnot g2531(.din(w_n3172_0[1]),.dout(n3173),.clk(gclk));
	jnot g2532(.din(w_n3171_0[0]),.dout(n3174),.clk(gclk));
	jand g2533(.dina(w_n3174_0[1]),.dinb(w_n3167_0[0]),.dout(n3175),.clk(gclk));
	jand g2534(.dina(w_n2803_52[0]),.dinb(w_n2467_0[0]),.dout(n3176),.clk(gclk));
	jand g2535(.dina(w_n2808_52[1]),.dinb(w_n2475_0[0]),.dout(n3177),.clk(gclk));
	jor g2536(.dina(n3177),.dinb(n3176),.dout(n3178),.clk(gclk));
	jnot g2537(.din(w_n3178_0[1]),.dout(n3179),.clk(gclk));
	jand g2538(.dina(w_n1721_52[2]),.dinb(w_n1374_0[0]),.dout(n3180),.clk(gclk));
	jand g2539(.dina(w_n1562_52[0]),.dinb(w_n1382_0[0]),.dout(n3181),.clk(gclk));
	jor g2540(.dina(n3181),.dinb(n3180),.dout(n3182),.clk(gclk));
	jand g2541(.dina(w_n3182_0[1]),.dinb(w_n3179_0[1]),.dout(n3183),.clk(gclk));
	jor g2542(.dina(n3183),.dinb(n3175),.dout(n3184),.clk(gclk));
	jand g2543(.dina(w_n1721_52[1]),.dinb(w_n800_0[0]),.dout(n3185),.clk(gclk));
	jand g2544(.dina(w_n1562_51[2]),.dinb(w_n1380_0[0]),.dout(n3186),.clk(gclk));
	jor g2545(.dina(n3186),.dinb(n3185),.dout(n3187),.clk(gclk));
	jand g2546(.dina(w_n2803_51[2]),.dinb(w_n1888_0[0]),.dout(n3188),.clk(gclk));
	jand g2547(.dina(w_n2808_52[0]),.dinb(w_n2473_0[0]),.dout(n3189),.clk(gclk));
	jor g2548(.dina(n3189),.dinb(n3188),.dout(n3190),.clk(gclk));
	jnot g2549(.din(w_n3190_0[1]),.dout(n3191),.clk(gclk));
	jand g2550(.dina(w_n3191_0[1]),.dinb(w_n3187_0[1]),.dout(n3192),.clk(gclk));
	jand g2551(.dina(w_n2803_51[1]),.dinb(w_n1890_0[0]),.dout(n3193),.clk(gclk));
	jand g2552(.dina(w_n2808_51[2]),.dinb(w_n2479_0[0]),.dout(n3194),.clk(gclk));
	jor g2553(.dina(n3194),.dinb(n3193),.dout(n3195),.clk(gclk));
	jnot g2554(.din(w_n3195_0[1]),.dout(n3196),.clk(gclk));
	jand g2555(.dina(w_n1721_52[0]),.dinb(w_n802_0[0]),.dout(n3197),.clk(gclk));
	jand g2556(.dina(w_n1562_51[1]),.dinb(w_n1386_0[0]),.dout(n3198),.clk(gclk));
	jor g2557(.dina(n3198),.dinb(n3197),.dout(n3199),.clk(gclk));
	jand g2558(.dina(w_n3199_0[1]),.dinb(w_n3196_0[1]),.dout(n3200),.clk(gclk));
	jor g2559(.dina(n3200),.dinb(w_n3192_0[1]),.dout(n3201),.clk(gclk));
	jor g2560(.dina(n3201),.dinb(w_n3184_0[1]),.dout(n3202),.clk(gclk));
	jand g2561(.dina(w_n1721_51[2]),.dinb(w_n1367_0[0]),.dout(n3203),.clk(gclk));
	jand g2562(.dina(w_n1562_51[0]),.dinb(w_n816_0[0]),.dout(n3204),.clk(gclk));
	jor g2563(.dina(n3204),.dinb(n3203),.dout(n3205),.clk(gclk));
	jand g2564(.dina(w_n2803_51[0]),.dinb(w_n2460_0[0]),.dout(n3206),.clk(gclk));
	jand g2565(.dina(w_n2808_51[1]),.dinb(w_n1904_0[0]),.dout(n3207),.clk(gclk));
	jor g2566(.dina(n3207),.dinb(n3206),.dout(n3208),.clk(gclk));
	jnot g2567(.din(w_n3208_0[1]),.dout(n3209),.clk(gclk));
	jand g2568(.dina(w_n3209_0[1]),.dinb(w_n3205_0[1]),.dout(n3210),.clk(gclk));
	jand g2569(.dina(w_n2803_50[2]),.dinb(w_n1893_0[0]),.dout(n3211),.clk(gclk));
	jand g2570(.dina(w_n2808_51[0]),.dinb(w_n1911_0[0]),.dout(n3212),.clk(gclk));
	jor g2571(.dina(n3212),.dinb(n3211),.dout(n3213),.clk(gclk));
	jnot g2572(.din(w_n3213_0[1]),.dout(n3214),.clk(gclk));
	jand g2573(.dina(w_n1721_51[1]),.dinb(w_n805_0[0]),.dout(n3215),.clk(gclk));
	jand g2574(.dina(w_n1562_50[2]),.dinb(w_n823_0[0]),.dout(n3216),.clk(gclk));
	jor g2575(.dina(n3216),.dinb(n3215),.dout(n3217),.clk(gclk));
	jand g2576(.dina(w_n3217_0[1]),.dinb(w_n3214_0[1]),.dout(n3218),.clk(gclk));
	jand g2577(.dina(w_n1721_51[0]),.dinb(w_n807_0[0]),.dout(n3219),.clk(gclk));
	jand g2578(.dina(w_n1562_50[1]),.dinb(w_n821_0[0]),.dout(n3220),.clk(gclk));
	jor g2579(.dina(n3220),.dinb(n3219),.dout(n3221),.clk(gclk));
	jand g2580(.dina(w_n2803_50[1]),.dinb(w_n1895_0[0]),.dout(n3222),.clk(gclk));
	jand g2581(.dina(w_n2808_50[2]),.dinb(w_n1909_0[0]),.dout(n3223),.clk(gclk));
	jor g2582(.dina(n3223),.dinb(n3222),.dout(n3224),.clk(gclk));
	jnot g2583(.din(w_n3224_0[1]),.dout(n3225),.clk(gclk));
	jand g2584(.dina(w_n3225_0[1]),.dinb(w_n3221_0[1]),.dout(n3226),.clk(gclk));
	jand g2585(.dina(w_n1721_50[2]),.dinb(w_n809_0[0]),.dout(n3227),.clk(gclk));
	jand g2586(.dina(w_n1562_50[0]),.dinb(w_n814_0[0]),.dout(n3228),.clk(gclk));
	jor g2587(.dina(n3228),.dinb(n3227),.dout(n3229),.clk(gclk));
	jand g2588(.dina(w_n2803_50[0]),.dinb(w_n1897_0[0]),.dout(n3230),.clk(gclk));
	jand g2589(.dina(w_n2808_50[1]),.dinb(w_n1902_0[0]),.dout(n3231),.clk(gclk));
	jor g2590(.dina(n3231),.dinb(n3230),.dout(n3232),.clk(gclk));
	jnot g2591(.din(w_n3232_0[1]),.dout(n3233),.clk(gclk));
	jand g2592(.dina(w_n3233_0[1]),.dinb(w_n3229_0[1]),.dout(n3234),.clk(gclk));
	jor g2593(.dina(n3234),.dinb(w_n3226_0[1]),.dout(n3235),.clk(gclk));
	jor g2594(.dina(n3235),.dinb(n3218),.dout(n3236),.clk(gclk));
	jor g2595(.dina(w_n3236_0[1]),.dinb(n3210),.dout(n3237),.clk(gclk));
	jand g2596(.dina(w_n2803_49[2]),.dinb(w_n1920_0[0]),.dout(n3238),.clk(gclk));
	jand g2597(.dina(w_n2808_50[0]),.dinb(w_n1938_0[0]),.dout(n3239),.clk(gclk));
	jor g2598(.dina(n3239),.dinb(n3238),.dout(n3240),.clk(gclk));
	jnot g2599(.din(w_n3240_0[1]),.dout(n3241),.clk(gclk));
	jand g2600(.dina(w_n1721_50[1]),.dinb(w_n837_0[0]),.dout(n3242),.clk(gclk));
	jand g2601(.dina(w_n1562_49[2]),.dinb(w_n855_0[0]),.dout(n3243),.clk(gclk));
	jor g2602(.dina(n3243),.dinb(n3242),.dout(n3244),.clk(gclk));
	jand g2603(.dina(w_n3244_0[1]),.dinb(w_n3241_0[1]),.dout(n3245),.clk(gclk));
	jand g2604(.dina(w_n1721_50[0]),.dinb(w_n839_0[0]),.dout(n3246),.clk(gclk));
	jand g2605(.dina(w_n1562_49[1]),.dinb(w_n853_0[0]),.dout(n3247),.clk(gclk));
	jor g2606(.dina(n3247),.dinb(n3246),.dout(n3248),.clk(gclk));
	jand g2607(.dina(w_n2803_49[1]),.dinb(w_n1922_0[0]),.dout(n3249),.clk(gclk));
	jand g2608(.dina(w_n2808_49[2]),.dinb(w_n1936_0[0]),.dout(n3250),.clk(gclk));
	jor g2609(.dina(n3250),.dinb(n3249),.dout(n3251),.clk(gclk));
	jnot g2610(.din(w_n3251_0[1]),.dout(n3252),.clk(gclk));
	jand g2611(.dina(w_n3252_0[1]),.dinb(w_n3248_0[1]),.dout(n3253),.clk(gclk));
	jand g2612(.dina(w_n1721_49[2]),.dinb(w_n841_0[0]),.dout(n3254),.clk(gclk));
	jand g2613(.dina(w_n1562_49[0]),.dinb(w_n846_0[0]),.dout(n3255),.clk(gclk));
	jor g2614(.dina(n3255),.dinb(n3254),.dout(n3256),.clk(gclk));
	jand g2615(.dina(w_n2803_49[0]),.dinb(w_n1924_0[0]),.dout(n3257),.clk(gclk));
	jand g2616(.dina(w_n2808_49[1]),.dinb(w_n1929_0[0]),.dout(n3258),.clk(gclk));
	jor g2617(.dina(n3258),.dinb(n3257),.dout(n3259),.clk(gclk));
	jnot g2618(.din(w_n3259_0[1]),.dout(n3260),.clk(gclk));
	jand g2619(.dina(w_n3260_0[1]),.dinb(w_n3256_0[1]),.dout(n3261),.clk(gclk));
	jor g2620(.dina(n3261),.dinb(w_n3253_0[1]),.dout(n3262),.clk(gclk));
	jor g2621(.dina(n3262),.dinb(n3245),.dout(n3263),.clk(gclk));
	jnot g2622(.din(w_n3263_0[1]),.dout(n3264),.clk(gclk));
	jnot g2623(.din(w_n3256_0[0]),.dout(n3265),.clk(gclk));
	jand g2624(.dina(w_n3259_0[0]),.dinb(w_n3265_0[1]),.dout(n3266),.clk(gclk));
	jand g2625(.dina(w_n1721_49[1]),.dinb(w_n1340_0[0]),.dout(n3267),.clk(gclk));
	jand g2626(.dina(w_n1562_48[2]),.dinb(w_n848_0[0]),.dout(n3268),.clk(gclk));
	jor g2627(.dina(n3268),.dinb(n3267),.dout(n3269),.clk(gclk));
	jnot g2628(.din(w_n3269_0[1]),.dout(n3270),.clk(gclk));
	jand g2629(.dina(w_n2803_48[2]),.dinb(w_n2428_0[0]),.dout(n3271),.clk(gclk));
	jand g2630(.dina(w_n2808_49[0]),.dinb(w_n1931_0[0]),.dout(n3272),.clk(gclk));
	jor g2631(.dina(n3272),.dinb(n3271),.dout(n3273),.clk(gclk));
	jand g2632(.dina(w_n3273_0[1]),.dinb(w_n3270_0[1]),.dout(n3274),.clk(gclk));
	jor g2633(.dina(n3274),.dinb(n3266),.dout(n3275),.clk(gclk));
	jand g2634(.dina(n3275),.dinb(n3264),.dout(n3276),.clk(gclk));
	jnot g2635(.din(w_n3253_0[0]),.dout(n3277),.clk(gclk));
	jnot g2636(.din(w_n3248_0[0]),.dout(n3278),.clk(gclk));
	jand g2637(.dina(w_n3251_0[0]),.dinb(w_n3278_0[1]),.dout(n3279),.clk(gclk));
	jnot g2638(.din(w_n3244_0[0]),.dout(n3280),.clk(gclk));
	jand g2639(.dina(w_n3280_0[1]),.dinb(w_n3240_0[0]),.dout(n3281),.clk(gclk));
	jor g2640(.dina(n3281),.dinb(n3279),.dout(n3282),.clk(gclk));
	jand g2641(.dina(n3282),.dinb(n3277),.dout(n3283),.clk(gclk));
	jor g2642(.dina(n3283),.dinb(n3276),.dout(n3284),.clk(gclk));
	jnot g2643(.din(w_n3284_0[1]),.dout(n3285),.clk(gclk));
	jand g2644(.dina(w_n1721_49[0]),.dinb(w_n1333_0[0]),.dout(n3286),.clk(gclk));
	jand g2645(.dina(w_n1562_48[1]),.dinb(w_n861_0[0]),.dout(n3287),.clk(gclk));
	jor g2646(.dina(n3287),.dinb(n3286),.dout(n3288),.clk(gclk));
	jnot g2647(.din(w_n3288_0[1]),.dout(n3289),.clk(gclk));
	jand g2648(.dina(w_n2803_48[1]),.dinb(w_n2421_0[0]),.dout(n3290),.clk(gclk));
	jand g2649(.dina(w_n2808_48[2]),.dinb(w_n1944_0[0]),.dout(n3291),.clk(gclk));
	jor g2650(.dina(n3291),.dinb(n3290),.dout(n3292),.clk(gclk));
	jand g2651(.dina(w_n3292_0[1]),.dinb(w_n3289_0[1]),.dout(n3293),.clk(gclk));
	jnot g2652(.din(w_n3293_0[1]),.dout(n3294),.clk(gclk));
	jand g2653(.dina(w_n2803_48[0]),.dinb(w_n2423_0[0]),.dout(n3295),.clk(gclk));
	jand g2654(.dina(w_n2808_48[1]),.dinb(w_n1953_0[0]),.dout(n3296),.clk(gclk));
	jor g2655(.dina(n3296),.dinb(n3295),.dout(n3297),.clk(gclk));
	jand g2656(.dina(w_n1721_48[2]),.dinb(w_n1335_0[0]),.dout(n3298),.clk(gclk));
	jand g2657(.dina(w_n1562_48[0]),.dinb(w_n870_0[0]),.dout(n3299),.clk(gclk));
	jor g2658(.dina(n3299),.dinb(n3298),.dout(n3300),.clk(gclk));
	jnot g2659(.din(w_n3300_0[1]),.dout(n3301),.clk(gclk));
	jand g2660(.dina(w_n3301_0[1]),.dinb(w_n3297_0[1]),.dout(n3302),.clk(gclk));
	jand g2661(.dina(w_n1721_48[1]),.dinb(w_n864_0[0]),.dout(n3303),.clk(gclk));
	jand g2662(.dina(w_n1562_47[2]),.dinb(w_n872_0[0]),.dout(n3304),.clk(gclk));
	jor g2663(.dina(n3304),.dinb(n3303),.dout(n3305),.clk(gclk));
	jnot g2664(.din(w_n3305_0[1]),.dout(n3306),.clk(gclk));
	jand g2665(.dina(w_n2803_47[2]),.dinb(w_n1947_0[0]),.dout(n3307),.clk(gclk));
	jand g2666(.dina(w_n2808_48[0]),.dinb(w_n1955_0[0]),.dout(n3308),.clk(gclk));
	jor g2667(.dina(n3308),.dinb(n3307),.dout(n3309),.clk(gclk));
	jand g2668(.dina(w_n3309_0[1]),.dinb(w_n3306_0[1]),.dout(n3310),.clk(gclk));
	jnot g2669(.din(w_n3309_0[0]),.dout(n3311),.clk(gclk));
	jand g2670(.dina(w_n3311_0[1]),.dinb(w_n3305_0[0]),.dout(n3312),.clk(gclk));
	jnot g2671(.din(w_n3312_0[1]),.dout(n3313),.clk(gclk));
	jand g2672(.dina(w_n2803_47[1]),.dinb(w_n2416_0[0]),.dout(n3314),.clk(gclk));
	jand g2673(.dina(w_n2808_47[2]),.dinb(w_n1950_0[0]),.dout(n3315),.clk(gclk));
	jor g2674(.dina(n3315),.dinb(n3314),.dout(n3316),.clk(gclk));
	jand g2675(.dina(w_n1721_48[0]),.dinb(w_n1328_0[0]),.dout(n3317),.clk(gclk));
	jand g2676(.dina(w_n1562_47[1]),.dinb(w_n867_0[0]),.dout(n3318),.clk(gclk));
	jor g2677(.dina(n3318),.dinb(n3317),.dout(n3319),.clk(gclk));
	jnot g2678(.din(w_n3319_0[1]),.dout(n3320),.clk(gclk));
	jand g2679(.dina(w_n3320_0[1]),.dinb(w_n3316_0[1]),.dout(n3321),.clk(gclk));
	jand g2680(.dina(n3321),.dinb(n3313),.dout(n3322),.clk(gclk));
	jor g2681(.dina(n3322),.dinb(n3310),.dout(n3323),.clk(gclk));
	jor g2682(.dina(n3323),.dinb(n3302),.dout(n3324),.clk(gclk));
	jnot g2683(.din(w_n3324_0[1]),.dout(n3325),.clk(gclk));
	jand g2684(.dina(w_n1721_47[2]),.dinb(w_n878_0[0]),.dout(n3326),.clk(gclk));
	jand g2685(.dina(w_n1562_47[0]),.dinb(w_n1312_0[0]),.dout(n3327),.clk(gclk));
	jor g2686(.dina(n3327),.dinb(n3326),.dout(n3328),.clk(gclk));
	jand g2687(.dina(w_n2803_47[0]),.dinb(w_n1961_0[0]),.dout(n3329),.clk(gclk));
	jand g2688(.dina(w_n2808_47[1]),.dinb(w_n2400_0[0]),.dout(n3330),.clk(gclk));
	jor g2689(.dina(n3330),.dinb(n3329),.dout(n3331),.clk(gclk));
	jnot g2690(.din(w_n3331_0[1]),.dout(n3332),.clk(gclk));
	jand g2691(.dina(w_n3332_0[1]),.dinb(w_n3328_0[1]),.dout(n3333),.clk(gclk));
	jand g2692(.dina(w_n2803_46[2]),.dinb(w_n1967_0[0]),.dout(n3334),.clk(gclk));
	jand g2693(.dina(w_n2808_47[0]),.dinb(w_n2407_0[0]),.dout(n3335),.clk(gclk));
	jor g2694(.dina(n3335),.dinb(n3334),.dout(n3336),.clk(gclk));
	jnot g2695(.din(w_n3336_0[1]),.dout(n3337),.clk(gclk));
	jand g2696(.dina(w_n1721_47[1]),.dinb(w_n884_0[0]),.dout(n3338),.clk(gclk));
	jand g2697(.dina(w_n1562_46[2]),.dinb(w_n1319_0[0]),.dout(n3339),.clk(gclk));
	jor g2698(.dina(n3339),.dinb(n3338),.dout(n3340),.clk(gclk));
	jand g2699(.dina(w_n3340_0[1]),.dinb(w_n3337_0[1]),.dout(n3341),.clk(gclk));
	jand g2700(.dina(w_n1721_47[0]),.dinb(w_n880_0[0]),.dout(n3342),.clk(gclk));
	jand g2701(.dina(w_n1562_46[1]),.dinb(w_n1317_0[0]),.dout(n3343),.clk(gclk));
	jor g2702(.dina(n3343),.dinb(n3342),.dout(n3344),.clk(gclk));
	jand g2703(.dina(w_n2803_46[1]),.dinb(w_n1963_0[0]),.dout(n3345),.clk(gclk));
	jand g2704(.dina(w_n2808_46[2]),.dinb(w_n2405_0[0]),.dout(n3346),.clk(gclk));
	jor g2705(.dina(n3346),.dinb(n3345),.dout(n3347),.clk(gclk));
	jnot g2706(.din(w_n3347_0[1]),.dout(n3348),.clk(gclk));
	jand g2707(.dina(w_n3348_0[1]),.dinb(w_n3344_0[1]),.dout(n3349),.clk(gclk));
	jand g2708(.dina(w_n1721_46[2]),.dinb(w_n882_0[0]),.dout(n3350),.clk(gclk));
	jand g2709(.dina(w_n1562_46[0]),.dinb(w_n1310_0[0]),.dout(n3351),.clk(gclk));
	jor g2710(.dina(n3351),.dinb(n3350),.dout(n3352),.clk(gclk));
	jand g2711(.dina(w_n2803_46[0]),.dinb(w_n1965_0[0]),.dout(n3353),.clk(gclk));
	jand g2712(.dina(w_n2808_46[1]),.dinb(w_n2398_0[0]),.dout(n3354),.clk(gclk));
	jor g2713(.dina(n3354),.dinb(n3353),.dout(n3355),.clk(gclk));
	jnot g2714(.din(w_n3355_0[1]),.dout(n3356),.clk(gclk));
	jand g2715(.dina(w_n3356_0[1]),.dinb(w_n3352_0[1]),.dout(n3357),.clk(gclk));
	jor g2716(.dina(n3357),.dinb(w_n3349_0[1]),.dout(n3358),.clk(gclk));
	jor g2717(.dina(n3358),.dinb(n3341),.dout(n3359),.clk(gclk));
	jor g2718(.dina(w_n3359_0[1]),.dinb(n3333),.dout(n3360),.clk(gclk));
	jnot g2719(.din(w_n3360_0[1]),.dout(n3361),.clk(gclk));
	jand g2720(.dina(w_n1721_46[1]),.dinb(w_n1290_0[0]),.dout(n3362),.clk(gclk));
	jand g2721(.dina(w_n1562_45[2]),.dinb(w_n877_0[0]),.dout(n3363),.clk(gclk));
	jor g2722(.dina(n3363),.dinb(n3362),.dout(n3364),.clk(gclk));
	jnot g2723(.din(w_n3364_0[1]),.dout(n3365),.clk(gclk));
	jand g2724(.dina(w_n2803_45[2]),.dinb(w_n2378_0[0]),.dout(n3366),.clk(gclk));
	jand g2725(.dina(w_n2808_46[0]),.dinb(w_n1960_0[0]),.dout(n3367),.clk(gclk));
	jor g2726(.dina(n3367),.dinb(n3366),.dout(n3368),.clk(gclk));
	jand g2727(.dina(w_n3368_0[1]),.dinb(w_n3365_0[1]),.dout(n3369),.clk(gclk));
	jnot g2728(.din(w_n3368_0[0]),.dout(n3370),.clk(gclk));
	jand g2729(.dina(w_n3370_0[1]),.dinb(w_n3364_0[0]),.dout(n3371),.clk(gclk));
	jand g2730(.dina(w_n1721_46[0]),.dinb(w_n1288_0[0]),.dout(n3372),.clk(gclk));
	jand g2731(.dina(w_n1562_45[1]),.dinb(w_n1301_0[0]),.dout(n3373),.clk(gclk));
	jor g2732(.dina(n3373),.dinb(n3372),.dout(n3374),.clk(gclk));
	jand g2733(.dina(w_n2803_45[1]),.dinb(w_n2376_0[0]),.dout(n3375),.clk(gclk));
	jand g2734(.dina(w_n2808_45[2]),.dinb(w_n2389_0[0]),.dout(n3376),.clk(gclk));
	jor g2735(.dina(n3376),.dinb(n3375),.dout(n3377),.clk(gclk));
	jnot g2736(.din(w_n3377_0[1]),.dout(n3378),.clk(gclk));
	jand g2737(.dina(w_n3378_0[1]),.dinb(w_n3374_0[1]),.dout(n3379),.clk(gclk));
	jor g2738(.dina(n3379),.dinb(n3371),.dout(n3380),.clk(gclk));
	jnot g2739(.din(w_n3380_0[1]),.dout(n3381),.clk(gclk));
	jnot g2740(.din(w_n3374_0[0]),.dout(n3382),.clk(gclk));
	jand g2741(.dina(w_n3377_0[0]),.dinb(w_n3382_0[1]),.dout(n3383),.clk(gclk));
	jand g2742(.dina(w_n1721_45[2]),.dinb(w_n1285_0[0]),.dout(n3384),.clk(gclk));
	jand g2743(.dina(w_n1562_45[0]),.dinb(w_n1299_0[0]),.dout(n3385),.clk(gclk));
	jor g2744(.dina(n3385),.dinb(n3384),.dout(n3386),.clk(gclk));
	jand g2745(.dina(w_n2803_45[0]),.dinb(w_n2373_0[0]),.dout(n3387),.clk(gclk));
	jand g2746(.dina(w_n2808_45[1]),.dinb(w_n2387_0[0]),.dout(n3388),.clk(gclk));
	jor g2747(.dina(n3388),.dinb(n3387),.dout(n3389),.clk(gclk));
	jnot g2748(.din(w_n3389_0[1]),.dout(n3390),.clk(gclk));
	jand g2749(.dina(w_n3390_0[1]),.dinb(w_n3386_0[1]),.dout(n3391),.clk(gclk));
	jnot g2750(.din(w_n3391_0[1]),.dout(n3392),.clk(gclk));
	jand g2751(.dina(w_n1721_45[1]),.dinb(w_n1282_0[0]),.dout(n3393),.clk(gclk));
	jand g2752(.dina(w_n1562_44[2]),.dinb(w_n1304_0[0]),.dout(n3394),.clk(gclk));
	jor g2753(.dina(n3394),.dinb(n3393),.dout(n3395),.clk(gclk));
	jnot g2754(.din(w_n3395_0[1]),.dout(n3396),.clk(gclk));
	jand g2755(.dina(w_n2803_44[2]),.dinb(w_n2370_0[0]),.dout(n3397),.clk(gclk));
	jand g2756(.dina(w_n2808_45[0]),.dinb(w_n2392_0[0]),.dout(n3398),.clk(gclk));
	jor g2757(.dina(n3398),.dinb(n3397),.dout(n3399),.clk(gclk));
	jand g2758(.dina(w_n3399_0[1]),.dinb(w_n3396_0[1]),.dout(n3400),.clk(gclk));
	jand g2759(.dina(n3400),.dinb(n3392),.dout(n3401),.clk(gclk));
	jnot g2760(.din(w_n3386_0[0]),.dout(n3402),.clk(gclk));
	jand g2761(.dina(w_n3389_0[0]),.dinb(w_n3402_0[1]),.dout(n3403),.clk(gclk));
	jor g2762(.dina(n3403),.dinb(n3401),.dout(n3404),.clk(gclk));
	jor g2763(.dina(n3404),.dinb(n3383),.dout(n3405),.clk(gclk));
	jand g2764(.dina(n3405),.dinb(n3381),.dout(n3406),.clk(gclk));
	jor g2765(.dina(n3406),.dinb(n3369),.dout(n3407),.clk(gclk));
	jand g2766(.dina(n3407),.dinb(n3361),.dout(n3408),.clk(gclk));
	jnot g2767(.din(w_n3408_0[1]),.dout(n3409),.clk(gclk));
	jand g2768(.dina(w_n1721_45[0]),.dinb(w_n896_0[0]),.dout(n3410),.clk(gclk));
	jand g2769(.dina(w_n1562_44[1]),.dinb(w_n1263_0[0]),.dout(n3411),.clk(gclk));
	jor g2770(.dina(n3411),.dinb(n3410),.dout(n3412),.clk(gclk));
	jnot g2771(.din(w_n3412_0[1]),.dout(n3413),.clk(gclk));
	jand g2772(.dina(w_n2803_44[1]),.dinb(w_n1979_0[0]),.dout(n3414),.clk(gclk));
	jand g2773(.dina(w_n2808_44[2]),.dinb(w_n2351_0[0]),.dout(n3415),.clk(gclk));
	jor g2774(.dina(n3415),.dinb(n3414),.dout(n3416),.clk(gclk));
	jand g2775(.dina(w_n3416_0[1]),.dinb(w_n3413_0[1]),.dout(n3417),.clk(gclk));
	jnot g2776(.din(w_n3417_0[1]),.dout(n3418),.clk(gclk));
	jand g2777(.dina(w_n2803_44[0]),.dinb(w_n2286_0[0]),.dout(n3419),.clk(gclk));
	jand g2778(.dina(w_n2808_44[1]),.dinb(w_n1992_0[0]),.dout(n3420),.clk(gclk));
	jor g2779(.dina(n3420),.dinb(n3419),.dout(n3421),.clk(gclk));
	jand g2780(.dina(w_n1721_44[2]),.dinb(w_n909_0[0]),.dout(n3422),.clk(gclk));
	jand g2781(.dina(w_n1562_44[0]),.dinb(w_n1218_0[0]),.dout(n3423),.clk(gclk));
	jor g2782(.dina(n3423),.dinb(n3422),.dout(n3424),.clk(gclk));
	jand g2783(.dina(w_n2803_43[2]),.dinb(w_n1993_0[0]),.dout(n3425),.clk(gclk));
	jand g2784(.dina(w_n2808_44[0]),.dinb(w_n2308_0[0]),.dout(n3426),.clk(gclk));
	jor g2785(.dina(n3426),.dinb(n3425),.dout(n3427),.clk(gclk));
	jnot g2786(.din(w_n3427_0[1]),.dout(n3428),.clk(gclk));
	jand g2787(.dina(w_n3428_0[1]),.dinb(w_n3424_0[1]),.dout(n3429),.clk(gclk));
	jnot g2788(.din(n3429),.dout(n3430),.clk(gclk));
	jand g2789(.dina(w_n1721_44[1]),.dinb(w_n911_0[0]),.dout(n3431),.clk(gclk));
	jand g2790(.dina(w_n1562_43[2]),.dinb(w_n1223_0[0]),.dout(n3432),.clk(gclk));
	jor g2791(.dina(n3432),.dinb(n3431),.dout(n3433),.clk(gclk));
	jand g2792(.dina(w_n2803_43[1]),.dinb(w_n1995_0[0]),.dout(n3434),.clk(gclk));
	jand g2793(.dina(w_n2808_43[2]),.dinb(w_n2313_0[0]),.dout(n3435),.clk(gclk));
	jor g2794(.dina(n3435),.dinb(n3434),.dout(n3436),.clk(gclk));
	jnot g2795(.din(w_n3436_0[1]),.dout(n3437),.clk(gclk));
	jand g2796(.dina(w_n3437_0[1]),.dinb(w_n3433_0[1]),.dout(n3438),.clk(gclk));
	jand g2797(.dina(w_n2803_43[0]),.dinb(w_n1999_0[0]),.dout(n3439),.clk(gclk));
	jand g2798(.dina(w_n2808_43[1]),.dinb(w_n2315_0[0]),.dout(n3440),.clk(gclk));
	jor g2799(.dina(n3440),.dinb(n3439),.dout(n3441),.clk(gclk));
	jnot g2800(.din(w_n3441_0[1]),.dout(n3442),.clk(gclk));
	jand g2801(.dina(w_n1721_44[0]),.dinb(w_n915_0[0]),.dout(n3443),.clk(gclk));
	jand g2802(.dina(w_n1562_43[1]),.dinb(w_n1225_0[0]),.dout(n3444),.clk(gclk));
	jor g2803(.dina(n3444),.dinb(n3443),.dout(n3445),.clk(gclk));
	jand g2804(.dina(w_n3445_0[1]),.dinb(w_n3442_0[1]),.dout(n3446),.clk(gclk));
	jor g2805(.dina(n3446),.dinb(w_n3438_0[1]),.dout(n3447),.clk(gclk));
	jnot g2806(.din(n3447),.dout(n3448),.clk(gclk));
	jand g2807(.dina(w_n1721_43[2]),.dinb(w_n913_0[0]),.dout(n3449),.clk(gclk));
	jand g2808(.dina(w_n1562_43[0]),.dinb(w_n1216_0[0]),.dout(n3450),.clk(gclk));
	jor g2809(.dina(n3450),.dinb(n3449),.dout(n3451),.clk(gclk));
	jand g2810(.dina(w_n2803_42[2]),.dinb(w_n1997_0[0]),.dout(n3452),.clk(gclk));
	jand g2811(.dina(w_n2808_43[0]),.dinb(w_n2306_0[0]),.dout(n3453),.clk(gclk));
	jor g2812(.dina(n3453),.dinb(n3452),.dout(n3454),.clk(gclk));
	jnot g2813(.din(w_n3454_0[1]),.dout(n3455),.clk(gclk));
	jand g2814(.dina(w_n3455_0[1]),.dinb(w_n3451_0[1]),.dout(n3456),.clk(gclk));
	jnot g2815(.din(n3456),.dout(n3457),.clk(gclk));
	jand g2816(.dina(w_n3457_0[1]),.dinb(w_n3448_0[1]),.dout(n3458),.clk(gclk));
	jand g2817(.dina(n3458),.dinb(n3430),.dout(n3459),.clk(gclk));
	jand g2818(.dina(w_n1721_43[1]),.dinb(w_n922_0[0]),.dout(n3460),.clk(gclk));
	jnot g2819(.din(n3460),.dout(n3461),.clk(gclk));
	jor g2820(.dina(w_n1721_43[0]),.dinb(w_in143_0[0]),.dout(n3462),.clk(gclk));
	jand g2821(.dina(n3462),.dinb(n3461),.dout(n3463),.clk(gclk));
	jand g2822(.dina(w_n3463_0[2]),.dinb(w_n3459_0[1]),.dout(n3464),.clk(gclk));
	jand g2823(.dina(n3464),.dinb(w_n3421_0[2]),.dout(n3465),.clk(gclk));
	jnot g2824(.din(w_n3465_0[1]),.dout(n3466),.clk(gclk));
	jand g2825(.dina(w_n1721_42[2]),.dinb(w_n962_0[0]),.dout(n3467),.clk(gclk));
	jand g2826(.dina(w_n1562_42[2]),.dinb(w_n1198_0[0]),.dout(n3468),.clk(gclk));
	jor g2827(.dina(n3468),.dinb(n3467),.dout(n3469),.clk(gclk));
	jand g2828(.dina(w_n2803_42[1]),.dinb(w_n2029_0[0]),.dout(n3470),.clk(gclk));
	jand g2829(.dina(w_n2808_42[2]),.dinb(w_n2266_0[0]),.dout(n3471),.clk(gclk));
	jor g2830(.dina(n3471),.dinb(n3470),.dout(n3472),.clk(gclk));
	jnot g2831(.din(w_n3472_0[1]),.dout(n3473),.clk(gclk));
	jand g2832(.dina(w_n3473_0[1]),.dinb(w_n3469_0[1]),.dout(n3474),.clk(gclk));
	jnot g2833(.din(n3474),.dout(n3475),.clk(gclk));
	jand g2834(.dina(w_n2803_42[0]),.dinb(w_n2027_0[0]),.dout(n3476),.clk(gclk));
	jand g2835(.dina(w_n2808_42[1]),.dinb(w_n2269_0[0]),.dout(n3477),.clk(gclk));
	jor g2836(.dina(n3477),.dinb(n3476),.dout(n3478),.clk(gclk));
	jnot g2837(.din(w_n3478_0[1]),.dout(n3479),.clk(gclk));
	jand g2838(.dina(w_n1721_42[1]),.dinb(w_n960_0[0]),.dout(n3480),.clk(gclk));
	jand g2839(.dina(w_n1562_42[1]),.dinb(w_n1201_0[0]),.dout(n3481),.clk(gclk));
	jor g2840(.dina(n3481),.dinb(n3480),.dout(n3482),.clk(gclk));
	jand g2841(.dina(w_n3482_0[1]),.dinb(w_n3479_0[1]),.dout(n3483),.clk(gclk));
	jand g2842(.dina(w_n1721_42[0]),.dinb(w_n964_0[0]),.dout(n3484),.clk(gclk));
	jand g2843(.dina(w_n1562_42[0]),.dinb(w_n1188_0[0]),.dout(n3485),.clk(gclk));
	jor g2844(.dina(n3485),.dinb(n3484),.dout(n3486),.clk(gclk));
	jand g2845(.dina(w_n2803_41[2]),.dinb(w_n2031_0[0]),.dout(n3487),.clk(gclk));
	jand g2846(.dina(w_n2808_42[0]),.dinb(w_n2256_0[0]),.dout(n3488),.clk(gclk));
	jor g2847(.dina(n3488),.dinb(n3487),.dout(n3489),.clk(gclk));
	jnot g2848(.din(w_n3489_0[1]),.dout(n3490),.clk(gclk));
	jand g2849(.dina(w_n3490_0[1]),.dinb(w_n3486_0[1]),.dout(n3491),.clk(gclk));
	jor g2850(.dina(n3491),.dinb(n3483),.dout(n3492),.clk(gclk));
	jnot g2851(.din(n3492),.dout(n3493),.clk(gclk));
	jnot g2852(.din(w_n3486_0[0]),.dout(n3494),.clk(gclk));
	jand g2853(.dina(w_n3489_0[0]),.dinb(w_n3494_0[1]),.dout(n3495),.clk(gclk));
	jand g2854(.dina(w_n1721_41[2]),.dinb(w_n958_0[0]),.dout(n3496),.clk(gclk));
	jand g2855(.dina(w_n1562_41[2]),.dinb(w_n1190_0[0]),.dout(n3497),.clk(gclk));
	jor g2856(.dina(n3497),.dinb(n3496),.dout(n3498),.clk(gclk));
	jnot g2857(.din(w_n3498_0[1]),.dout(n3499),.clk(gclk));
	jand g2858(.dina(w_n2803_41[1]),.dinb(w_n2025_0[0]),.dout(n3500),.clk(gclk));
	jand g2859(.dina(w_n2808_41[2]),.dinb(w_n2258_0[0]),.dout(n3501),.clk(gclk));
	jor g2860(.dina(n3501),.dinb(n3500),.dout(n3502),.clk(gclk));
	jand g2861(.dina(w_n3502_0[1]),.dinb(w_n3499_0[1]),.dout(n3503),.clk(gclk));
	jor g2862(.dina(n3503),.dinb(n3495),.dout(n3504),.clk(gclk));
	jnot g2863(.din(w_n3502_0[0]),.dout(n3505),.clk(gclk));
	jand g2864(.dina(w_n3505_0[1]),.dinb(w_n3498_0[0]),.dout(n3506),.clk(gclk));
	jnot g2865(.din(n3506),.dout(n3507),.clk(gclk));
	jand g2866(.dina(w_n1721_41[1]),.dinb(w_n953_0[0]),.dout(n3508),.clk(gclk));
	jand g2867(.dina(w_n1562_41[1]),.dinb(w_n1195_0[0]),.dout(n3509),.clk(gclk));
	jor g2868(.dina(n3509),.dinb(n3508),.dout(n3510),.clk(gclk));
	jand g2869(.dina(w_n2803_41[0]),.dinb(w_n2020_0[0]),.dout(n3511),.clk(gclk));
	jand g2870(.dina(w_n2808_41[1]),.dinb(w_n2263_0[0]),.dout(n3512),.clk(gclk));
	jor g2871(.dina(n3512),.dinb(n3511),.dout(n3513),.clk(gclk));
	jnot g2872(.din(w_n3513_0[1]),.dout(n3514),.clk(gclk));
	jand g2873(.dina(w_n3514_0[1]),.dinb(w_n3510_0[1]),.dout(n3515),.clk(gclk));
	jnot g2874(.din(w_n3515_0[1]),.dout(n3516),.clk(gclk));
	jand g2875(.dina(w_n1721_41[0]),.dinb(w_n946_0[0]),.dout(n3517),.clk(gclk));
	jand g2876(.dina(w_n1562_41[0]),.dinb(w_n941_0[0]),.dout(n3518),.clk(gclk));
	jor g2877(.dina(n3518),.dinb(n3517),.dout(n3519),.clk(gclk));
	jand g2878(.dina(w_n2803_40[2]),.dinb(w_n2013_0[0]),.dout(n3520),.clk(gclk));
	jand g2879(.dina(w_n2808_41[0]),.dinb(w_n2008_0[0]),.dout(n3521),.clk(gclk));
	jor g2880(.dina(n3521),.dinb(n3520),.dout(n3522),.clk(gclk));
	jnot g2881(.din(w_n3522_0[1]),.dout(n3523),.clk(gclk));
	jand g2882(.dina(w_n3523_0[1]),.dinb(w_n3519_0[1]),.dout(n3524),.clk(gclk));
	jand g2883(.dina(w_n2803_40[1]),.dinb(w_n2022_0[0]),.dout(n3525),.clk(gclk));
	jand g2884(.dina(w_n2808_40[2]),.dinb(w_n2010_0[0]),.dout(n3526),.clk(gclk));
	jor g2885(.dina(n3526),.dinb(n3525),.dout(n3527),.clk(gclk));
	jnot g2886(.din(w_n3527_0[1]),.dout(n3528),.clk(gclk));
	jand g2887(.dina(w_n1721_40[2]),.dinb(w_n955_0[0]),.dout(n3529),.clk(gclk));
	jand g2888(.dina(w_n1562_40[2]),.dinb(w_n943_0[0]),.dout(n3530),.clk(gclk));
	jor g2889(.dina(n3530),.dinb(n3529),.dout(n3531),.clk(gclk));
	jand g2890(.dina(w_n3531_0[1]),.dinb(w_n3528_0[1]),.dout(n3532),.clk(gclk));
	jor g2891(.dina(n3532),.dinb(n3524),.dout(n3533),.clk(gclk));
	jnot g2892(.din(w_n3533_0[1]),.dout(n3534),.clk(gclk));
	jand g2893(.dina(w_n2803_40[0]),.dinb(w_n2249_0[0]),.dout(n3535),.clk(gclk));
	jand g2894(.dina(w_n2808_40[1]),.dinb(w_n2016_0[0]),.dout(n3536),.clk(gclk));
	jor g2895(.dina(n3536),.dinb(n3535),.dout(n3537),.clk(gclk));
	jand g2896(.dina(w_n1721_40[1]),.dinb(w_n1181_0[0]),.dout(n3538),.clk(gclk));
	jand g2897(.dina(w_n1562_40[1]),.dinb(w_n949_0[0]),.dout(n3539),.clk(gclk));
	jor g2898(.dina(n3539),.dinb(n3538),.dout(n3540),.clk(gclk));
	jnot g2899(.din(w_n3540_0[1]),.dout(n3541),.clk(gclk));
	jand g2900(.dina(w_n3541_0[1]),.dinb(w_n3537_0[1]),.dout(n3542),.clk(gclk));
	jnot g2901(.din(w_n3519_0[0]),.dout(n3543),.clk(gclk));
	jand g2902(.dina(w_n3522_0[0]),.dinb(w_n3543_0[1]),.dout(n3544),.clk(gclk));
	jor g2903(.dina(n3544),.dinb(n3542),.dout(n3545),.clk(gclk));
	jand g2904(.dina(n3545),.dinb(w_n3534_0[1]),.dout(n3546),.clk(gclk));
	jnot g2905(.din(w_n3510_0[0]),.dout(n3547),.clk(gclk));
	jand g2906(.dina(w_n3513_0[0]),.dinb(w_n3547_0[1]),.dout(n3548),.clk(gclk));
	jnot g2907(.din(w_n3531_0[0]),.dout(n3549),.clk(gclk));
	jand g2908(.dina(w_n3549_0[1]),.dinb(w_n3527_0[0]),.dout(n3550),.clk(gclk));
	jor g2909(.dina(n3550),.dinb(n3548),.dout(n3551),.clk(gclk));
	jor g2910(.dina(n3551),.dinb(n3546),.dout(n3552),.clk(gclk));
	jand g2911(.dina(n3552),.dinb(n3516),.dout(n3553),.clk(gclk));
	jand g2912(.dina(n3553),.dinb(w_n3507_0[1]),.dout(n3554),.clk(gclk));
	jor g2913(.dina(n3554),.dinb(n3504),.dout(n3555),.clk(gclk));
	jand g2914(.dina(n3555),.dinb(w_n3493_0[1]),.dout(n3556),.clk(gclk));
	jnot g2915(.din(w_n3469_0[0]),.dout(n3557),.clk(gclk));
	jand g2916(.dina(w_n3472_0[0]),.dinb(w_n3557_0[1]),.dout(n3558),.clk(gclk));
	jnot g2917(.din(w_n3482_0[0]),.dout(n3559),.clk(gclk));
	jand g2918(.dina(w_n3559_0[1]),.dinb(w_n3478_0[0]),.dout(n3560),.clk(gclk));
	jor g2919(.dina(n3560),.dinb(n3558),.dout(n3561),.clk(gclk));
	jor g2920(.dina(n3561),.dinb(n3556),.dout(n3562),.clk(gclk));
	jand g2921(.dina(n3562),.dinb(w_n3475_0[1]),.dout(n3563),.clk(gclk));
	jnot g2922(.din(w_n3563_0[1]),.dout(n3564),.clk(gclk));
	jand g2923(.dina(w_n1721_40[0]),.dinb(w_n1179_0[0]),.dout(n3565),.clk(gclk));
	jand g2924(.dina(w_n1562_40[0]),.dinb(w_n1172_0[0]),.dout(n3566),.clk(gclk));
	jor g2925(.dina(n3566),.dinb(n3565),.dout(n3567),.clk(gclk));
	jnot g2926(.din(w_n3567_0[1]),.dout(n3568),.clk(gclk));
	jand g2927(.dina(w_n2803_39[2]),.dinb(w_n2247_0[0]),.dout(n3569),.clk(gclk));
	jand g2928(.dina(w_n2808_40[0]),.dinb(w_n2240_0[0]),.dout(n3570),.clk(gclk));
	jor g2929(.dina(n3570),.dinb(n3569),.dout(n3571),.clk(gclk));
	jand g2930(.dina(w_n3571_0[1]),.dinb(w_n3568_0[1]),.dout(n3572),.clk(gclk));
	jnot g2931(.din(w_n3572_0[1]),.dout(n3573),.clk(gclk));
	jand g2932(.dina(w_n1721_39[2]),.dinb(w_n978_0[0]),.dout(n3574),.clk(gclk));
	jand g2933(.dina(w_n1562_39[2]),.dinb(w_n975_0[0]),.dout(n3575),.clk(gclk));
	jor g2934(.dina(n3575),.dinb(n3574),.dout(n3576),.clk(gclk));
	jand g2935(.dina(w_n2803_39[1]),.dinb(w_n2045_0[0]),.dout(n3577),.clk(gclk));
	jand g2936(.dina(w_n2808_39[2]),.dinb(w_n2042_0[0]),.dout(n3578),.clk(gclk));
	jor g2937(.dina(n3578),.dinb(n3577),.dout(n3579),.clk(gclk));
	jnot g2938(.din(w_n3579_0[1]),.dout(n3580),.clk(gclk));
	jand g2939(.dina(w_n3580_0[1]),.dinb(w_n3576_0[1]),.dout(n3581),.clk(gclk));
	jand g2940(.dina(w_n1721_39[1]),.dinb(w_n983_0[0]),.dout(n3582),.clk(gclk));
	jand g2941(.dina(w_n1562_39[1]),.dinb(w_n980_0[0]),.dout(n3583),.clk(gclk));
	jor g2942(.dina(n3583),.dinb(n3582),.dout(n3584),.clk(gclk));
	jnot g2943(.din(w_n3584_0[1]),.dout(n3585),.clk(gclk));
	jand g2944(.dina(w_n2803_39[0]),.dinb(w_n2050_0[0]),.dout(n3586),.clk(gclk));
	jand g2945(.dina(w_n2808_39[1]),.dinb(w_n2047_0[0]),.dout(n3587),.clk(gclk));
	jor g2946(.dina(n3587),.dinb(n3586),.dout(n3588),.clk(gclk));
	jand g2947(.dina(w_n3588_0[1]),.dinb(w_n3585_0[1]),.dout(n3589),.clk(gclk));
	jnot g2948(.din(w_n3589_0[1]),.dout(n3590),.clk(gclk));
	jand g2949(.dina(w_n1721_39[0]),.dinb(w_n1158_0[0]),.dout(n3591),.clk(gclk));
	jand g2950(.dina(w_n1562_39[0]),.dinb(w_n990_0[0]),.dout(n3592),.clk(gclk));
	jor g2951(.dina(n3592),.dinb(n3591),.dout(n3593),.clk(gclk));
	jand g2952(.dina(w_n2803_38[2]),.dinb(w_n2226_0[0]),.dout(n3594),.clk(gclk));
	jand g2953(.dina(w_n2808_39[0]),.dinb(w_n2057_0[0]),.dout(n3595),.clk(gclk));
	jor g2954(.dina(n3595),.dinb(n3594),.dout(n3596),.clk(gclk));
	jnot g2955(.din(w_n3596_0[1]),.dout(n3597),.clk(gclk));
	jand g2956(.dina(w_n3597_0[1]),.dinb(w_n3593_0[1]),.dout(n3598),.clk(gclk));
	jand g2957(.dina(w_n2803_38[1]),.dinb(w_n2215_0[0]),.dout(n3599),.clk(gclk));
	jand g2958(.dina(w_n2808_38[2]),.dinb(w_n2219_0[0]),.dout(n3600),.clk(gclk));
	jor g2959(.dina(n3600),.dinb(n3599),.dout(n3601),.clk(gclk));
	jand g2960(.dina(w_n1721_38[2]),.dinb(w_n1147_0[0]),.dout(n3602),.clk(gclk));
	jand g2961(.dina(w_n1562_38[2]),.dinb(w_n1151_0[0]),.dout(n3603),.clk(gclk));
	jor g2962(.dina(n3603),.dinb(n3602),.dout(n3604),.clk(gclk));
	jnot g2963(.din(w_n3604_0[1]),.dout(n3605),.clk(gclk));
	jand g2964(.dina(w_n3605_0[1]),.dinb(w_n3601_0[1]),.dout(n3606),.clk(gclk));
	jand g2965(.dina(w_n2803_38[0]),.dinb(w_n2228_0[0]),.dout(n3607),.clk(gclk));
	jand g2966(.dina(w_n2808_38[1]),.dinb(w_n2221_0[0]),.dout(n3608),.clk(gclk));
	jor g2967(.dina(n3608),.dinb(n3607),.dout(n3609),.clk(gclk));
	jand g2968(.dina(w_n1721_38[1]),.dinb(w_n1160_0[0]),.dout(n3610),.clk(gclk));
	jand g2969(.dina(w_n1562_38[1]),.dinb(w_n1153_0[0]),.dout(n3611),.clk(gclk));
	jor g2970(.dina(n3611),.dinb(n3610),.dout(n3612),.clk(gclk));
	jnot g2971(.din(w_n3612_0[1]),.dout(n3613),.clk(gclk));
	jand g2972(.dina(w_n3613_0[1]),.dinb(w_n3609_0[1]),.dout(n3614),.clk(gclk));
	jor g2973(.dina(n3614),.dinb(n3606),.dout(n3615),.clk(gclk));
	jnot g2974(.din(w_n3615_0[1]),.dout(n3616),.clk(gclk));
	jand g2975(.dina(w_n1721_38[0]),.dinb(w_n993_0[0]),.dout(n3617),.clk(gclk));
	jand g2976(.dina(w_n1562_38[0]),.dinb(w_n1140_0[0]),.dout(n3618),.clk(gclk));
	jor g2977(.dina(n3618),.dinb(n3617),.dout(n3619),.clk(gclk));
	jnot g2978(.din(w_n3619_0[1]),.dout(n3620),.clk(gclk));
	jand g2979(.dina(w_n2803_37[2]),.dinb(w_n2060_0[0]),.dout(n3621),.clk(gclk));
	jand g2980(.dina(w_n2808_38[0]),.dinb(w_n2208_0[0]),.dout(n3622),.clk(gclk));
	jor g2981(.dina(n3622),.dinb(n3621),.dout(n3623),.clk(gclk));
	jand g2982(.dina(w_n3623_0[1]),.dinb(w_n3620_0[1]),.dout(n3624),.clk(gclk));
	jnot g2983(.din(w_n3624_0[1]),.dout(n3625),.clk(gclk));
	jand g2984(.dina(w_n1721_37[2]),.dinb(w_n995_0[0]),.dout(n3626),.clk(gclk));
	jand g2985(.dina(w_n1562_37[2]),.dinb(w_n1142_0[0]),.dout(n3627),.clk(gclk));
	jor g2986(.dina(n3627),.dinb(n3626),.dout(n3628),.clk(gclk));
	jand g2987(.dina(w_n2803_37[1]),.dinb(w_n2062_0[0]),.dout(n3629),.clk(gclk));
	jand g2988(.dina(w_n2808_37[2]),.dinb(w_n2210_0[0]),.dout(n3630),.clk(gclk));
	jor g2989(.dina(n3630),.dinb(n3629),.dout(n3631),.clk(gclk));
	jnot g2990(.din(w_n3631_0[1]),.dout(n3632),.clk(gclk));
	jand g2991(.dina(w_n3632_0[1]),.dinb(w_n3628_0[1]),.dout(n3633),.clk(gclk));
	jand g2992(.dina(w_n1721_37[1]),.dinb(w_n1005_0[0]),.dout(n3634),.clk(gclk));
	jand g2993(.dina(w_n1562_37[1]),.dinb(w_n1002_0[0]),.dout(n3635),.clk(gclk));
	jor g2994(.dina(n3635),.dinb(n3634),.dout(n3636),.clk(gclk));
	jand g2995(.dina(w_n2803_37[0]),.dinb(w_n2072_0[0]),.dout(n3637),.clk(gclk));
	jand g2996(.dina(w_n2808_37[1]),.dinb(w_n2069_0[0]),.dout(n3638),.clk(gclk));
	jor g2997(.dina(n3638),.dinb(n3637),.dout(n3639),.clk(gclk));
	jnot g2998(.din(w_n3639_0[1]),.dout(n3640),.clk(gclk));
	jand g2999(.dina(w_n3640_0[1]),.dinb(w_n3636_0[1]),.dout(n3641),.clk(gclk));
	jnot g3000(.din(w_n3636_0[0]),.dout(n3642),.clk(gclk));
	jand g3001(.dina(w_n3639_0[0]),.dinb(w_n3642_0[1]),.dout(n3643),.clk(gclk));
	jnot g3002(.din(w_n3643_0[1]),.dout(n3644),.clk(gclk));
	jand g3003(.dina(w_n1721_37[0]),.dinb(w_n1010_0[0]),.dout(n3645),.clk(gclk));
	jand g3004(.dina(w_n1562_37[0]),.dinb(w_n1007_0[0]),.dout(n3646),.clk(gclk));
	jor g3005(.dina(n3646),.dinb(n3645),.dout(n3647),.clk(gclk));
	jand g3006(.dina(w_n2803_36[2]),.dinb(w_n2077_0[0]),.dout(n3648),.clk(gclk));
	jand g3007(.dina(w_n2808_37[0]),.dinb(w_n2074_0[0]),.dout(n3649),.clk(gclk));
	jor g3008(.dina(n3649),.dinb(n3648),.dout(n3650),.clk(gclk));
	jnot g3009(.din(w_n3650_0[1]),.dout(n3651),.clk(gclk));
	jand g3010(.dina(w_n3651_0[1]),.dinb(w_n3647_0[1]),.dout(n3652),.clk(gclk));
	jand g3011(.dina(w_n1721_36[2]),.dinb(w_n1126_0[0]),.dout(n3653),.clk(gclk));
	jand g3012(.dina(w_n1562_36[2]),.dinb(w_n1012_0[0]),.dout(n3654),.clk(gclk));
	jor g3013(.dina(n3654),.dinb(n3653),.dout(n3655),.clk(gclk));
	jand g3014(.dina(w_n2803_36[1]),.dinb(w_n2194_0[0]),.dout(n3656),.clk(gclk));
	jand g3015(.dina(w_n2808_36[2]),.dinb(w_n2079_0[0]),.dout(n3657),.clk(gclk));
	jor g3016(.dina(n3657),.dinb(n3656),.dout(n3658),.clk(gclk));
	jnot g3017(.din(w_n3658_0[1]),.dout(n3659),.clk(gclk));
	jand g3018(.dina(w_n3659_0[1]),.dinb(w_n3655_0[1]),.dout(n3660),.clk(gclk));
	jand g3019(.dina(w_n2803_36[0]),.dinb(w_n2183_0[0]),.dout(n3661),.clk(gclk));
	jand g3020(.dina(w_n2808_36[1]),.dinb(w_n2187_0[0]),.dout(n3662),.clk(gclk));
	jor g3021(.dina(n3662),.dinb(n3661),.dout(n3663),.clk(gclk));
	jand g3022(.dina(w_n1721_36[1]),.dinb(w_n1115_0[0]),.dout(n3664),.clk(gclk));
	jand g3023(.dina(w_n1562_36[1]),.dinb(w_n1119_0[0]),.dout(n3665),.clk(gclk));
	jor g3024(.dina(n3665),.dinb(n3664),.dout(n3666),.clk(gclk));
	jnot g3025(.din(w_n3666_0[1]),.dout(n3667),.clk(gclk));
	jand g3026(.dina(w_n3667_0[1]),.dinb(w_n3663_0[1]),.dout(n3668),.clk(gclk));
	jnot g3027(.din(w_n3668_0[1]),.dout(n3669),.clk(gclk));
	jand g3028(.dina(w_n1721_36[0]),.dinb(w_n1015_0[0]),.dout(n3670),.clk(gclk));
	jand g3029(.dina(w_n1562_36[0]),.dinb(w_n1108_0[0]),.dout(n3671),.clk(gclk));
	jor g3030(.dina(n3671),.dinb(n3670),.dout(n3672),.clk(gclk));
	jand g3031(.dina(w_n2803_35[2]),.dinb(w_n2082_0[0]),.dout(n3673),.clk(gclk));
	jand g3032(.dina(w_n2808_36[0]),.dinb(w_n2176_0[0]),.dout(n3674),.clk(gclk));
	jor g3033(.dina(n3674),.dinb(n3673),.dout(n3675),.clk(gclk));
	jnot g3034(.din(w_n3675_0[1]),.dout(n3676),.clk(gclk));
	jand g3035(.dina(w_n3676_0[1]),.dinb(w_n3672_0[1]),.dout(n3677),.clk(gclk));
	jand g3036(.dina(w_n1721_35[2]),.dinb(w_n1017_0[0]),.dout(n3678),.clk(gclk));
	jand g3037(.dina(w_n1562_35[2]),.dinb(w_n1110_0[0]),.dout(n3679),.clk(gclk));
	jor g3038(.dina(n3679),.dinb(n3678),.dout(n3680),.clk(gclk));
	jand g3039(.dina(w_n2803_35[1]),.dinb(w_n2084_0[0]),.dout(n3681),.clk(gclk));
	jand g3040(.dina(w_n2808_35[2]),.dinb(w_n2178_0[0]),.dout(n3682),.clk(gclk));
	jor g3041(.dina(n3682),.dinb(n3681),.dout(n3683),.clk(gclk));
	jnot g3042(.din(w_n3683_0[1]),.dout(n3684),.clk(gclk));
	jand g3043(.dina(w_n3684_0[1]),.dinb(w_n3680_0[1]),.dout(n3685),.clk(gclk));
	jand g3044(.dina(w_n1721_35[1]),.dinb(w_n1022_0[0]),.dout(n3686),.clk(gclk));
	jand g3045(.dina(w_n1562_35[1]),.dinb(w_n1019_0[0]),.dout(n3687),.clk(gclk));
	jor g3046(.dina(n3687),.dinb(n3686),.dout(n3688),.clk(gclk));
	jnot g3047(.din(w_n3688_0[1]),.dout(n3689),.clk(gclk));
	jand g3048(.dina(w_n2803_35[0]),.dinb(w_n2089_0[0]),.dout(n3690),.clk(gclk));
	jand g3049(.dina(w_n2808_35[1]),.dinb(w_n2086_0[0]),.dout(n3691),.clk(gclk));
	jor g3050(.dina(n3691),.dinb(n3690),.dout(n3692),.clk(gclk));
	jand g3051(.dina(w_n3692_0[1]),.dinb(w_n3689_0[1]),.dout(n3693),.clk(gclk));
	jnot g3052(.din(w_n3693_0[1]),.dout(n3694),.clk(gclk));
	jnot g3053(.din(w_n3692_0[0]),.dout(n3695),.clk(gclk));
	jand g3054(.dina(w_n3695_0[1]),.dinb(w_n3688_0[0]),.dout(n3696),.clk(gclk));
	jand g3055(.dina(w_n1721_35[0]),.dinb(w_n1027_0[0]),.dout(n3697),.clk(gclk));
	jand g3056(.dina(w_n1562_35[0]),.dinb(w_n1024_0[0]),.dout(n3698),.clk(gclk));
	jor g3057(.dina(n3698),.dinb(n3697),.dout(n3699),.clk(gclk));
	jnot g3058(.din(w_n3699_0[1]),.dout(n3700),.clk(gclk));
	jand g3059(.dina(w_n2803_34[2]),.dinb(w_n2094_0[0]),.dout(n3701),.clk(gclk));
	jand g3060(.dina(w_n2808_35[0]),.dinb(w_n2091_0[0]),.dout(n3702),.clk(gclk));
	jor g3061(.dina(n3702),.dinb(n3701),.dout(n3703),.clk(gclk));
	jand g3062(.dina(w_n3703_0[1]),.dinb(w_n3700_0[1]),.dout(n3704),.clk(gclk));
	jnot g3063(.din(w_n3704_0[1]),.dout(n3705),.clk(gclk));
	jand g3064(.dina(w_n1721_34[2]),.dinb(w_n1094_0[0]),.dout(n3706),.clk(gclk));
	jand g3065(.dina(w_n1562_34[2]),.dinb(w_n1034_0[0]),.dout(n3707),.clk(gclk));
	jor g3066(.dina(n3707),.dinb(n3706),.dout(n3708),.clk(gclk));
	jand g3067(.dina(w_n2803_34[1]),.dinb(w_n2162_0[0]),.dout(n3709),.clk(gclk));
	jand g3068(.dina(w_n2808_34[2]),.dinb(w_n2101_0[0]),.dout(n3710),.clk(gclk));
	jor g3069(.dina(n3710),.dinb(n3709),.dout(n3711),.clk(gclk));
	jnot g3070(.din(w_n3711_0[1]),.dout(n3712),.clk(gclk));
	jand g3071(.dina(w_n3712_0[1]),.dinb(w_n3708_0[1]),.dout(n3713),.clk(gclk));
	jand g3072(.dina(w_n2803_34[0]),.dinb(w_n2151_0[0]),.dout(n3714),.clk(gclk));
	jand g3073(.dina(w_n2808_34[1]),.dinb(w_n2155_0[0]),.dout(n3715),.clk(gclk));
	jor g3074(.dina(n3715),.dinb(n3714),.dout(n3716),.clk(gclk));
	jand g3075(.dina(w_n1721_34[1]),.dinb(w_n1083_0[0]),.dout(n3717),.clk(gclk));
	jand g3076(.dina(w_n1562_34[1]),.dinb(w_n1087_0[0]),.dout(n3718),.clk(gclk));
	jor g3077(.dina(n3718),.dinb(n3717),.dout(n3719),.clk(gclk));
	jnot g3078(.din(w_n3719_0[1]),.dout(n3720),.clk(gclk));
	jand g3079(.dina(w_n3720_0[1]),.dinb(w_n3716_0[1]),.dout(n3721),.clk(gclk));
	jnot g3080(.din(w_n3721_0[1]),.dout(n3722),.clk(gclk));
	jand g3081(.dina(w_n1721_34[0]),.dinb(w_n1037_0[0]),.dout(n3723),.clk(gclk));
	jand g3082(.dina(w_n1562_34[0]),.dinb(w_n1076_0[0]),.dout(n3724),.clk(gclk));
	jor g3083(.dina(n3724),.dinb(n3723),.dout(n3725),.clk(gclk));
	jand g3084(.dina(w_n2803_33[2]),.dinb(w_n2104_0[0]),.dout(n3726),.clk(gclk));
	jand g3085(.dina(w_n2808_34[0]),.dinb(w_n2144_0[0]),.dout(n3727),.clk(gclk));
	jor g3086(.dina(n3727),.dinb(n3726),.dout(n3728),.clk(gclk));
	jnot g3087(.din(w_n3728_0[1]),.dout(n3729),.clk(gclk));
	jand g3088(.dina(w_n3729_0[1]),.dinb(w_n3725_0[1]),.dout(n3730),.clk(gclk));
	jand g3089(.dina(w_n2803_33[1]),.dinb(w_n2138_0[0]),.dout(n3731),.clk(gclk));
	jand g3090(.dina(w_n2808_33[2]),.dinb(w_n2146_0[0]),.dout(n3732),.clk(gclk));
	jor g3091(.dina(n3732),.dinb(n3731),.dout(n3733),.clk(gclk));
	jnot g3092(.din(w_n3733_0[1]),.dout(n3734),.clk(gclk));
	jand g3093(.dina(w_n1721_33[2]),.dinb(w_n1070_0[0]),.dout(n3735),.clk(gclk));
	jand g3094(.dina(w_n1562_33[2]),.dinb(w_n1078_0[0]),.dout(n3736),.clk(gclk));
	jor g3095(.dina(n3736),.dinb(n3735),.dout(n3737),.clk(gclk));
	jand g3096(.dina(w_n3737_0[1]),.dinb(w_n3734_0[1]),.dout(n3738),.clk(gclk));
	jand g3097(.dina(w_n2803_33[0]),.dinb(w_n2140_0[0]),.dout(n3739),.clk(gclk));
	jand g3098(.dina(w_n2808_33[1]),.dinb(w_n2133_0[0]),.dout(n3740),.clk(gclk));
	jor g3099(.dina(n3740),.dinb(n3739),.dout(n3741),.clk(gclk));
	jand g3100(.dina(w_n1721_33[1]),.dinb(w_n1072_0[0]),.dout(n3742),.clk(gclk));
	jand g3101(.dina(w_n1562_33[1]),.dinb(w_n1065_0[0]),.dout(n3743),.clk(gclk));
	jor g3102(.dina(n3743),.dinb(n3742),.dout(n3744),.clk(gclk));
	jnot g3103(.din(w_n3744_0[1]),.dout(n3745),.clk(gclk));
	jand g3104(.dina(w_n3745_0[1]),.dinb(w_n3741_0[1]),.dout(n3746),.clk(gclk));
	jnot g3105(.din(w_n3746_0[1]),.dout(n3747),.clk(gclk));
	jnot g3106(.din(w_n3741_0[0]),.dout(n3748),.clk(gclk));
	jand g3107(.dina(w_n3744_0[0]),.dinb(w_n3748_0[1]),.dout(n3749),.clk(gclk));
	jand g3108(.dina(w_n2803_32[2]),.dinb(w_n2127_0[0]),.dout(n3750),.clk(gclk));
	jand g3109(.dina(w_n2808_33[0]),.dinb(w_n2131_0[0]),.dout(n3751),.clk(gclk));
	jor g3110(.dina(n3751),.dinb(n3750),.dout(n3752),.clk(gclk));
	jand g3111(.dina(w_n1721_33[0]),.dinb(w_n1059_0[0]),.dout(n3753),.clk(gclk));
	jand g3112(.dina(w_n1562_33[0]),.dinb(w_n1063_0[0]),.dout(n3754),.clk(gclk));
	jor g3113(.dina(n3754),.dinb(n3753),.dout(n3755),.clk(gclk));
	jnot g3114(.din(w_n3755_0[1]),.dout(n3756),.clk(gclk));
	jand g3115(.dina(w_n3756_0[1]),.dinb(w_n3752_0[1]),.dout(n3757),.clk(gclk));
	jnot g3116(.din(w_n3757_0[1]),.dout(n3758),.clk(gclk));
	jor g3117(.dina(w_n2808_32[2]),.dinb(w_in21_0[1]),.dout(n3759),.clk(gclk));
	jor g3118(.dina(w_n2803_32[1]),.dinb(w_in31_0[0]),.dout(n3760),.clk(gclk));
	jand g3119(.dina(n3760),.dinb(n3759),.dout(n3761),.clk(gclk));
	jand g3120(.dina(w_n1721_32[2]),.dinb(w_n1044_0[0]),.dout(n3762),.clk(gclk));
	jand g3121(.dina(w_n1562_32[2]),.dinb(w_n1586_0[0]),.dout(n3763),.clk(gclk));
	jor g3122(.dina(n3763),.dinb(n3762),.dout(n3764),.clk(gclk));
	jor g3123(.dina(w_n3764_0[1]),.dinb(w_n3761_0[2]),.dout(n3765),.clk(gclk));
	jand g3124(.dina(w_n1721_32[1]),.dinb(w_n1046_0[0]),.dout(n3766),.clk(gclk));
	jand g3125(.dina(w_n1562_32[1]),.dinb(w_n1588_0[0]),.dout(n3767),.clk(gclk));
	jor g3126(.dina(n3767),.dinb(n3766),.dout(n3768),.clk(gclk));
	jor g3127(.dina(w_n2808_32[1]),.dinb(w_in20_0[0]),.dout(n3769),.clk(gclk));
	jor g3128(.dina(w_n2803_32[0]),.dinb(w_in30_0[0]),.dout(n3770),.clk(gclk));
	jand g3129(.dina(n3770),.dinb(n3769),.dout(n3771),.clk(gclk));
	jor g3130(.dina(w_n3771_0[1]),.dinb(n3768),.dout(n3772),.clk(gclk));
	jand g3131(.dina(n3772),.dinb(n3765),.dout(n3773),.clk(gclk));
	jand g3132(.dina(w_n1721_32[0]),.dinb(w_n1049_0[0]),.dout(n3774),.clk(gclk));
	jand g3133(.dina(w_n1562_32[0]),.dinb(w_n1041_0[0]),.dout(n3775),.clk(gclk));
	jor g3134(.dina(n3775),.dinb(n3774),.dout(n3776),.clk(gclk));
	jor g3135(.dina(w_n2808_32[0]),.dinb(w_in22_0[0]),.dout(n3777),.clk(gclk));
	jor g3136(.dina(w_n2803_31[2]),.dinb(w_in32_0[0]),.dout(n3778),.clk(gclk));
	jand g3137(.dina(n3778),.dinb(n3777),.dout(n3779),.clk(gclk));
	jand g3138(.dina(w_n3779_0[2]),.dinb(w_n3776_0[1]),.dout(n3780),.clk(gclk));
	jand g3139(.dina(w_n3764_0[0]),.dinb(w_n3761_0[1]),.dout(n3781),.clk(gclk));
	jor g3140(.dina(n3781),.dinb(n3780),.dout(n3782),.clk(gclk));
	jor g3141(.dina(n3782),.dinb(n3773),.dout(n3783),.clk(gclk));
	jor g3142(.dina(w_n3779_0[1]),.dinb(w_n3776_0[0]),.dout(n3784),.clk(gclk));
	jand g3143(.dina(w_n1721_31[2]),.dinb(w_n1039_0[0]),.dout(n3785),.clk(gclk));
	jand g3144(.dina(w_n1562_31[2]),.dinb(w_n1054_0[0]),.dout(n3786),.clk(gclk));
	jor g3145(.dina(n3786),.dinb(n3785),.dout(n3787),.clk(gclk));
	jand g3146(.dina(w_n2803_31[1]),.dinb(w_n2106_0[0]),.dout(n3788),.clk(gclk));
	jand g3147(.dina(w_n2808_31[2]),.dinb(w_n2120_0[0]),.dout(n3789),.clk(gclk));
	jor g3148(.dina(n3789),.dinb(n3788),.dout(n3790),.clk(gclk));
	jnot g3149(.din(w_n3790_0[1]),.dout(n3791),.clk(gclk));
	jor g3150(.dina(w_n3791_0[2]),.dinb(w_n3787_0[1]),.dout(n3792),.clk(gclk));
	jand g3151(.dina(n3792),.dinb(n3784),.dout(n3793),.clk(gclk));
	jand g3152(.dina(n3793),.dinb(n3783),.dout(n3794),.clk(gclk));
	jnot g3153(.din(w_n3752_0[0]),.dout(n3795),.clk(gclk));
	jand g3154(.dina(w_n3755_0[0]),.dinb(w_n3795_0[1]),.dout(n3796),.clk(gclk));
	jand g3155(.dina(w_n3791_0[1]),.dinb(w_n3787_0[0]),.dout(n3797),.clk(gclk));
	jor g3156(.dina(n3797),.dinb(n3796),.dout(n3798),.clk(gclk));
	jor g3157(.dina(w_n3798_0[1]),.dinb(n3794),.dout(n3799),.clk(gclk));
	jand g3158(.dina(n3799),.dinb(n3758),.dout(n3800),.clk(gclk));
	jor g3159(.dina(n3800),.dinb(w_n3749_0[1]),.dout(n3801),.clk(gclk));
	jand g3160(.dina(n3801),.dinb(n3747),.dout(n3802),.clk(gclk));
	jor g3161(.dina(n3802),.dinb(w_n3738_0[1]),.dout(n3803),.clk(gclk));
	jnot g3162(.din(w_n3725_0[0]),.dout(n3804),.clk(gclk));
	jand g3163(.dina(w_n3728_0[0]),.dinb(w_n3804_0[1]),.dout(n3805),.clk(gclk));
	jnot g3164(.din(w_n3737_0[0]),.dout(n3806),.clk(gclk));
	jand g3165(.dina(w_n3806_0[1]),.dinb(w_n3733_0[0]),.dout(n3807),.clk(gclk));
	jor g3166(.dina(n3807),.dinb(n3805),.dout(n3808),.clk(gclk));
	jnot g3167(.din(w_n3808_0[1]),.dout(n3809),.clk(gclk));
	jand g3168(.dina(n3809),.dinb(n3803),.dout(n3810),.clk(gclk));
	jnot g3169(.din(w_n3716_0[0]),.dout(n3811),.clk(gclk));
	jand g3170(.dina(w_n3719_0[0]),.dinb(w_n3811_0[1]),.dout(n3812),.clk(gclk));
	jor g3171(.dina(w_n3812_0[1]),.dinb(n3810),.dout(n3813),.clk(gclk));
	jor g3172(.dina(n3813),.dinb(w_n3730_0[1]),.dout(n3814),.clk(gclk));
	jand g3173(.dina(w_n2803_31[0]),.dinb(w_n2164_0[0]),.dout(n3815),.clk(gclk));
	jand g3174(.dina(w_n2808_31[1]),.dinb(w_n2157_0[0]),.dout(n3816),.clk(gclk));
	jor g3175(.dina(n3816),.dinb(n3815),.dout(n3817),.clk(gclk));
	jand g3176(.dina(w_n1721_31[1]),.dinb(w_n1096_0[0]),.dout(n3818),.clk(gclk));
	jand g3177(.dina(w_n1562_31[1]),.dinb(w_n1089_0[0]),.dout(n3819),.clk(gclk));
	jor g3178(.dina(n3819),.dinb(n3818),.dout(n3820),.clk(gclk));
	jnot g3179(.din(w_n3820_0[1]),.dout(n3821),.clk(gclk));
	jand g3180(.dina(w_n3821_0[1]),.dinb(w_n3817_0[1]),.dout(n3822),.clk(gclk));
	jnot g3181(.din(w_n3822_0[1]),.dout(n3823),.clk(gclk));
	jand g3182(.dina(n3823),.dinb(n3814),.dout(n3824),.clk(gclk));
	jand g3183(.dina(n3824),.dinb(n3722),.dout(n3825),.clk(gclk));
	jnot g3184(.din(w_n3817_0[0]),.dout(n3826),.clk(gclk));
	jand g3185(.dina(w_n3820_0[0]),.dinb(w_n3826_0[1]),.dout(n3827),.clk(gclk));
	jor g3186(.dina(w_n3827_0[1]),.dinb(n3825),.dout(n3828),.clk(gclk));
	jor g3187(.dina(n3828),.dinb(w_n3713_0[1]),.dout(n3829),.clk(gclk));
	jnot g3188(.din(w_n3708_0[0]),.dout(n3830),.clk(gclk));
	jand g3189(.dina(w_n3711_0[0]),.dinb(w_n3830_0[1]),.dout(n3831),.clk(gclk));
	jand g3190(.dina(w_n1721_31[0]),.dinb(w_n1032_0[0]),.dout(n3832),.clk(gclk));
	jand g3191(.dina(w_n1562_31[0]),.dinb(w_n1029_0[0]),.dout(n3833),.clk(gclk));
	jor g3192(.dina(n3833),.dinb(n3832),.dout(n3834),.clk(gclk));
	jnot g3193(.din(w_n3834_0[1]),.dout(n3835),.clk(gclk));
	jand g3194(.dina(w_n2803_30[2]),.dinb(w_n2099_0[0]),.dout(n3836),.clk(gclk));
	jand g3195(.dina(w_n2808_31[0]),.dinb(w_n2096_0[0]),.dout(n3837),.clk(gclk));
	jor g3196(.dina(n3837),.dinb(n3836),.dout(n3838),.clk(gclk));
	jand g3197(.dina(w_n3838_0[1]),.dinb(w_n3835_0[1]),.dout(n3839),.clk(gclk));
	jor g3198(.dina(n3839),.dinb(n3831),.dout(n3840),.clk(gclk));
	jnot g3199(.din(w_n3840_0[1]),.dout(n3841),.clk(gclk));
	jand g3200(.dina(n3841),.dinb(n3829),.dout(n3842),.clk(gclk));
	jnot g3201(.din(w_n3703_0[0]),.dout(n3843),.clk(gclk));
	jand g3202(.dina(w_n3843_0[1]),.dinb(w_n3699_0[0]),.dout(n3844),.clk(gclk));
	jnot g3203(.din(w_n3838_0[0]),.dout(n3845),.clk(gclk));
	jand g3204(.dina(w_n3845_0[1]),.dinb(w_n3834_0[0]),.dout(n3846),.clk(gclk));
	jor g3205(.dina(n3846),.dinb(n3844),.dout(n3847),.clk(gclk));
	jor g3206(.dina(w_n3847_0[1]),.dinb(n3842),.dout(n3848),.clk(gclk));
	jand g3207(.dina(n3848),.dinb(n3705),.dout(n3849),.clk(gclk));
	jor g3208(.dina(n3849),.dinb(w_n3696_0[1]),.dout(n3850),.clk(gclk));
	jand g3209(.dina(n3850),.dinb(n3694),.dout(n3851),.clk(gclk));
	jor g3210(.dina(n3851),.dinb(w_n3685_0[1]),.dout(n3852),.clk(gclk));
	jnot g3211(.din(w_n3672_0[0]),.dout(n3853),.clk(gclk));
	jand g3212(.dina(w_n3675_0[0]),.dinb(w_n3853_0[1]),.dout(n3854),.clk(gclk));
	jnot g3213(.din(w_n3680_0[0]),.dout(n3855),.clk(gclk));
	jand g3214(.dina(w_n3683_0[0]),.dinb(w_n3855_0[1]),.dout(n3856),.clk(gclk));
	jor g3215(.dina(n3856),.dinb(n3854),.dout(n3857),.clk(gclk));
	jnot g3216(.din(w_n3857_0[1]),.dout(n3858),.clk(gclk));
	jand g3217(.dina(n3858),.dinb(n3852),.dout(n3859),.clk(gclk));
	jnot g3218(.din(w_n3663_0[0]),.dout(n3860),.clk(gclk));
	jand g3219(.dina(w_n3666_0[0]),.dinb(w_n3860_0[1]),.dout(n3861),.clk(gclk));
	jor g3220(.dina(w_n3861_0[1]),.dinb(n3859),.dout(n3862),.clk(gclk));
	jor g3221(.dina(n3862),.dinb(w_n3677_0[1]),.dout(n3863),.clk(gclk));
	jand g3222(.dina(w_n2803_30[1]),.dinb(w_n2196_0[0]),.dout(n3864),.clk(gclk));
	jand g3223(.dina(w_n2808_30[2]),.dinb(w_n2189_0[0]),.dout(n3865),.clk(gclk));
	jor g3224(.dina(n3865),.dinb(n3864),.dout(n3866),.clk(gclk));
	jand g3225(.dina(w_n1721_30[2]),.dinb(w_n1128_0[0]),.dout(n3867),.clk(gclk));
	jand g3226(.dina(w_n1562_30[2]),.dinb(w_n1121_0[0]),.dout(n3868),.clk(gclk));
	jor g3227(.dina(n3868),.dinb(n3867),.dout(n3869),.clk(gclk));
	jnot g3228(.din(w_n3869_0[1]),.dout(n3870),.clk(gclk));
	jand g3229(.dina(w_n3870_0[1]),.dinb(w_n3866_0[1]),.dout(n3871),.clk(gclk));
	jnot g3230(.din(w_n3871_0[1]),.dout(n3872),.clk(gclk));
	jand g3231(.dina(n3872),.dinb(n3863),.dout(n3873),.clk(gclk));
	jand g3232(.dina(n3873),.dinb(n3669),.dout(n3874),.clk(gclk));
	jnot g3233(.din(w_n3866_0[0]),.dout(n3875),.clk(gclk));
	jand g3234(.dina(w_n3869_0[0]),.dinb(w_n3875_0[1]),.dout(n3876),.clk(gclk));
	jor g3235(.dina(w_n3876_0[1]),.dinb(n3874),.dout(n3877),.clk(gclk));
	jor g3236(.dina(n3877),.dinb(w_n3660_0[1]),.dout(n3878),.clk(gclk));
	jnot g3237(.din(w_n3655_0[0]),.dout(n3879),.clk(gclk));
	jand g3238(.dina(w_n3658_0[0]),.dinb(w_n3879_0[1]),.dout(n3880),.clk(gclk));
	jnot g3239(.din(w_n3647_0[0]),.dout(n3881),.clk(gclk));
	jand g3240(.dina(w_n3650_0[0]),.dinb(w_n3881_0[1]),.dout(n3882),.clk(gclk));
	jor g3241(.dina(n3882),.dinb(n3880),.dout(n3883),.clk(gclk));
	jnot g3242(.din(w_n3883_0[1]),.dout(n3884),.clk(gclk));
	jand g3243(.dina(n3884),.dinb(n3878),.dout(n3885),.clk(gclk));
	jor g3244(.dina(n3885),.dinb(w_n3652_0[1]),.dout(n3886),.clk(gclk));
	jand g3245(.dina(n3886),.dinb(n3644),.dout(n3887),.clk(gclk));
	jand g3246(.dina(w_n1721_30[1]),.dinb(w_n1000_0[0]),.dout(n3888),.clk(gclk));
	jand g3247(.dina(w_n1562_30[1]),.dinb(w_n997_0[0]),.dout(n3889),.clk(gclk));
	jor g3248(.dina(n3889),.dinb(n3888),.dout(n3890),.clk(gclk));
	jand g3249(.dina(w_n2803_30[0]),.dinb(w_n2067_0[0]),.dout(n3891),.clk(gclk));
	jand g3250(.dina(w_n2808_30[1]),.dinb(w_n2064_0[0]),.dout(n3892),.clk(gclk));
	jor g3251(.dina(n3892),.dinb(n3891),.dout(n3893),.clk(gclk));
	jnot g3252(.din(w_n3893_0[1]),.dout(n3894),.clk(gclk));
	jand g3253(.dina(w_n3894_0[1]),.dinb(w_n3890_0[1]),.dout(n3895),.clk(gclk));
	jor g3254(.dina(w_n3895_0[1]),.dinb(n3887),.dout(n3896),.clk(gclk));
	jor g3255(.dina(n3896),.dinb(w_n3641_0[1]),.dout(n3897),.clk(gclk));
	jnot g3256(.din(w_n3890_0[0]),.dout(n3898),.clk(gclk));
	jand g3257(.dina(w_n3893_0[0]),.dinb(w_n3898_0[1]),.dout(n3899),.clk(gclk));
	jnot g3258(.din(w_n3628_0[0]),.dout(n3900),.clk(gclk));
	jand g3259(.dina(w_n3631_0[0]),.dinb(w_n3900_0[1]),.dout(n3901),.clk(gclk));
	jor g3260(.dina(n3901),.dinb(n3899),.dout(n3902),.clk(gclk));
	jnot g3261(.din(w_n3902_0[1]),.dout(n3903),.clk(gclk));
	jand g3262(.dina(n3903),.dinb(n3897),.dout(n3904),.clk(gclk));
	jor g3263(.dina(n3904),.dinb(w_n3633_0[1]),.dout(n3905),.clk(gclk));
	jand g3264(.dina(n3905),.dinb(n3625),.dout(n3906),.clk(gclk));
	jnot g3265(.din(w_n3623_0[0]),.dout(n3907),.clk(gclk));
	jand g3266(.dina(w_n3907_0[1]),.dinb(w_n3619_0[0]),.dout(n3908),.clk(gclk));
	jnot g3267(.din(w_n3601_0[0]),.dout(n3909),.clk(gclk));
	jand g3268(.dina(w_n3604_0[0]),.dinb(w_n3909_0[1]),.dout(n3910),.clk(gclk));
	jor g3269(.dina(n3910),.dinb(n3908),.dout(n3911),.clk(gclk));
	jor g3270(.dina(w_n3911_0[1]),.dinb(n3906),.dout(n3912),.clk(gclk));
	jand g3271(.dina(n3912),.dinb(n3616),.dout(n3913),.clk(gclk));
	jnot g3272(.din(w_n3609_0[0]),.dout(n3914),.clk(gclk));
	jand g3273(.dina(w_n3612_0[0]),.dinb(w_n3914_0[1]),.dout(n3915),.clk(gclk));
	jor g3274(.dina(w_n3915_0[1]),.dinb(n3913),.dout(n3916),.clk(gclk));
	jor g3275(.dina(n3916),.dinb(w_n3598_0[1]),.dout(n3917),.clk(gclk));
	jnot g3276(.din(w_n3593_0[0]),.dout(n3918),.clk(gclk));
	jand g3277(.dina(w_n3596_0[0]),.dinb(w_n3918_0[1]),.dout(n3919),.clk(gclk));
	jand g3278(.dina(w_n1721_30[0]),.dinb(w_n988_0[0]),.dout(n3920),.clk(gclk));
	jand g3279(.dina(w_n1562_30[0]),.dinb(w_n985_0[0]),.dout(n3921),.clk(gclk));
	jor g3280(.dina(n3921),.dinb(n3920),.dout(n3922),.clk(gclk));
	jnot g3281(.din(w_n3922_0[1]),.dout(n3923),.clk(gclk));
	jand g3282(.dina(w_n2803_29[2]),.dinb(w_n2055_0[0]),.dout(n3924),.clk(gclk));
	jand g3283(.dina(w_n2808_30[0]),.dinb(w_n2052_0[0]),.dout(n3925),.clk(gclk));
	jor g3284(.dina(n3925),.dinb(n3924),.dout(n3926),.clk(gclk));
	jand g3285(.dina(w_n3926_0[1]),.dinb(w_n3923_0[1]),.dout(n3927),.clk(gclk));
	jor g3286(.dina(n3927),.dinb(n3919),.dout(n3928),.clk(gclk));
	jnot g3287(.din(w_n3928_0[1]),.dout(n3929),.clk(gclk));
	jand g3288(.dina(n3929),.dinb(n3917),.dout(n3930),.clk(gclk));
	jnot g3289(.din(w_n3588_0[0]),.dout(n3931),.clk(gclk));
	jand g3290(.dina(w_n3931_0[1]),.dinb(w_n3584_0[0]),.dout(n3932),.clk(gclk));
	jnot g3291(.din(w_n3926_0[0]),.dout(n3933),.clk(gclk));
	jand g3292(.dina(w_n3933_0[1]),.dinb(w_n3922_0[0]),.dout(n3934),.clk(gclk));
	jor g3293(.dina(n3934),.dinb(n3932),.dout(n3935),.clk(gclk));
	jor g3294(.dina(w_n3935_0[1]),.dinb(n3930),.dout(n3936),.clk(gclk));
	jand g3295(.dina(n3936),.dinb(n3590),.dout(n3937),.clk(gclk));
	jor g3296(.dina(n3937),.dinb(w_n3581_0[1]),.dout(n3938),.clk(gclk));
	jand g3297(.dina(w_n1721_29[2]),.dinb(w_n973_0[0]),.dout(n3939),.clk(gclk));
	jand g3298(.dina(w_n1562_29[2]),.dinb(w_n1174_0[0]),.dout(n3940),.clk(gclk));
	jor g3299(.dina(n3940),.dinb(n3939),.dout(n3941),.clk(gclk));
	jnot g3300(.din(w_n3941_0[1]),.dout(n3942),.clk(gclk));
	jand g3301(.dina(w_n2803_29[1]),.dinb(w_n2040_0[0]),.dout(n3943),.clk(gclk));
	jand g3302(.dina(w_n2808_29[2]),.dinb(w_n2242_0[0]),.dout(n3944),.clk(gclk));
	jor g3303(.dina(n3944),.dinb(n3943),.dout(n3945),.clk(gclk));
	jand g3304(.dina(w_n3945_0[1]),.dinb(w_n3942_0[1]),.dout(n3946),.clk(gclk));
	jnot g3305(.din(w_n3576_0[0]),.dout(n3947),.clk(gclk));
	jand g3306(.dina(w_n3579_0[0]),.dinb(w_n3947_0[1]),.dout(n3948),.clk(gclk));
	jor g3307(.dina(n3948),.dinb(n3946),.dout(n3949),.clk(gclk));
	jnot g3308(.din(w_n3949_0[1]),.dout(n3950),.clk(gclk));
	jand g3309(.dina(n3950),.dinb(n3938),.dout(n3951),.clk(gclk));
	jnot g3310(.din(w_n3571_0[0]),.dout(n3952),.clk(gclk));
	jand g3311(.dina(w_n3952_0[1]),.dinb(w_n3567_0[0]),.dout(n3953),.clk(gclk));
	jnot g3312(.din(w_n3945_0[0]),.dout(n3954),.clk(gclk));
	jand g3313(.dina(w_n3954_0[1]),.dinb(w_n3941_0[0]),.dout(n3955),.clk(gclk));
	jor g3314(.dina(n3955),.dinb(n3953),.dout(n3956),.clk(gclk));
	jor g3315(.dina(w_n3956_0[1]),.dinb(n3951),.dout(n3957),.clk(gclk));
	jand g3316(.dina(n3957),.dinb(n3573),.dout(n3958),.clk(gclk));
	jand g3317(.dina(w_n3507_0[0]),.dinb(w_n3475_0[0]),.dout(n3959),.clk(gclk));
	jnot g3318(.din(w_n3537_0[0]),.dout(n3960),.clk(gclk));
	jand g3319(.dina(w_n3540_0[0]),.dinb(w_n3960_0[1]),.dout(n3961),.clk(gclk));
	jor g3320(.dina(n3961),.dinb(w_n3515_0[0]),.dout(n3962),.clk(gclk));
	jnot g3321(.din(n3962),.dout(n3963),.clk(gclk));
	jand g3322(.dina(n3963),.dinb(n3959),.dout(n3964),.clk(gclk));
	jand g3323(.dina(n3964),.dinb(w_n3493_0[0]),.dout(n3965),.clk(gclk));
	jnot g3324(.din(w_n3965_0[1]),.dout(n3966),.clk(gclk));
	jor g3325(.dina(n3966),.dinb(n3958),.dout(n3967),.clk(gclk));
	jor g3326(.dina(n3967),.dinb(w_n3533_0[0]),.dout(n3968),.clk(gclk));
	jand g3327(.dina(n3968),.dinb(n3564),.dout(n3969),.clk(gclk));
	jand g3328(.dina(w_n1721_29[1]),.dinb(w_n931_0[0]),.dout(n3970),.clk(gclk));
	jand g3329(.dina(w_n1562_29[1]),.dinb(w_n929_0[0]),.dout(n3971),.clk(gclk));
	jor g3330(.dina(n3971),.dinb(n3970),.dout(n3972),.clk(gclk));
	jand g3331(.dina(w_n2803_29[0]),.dinb(w_n2281_0[0]),.dout(n3973),.clk(gclk));
	jand g3332(.dina(w_n2808_29[1]),.dinb(w_n2295_0[0]),.dout(n3974),.clk(gclk));
	jor g3333(.dina(n3974),.dinb(n3973),.dout(n3975),.clk(gclk));
	jnot g3334(.din(w_n3975_0[1]),.dout(n3976),.clk(gclk));
	jand g3335(.dina(w_n3976_0[1]),.dinb(w_n3972_0[1]),.dout(n3977),.clk(gclk));
	jand g3336(.dina(w_n1721_29[0]),.dinb(w_n1210_0[0]),.dout(n3978),.clk(gclk));
	jand g3337(.dina(w_n1562_29[0]),.dinb(w_n934_0[0]),.dout(n3979),.clk(gclk));
	jor g3338(.dina(n3979),.dinb(n3978),.dout(n3980),.clk(gclk));
	jand g3339(.dina(w_n2803_28[2]),.dinb(w_n2278_0[0]),.dout(n3981),.clk(gclk));
	jand g3340(.dina(w_n2808_29[0]),.dinb(w_n2300_0[0]),.dout(n3982),.clk(gclk));
	jor g3341(.dina(n3982),.dinb(n3981),.dout(n3983),.clk(gclk));
	jnot g3342(.din(w_n3983_0[1]),.dout(n3984),.clk(gclk));
	jand g3343(.dina(w_n3984_0[1]),.dinb(w_n3980_0[1]),.dout(n3985),.clk(gclk));
	jand g3344(.dina(w_n1721_28[2]),.dinb(w_n920_0[0]),.dout(n3986),.clk(gclk));
	jand g3345(.dina(w_n1562_28[2]),.dinb(w_n927_0[0]),.dout(n3987),.clk(gclk));
	jor g3346(.dina(n3987),.dinb(n3986),.dout(n3988),.clk(gclk));
	jand g3347(.dina(w_n2803_28[1]),.dinb(w_n2284_0[0]),.dout(n3989),.clk(gclk));
	jand g3348(.dina(w_n2808_28[2]),.dinb(w_n2297_0[0]),.dout(n3990),.clk(gclk));
	jor g3349(.dina(n3990),.dinb(n3989),.dout(n3991),.clk(gclk));
	jnot g3350(.din(w_n3991_0[1]),.dout(n3992),.clk(gclk));
	jand g3351(.dina(w_n3992_0[1]),.dinb(w_n3988_0[1]),.dout(n3993),.clk(gclk));
	jnot g3352(.din(n3993),.dout(n3994),.clk(gclk));
	jor g3353(.dina(w_n3463_0[1]),.dinb(w_n3421_0[1]),.dout(n3995),.clk(gclk));
	jand g3354(.dina(n3995),.dinb(n3994),.dout(n3996),.clk(gclk));
	jand g3355(.dina(n3996),.dinb(w_n3459_0[0]),.dout(n3997),.clk(gclk));
	jnot g3356(.din(w_n3997_0[1]),.dout(n3998),.clk(gclk));
	jor g3357(.dina(n3998),.dinb(n3985),.dout(n3999),.clk(gclk));
	jor g3358(.dina(n3999),.dinb(w_n3977_0[1]),.dout(n4000),.clk(gclk));
	jor g3359(.dina(w_n4000_0[1]),.dinb(n3969),.dout(n4001),.clk(gclk));
	jnot g3360(.din(w_n3988_0[0]),.dout(n4002),.clk(gclk));
	jand g3361(.dina(w_n3991_0[0]),.dinb(w_n4002_0[1]),.dout(n4003),.clk(gclk));
	jnot g3362(.din(w_n3977_0[0]),.dout(n4004),.clk(gclk));
	jnot g3363(.din(w_n3980_0[0]),.dout(n4005),.clk(gclk));
	jand g3364(.dina(w_n3983_0[0]),.dinb(w_n4005_0[1]),.dout(n4006),.clk(gclk));
	jand g3365(.dina(n4006),.dinb(n4004),.dout(n4007),.clk(gclk));
	jnot g3366(.din(w_n3972_0[0]),.dout(n4008),.clk(gclk));
	jand g3367(.dina(w_n3975_0[0]),.dinb(w_n4008_0[1]),.dout(n4009),.clk(gclk));
	jor g3368(.dina(n4009),.dinb(n4007),.dout(n4010),.clk(gclk));
	jor g3369(.dina(n4010),.dinb(n4003),.dout(n4011),.clk(gclk));
	jand g3370(.dina(n4011),.dinb(w_n3997_0[0]),.dout(n4012),.clk(gclk));
	jnot g3371(.din(w_n3451_0[0]),.dout(n4013),.clk(gclk));
	jand g3372(.dina(w_n3454_0[0]),.dinb(w_n4013_0[1]),.dout(n4014),.clk(gclk));
	jnot g3373(.din(w_n3424_0[0]),.dout(n4015),.clk(gclk));
	jand g3374(.dina(w_n3427_0[0]),.dinb(w_n4015_0[1]),.dout(n4016),.clk(gclk));
	jor g3375(.dina(n4016),.dinb(n4014),.dout(n4017),.clk(gclk));
	jand g3376(.dina(n4017),.dinb(w_n3457_0[0]),.dout(n4018),.clk(gclk));
	jand g3377(.dina(n4018),.dinb(w_n3448_0[0]),.dout(n4019),.clk(gclk));
	jnot g3378(.din(w_n3438_0[0]),.dout(n4020),.clk(gclk));
	jnot g3379(.din(w_n3433_0[0]),.dout(n4021),.clk(gclk));
	jand g3380(.dina(w_n3436_0[0]),.dinb(w_n4021_0[1]),.dout(n4022),.clk(gclk));
	jnot g3381(.din(w_n3445_0[0]),.dout(n4023),.clk(gclk));
	jand g3382(.dina(w_n4023_0[1]),.dinb(w_n3441_0[0]),.dout(n4024),.clk(gclk));
	jor g3383(.dina(n4024),.dinb(n4022),.dout(n4025),.clk(gclk));
	jand g3384(.dina(n4025),.dinb(n4020),.dout(n4026),.clk(gclk));
	jor g3385(.dina(n4026),.dinb(n4019),.dout(n4027),.clk(gclk));
	jor g3386(.dina(n4027),.dinb(n4012),.dout(n4028),.clk(gclk));
	jnot g3387(.din(w_n4028_0[1]),.dout(n4029),.clk(gclk));
	jand g3388(.dina(n4029),.dinb(n4001),.dout(n4030),.clk(gclk));
	jand g3389(.dina(n4030),.dinb(n3466),.dout(n4031),.clk(gclk));
	jand g3390(.dina(w_n1721_28[1]),.dinb(w_n1239_0[0]),.dout(n4032),.clk(gclk));
	jand g3391(.dina(w_n1562_28[1]),.dinb(w_n1253_0[0]),.dout(n4033),.clk(gclk));
	jor g3392(.dina(n4033),.dinb(n4032),.dout(n4034),.clk(gclk));
	jand g3393(.dina(w_n2803_28[0]),.dinb(w_n2327_0[0]),.dout(n4035),.clk(gclk));
	jand g3394(.dina(w_n2808_28[1]),.dinb(w_n2341_0[0]),.dout(n4036),.clk(gclk));
	jor g3395(.dina(n4036),.dinb(n4035),.dout(n4037),.clk(gclk));
	jnot g3396(.din(w_n4037_0[1]),.dout(n4038),.clk(gclk));
	jand g3397(.dina(w_n4038_0[1]),.dinb(w_n4034_0[1]),.dout(n4039),.clk(gclk));
	jand g3398(.dina(w_n2803_27[2]),.dinb(w_n2330_0[0]),.dout(n4040),.clk(gclk));
	jand g3399(.dina(w_n2808_28[0]),.dinb(w_n2343_0[0]),.dout(n4041),.clk(gclk));
	jor g3400(.dina(n4041),.dinb(n4040),.dout(n4042),.clk(gclk));
	jnot g3401(.din(w_n4042_0[1]),.dout(n4043),.clk(gclk));
	jand g3402(.dina(w_n1721_28[0]),.dinb(w_n1242_0[0]),.dout(n4044),.clk(gclk));
	jand g3403(.dina(w_n1562_28[0]),.dinb(w_n1255_0[0]),.dout(n4045),.clk(gclk));
	jor g3404(.dina(n4045),.dinb(n4044),.dout(n4046),.clk(gclk));
	jand g3405(.dina(w_n4046_0[1]),.dinb(w_n4043_0[1]),.dout(n4047),.clk(gclk));
	jor g3406(.dina(n4047),.dinb(n4039),.dout(n4048),.clk(gclk));
	jand g3407(.dina(w_n2803_27[1]),.dinb(w_n1984_0[0]),.dout(n4049),.clk(gclk));
	jand g3408(.dina(w_n2808_27[2]),.dinb(w_n2355_0[0]),.dout(n4050),.clk(gclk));
	jor g3409(.dina(n4050),.dinb(n4049),.dout(n4051),.clk(gclk));
	jnot g3410(.din(w_n4051_0[1]),.dout(n4052),.clk(gclk));
	jand g3411(.dina(w_n1721_27[2]),.dinb(w_n901_0[0]),.dout(n4053),.clk(gclk));
	jand g3412(.dina(w_n1562_27[2]),.dinb(w_n1267_0[0]),.dout(n4054),.clk(gclk));
	jor g3413(.dina(n4054),.dinb(n4053),.dout(n4055),.clk(gclk));
	jand g3414(.dina(w_n4055_0[1]),.dinb(w_n4052_0[1]),.dout(n4056),.clk(gclk));
	jand g3415(.dina(w_n1721_27[1]),.dinb(w_n894_0[0]),.dout(n4057),.clk(gclk));
	jand g3416(.dina(w_n1562_27[1]),.dinb(w_n1272_0[0]),.dout(n4058),.clk(gclk));
	jor g3417(.dina(n4058),.dinb(n4057),.dout(n4059),.clk(gclk));
	jand g3418(.dina(w_n2803_27[0]),.dinb(w_n1977_0[0]),.dout(n4060),.clk(gclk));
	jand g3419(.dina(w_n2808_27[1]),.dinb(w_n2360_0[0]),.dout(n4061),.clk(gclk));
	jor g3420(.dina(n4061),.dinb(n4060),.dout(n4062),.clk(gclk));
	jnot g3421(.din(w_n4062_0[1]),.dout(n4063),.clk(gclk));
	jand g3422(.dina(w_n4063_0[1]),.dinb(w_n4059_0[1]),.dout(n4064),.clk(gclk));
	jor g3423(.dina(n4064),.dinb(n4056),.dout(n4065),.clk(gclk));
	jnot g3424(.din(w_n3416_0[0]),.dout(n4066),.clk(gclk));
	jand g3425(.dina(w_n4066_0[1]),.dinb(w_n3412_0[0]),.dout(n4067),.clk(gclk));
	jand g3426(.dina(w_n2803_26[2]),.dinb(w_n1981_0[0]),.dout(n4068),.clk(gclk));
	jand g3427(.dina(w_n2808_27[0]),.dinb(w_n2358_0[0]),.dout(n4069),.clk(gclk));
	jor g3428(.dina(n4069),.dinb(n4068),.dout(n4070),.clk(gclk));
	jnot g3429(.din(w_n4070_0[1]),.dout(n4071),.clk(gclk));
	jand g3430(.dina(w_n1721_27[0]),.dinb(w_n898_0[0]),.dout(n4072),.clk(gclk));
	jand g3431(.dina(w_n1562_27[0]),.dinb(w_n1270_0[0]),.dout(n4073),.clk(gclk));
	jor g3432(.dina(n4073),.dinb(n4072),.dout(n4074),.clk(gclk));
	jand g3433(.dina(w_n4074_0[1]),.dinb(w_n4071_0[1]),.dout(n4075),.clk(gclk));
	jor g3434(.dina(n4075),.dinb(n4067),.dout(n4076),.clk(gclk));
	jand g3435(.dina(w_n2803_26[1]),.dinb(w_n2324_0[0]),.dout(n4077),.clk(gclk));
	jand g3436(.dina(w_n2808_26[2]),.dinb(w_n2346_0[0]),.dout(n4078),.clk(gclk));
	jor g3437(.dina(n4078),.dinb(n4077),.dout(n4079),.clk(gclk));
	jnot g3438(.din(w_n4079_0[1]),.dout(n4080),.clk(gclk));
	jand g3439(.dina(w_n1721_26[2]),.dinb(w_n1236_0[0]),.dout(n4081),.clk(gclk));
	jand g3440(.dina(w_n1562_26[2]),.dinb(w_n1258_0[0]),.dout(n4082),.clk(gclk));
	jor g3441(.dina(n4082),.dinb(n4081),.dout(n4083),.clk(gclk));
	jand g3442(.dina(w_n4083_0[1]),.dinb(w_n4080_0[1]),.dout(n4084),.clk(gclk));
	jand g3443(.dina(w_n1721_26[1]),.dinb(w_n1244_0[0]),.dout(n4085),.clk(gclk));
	jand g3444(.dina(w_n1562_26[1]),.dinb(w_n893_0[0]),.dout(n4086),.clk(gclk));
	jor g3445(.dina(n4086),.dinb(n4085),.dout(n4087),.clk(gclk));
	jand g3446(.dina(w_n2803_26[0]),.dinb(w_n2332_0[0]),.dout(n4088),.clk(gclk));
	jand g3447(.dina(w_n2808_26[1]),.dinb(w_n1976_0[0]),.dout(n4089),.clk(gclk));
	jor g3448(.dina(n4089),.dinb(n4088),.dout(n4090),.clk(gclk));
	jnot g3449(.din(w_n4090_0[1]),.dout(n4091),.clk(gclk));
	jand g3450(.dina(w_n4091_0[1]),.dinb(w_n4087_0[1]),.dout(n4092),.clk(gclk));
	jor g3451(.dina(w_n4092_0[1]),.dinb(n4084),.dout(n4093),.clk(gclk));
	jor g3452(.dina(n4093),.dinb(w_n4076_0[1]),.dout(n4094),.clk(gclk));
	jor g3453(.dina(n4094),.dinb(w_n4065_0[1]),.dout(n4095),.clk(gclk));
	jor g3454(.dina(n4095),.dinb(w_n4048_0[1]),.dout(n4096),.clk(gclk));
	jor g3455(.dina(w_n4096_0[1]),.dinb(n4031),.dout(n4097),.clk(gclk));
	jnot g3456(.din(w_n4076_0[0]),.dout(n4098),.clk(gclk));
	jnot g3457(.din(w_n4059_0[0]),.dout(n4099),.clk(gclk));
	jand g3458(.dina(w_n4062_0[0]),.dinb(w_n4099_0[1]),.dout(n4100),.clk(gclk));
	jnot g3459(.din(w_n4074_0[0]),.dout(n4101),.clk(gclk));
	jand g3460(.dina(w_n4101_0[1]),.dinb(w_n4070_0[0]),.dout(n4102),.clk(gclk));
	jnot g3461(.din(w_n4065_0[0]),.dout(n4103),.clk(gclk));
	jnot g3462(.din(w_n4055_0[0]),.dout(n4104),.clk(gclk));
	jand g3463(.dina(w_n4104_0[1]),.dinb(w_n4051_0[0]),.dout(n4105),.clk(gclk));
	jnot g3464(.din(w_n4092_0[0]),.dout(n4106),.clk(gclk));
	jnot g3465(.din(w_n4048_0[0]),.dout(n4107),.clk(gclk));
	jnot g3466(.din(w_n4083_0[0]),.dout(n4108),.clk(gclk));
	jand g3467(.dina(w_n4108_0[1]),.dinb(w_n4079_0[0]),.dout(n4109),.clk(gclk));
	jnot g3468(.din(w_n4034_0[0]),.dout(n4110),.clk(gclk));
	jand g3469(.dina(w_n4037_0[0]),.dinb(w_n4110_0[1]),.dout(n4111),.clk(gclk));
	jor g3470(.dina(n4111),.dinb(n4109),.dout(n4112),.clk(gclk));
	jand g3471(.dina(n4112),.dinb(n4107),.dout(n4113),.clk(gclk));
	jnot g3472(.din(w_n4087_0[0]),.dout(n4114),.clk(gclk));
	jand g3473(.dina(w_n4090_0[0]),.dinb(w_n4114_0[1]),.dout(n4115),.clk(gclk));
	jnot g3474(.din(w_n4046_0[0]),.dout(n4116),.clk(gclk));
	jand g3475(.dina(w_n4116_0[1]),.dinb(w_n4042_0[0]),.dout(n4117),.clk(gclk));
	jor g3476(.dina(n4117),.dinb(n4115),.dout(n4118),.clk(gclk));
	jor g3477(.dina(n4118),.dinb(n4113),.dout(n4119),.clk(gclk));
	jand g3478(.dina(n4119),.dinb(n4106),.dout(n4120),.clk(gclk));
	jor g3479(.dina(n4120),.dinb(n4105),.dout(n4121),.clk(gclk));
	jand g3480(.dina(n4121),.dinb(n4103),.dout(n4122),.clk(gclk));
	jor g3481(.dina(n4122),.dinb(n4102),.dout(n4123),.clk(gclk));
	jor g3482(.dina(n4123),.dinb(n4100),.dout(n4124),.clk(gclk));
	jand g3483(.dina(n4124),.dinb(n4098),.dout(n4125),.clk(gclk));
	jnot g3484(.din(w_n4125_0[1]),.dout(n4126),.clk(gclk));
	jand g3485(.dina(n4126),.dinb(n4097),.dout(n4127),.clk(gclk));
	jand g3486(.dina(n4127),.dinb(n3418),.dout(n4128),.clk(gclk));
	jnot g3487(.din(w_n3399_0[0]),.dout(n4129),.clk(gclk));
	jand g3488(.dina(w_n4129_0[1]),.dinb(w_n3395_0[0]),.dout(n4130),.clk(gclk));
	jor g3489(.dina(n4130),.dinb(w_n3391_0[0]),.dout(n4131),.clk(gclk));
	jor g3490(.dina(n4131),.dinb(w_n3380_0[0]),.dout(n4132),.clk(gclk));
	jor g3491(.dina(n4132),.dinb(w_n3360_0[0]),.dout(n4133),.clk(gclk));
	jor g3492(.dina(w_n4133_0[1]),.dinb(n4128),.dout(n4134),.clk(gclk));
	jnot g3493(.din(w_n3359_0[0]),.dout(n4135),.clk(gclk));
	jnot g3494(.din(w_n3352_0[0]),.dout(n4136),.clk(gclk));
	jand g3495(.dina(w_n3355_0[0]),.dinb(w_n4136_0[1]),.dout(n4137),.clk(gclk));
	jnot g3496(.din(w_n3328_0[0]),.dout(n4138),.clk(gclk));
	jand g3497(.dina(w_n3331_0[0]),.dinb(w_n4138_0[1]),.dout(n4139),.clk(gclk));
	jor g3498(.dina(n4139),.dinb(n4137),.dout(n4140),.clk(gclk));
	jand g3499(.dina(n4140),.dinb(n4135),.dout(n4141),.clk(gclk));
	jnot g3500(.din(w_n3349_0[0]),.dout(n4142),.clk(gclk));
	jnot g3501(.din(w_n3344_0[0]),.dout(n4143),.clk(gclk));
	jand g3502(.dina(w_n3347_0[0]),.dinb(w_n4143_0[1]),.dout(n4144),.clk(gclk));
	jnot g3503(.din(w_n3340_0[0]),.dout(n4145),.clk(gclk));
	jand g3504(.dina(w_n4145_0[1]),.dinb(w_n3336_0[0]),.dout(n4146),.clk(gclk));
	jor g3505(.dina(n4146),.dinb(n4144),.dout(n4147),.clk(gclk));
	jand g3506(.dina(n4147),.dinb(n4142),.dout(n4148),.clk(gclk));
	jor g3507(.dina(n4148),.dinb(n4141),.dout(n4149),.clk(gclk));
	jnot g3508(.din(w_n4149_0[1]),.dout(n4150),.clk(gclk));
	jand g3509(.dina(n4150),.dinb(n4134),.dout(n4151),.clk(gclk));
	jand g3510(.dina(n4151),.dinb(n3409),.dout(n4152),.clk(gclk));
	jnot g3511(.din(w_n3316_0[0]),.dout(n4153),.clk(gclk));
	jand g3512(.dina(w_n3319_0[0]),.dinb(w_n4153_0[1]),.dout(n4154),.clk(gclk));
	jor g3513(.dina(n4154),.dinb(w_n3312_0[0]),.dout(n4155),.clk(gclk));
	jor g3514(.dina(w_n4155_0[1]),.dinb(n4152),.dout(n4156),.clk(gclk));
	jand g3515(.dina(n4156),.dinb(n3325),.dout(n4157),.clk(gclk));
	jnot g3516(.din(w_n3292_0[0]),.dout(n4158),.clk(gclk));
	jand g3517(.dina(w_n4158_0[1]),.dinb(w_n3288_0[0]),.dout(n4159),.clk(gclk));
	jnot g3518(.din(w_n3297_0[0]),.dout(n4160),.clk(gclk));
	jand g3519(.dina(w_n3300_0[0]),.dinb(w_n4160_0[1]),.dout(n4161),.clk(gclk));
	jor g3520(.dina(n4161),.dinb(n4159),.dout(n4162),.clk(gclk));
	jor g3521(.dina(w_n4162_0[1]),.dinb(n4157),.dout(n4163),.clk(gclk));
	jand g3522(.dina(n4163),.dinb(n3294),.dout(n4164),.clk(gclk));
	jnot g3523(.din(w_n3273_0[0]),.dout(n4165),.clk(gclk));
	jand g3524(.dina(w_n4165_0[1]),.dinb(w_n3269_0[0]),.dout(n4166),.clk(gclk));
	jor g3525(.dina(n4166),.dinb(w_n3263_0[0]),.dout(n4167),.clk(gclk));
	jor g3526(.dina(w_n4167_0[1]),.dinb(n4164),.dout(n4168),.clk(gclk));
	jand g3527(.dina(n4168),.dinb(n3285),.dout(n4169),.clk(gclk));
	jand g3528(.dina(w_n2803_25[2]),.dinb(w_n2438_0[0]),.dout(n4170),.clk(gclk));
	jand g3529(.dina(w_n2808_26[0]),.dinb(w_n2452_0[0]),.dout(n4171),.clk(gclk));
	jor g3530(.dina(n4171),.dinb(n4170),.dout(n4172),.clk(gclk));
	jnot g3531(.din(w_n4172_0[1]),.dout(n4173),.clk(gclk));
	jand g3532(.dina(w_n1721_26[0]),.dinb(w_n832_0[0]),.dout(n4174),.clk(gclk));
	jand g3533(.dina(w_n1562_26[0]),.dinb(w_n1359_0[0]),.dout(n4175),.clk(gclk));
	jor g3534(.dina(n4175),.dinb(n4174),.dout(n4176),.clk(gclk));
	jand g3535(.dina(w_n4176_0[1]),.dinb(w_n4173_0[1]),.dout(n4177),.clk(gclk));
	jnot g3536(.din(n4177),.dout(n4178),.clk(gclk));
	jand g3537(.dina(w_n1721_25[2]),.dinb(w_n1345_0[0]),.dout(n4179),.clk(gclk));
	jand g3538(.dina(w_n1562_25[2]),.dinb(w_n829_0[0]),.dout(n4180),.clk(gclk));
	jor g3539(.dina(n4180),.dinb(n4179),.dout(n4181),.clk(gclk));
	jand g3540(.dina(w_n2803_25[1]),.dinb(w_n2433_0[0]),.dout(n4182),.clk(gclk));
	jand g3541(.dina(w_n2808_25[2]),.dinb(w_n1917_0[0]),.dout(n4183),.clk(gclk));
	jor g3542(.dina(n4183),.dinb(n4182),.dout(n4184),.clk(gclk));
	jnot g3543(.din(w_n4184_0[1]),.dout(n4185),.clk(gclk));
	jand g3544(.dina(w_n4185_0[1]),.dinb(w_n4181_0[1]),.dout(n4186),.clk(gclk));
	jand g3545(.dina(w_n2803_25[0]),.dinb(w_n2435_0[0]),.dout(n4187),.clk(gclk));
	jand g3546(.dina(w_n2808_25[1]),.dinb(w_n2448_0[0]),.dout(n4188),.clk(gclk));
	jor g3547(.dina(n4188),.dinb(n4187),.dout(n4189),.clk(gclk));
	jnot g3548(.din(w_n4189_0[1]),.dout(n4190),.clk(gclk));
	jand g3549(.dina(w_n1721_25[1]),.dinb(w_n1347_0[0]),.dout(n4191),.clk(gclk));
	jand g3550(.dina(w_n1562_25[1]),.dinb(w_n1355_0[0]),.dout(n4192),.clk(gclk));
	jor g3551(.dina(n4192),.dinb(n4191),.dout(n4193),.clk(gclk));
	jand g3552(.dina(w_n4193_0[1]),.dinb(w_n4190_0[1]),.dout(n4194),.clk(gclk));
	jor g3553(.dina(n4194),.dinb(n4186),.dout(n4195),.clk(gclk));
	jnot g3554(.din(n4195),.dout(n4196),.clk(gclk));
	jand g3555(.dina(w_n1721_25[0]),.dinb(w_n834_0[0]),.dout(n4197),.clk(gclk));
	jand g3556(.dina(w_n1562_25[0]),.dinb(w_n1353_0[0]),.dout(n4198),.clk(gclk));
	jor g3557(.dina(n4198),.dinb(n4197),.dout(n4199),.clk(gclk));
	jand g3558(.dina(w_n2803_24[2]),.dinb(w_n2440_0[0]),.dout(n4200),.clk(gclk));
	jand g3559(.dina(w_n2808_25[0]),.dinb(w_n2446_0[0]),.dout(n4201),.clk(gclk));
	jor g3560(.dina(n4201),.dinb(n4200),.dout(n4202),.clk(gclk));
	jnot g3561(.din(w_n4202_0[1]),.dout(n4203),.clk(gclk));
	jand g3562(.dina(w_n4203_0[1]),.dinb(w_n4199_0[1]),.dout(n4204),.clk(gclk));
	jnot g3563(.din(n4204),.dout(n4205),.clk(gclk));
	jand g3564(.dina(w_n4205_0[1]),.dinb(w_n4196_0[1]),.dout(n4206),.clk(gclk));
	jand g3565(.dina(n4206),.dinb(n4178),.dout(n4207),.clk(gclk));
	jnot g3566(.din(w_n4207_0[1]),.dout(n4208),.clk(gclk));
	jor g3567(.dina(n4208),.dinb(n4169),.dout(n4209),.clk(gclk));
	jnot g3568(.din(w_n4181_0[0]),.dout(n4210),.clk(gclk));
	jand g3569(.dina(w_n4184_0[0]),.dinb(w_n4210_0[1]),.dout(n4211),.clk(gclk));
	jnot g3570(.din(w_n4193_0[0]),.dout(n4212),.clk(gclk));
	jand g3571(.dina(w_n4212_0[1]),.dinb(w_n4189_0[0]),.dout(n4213),.clk(gclk));
	jnot g3572(.din(w_n4176_0[0]),.dout(n4214),.clk(gclk));
	jand g3573(.dina(w_n4214_0[1]),.dinb(w_n4172_0[0]),.dout(n4215),.clk(gclk));
	jand g3574(.dina(n4215),.dinb(w_n4205_0[0]),.dout(n4216),.clk(gclk));
	jnot g3575(.din(w_n4199_0[0]),.dout(n4217),.clk(gclk));
	jand g3576(.dina(w_n4202_0[0]),.dinb(w_n4217_0[1]),.dout(n4218),.clk(gclk));
	jor g3577(.dina(n4218),.dinb(n4216),.dout(n4219),.clk(gclk));
	jor g3578(.dina(n4219),.dinb(n4213),.dout(n4220),.clk(gclk));
	jand g3579(.dina(n4220),.dinb(w_n4196_0[0]),.dout(n4221),.clk(gclk));
	jor g3580(.dina(n4221),.dinb(n4211),.dout(n4222),.clk(gclk));
	jnot g3581(.din(w_n4222_0[1]),.dout(n4223),.clk(gclk));
	jand g3582(.dina(n4223),.dinb(n4209),.dout(n4224),.clk(gclk));
	jor g3583(.dina(n4224),.dinb(w_n3237_0[1]),.dout(n4225),.clk(gclk));
	jnot g3584(.din(w_n3236_0[0]),.dout(n4226),.clk(gclk));
	jnot g3585(.din(w_n3229_0[0]),.dout(n4227),.clk(gclk));
	jand g3586(.dina(w_n3232_0[0]),.dinb(w_n4227_0[1]),.dout(n4228),.clk(gclk));
	jnot g3587(.din(w_n3205_0[0]),.dout(n4229),.clk(gclk));
	jand g3588(.dina(w_n3208_0[0]),.dinb(w_n4229_0[1]),.dout(n4230),.clk(gclk));
	jor g3589(.dina(n4230),.dinb(n4228),.dout(n4231),.clk(gclk));
	jand g3590(.dina(n4231),.dinb(n4226),.dout(n4232),.clk(gclk));
	jnot g3591(.din(w_n3226_0[0]),.dout(n4233),.clk(gclk));
	jnot g3592(.din(w_n3221_0[0]),.dout(n4234),.clk(gclk));
	jand g3593(.dina(w_n3224_0[0]),.dinb(w_n4234_0[1]),.dout(n4235),.clk(gclk));
	jnot g3594(.din(w_n3217_0[0]),.dout(n4236),.clk(gclk));
	jand g3595(.dina(w_n4236_0[1]),.dinb(w_n3213_0[0]),.dout(n4237),.clk(gclk));
	jor g3596(.dina(n4237),.dinb(n4235),.dout(n4238),.clk(gclk));
	jand g3597(.dina(n4238),.dinb(n4233),.dout(n4239),.clk(gclk));
	jor g3598(.dina(n4239),.dinb(n4232),.dout(n4240),.clk(gclk));
	jnot g3599(.din(w_n4240_0[1]),.dout(n4241),.clk(gclk));
	jand g3600(.dina(n4241),.dinb(n4225),.dout(n4242),.clk(gclk));
	jor g3601(.dina(n4242),.dinb(w_n3202_0[1]),.dout(n4243),.clk(gclk));
	jnot g3602(.din(w_n3184_0[0]),.dout(n4244),.clk(gclk));
	jnot g3603(.din(w_n3182_0[0]),.dout(n4245),.clk(gclk));
	jand g3604(.dina(w_n4245_0[1]),.dinb(w_n3178_0[0]),.dout(n4246),.clk(gclk));
	jnot g3605(.din(w_n3192_0[0]),.dout(n4247),.clk(gclk));
	jnot g3606(.din(w_n3199_0[0]),.dout(n4248),.clk(gclk));
	jand g3607(.dina(w_n4248_0[1]),.dinb(w_n3195_0[0]),.dout(n4249),.clk(gclk));
	jand g3608(.dina(n4249),.dinb(n4247),.dout(n4250),.clk(gclk));
	jnot g3609(.din(w_n3187_0[0]),.dout(n4251),.clk(gclk));
	jand g3610(.dina(w_n3190_0[0]),.dinb(w_n4251_0[1]),.dout(n4252),.clk(gclk));
	jor g3611(.dina(n4252),.dinb(n4250),.dout(n4253),.clk(gclk));
	jor g3612(.dina(n4253),.dinb(n4246),.dout(n4254),.clk(gclk));
	jand g3613(.dina(n4254),.dinb(n4244),.dout(n4255),.clk(gclk));
	jnot g3614(.din(w_n4255_0[1]),.dout(n4256),.clk(gclk));
	jand g3615(.dina(n4256),.dinb(n4243),.dout(n4257),.clk(gclk));
	jand g3616(.dina(n4257),.dinb(n3173),.dout(n4258),.clk(gclk));
	jnot g3617(.din(w_n3152_0[0]),.dout(n4259),.clk(gclk));
	jand g3618(.dina(w_n4259_0[1]),.dinb(w_n3148_0[0]),.dout(n4260),.clk(gclk));
	jor g3619(.dina(n4260),.dinb(w_n3142_0[0]),.dout(n4261),.clk(gclk));
	jor g3620(.dina(w_n4261_0[1]),.dinb(n4258),.dout(n4262),.clk(gclk));
	jand g3621(.dina(n4262),.dinb(n3164),.dout(n4263),.clk(gclk));
	jand g3622(.dina(n4263),.dinb(n3156),.dout(n4264),.clk(gclk));
	jor g3623(.dina(n4264),.dinb(w_n3116_0[1]),.dout(n4265),.clk(gclk));
	jnot g3624(.din(w_n3084_0[0]),.dout(n4266),.clk(gclk));
	jand g3625(.dina(w_n3087_0[0]),.dinb(w_n4266_0[1]),.dout(n4267),.clk(gclk));
	jnot g3626(.din(w_n3098_0[0]),.dout(n4268),.clk(gclk));
	jnot g3627(.din(w_n3096_0[0]),.dout(n4269),.clk(gclk));
	jand g3628(.dina(w_n4269_0[1]),.dinb(w_n3092_0[0]),.dout(n4270),.clk(gclk));
	jnot g3629(.din(w_n3106_0[0]),.dout(n4271),.clk(gclk));
	jnot g3630(.din(w_n3113_0[0]),.dout(n4272),.clk(gclk));
	jand g3631(.dina(w_n4272_0[1]),.dinb(w_n3109_0[0]),.dout(n4273),.clk(gclk));
	jand g3632(.dina(n4273),.dinb(n4271),.dout(n4274),.clk(gclk));
	jnot g3633(.din(w_n3101_0[0]),.dout(n4275),.clk(gclk));
	jand g3634(.dina(w_n3104_0[0]),.dinb(w_n4275_0[1]),.dout(n4276),.clk(gclk));
	jor g3635(.dina(n4276),.dinb(n4274),.dout(n4277),.clk(gclk));
	jor g3636(.dina(n4277),.dinb(n4270),.dout(n4278),.clk(gclk));
	jand g3637(.dina(n4278),.dinb(n4268),.dout(n4279),.clk(gclk));
	jor g3638(.dina(n4279),.dinb(n4267),.dout(n4280),.clk(gclk));
	jnot g3639(.din(w_n4280_0[1]),.dout(n4281),.clk(gclk));
	jand g3640(.dina(n4281),.dinb(n4265),.dout(n4282),.clk(gclk));
	jor g3641(.dina(n4282),.dinb(w_n3081_0[1]),.dout(n4283),.clk(gclk));
	jnot g3642(.din(w_n3080_0[0]),.dout(n4284),.clk(gclk));
	jnot g3643(.din(w_n3073_0[0]),.dout(n4285),.clk(gclk));
	jand g3644(.dina(w_n3076_0[0]),.dinb(w_n4285_0[1]),.dout(n4286),.clk(gclk));
	jnot g3645(.din(w_n3049_0[0]),.dout(n4287),.clk(gclk));
	jand g3646(.dina(w_n3052_0[0]),.dinb(w_n4287_0[1]),.dout(n4288),.clk(gclk));
	jor g3647(.dina(n4288),.dinb(n4286),.dout(n4289),.clk(gclk));
	jand g3648(.dina(n4289),.dinb(n4284),.dout(n4290),.clk(gclk));
	jnot g3649(.din(w_n3070_0[0]),.dout(n4291),.clk(gclk));
	jnot g3650(.din(w_n3065_0[0]),.dout(n4292),.clk(gclk));
	jand g3651(.dina(w_n3068_0[0]),.dinb(w_n4292_0[1]),.dout(n4293),.clk(gclk));
	jnot g3652(.din(w_n3061_0[0]),.dout(n4294),.clk(gclk));
	jand g3653(.dina(w_n4294_0[1]),.dinb(w_n3057_0[0]),.dout(n4295),.clk(gclk));
	jor g3654(.dina(n4295),.dinb(n4293),.dout(n4296),.clk(gclk));
	jand g3655(.dina(n4296),.dinb(n4291),.dout(n4297),.clk(gclk));
	jor g3656(.dina(n4297),.dinb(n4290),.dout(n4298),.clk(gclk));
	jnot g3657(.din(w_n4298_0[1]),.dout(n4299),.clk(gclk));
	jand g3658(.dina(n4299),.dinb(n4283),.dout(n4300),.clk(gclk));
	jor g3659(.dina(n4300),.dinb(w_n3046_0[1]),.dout(n4301),.clk(gclk));
	jnot g3660(.din(w_n3014_0[0]),.dout(n4302),.clk(gclk));
	jand g3661(.dina(w_n3017_0[0]),.dinb(w_n4302_0[1]),.dout(n4303),.clk(gclk));
	jnot g3662(.din(w_n3028_0[0]),.dout(n4304),.clk(gclk));
	jnot g3663(.din(w_n3026_0[0]),.dout(n4305),.clk(gclk));
	jand g3664(.dina(w_n4305_0[1]),.dinb(w_n3022_0[0]),.dout(n4306),.clk(gclk));
	jnot g3665(.din(w_n3036_0[0]),.dout(n4307),.clk(gclk));
	jnot g3666(.din(w_n3043_0[0]),.dout(n4308),.clk(gclk));
	jand g3667(.dina(w_n4308_0[1]),.dinb(w_n3039_0[0]),.dout(n4309),.clk(gclk));
	jand g3668(.dina(n4309),.dinb(n4307),.dout(n4310),.clk(gclk));
	jnot g3669(.din(w_n3031_0[0]),.dout(n4311),.clk(gclk));
	jand g3670(.dina(w_n3034_0[0]),.dinb(w_n4311_0[1]),.dout(n4312),.clk(gclk));
	jor g3671(.dina(n4312),.dinb(n4310),.dout(n4313),.clk(gclk));
	jor g3672(.dina(n4313),.dinb(n4306),.dout(n4314),.clk(gclk));
	jand g3673(.dina(n4314),.dinb(n4304),.dout(n4315),.clk(gclk));
	jor g3674(.dina(n4315),.dinb(n4303),.dout(n4316),.clk(gclk));
	jnot g3675(.din(w_n4316_0[1]),.dout(n4317),.clk(gclk));
	jand g3676(.dina(n4317),.dinb(n4301),.dout(n4318),.clk(gclk));
	jor g3677(.dina(n4318),.dinb(w_n3011_0[1]),.dout(n4319),.clk(gclk));
	jnot g3678(.din(w_n3010_0[0]),.dout(n4320),.clk(gclk));
	jnot g3679(.din(w_n3003_0[0]),.dout(n4321),.clk(gclk));
	jand g3680(.dina(w_n3006_0[0]),.dinb(w_n4321_0[1]),.dout(n4322),.clk(gclk));
	jnot g3681(.din(w_n2979_0[0]),.dout(n4323),.clk(gclk));
	jand g3682(.dina(w_n2982_0[0]),.dinb(w_n4323_0[1]),.dout(n4324),.clk(gclk));
	jor g3683(.dina(n4324),.dinb(n4322),.dout(n4325),.clk(gclk));
	jand g3684(.dina(n4325),.dinb(n4320),.dout(n4326),.clk(gclk));
	jnot g3685(.din(w_n3000_0[0]),.dout(n4327),.clk(gclk));
	jnot g3686(.din(w_n2995_0[0]),.dout(n4328),.clk(gclk));
	jand g3687(.dina(w_n2998_0[0]),.dinb(w_n4328_0[1]),.dout(n4329),.clk(gclk));
	jnot g3688(.din(w_n2991_0[0]),.dout(n4330),.clk(gclk));
	jand g3689(.dina(w_n4330_0[1]),.dinb(w_n2987_0[0]),.dout(n4331),.clk(gclk));
	jor g3690(.dina(n4331),.dinb(n4329),.dout(n4332),.clk(gclk));
	jand g3691(.dina(n4332),.dinb(n4327),.dout(n4333),.clk(gclk));
	jor g3692(.dina(n4333),.dinb(n4326),.dout(n4334),.clk(gclk));
	jnot g3693(.din(w_n4334_0[1]),.dout(n4335),.clk(gclk));
	jand g3694(.dina(n4335),.dinb(n4319),.dout(n4336),.clk(gclk));
	jor g3695(.dina(n4336),.dinb(w_n2976_0[1]),.dout(n4337),.clk(gclk));
	jnot g3696(.din(w_n2944_0[0]),.dout(n4338),.clk(gclk));
	jand g3697(.dina(w_n2947_0[0]),.dinb(w_n4338_0[1]),.dout(n4339),.clk(gclk));
	jnot g3698(.din(w_n2958_0[0]),.dout(n4340),.clk(gclk));
	jnot g3699(.din(w_n2956_0[0]),.dout(n4341),.clk(gclk));
	jand g3700(.dina(w_n4341_0[1]),.dinb(w_n2952_0[0]),.dout(n4342),.clk(gclk));
	jnot g3701(.din(w_n2966_0[0]),.dout(n4343),.clk(gclk));
	jnot g3702(.din(w_n2973_0[0]),.dout(n4344),.clk(gclk));
	jand g3703(.dina(w_n4344_0[1]),.dinb(w_n2969_0[0]),.dout(n4345),.clk(gclk));
	jand g3704(.dina(n4345),.dinb(n4343),.dout(n4346),.clk(gclk));
	jnot g3705(.din(w_n2961_0[0]),.dout(n4347),.clk(gclk));
	jand g3706(.dina(w_n2964_0[0]),.dinb(w_n4347_0[1]),.dout(n4348),.clk(gclk));
	jor g3707(.dina(n4348),.dinb(n4346),.dout(n4349),.clk(gclk));
	jor g3708(.dina(n4349),.dinb(n4342),.dout(n4350),.clk(gclk));
	jand g3709(.dina(n4350),.dinb(n4340),.dout(n4351),.clk(gclk));
	jor g3710(.dina(n4351),.dinb(n4339),.dout(n4352),.clk(gclk));
	jnot g3711(.din(w_n4352_0[1]),.dout(n4353),.clk(gclk));
	jand g3712(.dina(n4353),.dinb(n4337),.dout(n4354),.clk(gclk));
	jor g3713(.dina(n4354),.dinb(w_n2941_0[1]),.dout(n4355),.clk(gclk));
	jnot g3714(.din(w_n2914_0[0]),.dout(n4356),.clk(gclk));
	jnot g3715(.din(w_n2909_0[0]),.dout(n4357),.clk(gclk));
	jand g3716(.dina(w_n2912_0[0]),.dinb(w_n4357_0[1]),.dout(n4358),.clk(gclk));
	jnot g3717(.din(w_n2905_0[0]),.dout(n4359),.clk(gclk));
	jand g3718(.dina(w_n4359_0[1]),.dinb(w_n2901_0[0]),.dout(n4360),.clk(gclk));
	jor g3719(.dina(n4360),.dinb(n4358),.dout(n4361),.clk(gclk));
	jand g3720(.dina(n4361),.dinb(n4356),.dout(n4362),.clk(gclk));
	jnot g3721(.din(w_n4362_0[1]),.dout(n4363),.clk(gclk));
	jand g3722(.dina(n4363),.dinb(n4355),.dout(n4364),.clk(gclk));
	jand g3723(.dina(n4364),.dinb(n2938),.dout(n4365),.clk(gclk));
	jand g3724(.dina(w_n1721_24[2]),.dinb(w_n677_0[0]),.dout(n4366),.clk(gclk));
	jand g3725(.dina(w_n1562_24[2]),.dinb(w_n1493_0[0]),.dout(n4367),.clk(gclk));
	jor g3726(.dina(n4367),.dinb(n4366),.dout(n4368),.clk(gclk));
	jand g3727(.dina(w_n2803_24[1]),.dinb(w_n1770_0[0]),.dout(n4369),.clk(gclk));
	jand g3728(.dina(w_n2808_24[2]),.dinb(w_n2591_0[0]),.dout(n4370),.clk(gclk));
	jor g3729(.dina(n4370),.dinb(n4369),.dout(n4371),.clk(gclk));
	jnot g3730(.din(w_n4371_0[1]),.dout(n4372),.clk(gclk));
	jand g3731(.dina(w_n4372_0[1]),.dinb(w_n4368_0[1]),.dout(n4373),.clk(gclk));
	jnot g3732(.din(w_n2896_0[0]),.dout(n4374),.clk(gclk));
	jand g3733(.dina(w_n4374_0[1]),.dinb(w_n2892_0[0]),.dout(n4375),.clk(gclk));
	jand g3734(.dina(w_n2803_24[0]),.dinb(w_n2585_0[0]),.dout(n4376),.clk(gclk));
	jand g3735(.dina(w_n2808_24[1]),.dinb(w_n2593_0[0]),.dout(n4377),.clk(gclk));
	jor g3736(.dina(n4377),.dinb(n4376),.dout(n4378),.clk(gclk));
	jnot g3737(.din(w_n4378_0[1]),.dout(n4379),.clk(gclk));
	jand g3738(.dina(w_n1721_24[1]),.dinb(w_n1487_0[0]),.dout(n4380),.clk(gclk));
	jand g3739(.dina(w_n1562_24[1]),.dinb(w_n1495_0[0]),.dout(n4381),.clk(gclk));
	jor g3740(.dina(n4381),.dinb(n4380),.dout(n4382),.clk(gclk));
	jand g3741(.dina(w_n4382_0[1]),.dinb(w_n4379_0[1]),.dout(n4383),.clk(gclk));
	jor g3742(.dina(n4383),.dinb(n4375),.dout(n4384),.clk(gclk));
	jand g3743(.dina(w_n2803_23[2]),.dinb(w_n1772_0[0]),.dout(n4385),.clk(gclk));
	jand g3744(.dina(w_n2808_24[0]),.dinb(w_n2597_0[0]),.dout(n4386),.clk(gclk));
	jor g3745(.dina(n4386),.dinb(n4385),.dout(n4387),.clk(gclk));
	jnot g3746(.din(w_n4387_0[1]),.dout(n4388),.clk(gclk));
	jand g3747(.dina(w_n1721_24[0]),.dinb(w_n679_0[0]),.dout(n4389),.clk(gclk));
	jand g3748(.dina(w_n1562_24[0]),.dinb(w_n1499_0[0]),.dout(n4390),.clk(gclk));
	jor g3749(.dina(n4390),.dinb(n4389),.dout(n4391),.clk(gclk));
	jand g3750(.dina(w_n4391_0[1]),.dinb(w_n4388_0[1]),.dout(n4392),.clk(gclk));
	jor g3751(.dina(n4392),.dinb(w_n4384_0[1]),.dout(n4393),.clk(gclk));
	jor g3752(.dina(n4393),.dinb(w_n4373_0[1]),.dout(n4394),.clk(gclk));
	jor g3753(.dina(w_n4394_0[1]),.dinb(n4365),.dout(n4395),.clk(gclk));
	jnot g3754(.din(w_n4384_0[0]),.dout(n4396),.clk(gclk));
	jnot g3755(.din(w_n4382_0[0]),.dout(n4397),.clk(gclk));
	jand g3756(.dina(w_n4397_0[1]),.dinb(w_n4378_0[0]),.dout(n4398),.clk(gclk));
	jnot g3757(.din(w_n4373_0[0]),.dout(n4399),.clk(gclk));
	jnot g3758(.din(w_n4391_0[0]),.dout(n4400),.clk(gclk));
	jand g3759(.dina(w_n4400_0[1]),.dinb(w_n4387_0[0]),.dout(n4401),.clk(gclk));
	jand g3760(.dina(n4401),.dinb(n4399),.dout(n4402),.clk(gclk));
	jnot g3761(.din(w_n4368_0[0]),.dout(n4403),.clk(gclk));
	jand g3762(.dina(w_n4371_0[0]),.dinb(w_n4403_0[1]),.dout(n4404),.clk(gclk));
	jor g3763(.dina(n4404),.dinb(n4402),.dout(n4405),.clk(gclk));
	jor g3764(.dina(n4405),.dinb(n4398),.dout(n4406),.clk(gclk));
	jand g3765(.dina(n4406),.dinb(n4396),.dout(n4407),.clk(gclk));
	jnot g3766(.din(w_n4407_0[1]),.dout(n4408),.clk(gclk));
	jand g3767(.dina(n4408),.dinb(n4395),.dout(n4409),.clk(gclk));
	jand g3768(.dina(n4409),.dinb(n2898),.dout(n4410),.clk(gclk));
	jnot g3769(.din(w_n2877_0[0]),.dout(n4411),.clk(gclk));
	jand g3770(.dina(w_n4411_0[1]),.dinb(w_n2873_0[0]),.dout(n4412),.clk(gclk));
	jor g3771(.dina(n4412),.dinb(w_n2867_0[0]),.dout(n4413),.clk(gclk));
	jor g3772(.dina(w_n4413_0[1]),.dinb(n4410),.dout(n4414),.clk(gclk));
	jand g3773(.dina(n4414),.dinb(n2889),.dout(n4415),.clk(gclk));
	jand g3774(.dina(w_n2803_23[1]),.dinb(w_n2615_0[0]),.dout(n4416),.clk(gclk));
	jand g3775(.dina(w_n2808_23[2]),.dinb(w_n2629_0[0]),.dout(n4417),.clk(gclk));
	jor g3776(.dina(n4417),.dinb(n4416),.dout(n4418),.clk(gclk));
	jnot g3777(.din(w_n4418_0[1]),.dout(n4419),.clk(gclk));
	jand g3778(.dina(w_n1721_23[2]),.dinb(w_n645_0[0]),.dout(n4420),.clk(gclk));
	jand g3779(.dina(w_n1562_23[2]),.dinb(w_n1526_0[0]),.dout(n4421),.clk(gclk));
	jor g3780(.dina(n4421),.dinb(n4420),.dout(n4422),.clk(gclk));
	jand g3781(.dina(w_n4422_0[1]),.dinb(w_n4419_0[1]),.dout(n4423),.clk(gclk));
	jnot g3782(.din(n4423),.dout(n4424),.clk(gclk));
	jand g3783(.dina(w_n1721_23[1]),.dinb(w_n1512_0[0]),.dout(n4425),.clk(gclk));
	jand g3784(.dina(w_n1562_23[1]),.dinb(w_n642_0[0]),.dout(n4426),.clk(gclk));
	jor g3785(.dina(n4426),.dinb(n4425),.dout(n4427),.clk(gclk));
	jand g3786(.dina(w_n2803_23[0]),.dinb(w_n2610_0[0]),.dout(n4428),.clk(gclk));
	jand g3787(.dina(w_n2808_23[1]),.dinb(w_n1740_0[0]),.dout(n4429),.clk(gclk));
	jor g3788(.dina(n4429),.dinb(n4428),.dout(n4430),.clk(gclk));
	jnot g3789(.din(w_n4430_0[1]),.dout(n4431),.clk(gclk));
	jand g3790(.dina(w_n4431_0[1]),.dinb(w_n4427_0[1]),.dout(n4432),.clk(gclk));
	jand g3791(.dina(w_n2803_22[2]),.dinb(w_n2612_0[0]),.dout(n4433),.clk(gclk));
	jand g3792(.dina(w_n2808_23[0]),.dinb(w_n2625_0[0]),.dout(n4434),.clk(gclk));
	jor g3793(.dina(n4434),.dinb(n4433),.dout(n4435),.clk(gclk));
	jnot g3794(.din(w_n4435_0[1]),.dout(n4436),.clk(gclk));
	jand g3795(.dina(w_n1721_23[0]),.dinb(w_n1514_0[0]),.dout(n4437),.clk(gclk));
	jand g3796(.dina(w_n1562_23[0]),.dinb(w_n1522_0[0]),.dout(n4438),.clk(gclk));
	jor g3797(.dina(n4438),.dinb(n4437),.dout(n4439),.clk(gclk));
	jand g3798(.dina(w_n4439_0[1]),.dinb(w_n4436_0[1]),.dout(n4440),.clk(gclk));
	jor g3799(.dina(n4440),.dinb(n4432),.dout(n4441),.clk(gclk));
	jnot g3800(.din(n4441),.dout(n4442),.clk(gclk));
	jand g3801(.dina(w_n1721_22[2]),.dinb(w_n647_0[0]),.dout(n4443),.clk(gclk));
	jand g3802(.dina(w_n1562_22[2]),.dinb(w_n1520_0[0]),.dout(n4444),.clk(gclk));
	jor g3803(.dina(n4444),.dinb(n4443),.dout(n4445),.clk(gclk));
	jand g3804(.dina(w_n2803_22[1]),.dinb(w_n2617_0[0]),.dout(n4446),.clk(gclk));
	jand g3805(.dina(w_n2808_22[2]),.dinb(w_n2623_0[0]),.dout(n4447),.clk(gclk));
	jor g3806(.dina(n4447),.dinb(n4446),.dout(n4448),.clk(gclk));
	jnot g3807(.din(w_n4448_0[1]),.dout(n4449),.clk(gclk));
	jand g3808(.dina(w_n4449_0[1]),.dinb(w_n4445_0[1]),.dout(n4450),.clk(gclk));
	jnot g3809(.din(n4450),.dout(n4451),.clk(gclk));
	jand g3810(.dina(w_n4451_0[1]),.dinb(w_n4442_0[1]),.dout(n4452),.clk(gclk));
	jand g3811(.dina(n4452),.dinb(n4424),.dout(n4453),.clk(gclk));
	jnot g3812(.din(w_n4453_0[1]),.dout(n4454),.clk(gclk));
	jor g3813(.dina(n4454),.dinb(n4415),.dout(n4455),.clk(gclk));
	jnot g3814(.din(w_n4427_0[0]),.dout(n4456),.clk(gclk));
	jand g3815(.dina(w_n4430_0[0]),.dinb(w_n4456_0[1]),.dout(n4457),.clk(gclk));
	jnot g3816(.din(w_n4439_0[0]),.dout(n4458),.clk(gclk));
	jand g3817(.dina(w_n4458_0[1]),.dinb(w_n4435_0[0]),.dout(n4459),.clk(gclk));
	jnot g3818(.din(w_n4422_0[0]),.dout(n4460),.clk(gclk));
	jand g3819(.dina(w_n4460_0[1]),.dinb(w_n4418_0[0]),.dout(n4461),.clk(gclk));
	jand g3820(.dina(n4461),.dinb(w_n4451_0[0]),.dout(n4462),.clk(gclk));
	jnot g3821(.din(w_n4445_0[0]),.dout(n4463),.clk(gclk));
	jand g3822(.dina(w_n4448_0[0]),.dinb(w_n4463_0[1]),.dout(n4464),.clk(gclk));
	jor g3823(.dina(n4464),.dinb(n4462),.dout(n4465),.clk(gclk));
	jor g3824(.dina(n4465),.dinb(n4459),.dout(n4466),.clk(gclk));
	jand g3825(.dina(n4466),.dinb(w_n4442_0[0]),.dout(n4467),.clk(gclk));
	jor g3826(.dina(n4467),.dinb(n4457),.dout(n4468),.clk(gclk));
	jnot g3827(.din(w_n4468_0[1]),.dout(n4469),.clk(gclk));
	jand g3828(.dina(n4469),.dinb(n4455),.dout(n4470),.clk(gclk));
	jor g3829(.dina(n4470),.dinb(w_n2841_0[1]),.dout(n4471),.clk(gclk));
	jand g3830(.dina(n4471),.dinb(n2838),.dout(n4472),.clk(gclk));
	jor g3831(.dina(n4472),.dinb(w_n2644_0[1]),.dout(n4473),.clk(gclk));
	jand g3832(.dina(w_n4473_0[1]),.dinb(w_n2642_0[0]),.dout(n4474),.clk(gclk));
	jand g3833(.dina(w_n4473_0[0]),.dinb(w_n2643_1[0]),.dout(n4475),.clk(gclk));
	jor g3834(.dina(n4475),.dinb(n4474),.dout(address1_fa_),.clk(gclk));
	jor g3835(.dina(w_address1_63[1]),.dinb(w_n1723_0[1]),.dout(n4477),.clk(gclk));
	jnot g3836(.din(w_n2644_0[0]),.dout(n4478),.clk(gclk));
	jnot g3837(.din(w_n2841_0[0]),.dout(n4479),.clk(gclk));
	jnot g3838(.din(w_n2941_0[0]),.dout(n4480),.clk(gclk));
	jnot g3839(.din(w_n2976_0[0]),.dout(n4481),.clk(gclk));
	jnot g3840(.din(w_n3011_0[0]),.dout(n4482),.clk(gclk));
	jnot g3841(.din(w_n3046_0[0]),.dout(n4483),.clk(gclk));
	jnot g3842(.din(w_n3081_0[0]),.dout(n4484),.clk(gclk));
	jnot g3843(.din(w_n3116_0[0]),.dout(n4485),.clk(gclk));
	jnot g3844(.din(w_n3202_0[0]),.dout(n4486),.clk(gclk));
	jnot g3845(.din(w_n3237_0[0]),.dout(n4487),.clk(gclk));
	jnot g3846(.din(w_n3581_0[0]),.dout(n4488),.clk(gclk));
	jnot g3847(.din(w_n3598_0[0]),.dout(n4489),.clk(gclk));
	jnot g3848(.din(w_n3633_0[0]),.dout(n4490),.clk(gclk));
	jnot g3849(.din(w_n3641_0[0]),.dout(n4491),.clk(gclk));
	jnot g3850(.din(w_n3652_0[0]),.dout(n4492),.clk(gclk));
	jnot g3851(.din(w_n3660_0[0]),.dout(n4493),.clk(gclk));
	jnot g3852(.din(w_n3677_0[0]),.dout(n4494),.clk(gclk));
	jnot g3853(.din(w_n3685_0[0]),.dout(n4495),.clk(gclk));
	jnot g3854(.din(w_n3696_0[0]),.dout(n4496),.clk(gclk));
	jnot g3855(.din(w_n3713_0[0]),.dout(n4497),.clk(gclk));
	jnot g3856(.din(w_n3730_0[0]),.dout(n4498),.clk(gclk));
	jnot g3857(.din(w_n3738_0[0]),.dout(n4499),.clk(gclk));
	jnot g3858(.din(w_n3749_0[0]),.dout(n4500),.clk(gclk));
	jand g3859(.dina(w_n2803_22[0]),.dinb(w_n2113_0[0]),.dout(n4501),.clk(gclk));
	jand g3860(.dina(w_n2808_22[1]),.dinb(w_n2110_0[0]),.dout(n4502),.clk(gclk));
	jor g3861(.dina(n4502),.dinb(n4501),.dout(n4503),.clk(gclk));
	jor g3862(.dina(w_n1562_22[1]),.dinb(w_in01_0[1]),.dout(n4504),.clk(gclk));
	jor g3863(.dina(w_n1721_22[1]),.dinb(w_in11_0[1]),.dout(n4505),.clk(gclk));
	jand g3864(.dina(n4505),.dinb(n4504),.dout(n4506),.clk(gclk));
	jand g3865(.dina(w_n4506_0[2]),.dinb(w_n4503_0[1]),.dout(n4507),.clk(gclk));
	jand g3866(.dina(w_n2803_21[2]),.dinb(w_n2115_0[0]),.dout(n4508),.clk(gclk));
	jand g3867(.dina(w_n2808_22[0]),.dinb(w_n2672_0[0]),.dout(n4509),.clk(gclk));
	jor g3868(.dina(n4509),.dinb(n4508),.dout(n4510),.clk(gclk));
	jand g3869(.dina(n4510),.dinb(w_n1723_0[0]),.dout(n4511),.clk(gclk));
	jor g3870(.dina(n4511),.dinb(n4507),.dout(n4512),.clk(gclk));
	jor g3871(.dina(w_n1562_22[0]),.dinb(w_in02_0[1]),.dout(n4513),.clk(gclk));
	jor g3872(.dina(w_n1721_22[0]),.dinb(w_in12_0[0]),.dout(n4514),.clk(gclk));
	jand g3873(.dina(n4514),.dinb(n4513),.dout(n4515),.clk(gclk));
	jand g3874(.dina(w_n2803_21[1]),.dinb(w_n2108_0[0]),.dout(n4516),.clk(gclk));
	jand g3875(.dina(w_n2808_21[2]),.dinb(w_n2122_0[0]),.dout(n4517),.clk(gclk));
	jor g3876(.dina(n4517),.dinb(n4516),.dout(n4518),.clk(gclk));
	jor g3877(.dina(w_n4518_0[1]),.dinb(w_n4515_0[2]),.dout(n4519),.clk(gclk));
	jor g3878(.dina(w_n4506_0[1]),.dinb(w_n4503_0[0]),.dout(n4520),.clk(gclk));
	jand g3879(.dina(n4520),.dinb(n4519),.dout(n4521),.clk(gclk));
	jand g3880(.dina(n4521),.dinb(n4512),.dout(n4522),.clk(gclk));
	jand g3881(.dina(w_n4518_0[0]),.dinb(w_n4515_0[1]),.dout(n4523),.clk(gclk));
	jor g3882(.dina(w_n1562_21[2]),.dinb(w_in03_0[0]),.dout(n4524),.clk(gclk));
	jor g3883(.dina(w_n1721_21[2]),.dinb(w_in13_0[0]),.dout(n4525),.clk(gclk));
	jand g3884(.dina(n4525),.dinb(n4524),.dout(n4526),.clk(gclk));
	jand g3885(.dina(w_n3790_0[0]),.dinb(w_n4526_0[1]),.dout(n4527),.clk(gclk));
	jor g3886(.dina(n4527),.dinb(n4523),.dout(n4528),.clk(gclk));
	jor g3887(.dina(n4528),.dinb(n4522),.dout(n4529),.clk(gclk));
	jnot g3888(.din(w_n3798_0[0]),.dout(n4530),.clk(gclk));
	jand g3889(.dina(n4530),.dinb(n4529),.dout(n4531),.clk(gclk));
	jor g3890(.dina(n4531),.dinb(w_n3757_0[0]),.dout(n4532),.clk(gclk));
	jand g3891(.dina(n4532),.dinb(n4500),.dout(n4533),.clk(gclk));
	jor g3892(.dina(n4533),.dinb(w_n3746_0[0]),.dout(n4534),.clk(gclk));
	jand g3893(.dina(n4534),.dinb(n4499),.dout(n4535),.clk(gclk));
	jor g3894(.dina(w_n3808_0[0]),.dinb(n4535),.dout(n4536),.clk(gclk));
	jnot g3895(.din(w_n3812_0[0]),.dout(n4537),.clk(gclk));
	jand g3896(.dina(n4537),.dinb(n4536),.dout(n4538),.clk(gclk));
	jand g3897(.dina(n4538),.dinb(n4498),.dout(n4539),.clk(gclk));
	jor g3898(.dina(w_n3822_0[0]),.dinb(n4539),.dout(n4540),.clk(gclk));
	jor g3899(.dina(n4540),.dinb(w_n3721_0[0]),.dout(n4541),.clk(gclk));
	jnot g3900(.din(w_n3827_0[0]),.dout(n4542),.clk(gclk));
	jand g3901(.dina(n4542),.dinb(n4541),.dout(n4543),.clk(gclk));
	jand g3902(.dina(n4543),.dinb(n4497),.dout(n4544),.clk(gclk));
	jor g3903(.dina(w_n3840_0[0]),.dinb(n4544),.dout(n4545),.clk(gclk));
	jnot g3904(.din(w_n3847_0[0]),.dout(n4546),.clk(gclk));
	jand g3905(.dina(n4546),.dinb(n4545),.dout(n4547),.clk(gclk));
	jor g3906(.dina(n4547),.dinb(w_n3704_0[0]),.dout(n4548),.clk(gclk));
	jand g3907(.dina(n4548),.dinb(n4496),.dout(n4549),.clk(gclk));
	jor g3908(.dina(n4549),.dinb(w_n3693_0[0]),.dout(n4550),.clk(gclk));
	jand g3909(.dina(n4550),.dinb(n4495),.dout(n4551),.clk(gclk));
	jor g3910(.dina(w_n3857_0[0]),.dinb(n4551),.dout(n4552),.clk(gclk));
	jnot g3911(.din(w_n3861_0[0]),.dout(n4553),.clk(gclk));
	jand g3912(.dina(n4553),.dinb(n4552),.dout(n4554),.clk(gclk));
	jand g3913(.dina(n4554),.dinb(n4494),.dout(n4555),.clk(gclk));
	jor g3914(.dina(w_n3871_0[0]),.dinb(n4555),.dout(n4556),.clk(gclk));
	jor g3915(.dina(n4556),.dinb(w_n3668_0[0]),.dout(n4557),.clk(gclk));
	jnot g3916(.din(w_n3876_0[0]),.dout(n4558),.clk(gclk));
	jand g3917(.dina(n4558),.dinb(n4557),.dout(n4559),.clk(gclk));
	jand g3918(.dina(n4559),.dinb(n4493),.dout(n4560),.clk(gclk));
	jor g3919(.dina(w_n3883_0[0]),.dinb(n4560),.dout(n4561),.clk(gclk));
	jand g3920(.dina(n4561),.dinb(n4492),.dout(n4562),.clk(gclk));
	jor g3921(.dina(n4562),.dinb(w_n3643_0[0]),.dout(n4563),.clk(gclk));
	jnot g3922(.din(w_n3895_0[0]),.dout(n4564),.clk(gclk));
	jand g3923(.dina(n4564),.dinb(n4563),.dout(n4565),.clk(gclk));
	jand g3924(.dina(n4565),.dinb(n4491),.dout(n4566),.clk(gclk));
	jor g3925(.dina(w_n3902_0[0]),.dinb(n4566),.dout(n4567),.clk(gclk));
	jand g3926(.dina(n4567),.dinb(n4490),.dout(n4568),.clk(gclk));
	jor g3927(.dina(n4568),.dinb(w_n3624_0[0]),.dout(n4569),.clk(gclk));
	jnot g3928(.din(w_n3911_0[0]),.dout(n4570),.clk(gclk));
	jand g3929(.dina(n4570),.dinb(n4569),.dout(n4571),.clk(gclk));
	jor g3930(.dina(n4571),.dinb(w_n3615_0[0]),.dout(n4572),.clk(gclk));
	jnot g3931(.din(w_n3915_0[0]),.dout(n4573),.clk(gclk));
	jand g3932(.dina(n4573),.dinb(n4572),.dout(n4574),.clk(gclk));
	jand g3933(.dina(n4574),.dinb(n4489),.dout(n4575),.clk(gclk));
	jor g3934(.dina(w_n3928_0[0]),.dinb(n4575),.dout(n4576),.clk(gclk));
	jnot g3935(.din(w_n3935_0[0]),.dout(n4577),.clk(gclk));
	jand g3936(.dina(n4577),.dinb(n4576),.dout(n4578),.clk(gclk));
	jor g3937(.dina(n4578),.dinb(w_n3589_0[0]),.dout(n4579),.clk(gclk));
	jand g3938(.dina(n4579),.dinb(n4488),.dout(n4580),.clk(gclk));
	jor g3939(.dina(w_n3949_0[0]),.dinb(n4580),.dout(n4581),.clk(gclk));
	jnot g3940(.din(w_n3956_0[0]),.dout(n4582),.clk(gclk));
	jand g3941(.dina(n4582),.dinb(n4581),.dout(n4583),.clk(gclk));
	jor g3942(.dina(n4583),.dinb(w_n3572_0[0]),.dout(n4584),.clk(gclk));
	jand g3943(.dina(w_n3965_0[0]),.dinb(n4584),.dout(n4585),.clk(gclk));
	jand g3944(.dina(n4585),.dinb(w_n3534_0[0]),.dout(n4586),.clk(gclk));
	jor g3945(.dina(n4586),.dinb(w_n3563_0[0]),.dout(n4587),.clk(gclk));
	jnot g3946(.din(w_n4000_0[0]),.dout(n4588),.clk(gclk));
	jand g3947(.dina(n4588),.dinb(n4587),.dout(n4589),.clk(gclk));
	jor g3948(.dina(w_n4028_0[0]),.dinb(n4589),.dout(n4590),.clk(gclk));
	jor g3949(.dina(n4590),.dinb(w_n3465_0[0]),.dout(n4591),.clk(gclk));
	jnot g3950(.din(w_n4096_0[0]),.dout(n4592),.clk(gclk));
	jand g3951(.dina(n4592),.dinb(n4591),.dout(n4593),.clk(gclk));
	jor g3952(.dina(w_n4125_0[0]),.dinb(n4593),.dout(n4594),.clk(gclk));
	jor g3953(.dina(n4594),.dinb(w_n3417_0[0]),.dout(n4595),.clk(gclk));
	jnot g3954(.din(w_n4133_0[0]),.dout(n4596),.clk(gclk));
	jand g3955(.dina(n4596),.dinb(n4595),.dout(n4597),.clk(gclk));
	jor g3956(.dina(w_n4149_0[0]),.dinb(n4597),.dout(n4598),.clk(gclk));
	jor g3957(.dina(n4598),.dinb(w_n3408_0[0]),.dout(n4599),.clk(gclk));
	jnot g3958(.din(w_n4155_0[0]),.dout(n4600),.clk(gclk));
	jand g3959(.dina(n4600),.dinb(n4599),.dout(n4601),.clk(gclk));
	jor g3960(.dina(n4601),.dinb(w_n3324_0[0]),.dout(n4602),.clk(gclk));
	jnot g3961(.din(w_n4162_0[0]),.dout(n4603),.clk(gclk));
	jand g3962(.dina(n4603),.dinb(n4602),.dout(n4604),.clk(gclk));
	jor g3963(.dina(n4604),.dinb(w_n3293_0[0]),.dout(n4605),.clk(gclk));
	jnot g3964(.din(w_n4167_0[0]),.dout(n4606),.clk(gclk));
	jand g3965(.dina(n4606),.dinb(n4605),.dout(n4607),.clk(gclk));
	jor g3966(.dina(n4607),.dinb(w_n3284_0[0]),.dout(n4608),.clk(gclk));
	jand g3967(.dina(w_n4207_0[0]),.dinb(n4608),.dout(n4609),.clk(gclk));
	jor g3968(.dina(w_n4222_0[0]),.dinb(n4609),.dout(n4610),.clk(gclk));
	jand g3969(.dina(n4610),.dinb(n4487),.dout(n4611),.clk(gclk));
	jor g3970(.dina(w_n4240_0[0]),.dinb(n4611),.dout(n4612),.clk(gclk));
	jand g3971(.dina(n4612),.dinb(n4486),.dout(n4613),.clk(gclk));
	jor g3972(.dina(w_n4255_0[0]),.dinb(n4613),.dout(n4614),.clk(gclk));
	jor g3973(.dina(n4614),.dinb(w_n3172_0[0]),.dout(n4615),.clk(gclk));
	jnot g3974(.din(w_n4261_0[0]),.dout(n4616),.clk(gclk));
	jand g3975(.dina(n4616),.dinb(n4615),.dout(n4617),.clk(gclk));
	jor g3976(.dina(n4617),.dinb(w_n3163_0[0]),.dout(n4618),.clk(gclk));
	jor g3977(.dina(n4618),.dinb(w_n3155_0[0]),.dout(n4619),.clk(gclk));
	jand g3978(.dina(n4619),.dinb(n4485),.dout(n4620),.clk(gclk));
	jor g3979(.dina(w_n4280_0[0]),.dinb(n4620),.dout(n4621),.clk(gclk));
	jand g3980(.dina(n4621),.dinb(n4484),.dout(n4622),.clk(gclk));
	jor g3981(.dina(w_n4298_0[0]),.dinb(n4622),.dout(n4623),.clk(gclk));
	jand g3982(.dina(n4623),.dinb(n4483),.dout(n4624),.clk(gclk));
	jor g3983(.dina(w_n4316_0[0]),.dinb(n4624),.dout(n4625),.clk(gclk));
	jand g3984(.dina(n4625),.dinb(n4482),.dout(n4626),.clk(gclk));
	jor g3985(.dina(w_n4334_0[0]),.dinb(n4626),.dout(n4627),.clk(gclk));
	jand g3986(.dina(n4627),.dinb(n4481),.dout(n4628),.clk(gclk));
	jor g3987(.dina(w_n4352_0[0]),.dinb(n4628),.dout(n4629),.clk(gclk));
	jand g3988(.dina(n4629),.dinb(n4480),.dout(n4630),.clk(gclk));
	jor g3989(.dina(w_n4362_0[0]),.dinb(n4630),.dout(n4631),.clk(gclk));
	jor g3990(.dina(n4631),.dinb(w_n2937_0[0]),.dout(n4632),.clk(gclk));
	jnot g3991(.din(w_n4394_0[0]),.dout(n4633),.clk(gclk));
	jand g3992(.dina(n4633),.dinb(n4632),.dout(n4634),.clk(gclk));
	jor g3993(.dina(w_n4407_0[0]),.dinb(n4634),.dout(n4635),.clk(gclk));
	jor g3994(.dina(n4635),.dinb(w_n2897_0[0]),.dout(n4636),.clk(gclk));
	jnot g3995(.din(w_n4413_0[0]),.dout(n4637),.clk(gclk));
	jand g3996(.dina(n4637),.dinb(n4636),.dout(n4638),.clk(gclk));
	jor g3997(.dina(n4638),.dinb(w_n2888_0[0]),.dout(n4639),.clk(gclk));
	jand g3998(.dina(w_n4453_0[0]),.dinb(n4639),.dout(n4640),.clk(gclk));
	jor g3999(.dina(w_n4468_0[0]),.dinb(n4640),.dout(n4641),.clk(gclk));
	jand g4000(.dina(n4641),.dinb(n4479),.dout(n4642),.clk(gclk));
	jor g4001(.dina(n4642),.dinb(w_n2837_0[0]),.dout(n4643),.clk(gclk));
	jand g4002(.dina(n4643),.dinb(n4478),.dout(n4644),.clk(gclk));
	jor g4003(.dina(w_n4644_0[1]),.dinb(w_n2641_0[1]),.dout(n4645),.clk(gclk));
	jnot g4004(.din(w_n2643_0[2]),.dout(n4646),.clk(gclk));
	jor g4005(.dina(w_n4644_0[0]),.dinb(n4646),.dout(n4647),.clk(gclk));
	jand g4006(.dina(n4647),.dinb(n4645),.dout(n4648),.clk(gclk));
	jor g4007(.dina(w_n4648_63[1]),.dinb(w_n3771_0[0]),.dout(n4649),.clk(gclk));
	jand g4008(.dina(n4649),.dinb(n4477),.dout(result0),.clk(gclk));
	jor g4009(.dina(w_address1_63[0]),.dinb(w_n4506_0[0]),.dout(n4651),.clk(gclk));
	jor g4010(.dina(w_n4648_63[0]),.dinb(w_n3761_0[0]),.dout(n4652),.clk(gclk));
	jand g4011(.dina(n4652),.dinb(n4651),.dout(result1),.clk(gclk));
	jor g4012(.dina(w_address1_62[2]),.dinb(w_n4515_0[0]),.dout(n4654),.clk(gclk));
	jor g4013(.dina(w_n4648_62[2]),.dinb(w_n3779_0[0]),.dout(n4655),.clk(gclk));
	jand g4014(.dina(n4655),.dinb(n4654),.dout(result2),.clk(gclk));
	jor g4015(.dina(w_address1_62[1]),.dinb(w_n4526_0[0]),.dout(n4657),.clk(gclk));
	jor g4016(.dina(w_n4648_62[1]),.dinb(w_n3791_0[0]),.dout(n4658),.clk(gclk));
	jand g4017(.dina(n4658),.dinb(n4657),.dout(result3),.clk(gclk));
	jor g4018(.dina(w_address1_62[0]),.dinb(w_n3756_0[0]),.dout(n4660),.clk(gclk));
	jor g4019(.dina(w_n4648_62[0]),.dinb(w_n3795_0[0]),.dout(n4661),.clk(gclk));
	jand g4020(.dina(n4661),.dinb(n4660),.dout(result4),.clk(gclk));
	jor g4021(.dina(w_address1_61[2]),.dinb(w_n3745_0[0]),.dout(n4663),.clk(gclk));
	jor g4022(.dina(w_n4648_61[2]),.dinb(w_n3748_0[0]),.dout(n4664),.clk(gclk));
	jand g4023(.dina(n4664),.dinb(n4663),.dout(result5),.clk(gclk));
	jor g4024(.dina(w_address1_61[1]),.dinb(w_n3806_0[0]),.dout(n4666),.clk(gclk));
	jor g4025(.dina(w_n4648_61[1]),.dinb(w_n3734_0[0]),.dout(n4667),.clk(gclk));
	jand g4026(.dina(n4667),.dinb(n4666),.dout(result6),.clk(gclk));
	jor g4027(.dina(w_address1_61[0]),.dinb(w_n3804_0[0]),.dout(n4669),.clk(gclk));
	jor g4028(.dina(w_n4648_61[0]),.dinb(w_n3729_0[0]),.dout(n4670),.clk(gclk));
	jand g4029(.dina(n4670),.dinb(n4669),.dout(result7),.clk(gclk));
	jor g4030(.dina(w_address1_60[2]),.dinb(w_n3720_0[0]),.dout(n4672),.clk(gclk));
	jor g4031(.dina(w_n4648_60[2]),.dinb(w_n3811_0[0]),.dout(n4673),.clk(gclk));
	jand g4032(.dina(n4673),.dinb(n4672),.dout(result8),.clk(gclk));
	jor g4033(.dina(w_address1_60[1]),.dinb(w_n3821_0[0]),.dout(n4675),.clk(gclk));
	jor g4034(.dina(w_n4648_60[1]),.dinb(w_n3826_0[0]),.dout(n4676),.clk(gclk));
	jand g4035(.dina(n4676),.dinb(n4675),.dout(result9),.clk(gclk));
	jor g4036(.dina(w_address1_60[0]),.dinb(w_n3830_0[0]),.dout(n4678),.clk(gclk));
	jor g4037(.dina(w_n4648_60[0]),.dinb(w_n3712_0[0]),.dout(n4679),.clk(gclk));
	jand g4038(.dina(n4679),.dinb(n4678),.dout(result10),.clk(gclk));
	jor g4039(.dina(w_address1_59[2]),.dinb(w_n3835_0[0]),.dout(n4681),.clk(gclk));
	jor g4040(.dina(w_n4648_59[2]),.dinb(w_n3845_0[0]),.dout(n4682),.clk(gclk));
	jand g4041(.dina(n4682),.dinb(n4681),.dout(result11),.clk(gclk));
	jor g4042(.dina(w_address1_59[1]),.dinb(w_n3700_0[0]),.dout(n4684),.clk(gclk));
	jor g4043(.dina(w_n4648_59[1]),.dinb(w_n3843_0[0]),.dout(n4685),.clk(gclk));
	jand g4044(.dina(n4685),.dinb(n4684),.dout(result12),.clk(gclk));
	jor g4045(.dina(w_address1_59[0]),.dinb(w_n3689_0[0]),.dout(n4687),.clk(gclk));
	jor g4046(.dina(w_n4648_59[0]),.dinb(w_n3695_0[0]),.dout(n4688),.clk(gclk));
	jand g4047(.dina(n4688),.dinb(n4687),.dout(result13),.clk(gclk));
	jor g4048(.dina(w_address1_58[2]),.dinb(w_n3855_0[0]),.dout(n4690),.clk(gclk));
	jor g4049(.dina(w_n4648_58[2]),.dinb(w_n3684_0[0]),.dout(n4691),.clk(gclk));
	jand g4050(.dina(n4691),.dinb(n4690),.dout(result14),.clk(gclk));
	jor g4051(.dina(w_address1_58[1]),.dinb(w_n3853_0[0]),.dout(n4693),.clk(gclk));
	jor g4052(.dina(w_n4648_58[1]),.dinb(w_n3676_0[0]),.dout(n4694),.clk(gclk));
	jand g4053(.dina(n4694),.dinb(n4693),.dout(result15),.clk(gclk));
	jor g4054(.dina(w_address1_58[0]),.dinb(w_n3667_0[0]),.dout(n4696),.clk(gclk));
	jor g4055(.dina(w_n4648_58[0]),.dinb(w_n3860_0[0]),.dout(n4697),.clk(gclk));
	jand g4056(.dina(n4697),.dinb(n4696),.dout(result16),.clk(gclk));
	jor g4057(.dina(w_address1_57[2]),.dinb(w_n3870_0[0]),.dout(n4699),.clk(gclk));
	jor g4058(.dina(w_n4648_57[2]),.dinb(w_n3875_0[0]),.dout(n4700),.clk(gclk));
	jand g4059(.dina(n4700),.dinb(n4699),.dout(result17),.clk(gclk));
	jor g4060(.dina(w_address1_57[1]),.dinb(w_n3879_0[0]),.dout(n4702),.clk(gclk));
	jor g4061(.dina(w_n4648_57[1]),.dinb(w_n3659_0[0]),.dout(n4703),.clk(gclk));
	jand g4062(.dina(n4703),.dinb(n4702),.dout(result18),.clk(gclk));
	jor g4063(.dina(w_address1_57[0]),.dinb(w_n3881_0[0]),.dout(n4705),.clk(gclk));
	jor g4064(.dina(w_n4648_57[0]),.dinb(w_n3651_0[0]),.dout(n4706),.clk(gclk));
	jand g4065(.dina(n4706),.dinb(n4705),.dout(result19),.clk(gclk));
	jor g4066(.dina(w_address1_56[2]),.dinb(w_n3642_0[0]),.dout(n4708),.clk(gclk));
	jor g4067(.dina(w_n4648_56[2]),.dinb(w_n3640_0[0]),.dout(n4709),.clk(gclk));
	jand g4068(.dina(n4709),.dinb(n4708),.dout(result20),.clk(gclk));
	jor g4069(.dina(w_address1_56[1]),.dinb(w_n3898_0[0]),.dout(n4711),.clk(gclk));
	jor g4070(.dina(w_n4648_56[1]),.dinb(w_n3894_0[0]),.dout(n4712),.clk(gclk));
	jand g4071(.dina(n4712),.dinb(n4711),.dout(result21),.clk(gclk));
	jor g4072(.dina(w_address1_56[0]),.dinb(w_n3900_0[0]),.dout(n4714),.clk(gclk));
	jor g4073(.dina(w_n4648_56[0]),.dinb(w_n3632_0[0]),.dout(n4715),.clk(gclk));
	jand g4074(.dina(n4715),.dinb(n4714),.dout(result22),.clk(gclk));
	jor g4075(.dina(w_address1_55[2]),.dinb(w_n3620_0[0]),.dout(n4717),.clk(gclk));
	jor g4076(.dina(w_n4648_55[2]),.dinb(w_n3907_0[0]),.dout(n4718),.clk(gclk));
	jand g4077(.dina(n4718),.dinb(n4717),.dout(result23),.clk(gclk));
	jor g4078(.dina(w_address1_55[1]),.dinb(w_n3605_0[0]),.dout(n4720),.clk(gclk));
	jor g4079(.dina(w_n4648_55[1]),.dinb(w_n3909_0[0]),.dout(n4721),.clk(gclk));
	jand g4080(.dina(n4721),.dinb(n4720),.dout(result24),.clk(gclk));
	jor g4081(.dina(w_address1_55[0]),.dinb(w_n3613_0[0]),.dout(n4723),.clk(gclk));
	jor g4082(.dina(w_n4648_55[0]),.dinb(w_n3914_0[0]),.dout(n4724),.clk(gclk));
	jand g4083(.dina(n4724),.dinb(n4723),.dout(result25),.clk(gclk));
	jor g4084(.dina(w_address1_54[2]),.dinb(w_n3918_0[0]),.dout(n4726),.clk(gclk));
	jor g4085(.dina(w_n4648_54[2]),.dinb(w_n3597_0[0]),.dout(n4727),.clk(gclk));
	jand g4086(.dina(n4727),.dinb(n4726),.dout(result26),.clk(gclk));
	jor g4087(.dina(w_address1_54[1]),.dinb(w_n3923_0[0]),.dout(n4729),.clk(gclk));
	jor g4088(.dina(w_n4648_54[1]),.dinb(w_n3933_0[0]),.dout(n4730),.clk(gclk));
	jand g4089(.dina(n4730),.dinb(n4729),.dout(result27),.clk(gclk));
	jor g4090(.dina(w_address1_54[0]),.dinb(w_n3585_0[0]),.dout(n4732),.clk(gclk));
	jor g4091(.dina(w_n4648_54[0]),.dinb(w_n3931_0[0]),.dout(n4733),.clk(gclk));
	jand g4092(.dina(n4733),.dinb(n4732),.dout(result28),.clk(gclk));
	jor g4093(.dina(w_address1_53[2]),.dinb(w_n3947_0[0]),.dout(n4735),.clk(gclk));
	jor g4094(.dina(w_n4648_53[2]),.dinb(w_n3580_0[0]),.dout(n4736),.clk(gclk));
	jand g4095(.dina(n4736),.dinb(n4735),.dout(result29),.clk(gclk));
	jor g4096(.dina(w_address1_53[1]),.dinb(w_n3942_0[0]),.dout(n4738),.clk(gclk));
	jor g4097(.dina(w_n4648_53[1]),.dinb(w_n3954_0[0]),.dout(n4739),.clk(gclk));
	jand g4098(.dina(n4739),.dinb(n4738),.dout(result30),.clk(gclk));
	jor g4099(.dina(w_address1_53[0]),.dinb(w_n3568_0[0]),.dout(n4741),.clk(gclk));
	jor g4100(.dina(w_n4648_53[0]),.dinb(w_n3952_0[0]),.dout(n4742),.clk(gclk));
	jand g4101(.dina(n4742),.dinb(n4741),.dout(result31),.clk(gclk));
	jor g4102(.dina(w_address1_52[2]),.dinb(w_n3541_0[0]),.dout(n4744),.clk(gclk));
	jor g4103(.dina(w_n4648_52[2]),.dinb(w_n3960_0[0]),.dout(n4745),.clk(gclk));
	jand g4104(.dina(n4745),.dinb(n4744),.dout(result32),.clk(gclk));
	jor g4105(.dina(w_address1_52[1]),.dinb(w_n3543_0[0]),.dout(n4747),.clk(gclk));
	jor g4106(.dina(w_n4648_52[1]),.dinb(w_n3523_0[0]),.dout(n4748),.clk(gclk));
	jand g4107(.dina(n4748),.dinb(n4747),.dout(result33),.clk(gclk));
	jor g4108(.dina(w_address1_52[0]),.dinb(w_n3549_0[0]),.dout(n4750),.clk(gclk));
	jor g4109(.dina(w_n4648_52[0]),.dinb(w_n3528_0[0]),.dout(n4751),.clk(gclk));
	jand g4110(.dina(n4751),.dinb(n4750),.dout(result34),.clk(gclk));
	jor g4111(.dina(w_address1_51[2]),.dinb(w_n3547_0[0]),.dout(n4753),.clk(gclk));
	jor g4112(.dina(w_n4648_51[2]),.dinb(w_n3514_0[0]),.dout(n4754),.clk(gclk));
	jand g4113(.dina(n4754),.dinb(n4753),.dout(result35),.clk(gclk));
	jor g4114(.dina(w_address1_51[1]),.dinb(w_n3499_0[0]),.dout(n4756),.clk(gclk));
	jor g4115(.dina(w_n4648_51[1]),.dinb(w_n3505_0[0]),.dout(n4757),.clk(gclk));
	jand g4116(.dina(n4757),.dinb(n4756),.dout(result36),.clk(gclk));
	jor g4117(.dina(w_address1_51[0]),.dinb(w_n3494_0[0]),.dout(n4759),.clk(gclk));
	jor g4118(.dina(w_n4648_51[0]),.dinb(w_n3490_0[0]),.dout(n4760),.clk(gclk));
	jand g4119(.dina(n4760),.dinb(n4759),.dout(result37),.clk(gclk));
	jor g4120(.dina(w_address1_50[2]),.dinb(w_n3559_0[0]),.dout(n4762),.clk(gclk));
	jor g4121(.dina(w_n4648_50[2]),.dinb(w_n3479_0[0]),.dout(n4763),.clk(gclk));
	jand g4122(.dina(n4763),.dinb(n4762),.dout(result38),.clk(gclk));
	jor g4123(.dina(w_address1_50[1]),.dinb(w_n3557_0[0]),.dout(n4765),.clk(gclk));
	jor g4124(.dina(w_n4648_50[1]),.dinb(w_n3473_0[0]),.dout(n4766),.clk(gclk));
	jand g4125(.dina(n4766),.dinb(n4765),.dout(result39),.clk(gclk));
	jor g4126(.dina(w_address1_50[0]),.dinb(w_n4005_0[0]),.dout(n4768),.clk(gclk));
	jor g4127(.dina(w_n4648_50[0]),.dinb(w_n3984_0[0]),.dout(n4769),.clk(gclk));
	jand g4128(.dina(n4769),.dinb(n4768),.dout(result40),.clk(gclk));
	jor g4129(.dina(w_address1_49[2]),.dinb(w_n4008_0[0]),.dout(n4771),.clk(gclk));
	jor g4130(.dina(w_n4648_49[2]),.dinb(w_n3976_0[0]),.dout(n4772),.clk(gclk));
	jand g4131(.dina(n4772),.dinb(n4771),.dout(result41),.clk(gclk));
	jor g4132(.dina(w_address1_49[1]),.dinb(w_n4002_0[0]),.dout(n4774),.clk(gclk));
	jor g4133(.dina(w_n4648_49[1]),.dinb(w_n3992_0[0]),.dout(n4775),.clk(gclk));
	jand g4134(.dina(n4775),.dinb(n4774),.dout(result42),.clk(gclk));
	jor g4135(.dina(w_address1_49[0]),.dinb(w_n3463_0[0]),.dout(n4777),.clk(gclk));
	jnot g4136(.din(w_n3421_0[0]),.dout(n4778),.clk(gclk));
	jor g4137(.dina(w_n4648_49[0]),.dinb(n4778),.dout(n4779),.clk(gclk));
	jand g4138(.dina(n4779),.dinb(n4777),.dout(result43),.clk(gclk));
	jor g4139(.dina(w_address1_48[2]),.dinb(w_n4015_0[0]),.dout(n4781),.clk(gclk));
	jor g4140(.dina(w_n4648_48[2]),.dinb(w_n3428_0[0]),.dout(n4782),.clk(gclk));
	jand g4141(.dina(n4782),.dinb(n4781),.dout(result44),.clk(gclk));
	jor g4142(.dina(w_address1_48[1]),.dinb(w_n4013_0[0]),.dout(n4784),.clk(gclk));
	jor g4143(.dina(w_n4648_48[1]),.dinb(w_n3455_0[0]),.dout(n4785),.clk(gclk));
	jand g4144(.dina(n4785),.dinb(n4784),.dout(result45),.clk(gclk));
	jor g4145(.dina(w_address1_48[0]),.dinb(w_n4023_0[0]),.dout(n4787),.clk(gclk));
	jor g4146(.dina(w_n4648_48[0]),.dinb(w_n3442_0[0]),.dout(n4788),.clk(gclk));
	jand g4147(.dina(n4788),.dinb(n4787),.dout(result46),.clk(gclk));
	jor g4148(.dina(w_address1_47[2]),.dinb(w_n4021_0[0]),.dout(n4790),.clk(gclk));
	jor g4149(.dina(w_n4648_47[2]),.dinb(w_n3437_0[0]),.dout(n4791),.clk(gclk));
	jand g4150(.dina(n4791),.dinb(n4790),.dout(result47),.clk(gclk));
	jor g4151(.dina(w_address1_47[1]),.dinb(w_n4108_0[0]),.dout(n4793),.clk(gclk));
	jor g4152(.dina(w_n4648_47[1]),.dinb(w_n4080_0[0]),.dout(n4794),.clk(gclk));
	jand g4153(.dina(n4794),.dinb(n4793),.dout(result48),.clk(gclk));
	jor g4154(.dina(w_address1_47[0]),.dinb(w_n4110_0[0]),.dout(n4796),.clk(gclk));
	jor g4155(.dina(w_n4648_47[0]),.dinb(w_n4038_0[0]),.dout(n4797),.clk(gclk));
	jand g4156(.dina(n4797),.dinb(n4796),.dout(result49),.clk(gclk));
	jor g4157(.dina(w_address1_46[2]),.dinb(w_n4116_0[0]),.dout(n4799),.clk(gclk));
	jor g4158(.dina(w_n4648_46[2]),.dinb(w_n4043_0[0]),.dout(n4800),.clk(gclk));
	jand g4159(.dina(n4800),.dinb(n4799),.dout(result50),.clk(gclk));
	jor g4160(.dina(w_address1_46[1]),.dinb(w_n4114_0[0]),.dout(n4802),.clk(gclk));
	jor g4161(.dina(w_n4648_46[1]),.dinb(w_n4091_0[0]),.dout(n4803),.clk(gclk));
	jand g4162(.dina(n4803),.dinb(n4802),.dout(result51),.clk(gclk));
	jor g4163(.dina(w_address1_46[0]),.dinb(w_n4104_0[0]),.dout(n4805),.clk(gclk));
	jor g4164(.dina(w_n4648_46[0]),.dinb(w_n4052_0[0]),.dout(n4806),.clk(gclk));
	jand g4165(.dina(n4806),.dinb(n4805),.dout(result52),.clk(gclk));
	jor g4166(.dina(w_address1_45[2]),.dinb(w_n4099_0[0]),.dout(n4808),.clk(gclk));
	jor g4167(.dina(w_n4648_45[2]),.dinb(w_n4063_0[0]),.dout(n4809),.clk(gclk));
	jand g4168(.dina(n4809),.dinb(n4808),.dout(result53),.clk(gclk));
	jor g4169(.dina(w_address1_45[1]),.dinb(w_n4101_0[0]),.dout(n4811),.clk(gclk));
	jor g4170(.dina(w_n4648_45[1]),.dinb(w_n4071_0[0]),.dout(n4812),.clk(gclk));
	jand g4171(.dina(n4812),.dinb(n4811),.dout(result54),.clk(gclk));
	jor g4172(.dina(w_address1_45[0]),.dinb(w_n3413_0[0]),.dout(n4814),.clk(gclk));
	jor g4173(.dina(w_n4648_45[0]),.dinb(w_n4066_0[0]),.dout(n4815),.clk(gclk));
	jand g4174(.dina(n4815),.dinb(n4814),.dout(result55),.clk(gclk));
	jor g4175(.dina(w_address1_44[2]),.dinb(w_n3396_0[0]),.dout(n4817),.clk(gclk));
	jor g4176(.dina(w_n4648_44[2]),.dinb(w_n4129_0[0]),.dout(n4818),.clk(gclk));
	jand g4177(.dina(n4818),.dinb(n4817),.dout(result56),.clk(gclk));
	jor g4178(.dina(w_address1_44[1]),.dinb(w_n3402_0[0]),.dout(n4820),.clk(gclk));
	jor g4179(.dina(w_n4648_44[1]),.dinb(w_n3390_0[0]),.dout(n4821),.clk(gclk));
	jand g4180(.dina(n4821),.dinb(n4820),.dout(result57),.clk(gclk));
	jor g4181(.dina(w_address1_44[0]),.dinb(w_n3382_0[0]),.dout(n4823),.clk(gclk));
	jor g4182(.dina(w_n4648_44[0]),.dinb(w_n3378_0[0]),.dout(n4824),.clk(gclk));
	jand g4183(.dina(n4824),.dinb(n4823),.dout(result58),.clk(gclk));
	jor g4184(.dina(w_address1_43[2]),.dinb(w_n3365_0[0]),.dout(n4826),.clk(gclk));
	jor g4185(.dina(w_n4648_43[2]),.dinb(w_n3370_0[0]),.dout(n4827),.clk(gclk));
	jand g4186(.dina(n4827),.dinb(n4826),.dout(result59),.clk(gclk));
	jor g4187(.dina(w_address1_43[1]),.dinb(w_n4138_0[0]),.dout(n4829),.clk(gclk));
	jor g4188(.dina(w_n4648_43[1]),.dinb(w_n3332_0[0]),.dout(n4830),.clk(gclk));
	jand g4189(.dina(n4830),.dinb(n4829),.dout(result60),.clk(gclk));
	jor g4190(.dina(w_address1_43[0]),.dinb(w_n4136_0[0]),.dout(n4832),.clk(gclk));
	jor g4191(.dina(w_n4648_43[0]),.dinb(w_n3356_0[0]),.dout(n4833),.clk(gclk));
	jand g4192(.dina(n4833),.dinb(n4832),.dout(result61),.clk(gclk));
	jor g4193(.dina(w_address1_42[2]),.dinb(w_n4145_0[0]),.dout(n4835),.clk(gclk));
	jor g4194(.dina(w_n4648_42[2]),.dinb(w_n3337_0[0]),.dout(n4836),.clk(gclk));
	jand g4195(.dina(n4836),.dinb(n4835),.dout(result62),.clk(gclk));
	jor g4196(.dina(w_address1_42[1]),.dinb(w_n4143_0[0]),.dout(n4838),.clk(gclk));
	jor g4197(.dina(w_n4648_42[1]),.dinb(w_n3348_0[0]),.dout(n4839),.clk(gclk));
	jand g4198(.dina(n4839),.dinb(n4838),.dout(result63),.clk(gclk));
	jor g4199(.dina(w_address1_42[0]),.dinb(w_n3320_0[0]),.dout(n4841),.clk(gclk));
	jor g4200(.dina(w_n4648_42[0]),.dinb(w_n4153_0[0]),.dout(n4842),.clk(gclk));
	jand g4201(.dina(n4842),.dinb(n4841),.dout(result64),.clk(gclk));
	jor g4202(.dina(w_address1_41[2]),.dinb(w_n3306_0[0]),.dout(n4844),.clk(gclk));
	jor g4203(.dina(w_n4648_41[2]),.dinb(w_n3311_0[0]),.dout(n4845),.clk(gclk));
	jand g4204(.dina(n4845),.dinb(n4844),.dout(result65),.clk(gclk));
	jor g4205(.dina(w_address1_41[1]),.dinb(w_n3301_0[0]),.dout(n4847),.clk(gclk));
	jor g4206(.dina(w_n4648_41[1]),.dinb(w_n4160_0[0]),.dout(n4848),.clk(gclk));
	jand g4207(.dina(n4848),.dinb(n4847),.dout(result66),.clk(gclk));
	jor g4208(.dina(w_address1_41[0]),.dinb(w_n3289_0[0]),.dout(n4850),.clk(gclk));
	jor g4209(.dina(w_n4648_41[0]),.dinb(w_n4158_0[0]),.dout(n4851),.clk(gclk));
	jand g4210(.dina(n4851),.dinb(n4850),.dout(result67),.clk(gclk));
	jor g4211(.dina(w_address1_40[2]),.dinb(w_n3270_0[0]),.dout(n4853),.clk(gclk));
	jor g4212(.dina(w_n4648_40[2]),.dinb(w_n4165_0[0]),.dout(n4854),.clk(gclk));
	jand g4213(.dina(n4854),.dinb(n4853),.dout(result68),.clk(gclk));
	jor g4214(.dina(w_address1_40[1]),.dinb(w_n3265_0[0]),.dout(n4856),.clk(gclk));
	jor g4215(.dina(w_n4648_40[1]),.dinb(w_n3260_0[0]),.dout(n4857),.clk(gclk));
	jand g4216(.dina(n4857),.dinb(n4856),.dout(result69),.clk(gclk));
	jor g4217(.dina(w_address1_40[0]),.dinb(w_n3280_0[0]),.dout(n4859),.clk(gclk));
	jor g4218(.dina(w_n4648_40[0]),.dinb(w_n3241_0[0]),.dout(n4860),.clk(gclk));
	jand g4219(.dina(n4860),.dinb(n4859),.dout(result70),.clk(gclk));
	jor g4220(.dina(w_address1_39[2]),.dinb(w_n3278_0[0]),.dout(n4862),.clk(gclk));
	jor g4221(.dina(w_n4648_39[2]),.dinb(w_n3252_0[0]),.dout(n4863),.clk(gclk));
	jand g4222(.dina(n4863),.dinb(n4862),.dout(result71),.clk(gclk));
	jor g4223(.dina(w_address1_39[1]),.dinb(w_n4214_0[0]),.dout(n4865),.clk(gclk));
	jor g4224(.dina(w_n4648_39[1]),.dinb(w_n4173_0[0]),.dout(n4866),.clk(gclk));
	jand g4225(.dina(n4866),.dinb(n4865),.dout(result72),.clk(gclk));
	jor g4226(.dina(w_address1_39[0]),.dinb(w_n4217_0[0]),.dout(n4868),.clk(gclk));
	jor g4227(.dina(w_n4648_39[0]),.dinb(w_n4203_0[0]),.dout(n4869),.clk(gclk));
	jand g4228(.dina(n4869),.dinb(n4868),.dout(result73),.clk(gclk));
	jor g4229(.dina(w_address1_38[2]),.dinb(w_n4212_0[0]),.dout(n4871),.clk(gclk));
	jor g4230(.dina(w_n4648_38[2]),.dinb(w_n4190_0[0]),.dout(n4872),.clk(gclk));
	jand g4231(.dina(n4872),.dinb(n4871),.dout(result74),.clk(gclk));
	jor g4232(.dina(w_address1_38[1]),.dinb(w_n4210_0[0]),.dout(n4874),.clk(gclk));
	jor g4233(.dina(w_n4648_38[1]),.dinb(w_n4185_0[0]),.dout(n4875),.clk(gclk));
	jand g4234(.dina(n4875),.dinb(n4874),.dout(result75),.clk(gclk));
	jor g4235(.dina(w_address1_38[0]),.dinb(w_n4229_0[0]),.dout(n4877),.clk(gclk));
	jor g4236(.dina(w_n4648_38[0]),.dinb(w_n3209_0[0]),.dout(n4878),.clk(gclk));
	jand g4237(.dina(n4878),.dinb(n4877),.dout(result76),.clk(gclk));
	jor g4238(.dina(w_address1_37[2]),.dinb(w_n4227_0[0]),.dout(n4880),.clk(gclk));
	jor g4239(.dina(w_n4648_37[2]),.dinb(w_n3233_0[0]),.dout(n4881),.clk(gclk));
	jand g4240(.dina(n4881),.dinb(n4880),.dout(result77),.clk(gclk));
	jor g4241(.dina(w_address1_37[1]),.dinb(w_n4236_0[0]),.dout(n4883),.clk(gclk));
	jor g4242(.dina(w_n4648_37[1]),.dinb(w_n3214_0[0]),.dout(n4884),.clk(gclk));
	jand g4243(.dina(n4884),.dinb(n4883),.dout(result78),.clk(gclk));
	jor g4244(.dina(w_address1_37[0]),.dinb(w_n4234_0[0]),.dout(n4886),.clk(gclk));
	jor g4245(.dina(w_n4648_37[0]),.dinb(w_n3225_0[0]),.dout(n4887),.clk(gclk));
	jand g4246(.dina(n4887),.dinb(n4886),.dout(result79),.clk(gclk));
	jor g4247(.dina(w_address1_36[2]),.dinb(w_n4248_0[0]),.dout(n4889),.clk(gclk));
	jor g4248(.dina(w_n4648_36[2]),.dinb(w_n3196_0[0]),.dout(n4890),.clk(gclk));
	jand g4249(.dina(n4890),.dinb(n4889),.dout(result80),.clk(gclk));
	jor g4250(.dina(w_address1_36[1]),.dinb(w_n4251_0[0]),.dout(n4892),.clk(gclk));
	jor g4251(.dina(w_n4648_36[1]),.dinb(w_n3191_0[0]),.dout(n4893),.clk(gclk));
	jand g4252(.dina(n4893),.dinb(n4892),.dout(result81),.clk(gclk));
	jor g4253(.dina(w_address1_36[0]),.dinb(w_n4245_0[0]),.dout(n4895),.clk(gclk));
	jor g4254(.dina(w_n4648_36[0]),.dinb(w_n3179_0[0]),.dout(n4896),.clk(gclk));
	jand g4255(.dina(n4896),.dinb(n4895),.dout(result82),.clk(gclk));
	jor g4256(.dina(w_address1_35[2]),.dinb(w_n3168_0[0]),.dout(n4898),.clk(gclk));
	jor g4257(.dina(w_n4648_35[2]),.dinb(w_n3174_0[0]),.dout(n4899),.clk(gclk));
	jand g4258(.dina(n4899),.dinb(n4898),.dout(result83),.clk(gclk));
	jor g4259(.dina(w_address1_35[1]),.dinb(w_n3149_0[0]),.dout(n4901),.clk(gclk));
	jor g4260(.dina(w_n4648_35[1]),.dinb(w_n4259_0[0]),.dout(n4902),.clk(gclk));
	jand g4261(.dina(n4902),.dinb(n4901),.dout(result84),.clk(gclk));
	jor g4262(.dina(w_address1_35[0]),.dinb(w_n3144_0[0]),.dout(n4904),.clk(gclk));
	jor g4263(.dina(w_n4648_35[0]),.dinb(w_n3139_0[0]),.dout(n4905),.clk(gclk));
	jand g4264(.dina(n4905),.dinb(n4904),.dout(result85),.clk(gclk));
	jor g4265(.dina(w_address1_34[2]),.dinb(w_n3160_0[0]),.dout(n4907),.clk(gclk));
	jor g4266(.dina(w_n4648_34[2]),.dinb(w_n3120_0[0]),.dout(n4908),.clk(gclk));
	jand g4267(.dina(n4908),.dinb(n4907),.dout(result86),.clk(gclk));
	jor g4268(.dina(w_address1_34[1]),.dinb(w_n3158_0[0]),.dout(n4910),.clk(gclk));
	jor g4269(.dina(w_n4648_34[1]),.dinb(w_n3131_0[0]),.dout(n4911),.clk(gclk));
	jand g4270(.dina(n4911),.dinb(n4910),.dout(result87),.clk(gclk));
	jor g4271(.dina(w_address1_34[0]),.dinb(w_n4272_0[0]),.dout(n4913),.clk(gclk));
	jor g4272(.dina(w_n4648_34[0]),.dinb(w_n3110_0[0]),.dout(n4914),.clk(gclk));
	jand g4273(.dina(n4914),.dinb(n4913),.dout(result88),.clk(gclk));
	jor g4274(.dina(w_address1_33[2]),.dinb(w_n4275_0[0]),.dout(n4916),.clk(gclk));
	jor g4275(.dina(w_n4648_33[2]),.dinb(w_n3105_0[0]),.dout(n4917),.clk(gclk));
	jand g4276(.dina(n4917),.dinb(n4916),.dout(result89),.clk(gclk));
	jor g4277(.dina(w_address1_33[1]),.dinb(w_n4269_0[0]),.dout(n4919),.clk(gclk));
	jor g4278(.dina(w_n4648_33[1]),.dinb(w_n3093_0[0]),.dout(n4920),.clk(gclk));
	jand g4279(.dina(n4920),.dinb(n4919),.dout(result90),.clk(gclk));
	jor g4280(.dina(w_address1_33[0]),.dinb(w_n4266_0[0]),.dout(n4922),.clk(gclk));
	jor g4281(.dina(w_n4648_33[0]),.dinb(w_n3088_0[0]),.dout(n4923),.clk(gclk));
	jand g4282(.dina(n4923),.dinb(n4922),.dout(result91),.clk(gclk));
	jor g4283(.dina(w_address1_32[2]),.dinb(w_n4287_0[0]),.dout(n4925),.clk(gclk));
	jor g4284(.dina(w_n4648_32[2]),.dinb(w_n3053_0[0]),.dout(n4926),.clk(gclk));
	jand g4285(.dina(n4926),.dinb(n4925),.dout(result92),.clk(gclk));
	jor g4286(.dina(w_address1_32[1]),.dinb(w_n4285_0[0]),.dout(n4928),.clk(gclk));
	jor g4287(.dina(w_n4648_32[1]),.dinb(w_n3077_0[0]),.dout(n4929),.clk(gclk));
	jand g4288(.dina(n4929),.dinb(n4928),.dout(result93),.clk(gclk));
	jor g4289(.dina(w_address1_32[0]),.dinb(w_n4294_0[0]),.dout(n4931),.clk(gclk));
	jor g4290(.dina(w_n4648_32[0]),.dinb(w_n3058_0[0]),.dout(n4932),.clk(gclk));
	jand g4291(.dina(n4932),.dinb(n4931),.dout(result94),.clk(gclk));
	jor g4292(.dina(w_address1_31[2]),.dinb(w_n4292_0[0]),.dout(n4934),.clk(gclk));
	jor g4293(.dina(w_n4648_31[2]),.dinb(w_n3069_0[0]),.dout(n4935),.clk(gclk));
	jand g4294(.dina(n4935),.dinb(n4934),.dout(result95),.clk(gclk));
	jor g4295(.dina(w_address1_31[1]),.dinb(w_n4308_0[0]),.dout(n4937),.clk(gclk));
	jor g4296(.dina(w_n4648_31[1]),.dinb(w_n3040_0[0]),.dout(n4938),.clk(gclk));
	jand g4297(.dina(n4938),.dinb(n4937),.dout(result96),.clk(gclk));
	jor g4298(.dina(w_address1_31[0]),.dinb(w_n4311_0[0]),.dout(n4940),.clk(gclk));
	jor g4299(.dina(w_n4648_31[0]),.dinb(w_n3035_0[0]),.dout(n4941),.clk(gclk));
	jand g4300(.dina(n4941),.dinb(n4940),.dout(result97),.clk(gclk));
	jor g4301(.dina(w_address1_30[2]),.dinb(w_n4305_0[0]),.dout(n4943),.clk(gclk));
	jor g4302(.dina(w_n4648_30[2]),.dinb(w_n3023_0[0]),.dout(n4944),.clk(gclk));
	jand g4303(.dina(n4944),.dinb(n4943),.dout(result98),.clk(gclk));
	jor g4304(.dina(w_address1_30[1]),.dinb(w_n4302_0[0]),.dout(n4946),.clk(gclk));
	jor g4305(.dina(w_n4648_30[1]),.dinb(w_n3018_0[0]),.dout(n4947),.clk(gclk));
	jand g4306(.dina(n4947),.dinb(n4946),.dout(result99),.clk(gclk));
	jor g4307(.dina(w_address1_30[0]),.dinb(w_n4323_0[0]),.dout(n4949),.clk(gclk));
	jor g4308(.dina(w_n4648_30[0]),.dinb(w_n2983_0[0]),.dout(n4950),.clk(gclk));
	jand g4309(.dina(n4950),.dinb(n4949),.dout(result100),.clk(gclk));
	jor g4310(.dina(w_address1_29[2]),.dinb(w_n4321_0[0]),.dout(n4952),.clk(gclk));
	jor g4311(.dina(w_n4648_29[2]),.dinb(w_n3007_0[0]),.dout(n4953),.clk(gclk));
	jand g4312(.dina(n4953),.dinb(n4952),.dout(result101),.clk(gclk));
	jor g4313(.dina(w_address1_29[1]),.dinb(w_n4330_0[0]),.dout(n4955),.clk(gclk));
	jor g4314(.dina(w_n4648_29[1]),.dinb(w_n2988_0[0]),.dout(n4956),.clk(gclk));
	jand g4315(.dina(n4956),.dinb(n4955),.dout(result102),.clk(gclk));
	jor g4316(.dina(w_address1_29[0]),.dinb(w_n4328_0[0]),.dout(n4958),.clk(gclk));
	jor g4317(.dina(w_n4648_29[0]),.dinb(w_n2999_0[0]),.dout(n4959),.clk(gclk));
	jand g4318(.dina(n4959),.dinb(n4958),.dout(result103),.clk(gclk));
	jor g4319(.dina(w_address1_28[2]),.dinb(w_n4344_0[0]),.dout(n4961),.clk(gclk));
	jor g4320(.dina(w_n4648_28[2]),.dinb(w_n2970_0[0]),.dout(n4962),.clk(gclk));
	jand g4321(.dina(n4962),.dinb(n4961),.dout(result104),.clk(gclk));
	jor g4322(.dina(w_address1_28[1]),.dinb(w_n4347_0[0]),.dout(n4964),.clk(gclk));
	jor g4323(.dina(w_n4648_28[1]),.dinb(w_n2965_0[0]),.dout(n4965),.clk(gclk));
	jand g4324(.dina(n4965),.dinb(n4964),.dout(result105),.clk(gclk));
	jor g4325(.dina(w_address1_28[0]),.dinb(w_n4341_0[0]),.dout(n4967),.clk(gclk));
	jor g4326(.dina(w_n4648_28[0]),.dinb(w_n2953_0[0]),.dout(n4968),.clk(gclk));
	jand g4327(.dina(n4968),.dinb(n4967),.dout(result106),.clk(gclk));
	jor g4328(.dina(w_address1_27[2]),.dinb(w_n4338_0[0]),.dout(n4970),.clk(gclk));
	jor g4329(.dina(w_n4648_27[2]),.dinb(w_n2948_0[0]),.dout(n4971),.clk(gclk));
	jand g4330(.dina(n4971),.dinb(n4970),.dout(result107),.clk(gclk));
	jor g4331(.dina(w_address1_27[1]),.dinb(w_n2931_0[0]),.dout(n4973),.clk(gclk));
	jor g4332(.dina(w_n4648_27[1]),.dinb(w_n2939_0[0]),.dout(n4974),.clk(gclk));
	jand g4333(.dina(n4974),.dinb(n4973),.dout(result108),.clk(gclk));
	jor g4334(.dina(w_address1_27[0]),.dinb(w_n2926_0[0]),.dout(n4976),.clk(gclk));
	jor g4335(.dina(w_n4648_27[0]),.dinb(w_n2921_0[0]),.dout(n4977),.clk(gclk));
	jand g4336(.dina(n4977),.dinb(n4976),.dout(result109),.clk(gclk));
	jor g4337(.dina(w_address1_26[2]),.dinb(w_n4359_0[0]),.dout(n4979),.clk(gclk));
	jor g4338(.dina(w_n4648_26[2]),.dinb(w_n2902_0[0]),.dout(n4980),.clk(gclk));
	jand g4339(.dina(n4980),.dinb(n4979),.dout(result110),.clk(gclk));
	jor g4340(.dina(w_address1_26[1]),.dinb(w_n4357_0[0]),.dout(n4982),.clk(gclk));
	jor g4341(.dina(w_n4648_26[1]),.dinb(w_n2913_0[0]),.dout(n4983),.clk(gclk));
	jand g4342(.dina(n4983),.dinb(n4982),.dout(result111),.clk(gclk));
	jor g4343(.dina(w_address1_26[0]),.dinb(w_n4400_0[0]),.dout(n4985),.clk(gclk));
	jor g4344(.dina(w_n4648_26[0]),.dinb(w_n4388_0[0]),.dout(n4986),.clk(gclk));
	jand g4345(.dina(n4986),.dinb(n4985),.dout(result112),.clk(gclk));
	jor g4346(.dina(w_address1_25[2]),.dinb(w_n4403_0[0]),.dout(n4988),.clk(gclk));
	jor g4347(.dina(w_n4648_25[2]),.dinb(w_n4372_0[0]),.dout(n4989),.clk(gclk));
	jand g4348(.dina(n4989),.dinb(n4988),.dout(result113),.clk(gclk));
	jor g4349(.dina(w_address1_25[1]),.dinb(w_n4397_0[0]),.dout(n4991),.clk(gclk));
	jor g4350(.dina(w_n4648_25[1]),.dinb(w_n4379_0[0]),.dout(n4992),.clk(gclk));
	jand g4351(.dina(n4992),.dinb(n4991),.dout(result114),.clk(gclk));
	jor g4352(.dina(w_address1_25[0]),.dinb(w_n2893_0[0]),.dout(n4994),.clk(gclk));
	jor g4353(.dina(w_n4648_25[0]),.dinb(w_n4374_0[0]),.dout(n4995),.clk(gclk));
	jand g4354(.dina(n4995),.dinb(n4994),.dout(result115),.clk(gclk));
	jor g4355(.dina(w_address1_24[2]),.dinb(w_n2874_0[0]),.dout(n4997),.clk(gclk));
	jor g4356(.dina(w_n4648_24[2]),.dinb(w_n4411_0[0]),.dout(n4998),.clk(gclk));
	jand g4357(.dina(n4998),.dinb(n4997),.dout(result116),.clk(gclk));
	jor g4358(.dina(w_address1_24[1]),.dinb(w_n2869_0[0]),.dout(n5000),.clk(gclk));
	jor g4359(.dina(w_n4648_24[1]),.dinb(w_n2864_0[0]),.dout(n5001),.clk(gclk));
	jand g4360(.dina(n5001),.dinb(n5000),.dout(result117),.clk(gclk));
	jor g4361(.dina(w_address1_24[0]),.dinb(w_n2884_0[0]),.dout(n5003),.clk(gclk));
	jor g4362(.dina(w_n4648_24[0]),.dinb(w_n2845_0[0]),.dout(n5004),.clk(gclk));
	jand g4363(.dina(n5004),.dinb(n5003),.dout(result118),.clk(gclk));
	jor g4364(.dina(w_address1_23[2]),.dinb(w_n2882_0[0]),.dout(n5006),.clk(gclk));
	jor g4365(.dina(w_n4648_23[2]),.dinb(w_n2856_0[0]),.dout(n5007),.clk(gclk));
	jand g4366(.dina(n5007),.dinb(n5006),.dout(result119),.clk(gclk));
	jor g4367(.dina(w_address1_23[1]),.dinb(w_n4460_0[0]),.dout(n5009),.clk(gclk));
	jor g4368(.dina(w_n4648_23[1]),.dinb(w_n4419_0[0]),.dout(n5010),.clk(gclk));
	jand g4369(.dina(n5010),.dinb(n5009),.dout(result120),.clk(gclk));
	jor g4370(.dina(w_address1_23[0]),.dinb(w_n4463_0[0]),.dout(n5012),.clk(gclk));
	jor g4371(.dina(w_n4648_23[0]),.dinb(w_n4449_0[0]),.dout(n5013),.clk(gclk));
	jand g4372(.dina(n5013),.dinb(n5012),.dout(result121),.clk(gclk));
	jor g4373(.dina(w_address1_22[2]),.dinb(w_n4458_0[0]),.dout(n5015),.clk(gclk));
	jor g4374(.dina(w_n4648_22[2]),.dinb(w_n4436_0[0]),.dout(n5016),.clk(gclk));
	jand g4375(.dina(n5016),.dinb(n5015),.dout(result122),.clk(gclk));
	jor g4376(.dina(w_address1_22[1]),.dinb(w_n4456_0[0]),.dout(n5018),.clk(gclk));
	jor g4377(.dina(w_n4648_22[1]),.dinb(w_n4431_0[0]),.dout(n5019),.clk(gclk));
	jand g4378(.dina(n5019),.dinb(n5018),.dout(result123),.clk(gclk));
	jor g4379(.dina(w_address1_22[0]),.dinb(w_n2826_0[0]),.dout(n5021),.clk(gclk));
	jor g4380(.dina(w_n4648_22[0]),.dinb(w_n2839_0[0]),.dout(n5022),.clk(gclk));
	jand g4381(.dina(n5022),.dinb(n5021),.dout(result124),.clk(gclk));
	jor g4382(.dina(w_address1_21[2]),.dinb(w_n2831_0[0]),.dout(n5024),.clk(gclk));
	jor g4383(.dina(w_n4648_21[2]),.dinb(w_n2819_0[0]),.dout(n5025),.clk(gclk));
	jand g4384(.dina(n5025),.dinb(n5024),.dout(result125),.clk(gclk));
	jor g4385(.dina(w_address1_21[1]),.dinb(w_n2835_0[0]),.dout(n5027),.clk(gclk));
	jor g4386(.dina(w_n4648_21[1]),.dinb(w_n2811_0[0]),.dout(n5028),.clk(gclk));
	jand g4387(.dina(n5028),.dinb(n5027),.dout(result126),.clk(gclk));
	jand g4388(.dina(w_n2643_0[1]),.dinb(w_n2641_0[0]),.dout(w_dff_A_4jf92R4g9_2),.clk(gclk));
	jor g4389(.dina(w_address1_21[0]),.dinb(w_n1562_21[1]),.dout(n5031),.clk(gclk));
	jor g4390(.dina(w_n4648_21[0]),.dinb(w_n2808_21[1]),.dout(n5032),.clk(gclk));
	jand g4391(.dina(n5032),.dinb(n5031),.dout(address0),.clk(gclk));
	jspl3 jspl3_w_in00_0(.douta(w_in00_0[0]),.doutb(w_in00_0[1]),.doutc(w_in00_0[2]),.din(in00));
	jspl3 jspl3_w_in01_0(.douta(w_in01_0[0]),.doutb(w_in01_0[1]),.doutc(w_in01_0[2]),.din(in01));
	jspl jspl_w_in01_1(.douta(w_in01_1[0]),.doutb(w_in01_1[1]),.din(w_in01_0[0]));
	jspl3 jspl3_w_in02_0(.douta(w_in02_0[0]),.doutb(w_in02_0[1]),.doutc(w_in02_0[2]),.din(in02));
	jspl jspl_w_in02_1(.douta(w_in02_1[0]),.doutb(w_in02_1[1]),.din(w_in02_0[0]));
	jspl3 jspl3_w_in03_0(.douta(w_in03_0[0]),.doutb(w_in03_0[1]),.doutc(w_in03_0[2]),.din(in03));
	jspl jspl_w_in04_0(.douta(w_in04_0[0]),.doutb(w_in04_0[1]),.din(in04));
	jspl jspl_w_in05_0(.douta(w_in05_0[0]),.doutb(w_in05_0[1]),.din(in05));
	jspl jspl_w_in06_0(.douta(w_in06_0[0]),.doutb(w_in06_0[1]),.din(in06));
	jspl jspl_w_in07_0(.douta(w_in07_0[0]),.doutb(w_in07_0[1]),.din(in07));
	jspl jspl_w_in08_0(.douta(w_in08_0[0]),.doutb(w_in08_0[1]),.din(in08));
	jspl jspl_w_in09_0(.douta(w_in09_0[0]),.doutb(w_in09_0[1]),.din(in09));
	jspl jspl_w_in010_0(.douta(w_in010_0[0]),.doutb(w_in010_0[1]),.din(in010));
	jspl jspl_w_in011_0(.douta(w_in011_0[0]),.doutb(w_in011_0[1]),.din(in011));
	jspl jspl_w_in012_0(.douta(w_in012_0[0]),.doutb(w_in012_0[1]),.din(in012));
	jspl jspl_w_in013_0(.douta(w_in013_0[0]),.doutb(w_in013_0[1]),.din(in013));
	jspl jspl_w_in014_0(.douta(w_in014_0[0]),.doutb(w_in014_0[1]),.din(in014));
	jspl jspl_w_in015_0(.douta(w_in015_0[0]),.doutb(w_in015_0[1]),.din(in015));
	jspl jspl_w_in016_0(.douta(w_in016_0[0]),.doutb(w_in016_0[1]),.din(in016));
	jspl jspl_w_in017_0(.douta(w_in017_0[0]),.doutb(w_in017_0[1]),.din(in017));
	jspl jspl_w_in018_0(.douta(w_in018_0[0]),.doutb(w_in018_0[1]),.din(in018));
	jspl jspl_w_in019_0(.douta(w_in019_0[0]),.doutb(w_in019_0[1]),.din(in019));
	jspl jspl_w_in020_0(.douta(w_in020_0[0]),.doutb(w_in020_0[1]),.din(in020));
	jspl jspl_w_in021_0(.douta(w_in021_0[0]),.doutb(w_in021_0[1]),.din(in021));
	jspl jspl_w_in022_0(.douta(w_in022_0[0]),.doutb(w_in022_0[1]),.din(in022));
	jspl jspl_w_in023_0(.douta(w_in023_0[0]),.doutb(w_in023_0[1]),.din(in023));
	jspl jspl_w_in024_0(.douta(w_in024_0[0]),.doutb(w_in024_0[1]),.din(in024));
	jspl jspl_w_in025_0(.douta(w_in025_0[0]),.doutb(w_in025_0[1]),.din(in025));
	jspl jspl_w_in026_0(.douta(w_in026_0[0]),.doutb(w_in026_0[1]),.din(in026));
	jspl jspl_w_in027_0(.douta(w_in027_0[0]),.doutb(w_in027_0[1]),.din(in027));
	jspl jspl_w_in028_0(.douta(w_in028_0[0]),.doutb(w_in028_0[1]),.din(in028));
	jspl jspl_w_in029_0(.douta(w_in029_0[0]),.doutb(w_in029_0[1]),.din(in029));
	jspl jspl_w_in030_0(.douta(w_in030_0[0]),.doutb(w_in030_0[1]),.din(in030));
	jspl jspl_w_in031_0(.douta(w_in031_0[0]),.doutb(w_in031_0[1]),.din(in031));
	jspl jspl_w_in032_0(.douta(w_in032_0[0]),.doutb(w_in032_0[1]),.din(in032));
	jspl jspl_w_in033_0(.douta(w_in033_0[0]),.doutb(w_in033_0[1]),.din(in033));
	jspl jspl_w_in034_0(.douta(w_in034_0[0]),.doutb(w_in034_0[1]),.din(in034));
	jspl jspl_w_in035_0(.douta(w_in035_0[0]),.doutb(w_in035_0[1]),.din(in035));
	jspl jspl_w_in036_0(.douta(w_in036_0[0]),.doutb(w_in036_0[1]),.din(in036));
	jspl jspl_w_in037_0(.douta(w_in037_0[0]),.doutb(w_in037_0[1]),.din(in037));
	jspl jspl_w_in038_0(.douta(w_in038_0[0]),.doutb(w_in038_0[1]),.din(in038));
	jspl jspl_w_in039_0(.douta(w_in039_0[0]),.doutb(w_in039_0[1]),.din(in039));
	jspl jspl_w_in040_0(.douta(w_in040_0[0]),.doutb(w_in040_0[1]),.din(in040));
	jspl jspl_w_in041_0(.douta(w_in041_0[0]),.doutb(w_in041_0[1]),.din(in041));
	jspl jspl_w_in042_0(.douta(w_in042_0[0]),.doutb(w_in042_0[1]),.din(in042));
	jspl jspl_w_in044_0(.douta(w_in044_0[0]),.doutb(w_in044_0[1]),.din(in044));
	jspl jspl_w_in045_0(.douta(w_in045_0[0]),.doutb(w_in045_0[1]),.din(in045));
	jspl jspl_w_in046_0(.douta(w_in046_0[0]),.doutb(w_in046_0[1]),.din(in046));
	jspl jspl_w_in047_0(.douta(w_in047_0[0]),.doutb(w_in047_0[1]),.din(in047));
	jspl jspl_w_in048_0(.douta(w_in048_0[0]),.doutb(w_in048_0[1]),.din(in048));
	jspl jspl_w_in049_0(.douta(w_in049_0[0]),.doutb(w_in049_0[1]),.din(in049));
	jspl jspl_w_in050_0(.douta(w_in050_0[0]),.doutb(w_in050_0[1]),.din(in050));
	jspl jspl_w_in051_0(.douta(w_in051_0[0]),.doutb(w_in051_0[1]),.din(in051));
	jspl jspl_w_in052_0(.douta(w_in052_0[0]),.doutb(w_in052_0[1]),.din(in052));
	jspl jspl_w_in053_0(.douta(w_in053_0[0]),.doutb(w_in053_0[1]),.din(in053));
	jspl jspl_w_in054_0(.douta(w_in054_0[0]),.doutb(w_in054_0[1]),.din(in054));
	jspl jspl_w_in055_0(.douta(w_in055_0[0]),.doutb(w_in055_0[1]),.din(in055));
	jspl jspl_w_in056_0(.douta(w_in056_0[0]),.doutb(w_in056_0[1]),.din(in056));
	jspl jspl_w_in057_0(.douta(w_in057_0[0]),.doutb(w_in057_0[1]),.din(in057));
	jspl jspl_w_in058_0(.douta(w_in058_0[0]),.doutb(w_in058_0[1]),.din(in058));
	jspl jspl_w_in059_0(.douta(w_in059_0[0]),.doutb(w_in059_0[1]),.din(in059));
	jspl jspl_w_in060_0(.douta(w_in060_0[0]),.doutb(w_in060_0[1]),.din(in060));
	jspl jspl_w_in061_0(.douta(w_in061_0[0]),.doutb(w_in061_0[1]),.din(in061));
	jspl jspl_w_in062_0(.douta(w_in062_0[0]),.doutb(w_in062_0[1]),.din(in062));
	jspl jspl_w_in063_0(.douta(w_in063_0[0]),.doutb(w_in063_0[1]),.din(in063));
	jspl jspl_w_in064_0(.douta(w_in064_0[0]),.doutb(w_in064_0[1]),.din(in064));
	jspl jspl_w_in065_0(.douta(w_in065_0[0]),.doutb(w_in065_0[1]),.din(in065));
	jspl jspl_w_in066_0(.douta(w_in066_0[0]),.doutb(w_in066_0[1]),.din(in066));
	jspl jspl_w_in067_0(.douta(w_in067_0[0]),.doutb(w_in067_0[1]),.din(in067));
	jspl jspl_w_in068_0(.douta(w_in068_0[0]),.doutb(w_in068_0[1]),.din(in068));
	jspl jspl_w_in069_0(.douta(w_in069_0[0]),.doutb(w_in069_0[1]),.din(in069));
	jspl jspl_w_in070_0(.douta(w_in070_0[0]),.doutb(w_in070_0[1]),.din(in070));
	jspl jspl_w_in071_0(.douta(w_in071_0[0]),.doutb(w_in071_0[1]),.din(in071));
	jspl jspl_w_in072_0(.douta(w_in072_0[0]),.doutb(w_in072_0[1]),.din(in072));
	jspl jspl_w_in073_0(.douta(w_in073_0[0]),.doutb(w_in073_0[1]),.din(in073));
	jspl jspl_w_in074_0(.douta(w_in074_0[0]),.doutb(w_in074_0[1]),.din(in074));
	jspl jspl_w_in075_0(.douta(w_in075_0[0]),.doutb(w_in075_0[1]),.din(in075));
	jspl jspl_w_in076_0(.douta(w_in076_0[0]),.doutb(w_in076_0[1]),.din(in076));
	jspl jspl_w_in077_0(.douta(w_in077_0[0]),.doutb(w_in077_0[1]),.din(in077));
	jspl jspl_w_in078_0(.douta(w_in078_0[0]),.doutb(w_in078_0[1]),.din(in078));
	jspl jspl_w_in079_0(.douta(w_in079_0[0]),.doutb(w_in079_0[1]),.din(in079));
	jspl jspl_w_in080_0(.douta(w_in080_0[0]),.doutb(w_in080_0[1]),.din(in080));
	jspl jspl_w_in081_0(.douta(w_in081_0[0]),.doutb(w_in081_0[1]),.din(in081));
	jspl jspl_w_in082_0(.douta(w_in082_0[0]),.doutb(w_in082_0[1]),.din(in082));
	jspl jspl_w_in083_0(.douta(w_in083_0[0]),.doutb(w_in083_0[1]),.din(in083));
	jspl jspl_w_in084_0(.douta(w_in084_0[0]),.doutb(w_in084_0[1]),.din(in084));
	jspl jspl_w_in085_0(.douta(w_in085_0[0]),.doutb(w_in085_0[1]),.din(in085));
	jspl jspl_w_in086_0(.douta(w_in086_0[0]),.doutb(w_in086_0[1]),.din(in086));
	jspl jspl_w_in087_0(.douta(w_in087_0[0]),.doutb(w_in087_0[1]),.din(in087));
	jspl jspl_w_in088_0(.douta(w_in088_0[0]),.doutb(w_in088_0[1]),.din(in088));
	jspl jspl_w_in089_0(.douta(w_in089_0[0]),.doutb(w_in089_0[1]),.din(in089));
	jspl jspl_w_in090_0(.douta(w_in090_0[0]),.doutb(w_in090_0[1]),.din(in090));
	jspl jspl_w_in091_0(.douta(w_in091_0[0]),.doutb(w_in091_0[1]),.din(in091));
	jspl jspl_w_in092_0(.douta(w_in092_0[0]),.doutb(w_in092_0[1]),.din(in092));
	jspl jspl_w_in093_0(.douta(w_in093_0[0]),.doutb(w_in093_0[1]),.din(in093));
	jspl jspl_w_in094_0(.douta(w_in094_0[0]),.doutb(w_in094_0[1]),.din(in094));
	jspl jspl_w_in095_0(.douta(w_in095_0[0]),.doutb(w_in095_0[1]),.din(in095));
	jspl jspl_w_in096_0(.douta(w_in096_0[0]),.doutb(w_in096_0[1]),.din(in096));
	jspl jspl_w_in097_0(.douta(w_in097_0[0]),.doutb(w_in097_0[1]),.din(in097));
	jspl jspl_w_in098_0(.douta(w_in098_0[0]),.doutb(w_in098_0[1]),.din(in098));
	jspl jspl_w_in099_0(.douta(w_in099_0[0]),.doutb(w_in099_0[1]),.din(in099));
	jspl jspl_w_in0100_0(.douta(w_in0100_0[0]),.doutb(w_in0100_0[1]),.din(in0100));
	jspl jspl_w_in0101_0(.douta(w_in0101_0[0]),.doutb(w_in0101_0[1]),.din(in0101));
	jspl jspl_w_in0102_0(.douta(w_in0102_0[0]),.doutb(w_in0102_0[1]),.din(in0102));
	jspl jspl_w_in0103_0(.douta(w_in0103_0[0]),.doutb(w_in0103_0[1]),.din(in0103));
	jspl jspl_w_in0104_0(.douta(w_in0104_0[0]),.doutb(w_in0104_0[1]),.din(in0104));
	jspl jspl_w_in0105_0(.douta(w_in0105_0[0]),.doutb(w_in0105_0[1]),.din(in0105));
	jspl jspl_w_in0106_0(.douta(w_in0106_0[0]),.doutb(w_in0106_0[1]),.din(in0106));
	jspl jspl_w_in0107_0(.douta(w_in0107_0[0]),.doutb(w_in0107_0[1]),.din(in0107));
	jspl jspl_w_in0108_0(.douta(w_in0108_0[0]),.doutb(w_in0108_0[1]),.din(in0108));
	jspl jspl_w_in0109_0(.douta(w_in0109_0[0]),.doutb(w_in0109_0[1]),.din(in0109));
	jspl jspl_w_in0110_0(.douta(w_in0110_0[0]),.doutb(w_in0110_0[1]),.din(in0110));
	jspl jspl_w_in0111_0(.douta(w_in0111_0[0]),.doutb(w_in0111_0[1]),.din(in0111));
	jspl jspl_w_in0112_0(.douta(w_in0112_0[0]),.doutb(w_in0112_0[1]),.din(in0112));
	jspl jspl_w_in0113_0(.douta(w_in0113_0[0]),.doutb(w_in0113_0[1]),.din(in0113));
	jspl jspl_w_in0114_0(.douta(w_in0114_0[0]),.doutb(w_in0114_0[1]),.din(in0114));
	jspl jspl_w_in0115_0(.douta(w_in0115_0[0]),.doutb(w_in0115_0[1]),.din(in0115));
	jspl jspl_w_in0116_0(.douta(w_in0116_0[0]),.doutb(w_in0116_0[1]),.din(in0116));
	jspl jspl_w_in0117_0(.douta(w_in0117_0[0]),.doutb(w_in0117_0[1]),.din(in0117));
	jspl jspl_w_in0118_0(.douta(w_in0118_0[0]),.doutb(w_in0118_0[1]),.din(in0118));
	jspl jspl_w_in0119_0(.douta(w_in0119_0[0]),.doutb(w_in0119_0[1]),.din(in0119));
	jspl jspl_w_in0120_0(.douta(w_in0120_0[0]),.doutb(w_in0120_0[1]),.din(in0120));
	jspl jspl_w_in0121_0(.douta(w_in0121_0[0]),.doutb(w_in0121_0[1]),.din(in0121));
	jspl jspl_w_in0122_0(.douta(w_in0122_0[0]),.doutb(w_in0122_0[1]),.din(in0122));
	jspl jspl_w_in0123_0(.douta(w_in0123_0[0]),.doutb(w_in0123_0[1]),.din(in0123));
	jspl jspl_w_in0124_0(.douta(w_in0124_0[0]),.doutb(w_in0124_0[1]),.din(in0124));
	jspl jspl_w_in0125_0(.douta(w_in0125_0[0]),.doutb(w_in0125_0[1]),.din(in0125));
	jspl jspl_w_in0126_0(.douta(w_in0126_0[0]),.doutb(w_in0126_0[1]),.din(in0126));
	jspl3 jspl3_w_in0127_0(.douta(w_in0127_0[0]),.doutb(w_in0127_0[1]),.doutc(w_in0127_0[2]),.din(in0127));
	jspl3 jspl3_w_in10_0(.douta(w_in10_0[0]),.doutb(w_in10_0[1]),.doutc(w_in10_0[2]),.din(in10));
	jspl3 jspl3_w_in11_0(.douta(w_in11_0[0]),.doutb(w_in11_0[1]),.doutc(w_in11_0[2]),.din(in11));
	jspl jspl_w_in11_1(.douta(w_in11_1[0]),.doutb(w_in11_1[1]),.din(w_in11_0[0]));
	jspl3 jspl3_w_in12_0(.douta(w_in12_0[0]),.doutb(w_in12_0[1]),.doutc(w_in12_0[2]),.din(in12));
	jspl3 jspl3_w_in13_0(.douta(w_in13_0[0]),.doutb(w_in13_0[1]),.doutc(w_in13_0[2]),.din(in13));
	jspl jspl_w_in14_0(.douta(w_in14_0[0]),.doutb(w_in14_0[1]),.din(in14));
	jspl jspl_w_in15_0(.douta(w_in15_0[0]),.doutb(w_in15_0[1]),.din(in15));
	jspl jspl_w_in16_0(.douta(w_in16_0[0]),.doutb(w_in16_0[1]),.din(in16));
	jspl jspl_w_in17_0(.douta(w_in17_0[0]),.doutb(w_in17_0[1]),.din(in17));
	jspl jspl_w_in18_0(.douta(w_in18_0[0]),.doutb(w_in18_0[1]),.din(in18));
	jspl jspl_w_in19_0(.douta(w_in19_0[0]),.doutb(w_in19_0[1]),.din(in19));
	jspl jspl_w_in110_0(.douta(w_in110_0[0]),.doutb(w_in110_0[1]),.din(in110));
	jspl jspl_w_in111_0(.douta(w_in111_0[0]),.doutb(w_in111_0[1]),.din(in111));
	jspl jspl_w_in112_0(.douta(w_in112_0[0]),.doutb(w_in112_0[1]),.din(in112));
	jspl jspl_w_in113_0(.douta(w_in113_0[0]),.doutb(w_in113_0[1]),.din(in113));
	jspl jspl_w_in114_0(.douta(w_in114_0[0]),.doutb(w_in114_0[1]),.din(in114));
	jspl jspl_w_in115_0(.douta(w_in115_0[0]),.doutb(w_in115_0[1]),.din(in115));
	jspl jspl_w_in116_0(.douta(w_in116_0[0]),.doutb(w_in116_0[1]),.din(in116));
	jspl jspl_w_in117_0(.douta(w_in117_0[0]),.doutb(w_in117_0[1]),.din(in117));
	jspl jspl_w_in118_0(.douta(w_in118_0[0]),.doutb(w_in118_0[1]),.din(in118));
	jspl jspl_w_in119_0(.douta(w_in119_0[0]),.doutb(w_in119_0[1]),.din(in119));
	jspl jspl_w_in120_0(.douta(w_in120_0[0]),.doutb(w_in120_0[1]),.din(in120));
	jspl jspl_w_in121_0(.douta(w_in121_0[0]),.doutb(w_in121_0[1]),.din(in121));
	jspl jspl_w_in122_0(.douta(w_in122_0[0]),.doutb(w_in122_0[1]),.din(in122));
	jspl jspl_w_in123_0(.douta(w_in123_0[0]),.doutb(w_in123_0[1]),.din(in123));
	jspl jspl_w_in124_0(.douta(w_in124_0[0]),.doutb(w_in124_0[1]),.din(in124));
	jspl jspl_w_in125_0(.douta(w_in125_0[0]),.doutb(w_in125_0[1]),.din(in125));
	jspl jspl_w_in126_0(.douta(w_in126_0[0]),.doutb(w_in126_0[1]),.din(in126));
	jspl jspl_w_in127_0(.douta(w_in127_0[0]),.doutb(w_in127_0[1]),.din(in127));
	jspl jspl_w_in128_0(.douta(w_in128_0[0]),.doutb(w_in128_0[1]),.din(in128));
	jspl jspl_w_in129_0(.douta(w_in129_0[0]),.doutb(w_in129_0[1]),.din(in129));
	jspl jspl_w_in130_0(.douta(w_in130_0[0]),.doutb(w_in130_0[1]),.din(in130));
	jspl jspl_w_in131_0(.douta(w_in131_0[0]),.doutb(w_in131_0[1]),.din(in131));
	jspl jspl_w_in132_0(.douta(w_in132_0[0]),.doutb(w_in132_0[1]),.din(in132));
	jspl jspl_w_in133_0(.douta(w_in133_0[0]),.doutb(w_in133_0[1]),.din(in133));
	jspl jspl_w_in134_0(.douta(w_in134_0[0]),.doutb(w_in134_0[1]),.din(in134));
	jspl jspl_w_in135_0(.douta(w_in135_0[0]),.doutb(w_in135_0[1]),.din(in135));
	jspl jspl_w_in136_0(.douta(w_in136_0[0]),.doutb(w_in136_0[1]),.din(in136));
	jspl jspl_w_in137_0(.douta(w_in137_0[0]),.doutb(w_in137_0[1]),.din(in137));
	jspl jspl_w_in138_0(.douta(w_in138_0[0]),.doutb(w_in138_0[1]),.din(in138));
	jspl jspl_w_in139_0(.douta(w_in139_0[0]),.doutb(w_in139_0[1]),.din(in139));
	jspl jspl_w_in140_0(.douta(w_in140_0[0]),.doutb(w_in140_0[1]),.din(in140));
	jspl jspl_w_in141_0(.douta(w_in141_0[0]),.doutb(w_in141_0[1]),.din(in141));
	jspl jspl_w_in142_0(.douta(w_in142_0[0]),.doutb(w_in142_0[1]),.din(in142));
	jspl3 jspl3_w_in143_0(.douta(w_in143_0[0]),.doutb(w_in143_0[1]),.doutc(w_in143_0[2]),.din(in143));
	jspl jspl_w_in144_0(.douta(w_in144_0[0]),.doutb(w_in144_0[1]),.din(in144));
	jspl jspl_w_in145_0(.douta(w_in145_0[0]),.doutb(w_in145_0[1]),.din(in145));
	jspl jspl_w_in146_0(.douta(w_in146_0[0]),.doutb(w_in146_0[1]),.din(in146));
	jspl jspl_w_in147_0(.douta(w_in147_0[0]),.doutb(w_in147_0[1]),.din(in147));
	jspl jspl_w_in148_0(.douta(w_in148_0[0]),.doutb(w_in148_0[1]),.din(in148));
	jspl jspl_w_in149_0(.douta(w_in149_0[0]),.doutb(w_in149_0[1]),.din(in149));
	jspl jspl_w_in150_0(.douta(w_in150_0[0]),.doutb(w_in150_0[1]),.din(in150));
	jspl jspl_w_in151_0(.douta(w_in151_0[0]),.doutb(w_in151_0[1]),.din(in151));
	jspl jspl_w_in152_0(.douta(w_in152_0[0]),.doutb(w_in152_0[1]),.din(in152));
	jspl jspl_w_in153_0(.douta(w_in153_0[0]),.doutb(w_in153_0[1]),.din(in153));
	jspl jspl_w_in154_0(.douta(w_in154_0[0]),.doutb(w_in154_0[1]),.din(in154));
	jspl jspl_w_in155_0(.douta(w_in155_0[0]),.doutb(w_in155_0[1]),.din(in155));
	jspl jspl_w_in156_0(.douta(w_in156_0[0]),.doutb(w_in156_0[1]),.din(in156));
	jspl jspl_w_in157_0(.douta(w_in157_0[0]),.doutb(w_in157_0[1]),.din(in157));
	jspl jspl_w_in158_0(.douta(w_in158_0[0]),.doutb(w_in158_0[1]),.din(in158));
	jspl jspl_w_in159_0(.douta(w_in159_0[0]),.doutb(w_in159_0[1]),.din(in159));
	jspl jspl_w_in160_0(.douta(w_in160_0[0]),.doutb(w_in160_0[1]),.din(in160));
	jspl jspl_w_in161_0(.douta(w_in161_0[0]),.doutb(w_in161_0[1]),.din(in161));
	jspl jspl_w_in162_0(.douta(w_in162_0[0]),.doutb(w_in162_0[1]),.din(in162));
	jspl jspl_w_in163_0(.douta(w_in163_0[0]),.doutb(w_in163_0[1]),.din(in163));
	jspl jspl_w_in164_0(.douta(w_in164_0[0]),.doutb(w_in164_0[1]),.din(in164));
	jspl jspl_w_in165_0(.douta(w_in165_0[0]),.doutb(w_in165_0[1]),.din(in165));
	jspl jspl_w_in166_0(.douta(w_in166_0[0]),.doutb(w_in166_0[1]),.din(in166));
	jspl jspl_w_in167_0(.douta(w_in167_0[0]),.doutb(w_in167_0[1]),.din(in167));
	jspl jspl_w_in168_0(.douta(w_in168_0[0]),.doutb(w_in168_0[1]),.din(in168));
	jspl jspl_w_in169_0(.douta(w_in169_0[0]),.doutb(w_in169_0[1]),.din(in169));
	jspl jspl_w_in170_0(.douta(w_in170_0[0]),.doutb(w_in170_0[1]),.din(in170));
	jspl jspl_w_in171_0(.douta(w_in171_0[0]),.doutb(w_in171_0[1]),.din(in171));
	jspl jspl_w_in172_0(.douta(w_in172_0[0]),.doutb(w_in172_0[1]),.din(in172));
	jspl jspl_w_in173_0(.douta(w_in173_0[0]),.doutb(w_in173_0[1]),.din(in173));
	jspl jspl_w_in174_0(.douta(w_in174_0[0]),.doutb(w_in174_0[1]),.din(in174));
	jspl jspl_w_in175_0(.douta(w_in175_0[0]),.doutb(w_in175_0[1]),.din(in175));
	jspl jspl_w_in176_0(.douta(w_in176_0[0]),.doutb(w_in176_0[1]),.din(in176));
	jspl jspl_w_in177_0(.douta(w_in177_0[0]),.doutb(w_in177_0[1]),.din(in177));
	jspl jspl_w_in178_0(.douta(w_in178_0[0]),.doutb(w_in178_0[1]),.din(in178));
	jspl jspl_w_in179_0(.douta(w_in179_0[0]),.doutb(w_in179_0[1]),.din(in179));
	jspl jspl_w_in180_0(.douta(w_in180_0[0]),.doutb(w_in180_0[1]),.din(in180));
	jspl jspl_w_in181_0(.douta(w_in181_0[0]),.doutb(w_in181_0[1]),.din(in181));
	jspl jspl_w_in182_0(.douta(w_in182_0[0]),.doutb(w_in182_0[1]),.din(in182));
	jspl jspl_w_in183_0(.douta(w_in183_0[0]),.doutb(w_in183_0[1]),.din(in183));
	jspl jspl_w_in184_0(.douta(w_in184_0[0]),.doutb(w_in184_0[1]),.din(in184));
	jspl jspl_w_in185_0(.douta(w_in185_0[0]),.doutb(w_in185_0[1]),.din(in185));
	jspl jspl_w_in186_0(.douta(w_in186_0[0]),.doutb(w_in186_0[1]),.din(in186));
	jspl jspl_w_in187_0(.douta(w_in187_0[0]),.doutb(w_in187_0[1]),.din(in187));
	jspl jspl_w_in188_0(.douta(w_in188_0[0]),.doutb(w_in188_0[1]),.din(in188));
	jspl jspl_w_in189_0(.douta(w_in189_0[0]),.doutb(w_in189_0[1]),.din(in189));
	jspl jspl_w_in190_0(.douta(w_in190_0[0]),.doutb(w_in190_0[1]),.din(in190));
	jspl jspl_w_in191_0(.douta(w_in191_0[0]),.doutb(w_in191_0[1]),.din(in191));
	jspl jspl_w_in192_0(.douta(w_in192_0[0]),.doutb(w_in192_0[1]),.din(in192));
	jspl jspl_w_in193_0(.douta(w_in193_0[0]),.doutb(w_in193_0[1]),.din(in193));
	jspl jspl_w_in194_0(.douta(w_in194_0[0]),.doutb(w_in194_0[1]),.din(in194));
	jspl jspl_w_in195_0(.douta(w_in195_0[0]),.doutb(w_in195_0[1]),.din(in195));
	jspl jspl_w_in196_0(.douta(w_in196_0[0]),.doutb(w_in196_0[1]),.din(in196));
	jspl jspl_w_in197_0(.douta(w_in197_0[0]),.doutb(w_in197_0[1]),.din(in197));
	jspl jspl_w_in198_0(.douta(w_in198_0[0]),.doutb(w_in198_0[1]),.din(in198));
	jspl jspl_w_in199_0(.douta(w_in199_0[0]),.doutb(w_in199_0[1]),.din(in199));
	jspl jspl_w_in1100_0(.douta(w_in1100_0[0]),.doutb(w_in1100_0[1]),.din(in1100));
	jspl jspl_w_in1101_0(.douta(w_in1101_0[0]),.doutb(w_in1101_0[1]),.din(in1101));
	jspl jspl_w_in1102_0(.douta(w_in1102_0[0]),.doutb(w_in1102_0[1]),.din(in1102));
	jspl jspl_w_in1103_0(.douta(w_in1103_0[0]),.doutb(w_in1103_0[1]),.din(in1103));
	jspl jspl_w_in1104_0(.douta(w_in1104_0[0]),.doutb(w_in1104_0[1]),.din(in1104));
	jspl jspl_w_in1105_0(.douta(w_in1105_0[0]),.doutb(w_in1105_0[1]),.din(in1105));
	jspl jspl_w_in1106_0(.douta(w_in1106_0[0]),.doutb(w_in1106_0[1]),.din(in1106));
	jspl jspl_w_in1107_0(.douta(w_in1107_0[0]),.doutb(w_in1107_0[1]),.din(in1107));
	jspl jspl_w_in1108_0(.douta(w_in1108_0[0]),.doutb(w_in1108_0[1]),.din(in1108));
	jspl jspl_w_in1109_0(.douta(w_in1109_0[0]),.doutb(w_in1109_0[1]),.din(in1109));
	jspl jspl_w_in1110_0(.douta(w_in1110_0[0]),.doutb(w_in1110_0[1]),.din(in1110));
	jspl jspl_w_in1111_0(.douta(w_in1111_0[0]),.doutb(w_in1111_0[1]),.din(in1111));
	jspl jspl_w_in1112_0(.douta(w_in1112_0[0]),.doutb(w_in1112_0[1]),.din(in1112));
	jspl jspl_w_in1113_0(.douta(w_in1113_0[0]),.doutb(w_in1113_0[1]),.din(in1113));
	jspl jspl_w_in1114_0(.douta(w_in1114_0[0]),.doutb(w_in1114_0[1]),.din(in1114));
	jspl jspl_w_in1115_0(.douta(w_in1115_0[0]),.doutb(w_in1115_0[1]),.din(in1115));
	jspl jspl_w_in1116_0(.douta(w_in1116_0[0]),.doutb(w_in1116_0[1]),.din(in1116));
	jspl jspl_w_in1117_0(.douta(w_in1117_0[0]),.doutb(w_in1117_0[1]),.din(in1117));
	jspl jspl_w_in1118_0(.douta(w_in1118_0[0]),.doutb(w_in1118_0[1]),.din(in1118));
	jspl jspl_w_in1119_0(.douta(w_in1119_0[0]),.doutb(w_in1119_0[1]),.din(in1119));
	jspl jspl_w_in1120_0(.douta(w_in1120_0[0]),.doutb(w_in1120_0[1]),.din(in1120));
	jspl jspl_w_in1121_0(.douta(w_in1121_0[0]),.doutb(w_in1121_0[1]),.din(in1121));
	jspl jspl_w_in1122_0(.douta(w_in1122_0[0]),.doutb(w_in1122_0[1]),.din(in1122));
	jspl jspl_w_in1123_0(.douta(w_in1123_0[0]),.doutb(w_in1123_0[1]),.din(in1123));
	jspl jspl_w_in1124_0(.douta(w_in1124_0[0]),.doutb(w_in1124_0[1]),.din(in1124));
	jspl jspl_w_in1125_0(.douta(w_in1125_0[0]),.doutb(w_in1125_0[1]),.din(in1125));
	jspl jspl_w_in1126_0(.douta(w_in1126_0[0]),.doutb(w_in1126_0[1]),.din(in1126));
	jspl3 jspl3_w_in1127_0(.douta(w_in1127_0[0]),.doutb(w_in1127_0[1]),.doutc(w_in1127_0[2]),.din(in1127));
	jspl3 jspl3_w_in20_0(.douta(w_in20_0[0]),.doutb(w_in20_0[1]),.doutc(w_in20_0[2]),.din(in20));
	jspl3 jspl3_w_in21_0(.douta(w_in21_0[0]),.doutb(w_in21_0[1]),.doutc(w_in21_0[2]),.din(in21));
	jspl jspl_w_in21_1(.douta(w_in21_1[0]),.doutb(w_in21_1[1]),.din(w_in21_0[0]));
	jspl3 jspl3_w_in22_0(.douta(w_in22_0[0]),.doutb(w_in22_0[1]),.doutc(w_in22_0[2]),.din(in22));
	jspl jspl_w_in23_0(.douta(w_in23_0[0]),.doutb(w_in23_0[1]),.din(in23));
	jspl jspl_w_in24_0(.douta(w_in24_0[0]),.doutb(w_in24_0[1]),.din(in24));
	jspl jspl_w_in25_0(.douta(w_in25_0[0]),.doutb(w_in25_0[1]),.din(in25));
	jspl jspl_w_in26_0(.douta(w_in26_0[0]),.doutb(w_in26_0[1]),.din(in26));
	jspl jspl_w_in27_0(.douta(w_in27_0[0]),.doutb(w_in27_0[1]),.din(in27));
	jspl jspl_w_in28_0(.douta(w_in28_0[0]),.doutb(w_in28_0[1]),.din(in28));
	jspl jspl_w_in29_0(.douta(w_in29_0[0]),.doutb(w_in29_0[1]),.din(in29));
	jspl jspl_w_in210_0(.douta(w_in210_0[0]),.doutb(w_in210_0[1]),.din(in210));
	jspl jspl_w_in211_0(.douta(w_in211_0[0]),.doutb(w_in211_0[1]),.din(in211));
	jspl jspl_w_in212_0(.douta(w_in212_0[0]),.doutb(w_in212_0[1]),.din(in212));
	jspl jspl_w_in213_0(.douta(w_in213_0[0]),.doutb(w_in213_0[1]),.din(in213));
	jspl jspl_w_in214_0(.douta(w_in214_0[0]),.doutb(w_in214_0[1]),.din(in214));
	jspl jspl_w_in215_0(.douta(w_in215_0[0]),.doutb(w_in215_0[1]),.din(in215));
	jspl jspl_w_in216_0(.douta(w_in216_0[0]),.doutb(w_in216_0[1]),.din(in216));
	jspl jspl_w_in217_0(.douta(w_in217_0[0]),.doutb(w_in217_0[1]),.din(in217));
	jspl jspl_w_in218_0(.douta(w_in218_0[0]),.doutb(w_in218_0[1]),.din(in218));
	jspl jspl_w_in219_0(.douta(w_in219_0[0]),.doutb(w_in219_0[1]),.din(in219));
	jspl jspl_w_in220_0(.douta(w_in220_0[0]),.doutb(w_in220_0[1]),.din(in220));
	jspl jspl_w_in221_0(.douta(w_in221_0[0]),.doutb(w_in221_0[1]),.din(in221));
	jspl jspl_w_in222_0(.douta(w_in222_0[0]),.doutb(w_in222_0[1]),.din(in222));
	jspl jspl_w_in223_0(.douta(w_in223_0[0]),.doutb(w_in223_0[1]),.din(in223));
	jspl jspl_w_in224_0(.douta(w_in224_0[0]),.doutb(w_in224_0[1]),.din(in224));
	jspl jspl_w_in225_0(.douta(w_in225_0[0]),.doutb(w_in225_0[1]),.din(in225));
	jspl jspl_w_in226_0(.douta(w_in226_0[0]),.doutb(w_in226_0[1]),.din(in226));
	jspl jspl_w_in227_0(.douta(w_in227_0[0]),.doutb(w_in227_0[1]),.din(in227));
	jspl jspl_w_in228_0(.douta(w_in228_0[0]),.doutb(w_in228_0[1]),.din(in228));
	jspl jspl_w_in229_0(.douta(w_in229_0[0]),.doutb(w_in229_0[1]),.din(in229));
	jspl jspl_w_in230_0(.douta(w_in230_0[0]),.doutb(w_in230_0[1]),.din(in230));
	jspl jspl_w_in231_0(.douta(w_in231_0[0]),.doutb(w_in231_0[1]),.din(in231));
	jspl jspl_w_in232_0(.douta(w_in232_0[0]),.doutb(w_in232_0[1]),.din(in232));
	jspl jspl_w_in233_0(.douta(w_in233_0[0]),.doutb(w_in233_0[1]),.din(in233));
	jspl jspl_w_in234_0(.douta(w_in234_0[0]),.doutb(w_in234_0[1]),.din(in234));
	jspl jspl_w_in235_0(.douta(w_in235_0[0]),.doutb(w_in235_0[1]),.din(in235));
	jspl jspl_w_in236_0(.douta(w_in236_0[0]),.doutb(w_in236_0[1]),.din(in236));
	jspl jspl_w_in237_0(.douta(w_in237_0[0]),.doutb(w_in237_0[1]),.din(in237));
	jspl jspl_w_in238_0(.douta(w_in238_0[0]),.doutb(w_in238_0[1]),.din(in238));
	jspl jspl_w_in239_0(.douta(w_in239_0[0]),.doutb(w_in239_0[1]),.din(in239));
	jspl jspl_w_in240_0(.douta(w_in240_0[0]),.doutb(w_in240_0[1]),.din(in240));
	jspl jspl_w_in241_0(.douta(w_in241_0[0]),.doutb(w_in241_0[1]),.din(in241));
	jspl jspl_w_in242_0(.douta(w_in242_0[0]),.doutb(w_in242_0[1]),.din(in242));
	jspl jspl_w_in243_0(.douta(w_in243_0[0]),.doutb(w_in243_0[1]),.din(in243));
	jspl jspl_w_in244_0(.douta(w_in244_0[0]),.doutb(w_in244_0[1]),.din(in244));
	jspl jspl_w_in245_0(.douta(w_in245_0[0]),.doutb(w_in245_0[1]),.din(in245));
	jspl jspl_w_in246_0(.douta(w_in246_0[0]),.doutb(w_in246_0[1]),.din(in246));
	jspl jspl_w_in247_0(.douta(w_in247_0[0]),.doutb(w_in247_0[1]),.din(in247));
	jspl jspl_w_in248_0(.douta(w_in248_0[0]),.doutb(w_in248_0[1]),.din(in248));
	jspl jspl_w_in249_0(.douta(w_in249_0[0]),.doutb(w_in249_0[1]),.din(in249));
	jspl jspl_w_in250_0(.douta(w_in250_0[0]),.doutb(w_in250_0[1]),.din(in250));
	jspl jspl_w_in251_0(.douta(w_in251_0[0]),.doutb(w_in251_0[1]),.din(in251));
	jspl jspl_w_in252_0(.douta(w_in252_0[0]),.doutb(w_in252_0[1]),.din(in252));
	jspl jspl_w_in253_0(.douta(w_in253_0[0]),.doutb(w_in253_0[1]),.din(in253));
	jspl jspl_w_in254_0(.douta(w_in254_0[0]),.doutb(w_in254_0[1]),.din(in254));
	jspl jspl_w_in255_0(.douta(w_in255_0[0]),.doutb(w_in255_0[1]),.din(in255));
	jspl jspl_w_in256_0(.douta(w_in256_0[0]),.doutb(w_in256_0[1]),.din(in256));
	jspl jspl_w_in257_0(.douta(w_in257_0[0]),.doutb(w_in257_0[1]),.din(in257));
	jspl jspl_w_in258_0(.douta(w_in258_0[0]),.doutb(w_in258_0[1]),.din(in258));
	jspl jspl_w_in259_0(.douta(w_in259_0[0]),.doutb(w_in259_0[1]),.din(in259));
	jspl jspl_w_in260_0(.douta(w_in260_0[0]),.doutb(w_in260_0[1]),.din(in260));
	jspl jspl_w_in261_0(.douta(w_in261_0[0]),.doutb(w_in261_0[1]),.din(in261));
	jspl jspl_w_in262_0(.douta(w_in262_0[0]),.doutb(w_in262_0[1]),.din(in262));
	jspl jspl_w_in263_0(.douta(w_in263_0[0]),.doutb(w_in263_0[1]),.din(in263));
	jspl jspl_w_in264_0(.douta(w_in264_0[0]),.doutb(w_in264_0[1]),.din(in264));
	jspl jspl_w_in265_0(.douta(w_in265_0[0]),.doutb(w_in265_0[1]),.din(in265));
	jspl jspl_w_in266_0(.douta(w_in266_0[0]),.doutb(w_in266_0[1]),.din(in266));
	jspl jspl_w_in267_0(.douta(w_in267_0[0]),.doutb(w_in267_0[1]),.din(in267));
	jspl jspl_w_in268_0(.douta(w_in268_0[0]),.doutb(w_in268_0[1]),.din(in268));
	jspl jspl_w_in269_0(.douta(w_in269_0[0]),.doutb(w_in269_0[1]),.din(in269));
	jspl jspl_w_in270_0(.douta(w_in270_0[0]),.doutb(w_in270_0[1]),.din(in270));
	jspl jspl_w_in271_0(.douta(w_in271_0[0]),.doutb(w_in271_0[1]),.din(in271));
	jspl jspl_w_in272_0(.douta(w_in272_0[0]),.doutb(w_in272_0[1]),.din(in272));
	jspl jspl_w_in273_0(.douta(w_in273_0[0]),.doutb(w_in273_0[1]),.din(in273));
	jspl jspl_w_in274_0(.douta(w_in274_0[0]),.doutb(w_in274_0[1]),.din(in274));
	jspl jspl_w_in275_0(.douta(w_in275_0[0]),.doutb(w_in275_0[1]),.din(in275));
	jspl jspl_w_in276_0(.douta(w_in276_0[0]),.doutb(w_in276_0[1]),.din(in276));
	jspl jspl_w_in277_0(.douta(w_in277_0[0]),.doutb(w_in277_0[1]),.din(in277));
	jspl jspl_w_in278_0(.douta(w_in278_0[0]),.doutb(w_in278_0[1]),.din(in278));
	jspl jspl_w_in279_0(.douta(w_in279_0[0]),.doutb(w_in279_0[1]),.din(in279));
	jspl jspl_w_in280_0(.douta(w_in280_0[0]),.doutb(w_in280_0[1]),.din(in280));
	jspl jspl_w_in281_0(.douta(w_in281_0[0]),.doutb(w_in281_0[1]),.din(in281));
	jspl jspl_w_in282_0(.douta(w_in282_0[0]),.doutb(w_in282_0[1]),.din(in282));
	jspl jspl_w_in283_0(.douta(w_in283_0[0]),.doutb(w_in283_0[1]),.din(in283));
	jspl jspl_w_in284_0(.douta(w_in284_0[0]),.doutb(w_in284_0[1]),.din(in284));
	jspl jspl_w_in285_0(.douta(w_in285_0[0]),.doutb(w_in285_0[1]),.din(in285));
	jspl jspl_w_in286_0(.douta(w_in286_0[0]),.doutb(w_in286_0[1]),.din(in286));
	jspl jspl_w_in287_0(.douta(w_in287_0[0]),.doutb(w_in287_0[1]),.din(in287));
	jspl jspl_w_in288_0(.douta(w_in288_0[0]),.doutb(w_in288_0[1]),.din(in288));
	jspl jspl_w_in289_0(.douta(w_in289_0[0]),.doutb(w_in289_0[1]),.din(in289));
	jspl jspl_w_in290_0(.douta(w_in290_0[0]),.doutb(w_in290_0[1]),.din(in290));
	jspl jspl_w_in291_0(.douta(w_in291_0[0]),.doutb(w_in291_0[1]),.din(in291));
	jspl jspl_w_in292_0(.douta(w_in292_0[0]),.doutb(w_in292_0[1]),.din(in292));
	jspl jspl_w_in293_0(.douta(w_in293_0[0]),.doutb(w_in293_0[1]),.din(in293));
	jspl jspl_w_in294_0(.douta(w_in294_0[0]),.doutb(w_in294_0[1]),.din(in294));
	jspl jspl_w_in295_0(.douta(w_in295_0[0]),.doutb(w_in295_0[1]),.din(in295));
	jspl jspl_w_in296_0(.douta(w_in296_0[0]),.doutb(w_in296_0[1]),.din(in296));
	jspl jspl_w_in297_0(.douta(w_in297_0[0]),.doutb(w_in297_0[1]),.din(in297));
	jspl jspl_w_in298_0(.douta(w_in298_0[0]),.doutb(w_in298_0[1]),.din(in298));
	jspl jspl_w_in299_0(.douta(w_in299_0[0]),.doutb(w_in299_0[1]),.din(in299));
	jspl jspl_w_in2100_0(.douta(w_in2100_0[0]),.doutb(w_in2100_0[1]),.din(in2100));
	jspl jspl_w_in2101_0(.douta(w_in2101_0[0]),.doutb(w_in2101_0[1]),.din(in2101));
	jspl jspl_w_in2102_0(.douta(w_in2102_0[0]),.doutb(w_in2102_0[1]),.din(in2102));
	jspl jspl_w_in2103_0(.douta(w_in2103_0[0]),.doutb(w_in2103_0[1]),.din(in2103));
	jspl jspl_w_in2104_0(.douta(w_in2104_0[0]),.doutb(w_in2104_0[1]),.din(in2104));
	jspl jspl_w_in2105_0(.douta(w_in2105_0[0]),.doutb(w_in2105_0[1]),.din(in2105));
	jspl jspl_w_in2106_0(.douta(w_in2106_0[0]),.doutb(w_in2106_0[1]),.din(in2106));
	jspl jspl_w_in2107_0(.douta(w_in2107_0[0]),.doutb(w_in2107_0[1]),.din(in2107));
	jspl jspl_w_in2108_0(.douta(w_in2108_0[0]),.doutb(w_in2108_0[1]),.din(in2108));
	jspl jspl_w_in2109_0(.douta(w_in2109_0[0]),.doutb(w_in2109_0[1]),.din(in2109));
	jspl jspl_w_in2110_0(.douta(w_in2110_0[0]),.doutb(w_in2110_0[1]),.din(in2110));
	jspl jspl_w_in2111_0(.douta(w_in2111_0[0]),.doutb(w_in2111_0[1]),.din(in2111));
	jspl jspl_w_in2112_0(.douta(w_in2112_0[0]),.doutb(w_in2112_0[1]),.din(in2112));
	jspl jspl_w_in2113_0(.douta(w_in2113_0[0]),.doutb(w_in2113_0[1]),.din(in2113));
	jspl jspl_w_in2114_0(.douta(w_in2114_0[0]),.doutb(w_in2114_0[1]),.din(in2114));
	jspl jspl_w_in2115_0(.douta(w_in2115_0[0]),.doutb(w_in2115_0[1]),.din(in2115));
	jspl jspl_w_in2116_0(.douta(w_in2116_0[0]),.doutb(w_in2116_0[1]),.din(in2116));
	jspl jspl_w_in2117_0(.douta(w_in2117_0[0]),.doutb(w_in2117_0[1]),.din(in2117));
	jspl jspl_w_in2118_0(.douta(w_in2118_0[0]),.doutb(w_in2118_0[1]),.din(in2118));
	jspl jspl_w_in2119_0(.douta(w_in2119_0[0]),.doutb(w_in2119_0[1]),.din(in2119));
	jspl jspl_w_in2120_0(.douta(w_in2120_0[0]),.doutb(w_in2120_0[1]),.din(in2120));
	jspl jspl_w_in2121_0(.douta(w_in2121_0[0]),.doutb(w_in2121_0[1]),.din(in2121));
	jspl jspl_w_in2122_0(.douta(w_in2122_0[0]),.doutb(w_in2122_0[1]),.din(in2122));
	jspl jspl_w_in2123_0(.douta(w_in2123_0[0]),.doutb(w_in2123_0[1]),.din(in2123));
	jspl jspl_w_in2124_0(.douta(w_in2124_0[0]),.doutb(w_in2124_0[1]),.din(in2124));
	jspl jspl_w_in2125_0(.douta(w_in2125_0[0]),.doutb(w_in2125_0[1]),.din(in2125));
	jspl jspl_w_in2126_0(.douta(w_in2126_0[0]),.doutb(w_in2126_0[1]),.din(in2126));
	jspl3 jspl3_w_in2127_0(.douta(w_in2127_0[0]),.doutb(w_in2127_0[1]),.doutc(w_in2127_0[2]),.din(in2127));
	jspl3 jspl3_w_in30_0(.douta(w_in30_0[0]),.doutb(w_in30_0[1]),.doutc(w_in30_0[2]),.din(in30));
	jspl3 jspl3_w_in31_0(.douta(w_in31_0[0]),.doutb(w_in31_0[1]),.doutc(w_in31_0[2]),.din(in31));
	jspl3 jspl3_w_in32_0(.douta(w_in32_0[0]),.doutb(w_in32_0[1]),.doutc(w_in32_0[2]),.din(in32));
	jspl jspl_w_in33_0(.douta(w_in33_0[0]),.doutb(w_in33_0[1]),.din(in33));
	jspl jspl_w_in34_0(.douta(w_in34_0[0]),.doutb(w_in34_0[1]),.din(in34));
	jspl jspl_w_in35_0(.douta(w_in35_0[0]),.doutb(w_in35_0[1]),.din(in35));
	jspl jspl_w_in36_0(.douta(w_in36_0[0]),.doutb(w_in36_0[1]),.din(in36));
	jspl jspl_w_in37_0(.douta(w_in37_0[0]),.doutb(w_in37_0[1]),.din(in37));
	jspl jspl_w_in38_0(.douta(w_in38_0[0]),.doutb(w_in38_0[1]),.din(in38));
	jspl jspl_w_in39_0(.douta(w_in39_0[0]),.doutb(w_in39_0[1]),.din(in39));
	jspl jspl_w_in310_0(.douta(w_in310_0[0]),.doutb(w_in310_0[1]),.din(in310));
	jspl jspl_w_in311_0(.douta(w_in311_0[0]),.doutb(w_in311_0[1]),.din(in311));
	jspl jspl_w_in312_0(.douta(w_in312_0[0]),.doutb(w_in312_0[1]),.din(in312));
	jspl jspl_w_in313_0(.douta(w_in313_0[0]),.doutb(w_in313_0[1]),.din(in313));
	jspl jspl_w_in314_0(.douta(w_in314_0[0]),.doutb(w_in314_0[1]),.din(in314));
	jspl jspl_w_in315_0(.douta(w_in315_0[0]),.doutb(w_in315_0[1]),.din(in315));
	jspl jspl_w_in316_0(.douta(w_in316_0[0]),.doutb(w_in316_0[1]),.din(in316));
	jspl jspl_w_in317_0(.douta(w_in317_0[0]),.doutb(w_in317_0[1]),.din(in317));
	jspl jspl_w_in318_0(.douta(w_in318_0[0]),.doutb(w_in318_0[1]),.din(in318));
	jspl jspl_w_in319_0(.douta(w_in319_0[0]),.doutb(w_in319_0[1]),.din(in319));
	jspl jspl_w_in320_0(.douta(w_in320_0[0]),.doutb(w_in320_0[1]),.din(in320));
	jspl jspl_w_in321_0(.douta(w_in321_0[0]),.doutb(w_in321_0[1]),.din(in321));
	jspl jspl_w_in322_0(.douta(w_in322_0[0]),.doutb(w_in322_0[1]),.din(in322));
	jspl jspl_w_in323_0(.douta(w_in323_0[0]),.doutb(w_in323_0[1]),.din(in323));
	jspl jspl_w_in324_0(.douta(w_in324_0[0]),.doutb(w_in324_0[1]),.din(in324));
	jspl jspl_w_in325_0(.douta(w_in325_0[0]),.doutb(w_in325_0[1]),.din(in325));
	jspl jspl_w_in326_0(.douta(w_in326_0[0]),.doutb(w_in326_0[1]),.din(in326));
	jspl jspl_w_in327_0(.douta(w_in327_0[0]),.doutb(w_in327_0[1]),.din(in327));
	jspl jspl_w_in328_0(.douta(w_in328_0[0]),.doutb(w_in328_0[1]),.din(in328));
	jspl jspl_w_in329_0(.douta(w_in329_0[0]),.doutb(w_in329_0[1]),.din(in329));
	jspl jspl_w_in330_0(.douta(w_in330_0[0]),.doutb(w_in330_0[1]),.din(in330));
	jspl jspl_w_in331_0(.douta(w_in331_0[0]),.doutb(w_in331_0[1]),.din(in331));
	jspl jspl_w_in332_0(.douta(w_in332_0[0]),.doutb(w_in332_0[1]),.din(in332));
	jspl jspl_w_in333_0(.douta(w_in333_0[0]),.doutb(w_in333_0[1]),.din(in333));
	jspl jspl_w_in334_0(.douta(w_in334_0[0]),.doutb(w_in334_0[1]),.din(in334));
	jspl jspl_w_in335_0(.douta(w_in335_0[0]),.doutb(w_in335_0[1]),.din(in335));
	jspl jspl_w_in336_0(.douta(w_in336_0[0]),.doutb(w_in336_0[1]),.din(in336));
	jspl jspl_w_in337_0(.douta(w_in337_0[0]),.doutb(w_in337_0[1]),.din(in337));
	jspl jspl_w_in338_0(.douta(w_in338_0[0]),.doutb(w_in338_0[1]),.din(in338));
	jspl jspl_w_in339_0(.douta(w_in339_0[0]),.doutb(w_in339_0[1]),.din(in339));
	jspl jspl_w_in340_0(.douta(w_in340_0[0]),.doutb(w_in340_0[1]),.din(in340));
	jspl jspl_w_in341_0(.douta(w_in341_0[0]),.doutb(w_in341_0[1]),.din(in341));
	jspl jspl_w_in342_0(.douta(w_in342_0[0]),.doutb(w_in342_0[1]),.din(in342));
	jspl jspl_w_in343_0(.douta(w_in343_0[0]),.doutb(w_in343_0[1]),.din(in343));
	jspl jspl_w_in344_0(.douta(w_in344_0[0]),.doutb(w_in344_0[1]),.din(in344));
	jspl jspl_w_in345_0(.douta(w_in345_0[0]),.doutb(w_in345_0[1]),.din(in345));
	jspl jspl_w_in346_0(.douta(w_in346_0[0]),.doutb(w_in346_0[1]),.din(in346));
	jspl jspl_w_in347_0(.douta(w_in347_0[0]),.doutb(w_in347_0[1]),.din(in347));
	jspl jspl_w_in348_0(.douta(w_in348_0[0]),.doutb(w_in348_0[1]),.din(in348));
	jspl jspl_w_in349_0(.douta(w_in349_0[0]),.doutb(w_in349_0[1]),.din(in349));
	jspl jspl_w_in350_0(.douta(w_in350_0[0]),.doutb(w_in350_0[1]),.din(in350));
	jspl jspl_w_in351_0(.douta(w_in351_0[0]),.doutb(w_in351_0[1]),.din(in351));
	jspl jspl_w_in352_0(.douta(w_in352_0[0]),.doutb(w_in352_0[1]),.din(in352));
	jspl jspl_w_in353_0(.douta(w_in353_0[0]),.doutb(w_in353_0[1]),.din(in353));
	jspl jspl_w_in354_0(.douta(w_in354_0[0]),.doutb(w_in354_0[1]),.din(in354));
	jspl jspl_w_in355_0(.douta(w_in355_0[0]),.doutb(w_in355_0[1]),.din(in355));
	jspl jspl_w_in356_0(.douta(w_in356_0[0]),.doutb(w_in356_0[1]),.din(in356));
	jspl jspl_w_in357_0(.douta(w_in357_0[0]),.doutb(w_in357_0[1]),.din(in357));
	jspl jspl_w_in358_0(.douta(w_in358_0[0]),.doutb(w_in358_0[1]),.din(in358));
	jspl jspl_w_in359_0(.douta(w_in359_0[0]),.doutb(w_in359_0[1]),.din(in359));
	jspl jspl_w_in360_0(.douta(w_in360_0[0]),.doutb(w_in360_0[1]),.din(in360));
	jspl jspl_w_in361_0(.douta(w_in361_0[0]),.doutb(w_in361_0[1]),.din(in361));
	jspl jspl_w_in362_0(.douta(w_in362_0[0]),.doutb(w_in362_0[1]),.din(in362));
	jspl jspl_w_in363_0(.douta(w_in363_0[0]),.doutb(w_in363_0[1]),.din(in363));
	jspl jspl_w_in364_0(.douta(w_in364_0[0]),.doutb(w_in364_0[1]),.din(in364));
	jspl jspl_w_in365_0(.douta(w_in365_0[0]),.doutb(w_in365_0[1]),.din(in365));
	jspl jspl_w_in366_0(.douta(w_in366_0[0]),.doutb(w_in366_0[1]),.din(in366));
	jspl jspl_w_in367_0(.douta(w_in367_0[0]),.doutb(w_in367_0[1]),.din(in367));
	jspl jspl_w_in368_0(.douta(w_in368_0[0]),.doutb(w_in368_0[1]),.din(in368));
	jspl jspl_w_in369_0(.douta(w_in369_0[0]),.doutb(w_in369_0[1]),.din(in369));
	jspl jspl_w_in370_0(.douta(w_in370_0[0]),.doutb(w_in370_0[1]),.din(in370));
	jspl jspl_w_in371_0(.douta(w_in371_0[0]),.doutb(w_in371_0[1]),.din(in371));
	jspl jspl_w_in372_0(.douta(w_in372_0[0]),.doutb(w_in372_0[1]),.din(in372));
	jspl jspl_w_in373_0(.douta(w_in373_0[0]),.doutb(w_in373_0[1]),.din(in373));
	jspl jspl_w_in374_0(.douta(w_in374_0[0]),.doutb(w_in374_0[1]),.din(in374));
	jspl jspl_w_in375_0(.douta(w_in375_0[0]),.doutb(w_in375_0[1]),.din(in375));
	jspl jspl_w_in376_0(.douta(w_in376_0[0]),.doutb(w_in376_0[1]),.din(in376));
	jspl jspl_w_in377_0(.douta(w_in377_0[0]),.doutb(w_in377_0[1]),.din(in377));
	jspl jspl_w_in378_0(.douta(w_in378_0[0]),.doutb(w_in378_0[1]),.din(in378));
	jspl jspl_w_in379_0(.douta(w_in379_0[0]),.doutb(w_in379_0[1]),.din(in379));
	jspl jspl_w_in380_0(.douta(w_in380_0[0]),.doutb(w_in380_0[1]),.din(in380));
	jspl jspl_w_in381_0(.douta(w_in381_0[0]),.doutb(w_in381_0[1]),.din(in381));
	jspl jspl_w_in382_0(.douta(w_in382_0[0]),.doutb(w_in382_0[1]),.din(in382));
	jspl jspl_w_in383_0(.douta(w_in383_0[0]),.doutb(w_in383_0[1]),.din(in383));
	jspl jspl_w_in384_0(.douta(w_in384_0[0]),.doutb(w_in384_0[1]),.din(in384));
	jspl jspl_w_in385_0(.douta(w_in385_0[0]),.doutb(w_in385_0[1]),.din(in385));
	jspl jspl_w_in386_0(.douta(w_in386_0[0]),.doutb(w_in386_0[1]),.din(in386));
	jspl jspl_w_in387_0(.douta(w_in387_0[0]),.doutb(w_in387_0[1]),.din(in387));
	jspl jspl_w_in388_0(.douta(w_in388_0[0]),.doutb(w_in388_0[1]),.din(in388));
	jspl jspl_w_in389_0(.douta(w_in389_0[0]),.doutb(w_in389_0[1]),.din(in389));
	jspl jspl_w_in390_0(.douta(w_in390_0[0]),.doutb(w_in390_0[1]),.din(in390));
	jspl jspl_w_in391_0(.douta(w_in391_0[0]),.doutb(w_in391_0[1]),.din(in391));
	jspl jspl_w_in392_0(.douta(w_in392_0[0]),.doutb(w_in392_0[1]),.din(in392));
	jspl jspl_w_in393_0(.douta(w_in393_0[0]),.doutb(w_in393_0[1]),.din(in393));
	jspl jspl_w_in394_0(.douta(w_in394_0[0]),.doutb(w_in394_0[1]),.din(in394));
	jspl jspl_w_in395_0(.douta(w_in395_0[0]),.doutb(w_in395_0[1]),.din(in395));
	jspl jspl_w_in396_0(.douta(w_in396_0[0]),.doutb(w_in396_0[1]),.din(in396));
	jspl jspl_w_in397_0(.douta(w_in397_0[0]),.doutb(w_in397_0[1]),.din(in397));
	jspl jspl_w_in398_0(.douta(w_in398_0[0]),.doutb(w_in398_0[1]),.din(in398));
	jspl jspl_w_in399_0(.douta(w_in399_0[0]),.doutb(w_in399_0[1]),.din(in399));
	jspl jspl_w_in3100_0(.douta(w_in3100_0[0]),.doutb(w_in3100_0[1]),.din(in3100));
	jspl jspl_w_in3101_0(.douta(w_in3101_0[0]),.doutb(w_in3101_0[1]),.din(in3101));
	jspl jspl_w_in3102_0(.douta(w_in3102_0[0]),.doutb(w_in3102_0[1]),.din(in3102));
	jspl jspl_w_in3103_0(.douta(w_in3103_0[0]),.doutb(w_in3103_0[1]),.din(in3103));
	jspl jspl_w_in3104_0(.douta(w_in3104_0[0]),.doutb(w_in3104_0[1]),.din(in3104));
	jspl jspl_w_in3105_0(.douta(w_in3105_0[0]),.doutb(w_in3105_0[1]),.din(in3105));
	jspl jspl_w_in3106_0(.douta(w_in3106_0[0]),.doutb(w_in3106_0[1]),.din(in3106));
	jspl jspl_w_in3107_0(.douta(w_in3107_0[0]),.doutb(w_in3107_0[1]),.din(in3107));
	jspl jspl_w_in3108_0(.douta(w_in3108_0[0]),.doutb(w_in3108_0[1]),.din(in3108));
	jspl jspl_w_in3109_0(.douta(w_in3109_0[0]),.doutb(w_in3109_0[1]),.din(in3109));
	jspl jspl_w_in3110_0(.douta(w_in3110_0[0]),.doutb(w_in3110_0[1]),.din(in3110));
	jspl jspl_w_in3111_0(.douta(w_in3111_0[0]),.doutb(w_in3111_0[1]),.din(in3111));
	jspl jspl_w_in3112_0(.douta(w_in3112_0[0]),.doutb(w_in3112_0[1]),.din(in3112));
	jspl jspl_w_in3113_0(.douta(w_in3113_0[0]),.doutb(w_in3113_0[1]),.din(in3113));
	jspl jspl_w_in3114_0(.douta(w_in3114_0[0]),.doutb(w_in3114_0[1]),.din(in3114));
	jspl jspl_w_in3115_0(.douta(w_in3115_0[0]),.doutb(w_in3115_0[1]),.din(in3115));
	jspl jspl_w_in3116_0(.douta(w_in3116_0[0]),.doutb(w_in3116_0[1]),.din(in3116));
	jspl jspl_w_in3117_0(.douta(w_in3117_0[0]),.doutb(w_in3117_0[1]),.din(in3117));
	jspl jspl_w_in3118_0(.douta(w_in3118_0[0]),.doutb(w_in3118_0[1]),.din(in3118));
	jspl jspl_w_in3119_0(.douta(w_in3119_0[0]),.doutb(w_in3119_0[1]),.din(in3119));
	jspl jspl_w_in3120_0(.douta(w_in3120_0[0]),.doutb(w_in3120_0[1]),.din(in3120));
	jspl jspl_w_in3121_0(.douta(w_in3121_0[0]),.doutb(w_in3121_0[1]),.din(in3121));
	jspl jspl_w_in3122_0(.douta(w_in3122_0[0]),.doutb(w_in3122_0[1]),.din(in3122));
	jspl jspl_w_in3123_0(.douta(w_in3123_0[0]),.doutb(w_in3123_0[1]),.din(in3123));
	jspl jspl_w_in3124_0(.douta(w_in3124_0[0]),.doutb(w_in3124_0[1]),.din(in3124));
	jspl jspl_w_in3125_0(.douta(w_in3125_0[0]),.doutb(w_in3125_0[1]),.din(in3125));
	jspl jspl_w_in3126_0(.douta(w_in3126_0[0]),.doutb(w_in3126_0[1]),.din(in3126));
	jspl jspl_w_in3127_0(.douta(w_in3127_0[0]),.doutb(w_in3127_0[1]),.din(in3127));
	jspl3 jspl3_w_address1_0(.douta(w_address1_0[0]),.doutb(w_address1_0[1]),.doutc(w_address1_0[2]),.din(address1_fa_));
	jspl3 jspl3_w_address1_1(.douta(w_address1_1[0]),.doutb(w_address1_1[1]),.doutc(w_address1_1[2]),.din(w_address1_0[0]));
	jspl3 jspl3_w_address1_2(.douta(w_address1_2[0]),.doutb(w_address1_2[1]),.doutc(w_address1_2[2]),.din(w_address1_0[1]));
	jspl3 jspl3_w_address1_3(.douta(w_address1_3[0]),.doutb(w_address1_3[1]),.doutc(w_address1_3[2]),.din(w_address1_0[2]));
	jspl3 jspl3_w_address1_4(.douta(w_address1_4[0]),.doutb(w_address1_4[1]),.doutc(w_address1_4[2]),.din(w_address1_1[0]));
	jspl3 jspl3_w_address1_5(.douta(w_address1_5[0]),.doutb(w_address1_5[1]),.doutc(w_address1_5[2]),.din(w_address1_1[1]));
	jspl3 jspl3_w_address1_6(.douta(w_address1_6[0]),.doutb(w_address1_6[1]),.doutc(w_address1_6[2]),.din(w_address1_1[2]));
	jspl3 jspl3_w_address1_7(.douta(w_address1_7[0]),.doutb(w_address1_7[1]),.doutc(w_address1_7[2]),.din(w_address1_2[0]));
	jspl3 jspl3_w_address1_8(.douta(w_address1_8[0]),.doutb(w_address1_8[1]),.doutc(w_address1_8[2]),.din(w_address1_2[1]));
	jspl3 jspl3_w_address1_9(.douta(w_address1_9[0]),.doutb(w_address1_9[1]),.doutc(w_address1_9[2]),.din(w_address1_2[2]));
	jspl3 jspl3_w_address1_10(.douta(w_address1_10[0]),.doutb(w_address1_10[1]),.doutc(w_address1_10[2]),.din(w_address1_3[0]));
	jspl3 jspl3_w_address1_11(.douta(w_address1_11[0]),.doutb(w_address1_11[1]),.doutc(w_address1_11[2]),.din(w_address1_3[1]));
	jspl3 jspl3_w_address1_12(.douta(w_address1_12[0]),.doutb(w_address1_12[1]),.doutc(w_address1_12[2]),.din(w_address1_3[2]));
	jspl3 jspl3_w_address1_13(.douta(w_address1_13[0]),.doutb(w_address1_13[1]),.doutc(w_address1_13[2]),.din(w_address1_4[0]));
	jspl3 jspl3_w_address1_14(.douta(w_address1_14[0]),.doutb(w_address1_14[1]),.doutc(w_address1_14[2]),.din(w_address1_4[1]));
	jspl3 jspl3_w_address1_15(.douta(w_address1_15[0]),.doutb(w_address1_15[1]),.doutc(w_address1_15[2]),.din(w_address1_4[2]));
	jspl3 jspl3_w_address1_16(.douta(w_address1_16[0]),.doutb(w_address1_16[1]),.doutc(w_address1_16[2]),.din(w_address1_5[0]));
	jspl3 jspl3_w_address1_17(.douta(w_address1_17[0]),.doutb(w_address1_17[1]),.doutc(w_address1_17[2]),.din(w_address1_5[1]));
	jspl3 jspl3_w_address1_18(.douta(w_address1_18[0]),.doutb(w_address1_18[1]),.doutc(w_address1_18[2]),.din(w_address1_5[2]));
	jspl3 jspl3_w_address1_19(.douta(w_address1_19[0]),.doutb(w_address1_19[1]),.doutc(w_address1_19[2]),.din(w_address1_6[0]));
	jspl3 jspl3_w_address1_20(.douta(w_address1_20[0]),.doutb(w_address1_20[1]),.doutc(w_address1_20[2]),.din(w_address1_6[1]));
	jspl3 jspl3_w_address1_21(.douta(w_address1_21[0]),.doutb(w_address1_21[1]),.doutc(w_address1_21[2]),.din(w_address1_6[2]));
	jspl3 jspl3_w_address1_22(.douta(w_address1_22[0]),.doutb(w_address1_22[1]),.doutc(w_address1_22[2]),.din(w_address1_7[0]));
	jspl3 jspl3_w_address1_23(.douta(w_address1_23[0]),.doutb(w_address1_23[1]),.doutc(w_address1_23[2]),.din(w_address1_7[1]));
	jspl3 jspl3_w_address1_24(.douta(w_address1_24[0]),.doutb(w_address1_24[1]),.doutc(w_address1_24[2]),.din(w_address1_7[2]));
	jspl3 jspl3_w_address1_25(.douta(w_address1_25[0]),.doutb(w_address1_25[1]),.doutc(w_address1_25[2]),.din(w_address1_8[0]));
	jspl3 jspl3_w_address1_26(.douta(w_address1_26[0]),.doutb(w_address1_26[1]),.doutc(w_address1_26[2]),.din(w_address1_8[1]));
	jspl3 jspl3_w_address1_27(.douta(w_address1_27[0]),.doutb(w_address1_27[1]),.doutc(w_address1_27[2]),.din(w_address1_8[2]));
	jspl3 jspl3_w_address1_28(.douta(w_address1_28[0]),.doutb(w_address1_28[1]),.doutc(w_address1_28[2]),.din(w_address1_9[0]));
	jspl3 jspl3_w_address1_29(.douta(w_address1_29[0]),.doutb(w_address1_29[1]),.doutc(w_address1_29[2]),.din(w_address1_9[1]));
	jspl3 jspl3_w_address1_30(.douta(w_address1_30[0]),.doutb(w_address1_30[1]),.doutc(w_address1_30[2]),.din(w_address1_9[2]));
	jspl3 jspl3_w_address1_31(.douta(w_address1_31[0]),.doutb(w_address1_31[1]),.doutc(w_address1_31[2]),.din(w_address1_10[0]));
	jspl3 jspl3_w_address1_32(.douta(w_address1_32[0]),.doutb(w_address1_32[1]),.doutc(w_address1_32[2]),.din(w_address1_10[1]));
	jspl3 jspl3_w_address1_33(.douta(w_address1_33[0]),.doutb(w_address1_33[1]),.doutc(w_address1_33[2]),.din(w_address1_10[2]));
	jspl3 jspl3_w_address1_34(.douta(w_address1_34[0]),.doutb(w_address1_34[1]),.doutc(w_address1_34[2]),.din(w_address1_11[0]));
	jspl3 jspl3_w_address1_35(.douta(w_address1_35[0]),.doutb(w_address1_35[1]),.doutc(w_address1_35[2]),.din(w_address1_11[1]));
	jspl3 jspl3_w_address1_36(.douta(w_address1_36[0]),.doutb(w_address1_36[1]),.doutc(w_address1_36[2]),.din(w_address1_11[2]));
	jspl3 jspl3_w_address1_37(.douta(w_address1_37[0]),.doutb(w_address1_37[1]),.doutc(w_address1_37[2]),.din(w_address1_12[0]));
	jspl3 jspl3_w_address1_38(.douta(w_address1_38[0]),.doutb(w_address1_38[1]),.doutc(w_address1_38[2]),.din(w_address1_12[1]));
	jspl3 jspl3_w_address1_39(.douta(w_address1_39[0]),.doutb(w_address1_39[1]),.doutc(w_address1_39[2]),.din(w_address1_12[2]));
	jspl3 jspl3_w_address1_40(.douta(w_address1_40[0]),.doutb(w_address1_40[1]),.doutc(w_address1_40[2]),.din(w_address1_13[0]));
	jspl3 jspl3_w_address1_41(.douta(w_address1_41[0]),.doutb(w_address1_41[1]),.doutc(w_address1_41[2]),.din(w_address1_13[1]));
	jspl3 jspl3_w_address1_42(.douta(w_address1_42[0]),.doutb(w_address1_42[1]),.doutc(w_address1_42[2]),.din(w_address1_13[2]));
	jspl3 jspl3_w_address1_43(.douta(w_address1_43[0]),.doutb(w_address1_43[1]),.doutc(w_address1_43[2]),.din(w_address1_14[0]));
	jspl3 jspl3_w_address1_44(.douta(w_address1_44[0]),.doutb(w_address1_44[1]),.doutc(w_address1_44[2]),.din(w_address1_14[1]));
	jspl3 jspl3_w_address1_45(.douta(w_address1_45[0]),.doutb(w_address1_45[1]),.doutc(w_address1_45[2]),.din(w_address1_14[2]));
	jspl3 jspl3_w_address1_46(.douta(w_address1_46[0]),.doutb(w_address1_46[1]),.doutc(w_address1_46[2]),.din(w_address1_15[0]));
	jspl3 jspl3_w_address1_47(.douta(w_address1_47[0]),.doutb(w_address1_47[1]),.doutc(w_address1_47[2]),.din(w_address1_15[1]));
	jspl3 jspl3_w_address1_48(.douta(w_address1_48[0]),.doutb(w_address1_48[1]),.doutc(w_address1_48[2]),.din(w_address1_15[2]));
	jspl3 jspl3_w_address1_49(.douta(w_address1_49[0]),.doutb(w_address1_49[1]),.doutc(w_address1_49[2]),.din(w_address1_16[0]));
	jspl3 jspl3_w_address1_50(.douta(w_address1_50[0]),.doutb(w_address1_50[1]),.doutc(w_address1_50[2]),.din(w_address1_16[1]));
	jspl3 jspl3_w_address1_51(.douta(w_address1_51[0]),.doutb(w_address1_51[1]),.doutc(w_address1_51[2]),.din(w_address1_16[2]));
	jspl3 jspl3_w_address1_52(.douta(w_address1_52[0]),.doutb(w_address1_52[1]),.doutc(w_address1_52[2]),.din(w_address1_17[0]));
	jspl3 jspl3_w_address1_53(.douta(w_address1_53[0]),.doutb(w_address1_53[1]),.doutc(w_address1_53[2]),.din(w_address1_17[1]));
	jspl3 jspl3_w_address1_54(.douta(w_address1_54[0]),.doutb(w_address1_54[1]),.doutc(w_address1_54[2]),.din(w_address1_17[2]));
	jspl3 jspl3_w_address1_55(.douta(w_address1_55[0]),.doutb(w_address1_55[1]),.doutc(w_address1_55[2]),.din(w_address1_18[0]));
	jspl3 jspl3_w_address1_56(.douta(w_address1_56[0]),.doutb(w_address1_56[1]),.doutc(w_address1_56[2]),.din(w_address1_18[1]));
	jspl3 jspl3_w_address1_57(.douta(w_address1_57[0]),.doutb(w_address1_57[1]),.doutc(w_address1_57[2]),.din(w_address1_18[2]));
	jspl3 jspl3_w_address1_58(.douta(w_address1_58[0]),.doutb(w_address1_58[1]),.doutc(w_address1_58[2]),.din(w_address1_19[0]));
	jspl3 jspl3_w_address1_59(.douta(w_address1_59[0]),.doutb(w_address1_59[1]),.doutc(w_address1_59[2]),.din(w_address1_19[1]));
	jspl3 jspl3_w_address1_60(.douta(w_address1_60[0]),.doutb(w_address1_60[1]),.doutc(w_address1_60[2]),.din(w_address1_19[2]));
	jspl3 jspl3_w_address1_61(.douta(w_address1_61[0]),.doutb(w_address1_61[1]),.doutc(w_address1_61[2]),.din(w_address1_20[0]));
	jspl3 jspl3_w_address1_62(.douta(w_address1_62[0]),.doutb(w_address1_62[1]),.doutc(w_address1_62[2]),.din(w_address1_20[1]));
	jspl3 jspl3_w_address1_63(.douta(w_address1_63[0]),.doutb(w_address1_63[1]),.doutc(w_dff_A_J7blzP2R6_2),.din(w_address1_20[2]));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl jspl_w_n643_0(.douta(w_n643_0[0]),.doutb(w_n643_0[1]),.din(n643));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl jspl_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.din(n648));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.din(n653));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(n654));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n668_0(.douta(w_n668_0[0]),.doutb(w_n668_0[1]),.din(n668));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(n674));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.din(n679));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.din(n707));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(n709));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.din(n725));
	jspl jspl_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.din(n730));
	jspl jspl_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.din(n732));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(n739));
	jspl jspl_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl jspl_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.din(n743));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl jspl_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.din(n746));
	jspl jspl_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.din(n748));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(n749));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.din(n753));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(n764));
	jspl jspl_w_n768_0(.douta(w_n768_0[0]),.doutb(w_n768_0[1]),.din(n768));
	jspl jspl_w_n770_0(.douta(w_n770_0[0]),.doutb(w_n770_0[1]),.din(n770));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n776_0(.douta(w_n776_0[0]),.doutb(w_n776_0[1]),.din(n776));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.din(n789));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl jspl_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.din(n801));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.din(n804));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(n807));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.din(n812));
	jspl jspl_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.din(n814));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n836_0(.douta(w_n836_0[0]),.doutb(w_n836_0[1]),.din(n836));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(n837));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl jspl_w_n841_0(.douta(w_n841_0[0]),.doutb(w_n841_0[1]),.din(n841));
	jspl jspl_w_n844_0(.douta(w_n844_0[0]),.doutb(w_n844_0[1]),.din(n844));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(n846));
	jspl jspl_w_n848_0(.douta(w_n848_0[0]),.doutb(w_n848_0[1]),.din(n848));
	jspl jspl_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.din(n853));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(n861));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.din(n870));
	jspl jspl_w_n872_0(.douta(w_n872_0[0]),.doutb(w_n872_0[1]),.din(n872));
	jspl jspl_w_n875_0(.douta(w_n875_0[0]),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl jspl_w_n878_0(.douta(w_n878_0[0]),.doutb(w_n878_0[1]),.din(n878));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.din(n882));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl jspl_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.din(n888));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(n898));
	jspl jspl_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.din(n900));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_n901_0[1]),.din(n901));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_n904_0[1]),.din(n904));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(n907));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(n911));
	jspl jspl_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.din(n912));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(n915));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl3 jspl3_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.doutc(w_n922_0[2]),.din(n922));
	jspl jspl_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.din(n925));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_n931_0[1]),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n934_0(.douta(w_n934_0[0]),.doutb(w_n934_0[1]),.din(n934));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(n939));
	jspl jspl_w_n941_0(.douta(w_n941_0[0]),.doutb(w_n941_0[1]),.din(n941));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(n943));
	jspl jspl_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.din(n946));
	jspl jspl_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.din(n947));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl jspl_w_n955_0(.douta(w_n955_0[0]),.doutb(w_n955_0[1]),.din(n955));
	jspl jspl_w_n958_0(.douta(w_n958_0[0]),.doutb(w_n958_0[1]),.din(n958));
	jspl jspl_w_n960_0(.douta(w_n960_0[0]),.doutb(w_n960_0[1]),.din(n960));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n963_0(.douta(w_n963_0[0]),.doutb(w_n963_0[1]),.din(n963));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n967_0(.douta(w_n967_0[0]),.doutb(w_n967_0[1]),.din(n967));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_n968_0[1]),.din(n968));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_n971_0[1]),.din(n971));
	jspl jspl_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.din(n973));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n975_0(.douta(w_n975_0[0]),.doutb(w_n975_0[1]),.din(n975));
	jspl jspl_w_n976_0(.douta(w_n976_0[0]),.doutb(w_n976_0[1]),.din(n976));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.din(n980));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.din(n983));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(n988));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(n990));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.din(n995));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(n996));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.din(n1006));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.din(n1010));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.din(n1012));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(n1016));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(n1018));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(n1020));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.din(n1025));
	jspl jspl_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(n1028));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.din(n1030));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.din(n1032));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1034_0(.douta(w_n1034_0[0]),.doutb(w_n1034_0[1]),.din(n1034));
	jspl jspl_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.din(n1035));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(n1037));
	jspl jspl_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.din(n1038));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.din(n1039));
	jspl jspl_w_n1040_0(.douta(w_n1040_0[0]),.doutb(w_n1040_0[1]),.din(n1040));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1042_0(.douta(w_n1042_0[0]),.doutb(w_n1042_0[1]),.din(n1042));
	jspl3 jspl3_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.doutc(w_n1044_0[2]),.din(n1044));
	jspl jspl_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.din(n1046));
	jspl jspl_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.din(n1049));
	jspl jspl_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.din(n1054));
	jspl jspl_w_n1055_0(.douta(w_n1055_0[0]),.doutb(w_n1055_0[1]),.din(n1055));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1060_0(.douta(w_n1060_0[0]),.doutb(w_n1060_0[1]),.din(n1060));
	jspl jspl_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.din(n1063));
	jspl jspl_w_n1065_0(.douta(w_n1065_0[0]),.doutb(w_n1065_0[1]),.din(n1065));
	jspl jspl_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.din(n1067));
	jspl jspl_w_n1070_0(.douta(w_n1070_0[0]),.doutb(w_n1070_0[1]),.din(n1070));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(n1072));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(n1074));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(n1083));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(n1084));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(n1089));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(n1091));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1098_0(.douta(w_n1098_0[0]),.doutb(w_n1098_0[1]),.din(n1098));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_n1108_0[1]),.din(n1108));
	jspl jspl_w_n1110_0(.douta(w_n1110_0[0]),.doutb(w_n1110_0[1]),.din(n1110));
	jspl jspl_w_n1112_0(.douta(w_n1112_0[0]),.doutb(w_n1112_0[1]),.din(n1112));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(n1119));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(n1121));
	jspl jspl_w_n1123_0(.douta(w_n1123_0[0]),.doutb(w_n1123_0[1]),.din(n1123));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(n1126));
	jspl jspl_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.din(n1128));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_n1140_0[1]),.din(n1140));
	jspl jspl_w_n1142_0(.douta(w_n1142_0[0]),.doutb(w_n1142_0[1]),.din(n1142));
	jspl jspl_w_n1144_0(.douta(w_n1144_0[0]),.doutb(w_n1144_0[1]),.din(n1144));
	jspl jspl_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_n1147_0[1]),.din(n1147));
	jspl jspl_w_n1148_0(.douta(w_n1148_0[0]),.doutb(w_n1148_0[1]),.din(n1148));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl jspl_w_n1153_0(.douta(w_n1153_0[0]),.doutb(w_n1153_0[1]),.din(n1153));
	jspl jspl_w_n1155_0(.douta(w_n1155_0[0]),.doutb(w_n1155_0[1]),.din(n1155));
	jspl jspl_w_n1158_0(.douta(w_n1158_0[0]),.doutb(w_n1158_0[1]),.din(n1158));
	jspl jspl_w_n1160_0(.douta(w_n1160_0[0]),.doutb(w_n1160_0[1]),.din(n1160));
	jspl jspl_w_n1162_0(.douta(w_n1162_0[0]),.doutb(w_n1162_0[1]),.din(n1162));
	jspl jspl_w_n1172_0(.douta(w_n1172_0[0]),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1174_0(.douta(w_n1174_0[0]),.doutb(w_n1174_0[1]),.din(n1174));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(n1188));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(n1190));
	jspl jspl_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.din(n1195));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(n1206));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1218_0(.douta(w_n1218_0[0]),.doutb(w_n1218_0[1]),.din(n1218));
	jspl jspl_w_n1223_0(.douta(w_n1223_0[0]),.doutb(w_n1223_0[1]),.din(n1223));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1233_0(.douta(w_n1233_0[0]),.doutb(w_n1233_0[1]),.din(n1233));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1239_0(.douta(w_n1239_0[0]),.doutb(w_n1239_0[1]),.din(n1239));
	jspl jspl_w_n1241_0(.douta(w_n1241_0[0]),.doutb(w_n1241_0[1]),.din(n1241));
	jspl jspl_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.din(n1242));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(n1248));
	jspl jspl_w_n1250_0(.douta(w_n1250_0[0]),.doutb(w_n1250_0[1]),.din(n1250));
	jspl jspl_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.din(n1253));
	jspl jspl_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.din(n1255));
	jspl jspl_w_n1258_0(.douta(w_n1258_0[0]),.doutb(w_n1258_0[1]),.din(n1258));
	jspl jspl_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.din(n1263));
	jspl jspl_w_n1267_0(.douta(w_n1267_0[0]),.doutb(w_n1267_0[1]),.din(n1267));
	jspl jspl_w_n1270_0(.douta(w_n1270_0[0]),.doutb(w_n1270_0[1]),.din(n1270));
	jspl jspl_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.din(n1272));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(n1278));
	jspl jspl_w_n1282_0(.douta(w_n1282_0[0]),.doutb(w_n1282_0[1]),.din(n1282));
	jspl jspl_w_n1285_0(.douta(w_n1285_0[0]),.doutb(w_n1285_0[1]),.din(n1285));
	jspl jspl_w_n1287_0(.douta(w_n1287_0[0]),.doutb(w_n1287_0[1]),.din(n1287));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1290_0(.douta(w_n1290_0[0]),.doutb(w_n1290_0[1]),.din(n1290));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_n1294_0[1]),.din(n1294));
	jspl jspl_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.din(n1296));
	jspl jspl_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.din(n1299));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1304_0(.douta(w_n1304_0[0]),.doutb(w_n1304_0[1]),.din(n1304));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(n1312));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl jspl_w_n1324_0(.douta(w_n1324_0[0]),.doutb(w_n1324_0[1]),.din(n1324));
	jspl jspl_w_n1328_0(.douta(w_n1328_0[0]),.doutb(w_n1328_0[1]),.din(n1328));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl jspl_w_n1333_0(.douta(w_n1333_0[0]),.doutb(w_n1333_0[1]),.din(n1333));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(n1337));
	jspl jspl_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.din(n1340));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(n1342));
	jspl jspl_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.din(n1345));
	jspl jspl_w_n1347_0(.douta(w_n1347_0[0]),.doutb(w_n1347_0[1]),.din(n1347));
	jspl jspl_w_n1349_0(.douta(w_n1349_0[0]),.doutb(w_n1349_0[1]),.din(n1349));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(n1352));
	jspl jspl_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.din(n1353));
	jspl jspl_w_n1355_0(.douta(w_n1355_0[0]),.doutb(w_n1355_0[1]),.din(n1355));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1374_0(.douta(w_n1374_0[0]),.doutb(w_n1374_0[1]),.din(n1374));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_n1379_0[1]),.din(n1379));
	jspl jspl_w_n1380_0(.douta(w_n1380_0[0]),.doutb(w_n1380_0[1]),.din(n1380));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(n1382));
	jspl jspl_w_n1386_0(.douta(w_n1386_0[0]),.doutb(w_n1386_0[1]),.din(n1386));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.din(n1401));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.din(n1404));
	jspl jspl_w_n1406_0(.douta(w_n1406_0[0]),.doutb(w_n1406_0[1]),.din(n1406));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1412_0(.douta(w_n1412_0[0]),.doutb(w_n1412_0[1]),.din(n1412));
	jspl jspl_w_n1414_0(.douta(w_n1414_0[0]),.doutb(w_n1414_0[1]),.din(n1414));
	jspl jspl_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.din(n1418));
	jspl jspl_w_n1422_0(.douta(w_n1422_0[0]),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(n1426));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(n1428));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(n1431));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_n1438_0[1]),.din(n1438));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(n1449));
	jspl jspl_w_n1453_0(.douta(w_n1453_0[0]),.doutb(w_n1453_0[1]),.din(n1453));
	jspl jspl_w_n1455_0(.douta(w_n1455_0[0]),.doutb(w_n1455_0[1]),.din(n1455));
	jspl jspl_w_n1458_0(.douta(w_n1458_0[0]),.doutb(w_n1458_0[1]),.din(n1458));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(n1460));
	jspl jspl_w_n1462_0(.douta(w_n1462_0[0]),.doutb(w_n1462_0[1]),.din(n1462));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(n1465));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(n1466));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1482_0(.douta(w_n1482_0[0]),.doutb(w_n1482_0[1]),.din(n1482));
	jspl jspl_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.din(n1485));
	jspl jspl_w_n1487_0(.douta(w_n1487_0[0]),.doutb(w_n1487_0[1]),.din(n1487));
	jspl jspl_w_n1489_0(.douta(w_n1489_0[0]),.doutb(w_n1489_0[1]),.din(n1489));
	jspl jspl_w_n1492_0(.douta(w_n1492_0[0]),.doutb(w_n1492_0[1]),.din(n1492));
	jspl jspl_w_n1493_0(.douta(w_n1493_0[0]),.doutb(w_n1493_0[1]),.din(n1493));
	jspl jspl_w_n1495_0(.douta(w_n1495_0[0]),.doutb(w_n1495_0[1]),.din(n1495));
	jspl jspl_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.din(n1499));
	jspl jspl_w_n1503_0(.douta(w_n1503_0[0]),.doutb(w_n1503_0[1]),.din(n1503));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(n1507));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(n1512));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl jspl_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.din(n1516));
	jspl jspl_w_n1519_0(.douta(w_n1519_0[0]),.doutb(w_n1519_0[1]),.din(n1519));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(n1520));
	jspl jspl_w_n1522_0(.douta(w_n1522_0[0]),.doutb(w_n1522_0[1]),.din(n1522));
	jspl jspl_w_n1526_0(.douta(w_n1526_0[0]),.doutb(w_n1526_0[1]),.din(n1526));
	jspl jspl_w_n1530_0(.douta(w_n1530_0[0]),.doutb(w_n1530_0[1]),.din(n1530));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1536_0(.douta(w_n1536_0[0]),.doutb(w_n1536_0[1]),.din(n1536));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.din(n1542));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(n1550));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl3 jspl3_w_n1562_0(.douta(w_n1562_0[0]),.doutb(w_n1562_0[1]),.doutc(w_n1562_0[2]),.din(n1562));
	jspl3 jspl3_w_n1562_1(.douta(w_n1562_1[0]),.doutb(w_n1562_1[1]),.doutc(w_n1562_1[2]),.din(w_n1562_0[0]));
	jspl3 jspl3_w_n1562_2(.douta(w_n1562_2[0]),.doutb(w_n1562_2[1]),.doutc(w_n1562_2[2]),.din(w_n1562_0[1]));
	jspl3 jspl3_w_n1562_3(.douta(w_n1562_3[0]),.doutb(w_n1562_3[1]),.doutc(w_n1562_3[2]),.din(w_n1562_0[2]));
	jspl3 jspl3_w_n1562_4(.douta(w_n1562_4[0]),.doutb(w_n1562_4[1]),.doutc(w_n1562_4[2]),.din(w_n1562_1[0]));
	jspl3 jspl3_w_n1562_5(.douta(w_n1562_5[0]),.doutb(w_n1562_5[1]),.doutc(w_n1562_5[2]),.din(w_n1562_1[1]));
	jspl3 jspl3_w_n1562_6(.douta(w_n1562_6[0]),.doutb(w_n1562_6[1]),.doutc(w_n1562_6[2]),.din(w_n1562_1[2]));
	jspl3 jspl3_w_n1562_7(.douta(w_n1562_7[0]),.doutb(w_n1562_7[1]),.doutc(w_n1562_7[2]),.din(w_n1562_2[0]));
	jspl3 jspl3_w_n1562_8(.douta(w_n1562_8[0]),.doutb(w_n1562_8[1]),.doutc(w_n1562_8[2]),.din(w_n1562_2[1]));
	jspl3 jspl3_w_n1562_9(.douta(w_n1562_9[0]),.doutb(w_n1562_9[1]),.doutc(w_n1562_9[2]),.din(w_n1562_2[2]));
	jspl3 jspl3_w_n1562_10(.douta(w_n1562_10[0]),.doutb(w_n1562_10[1]),.doutc(w_n1562_10[2]),.din(w_n1562_3[0]));
	jspl3 jspl3_w_n1562_11(.douta(w_n1562_11[0]),.doutb(w_n1562_11[1]),.doutc(w_n1562_11[2]),.din(w_n1562_3[1]));
	jspl3 jspl3_w_n1562_12(.douta(w_n1562_12[0]),.doutb(w_n1562_12[1]),.doutc(w_n1562_12[2]),.din(w_n1562_3[2]));
	jspl3 jspl3_w_n1562_13(.douta(w_n1562_13[0]),.doutb(w_n1562_13[1]),.doutc(w_n1562_13[2]),.din(w_n1562_4[0]));
	jspl3 jspl3_w_n1562_14(.douta(w_n1562_14[0]),.doutb(w_n1562_14[1]),.doutc(w_n1562_14[2]),.din(w_n1562_4[1]));
	jspl3 jspl3_w_n1562_15(.douta(w_n1562_15[0]),.doutb(w_n1562_15[1]),.doutc(w_n1562_15[2]),.din(w_n1562_4[2]));
	jspl3 jspl3_w_n1562_16(.douta(w_n1562_16[0]),.doutb(w_n1562_16[1]),.doutc(w_n1562_16[2]),.din(w_n1562_5[0]));
	jspl3 jspl3_w_n1562_17(.douta(w_n1562_17[0]),.doutb(w_n1562_17[1]),.doutc(w_n1562_17[2]),.din(w_n1562_5[1]));
	jspl3 jspl3_w_n1562_18(.douta(w_n1562_18[0]),.doutb(w_n1562_18[1]),.doutc(w_n1562_18[2]),.din(w_n1562_5[2]));
	jspl3 jspl3_w_n1562_19(.douta(w_n1562_19[0]),.doutb(w_n1562_19[1]),.doutc(w_n1562_19[2]),.din(w_n1562_6[0]));
	jspl3 jspl3_w_n1562_20(.douta(w_n1562_20[0]),.doutb(w_n1562_20[1]),.doutc(w_n1562_20[2]),.din(w_n1562_6[1]));
	jspl3 jspl3_w_n1562_21(.douta(w_n1562_21[0]),.doutb(w_n1562_21[1]),.doutc(w_n1562_21[2]),.din(w_n1562_6[2]));
	jspl3 jspl3_w_n1562_22(.douta(w_n1562_22[0]),.doutb(w_n1562_22[1]),.doutc(w_n1562_22[2]),.din(w_n1562_7[0]));
	jspl3 jspl3_w_n1562_23(.douta(w_n1562_23[0]),.doutb(w_n1562_23[1]),.doutc(w_n1562_23[2]),.din(w_n1562_7[1]));
	jspl3 jspl3_w_n1562_24(.douta(w_n1562_24[0]),.doutb(w_n1562_24[1]),.doutc(w_n1562_24[2]),.din(w_n1562_7[2]));
	jspl3 jspl3_w_n1562_25(.douta(w_n1562_25[0]),.doutb(w_n1562_25[1]),.doutc(w_n1562_25[2]),.din(w_n1562_8[0]));
	jspl3 jspl3_w_n1562_26(.douta(w_n1562_26[0]),.doutb(w_n1562_26[1]),.doutc(w_n1562_26[2]),.din(w_n1562_8[1]));
	jspl3 jspl3_w_n1562_27(.douta(w_n1562_27[0]),.doutb(w_n1562_27[1]),.doutc(w_n1562_27[2]),.din(w_n1562_8[2]));
	jspl3 jspl3_w_n1562_28(.douta(w_n1562_28[0]),.doutb(w_n1562_28[1]),.doutc(w_n1562_28[2]),.din(w_n1562_9[0]));
	jspl3 jspl3_w_n1562_29(.douta(w_n1562_29[0]),.doutb(w_n1562_29[1]),.doutc(w_n1562_29[2]),.din(w_n1562_9[1]));
	jspl3 jspl3_w_n1562_30(.douta(w_n1562_30[0]),.doutb(w_n1562_30[1]),.doutc(w_n1562_30[2]),.din(w_n1562_9[2]));
	jspl3 jspl3_w_n1562_31(.douta(w_n1562_31[0]),.doutb(w_n1562_31[1]),.doutc(w_n1562_31[2]),.din(w_n1562_10[0]));
	jspl3 jspl3_w_n1562_32(.douta(w_n1562_32[0]),.doutb(w_n1562_32[1]),.doutc(w_n1562_32[2]),.din(w_n1562_10[1]));
	jspl3 jspl3_w_n1562_33(.douta(w_n1562_33[0]),.doutb(w_n1562_33[1]),.doutc(w_n1562_33[2]),.din(w_n1562_10[2]));
	jspl3 jspl3_w_n1562_34(.douta(w_n1562_34[0]),.doutb(w_n1562_34[1]),.doutc(w_n1562_34[2]),.din(w_n1562_11[0]));
	jspl3 jspl3_w_n1562_35(.douta(w_n1562_35[0]),.doutb(w_n1562_35[1]),.doutc(w_n1562_35[2]),.din(w_n1562_11[1]));
	jspl3 jspl3_w_n1562_36(.douta(w_n1562_36[0]),.doutb(w_n1562_36[1]),.doutc(w_n1562_36[2]),.din(w_n1562_11[2]));
	jspl3 jspl3_w_n1562_37(.douta(w_n1562_37[0]),.doutb(w_n1562_37[1]),.doutc(w_n1562_37[2]),.din(w_n1562_12[0]));
	jspl3 jspl3_w_n1562_38(.douta(w_n1562_38[0]),.doutb(w_n1562_38[1]),.doutc(w_n1562_38[2]),.din(w_n1562_12[1]));
	jspl3 jspl3_w_n1562_39(.douta(w_n1562_39[0]),.doutb(w_n1562_39[1]),.doutc(w_n1562_39[2]),.din(w_n1562_12[2]));
	jspl3 jspl3_w_n1562_40(.douta(w_n1562_40[0]),.doutb(w_n1562_40[1]),.doutc(w_n1562_40[2]),.din(w_n1562_13[0]));
	jspl3 jspl3_w_n1562_41(.douta(w_n1562_41[0]),.doutb(w_n1562_41[1]),.doutc(w_n1562_41[2]),.din(w_n1562_13[1]));
	jspl3 jspl3_w_n1562_42(.douta(w_n1562_42[0]),.doutb(w_n1562_42[1]),.doutc(w_n1562_42[2]),.din(w_n1562_13[2]));
	jspl3 jspl3_w_n1562_43(.douta(w_n1562_43[0]),.doutb(w_n1562_43[1]),.doutc(w_n1562_43[2]),.din(w_n1562_14[0]));
	jspl3 jspl3_w_n1562_44(.douta(w_n1562_44[0]),.doutb(w_n1562_44[1]),.doutc(w_n1562_44[2]),.din(w_n1562_14[1]));
	jspl3 jspl3_w_n1562_45(.douta(w_n1562_45[0]),.doutb(w_n1562_45[1]),.doutc(w_n1562_45[2]),.din(w_n1562_14[2]));
	jspl3 jspl3_w_n1562_46(.douta(w_n1562_46[0]),.doutb(w_n1562_46[1]),.doutc(w_n1562_46[2]),.din(w_n1562_15[0]));
	jspl3 jspl3_w_n1562_47(.douta(w_n1562_47[0]),.doutb(w_n1562_47[1]),.doutc(w_n1562_47[2]),.din(w_n1562_15[1]));
	jspl3 jspl3_w_n1562_48(.douta(w_n1562_48[0]),.doutb(w_n1562_48[1]),.doutc(w_n1562_48[2]),.din(w_n1562_15[2]));
	jspl3 jspl3_w_n1562_49(.douta(w_n1562_49[0]),.doutb(w_n1562_49[1]),.doutc(w_n1562_49[2]),.din(w_n1562_16[0]));
	jspl3 jspl3_w_n1562_50(.douta(w_n1562_50[0]),.doutb(w_n1562_50[1]),.doutc(w_n1562_50[2]),.din(w_n1562_16[1]));
	jspl3 jspl3_w_n1562_51(.douta(w_n1562_51[0]),.doutb(w_n1562_51[1]),.doutc(w_n1562_51[2]),.din(w_n1562_16[2]));
	jspl3 jspl3_w_n1562_52(.douta(w_n1562_52[0]),.doutb(w_n1562_52[1]),.doutc(w_n1562_52[2]),.din(w_n1562_17[0]));
	jspl3 jspl3_w_n1562_53(.douta(w_n1562_53[0]),.doutb(w_n1562_53[1]),.doutc(w_n1562_53[2]),.din(w_n1562_17[1]));
	jspl3 jspl3_w_n1562_54(.douta(w_n1562_54[0]),.doutb(w_n1562_54[1]),.doutc(w_n1562_54[2]),.din(w_n1562_17[2]));
	jspl3 jspl3_w_n1562_55(.douta(w_n1562_55[0]),.doutb(w_n1562_55[1]),.doutc(w_n1562_55[2]),.din(w_n1562_18[0]));
	jspl3 jspl3_w_n1562_56(.douta(w_n1562_56[0]),.doutb(w_n1562_56[1]),.doutc(w_n1562_56[2]),.din(w_n1562_18[1]));
	jspl3 jspl3_w_n1562_57(.douta(w_n1562_57[0]),.doutb(w_n1562_57[1]),.doutc(w_n1562_57[2]),.din(w_n1562_18[2]));
	jspl3 jspl3_w_n1562_58(.douta(w_n1562_58[0]),.doutb(w_n1562_58[1]),.doutc(w_n1562_58[2]),.din(w_n1562_19[0]));
	jspl3 jspl3_w_n1562_59(.douta(w_n1562_59[0]),.doutb(w_n1562_59[1]),.doutc(w_n1562_59[2]),.din(w_n1562_19[1]));
	jspl3 jspl3_w_n1562_60(.douta(w_n1562_60[0]),.doutb(w_n1562_60[1]),.doutc(w_n1562_60[2]),.din(w_n1562_19[2]));
	jspl3 jspl3_w_n1562_61(.douta(w_n1562_61[0]),.doutb(w_n1562_61[1]),.doutc(w_n1562_61[2]),.din(w_n1562_20[0]));
	jspl3 jspl3_w_n1562_62(.douta(w_n1562_62[0]),.doutb(w_n1562_62[1]),.doutc(w_n1562_62[2]),.din(w_n1562_20[1]));
	jspl3 jspl3_w_n1562_63(.douta(w_n1562_63[0]),.doutb(w_n1562_63[1]),.doutc(w_n1562_63[2]),.din(w_n1562_20[2]));
	jspl3 jspl3_w_n1562_64(.douta(w_n1562_64[0]),.doutb(w_n1562_64[1]),.doutc(w_n1562_64[2]),.din(w_n1562_21[0]));
	jspl3 jspl3_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.doutc(w_n1586_0[2]),.din(n1586));
	jspl jspl_w_n1588_0(.douta(w_n1588_0[0]),.doutb(w_n1588_0[1]),.din(n1588));
	jspl3 jspl3_w_n1721_0(.douta(w_n1721_0[0]),.doutb(w_n1721_0[1]),.doutc(w_n1721_0[2]),.din(n1721));
	jspl3 jspl3_w_n1721_1(.douta(w_n1721_1[0]),.doutb(w_n1721_1[1]),.doutc(w_n1721_1[2]),.din(w_n1721_0[0]));
	jspl3 jspl3_w_n1721_2(.douta(w_n1721_2[0]),.doutb(w_n1721_2[1]),.doutc(w_n1721_2[2]),.din(w_n1721_0[1]));
	jspl3 jspl3_w_n1721_3(.douta(w_n1721_3[0]),.doutb(w_n1721_3[1]),.doutc(w_n1721_3[2]),.din(w_n1721_0[2]));
	jspl3 jspl3_w_n1721_4(.douta(w_n1721_4[0]),.doutb(w_n1721_4[1]),.doutc(w_n1721_4[2]),.din(w_n1721_1[0]));
	jspl3 jspl3_w_n1721_5(.douta(w_n1721_5[0]),.doutb(w_n1721_5[1]),.doutc(w_n1721_5[2]),.din(w_n1721_1[1]));
	jspl3 jspl3_w_n1721_6(.douta(w_n1721_6[0]),.doutb(w_n1721_6[1]),.doutc(w_n1721_6[2]),.din(w_n1721_1[2]));
	jspl3 jspl3_w_n1721_7(.douta(w_n1721_7[0]),.doutb(w_n1721_7[1]),.doutc(w_n1721_7[2]),.din(w_n1721_2[0]));
	jspl3 jspl3_w_n1721_8(.douta(w_n1721_8[0]),.doutb(w_n1721_8[1]),.doutc(w_n1721_8[2]),.din(w_n1721_2[1]));
	jspl3 jspl3_w_n1721_9(.douta(w_n1721_9[0]),.doutb(w_n1721_9[1]),.doutc(w_n1721_9[2]),.din(w_n1721_2[2]));
	jspl3 jspl3_w_n1721_10(.douta(w_n1721_10[0]),.doutb(w_n1721_10[1]),.doutc(w_n1721_10[2]),.din(w_n1721_3[0]));
	jspl3 jspl3_w_n1721_11(.douta(w_n1721_11[0]),.doutb(w_n1721_11[1]),.doutc(w_n1721_11[2]),.din(w_n1721_3[1]));
	jspl3 jspl3_w_n1721_12(.douta(w_n1721_12[0]),.doutb(w_n1721_12[1]),.doutc(w_n1721_12[2]),.din(w_n1721_3[2]));
	jspl3 jspl3_w_n1721_13(.douta(w_n1721_13[0]),.doutb(w_n1721_13[1]),.doutc(w_n1721_13[2]),.din(w_n1721_4[0]));
	jspl3 jspl3_w_n1721_14(.douta(w_n1721_14[0]),.doutb(w_n1721_14[1]),.doutc(w_n1721_14[2]),.din(w_n1721_4[1]));
	jspl3 jspl3_w_n1721_15(.douta(w_n1721_15[0]),.doutb(w_n1721_15[1]),.doutc(w_n1721_15[2]),.din(w_n1721_4[2]));
	jspl3 jspl3_w_n1721_16(.douta(w_n1721_16[0]),.doutb(w_n1721_16[1]),.doutc(w_n1721_16[2]),.din(w_n1721_5[0]));
	jspl3 jspl3_w_n1721_17(.douta(w_n1721_17[0]),.doutb(w_n1721_17[1]),.doutc(w_n1721_17[2]),.din(w_n1721_5[1]));
	jspl3 jspl3_w_n1721_18(.douta(w_n1721_18[0]),.doutb(w_n1721_18[1]),.doutc(w_n1721_18[2]),.din(w_n1721_5[2]));
	jspl3 jspl3_w_n1721_19(.douta(w_n1721_19[0]),.doutb(w_n1721_19[1]),.doutc(w_n1721_19[2]),.din(w_n1721_6[0]));
	jspl3 jspl3_w_n1721_20(.douta(w_n1721_20[0]),.doutb(w_n1721_20[1]),.doutc(w_n1721_20[2]),.din(w_n1721_6[1]));
	jspl3 jspl3_w_n1721_21(.douta(w_n1721_21[0]),.doutb(w_n1721_21[1]),.doutc(w_n1721_21[2]),.din(w_n1721_6[2]));
	jspl3 jspl3_w_n1721_22(.douta(w_n1721_22[0]),.doutb(w_n1721_22[1]),.doutc(w_n1721_22[2]),.din(w_n1721_7[0]));
	jspl3 jspl3_w_n1721_23(.douta(w_n1721_23[0]),.doutb(w_n1721_23[1]),.doutc(w_n1721_23[2]),.din(w_n1721_7[1]));
	jspl3 jspl3_w_n1721_24(.douta(w_n1721_24[0]),.doutb(w_n1721_24[1]),.doutc(w_n1721_24[2]),.din(w_n1721_7[2]));
	jspl3 jspl3_w_n1721_25(.douta(w_n1721_25[0]),.doutb(w_n1721_25[1]),.doutc(w_n1721_25[2]),.din(w_n1721_8[0]));
	jspl3 jspl3_w_n1721_26(.douta(w_n1721_26[0]),.doutb(w_n1721_26[1]),.doutc(w_n1721_26[2]),.din(w_n1721_8[1]));
	jspl3 jspl3_w_n1721_27(.douta(w_n1721_27[0]),.doutb(w_n1721_27[1]),.doutc(w_n1721_27[2]),.din(w_n1721_8[2]));
	jspl3 jspl3_w_n1721_28(.douta(w_n1721_28[0]),.doutb(w_n1721_28[1]),.doutc(w_n1721_28[2]),.din(w_n1721_9[0]));
	jspl3 jspl3_w_n1721_29(.douta(w_n1721_29[0]),.doutb(w_n1721_29[1]),.doutc(w_n1721_29[2]),.din(w_n1721_9[1]));
	jspl3 jspl3_w_n1721_30(.douta(w_n1721_30[0]),.doutb(w_n1721_30[1]),.doutc(w_n1721_30[2]),.din(w_n1721_9[2]));
	jspl3 jspl3_w_n1721_31(.douta(w_n1721_31[0]),.doutb(w_n1721_31[1]),.doutc(w_n1721_31[2]),.din(w_n1721_10[0]));
	jspl3 jspl3_w_n1721_32(.douta(w_n1721_32[0]),.doutb(w_n1721_32[1]),.doutc(w_n1721_32[2]),.din(w_n1721_10[1]));
	jspl3 jspl3_w_n1721_33(.douta(w_n1721_33[0]),.doutb(w_n1721_33[1]),.doutc(w_n1721_33[2]),.din(w_n1721_10[2]));
	jspl3 jspl3_w_n1721_34(.douta(w_n1721_34[0]),.doutb(w_n1721_34[1]),.doutc(w_n1721_34[2]),.din(w_n1721_11[0]));
	jspl3 jspl3_w_n1721_35(.douta(w_n1721_35[0]),.doutb(w_n1721_35[1]),.doutc(w_n1721_35[2]),.din(w_n1721_11[1]));
	jspl3 jspl3_w_n1721_36(.douta(w_n1721_36[0]),.doutb(w_n1721_36[1]),.doutc(w_n1721_36[2]),.din(w_n1721_11[2]));
	jspl3 jspl3_w_n1721_37(.douta(w_n1721_37[0]),.doutb(w_n1721_37[1]),.doutc(w_n1721_37[2]),.din(w_n1721_12[0]));
	jspl3 jspl3_w_n1721_38(.douta(w_n1721_38[0]),.doutb(w_n1721_38[1]),.doutc(w_n1721_38[2]),.din(w_n1721_12[1]));
	jspl3 jspl3_w_n1721_39(.douta(w_n1721_39[0]),.doutb(w_n1721_39[1]),.doutc(w_n1721_39[2]),.din(w_n1721_12[2]));
	jspl3 jspl3_w_n1721_40(.douta(w_n1721_40[0]),.doutb(w_n1721_40[1]),.doutc(w_n1721_40[2]),.din(w_n1721_13[0]));
	jspl3 jspl3_w_n1721_41(.douta(w_n1721_41[0]),.doutb(w_n1721_41[1]),.doutc(w_n1721_41[2]),.din(w_n1721_13[1]));
	jspl3 jspl3_w_n1721_42(.douta(w_n1721_42[0]),.doutb(w_n1721_42[1]),.doutc(w_n1721_42[2]),.din(w_n1721_13[2]));
	jspl3 jspl3_w_n1721_43(.douta(w_n1721_43[0]),.doutb(w_n1721_43[1]),.doutc(w_n1721_43[2]),.din(w_n1721_14[0]));
	jspl3 jspl3_w_n1721_44(.douta(w_n1721_44[0]),.doutb(w_n1721_44[1]),.doutc(w_n1721_44[2]),.din(w_n1721_14[1]));
	jspl3 jspl3_w_n1721_45(.douta(w_n1721_45[0]),.doutb(w_n1721_45[1]),.doutc(w_n1721_45[2]),.din(w_n1721_14[2]));
	jspl3 jspl3_w_n1721_46(.douta(w_n1721_46[0]),.doutb(w_n1721_46[1]),.doutc(w_n1721_46[2]),.din(w_n1721_15[0]));
	jspl3 jspl3_w_n1721_47(.douta(w_n1721_47[0]),.doutb(w_n1721_47[1]),.doutc(w_n1721_47[2]),.din(w_n1721_15[1]));
	jspl3 jspl3_w_n1721_48(.douta(w_n1721_48[0]),.doutb(w_n1721_48[1]),.doutc(w_n1721_48[2]),.din(w_n1721_15[2]));
	jspl3 jspl3_w_n1721_49(.douta(w_n1721_49[0]),.doutb(w_n1721_49[1]),.doutc(w_n1721_49[2]),.din(w_n1721_16[0]));
	jspl3 jspl3_w_n1721_50(.douta(w_n1721_50[0]),.doutb(w_n1721_50[1]),.doutc(w_n1721_50[2]),.din(w_n1721_16[1]));
	jspl3 jspl3_w_n1721_51(.douta(w_n1721_51[0]),.doutb(w_n1721_51[1]),.doutc(w_n1721_51[2]),.din(w_n1721_16[2]));
	jspl3 jspl3_w_n1721_52(.douta(w_n1721_52[0]),.doutb(w_n1721_52[1]),.doutc(w_n1721_52[2]),.din(w_n1721_17[0]));
	jspl3 jspl3_w_n1721_53(.douta(w_n1721_53[0]),.doutb(w_n1721_53[1]),.doutc(w_n1721_53[2]),.din(w_n1721_17[1]));
	jspl3 jspl3_w_n1721_54(.douta(w_n1721_54[0]),.doutb(w_n1721_54[1]),.doutc(w_n1721_54[2]),.din(w_n1721_17[2]));
	jspl3 jspl3_w_n1721_55(.douta(w_n1721_55[0]),.doutb(w_n1721_55[1]),.doutc(w_n1721_55[2]),.din(w_n1721_18[0]));
	jspl3 jspl3_w_n1721_56(.douta(w_n1721_56[0]),.doutb(w_n1721_56[1]),.doutc(w_n1721_56[2]),.din(w_n1721_18[1]));
	jspl3 jspl3_w_n1721_57(.douta(w_n1721_57[0]),.doutb(w_n1721_57[1]),.doutc(w_n1721_57[2]),.din(w_n1721_18[2]));
	jspl3 jspl3_w_n1721_58(.douta(w_n1721_58[0]),.doutb(w_n1721_58[1]),.doutc(w_n1721_58[2]),.din(w_n1721_19[0]));
	jspl3 jspl3_w_n1721_59(.douta(w_n1721_59[0]),.doutb(w_n1721_59[1]),.doutc(w_n1721_59[2]),.din(w_n1721_19[1]));
	jspl3 jspl3_w_n1721_60(.douta(w_n1721_60[0]),.doutb(w_n1721_60[1]),.doutc(w_n1721_60[2]),.din(w_n1721_19[2]));
	jspl3 jspl3_w_n1721_61(.douta(w_n1721_61[0]),.doutb(w_n1721_61[1]),.doutc(w_n1721_61[2]),.din(w_n1721_20[0]));
	jspl3 jspl3_w_n1721_62(.douta(w_n1721_62[0]),.doutb(w_n1721_62[1]),.doutc(w_n1721_62[2]),.din(w_n1721_20[1]));
	jspl3 jspl3_w_n1721_63(.douta(w_n1721_63[0]),.doutb(w_n1721_63[1]),.doutc(w_n1721_63[2]),.din(w_n1721_20[2]));
	jspl3 jspl3_w_n1721_64(.douta(w_n1721_64[0]),.doutb(w_n1721_64[1]),.doutc(w_n1721_64[2]),.din(w_n1721_21[0]));
	jspl jspl_w_n1721_65(.douta(w_n1721_65[0]),.doutb(w_n1721_65[1]),.din(w_n1721_21[1]));
	jspl jspl_w_n1723_0(.douta(w_n1723_0[0]),.doutb(w_n1723_0[1]),.din(n1723));
	jspl jspl_w_n1724_0(.douta(w_n1724_0[0]),.doutb(w_n1724_0[1]),.din(n1724));
	jspl jspl_w_n1726_0(.douta(w_n1726_0[0]),.doutb(w_n1726_0[1]),.din(n1726));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_n1728_0[1]),.din(n1728));
	jspl jspl_w_n1730_0(.douta(w_n1730_0[0]),.doutb(w_n1730_0[1]),.din(n1730));
	jspl jspl_w_n1732_0(.douta(w_n1732_0[0]),.doutb(w_n1732_0[1]),.din(n1732));
	jspl jspl_w_n1736_0(.douta(w_n1736_0[0]),.doutb(w_n1736_0[1]),.din(n1736));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(n1738));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(n1740));
	jspl jspl_w_n1741_0(.douta(w_n1741_0[0]),.doutb(w_n1741_0[1]),.din(n1741));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(n1743));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(n1745));
	jspl jspl_w_n1746_0(.douta(w_n1746_0[0]),.doutb(w_n1746_0[1]),.din(n1746));
	jspl jspl_w_n1747_0(.douta(w_n1747_0[0]),.doutb(w_n1747_0[1]),.din(n1747));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1759_0(.douta(w_n1759_0[0]),.doutb(w_n1759_0[1]),.din(n1759));
	jspl jspl_w_n1761_0(.douta(w_n1761_0[0]),.doutb(w_n1761_0[1]),.din(n1761));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.din(n1767));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_n1768_0[1]),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(n1770));
	jspl jspl_w_n1771_0(.douta(w_n1771_0[0]),.doutb(w_n1771_0[1]),.din(n1771));
	jspl jspl_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.din(n1772));
	jspl jspl_w_n1774_0(.douta(w_n1774_0[0]),.doutb(w_n1774_0[1]),.din(n1774));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(n1775));
	jspl jspl_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.din(n1777));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(n1778));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(n1779));
	jspl jspl_w_n1782_0(.douta(w_n1782_0[0]),.doutb(w_n1782_0[1]),.din(n1782));
	jspl jspl_w_n1784_0(.douta(w_n1784_0[0]),.doutb(w_n1784_0[1]),.din(n1784));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.din(n1786));
	jspl jspl_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_n1791_0[1]),.din(n1791));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1797_0(.douta(w_n1797_0[0]),.doutb(w_n1797_0[1]),.din(n1797));
	jspl jspl_w_n1799_0(.douta(w_n1799_0[0]),.doutb(w_n1799_0[1]),.din(n1799));
	jspl jspl_w_n1800_0(.douta(w_n1800_0[0]),.doutb(w_n1800_0[1]),.din(n1800));
	jspl jspl_w_n1802_0(.douta(w_n1802_0[0]),.doutb(w_n1802_0[1]),.din(n1802));
	jspl jspl_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.din(n1804));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_n1805_0[1]),.din(n1805));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(n1806));
	jspl jspl_w_n1809_0(.douta(w_n1809_0[0]),.doutb(w_n1809_0[1]),.din(n1809));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1818_0(.douta(w_n1818_0[0]),.doutb(w_n1818_0[1]),.din(n1818));
	jspl jspl_w_n1820_0(.douta(w_n1820_0[0]),.doutb(w_n1820_0[1]),.din(n1820));
	jspl jspl_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.din(n1824));
	jspl jspl_w_n1826_0(.douta(w_n1826_0[0]),.doutb(w_n1826_0[1]),.din(n1826));
	jspl jspl_w_n1827_0(.douta(w_n1827_0[0]),.doutb(w_n1827_0[1]),.din(n1827));
	jspl jspl_w_n1829_0(.douta(w_n1829_0[0]),.doutb(w_n1829_0[1]),.din(n1829));
	jspl jspl_w_n1830_0(.douta(w_n1830_0[0]),.doutb(w_n1830_0[1]),.din(n1830));
	jspl jspl_w_n1831_0(.douta(w_n1831_0[0]),.doutb(w_n1831_0[1]),.din(n1831));
	jspl jspl_w_n1833_0(.douta(w_n1833_0[0]),.doutb(w_n1833_0[1]),.din(n1833));
	jspl jspl_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.din(n1834));
	jspl jspl_w_n1836_0(.douta(w_n1836_0[0]),.doutb(w_n1836_0[1]),.din(n1836));
	jspl jspl_w_n1837_0(.douta(w_n1837_0[0]),.doutb(w_n1837_0[1]),.din(n1837));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(n1838));
	jspl jspl_w_n1841_0(.douta(w_n1841_0[0]),.doutb(w_n1841_0[1]),.din(n1841));
	jspl jspl_w_n1843_0(.douta(w_n1843_0[0]),.doutb(w_n1843_0[1]),.din(n1843));
	jspl jspl_w_n1845_0(.douta(w_n1845_0[0]),.doutb(w_n1845_0[1]),.din(n1845));
	jspl jspl_w_n1850_0(.douta(w_n1850_0[0]),.doutb(w_n1850_0[1]),.din(n1850));
	jspl jspl_w_n1852_0(.douta(w_n1852_0[0]),.doutb(w_n1852_0[1]),.din(n1852));
	jspl jspl_w_n1856_0(.douta(w_n1856_0[0]),.doutb(w_n1856_0[1]),.din(n1856));
	jspl jspl_w_n1858_0(.douta(w_n1858_0[0]),.doutb(w_n1858_0[1]),.din(n1858));
	jspl jspl_w_n1859_0(.douta(w_n1859_0[0]),.doutb(w_n1859_0[1]),.din(n1859));
	jspl jspl_w_n1861_0(.douta(w_n1861_0[0]),.doutb(w_n1861_0[1]),.din(n1861));
	jspl jspl_w_n1863_0(.douta(w_n1863_0[0]),.doutb(w_n1863_0[1]),.din(n1863));
	jspl jspl_w_n1864_0(.douta(w_n1864_0[0]),.doutb(w_n1864_0[1]),.din(n1864));
	jspl jspl_w_n1865_0(.douta(w_n1865_0[0]),.doutb(w_n1865_0[1]),.din(n1865));
	jspl jspl_w_n1868_0(.douta(w_n1868_0[0]),.doutb(w_n1868_0[1]),.din(n1868));
	jspl jspl_w_n1870_0(.douta(w_n1870_0[0]),.doutb(w_n1870_0[1]),.din(n1870));
	jspl jspl_w_n1872_0(.douta(w_n1872_0[0]),.doutb(w_n1872_0[1]),.din(n1872));
	jspl jspl_w_n1877_0(.douta(w_n1877_0[0]),.doutb(w_n1877_0[1]),.din(n1877));
	jspl jspl_w_n1879_0(.douta(w_n1879_0[0]),.doutb(w_n1879_0[1]),.din(n1879));
	jspl jspl_w_n1883_0(.douta(w_n1883_0[0]),.doutb(w_n1883_0[1]),.din(n1883));
	jspl jspl_w_n1885_0(.douta(w_n1885_0[0]),.doutb(w_n1885_0[1]),.din(n1885));
	jspl jspl_w_n1886_0(.douta(w_n1886_0[0]),.doutb(w_n1886_0[1]),.din(n1886));
	jspl jspl_w_n1888_0(.douta(w_n1888_0[0]),.doutb(w_n1888_0[1]),.din(n1888));
	jspl jspl_w_n1889_0(.douta(w_n1889_0[0]),.doutb(w_n1889_0[1]),.din(n1889));
	jspl jspl_w_n1890_0(.douta(w_n1890_0[0]),.doutb(w_n1890_0[1]),.din(n1890));
	jspl jspl_w_n1892_0(.douta(w_n1892_0[0]),.doutb(w_n1892_0[1]),.din(n1892));
	jspl jspl_w_n1893_0(.douta(w_n1893_0[0]),.doutb(w_n1893_0[1]),.din(n1893));
	jspl jspl_w_n1895_0(.douta(w_n1895_0[0]),.doutb(w_n1895_0[1]),.din(n1895));
	jspl jspl_w_n1896_0(.douta(w_n1896_0[0]),.doutb(w_n1896_0[1]),.din(n1896));
	jspl jspl_w_n1897_0(.douta(w_n1897_0[0]),.doutb(w_n1897_0[1]),.din(n1897));
	jspl jspl_w_n1900_0(.douta(w_n1900_0[0]),.doutb(w_n1900_0[1]),.din(n1900));
	jspl jspl_w_n1902_0(.douta(w_n1902_0[0]),.doutb(w_n1902_0[1]),.din(n1902));
	jspl jspl_w_n1904_0(.douta(w_n1904_0[0]),.doutb(w_n1904_0[1]),.din(n1904));
	jspl jspl_w_n1909_0(.douta(w_n1909_0[0]),.doutb(w_n1909_0[1]),.din(n1909));
	jspl jspl_w_n1911_0(.douta(w_n1911_0[0]),.doutb(w_n1911_0[1]),.din(n1911));
	jspl jspl_w_n1915_0(.douta(w_n1915_0[0]),.doutb(w_n1915_0[1]),.din(n1915));
	jspl jspl_w_n1917_0(.douta(w_n1917_0[0]),.doutb(w_n1917_0[1]),.din(n1917));
	jspl jspl_w_n1918_0(.douta(w_n1918_0[0]),.doutb(w_n1918_0[1]),.din(n1918));
	jspl jspl_w_n1920_0(.douta(w_n1920_0[0]),.doutb(w_n1920_0[1]),.din(n1920));
	jspl jspl_w_n1922_0(.douta(w_n1922_0[0]),.doutb(w_n1922_0[1]),.din(n1922));
	jspl jspl_w_n1923_0(.douta(w_n1923_0[0]),.doutb(w_n1923_0[1]),.din(n1923));
	jspl jspl_w_n1924_0(.douta(w_n1924_0[0]),.doutb(w_n1924_0[1]),.din(n1924));
	jspl jspl_w_n1927_0(.douta(w_n1927_0[0]),.doutb(w_n1927_0[1]),.din(n1927));
	jspl jspl_w_n1929_0(.douta(w_n1929_0[0]),.doutb(w_n1929_0[1]),.din(n1929));
	jspl jspl_w_n1931_0(.douta(w_n1931_0[0]),.doutb(w_n1931_0[1]),.din(n1931));
	jspl jspl_w_n1936_0(.douta(w_n1936_0[0]),.doutb(w_n1936_0[1]),.din(n1936));
	jspl jspl_w_n1938_0(.douta(w_n1938_0[0]),.doutb(w_n1938_0[1]),.din(n1938));
	jspl jspl_w_n1942_0(.douta(w_n1942_0[0]),.doutb(w_n1942_0[1]),.din(n1942));
	jspl jspl_w_n1944_0(.douta(w_n1944_0[0]),.doutb(w_n1944_0[1]),.din(n1944));
	jspl jspl_w_n1945_0(.douta(w_n1945_0[0]),.doutb(w_n1945_0[1]),.din(n1945));
	jspl jspl_w_n1947_0(.douta(w_n1947_0[0]),.doutb(w_n1947_0[1]),.din(n1947));
	jspl jspl_w_n1948_0(.douta(w_n1948_0[0]),.doutb(w_n1948_0[1]),.din(n1948));
	jspl jspl_w_n1950_0(.douta(w_n1950_0[0]),.doutb(w_n1950_0[1]),.din(n1950));
	jspl jspl_w_n1953_0(.douta(w_n1953_0[0]),.doutb(w_n1953_0[1]),.din(n1953));
	jspl jspl_w_n1955_0(.douta(w_n1955_0[0]),.doutb(w_n1955_0[1]),.din(n1955));
	jspl jspl_w_n1958_0(.douta(w_n1958_0[0]),.doutb(w_n1958_0[1]),.din(n1958));
	jspl jspl_w_n1960_0(.douta(w_n1960_0[0]),.doutb(w_n1960_0[1]),.din(n1960));
	jspl jspl_w_n1961_0(.douta(w_n1961_0[0]),.doutb(w_n1961_0[1]),.din(n1961));
	jspl jspl_w_n1963_0(.douta(w_n1963_0[0]),.doutb(w_n1963_0[1]),.din(n1963));
	jspl jspl_w_n1964_0(.douta(w_n1964_0[0]),.doutb(w_n1964_0[1]),.din(n1964));
	jspl jspl_w_n1965_0(.douta(w_n1965_0[0]),.doutb(w_n1965_0[1]),.din(n1965));
	jspl jspl_w_n1967_0(.douta(w_n1967_0[0]),.doutb(w_n1967_0[1]),.din(n1967));
	jspl jspl_w_n1970_0(.douta(w_n1970_0[0]),.doutb(w_n1970_0[1]),.din(n1970));
	jspl jspl_w_n1971_0(.douta(w_n1971_0[0]),.doutb(w_n1971_0[1]),.din(n1971));
	jspl jspl_w_n1974_0(.douta(w_n1974_0[0]),.doutb(w_n1974_0[1]),.din(n1974));
	jspl jspl_w_n1976_0(.douta(w_n1976_0[0]),.doutb(w_n1976_0[1]),.din(n1976));
	jspl jspl_w_n1977_0(.douta(w_n1977_0[0]),.doutb(w_n1977_0[1]),.din(n1977));
	jspl jspl_w_n1978_0(.douta(w_n1978_0[0]),.doutb(w_n1978_0[1]),.din(n1978));
	jspl jspl_w_n1979_0(.douta(w_n1979_0[0]),.doutb(w_n1979_0[1]),.din(n1979));
	jspl jspl_w_n1981_0(.douta(w_n1981_0[0]),.doutb(w_n1981_0[1]),.din(n1981));
	jspl jspl_w_n1983_0(.douta(w_n1983_0[0]),.doutb(w_n1983_0[1]),.din(n1983));
	jspl jspl_w_n1984_0(.douta(w_n1984_0[0]),.doutb(w_n1984_0[1]),.din(n1984));
	jspl jspl_w_n1987_0(.douta(w_n1987_0[0]),.doutb(w_n1987_0[1]),.din(n1987));
	jspl jspl_w_n1990_0(.douta(w_n1990_0[0]),.doutb(w_n1990_0[1]),.din(n1990));
	jspl jspl_w_n1992_0(.douta(w_n1992_0[0]),.doutb(w_n1992_0[1]),.din(n1992));
	jspl jspl_w_n1993_0(.douta(w_n1993_0[0]),.doutb(w_n1993_0[1]),.din(n1993));
	jspl jspl_w_n1995_0(.douta(w_n1995_0[0]),.doutb(w_n1995_0[1]),.din(n1995));
	jspl jspl_w_n1996_0(.douta(w_n1996_0[0]),.doutb(w_n1996_0[1]),.din(n1996));
	jspl jspl_w_n1997_0(.douta(w_n1997_0[0]),.doutb(w_n1997_0[1]),.din(n1997));
	jspl jspl_w_n1999_0(.douta(w_n1999_0[0]),.doutb(w_n1999_0[1]),.din(n1999));
	jspl jspl_w_n2002_0(.douta(w_n2002_0[0]),.doutb(w_n2002_0[1]),.din(n2002));
	jspl jspl_w_n2003_0(.douta(w_n2003_0[0]),.doutb(w_n2003_0[1]),.din(n2003));
	jspl jspl_w_n2006_0(.douta(w_n2006_0[0]),.doutb(w_n2006_0[1]),.din(n2006));
	jspl jspl_w_n2008_0(.douta(w_n2008_0[0]),.doutb(w_n2008_0[1]),.din(n2008));
	jspl jspl_w_n2010_0(.douta(w_n2010_0[0]),.doutb(w_n2010_0[1]),.din(n2010));
	jspl jspl_w_n2013_0(.douta(w_n2013_0[0]),.doutb(w_n2013_0[1]),.din(n2013));
	jspl jspl_w_n2014_0(.douta(w_n2014_0[0]),.doutb(w_n2014_0[1]),.din(n2014));
	jspl jspl_w_n2016_0(.douta(w_n2016_0[0]),.doutb(w_n2016_0[1]),.din(n2016));
	jspl jspl_w_n2020_0(.douta(w_n2020_0[0]),.doutb(w_n2020_0[1]),.din(n2020));
	jspl jspl_w_n2022_0(.douta(w_n2022_0[0]),.doutb(w_n2022_0[1]),.din(n2022));
	jspl jspl_w_n2025_0(.douta(w_n2025_0[0]),.doutb(w_n2025_0[1]),.din(n2025));
	jspl jspl_w_n2027_0(.douta(w_n2027_0[0]),.doutb(w_n2027_0[1]),.din(n2027));
	jspl jspl_w_n2029_0(.douta(w_n2029_0[0]),.doutb(w_n2029_0[1]),.din(n2029));
	jspl jspl_w_n2030_0(.douta(w_n2030_0[0]),.doutb(w_n2030_0[1]),.din(n2030));
	jspl jspl_w_n2031_0(.douta(w_n2031_0[0]),.doutb(w_n2031_0[1]),.din(n2031));
	jspl jspl_w_n2034_0(.douta(w_n2034_0[0]),.doutb(w_n2034_0[1]),.din(n2034));
	jspl jspl_w_n2035_0(.douta(w_n2035_0[0]),.doutb(w_n2035_0[1]),.din(n2035));
	jspl jspl_w_n2036_0(.douta(w_n2036_0[0]),.doutb(w_n2036_0[1]),.din(n2036));
	jspl jspl_w_n2038_0(.douta(w_n2038_0[0]),.doutb(w_n2038_0[1]),.din(n2038));
	jspl jspl_w_n2040_0(.douta(w_n2040_0[0]),.doutb(w_n2040_0[1]),.din(n2040));
	jspl jspl_w_n2041_0(.douta(w_n2041_0[0]),.doutb(w_n2041_0[1]),.din(n2041));
	jspl jspl_w_n2042_0(.douta(w_n2042_0[0]),.doutb(w_n2042_0[1]),.din(n2042));
	jspl jspl_w_n2043_0(.douta(w_n2043_0[0]),.doutb(w_n2043_0[1]),.din(n2043));
	jspl jspl_w_n2045_0(.douta(w_n2045_0[0]),.doutb(w_n2045_0[1]),.din(n2045));
	jspl jspl_w_n2046_0(.douta(w_n2046_0[0]),.doutb(w_n2046_0[1]),.din(n2046));
	jspl jspl_w_n2047_0(.douta(w_n2047_0[0]),.doutb(w_n2047_0[1]),.din(n2047));
	jspl jspl_w_n2048_0(.douta(w_n2048_0[0]),.doutb(w_n2048_0[1]),.din(n2048));
	jspl jspl_w_n2050_0(.douta(w_n2050_0[0]),.doutb(w_n2050_0[1]),.din(n2050));
	jspl jspl_w_n2051_0(.douta(w_n2051_0[0]),.doutb(w_n2051_0[1]),.din(n2051));
	jspl jspl_w_n2052_0(.douta(w_n2052_0[0]),.doutb(w_n2052_0[1]),.din(n2052));
	jspl jspl_w_n2053_0(.douta(w_n2053_0[0]),.doutb(w_n2053_0[1]),.din(n2053));
	jspl jspl_w_n2055_0(.douta(w_n2055_0[0]),.doutb(w_n2055_0[1]),.din(n2055));
	jspl jspl_w_n2056_0(.douta(w_n2056_0[0]),.doutb(w_n2056_0[1]),.din(n2056));
	jspl jspl_w_n2057_0(.douta(w_n2057_0[0]),.doutb(w_n2057_0[1]),.din(n2057));
	jspl jspl_w_n2058_0(.douta(w_n2058_0[0]),.doutb(w_n2058_0[1]),.din(n2058));
	jspl jspl_w_n2060_0(.douta(w_n2060_0[0]),.doutb(w_n2060_0[1]),.din(n2060));
	jspl jspl_w_n2061_0(.douta(w_n2061_0[0]),.doutb(w_n2061_0[1]),.din(n2061));
	jspl jspl_w_n2062_0(.douta(w_n2062_0[0]),.doutb(w_n2062_0[1]),.din(n2062));
	jspl jspl_w_n2063_0(.douta(w_n2063_0[0]),.doutb(w_n2063_0[1]),.din(n2063));
	jspl jspl_w_n2064_0(.douta(w_n2064_0[0]),.doutb(w_n2064_0[1]),.din(n2064));
	jspl jspl_w_n2065_0(.douta(w_n2065_0[0]),.doutb(w_n2065_0[1]),.din(n2065));
	jspl jspl_w_n2067_0(.douta(w_n2067_0[0]),.doutb(w_n2067_0[1]),.din(n2067));
	jspl jspl_w_n2068_0(.douta(w_n2068_0[0]),.doutb(w_n2068_0[1]),.din(n2068));
	jspl jspl_w_n2069_0(.douta(w_n2069_0[0]),.doutb(w_n2069_0[1]),.din(n2069));
	jspl jspl_w_n2070_0(.douta(w_n2070_0[0]),.doutb(w_n2070_0[1]),.din(n2070));
	jspl jspl_w_n2072_0(.douta(w_n2072_0[0]),.doutb(w_n2072_0[1]),.din(n2072));
	jspl jspl_w_n2073_0(.douta(w_n2073_0[0]),.doutb(w_n2073_0[1]),.din(n2073));
	jspl jspl_w_n2074_0(.douta(w_n2074_0[0]),.doutb(w_n2074_0[1]),.din(n2074));
	jspl jspl_w_n2075_0(.douta(w_n2075_0[0]),.doutb(w_n2075_0[1]),.din(n2075));
	jspl jspl_w_n2077_0(.douta(w_n2077_0[0]),.doutb(w_n2077_0[1]),.din(n2077));
	jspl jspl_w_n2078_0(.douta(w_n2078_0[0]),.doutb(w_n2078_0[1]),.din(n2078));
	jspl jspl_w_n2079_0(.douta(w_n2079_0[0]),.doutb(w_n2079_0[1]),.din(n2079));
	jspl jspl_w_n2080_0(.douta(w_n2080_0[0]),.doutb(w_n2080_0[1]),.din(n2080));
	jspl jspl_w_n2082_0(.douta(w_n2082_0[0]),.doutb(w_n2082_0[1]),.din(n2082));
	jspl jspl_w_n2083_0(.douta(w_n2083_0[0]),.doutb(w_n2083_0[1]),.din(n2083));
	jspl jspl_w_n2084_0(.douta(w_n2084_0[0]),.doutb(w_n2084_0[1]),.din(n2084));
	jspl jspl_w_n2085_0(.douta(w_n2085_0[0]),.doutb(w_n2085_0[1]),.din(n2085));
	jspl jspl_w_n2086_0(.douta(w_n2086_0[0]),.doutb(w_n2086_0[1]),.din(n2086));
	jspl jspl_w_n2087_0(.douta(w_n2087_0[0]),.doutb(w_n2087_0[1]),.din(n2087));
	jspl jspl_w_n2089_0(.douta(w_n2089_0[0]),.doutb(w_n2089_0[1]),.din(n2089));
	jspl jspl_w_n2090_0(.douta(w_n2090_0[0]),.doutb(w_n2090_0[1]),.din(n2090));
	jspl jspl_w_n2091_0(.douta(w_n2091_0[0]),.doutb(w_n2091_0[1]),.din(n2091));
	jspl jspl_w_n2092_0(.douta(w_n2092_0[0]),.doutb(w_n2092_0[1]),.din(n2092));
	jspl jspl_w_n2094_0(.douta(w_n2094_0[0]),.doutb(w_n2094_0[1]),.din(n2094));
	jspl jspl_w_n2095_0(.douta(w_n2095_0[0]),.doutb(w_n2095_0[1]),.din(n2095));
	jspl jspl_w_n2096_0(.douta(w_n2096_0[0]),.doutb(w_n2096_0[1]),.din(n2096));
	jspl jspl_w_n2097_0(.douta(w_n2097_0[0]),.doutb(w_n2097_0[1]),.din(n2097));
	jspl jspl_w_n2099_0(.douta(w_n2099_0[0]),.doutb(w_n2099_0[1]),.din(n2099));
	jspl jspl_w_n2100_0(.douta(w_n2100_0[0]),.doutb(w_n2100_0[1]),.din(n2100));
	jspl jspl_w_n2101_0(.douta(w_n2101_0[0]),.doutb(w_n2101_0[1]),.din(n2101));
	jspl jspl_w_n2102_0(.douta(w_n2102_0[0]),.doutb(w_n2102_0[1]),.din(n2102));
	jspl jspl_w_n2104_0(.douta(w_n2104_0[0]),.doutb(w_n2104_0[1]),.din(n2104));
	jspl jspl_w_n2105_0(.douta(w_n2105_0[0]),.doutb(w_n2105_0[1]),.din(n2105));
	jspl jspl_w_n2106_0(.douta(w_n2106_0[0]),.doutb(w_n2106_0[1]),.din(n2106));
	jspl jspl_w_n2107_0(.douta(w_n2107_0[0]),.doutb(w_n2107_0[1]),.din(n2107));
	jspl jspl_w_n2108_0(.douta(w_n2108_0[0]),.doutb(w_n2108_0[1]),.din(n2108));
	jspl jspl_w_n2109_0(.douta(w_n2109_0[0]),.doutb(w_n2109_0[1]),.din(n2109));
	jspl3 jspl3_w_n2110_0(.douta(w_n2110_0[0]),.doutb(w_n2110_0[1]),.doutc(w_n2110_0[2]),.din(n2110));
	jspl jspl_w_n2111_0(.douta(w_n2111_0[0]),.doutb(w_n2111_0[1]),.din(n2111));
	jspl jspl_w_n2113_0(.douta(w_n2113_0[0]),.doutb(w_n2113_0[1]),.din(n2113));
	jspl jspl_w_n2115_0(.douta(w_n2115_0[0]),.doutb(w_n2115_0[1]),.din(n2115));
	jspl jspl_w_n2120_0(.douta(w_n2120_0[0]),.doutb(w_n2120_0[1]),.din(n2120));
	jspl jspl_w_n2122_0(.douta(w_n2122_0[0]),.doutb(w_n2122_0[1]),.din(n2122));
	jspl jspl_w_n2124_0(.douta(w_n2124_0[0]),.doutb(w_n2124_0[1]),.din(n2124));
	jspl jspl_w_n2127_0(.douta(w_n2127_0[0]),.doutb(w_n2127_0[1]),.din(n2127));
	jspl jspl_w_n2128_0(.douta(w_n2128_0[0]),.doutb(w_n2128_0[1]),.din(n2128));
	jspl jspl_w_n2131_0(.douta(w_n2131_0[0]),.doutb(w_n2131_0[1]),.din(n2131));
	jspl jspl_w_n2133_0(.douta(w_n2133_0[0]),.doutb(w_n2133_0[1]),.din(n2133));
	jspl jspl_w_n2135_0(.douta(w_n2135_0[0]),.doutb(w_n2135_0[1]),.din(n2135));
	jspl jspl_w_n2138_0(.douta(w_n2138_0[0]),.doutb(w_n2138_0[1]),.din(n2138));
	jspl jspl_w_n2140_0(.douta(w_n2140_0[0]),.doutb(w_n2140_0[1]),.din(n2140));
	jspl jspl_w_n2142_0(.douta(w_n2142_0[0]),.doutb(w_n2142_0[1]),.din(n2142));
	jspl jspl_w_n2144_0(.douta(w_n2144_0[0]),.doutb(w_n2144_0[1]),.din(n2144));
	jspl jspl_w_n2146_0(.douta(w_n2146_0[0]),.doutb(w_n2146_0[1]),.din(n2146));
	jspl jspl_w_n2148_0(.douta(w_n2148_0[0]),.doutb(w_n2148_0[1]),.din(n2148));
	jspl jspl_w_n2151_0(.douta(w_n2151_0[0]),.doutb(w_n2151_0[1]),.din(n2151));
	jspl jspl_w_n2152_0(.douta(w_n2152_0[0]),.doutb(w_n2152_0[1]),.din(n2152));
	jspl jspl_w_n2155_0(.douta(w_n2155_0[0]),.doutb(w_n2155_0[1]),.din(n2155));
	jspl jspl_w_n2157_0(.douta(w_n2157_0[0]),.doutb(w_n2157_0[1]),.din(n2157));
	jspl jspl_w_n2159_0(.douta(w_n2159_0[0]),.doutb(w_n2159_0[1]),.din(n2159));
	jspl jspl_w_n2162_0(.douta(w_n2162_0[0]),.doutb(w_n2162_0[1]),.din(n2162));
	jspl jspl_w_n2164_0(.douta(w_n2164_0[0]),.doutb(w_n2164_0[1]),.din(n2164));
	jspl jspl_w_n2166_0(.douta(w_n2166_0[0]),.doutb(w_n2166_0[1]),.din(n2166));
	jspl jspl_w_n2176_0(.douta(w_n2176_0[0]),.doutb(w_n2176_0[1]),.din(n2176));
	jspl jspl_w_n2178_0(.douta(w_n2178_0[0]),.doutb(w_n2178_0[1]),.din(n2178));
	jspl jspl_w_n2180_0(.douta(w_n2180_0[0]),.doutb(w_n2180_0[1]),.din(n2180));
	jspl jspl_w_n2183_0(.douta(w_n2183_0[0]),.doutb(w_n2183_0[1]),.din(n2183));
	jspl jspl_w_n2184_0(.douta(w_n2184_0[0]),.doutb(w_n2184_0[1]),.din(n2184));
	jspl jspl_w_n2187_0(.douta(w_n2187_0[0]),.doutb(w_n2187_0[1]),.din(n2187));
	jspl jspl_w_n2189_0(.douta(w_n2189_0[0]),.doutb(w_n2189_0[1]),.din(n2189));
	jspl jspl_w_n2191_0(.douta(w_n2191_0[0]),.doutb(w_n2191_0[1]),.din(n2191));
	jspl jspl_w_n2194_0(.douta(w_n2194_0[0]),.doutb(w_n2194_0[1]),.din(n2194));
	jspl jspl_w_n2196_0(.douta(w_n2196_0[0]),.doutb(w_n2196_0[1]),.din(n2196));
	jspl jspl_w_n2198_0(.douta(w_n2198_0[0]),.doutb(w_n2198_0[1]),.din(n2198));
	jspl jspl_w_n2208_0(.douta(w_n2208_0[0]),.doutb(w_n2208_0[1]),.din(n2208));
	jspl jspl_w_n2210_0(.douta(w_n2210_0[0]),.doutb(w_n2210_0[1]),.din(n2210));
	jspl jspl_w_n2212_0(.douta(w_n2212_0[0]),.doutb(w_n2212_0[1]),.din(n2212));
	jspl jspl_w_n2215_0(.douta(w_n2215_0[0]),.doutb(w_n2215_0[1]),.din(n2215));
	jspl jspl_w_n2216_0(.douta(w_n2216_0[0]),.doutb(w_n2216_0[1]),.din(n2216));
	jspl jspl_w_n2219_0(.douta(w_n2219_0[0]),.doutb(w_n2219_0[1]),.din(n2219));
	jspl jspl_w_n2221_0(.douta(w_n2221_0[0]),.doutb(w_n2221_0[1]),.din(n2221));
	jspl jspl_w_n2223_0(.douta(w_n2223_0[0]),.doutb(w_n2223_0[1]),.din(n2223));
	jspl jspl_w_n2226_0(.douta(w_n2226_0[0]),.doutb(w_n2226_0[1]),.din(n2226));
	jspl jspl_w_n2228_0(.douta(w_n2228_0[0]),.doutb(w_n2228_0[1]),.din(n2228));
	jspl jspl_w_n2230_0(.douta(w_n2230_0[0]),.doutb(w_n2230_0[1]),.din(n2230));
	jspl jspl_w_n2240_0(.douta(w_n2240_0[0]),.doutb(w_n2240_0[1]),.din(n2240));
	jspl jspl_w_n2242_0(.douta(w_n2242_0[0]),.doutb(w_n2242_0[1]),.din(n2242));
	jspl jspl_w_n2244_0(.douta(w_n2244_0[0]),.doutb(w_n2244_0[1]),.din(n2244));
	jspl jspl_w_n2247_0(.douta(w_n2247_0[0]),.doutb(w_n2247_0[1]),.din(n2247));
	jspl jspl_w_n2249_0(.douta(w_n2249_0[0]),.doutb(w_n2249_0[1]),.din(n2249));
	jspl jspl_w_n2253_0(.douta(w_n2253_0[0]),.doutb(w_n2253_0[1]),.din(n2253));
	jspl jspl_w_n2256_0(.douta(w_n2256_0[0]),.doutb(w_n2256_0[1]),.din(n2256));
	jspl jspl_w_n2258_0(.douta(w_n2258_0[0]),.doutb(w_n2258_0[1]),.din(n2258));
	jspl jspl_w_n2263_0(.douta(w_n2263_0[0]),.doutb(w_n2263_0[1]),.din(n2263));
	jspl jspl_w_n2266_0(.douta(w_n2266_0[0]),.doutb(w_n2266_0[1]),.din(n2266));
	jspl jspl_w_n2269_0(.douta(w_n2269_0[0]),.doutb(w_n2269_0[1]),.din(n2269));
	jspl jspl_w_n2274_0(.douta(w_n2274_0[0]),.doutb(w_n2274_0[1]),.din(n2274));
	jspl jspl_w_n2278_0(.douta(w_n2278_0[0]),.doutb(w_n2278_0[1]),.din(n2278));
	jspl jspl_w_n2281_0(.douta(w_n2281_0[0]),.doutb(w_n2281_0[1]),.din(n2281));
	jspl jspl_w_n2283_0(.douta(w_n2283_0[0]),.doutb(w_n2283_0[1]),.din(n2283));
	jspl jspl_w_n2284_0(.douta(w_n2284_0[0]),.doutb(w_n2284_0[1]),.din(n2284));
	jspl jspl_w_n2286_0(.douta(w_n2286_0[0]),.doutb(w_n2286_0[1]),.din(n2286));
	jspl jspl_w_n2290_0(.douta(w_n2290_0[0]),.doutb(w_n2290_0[1]),.din(n2290));
	jspl jspl_w_n2292_0(.douta(w_n2292_0[0]),.doutb(w_n2292_0[1]),.din(n2292));
	jspl jspl_w_n2295_0(.douta(w_n2295_0[0]),.doutb(w_n2295_0[1]),.din(n2295));
	jspl jspl_w_n2297_0(.douta(w_n2297_0[0]),.doutb(w_n2297_0[1]),.din(n2297));
	jspl jspl_w_n2300_0(.douta(w_n2300_0[0]),.doutb(w_n2300_0[1]),.din(n2300));
	jspl jspl_w_n2306_0(.douta(w_n2306_0[0]),.doutb(w_n2306_0[1]),.din(n2306));
	jspl jspl_w_n2308_0(.douta(w_n2308_0[0]),.doutb(w_n2308_0[1]),.din(n2308));
	jspl jspl_w_n2313_0(.douta(w_n2313_0[0]),.doutb(w_n2313_0[1]),.din(n2313));
	jspl jspl_w_n2315_0(.douta(w_n2315_0[0]),.doutb(w_n2315_0[1]),.din(n2315));
	jspl jspl_w_n2320_0(.douta(w_n2320_0[0]),.doutb(w_n2320_0[1]),.din(n2320));
	jspl jspl_w_n2324_0(.douta(w_n2324_0[0]),.doutb(w_n2324_0[1]),.din(n2324));
	jspl jspl_w_n2327_0(.douta(w_n2327_0[0]),.doutb(w_n2327_0[1]),.din(n2327));
	jspl jspl_w_n2329_0(.douta(w_n2329_0[0]),.doutb(w_n2329_0[1]),.din(n2329));
	jspl jspl_w_n2330_0(.douta(w_n2330_0[0]),.doutb(w_n2330_0[1]),.din(n2330));
	jspl jspl_w_n2332_0(.douta(w_n2332_0[0]),.doutb(w_n2332_0[1]),.din(n2332));
	jspl jspl_w_n2336_0(.douta(w_n2336_0[0]),.doutb(w_n2336_0[1]),.din(n2336));
	jspl jspl_w_n2338_0(.douta(w_n2338_0[0]),.doutb(w_n2338_0[1]),.din(n2338));
	jspl jspl_w_n2341_0(.douta(w_n2341_0[0]),.doutb(w_n2341_0[1]),.din(n2341));
	jspl jspl_w_n2343_0(.douta(w_n2343_0[0]),.doutb(w_n2343_0[1]),.din(n2343));
	jspl jspl_w_n2346_0(.douta(w_n2346_0[0]),.doutb(w_n2346_0[1]),.din(n2346));
	jspl jspl_w_n2351_0(.douta(w_n2351_0[0]),.doutb(w_n2351_0[1]),.din(n2351));
	jspl jspl_w_n2355_0(.douta(w_n2355_0[0]),.doutb(w_n2355_0[1]),.din(n2355));
	jspl jspl_w_n2358_0(.douta(w_n2358_0[0]),.doutb(w_n2358_0[1]),.din(n2358));
	jspl jspl_w_n2360_0(.douta(w_n2360_0[0]),.doutb(w_n2360_0[1]),.din(n2360));
	jspl jspl_w_n2366_0(.douta(w_n2366_0[0]),.doutb(w_n2366_0[1]),.din(n2366));
	jspl jspl_w_n2370_0(.douta(w_n2370_0[0]),.doutb(w_n2370_0[1]),.din(n2370));
	jspl jspl_w_n2373_0(.douta(w_n2373_0[0]),.doutb(w_n2373_0[1]),.din(n2373));
	jspl jspl_w_n2375_0(.douta(w_n2375_0[0]),.doutb(w_n2375_0[1]),.din(n2375));
	jspl jspl_w_n2376_0(.douta(w_n2376_0[0]),.doutb(w_n2376_0[1]),.din(n2376));
	jspl jspl_w_n2378_0(.douta(w_n2378_0[0]),.doutb(w_n2378_0[1]),.din(n2378));
	jspl jspl_w_n2382_0(.douta(w_n2382_0[0]),.doutb(w_n2382_0[1]),.din(n2382));
	jspl jspl_w_n2384_0(.douta(w_n2384_0[0]),.doutb(w_n2384_0[1]),.din(n2384));
	jspl jspl_w_n2387_0(.douta(w_n2387_0[0]),.doutb(w_n2387_0[1]),.din(n2387));
	jspl jspl_w_n2389_0(.douta(w_n2389_0[0]),.doutb(w_n2389_0[1]),.din(n2389));
	jspl jspl_w_n2392_0(.douta(w_n2392_0[0]),.doutb(w_n2392_0[1]),.din(n2392));
	jspl jspl_w_n2398_0(.douta(w_n2398_0[0]),.doutb(w_n2398_0[1]),.din(n2398));
	jspl jspl_w_n2400_0(.douta(w_n2400_0[0]),.doutb(w_n2400_0[1]),.din(n2400));
	jspl jspl_w_n2405_0(.douta(w_n2405_0[0]),.doutb(w_n2405_0[1]),.din(n2405));
	jspl jspl_w_n2407_0(.douta(w_n2407_0[0]),.doutb(w_n2407_0[1]),.din(n2407));
	jspl jspl_w_n2412_0(.douta(w_n2412_0[0]),.doutb(w_n2412_0[1]),.din(n2412));
	jspl jspl_w_n2416_0(.douta(w_n2416_0[0]),.doutb(w_n2416_0[1]),.din(n2416));
	jspl jspl_w_n2418_0(.douta(w_n2418_0[0]),.doutb(w_n2418_0[1]),.din(n2418));
	jspl jspl_w_n2421_0(.douta(w_n2421_0[0]),.doutb(w_n2421_0[1]),.din(n2421));
	jspl jspl_w_n2423_0(.douta(w_n2423_0[0]),.doutb(w_n2423_0[1]),.din(n2423));
	jspl jspl_w_n2425_0(.douta(w_n2425_0[0]),.doutb(w_n2425_0[1]),.din(n2425));
	jspl jspl_w_n2428_0(.douta(w_n2428_0[0]),.doutb(w_n2428_0[1]),.din(n2428));
	jspl jspl_w_n2430_0(.douta(w_n2430_0[0]),.doutb(w_n2430_0[1]),.din(n2430));
	jspl jspl_w_n2433_0(.douta(w_n2433_0[0]),.doutb(w_n2433_0[1]),.din(n2433));
	jspl jspl_w_n2435_0(.douta(w_n2435_0[0]),.doutb(w_n2435_0[1]),.din(n2435));
	jspl jspl_w_n2437_0(.douta(w_n2437_0[0]),.doutb(w_n2437_0[1]),.din(n2437));
	jspl jspl_w_n2438_0(.douta(w_n2438_0[0]),.doutb(w_n2438_0[1]),.din(n2438));
	jspl jspl_w_n2440_0(.douta(w_n2440_0[0]),.doutb(w_n2440_0[1]),.din(n2440));
	jspl jspl_w_n2441_0(.douta(w_n2441_0[0]),.doutb(w_n2441_0[1]),.din(n2441));
	jspl jspl_w_n2443_0(.douta(w_n2443_0[0]),.doutb(w_n2443_0[1]),.din(n2443));
	jspl jspl_w_n2446_0(.douta(w_n2446_0[0]),.doutb(w_n2446_0[1]),.din(n2446));
	jspl jspl_w_n2448_0(.douta(w_n2448_0[0]),.doutb(w_n2448_0[1]),.din(n2448));
	jspl jspl_w_n2452_0(.douta(w_n2452_0[0]),.doutb(w_n2452_0[1]),.din(n2452));
	jspl jspl_w_n2456_0(.douta(w_n2456_0[0]),.doutb(w_n2456_0[1]),.din(n2456));
	jspl jspl_w_n2460_0(.douta(w_n2460_0[0]),.doutb(w_n2460_0[1]),.din(n2460));
	jspl jspl_w_n2462_0(.douta(w_n2462_0[0]),.doutb(w_n2462_0[1]),.din(n2462));
	jspl jspl_w_n2465_0(.douta(w_n2465_0[0]),.doutb(w_n2465_0[1]),.din(n2465));
	jspl jspl_w_n2467_0(.douta(w_n2467_0[0]),.doutb(w_n2467_0[1]),.din(n2467));
	jspl jspl_w_n2469_0(.douta(w_n2469_0[0]),.doutb(w_n2469_0[1]),.din(n2469));
	jspl jspl_w_n2472_0(.douta(w_n2472_0[0]),.doutb(w_n2472_0[1]),.din(n2472));
	jspl jspl_w_n2473_0(.douta(w_n2473_0[0]),.doutb(w_n2473_0[1]),.din(n2473));
	jspl jspl_w_n2475_0(.douta(w_n2475_0[0]),.doutb(w_n2475_0[1]),.din(n2475));
	jspl jspl_w_n2479_0(.douta(w_n2479_0[0]),.doutb(w_n2479_0[1]),.din(n2479));
	jspl jspl_w_n2483_0(.douta(w_n2483_0[0]),.doutb(w_n2483_0[1]),.din(n2483));
	jspl jspl_w_n2487_0(.douta(w_n2487_0[0]),.doutb(w_n2487_0[1]),.din(n2487));
	jspl jspl_w_n2489_0(.douta(w_n2489_0[0]),.doutb(w_n2489_0[1]),.din(n2489));
	jspl jspl_w_n2492_0(.douta(w_n2492_0[0]),.doutb(w_n2492_0[1]),.din(n2492));
	jspl jspl_w_n2494_0(.douta(w_n2494_0[0]),.doutb(w_n2494_0[1]),.din(n2494));
	jspl jspl_w_n2496_0(.douta(w_n2496_0[0]),.doutb(w_n2496_0[1]),.din(n2496));
	jspl jspl_w_n2497_0(.douta(w_n2497_0[0]),.doutb(w_n2497_0[1]),.din(n2497));
	jspl jspl_w_n2499_0(.douta(w_n2499_0[0]),.doutb(w_n2499_0[1]),.din(n2499));
	jspl jspl_w_n2500_0(.douta(w_n2500_0[0]),.doutb(w_n2500_0[1]),.din(n2500));
	jspl jspl_w_n2502_0(.douta(w_n2502_0[0]),.doutb(w_n2502_0[1]),.din(n2502));
	jspl jspl_w_n2505_0(.douta(w_n2505_0[0]),.doutb(w_n2505_0[1]),.din(n2505));
	jspl jspl_w_n2507_0(.douta(w_n2507_0[0]),.doutb(w_n2507_0[1]),.din(n2507));
	jspl jspl_w_n2511_0(.douta(w_n2511_0[0]),.doutb(w_n2511_0[1]),.din(n2511));
	jspl jspl_w_n2515_0(.douta(w_n2515_0[0]),.doutb(w_n2515_0[1]),.din(n2515));
	jspl jspl_w_n2519_0(.douta(w_n2519_0[0]),.doutb(w_n2519_0[1]),.din(n2519));
	jspl jspl_w_n2521_0(.douta(w_n2521_0[0]),.doutb(w_n2521_0[1]),.din(n2521));
	jspl jspl_w_n2524_0(.douta(w_n2524_0[0]),.doutb(w_n2524_0[1]),.din(n2524));
	jspl jspl_w_n2526_0(.douta(w_n2526_0[0]),.doutb(w_n2526_0[1]),.din(n2526));
	jspl jspl_w_n2528_0(.douta(w_n2528_0[0]),.doutb(w_n2528_0[1]),.din(n2528));
	jspl jspl_w_n2531_0(.douta(w_n2531_0[0]),.doutb(w_n2531_0[1]),.din(n2531));
	jspl jspl_w_n2532_0(.douta(w_n2532_0[0]),.doutb(w_n2532_0[1]),.din(n2532));
	jspl jspl_w_n2534_0(.douta(w_n2534_0[0]),.doutb(w_n2534_0[1]),.din(n2534));
	jspl jspl_w_n2538_0(.douta(w_n2538_0[0]),.doutb(w_n2538_0[1]),.din(n2538));
	jspl jspl_w_n2542_0(.douta(w_n2542_0[0]),.doutb(w_n2542_0[1]),.din(n2542));
	jspl jspl_w_n2546_0(.douta(w_n2546_0[0]),.doutb(w_n2546_0[1]),.din(n2546));
	jspl jspl_w_n2548_0(.douta(w_n2548_0[0]),.doutb(w_n2548_0[1]),.din(n2548));
	jspl jspl_w_n2551_0(.douta(w_n2551_0[0]),.doutb(w_n2551_0[1]),.din(n2551));
	jspl jspl_w_n2553_0(.douta(w_n2553_0[0]),.doutb(w_n2553_0[1]),.din(n2553));
	jspl jspl_w_n2555_0(.douta(w_n2555_0[0]),.doutb(w_n2555_0[1]),.din(n2555));
	jspl jspl_w_n2556_0(.douta(w_n2556_0[0]),.doutb(w_n2556_0[1]),.din(n2556));
	jspl jspl_w_n2558_0(.douta(w_n2558_0[0]),.doutb(w_n2558_0[1]),.din(n2558));
	jspl jspl_w_n2559_0(.douta(w_n2559_0[0]),.doutb(w_n2559_0[1]),.din(n2559));
	jspl jspl_w_n2561_0(.douta(w_n2561_0[0]),.doutb(w_n2561_0[1]),.din(n2561));
	jspl jspl_w_n2564_0(.douta(w_n2564_0[0]),.doutb(w_n2564_0[1]),.din(n2564));
	jspl jspl_w_n2566_0(.douta(w_n2566_0[0]),.doutb(w_n2566_0[1]),.din(n2566));
	jspl jspl_w_n2570_0(.douta(w_n2570_0[0]),.doutb(w_n2570_0[1]),.din(n2570));
	jspl jspl_w_n2574_0(.douta(w_n2574_0[0]),.doutb(w_n2574_0[1]),.din(n2574));
	jspl jspl_w_n2578_0(.douta(w_n2578_0[0]),.doutb(w_n2578_0[1]),.din(n2578));
	jspl jspl_w_n2580_0(.douta(w_n2580_0[0]),.doutb(w_n2580_0[1]),.din(n2580));
	jspl jspl_w_n2583_0(.douta(w_n2583_0[0]),.doutb(w_n2583_0[1]),.din(n2583));
	jspl jspl_w_n2585_0(.douta(w_n2585_0[0]),.doutb(w_n2585_0[1]),.din(n2585));
	jspl jspl_w_n2587_0(.douta(w_n2587_0[0]),.doutb(w_n2587_0[1]),.din(n2587));
	jspl jspl_w_n2590_0(.douta(w_n2590_0[0]),.doutb(w_n2590_0[1]),.din(n2590));
	jspl jspl_w_n2591_0(.douta(w_n2591_0[0]),.doutb(w_n2591_0[1]),.din(n2591));
	jspl jspl_w_n2593_0(.douta(w_n2593_0[0]),.doutb(w_n2593_0[1]),.din(n2593));
	jspl jspl_w_n2597_0(.douta(w_n2597_0[0]),.doutb(w_n2597_0[1]),.din(n2597));
	jspl jspl_w_n2601_0(.douta(w_n2601_0[0]),.doutb(w_n2601_0[1]),.din(n2601));
	jspl jspl_w_n2605_0(.douta(w_n2605_0[0]),.doutb(w_n2605_0[1]),.din(n2605));
	jspl jspl_w_n2607_0(.douta(w_n2607_0[0]),.doutb(w_n2607_0[1]),.din(n2607));
	jspl jspl_w_n2610_0(.douta(w_n2610_0[0]),.doutb(w_n2610_0[1]),.din(n2610));
	jspl jspl_w_n2612_0(.douta(w_n2612_0[0]),.doutb(w_n2612_0[1]),.din(n2612));
	jspl jspl_w_n2614_0(.douta(w_n2614_0[0]),.doutb(w_n2614_0[1]),.din(n2614));
	jspl jspl_w_n2615_0(.douta(w_n2615_0[0]),.doutb(w_n2615_0[1]),.din(n2615));
	jspl jspl_w_n2617_0(.douta(w_n2617_0[0]),.doutb(w_n2617_0[1]),.din(n2617));
	jspl jspl_w_n2618_0(.douta(w_n2618_0[0]),.doutb(w_n2618_0[1]),.din(n2618));
	jspl jspl_w_n2620_0(.douta(w_n2620_0[0]),.doutb(w_n2620_0[1]),.din(n2620));
	jspl jspl_w_n2623_0(.douta(w_n2623_0[0]),.doutb(w_n2623_0[1]),.din(n2623));
	jspl jspl_w_n2625_0(.douta(w_n2625_0[0]),.doutb(w_n2625_0[1]),.din(n2625));
	jspl jspl_w_n2629_0(.douta(w_n2629_0[0]),.doutb(w_n2629_0[1]),.din(n2629));
	jspl jspl_w_n2633_0(.douta(w_n2633_0[0]),.doutb(w_n2633_0[1]),.din(n2633));
	jspl jspl_w_n2637_0(.douta(w_n2637_0[0]),.doutb(w_n2637_0[1]),.din(n2637));
	jspl jspl_w_n2639_0(.douta(w_n2639_0[0]),.doutb(w_n2639_0[1]),.din(n2639));
	jspl3 jspl3_w_n2641_0(.douta(w_n2641_0[0]),.doutb(w_n2641_0[1]),.doutc(w_n2641_0[2]),.din(n2641));
	jspl jspl_w_n2642_0(.douta(w_n2642_0[0]),.doutb(w_n2642_0[1]),.din(n2642));
	jspl3 jspl3_w_n2643_0(.douta(w_n2643_0[0]),.doutb(w_n2643_0[1]),.doutc(w_n2643_0[2]),.din(n2643));
	jspl jspl_w_n2643_1(.douta(w_n2643_1[0]),.doutb(w_n2643_1[1]),.din(w_n2643_0[0]));
	jspl jspl_w_n2644_0(.douta(w_n2644_0[0]),.doutb(w_n2644_0[1]),.din(n2644));
	jspl jspl_w_n2647_0(.douta(w_n2647_0[0]),.doutb(w_n2647_0[1]),.din(n2647));
	jspl jspl_w_n2648_0(.douta(w_n2648_0[0]),.doutb(w_n2648_0[1]),.din(n2648));
	jspl jspl_w_n2649_0(.douta(w_n2649_0[0]),.doutb(w_n2649_0[1]),.din(n2649));
	jspl jspl_w_n2672_0(.douta(w_n2672_0[0]),.doutb(w_n2672_0[1]),.din(n2672));
	jspl jspl_w_n2801_0(.douta(w_n2801_0[0]),.doutb(w_n2801_0[1]),.din(n2801));
	jspl3 jspl3_w_n2803_0(.douta(w_n2803_0[0]),.doutb(w_n2803_0[1]),.doutc(w_n2803_0[2]),.din(n2803));
	jspl3 jspl3_w_n2803_1(.douta(w_n2803_1[0]),.doutb(w_n2803_1[1]),.doutc(w_n2803_1[2]),.din(w_n2803_0[0]));
	jspl3 jspl3_w_n2803_2(.douta(w_n2803_2[0]),.doutb(w_n2803_2[1]),.doutc(w_n2803_2[2]),.din(w_n2803_0[1]));
	jspl3 jspl3_w_n2803_3(.douta(w_n2803_3[0]),.doutb(w_n2803_3[1]),.doutc(w_n2803_3[2]),.din(w_n2803_0[2]));
	jspl3 jspl3_w_n2803_4(.douta(w_n2803_4[0]),.doutb(w_n2803_4[1]),.doutc(w_n2803_4[2]),.din(w_n2803_1[0]));
	jspl3 jspl3_w_n2803_5(.douta(w_n2803_5[0]),.doutb(w_n2803_5[1]),.doutc(w_n2803_5[2]),.din(w_n2803_1[1]));
	jspl3 jspl3_w_n2803_6(.douta(w_n2803_6[0]),.doutb(w_n2803_6[1]),.doutc(w_n2803_6[2]),.din(w_n2803_1[2]));
	jspl3 jspl3_w_n2803_7(.douta(w_n2803_7[0]),.doutb(w_n2803_7[1]),.doutc(w_n2803_7[2]),.din(w_n2803_2[0]));
	jspl3 jspl3_w_n2803_8(.douta(w_n2803_8[0]),.doutb(w_n2803_8[1]),.doutc(w_n2803_8[2]),.din(w_n2803_2[1]));
	jspl3 jspl3_w_n2803_9(.douta(w_n2803_9[0]),.doutb(w_n2803_9[1]),.doutc(w_n2803_9[2]),.din(w_n2803_2[2]));
	jspl3 jspl3_w_n2803_10(.douta(w_n2803_10[0]),.doutb(w_n2803_10[1]),.doutc(w_n2803_10[2]),.din(w_n2803_3[0]));
	jspl3 jspl3_w_n2803_11(.douta(w_n2803_11[0]),.doutb(w_n2803_11[1]),.doutc(w_n2803_11[2]),.din(w_n2803_3[1]));
	jspl3 jspl3_w_n2803_12(.douta(w_n2803_12[0]),.doutb(w_n2803_12[1]),.doutc(w_n2803_12[2]),.din(w_n2803_3[2]));
	jspl3 jspl3_w_n2803_13(.douta(w_n2803_13[0]),.doutb(w_n2803_13[1]),.doutc(w_n2803_13[2]),.din(w_n2803_4[0]));
	jspl3 jspl3_w_n2803_14(.douta(w_n2803_14[0]),.doutb(w_n2803_14[1]),.doutc(w_n2803_14[2]),.din(w_n2803_4[1]));
	jspl3 jspl3_w_n2803_15(.douta(w_n2803_15[0]),.doutb(w_n2803_15[1]),.doutc(w_n2803_15[2]),.din(w_n2803_4[2]));
	jspl3 jspl3_w_n2803_16(.douta(w_n2803_16[0]),.doutb(w_n2803_16[1]),.doutc(w_n2803_16[2]),.din(w_n2803_5[0]));
	jspl3 jspl3_w_n2803_17(.douta(w_n2803_17[0]),.doutb(w_n2803_17[1]),.doutc(w_n2803_17[2]),.din(w_n2803_5[1]));
	jspl3 jspl3_w_n2803_18(.douta(w_n2803_18[0]),.doutb(w_n2803_18[1]),.doutc(w_n2803_18[2]),.din(w_n2803_5[2]));
	jspl3 jspl3_w_n2803_19(.douta(w_n2803_19[0]),.doutb(w_n2803_19[1]),.doutc(w_n2803_19[2]),.din(w_n2803_6[0]));
	jspl3 jspl3_w_n2803_20(.douta(w_n2803_20[0]),.doutb(w_n2803_20[1]),.doutc(w_n2803_20[2]),.din(w_n2803_6[1]));
	jspl3 jspl3_w_n2803_21(.douta(w_n2803_21[0]),.doutb(w_n2803_21[1]),.doutc(w_n2803_21[2]),.din(w_n2803_6[2]));
	jspl3 jspl3_w_n2803_22(.douta(w_n2803_22[0]),.doutb(w_n2803_22[1]),.doutc(w_n2803_22[2]),.din(w_n2803_7[0]));
	jspl3 jspl3_w_n2803_23(.douta(w_n2803_23[0]),.doutb(w_n2803_23[1]),.doutc(w_n2803_23[2]),.din(w_n2803_7[1]));
	jspl3 jspl3_w_n2803_24(.douta(w_n2803_24[0]),.doutb(w_n2803_24[1]),.doutc(w_n2803_24[2]),.din(w_n2803_7[2]));
	jspl3 jspl3_w_n2803_25(.douta(w_n2803_25[0]),.doutb(w_n2803_25[1]),.doutc(w_n2803_25[2]),.din(w_n2803_8[0]));
	jspl3 jspl3_w_n2803_26(.douta(w_n2803_26[0]),.doutb(w_n2803_26[1]),.doutc(w_n2803_26[2]),.din(w_n2803_8[1]));
	jspl3 jspl3_w_n2803_27(.douta(w_n2803_27[0]),.doutb(w_n2803_27[1]),.doutc(w_n2803_27[2]),.din(w_n2803_8[2]));
	jspl3 jspl3_w_n2803_28(.douta(w_n2803_28[0]),.doutb(w_n2803_28[1]),.doutc(w_n2803_28[2]),.din(w_n2803_9[0]));
	jspl3 jspl3_w_n2803_29(.douta(w_n2803_29[0]),.doutb(w_n2803_29[1]),.doutc(w_n2803_29[2]),.din(w_n2803_9[1]));
	jspl3 jspl3_w_n2803_30(.douta(w_n2803_30[0]),.doutb(w_n2803_30[1]),.doutc(w_n2803_30[2]),.din(w_n2803_9[2]));
	jspl3 jspl3_w_n2803_31(.douta(w_n2803_31[0]),.doutb(w_n2803_31[1]),.doutc(w_n2803_31[2]),.din(w_n2803_10[0]));
	jspl3 jspl3_w_n2803_32(.douta(w_n2803_32[0]),.doutb(w_n2803_32[1]),.doutc(w_n2803_32[2]),.din(w_n2803_10[1]));
	jspl3 jspl3_w_n2803_33(.douta(w_n2803_33[0]),.doutb(w_n2803_33[1]),.doutc(w_n2803_33[2]),.din(w_n2803_10[2]));
	jspl3 jspl3_w_n2803_34(.douta(w_n2803_34[0]),.doutb(w_n2803_34[1]),.doutc(w_n2803_34[2]),.din(w_n2803_11[0]));
	jspl3 jspl3_w_n2803_35(.douta(w_n2803_35[0]),.doutb(w_n2803_35[1]),.doutc(w_n2803_35[2]),.din(w_n2803_11[1]));
	jspl3 jspl3_w_n2803_36(.douta(w_n2803_36[0]),.doutb(w_n2803_36[1]),.doutc(w_n2803_36[2]),.din(w_n2803_11[2]));
	jspl3 jspl3_w_n2803_37(.douta(w_n2803_37[0]),.doutb(w_n2803_37[1]),.doutc(w_n2803_37[2]),.din(w_n2803_12[0]));
	jspl3 jspl3_w_n2803_38(.douta(w_n2803_38[0]),.doutb(w_n2803_38[1]),.doutc(w_n2803_38[2]),.din(w_n2803_12[1]));
	jspl3 jspl3_w_n2803_39(.douta(w_n2803_39[0]),.doutb(w_n2803_39[1]),.doutc(w_n2803_39[2]),.din(w_n2803_12[2]));
	jspl3 jspl3_w_n2803_40(.douta(w_n2803_40[0]),.doutb(w_n2803_40[1]),.doutc(w_n2803_40[2]),.din(w_n2803_13[0]));
	jspl3 jspl3_w_n2803_41(.douta(w_n2803_41[0]),.doutb(w_n2803_41[1]),.doutc(w_n2803_41[2]),.din(w_n2803_13[1]));
	jspl3 jspl3_w_n2803_42(.douta(w_n2803_42[0]),.doutb(w_n2803_42[1]),.doutc(w_n2803_42[2]),.din(w_n2803_13[2]));
	jspl3 jspl3_w_n2803_43(.douta(w_n2803_43[0]),.doutb(w_n2803_43[1]),.doutc(w_n2803_43[2]),.din(w_n2803_14[0]));
	jspl3 jspl3_w_n2803_44(.douta(w_n2803_44[0]),.doutb(w_n2803_44[1]),.doutc(w_n2803_44[2]),.din(w_n2803_14[1]));
	jspl3 jspl3_w_n2803_45(.douta(w_n2803_45[0]),.doutb(w_n2803_45[1]),.doutc(w_n2803_45[2]),.din(w_n2803_14[2]));
	jspl3 jspl3_w_n2803_46(.douta(w_n2803_46[0]),.doutb(w_n2803_46[1]),.doutc(w_n2803_46[2]),.din(w_n2803_15[0]));
	jspl3 jspl3_w_n2803_47(.douta(w_n2803_47[0]),.doutb(w_n2803_47[1]),.doutc(w_n2803_47[2]),.din(w_n2803_15[1]));
	jspl3 jspl3_w_n2803_48(.douta(w_n2803_48[0]),.doutb(w_n2803_48[1]),.doutc(w_n2803_48[2]),.din(w_n2803_15[2]));
	jspl3 jspl3_w_n2803_49(.douta(w_n2803_49[0]),.doutb(w_n2803_49[1]),.doutc(w_n2803_49[2]),.din(w_n2803_16[0]));
	jspl3 jspl3_w_n2803_50(.douta(w_n2803_50[0]),.doutb(w_n2803_50[1]),.doutc(w_n2803_50[2]),.din(w_n2803_16[1]));
	jspl3 jspl3_w_n2803_51(.douta(w_n2803_51[0]),.doutb(w_n2803_51[1]),.doutc(w_n2803_51[2]),.din(w_n2803_16[2]));
	jspl3 jspl3_w_n2803_52(.douta(w_n2803_52[0]),.doutb(w_n2803_52[1]),.doutc(w_n2803_52[2]),.din(w_n2803_17[0]));
	jspl3 jspl3_w_n2803_53(.douta(w_n2803_53[0]),.doutb(w_n2803_53[1]),.doutc(w_n2803_53[2]),.din(w_n2803_17[1]));
	jspl3 jspl3_w_n2803_54(.douta(w_n2803_54[0]),.doutb(w_n2803_54[1]),.doutc(w_n2803_54[2]),.din(w_n2803_17[2]));
	jspl3 jspl3_w_n2803_55(.douta(w_n2803_55[0]),.doutb(w_n2803_55[1]),.doutc(w_n2803_55[2]),.din(w_n2803_18[0]));
	jspl3 jspl3_w_n2803_56(.douta(w_n2803_56[0]),.doutb(w_n2803_56[1]),.doutc(w_n2803_56[2]),.din(w_n2803_18[1]));
	jspl3 jspl3_w_n2803_57(.douta(w_n2803_57[0]),.doutb(w_n2803_57[1]),.doutc(w_n2803_57[2]),.din(w_n2803_18[2]));
	jspl3 jspl3_w_n2803_58(.douta(w_n2803_58[0]),.doutb(w_n2803_58[1]),.doutc(w_n2803_58[2]),.din(w_n2803_19[0]));
	jspl3 jspl3_w_n2803_59(.douta(w_n2803_59[0]),.doutb(w_n2803_59[1]),.doutc(w_n2803_59[2]),.din(w_n2803_19[1]));
	jspl3 jspl3_w_n2803_60(.douta(w_n2803_60[0]),.doutb(w_n2803_60[1]),.doutc(w_n2803_60[2]),.din(w_n2803_19[2]));
	jspl3 jspl3_w_n2803_61(.douta(w_n2803_61[0]),.doutb(w_n2803_61[1]),.doutc(w_n2803_61[2]),.din(w_n2803_20[0]));
	jspl3 jspl3_w_n2803_62(.douta(w_n2803_62[0]),.doutb(w_n2803_62[1]),.doutc(w_n2803_62[2]),.din(w_n2803_20[1]));
	jspl3 jspl3_w_n2803_63(.douta(w_n2803_63[0]),.doutb(w_n2803_63[1]),.doutc(w_n2803_63[2]),.din(w_n2803_20[2]));
	jspl jspl_w_n2803_64(.douta(w_n2803_64[0]),.doutb(w_n2803_64[1]),.din(w_n2803_21[0]));
	jspl3 jspl3_w_n2808_0(.douta(w_n2808_0[0]),.doutb(w_n2808_0[1]),.doutc(w_n2808_0[2]),.din(n2808));
	jspl3 jspl3_w_n2808_1(.douta(w_n2808_1[0]),.doutb(w_n2808_1[1]),.doutc(w_n2808_1[2]),.din(w_n2808_0[0]));
	jspl3 jspl3_w_n2808_2(.douta(w_n2808_2[0]),.doutb(w_n2808_2[1]),.doutc(w_n2808_2[2]),.din(w_n2808_0[1]));
	jspl3 jspl3_w_n2808_3(.douta(w_n2808_3[0]),.doutb(w_n2808_3[1]),.doutc(w_n2808_3[2]),.din(w_n2808_0[2]));
	jspl3 jspl3_w_n2808_4(.douta(w_n2808_4[0]),.doutb(w_n2808_4[1]),.doutc(w_n2808_4[2]),.din(w_n2808_1[0]));
	jspl3 jspl3_w_n2808_5(.douta(w_n2808_5[0]),.doutb(w_n2808_5[1]),.doutc(w_n2808_5[2]),.din(w_n2808_1[1]));
	jspl3 jspl3_w_n2808_6(.douta(w_n2808_6[0]),.doutb(w_n2808_6[1]),.doutc(w_n2808_6[2]),.din(w_n2808_1[2]));
	jspl3 jspl3_w_n2808_7(.douta(w_n2808_7[0]),.doutb(w_n2808_7[1]),.doutc(w_n2808_7[2]),.din(w_n2808_2[0]));
	jspl3 jspl3_w_n2808_8(.douta(w_n2808_8[0]),.doutb(w_n2808_8[1]),.doutc(w_n2808_8[2]),.din(w_n2808_2[1]));
	jspl3 jspl3_w_n2808_9(.douta(w_n2808_9[0]),.doutb(w_n2808_9[1]),.doutc(w_n2808_9[2]),.din(w_n2808_2[2]));
	jspl3 jspl3_w_n2808_10(.douta(w_n2808_10[0]),.doutb(w_n2808_10[1]),.doutc(w_n2808_10[2]),.din(w_n2808_3[0]));
	jspl3 jspl3_w_n2808_11(.douta(w_n2808_11[0]),.doutb(w_n2808_11[1]),.doutc(w_n2808_11[2]),.din(w_n2808_3[1]));
	jspl3 jspl3_w_n2808_12(.douta(w_n2808_12[0]),.doutb(w_n2808_12[1]),.doutc(w_n2808_12[2]),.din(w_n2808_3[2]));
	jspl3 jspl3_w_n2808_13(.douta(w_n2808_13[0]),.doutb(w_n2808_13[1]),.doutc(w_n2808_13[2]),.din(w_n2808_4[0]));
	jspl3 jspl3_w_n2808_14(.douta(w_n2808_14[0]),.doutb(w_n2808_14[1]),.doutc(w_n2808_14[2]),.din(w_n2808_4[1]));
	jspl3 jspl3_w_n2808_15(.douta(w_n2808_15[0]),.doutb(w_n2808_15[1]),.doutc(w_n2808_15[2]),.din(w_n2808_4[2]));
	jspl3 jspl3_w_n2808_16(.douta(w_n2808_16[0]),.doutb(w_n2808_16[1]),.doutc(w_n2808_16[2]),.din(w_n2808_5[0]));
	jspl3 jspl3_w_n2808_17(.douta(w_n2808_17[0]),.doutb(w_n2808_17[1]),.doutc(w_n2808_17[2]),.din(w_n2808_5[1]));
	jspl3 jspl3_w_n2808_18(.douta(w_n2808_18[0]),.doutb(w_n2808_18[1]),.doutc(w_n2808_18[2]),.din(w_n2808_5[2]));
	jspl3 jspl3_w_n2808_19(.douta(w_n2808_19[0]),.doutb(w_n2808_19[1]),.doutc(w_n2808_19[2]),.din(w_n2808_6[0]));
	jspl3 jspl3_w_n2808_20(.douta(w_n2808_20[0]),.doutb(w_n2808_20[1]),.doutc(w_n2808_20[2]),.din(w_n2808_6[1]));
	jspl3 jspl3_w_n2808_21(.douta(w_n2808_21[0]),.doutb(w_n2808_21[1]),.doutc(w_n2808_21[2]),.din(w_n2808_6[2]));
	jspl3 jspl3_w_n2808_22(.douta(w_n2808_22[0]),.doutb(w_n2808_22[1]),.doutc(w_n2808_22[2]),.din(w_n2808_7[0]));
	jspl3 jspl3_w_n2808_23(.douta(w_n2808_23[0]),.doutb(w_n2808_23[1]),.doutc(w_n2808_23[2]),.din(w_n2808_7[1]));
	jspl3 jspl3_w_n2808_24(.douta(w_n2808_24[0]),.doutb(w_n2808_24[1]),.doutc(w_n2808_24[2]),.din(w_n2808_7[2]));
	jspl3 jspl3_w_n2808_25(.douta(w_n2808_25[0]),.doutb(w_n2808_25[1]),.doutc(w_n2808_25[2]),.din(w_n2808_8[0]));
	jspl3 jspl3_w_n2808_26(.douta(w_n2808_26[0]),.doutb(w_n2808_26[1]),.doutc(w_n2808_26[2]),.din(w_n2808_8[1]));
	jspl3 jspl3_w_n2808_27(.douta(w_n2808_27[0]),.doutb(w_n2808_27[1]),.doutc(w_n2808_27[2]),.din(w_n2808_8[2]));
	jspl3 jspl3_w_n2808_28(.douta(w_n2808_28[0]),.doutb(w_n2808_28[1]),.doutc(w_n2808_28[2]),.din(w_n2808_9[0]));
	jspl3 jspl3_w_n2808_29(.douta(w_n2808_29[0]),.doutb(w_n2808_29[1]),.doutc(w_n2808_29[2]),.din(w_n2808_9[1]));
	jspl3 jspl3_w_n2808_30(.douta(w_n2808_30[0]),.doutb(w_n2808_30[1]),.doutc(w_n2808_30[2]),.din(w_n2808_9[2]));
	jspl3 jspl3_w_n2808_31(.douta(w_n2808_31[0]),.doutb(w_n2808_31[1]),.doutc(w_n2808_31[2]),.din(w_n2808_10[0]));
	jspl3 jspl3_w_n2808_32(.douta(w_n2808_32[0]),.doutb(w_n2808_32[1]),.doutc(w_n2808_32[2]),.din(w_n2808_10[1]));
	jspl3 jspl3_w_n2808_33(.douta(w_n2808_33[0]),.doutb(w_n2808_33[1]),.doutc(w_n2808_33[2]),.din(w_n2808_10[2]));
	jspl3 jspl3_w_n2808_34(.douta(w_n2808_34[0]),.doutb(w_n2808_34[1]),.doutc(w_n2808_34[2]),.din(w_n2808_11[0]));
	jspl3 jspl3_w_n2808_35(.douta(w_n2808_35[0]),.doutb(w_n2808_35[1]),.doutc(w_n2808_35[2]),.din(w_n2808_11[1]));
	jspl3 jspl3_w_n2808_36(.douta(w_n2808_36[0]),.doutb(w_n2808_36[1]),.doutc(w_n2808_36[2]),.din(w_n2808_11[2]));
	jspl3 jspl3_w_n2808_37(.douta(w_n2808_37[0]),.doutb(w_n2808_37[1]),.doutc(w_n2808_37[2]),.din(w_n2808_12[0]));
	jspl3 jspl3_w_n2808_38(.douta(w_n2808_38[0]),.doutb(w_n2808_38[1]),.doutc(w_n2808_38[2]),.din(w_n2808_12[1]));
	jspl3 jspl3_w_n2808_39(.douta(w_n2808_39[0]),.doutb(w_n2808_39[1]),.doutc(w_n2808_39[2]),.din(w_n2808_12[2]));
	jspl3 jspl3_w_n2808_40(.douta(w_n2808_40[0]),.doutb(w_n2808_40[1]),.doutc(w_n2808_40[2]),.din(w_n2808_13[0]));
	jspl3 jspl3_w_n2808_41(.douta(w_n2808_41[0]),.doutb(w_n2808_41[1]),.doutc(w_n2808_41[2]),.din(w_n2808_13[1]));
	jspl3 jspl3_w_n2808_42(.douta(w_n2808_42[0]),.doutb(w_n2808_42[1]),.doutc(w_n2808_42[2]),.din(w_n2808_13[2]));
	jspl3 jspl3_w_n2808_43(.douta(w_n2808_43[0]),.doutb(w_n2808_43[1]),.doutc(w_n2808_43[2]),.din(w_n2808_14[0]));
	jspl3 jspl3_w_n2808_44(.douta(w_n2808_44[0]),.doutb(w_n2808_44[1]),.doutc(w_n2808_44[2]),.din(w_n2808_14[1]));
	jspl3 jspl3_w_n2808_45(.douta(w_n2808_45[0]),.doutb(w_n2808_45[1]),.doutc(w_n2808_45[2]),.din(w_n2808_14[2]));
	jspl3 jspl3_w_n2808_46(.douta(w_n2808_46[0]),.doutb(w_n2808_46[1]),.doutc(w_n2808_46[2]),.din(w_n2808_15[0]));
	jspl3 jspl3_w_n2808_47(.douta(w_n2808_47[0]),.doutb(w_n2808_47[1]),.doutc(w_n2808_47[2]),.din(w_n2808_15[1]));
	jspl3 jspl3_w_n2808_48(.douta(w_n2808_48[0]),.doutb(w_n2808_48[1]),.doutc(w_n2808_48[2]),.din(w_n2808_15[2]));
	jspl3 jspl3_w_n2808_49(.douta(w_n2808_49[0]),.doutb(w_n2808_49[1]),.doutc(w_n2808_49[2]),.din(w_n2808_16[0]));
	jspl3 jspl3_w_n2808_50(.douta(w_n2808_50[0]),.doutb(w_n2808_50[1]),.doutc(w_n2808_50[2]),.din(w_n2808_16[1]));
	jspl3 jspl3_w_n2808_51(.douta(w_n2808_51[0]),.doutb(w_n2808_51[1]),.doutc(w_n2808_51[2]),.din(w_n2808_16[2]));
	jspl3 jspl3_w_n2808_52(.douta(w_n2808_52[0]),.doutb(w_n2808_52[1]),.doutc(w_n2808_52[2]),.din(w_n2808_17[0]));
	jspl3 jspl3_w_n2808_53(.douta(w_n2808_53[0]),.doutb(w_n2808_53[1]),.doutc(w_n2808_53[2]),.din(w_n2808_17[1]));
	jspl3 jspl3_w_n2808_54(.douta(w_n2808_54[0]),.doutb(w_n2808_54[1]),.doutc(w_n2808_54[2]),.din(w_n2808_17[2]));
	jspl3 jspl3_w_n2808_55(.douta(w_n2808_55[0]),.doutb(w_n2808_55[1]),.doutc(w_n2808_55[2]),.din(w_n2808_18[0]));
	jspl3 jspl3_w_n2808_56(.douta(w_n2808_56[0]),.doutb(w_n2808_56[1]),.doutc(w_n2808_56[2]),.din(w_n2808_18[1]));
	jspl3 jspl3_w_n2808_57(.douta(w_n2808_57[0]),.doutb(w_n2808_57[1]),.doutc(w_n2808_57[2]),.din(w_n2808_18[2]));
	jspl3 jspl3_w_n2808_58(.douta(w_n2808_58[0]),.doutb(w_n2808_58[1]),.doutc(w_n2808_58[2]),.din(w_n2808_19[0]));
	jspl3 jspl3_w_n2808_59(.douta(w_n2808_59[0]),.doutb(w_n2808_59[1]),.doutc(w_n2808_59[2]),.din(w_n2808_19[1]));
	jspl3 jspl3_w_n2808_60(.douta(w_n2808_60[0]),.doutb(w_n2808_60[1]),.doutc(w_n2808_60[2]),.din(w_n2808_19[2]));
	jspl3 jspl3_w_n2808_61(.douta(w_n2808_61[0]),.doutb(w_n2808_61[1]),.doutc(w_n2808_61[2]),.din(w_n2808_20[0]));
	jspl3 jspl3_w_n2808_62(.douta(w_n2808_62[0]),.doutb(w_n2808_62[1]),.doutc(w_n2808_62[2]),.din(w_n2808_20[1]));
	jspl3 jspl3_w_n2808_63(.douta(w_n2808_63[0]),.doutb(w_n2808_63[1]),.doutc(w_n2808_63[2]),.din(w_n2808_20[2]));
	jspl3 jspl3_w_n2808_64(.douta(w_n2808_64[0]),.doutb(w_n2808_64[1]),.doutc(w_n2808_64[2]),.din(w_n2808_21[0]));
	jspl jspl_w_n2810_0(.douta(w_n2810_0[0]),.doutb(w_n2810_0[1]),.din(n2810));
	jspl jspl_w_n2811_0(.douta(w_n2811_0[0]),.doutb(w_n2811_0[1]),.din(n2811));
	jspl jspl_w_n2815_0(.douta(w_n2815_0[0]),.doutb(w_n2815_0[1]),.din(n2815));
	jspl jspl_w_n2818_0(.douta(w_n2818_0[0]),.doutb(w_n2818_0[1]),.din(n2818));
	jspl jspl_w_n2819_0(.douta(w_n2819_0[0]),.doutb(w_n2819_0[1]),.din(n2819));
	jspl jspl_w_n2821_0(.douta(w_n2821_0[0]),.doutb(w_n2821_0[1]),.din(n2821));
	jspl jspl_w_n2825_0(.douta(w_n2825_0[0]),.doutb(w_n2825_0[1]),.din(n2825));
	jspl jspl_w_n2826_0(.douta(w_n2826_0[0]),.doutb(w_n2826_0[1]),.din(n2826));
	jspl jspl_w_n2829_0(.douta(w_n2829_0[0]),.doutb(w_n2829_0[1]),.din(n2829));
	jspl jspl_w_n2831_0(.douta(w_n2831_0[0]),.doutb(w_n2831_0[1]),.din(n2831));
	jspl jspl_w_n2835_0(.douta(w_n2835_0[0]),.doutb(w_n2835_0[1]),.din(n2835));
	jspl jspl_w_n2837_0(.douta(w_n2837_0[0]),.doutb(w_n2837_0[1]),.din(n2837));
	jspl jspl_w_n2839_0(.douta(w_n2839_0[0]),.doutb(w_n2839_0[1]),.din(n2839));
	jspl jspl_w_n2841_0(.douta(w_n2841_0[0]),.doutb(w_n2841_0[1]),.din(n2841));
	jspl jspl_w_n2844_0(.douta(w_n2844_0[0]),.doutb(w_n2844_0[1]),.din(n2844));
	jspl jspl_w_n2845_0(.douta(w_n2845_0[0]),.doutb(w_n2845_0[1]),.din(n2845));
	jspl jspl_w_n2848_0(.douta(w_n2848_0[0]),.doutb(w_n2848_0[1]),.din(n2848));
	jspl jspl_w_n2852_0(.douta(w_n2852_0[0]),.doutb(w_n2852_0[1]),.din(n2852));
	jspl jspl_w_n2855_0(.douta(w_n2855_0[0]),.doutb(w_n2855_0[1]),.din(n2855));
	jspl jspl_w_n2856_0(.douta(w_n2856_0[0]),.doutb(w_n2856_0[1]),.din(n2856));
	jspl jspl_w_n2857_0(.douta(w_n2857_0[0]),.doutb(w_n2857_0[1]),.din(n2857));
	jspl jspl_w_n2860_0(.douta(w_n2860_0[0]),.doutb(w_n2860_0[1]),.din(n2860));
	jspl jspl_w_n2863_0(.douta(w_n2863_0[0]),.doutb(w_n2863_0[1]),.din(n2863));
	jspl jspl_w_n2864_0(.douta(w_n2864_0[0]),.doutb(w_n2864_0[1]),.din(n2864));
	jspl jspl_w_n2867_0(.douta(w_n2867_0[0]),.doutb(w_n2867_0[1]),.din(n2867));
	jspl jspl_w_n2869_0(.douta(w_n2869_0[0]),.doutb(w_n2869_0[1]),.din(n2869));
	jspl jspl_w_n2873_0(.douta(w_n2873_0[0]),.doutb(w_n2873_0[1]),.din(n2873));
	jspl jspl_w_n2874_0(.douta(w_n2874_0[0]),.doutb(w_n2874_0[1]),.din(n2874));
	jspl jspl_w_n2877_0(.douta(w_n2877_0[0]),.doutb(w_n2877_0[1]),.din(n2877));
	jspl jspl_w_n2882_0(.douta(w_n2882_0[0]),.doutb(w_n2882_0[1]),.din(n2882));
	jspl jspl_w_n2884_0(.douta(w_n2884_0[0]),.doutb(w_n2884_0[1]),.din(n2884));
	jspl jspl_w_n2888_0(.douta(w_n2888_0[0]),.doutb(w_n2888_0[1]),.din(n2888));
	jspl jspl_w_n2892_0(.douta(w_n2892_0[0]),.doutb(w_n2892_0[1]),.din(n2892));
	jspl jspl_w_n2893_0(.douta(w_n2893_0[0]),.doutb(w_n2893_0[1]),.din(n2893));
	jspl jspl_w_n2896_0(.douta(w_n2896_0[0]),.doutb(w_n2896_0[1]),.din(n2896));
	jspl jspl_w_n2897_0(.douta(w_n2897_0[0]),.doutb(w_n2897_0[1]),.din(n2897));
	jspl jspl_w_n2901_0(.douta(w_n2901_0[0]),.doutb(w_n2901_0[1]),.din(n2901));
	jspl jspl_w_n2902_0(.douta(w_n2902_0[0]),.doutb(w_n2902_0[1]),.din(n2902));
	jspl jspl_w_n2905_0(.douta(w_n2905_0[0]),.doutb(w_n2905_0[1]),.din(n2905));
	jspl jspl_w_n2909_0(.douta(w_n2909_0[0]),.doutb(w_n2909_0[1]),.din(n2909));
	jspl jspl_w_n2912_0(.douta(w_n2912_0[0]),.doutb(w_n2912_0[1]),.din(n2912));
	jspl jspl_w_n2913_0(.douta(w_n2913_0[0]),.doutb(w_n2913_0[1]),.din(n2913));
	jspl jspl_w_n2914_0(.douta(w_n2914_0[0]),.doutb(w_n2914_0[1]),.din(n2914));
	jspl jspl_w_n2917_0(.douta(w_n2917_0[0]),.doutb(w_n2917_0[1]),.din(n2917));
	jspl jspl_w_n2920_0(.douta(w_n2920_0[0]),.doutb(w_n2920_0[1]),.din(n2920));
	jspl jspl_w_n2921_0(.douta(w_n2921_0[0]),.doutb(w_n2921_0[1]),.din(n2921));
	jspl jspl_w_n2924_0(.douta(w_n2924_0[0]),.doutb(w_n2924_0[1]),.din(n2924));
	jspl jspl_w_n2926_0(.douta(w_n2926_0[0]),.doutb(w_n2926_0[1]),.din(n2926));
	jspl jspl_w_n2930_0(.douta(w_n2930_0[0]),.doutb(w_n2930_0[1]),.din(n2930));
	jspl jspl_w_n2931_0(.douta(w_n2931_0[0]),.doutb(w_n2931_0[1]),.din(n2931));
	jspl jspl_w_n2934_0(.douta(w_n2934_0[0]),.doutb(w_n2934_0[1]),.din(n2934));
	jspl jspl_w_n2937_0(.douta(w_n2937_0[0]),.doutb(w_n2937_0[1]),.din(n2937));
	jspl jspl_w_n2939_0(.douta(w_n2939_0[0]),.doutb(w_n2939_0[1]),.din(n2939));
	jspl jspl_w_n2941_0(.douta(w_n2941_0[0]),.doutb(w_n2941_0[1]),.din(n2941));
	jspl jspl_w_n2944_0(.douta(w_n2944_0[0]),.doutb(w_n2944_0[1]),.din(n2944));
	jspl jspl_w_n2947_0(.douta(w_n2947_0[0]),.doutb(w_n2947_0[1]),.din(n2947));
	jspl jspl_w_n2948_0(.douta(w_n2948_0[0]),.doutb(w_n2948_0[1]),.din(n2948));
	jspl jspl_w_n2952_0(.douta(w_n2952_0[0]),.doutb(w_n2952_0[1]),.din(n2952));
	jspl jspl_w_n2953_0(.douta(w_n2953_0[0]),.doutb(w_n2953_0[1]),.din(n2953));
	jspl jspl_w_n2956_0(.douta(w_n2956_0[0]),.doutb(w_n2956_0[1]),.din(n2956));
	jspl jspl_w_n2958_0(.douta(w_n2958_0[0]),.doutb(w_n2958_0[1]),.din(n2958));
	jspl jspl_w_n2961_0(.douta(w_n2961_0[0]),.doutb(w_n2961_0[1]),.din(n2961));
	jspl jspl_w_n2964_0(.douta(w_n2964_0[0]),.doutb(w_n2964_0[1]),.din(n2964));
	jspl jspl_w_n2965_0(.douta(w_n2965_0[0]),.doutb(w_n2965_0[1]),.din(n2965));
	jspl jspl_w_n2966_0(.douta(w_n2966_0[0]),.doutb(w_n2966_0[1]),.din(n2966));
	jspl jspl_w_n2969_0(.douta(w_n2969_0[0]),.doutb(w_n2969_0[1]),.din(n2969));
	jspl jspl_w_n2970_0(.douta(w_n2970_0[0]),.doutb(w_n2970_0[1]),.din(n2970));
	jspl jspl_w_n2973_0(.douta(w_n2973_0[0]),.doutb(w_n2973_0[1]),.din(n2973));
	jspl jspl_w_n2976_0(.douta(w_n2976_0[0]),.doutb(w_n2976_0[1]),.din(n2976));
	jspl jspl_w_n2979_0(.douta(w_n2979_0[0]),.doutb(w_n2979_0[1]),.din(n2979));
	jspl jspl_w_n2982_0(.douta(w_n2982_0[0]),.doutb(w_n2982_0[1]),.din(n2982));
	jspl jspl_w_n2983_0(.douta(w_n2983_0[0]),.doutb(w_n2983_0[1]),.din(n2983));
	jspl jspl_w_n2987_0(.douta(w_n2987_0[0]),.doutb(w_n2987_0[1]),.din(n2987));
	jspl jspl_w_n2988_0(.douta(w_n2988_0[0]),.doutb(w_n2988_0[1]),.din(n2988));
	jspl jspl_w_n2991_0(.douta(w_n2991_0[0]),.doutb(w_n2991_0[1]),.din(n2991));
	jspl jspl_w_n2995_0(.douta(w_n2995_0[0]),.doutb(w_n2995_0[1]),.din(n2995));
	jspl jspl_w_n2998_0(.douta(w_n2998_0[0]),.doutb(w_n2998_0[1]),.din(n2998));
	jspl jspl_w_n2999_0(.douta(w_n2999_0[0]),.doutb(w_n2999_0[1]),.din(n2999));
	jspl jspl_w_n3000_0(.douta(w_n3000_0[0]),.doutb(w_n3000_0[1]),.din(n3000));
	jspl jspl_w_n3003_0(.douta(w_n3003_0[0]),.doutb(w_n3003_0[1]),.din(n3003));
	jspl jspl_w_n3006_0(.douta(w_n3006_0[0]),.doutb(w_n3006_0[1]),.din(n3006));
	jspl jspl_w_n3007_0(.douta(w_n3007_0[0]),.doutb(w_n3007_0[1]),.din(n3007));
	jspl jspl_w_n3010_0(.douta(w_n3010_0[0]),.doutb(w_n3010_0[1]),.din(n3010));
	jspl jspl_w_n3011_0(.douta(w_n3011_0[0]),.doutb(w_n3011_0[1]),.din(n3011));
	jspl jspl_w_n3014_0(.douta(w_n3014_0[0]),.doutb(w_n3014_0[1]),.din(n3014));
	jspl jspl_w_n3017_0(.douta(w_n3017_0[0]),.doutb(w_n3017_0[1]),.din(n3017));
	jspl jspl_w_n3018_0(.douta(w_n3018_0[0]),.doutb(w_n3018_0[1]),.din(n3018));
	jspl jspl_w_n3022_0(.douta(w_n3022_0[0]),.doutb(w_n3022_0[1]),.din(n3022));
	jspl jspl_w_n3023_0(.douta(w_n3023_0[0]),.doutb(w_n3023_0[1]),.din(n3023));
	jspl jspl_w_n3026_0(.douta(w_n3026_0[0]),.doutb(w_n3026_0[1]),.din(n3026));
	jspl jspl_w_n3028_0(.douta(w_n3028_0[0]),.doutb(w_n3028_0[1]),.din(n3028));
	jspl jspl_w_n3031_0(.douta(w_n3031_0[0]),.doutb(w_n3031_0[1]),.din(n3031));
	jspl jspl_w_n3034_0(.douta(w_n3034_0[0]),.doutb(w_n3034_0[1]),.din(n3034));
	jspl jspl_w_n3035_0(.douta(w_n3035_0[0]),.doutb(w_n3035_0[1]),.din(n3035));
	jspl jspl_w_n3036_0(.douta(w_n3036_0[0]),.doutb(w_n3036_0[1]),.din(n3036));
	jspl jspl_w_n3039_0(.douta(w_n3039_0[0]),.doutb(w_n3039_0[1]),.din(n3039));
	jspl jspl_w_n3040_0(.douta(w_n3040_0[0]),.doutb(w_n3040_0[1]),.din(n3040));
	jspl jspl_w_n3043_0(.douta(w_n3043_0[0]),.doutb(w_n3043_0[1]),.din(n3043));
	jspl jspl_w_n3046_0(.douta(w_n3046_0[0]),.doutb(w_n3046_0[1]),.din(n3046));
	jspl jspl_w_n3049_0(.douta(w_n3049_0[0]),.doutb(w_n3049_0[1]),.din(n3049));
	jspl jspl_w_n3052_0(.douta(w_n3052_0[0]),.doutb(w_n3052_0[1]),.din(n3052));
	jspl jspl_w_n3053_0(.douta(w_n3053_0[0]),.doutb(w_n3053_0[1]),.din(n3053));
	jspl jspl_w_n3057_0(.douta(w_n3057_0[0]),.doutb(w_n3057_0[1]),.din(n3057));
	jspl jspl_w_n3058_0(.douta(w_n3058_0[0]),.doutb(w_n3058_0[1]),.din(n3058));
	jspl jspl_w_n3061_0(.douta(w_n3061_0[0]),.doutb(w_n3061_0[1]),.din(n3061));
	jspl jspl_w_n3065_0(.douta(w_n3065_0[0]),.doutb(w_n3065_0[1]),.din(n3065));
	jspl jspl_w_n3068_0(.douta(w_n3068_0[0]),.doutb(w_n3068_0[1]),.din(n3068));
	jspl jspl_w_n3069_0(.douta(w_n3069_0[0]),.doutb(w_n3069_0[1]),.din(n3069));
	jspl jspl_w_n3070_0(.douta(w_n3070_0[0]),.doutb(w_n3070_0[1]),.din(n3070));
	jspl jspl_w_n3073_0(.douta(w_n3073_0[0]),.doutb(w_n3073_0[1]),.din(n3073));
	jspl jspl_w_n3076_0(.douta(w_n3076_0[0]),.doutb(w_n3076_0[1]),.din(n3076));
	jspl jspl_w_n3077_0(.douta(w_n3077_0[0]),.doutb(w_n3077_0[1]),.din(n3077));
	jspl jspl_w_n3080_0(.douta(w_n3080_0[0]),.doutb(w_n3080_0[1]),.din(n3080));
	jspl jspl_w_n3081_0(.douta(w_n3081_0[0]),.doutb(w_n3081_0[1]),.din(n3081));
	jspl jspl_w_n3084_0(.douta(w_n3084_0[0]),.doutb(w_n3084_0[1]),.din(n3084));
	jspl jspl_w_n3087_0(.douta(w_n3087_0[0]),.doutb(w_n3087_0[1]),.din(n3087));
	jspl jspl_w_n3088_0(.douta(w_n3088_0[0]),.doutb(w_n3088_0[1]),.din(n3088));
	jspl jspl_w_n3092_0(.douta(w_n3092_0[0]),.doutb(w_n3092_0[1]),.din(n3092));
	jspl jspl_w_n3093_0(.douta(w_n3093_0[0]),.doutb(w_n3093_0[1]),.din(n3093));
	jspl jspl_w_n3096_0(.douta(w_n3096_0[0]),.doutb(w_n3096_0[1]),.din(n3096));
	jspl jspl_w_n3098_0(.douta(w_n3098_0[0]),.doutb(w_n3098_0[1]),.din(n3098));
	jspl jspl_w_n3101_0(.douta(w_n3101_0[0]),.doutb(w_n3101_0[1]),.din(n3101));
	jspl jspl_w_n3104_0(.douta(w_n3104_0[0]),.doutb(w_n3104_0[1]),.din(n3104));
	jspl jspl_w_n3105_0(.douta(w_n3105_0[0]),.doutb(w_n3105_0[1]),.din(n3105));
	jspl jspl_w_n3106_0(.douta(w_n3106_0[0]),.doutb(w_n3106_0[1]),.din(n3106));
	jspl jspl_w_n3109_0(.douta(w_n3109_0[0]),.doutb(w_n3109_0[1]),.din(n3109));
	jspl jspl_w_n3110_0(.douta(w_n3110_0[0]),.doutb(w_n3110_0[1]),.din(n3110));
	jspl jspl_w_n3113_0(.douta(w_n3113_0[0]),.doutb(w_n3113_0[1]),.din(n3113));
	jspl jspl_w_n3116_0(.douta(w_n3116_0[0]),.doutb(w_n3116_0[1]),.din(n3116));
	jspl jspl_w_n3119_0(.douta(w_n3119_0[0]),.doutb(w_n3119_0[1]),.din(n3119));
	jspl jspl_w_n3120_0(.douta(w_n3120_0[0]),.doutb(w_n3120_0[1]),.din(n3120));
	jspl jspl_w_n3123_0(.douta(w_n3123_0[0]),.doutb(w_n3123_0[1]),.din(n3123));
	jspl jspl_w_n3127_0(.douta(w_n3127_0[0]),.doutb(w_n3127_0[1]),.din(n3127));
	jspl jspl_w_n3130_0(.douta(w_n3130_0[0]),.doutb(w_n3130_0[1]),.din(n3130));
	jspl jspl_w_n3131_0(.douta(w_n3131_0[0]),.doutb(w_n3131_0[1]),.din(n3131));
	jspl jspl_w_n3132_0(.douta(w_n3132_0[0]),.doutb(w_n3132_0[1]),.din(n3132));
	jspl jspl_w_n3135_0(.douta(w_n3135_0[0]),.doutb(w_n3135_0[1]),.din(n3135));
	jspl jspl_w_n3138_0(.douta(w_n3138_0[0]),.doutb(w_n3138_0[1]),.din(n3138));
	jspl jspl_w_n3139_0(.douta(w_n3139_0[0]),.doutb(w_n3139_0[1]),.din(n3139));
	jspl jspl_w_n3142_0(.douta(w_n3142_0[0]),.doutb(w_n3142_0[1]),.din(n3142));
	jspl jspl_w_n3144_0(.douta(w_n3144_0[0]),.doutb(w_n3144_0[1]),.din(n3144));
	jspl jspl_w_n3148_0(.douta(w_n3148_0[0]),.doutb(w_n3148_0[1]),.din(n3148));
	jspl jspl_w_n3149_0(.douta(w_n3149_0[0]),.doutb(w_n3149_0[1]),.din(n3149));
	jspl jspl_w_n3152_0(.douta(w_n3152_0[0]),.doutb(w_n3152_0[1]),.din(n3152));
	jspl jspl_w_n3155_0(.douta(w_n3155_0[0]),.doutb(w_n3155_0[1]),.din(n3155));
	jspl jspl_w_n3158_0(.douta(w_n3158_0[0]),.doutb(w_n3158_0[1]),.din(n3158));
	jspl jspl_w_n3160_0(.douta(w_n3160_0[0]),.doutb(w_n3160_0[1]),.din(n3160));
	jspl jspl_w_n3163_0(.douta(w_n3163_0[0]),.doutb(w_n3163_0[1]),.din(n3163));
	jspl jspl_w_n3167_0(.douta(w_n3167_0[0]),.doutb(w_n3167_0[1]),.din(n3167));
	jspl jspl_w_n3168_0(.douta(w_n3168_0[0]),.doutb(w_n3168_0[1]),.din(n3168));
	jspl jspl_w_n3171_0(.douta(w_n3171_0[0]),.doutb(w_n3171_0[1]),.din(n3171));
	jspl jspl_w_n3172_0(.douta(w_n3172_0[0]),.doutb(w_n3172_0[1]),.din(n3172));
	jspl jspl_w_n3174_0(.douta(w_n3174_0[0]),.doutb(w_n3174_0[1]),.din(n3174));
	jspl jspl_w_n3178_0(.douta(w_n3178_0[0]),.doutb(w_n3178_0[1]),.din(n3178));
	jspl jspl_w_n3179_0(.douta(w_n3179_0[0]),.doutb(w_n3179_0[1]),.din(n3179));
	jspl jspl_w_n3182_0(.douta(w_n3182_0[0]),.doutb(w_n3182_0[1]),.din(n3182));
	jspl jspl_w_n3184_0(.douta(w_n3184_0[0]),.doutb(w_n3184_0[1]),.din(n3184));
	jspl jspl_w_n3187_0(.douta(w_n3187_0[0]),.doutb(w_n3187_0[1]),.din(n3187));
	jspl jspl_w_n3190_0(.douta(w_n3190_0[0]),.doutb(w_n3190_0[1]),.din(n3190));
	jspl jspl_w_n3191_0(.douta(w_n3191_0[0]),.doutb(w_n3191_0[1]),.din(n3191));
	jspl jspl_w_n3192_0(.douta(w_n3192_0[0]),.doutb(w_n3192_0[1]),.din(n3192));
	jspl jspl_w_n3195_0(.douta(w_n3195_0[0]),.doutb(w_n3195_0[1]),.din(n3195));
	jspl jspl_w_n3196_0(.douta(w_n3196_0[0]),.doutb(w_n3196_0[1]),.din(n3196));
	jspl jspl_w_n3199_0(.douta(w_n3199_0[0]),.doutb(w_n3199_0[1]),.din(n3199));
	jspl jspl_w_n3202_0(.douta(w_n3202_0[0]),.doutb(w_n3202_0[1]),.din(n3202));
	jspl jspl_w_n3205_0(.douta(w_n3205_0[0]),.doutb(w_n3205_0[1]),.din(n3205));
	jspl jspl_w_n3208_0(.douta(w_n3208_0[0]),.doutb(w_n3208_0[1]),.din(n3208));
	jspl jspl_w_n3209_0(.douta(w_n3209_0[0]),.doutb(w_n3209_0[1]),.din(n3209));
	jspl jspl_w_n3213_0(.douta(w_n3213_0[0]),.doutb(w_n3213_0[1]),.din(n3213));
	jspl jspl_w_n3214_0(.douta(w_n3214_0[0]),.doutb(w_n3214_0[1]),.din(n3214));
	jspl jspl_w_n3217_0(.douta(w_n3217_0[0]),.doutb(w_n3217_0[1]),.din(n3217));
	jspl jspl_w_n3221_0(.douta(w_n3221_0[0]),.doutb(w_n3221_0[1]),.din(n3221));
	jspl jspl_w_n3224_0(.douta(w_n3224_0[0]),.doutb(w_n3224_0[1]),.din(n3224));
	jspl jspl_w_n3225_0(.douta(w_n3225_0[0]),.doutb(w_n3225_0[1]),.din(n3225));
	jspl jspl_w_n3226_0(.douta(w_n3226_0[0]),.doutb(w_n3226_0[1]),.din(n3226));
	jspl jspl_w_n3229_0(.douta(w_n3229_0[0]),.doutb(w_n3229_0[1]),.din(n3229));
	jspl jspl_w_n3232_0(.douta(w_n3232_0[0]),.doutb(w_n3232_0[1]),.din(n3232));
	jspl jspl_w_n3233_0(.douta(w_n3233_0[0]),.doutb(w_n3233_0[1]),.din(n3233));
	jspl jspl_w_n3236_0(.douta(w_n3236_0[0]),.doutb(w_n3236_0[1]),.din(n3236));
	jspl jspl_w_n3237_0(.douta(w_n3237_0[0]),.doutb(w_n3237_0[1]),.din(n3237));
	jspl jspl_w_n3240_0(.douta(w_n3240_0[0]),.doutb(w_n3240_0[1]),.din(n3240));
	jspl jspl_w_n3241_0(.douta(w_n3241_0[0]),.doutb(w_n3241_0[1]),.din(n3241));
	jspl jspl_w_n3244_0(.douta(w_n3244_0[0]),.doutb(w_n3244_0[1]),.din(n3244));
	jspl jspl_w_n3248_0(.douta(w_n3248_0[0]),.doutb(w_n3248_0[1]),.din(n3248));
	jspl jspl_w_n3251_0(.douta(w_n3251_0[0]),.doutb(w_n3251_0[1]),.din(n3251));
	jspl jspl_w_n3252_0(.douta(w_n3252_0[0]),.doutb(w_n3252_0[1]),.din(n3252));
	jspl jspl_w_n3253_0(.douta(w_n3253_0[0]),.doutb(w_n3253_0[1]),.din(n3253));
	jspl jspl_w_n3256_0(.douta(w_n3256_0[0]),.doutb(w_n3256_0[1]),.din(n3256));
	jspl jspl_w_n3259_0(.douta(w_n3259_0[0]),.doutb(w_n3259_0[1]),.din(n3259));
	jspl jspl_w_n3260_0(.douta(w_n3260_0[0]),.doutb(w_n3260_0[1]),.din(n3260));
	jspl jspl_w_n3263_0(.douta(w_n3263_0[0]),.doutb(w_n3263_0[1]),.din(n3263));
	jspl jspl_w_n3265_0(.douta(w_n3265_0[0]),.doutb(w_n3265_0[1]),.din(n3265));
	jspl jspl_w_n3269_0(.douta(w_n3269_0[0]),.doutb(w_n3269_0[1]),.din(n3269));
	jspl jspl_w_n3270_0(.douta(w_n3270_0[0]),.doutb(w_n3270_0[1]),.din(n3270));
	jspl jspl_w_n3273_0(.douta(w_n3273_0[0]),.doutb(w_n3273_0[1]),.din(n3273));
	jspl jspl_w_n3278_0(.douta(w_n3278_0[0]),.doutb(w_n3278_0[1]),.din(n3278));
	jspl jspl_w_n3280_0(.douta(w_n3280_0[0]),.doutb(w_n3280_0[1]),.din(n3280));
	jspl jspl_w_n3284_0(.douta(w_n3284_0[0]),.doutb(w_n3284_0[1]),.din(n3284));
	jspl jspl_w_n3288_0(.douta(w_n3288_0[0]),.doutb(w_n3288_0[1]),.din(n3288));
	jspl jspl_w_n3289_0(.douta(w_n3289_0[0]),.doutb(w_n3289_0[1]),.din(n3289));
	jspl jspl_w_n3292_0(.douta(w_n3292_0[0]),.doutb(w_n3292_0[1]),.din(n3292));
	jspl jspl_w_n3293_0(.douta(w_n3293_0[0]),.doutb(w_n3293_0[1]),.din(n3293));
	jspl jspl_w_n3297_0(.douta(w_n3297_0[0]),.doutb(w_n3297_0[1]),.din(n3297));
	jspl jspl_w_n3300_0(.douta(w_n3300_0[0]),.doutb(w_n3300_0[1]),.din(n3300));
	jspl jspl_w_n3301_0(.douta(w_n3301_0[0]),.doutb(w_n3301_0[1]),.din(n3301));
	jspl jspl_w_n3305_0(.douta(w_n3305_0[0]),.doutb(w_n3305_0[1]),.din(n3305));
	jspl jspl_w_n3306_0(.douta(w_n3306_0[0]),.doutb(w_n3306_0[1]),.din(n3306));
	jspl jspl_w_n3309_0(.douta(w_n3309_0[0]),.doutb(w_n3309_0[1]),.din(n3309));
	jspl jspl_w_n3311_0(.douta(w_n3311_0[0]),.doutb(w_n3311_0[1]),.din(n3311));
	jspl jspl_w_n3312_0(.douta(w_n3312_0[0]),.doutb(w_n3312_0[1]),.din(n3312));
	jspl jspl_w_n3316_0(.douta(w_n3316_0[0]),.doutb(w_n3316_0[1]),.din(n3316));
	jspl jspl_w_n3319_0(.douta(w_n3319_0[0]),.doutb(w_n3319_0[1]),.din(n3319));
	jspl jspl_w_n3320_0(.douta(w_n3320_0[0]),.doutb(w_n3320_0[1]),.din(n3320));
	jspl jspl_w_n3324_0(.douta(w_n3324_0[0]),.doutb(w_n3324_0[1]),.din(n3324));
	jspl jspl_w_n3328_0(.douta(w_n3328_0[0]),.doutb(w_n3328_0[1]),.din(n3328));
	jspl jspl_w_n3331_0(.douta(w_n3331_0[0]),.doutb(w_n3331_0[1]),.din(n3331));
	jspl jspl_w_n3332_0(.douta(w_n3332_0[0]),.doutb(w_n3332_0[1]),.din(n3332));
	jspl jspl_w_n3336_0(.douta(w_n3336_0[0]),.doutb(w_n3336_0[1]),.din(n3336));
	jspl jspl_w_n3337_0(.douta(w_n3337_0[0]),.doutb(w_n3337_0[1]),.din(n3337));
	jspl jspl_w_n3340_0(.douta(w_n3340_0[0]),.doutb(w_n3340_0[1]),.din(n3340));
	jspl jspl_w_n3344_0(.douta(w_n3344_0[0]),.doutb(w_n3344_0[1]),.din(n3344));
	jspl jspl_w_n3347_0(.douta(w_n3347_0[0]),.doutb(w_n3347_0[1]),.din(n3347));
	jspl jspl_w_n3348_0(.douta(w_n3348_0[0]),.doutb(w_n3348_0[1]),.din(n3348));
	jspl jspl_w_n3349_0(.douta(w_n3349_0[0]),.doutb(w_n3349_0[1]),.din(n3349));
	jspl jspl_w_n3352_0(.douta(w_n3352_0[0]),.doutb(w_n3352_0[1]),.din(n3352));
	jspl jspl_w_n3355_0(.douta(w_n3355_0[0]),.doutb(w_n3355_0[1]),.din(n3355));
	jspl jspl_w_n3356_0(.douta(w_n3356_0[0]),.doutb(w_n3356_0[1]),.din(n3356));
	jspl jspl_w_n3359_0(.douta(w_n3359_0[0]),.doutb(w_n3359_0[1]),.din(n3359));
	jspl jspl_w_n3360_0(.douta(w_n3360_0[0]),.doutb(w_n3360_0[1]),.din(n3360));
	jspl jspl_w_n3364_0(.douta(w_n3364_0[0]),.doutb(w_n3364_0[1]),.din(n3364));
	jspl jspl_w_n3365_0(.douta(w_n3365_0[0]),.doutb(w_n3365_0[1]),.din(n3365));
	jspl jspl_w_n3368_0(.douta(w_n3368_0[0]),.doutb(w_n3368_0[1]),.din(n3368));
	jspl jspl_w_n3370_0(.douta(w_n3370_0[0]),.doutb(w_n3370_0[1]),.din(n3370));
	jspl jspl_w_n3374_0(.douta(w_n3374_0[0]),.doutb(w_n3374_0[1]),.din(n3374));
	jspl jspl_w_n3377_0(.douta(w_n3377_0[0]),.doutb(w_n3377_0[1]),.din(n3377));
	jspl jspl_w_n3378_0(.douta(w_n3378_0[0]),.doutb(w_n3378_0[1]),.din(n3378));
	jspl jspl_w_n3380_0(.douta(w_n3380_0[0]),.doutb(w_n3380_0[1]),.din(n3380));
	jspl jspl_w_n3382_0(.douta(w_n3382_0[0]),.doutb(w_n3382_0[1]),.din(n3382));
	jspl jspl_w_n3386_0(.douta(w_n3386_0[0]),.doutb(w_n3386_0[1]),.din(n3386));
	jspl jspl_w_n3389_0(.douta(w_n3389_0[0]),.doutb(w_n3389_0[1]),.din(n3389));
	jspl jspl_w_n3390_0(.douta(w_n3390_0[0]),.doutb(w_n3390_0[1]),.din(n3390));
	jspl jspl_w_n3391_0(.douta(w_n3391_0[0]),.doutb(w_n3391_0[1]),.din(n3391));
	jspl jspl_w_n3395_0(.douta(w_n3395_0[0]),.doutb(w_n3395_0[1]),.din(n3395));
	jspl jspl_w_n3396_0(.douta(w_n3396_0[0]),.doutb(w_n3396_0[1]),.din(n3396));
	jspl jspl_w_n3399_0(.douta(w_n3399_0[0]),.doutb(w_n3399_0[1]),.din(n3399));
	jspl jspl_w_n3402_0(.douta(w_n3402_0[0]),.doutb(w_n3402_0[1]),.din(n3402));
	jspl jspl_w_n3408_0(.douta(w_n3408_0[0]),.doutb(w_n3408_0[1]),.din(n3408));
	jspl jspl_w_n3412_0(.douta(w_n3412_0[0]),.doutb(w_n3412_0[1]),.din(n3412));
	jspl jspl_w_n3413_0(.douta(w_n3413_0[0]),.doutb(w_n3413_0[1]),.din(n3413));
	jspl jspl_w_n3416_0(.douta(w_n3416_0[0]),.doutb(w_n3416_0[1]),.din(n3416));
	jspl jspl_w_n3417_0(.douta(w_n3417_0[0]),.doutb(w_n3417_0[1]),.din(n3417));
	jspl3 jspl3_w_n3421_0(.douta(w_n3421_0[0]),.doutb(w_n3421_0[1]),.doutc(w_n3421_0[2]),.din(n3421));
	jspl jspl_w_n3424_0(.douta(w_n3424_0[0]),.doutb(w_n3424_0[1]),.din(n3424));
	jspl jspl_w_n3427_0(.douta(w_n3427_0[0]),.doutb(w_n3427_0[1]),.din(n3427));
	jspl jspl_w_n3428_0(.douta(w_n3428_0[0]),.doutb(w_n3428_0[1]),.din(n3428));
	jspl jspl_w_n3433_0(.douta(w_n3433_0[0]),.doutb(w_n3433_0[1]),.din(n3433));
	jspl jspl_w_n3436_0(.douta(w_n3436_0[0]),.doutb(w_n3436_0[1]),.din(n3436));
	jspl jspl_w_n3437_0(.douta(w_n3437_0[0]),.doutb(w_n3437_0[1]),.din(n3437));
	jspl jspl_w_n3438_0(.douta(w_n3438_0[0]),.doutb(w_n3438_0[1]),.din(n3438));
	jspl jspl_w_n3441_0(.douta(w_n3441_0[0]),.doutb(w_n3441_0[1]),.din(n3441));
	jspl jspl_w_n3442_0(.douta(w_n3442_0[0]),.doutb(w_n3442_0[1]),.din(n3442));
	jspl jspl_w_n3445_0(.douta(w_n3445_0[0]),.doutb(w_n3445_0[1]),.din(n3445));
	jspl jspl_w_n3448_0(.douta(w_n3448_0[0]),.doutb(w_n3448_0[1]),.din(n3448));
	jspl jspl_w_n3451_0(.douta(w_n3451_0[0]),.doutb(w_n3451_0[1]),.din(n3451));
	jspl jspl_w_n3454_0(.douta(w_n3454_0[0]),.doutb(w_n3454_0[1]),.din(n3454));
	jspl jspl_w_n3455_0(.douta(w_n3455_0[0]),.doutb(w_n3455_0[1]),.din(n3455));
	jspl jspl_w_n3457_0(.douta(w_n3457_0[0]),.doutb(w_n3457_0[1]),.din(n3457));
	jspl jspl_w_n3459_0(.douta(w_n3459_0[0]),.doutb(w_n3459_0[1]),.din(n3459));
	jspl3 jspl3_w_n3463_0(.douta(w_n3463_0[0]),.doutb(w_n3463_0[1]),.doutc(w_n3463_0[2]),.din(n3463));
	jspl jspl_w_n3465_0(.douta(w_n3465_0[0]),.doutb(w_n3465_0[1]),.din(n3465));
	jspl jspl_w_n3469_0(.douta(w_n3469_0[0]),.doutb(w_n3469_0[1]),.din(n3469));
	jspl jspl_w_n3472_0(.douta(w_n3472_0[0]),.doutb(w_n3472_0[1]),.din(n3472));
	jspl jspl_w_n3473_0(.douta(w_n3473_0[0]),.doutb(w_n3473_0[1]),.din(n3473));
	jspl jspl_w_n3475_0(.douta(w_n3475_0[0]),.doutb(w_n3475_0[1]),.din(n3475));
	jspl jspl_w_n3478_0(.douta(w_n3478_0[0]),.doutb(w_n3478_0[1]),.din(n3478));
	jspl jspl_w_n3479_0(.douta(w_n3479_0[0]),.doutb(w_n3479_0[1]),.din(n3479));
	jspl jspl_w_n3482_0(.douta(w_n3482_0[0]),.doutb(w_n3482_0[1]),.din(n3482));
	jspl jspl_w_n3486_0(.douta(w_n3486_0[0]),.doutb(w_n3486_0[1]),.din(n3486));
	jspl jspl_w_n3489_0(.douta(w_n3489_0[0]),.doutb(w_n3489_0[1]),.din(n3489));
	jspl jspl_w_n3490_0(.douta(w_n3490_0[0]),.doutb(w_n3490_0[1]),.din(n3490));
	jspl jspl_w_n3493_0(.douta(w_n3493_0[0]),.doutb(w_n3493_0[1]),.din(n3493));
	jspl jspl_w_n3494_0(.douta(w_n3494_0[0]),.doutb(w_n3494_0[1]),.din(n3494));
	jspl jspl_w_n3498_0(.douta(w_n3498_0[0]),.doutb(w_n3498_0[1]),.din(n3498));
	jspl jspl_w_n3499_0(.douta(w_n3499_0[0]),.doutb(w_n3499_0[1]),.din(n3499));
	jspl jspl_w_n3502_0(.douta(w_n3502_0[0]),.doutb(w_n3502_0[1]),.din(n3502));
	jspl jspl_w_n3505_0(.douta(w_n3505_0[0]),.doutb(w_n3505_0[1]),.din(n3505));
	jspl jspl_w_n3507_0(.douta(w_n3507_0[0]),.doutb(w_n3507_0[1]),.din(n3507));
	jspl jspl_w_n3510_0(.douta(w_n3510_0[0]),.doutb(w_n3510_0[1]),.din(n3510));
	jspl jspl_w_n3513_0(.douta(w_n3513_0[0]),.doutb(w_n3513_0[1]),.din(n3513));
	jspl jspl_w_n3514_0(.douta(w_n3514_0[0]),.doutb(w_n3514_0[1]),.din(n3514));
	jspl jspl_w_n3515_0(.douta(w_n3515_0[0]),.doutb(w_n3515_0[1]),.din(n3515));
	jspl jspl_w_n3519_0(.douta(w_n3519_0[0]),.doutb(w_n3519_0[1]),.din(n3519));
	jspl jspl_w_n3522_0(.douta(w_n3522_0[0]),.doutb(w_n3522_0[1]),.din(n3522));
	jspl jspl_w_n3523_0(.douta(w_n3523_0[0]),.doutb(w_n3523_0[1]),.din(n3523));
	jspl jspl_w_n3527_0(.douta(w_n3527_0[0]),.doutb(w_n3527_0[1]),.din(n3527));
	jspl jspl_w_n3528_0(.douta(w_n3528_0[0]),.doutb(w_n3528_0[1]),.din(n3528));
	jspl jspl_w_n3531_0(.douta(w_n3531_0[0]),.doutb(w_n3531_0[1]),.din(n3531));
	jspl jspl_w_n3533_0(.douta(w_n3533_0[0]),.doutb(w_n3533_0[1]),.din(n3533));
	jspl jspl_w_n3534_0(.douta(w_n3534_0[0]),.doutb(w_n3534_0[1]),.din(n3534));
	jspl jspl_w_n3537_0(.douta(w_n3537_0[0]),.doutb(w_n3537_0[1]),.din(n3537));
	jspl jspl_w_n3540_0(.douta(w_n3540_0[0]),.doutb(w_n3540_0[1]),.din(n3540));
	jspl jspl_w_n3541_0(.douta(w_n3541_0[0]),.doutb(w_n3541_0[1]),.din(n3541));
	jspl jspl_w_n3543_0(.douta(w_n3543_0[0]),.doutb(w_n3543_0[1]),.din(n3543));
	jspl jspl_w_n3547_0(.douta(w_n3547_0[0]),.doutb(w_n3547_0[1]),.din(n3547));
	jspl jspl_w_n3549_0(.douta(w_n3549_0[0]),.doutb(w_n3549_0[1]),.din(n3549));
	jspl jspl_w_n3557_0(.douta(w_n3557_0[0]),.doutb(w_n3557_0[1]),.din(n3557));
	jspl jspl_w_n3559_0(.douta(w_n3559_0[0]),.doutb(w_n3559_0[1]),.din(n3559));
	jspl jspl_w_n3563_0(.douta(w_n3563_0[0]),.doutb(w_n3563_0[1]),.din(n3563));
	jspl jspl_w_n3567_0(.douta(w_n3567_0[0]),.doutb(w_n3567_0[1]),.din(n3567));
	jspl jspl_w_n3568_0(.douta(w_n3568_0[0]),.doutb(w_n3568_0[1]),.din(n3568));
	jspl jspl_w_n3571_0(.douta(w_n3571_0[0]),.doutb(w_n3571_0[1]),.din(n3571));
	jspl jspl_w_n3572_0(.douta(w_n3572_0[0]),.doutb(w_n3572_0[1]),.din(n3572));
	jspl jspl_w_n3576_0(.douta(w_n3576_0[0]),.doutb(w_n3576_0[1]),.din(n3576));
	jspl jspl_w_n3579_0(.douta(w_n3579_0[0]),.doutb(w_n3579_0[1]),.din(n3579));
	jspl jspl_w_n3580_0(.douta(w_n3580_0[0]),.doutb(w_n3580_0[1]),.din(n3580));
	jspl jspl_w_n3581_0(.douta(w_n3581_0[0]),.doutb(w_n3581_0[1]),.din(n3581));
	jspl jspl_w_n3584_0(.douta(w_n3584_0[0]),.doutb(w_n3584_0[1]),.din(n3584));
	jspl jspl_w_n3585_0(.douta(w_n3585_0[0]),.doutb(w_n3585_0[1]),.din(n3585));
	jspl jspl_w_n3588_0(.douta(w_n3588_0[0]),.doutb(w_n3588_0[1]),.din(n3588));
	jspl jspl_w_n3589_0(.douta(w_n3589_0[0]),.doutb(w_n3589_0[1]),.din(n3589));
	jspl jspl_w_n3593_0(.douta(w_n3593_0[0]),.doutb(w_n3593_0[1]),.din(n3593));
	jspl jspl_w_n3596_0(.douta(w_n3596_0[0]),.doutb(w_n3596_0[1]),.din(n3596));
	jspl jspl_w_n3597_0(.douta(w_n3597_0[0]),.doutb(w_n3597_0[1]),.din(n3597));
	jspl jspl_w_n3598_0(.douta(w_n3598_0[0]),.doutb(w_n3598_0[1]),.din(n3598));
	jspl jspl_w_n3601_0(.douta(w_n3601_0[0]),.doutb(w_n3601_0[1]),.din(n3601));
	jspl jspl_w_n3604_0(.douta(w_n3604_0[0]),.doutb(w_n3604_0[1]),.din(n3604));
	jspl jspl_w_n3605_0(.douta(w_n3605_0[0]),.doutb(w_n3605_0[1]),.din(n3605));
	jspl jspl_w_n3609_0(.douta(w_n3609_0[0]),.doutb(w_n3609_0[1]),.din(n3609));
	jspl jspl_w_n3612_0(.douta(w_n3612_0[0]),.doutb(w_n3612_0[1]),.din(n3612));
	jspl jspl_w_n3613_0(.douta(w_n3613_0[0]),.doutb(w_n3613_0[1]),.din(n3613));
	jspl jspl_w_n3615_0(.douta(w_n3615_0[0]),.doutb(w_n3615_0[1]),.din(n3615));
	jspl jspl_w_n3619_0(.douta(w_n3619_0[0]),.doutb(w_n3619_0[1]),.din(n3619));
	jspl jspl_w_n3620_0(.douta(w_n3620_0[0]),.doutb(w_n3620_0[1]),.din(n3620));
	jspl jspl_w_n3623_0(.douta(w_n3623_0[0]),.doutb(w_n3623_0[1]),.din(n3623));
	jspl jspl_w_n3624_0(.douta(w_n3624_0[0]),.doutb(w_n3624_0[1]),.din(n3624));
	jspl jspl_w_n3628_0(.douta(w_n3628_0[0]),.doutb(w_n3628_0[1]),.din(n3628));
	jspl jspl_w_n3631_0(.douta(w_n3631_0[0]),.doutb(w_n3631_0[1]),.din(n3631));
	jspl jspl_w_n3632_0(.douta(w_n3632_0[0]),.doutb(w_n3632_0[1]),.din(n3632));
	jspl jspl_w_n3633_0(.douta(w_n3633_0[0]),.doutb(w_n3633_0[1]),.din(n3633));
	jspl jspl_w_n3636_0(.douta(w_n3636_0[0]),.doutb(w_n3636_0[1]),.din(n3636));
	jspl jspl_w_n3639_0(.douta(w_n3639_0[0]),.doutb(w_n3639_0[1]),.din(n3639));
	jspl jspl_w_n3640_0(.douta(w_n3640_0[0]),.doutb(w_n3640_0[1]),.din(n3640));
	jspl jspl_w_n3641_0(.douta(w_n3641_0[0]),.doutb(w_n3641_0[1]),.din(n3641));
	jspl jspl_w_n3642_0(.douta(w_n3642_0[0]),.doutb(w_n3642_0[1]),.din(n3642));
	jspl jspl_w_n3643_0(.douta(w_n3643_0[0]),.doutb(w_n3643_0[1]),.din(n3643));
	jspl jspl_w_n3647_0(.douta(w_n3647_0[0]),.doutb(w_n3647_0[1]),.din(n3647));
	jspl jspl_w_n3650_0(.douta(w_n3650_0[0]),.doutb(w_n3650_0[1]),.din(n3650));
	jspl jspl_w_n3651_0(.douta(w_n3651_0[0]),.doutb(w_n3651_0[1]),.din(n3651));
	jspl jspl_w_n3652_0(.douta(w_n3652_0[0]),.doutb(w_n3652_0[1]),.din(n3652));
	jspl jspl_w_n3655_0(.douta(w_n3655_0[0]),.doutb(w_n3655_0[1]),.din(n3655));
	jspl jspl_w_n3658_0(.douta(w_n3658_0[0]),.doutb(w_n3658_0[1]),.din(n3658));
	jspl jspl_w_n3659_0(.douta(w_n3659_0[0]),.doutb(w_n3659_0[1]),.din(n3659));
	jspl jspl_w_n3660_0(.douta(w_n3660_0[0]),.doutb(w_n3660_0[1]),.din(n3660));
	jspl jspl_w_n3663_0(.douta(w_n3663_0[0]),.doutb(w_n3663_0[1]),.din(n3663));
	jspl jspl_w_n3666_0(.douta(w_n3666_0[0]),.doutb(w_n3666_0[1]),.din(n3666));
	jspl jspl_w_n3667_0(.douta(w_n3667_0[0]),.doutb(w_n3667_0[1]),.din(n3667));
	jspl jspl_w_n3668_0(.douta(w_n3668_0[0]),.doutb(w_n3668_0[1]),.din(n3668));
	jspl jspl_w_n3672_0(.douta(w_n3672_0[0]),.doutb(w_n3672_0[1]),.din(n3672));
	jspl jspl_w_n3675_0(.douta(w_n3675_0[0]),.doutb(w_n3675_0[1]),.din(n3675));
	jspl jspl_w_n3676_0(.douta(w_n3676_0[0]),.doutb(w_n3676_0[1]),.din(n3676));
	jspl jspl_w_n3677_0(.douta(w_n3677_0[0]),.doutb(w_n3677_0[1]),.din(n3677));
	jspl jspl_w_n3680_0(.douta(w_n3680_0[0]),.doutb(w_n3680_0[1]),.din(n3680));
	jspl jspl_w_n3683_0(.douta(w_n3683_0[0]),.doutb(w_n3683_0[1]),.din(n3683));
	jspl jspl_w_n3684_0(.douta(w_n3684_0[0]),.doutb(w_n3684_0[1]),.din(n3684));
	jspl jspl_w_n3685_0(.douta(w_n3685_0[0]),.doutb(w_n3685_0[1]),.din(n3685));
	jspl jspl_w_n3688_0(.douta(w_n3688_0[0]),.doutb(w_n3688_0[1]),.din(n3688));
	jspl jspl_w_n3689_0(.douta(w_n3689_0[0]),.doutb(w_n3689_0[1]),.din(n3689));
	jspl jspl_w_n3692_0(.douta(w_n3692_0[0]),.doutb(w_n3692_0[1]),.din(n3692));
	jspl jspl_w_n3693_0(.douta(w_n3693_0[0]),.doutb(w_n3693_0[1]),.din(n3693));
	jspl jspl_w_n3695_0(.douta(w_n3695_0[0]),.doutb(w_n3695_0[1]),.din(n3695));
	jspl jspl_w_n3696_0(.douta(w_n3696_0[0]),.doutb(w_n3696_0[1]),.din(n3696));
	jspl jspl_w_n3699_0(.douta(w_n3699_0[0]),.doutb(w_n3699_0[1]),.din(n3699));
	jspl jspl_w_n3700_0(.douta(w_n3700_0[0]),.doutb(w_n3700_0[1]),.din(n3700));
	jspl jspl_w_n3703_0(.douta(w_n3703_0[0]),.doutb(w_n3703_0[1]),.din(n3703));
	jspl jspl_w_n3704_0(.douta(w_n3704_0[0]),.doutb(w_n3704_0[1]),.din(n3704));
	jspl jspl_w_n3708_0(.douta(w_n3708_0[0]),.doutb(w_n3708_0[1]),.din(n3708));
	jspl jspl_w_n3711_0(.douta(w_n3711_0[0]),.doutb(w_n3711_0[1]),.din(n3711));
	jspl jspl_w_n3712_0(.douta(w_n3712_0[0]),.doutb(w_n3712_0[1]),.din(n3712));
	jspl jspl_w_n3713_0(.douta(w_n3713_0[0]),.doutb(w_n3713_0[1]),.din(n3713));
	jspl jspl_w_n3716_0(.douta(w_n3716_0[0]),.doutb(w_n3716_0[1]),.din(n3716));
	jspl jspl_w_n3719_0(.douta(w_n3719_0[0]),.doutb(w_n3719_0[1]),.din(n3719));
	jspl jspl_w_n3720_0(.douta(w_n3720_0[0]),.doutb(w_n3720_0[1]),.din(n3720));
	jspl jspl_w_n3721_0(.douta(w_n3721_0[0]),.doutb(w_n3721_0[1]),.din(n3721));
	jspl jspl_w_n3725_0(.douta(w_n3725_0[0]),.doutb(w_n3725_0[1]),.din(n3725));
	jspl jspl_w_n3728_0(.douta(w_n3728_0[0]),.doutb(w_n3728_0[1]),.din(n3728));
	jspl jspl_w_n3729_0(.douta(w_n3729_0[0]),.doutb(w_n3729_0[1]),.din(n3729));
	jspl jspl_w_n3730_0(.douta(w_n3730_0[0]),.doutb(w_n3730_0[1]),.din(n3730));
	jspl jspl_w_n3733_0(.douta(w_n3733_0[0]),.doutb(w_n3733_0[1]),.din(n3733));
	jspl jspl_w_n3734_0(.douta(w_n3734_0[0]),.doutb(w_n3734_0[1]),.din(n3734));
	jspl jspl_w_n3737_0(.douta(w_n3737_0[0]),.doutb(w_n3737_0[1]),.din(n3737));
	jspl jspl_w_n3738_0(.douta(w_n3738_0[0]),.doutb(w_n3738_0[1]),.din(n3738));
	jspl jspl_w_n3741_0(.douta(w_n3741_0[0]),.doutb(w_n3741_0[1]),.din(n3741));
	jspl jspl_w_n3744_0(.douta(w_n3744_0[0]),.doutb(w_n3744_0[1]),.din(n3744));
	jspl jspl_w_n3745_0(.douta(w_n3745_0[0]),.doutb(w_n3745_0[1]),.din(n3745));
	jspl jspl_w_n3746_0(.douta(w_n3746_0[0]),.doutb(w_n3746_0[1]),.din(n3746));
	jspl jspl_w_n3748_0(.douta(w_n3748_0[0]),.doutb(w_n3748_0[1]),.din(n3748));
	jspl jspl_w_n3749_0(.douta(w_n3749_0[0]),.doutb(w_n3749_0[1]),.din(n3749));
	jspl jspl_w_n3752_0(.douta(w_n3752_0[0]),.doutb(w_n3752_0[1]),.din(n3752));
	jspl jspl_w_n3755_0(.douta(w_n3755_0[0]),.doutb(w_n3755_0[1]),.din(n3755));
	jspl jspl_w_n3756_0(.douta(w_n3756_0[0]),.doutb(w_n3756_0[1]),.din(n3756));
	jspl jspl_w_n3757_0(.douta(w_n3757_0[0]),.doutb(w_n3757_0[1]),.din(n3757));
	jspl3 jspl3_w_n3761_0(.douta(w_n3761_0[0]),.doutb(w_n3761_0[1]),.doutc(w_n3761_0[2]),.din(n3761));
	jspl jspl_w_n3764_0(.douta(w_n3764_0[0]),.doutb(w_n3764_0[1]),.din(n3764));
	jspl jspl_w_n3771_0(.douta(w_n3771_0[0]),.doutb(w_n3771_0[1]),.din(n3771));
	jspl jspl_w_n3776_0(.douta(w_n3776_0[0]),.doutb(w_n3776_0[1]),.din(n3776));
	jspl3 jspl3_w_n3779_0(.douta(w_n3779_0[0]),.doutb(w_n3779_0[1]),.doutc(w_n3779_0[2]),.din(n3779));
	jspl jspl_w_n3787_0(.douta(w_n3787_0[0]),.doutb(w_n3787_0[1]),.din(n3787));
	jspl jspl_w_n3790_0(.douta(w_n3790_0[0]),.doutb(w_n3790_0[1]),.din(n3790));
	jspl3 jspl3_w_n3791_0(.douta(w_n3791_0[0]),.doutb(w_n3791_0[1]),.doutc(w_n3791_0[2]),.din(n3791));
	jspl jspl_w_n3795_0(.douta(w_n3795_0[0]),.doutb(w_n3795_0[1]),.din(n3795));
	jspl jspl_w_n3798_0(.douta(w_n3798_0[0]),.doutb(w_n3798_0[1]),.din(n3798));
	jspl jspl_w_n3804_0(.douta(w_n3804_0[0]),.doutb(w_n3804_0[1]),.din(n3804));
	jspl jspl_w_n3806_0(.douta(w_n3806_0[0]),.doutb(w_n3806_0[1]),.din(n3806));
	jspl jspl_w_n3808_0(.douta(w_n3808_0[0]),.doutb(w_n3808_0[1]),.din(n3808));
	jspl jspl_w_n3811_0(.douta(w_n3811_0[0]),.doutb(w_n3811_0[1]),.din(n3811));
	jspl jspl_w_n3812_0(.douta(w_n3812_0[0]),.doutb(w_n3812_0[1]),.din(n3812));
	jspl jspl_w_n3817_0(.douta(w_n3817_0[0]),.doutb(w_n3817_0[1]),.din(n3817));
	jspl jspl_w_n3820_0(.douta(w_n3820_0[0]),.doutb(w_n3820_0[1]),.din(n3820));
	jspl jspl_w_n3821_0(.douta(w_n3821_0[0]),.doutb(w_n3821_0[1]),.din(n3821));
	jspl jspl_w_n3822_0(.douta(w_n3822_0[0]),.doutb(w_n3822_0[1]),.din(n3822));
	jspl jspl_w_n3826_0(.douta(w_n3826_0[0]),.doutb(w_n3826_0[1]),.din(n3826));
	jspl jspl_w_n3827_0(.douta(w_n3827_0[0]),.doutb(w_n3827_0[1]),.din(n3827));
	jspl jspl_w_n3830_0(.douta(w_n3830_0[0]),.doutb(w_n3830_0[1]),.din(n3830));
	jspl jspl_w_n3834_0(.douta(w_n3834_0[0]),.doutb(w_n3834_0[1]),.din(n3834));
	jspl jspl_w_n3835_0(.douta(w_n3835_0[0]),.doutb(w_n3835_0[1]),.din(n3835));
	jspl jspl_w_n3838_0(.douta(w_n3838_0[0]),.doutb(w_n3838_0[1]),.din(n3838));
	jspl jspl_w_n3840_0(.douta(w_n3840_0[0]),.doutb(w_n3840_0[1]),.din(n3840));
	jspl jspl_w_n3843_0(.douta(w_n3843_0[0]),.doutb(w_n3843_0[1]),.din(n3843));
	jspl jspl_w_n3845_0(.douta(w_n3845_0[0]),.doutb(w_n3845_0[1]),.din(n3845));
	jspl jspl_w_n3847_0(.douta(w_n3847_0[0]),.doutb(w_n3847_0[1]),.din(n3847));
	jspl jspl_w_n3853_0(.douta(w_n3853_0[0]),.doutb(w_n3853_0[1]),.din(n3853));
	jspl jspl_w_n3855_0(.douta(w_n3855_0[0]),.doutb(w_n3855_0[1]),.din(n3855));
	jspl jspl_w_n3857_0(.douta(w_n3857_0[0]),.doutb(w_n3857_0[1]),.din(n3857));
	jspl jspl_w_n3860_0(.douta(w_n3860_0[0]),.doutb(w_n3860_0[1]),.din(n3860));
	jspl jspl_w_n3861_0(.douta(w_n3861_0[0]),.doutb(w_n3861_0[1]),.din(n3861));
	jspl jspl_w_n3866_0(.douta(w_n3866_0[0]),.doutb(w_n3866_0[1]),.din(n3866));
	jspl jspl_w_n3869_0(.douta(w_n3869_0[0]),.doutb(w_n3869_0[1]),.din(n3869));
	jspl jspl_w_n3870_0(.douta(w_n3870_0[0]),.doutb(w_n3870_0[1]),.din(n3870));
	jspl jspl_w_n3871_0(.douta(w_n3871_0[0]),.doutb(w_n3871_0[1]),.din(n3871));
	jspl jspl_w_n3875_0(.douta(w_n3875_0[0]),.doutb(w_n3875_0[1]),.din(n3875));
	jspl jspl_w_n3876_0(.douta(w_n3876_0[0]),.doutb(w_n3876_0[1]),.din(n3876));
	jspl jspl_w_n3879_0(.douta(w_n3879_0[0]),.doutb(w_n3879_0[1]),.din(n3879));
	jspl jspl_w_n3881_0(.douta(w_n3881_0[0]),.doutb(w_n3881_0[1]),.din(n3881));
	jspl jspl_w_n3883_0(.douta(w_n3883_0[0]),.doutb(w_n3883_0[1]),.din(n3883));
	jspl jspl_w_n3890_0(.douta(w_n3890_0[0]),.doutb(w_n3890_0[1]),.din(n3890));
	jspl jspl_w_n3893_0(.douta(w_n3893_0[0]),.doutb(w_n3893_0[1]),.din(n3893));
	jspl jspl_w_n3894_0(.douta(w_n3894_0[0]),.doutb(w_n3894_0[1]),.din(n3894));
	jspl jspl_w_n3895_0(.douta(w_n3895_0[0]),.doutb(w_n3895_0[1]),.din(n3895));
	jspl jspl_w_n3898_0(.douta(w_n3898_0[0]),.doutb(w_n3898_0[1]),.din(n3898));
	jspl jspl_w_n3900_0(.douta(w_n3900_0[0]),.doutb(w_n3900_0[1]),.din(n3900));
	jspl jspl_w_n3902_0(.douta(w_n3902_0[0]),.doutb(w_n3902_0[1]),.din(n3902));
	jspl jspl_w_n3907_0(.douta(w_n3907_0[0]),.doutb(w_n3907_0[1]),.din(n3907));
	jspl jspl_w_n3909_0(.douta(w_n3909_0[0]),.doutb(w_n3909_0[1]),.din(n3909));
	jspl jspl_w_n3911_0(.douta(w_n3911_0[0]),.doutb(w_n3911_0[1]),.din(n3911));
	jspl jspl_w_n3914_0(.douta(w_n3914_0[0]),.doutb(w_n3914_0[1]),.din(n3914));
	jspl jspl_w_n3915_0(.douta(w_n3915_0[0]),.doutb(w_n3915_0[1]),.din(n3915));
	jspl jspl_w_n3918_0(.douta(w_n3918_0[0]),.doutb(w_n3918_0[1]),.din(n3918));
	jspl jspl_w_n3922_0(.douta(w_n3922_0[0]),.doutb(w_n3922_0[1]),.din(n3922));
	jspl jspl_w_n3923_0(.douta(w_n3923_0[0]),.doutb(w_n3923_0[1]),.din(n3923));
	jspl jspl_w_n3926_0(.douta(w_n3926_0[0]),.doutb(w_n3926_0[1]),.din(n3926));
	jspl jspl_w_n3928_0(.douta(w_n3928_0[0]),.doutb(w_n3928_0[1]),.din(n3928));
	jspl jspl_w_n3931_0(.douta(w_n3931_0[0]),.doutb(w_n3931_0[1]),.din(n3931));
	jspl jspl_w_n3933_0(.douta(w_n3933_0[0]),.doutb(w_n3933_0[1]),.din(n3933));
	jspl jspl_w_n3935_0(.douta(w_n3935_0[0]),.doutb(w_n3935_0[1]),.din(n3935));
	jspl jspl_w_n3941_0(.douta(w_n3941_0[0]),.doutb(w_n3941_0[1]),.din(n3941));
	jspl jspl_w_n3942_0(.douta(w_n3942_0[0]),.doutb(w_n3942_0[1]),.din(n3942));
	jspl jspl_w_n3945_0(.douta(w_n3945_0[0]),.doutb(w_n3945_0[1]),.din(n3945));
	jspl jspl_w_n3947_0(.douta(w_n3947_0[0]),.doutb(w_n3947_0[1]),.din(n3947));
	jspl jspl_w_n3949_0(.douta(w_n3949_0[0]),.doutb(w_n3949_0[1]),.din(n3949));
	jspl jspl_w_n3952_0(.douta(w_n3952_0[0]),.doutb(w_n3952_0[1]),.din(n3952));
	jspl jspl_w_n3954_0(.douta(w_n3954_0[0]),.doutb(w_n3954_0[1]),.din(n3954));
	jspl jspl_w_n3956_0(.douta(w_n3956_0[0]),.doutb(w_n3956_0[1]),.din(n3956));
	jspl jspl_w_n3960_0(.douta(w_n3960_0[0]),.doutb(w_n3960_0[1]),.din(n3960));
	jspl jspl_w_n3965_0(.douta(w_n3965_0[0]),.doutb(w_n3965_0[1]),.din(n3965));
	jspl jspl_w_n3972_0(.douta(w_n3972_0[0]),.doutb(w_n3972_0[1]),.din(n3972));
	jspl jspl_w_n3975_0(.douta(w_n3975_0[0]),.doutb(w_n3975_0[1]),.din(n3975));
	jspl jspl_w_n3976_0(.douta(w_n3976_0[0]),.doutb(w_n3976_0[1]),.din(n3976));
	jspl jspl_w_n3977_0(.douta(w_n3977_0[0]),.doutb(w_n3977_0[1]),.din(n3977));
	jspl jspl_w_n3980_0(.douta(w_n3980_0[0]),.doutb(w_n3980_0[1]),.din(n3980));
	jspl jspl_w_n3983_0(.douta(w_n3983_0[0]),.doutb(w_n3983_0[1]),.din(n3983));
	jspl jspl_w_n3984_0(.douta(w_n3984_0[0]),.doutb(w_n3984_0[1]),.din(n3984));
	jspl jspl_w_n3988_0(.douta(w_n3988_0[0]),.doutb(w_n3988_0[1]),.din(n3988));
	jspl jspl_w_n3991_0(.douta(w_n3991_0[0]),.doutb(w_n3991_0[1]),.din(n3991));
	jspl jspl_w_n3992_0(.douta(w_n3992_0[0]),.doutb(w_n3992_0[1]),.din(n3992));
	jspl jspl_w_n3997_0(.douta(w_n3997_0[0]),.doutb(w_n3997_0[1]),.din(n3997));
	jspl jspl_w_n4000_0(.douta(w_n4000_0[0]),.doutb(w_n4000_0[1]),.din(n4000));
	jspl jspl_w_n4002_0(.douta(w_n4002_0[0]),.doutb(w_n4002_0[1]),.din(n4002));
	jspl jspl_w_n4005_0(.douta(w_n4005_0[0]),.doutb(w_n4005_0[1]),.din(n4005));
	jspl jspl_w_n4008_0(.douta(w_n4008_0[0]),.doutb(w_n4008_0[1]),.din(n4008));
	jspl jspl_w_n4013_0(.douta(w_n4013_0[0]),.doutb(w_n4013_0[1]),.din(n4013));
	jspl jspl_w_n4015_0(.douta(w_n4015_0[0]),.doutb(w_n4015_0[1]),.din(n4015));
	jspl jspl_w_n4021_0(.douta(w_n4021_0[0]),.doutb(w_n4021_0[1]),.din(n4021));
	jspl jspl_w_n4023_0(.douta(w_n4023_0[0]),.doutb(w_n4023_0[1]),.din(n4023));
	jspl jspl_w_n4028_0(.douta(w_n4028_0[0]),.doutb(w_n4028_0[1]),.din(n4028));
	jspl jspl_w_n4034_0(.douta(w_n4034_0[0]),.doutb(w_n4034_0[1]),.din(n4034));
	jspl jspl_w_n4037_0(.douta(w_n4037_0[0]),.doutb(w_n4037_0[1]),.din(n4037));
	jspl jspl_w_n4038_0(.douta(w_n4038_0[0]),.doutb(w_n4038_0[1]),.din(n4038));
	jspl jspl_w_n4042_0(.douta(w_n4042_0[0]),.doutb(w_n4042_0[1]),.din(n4042));
	jspl jspl_w_n4043_0(.douta(w_n4043_0[0]),.doutb(w_n4043_0[1]),.din(n4043));
	jspl jspl_w_n4046_0(.douta(w_n4046_0[0]),.doutb(w_n4046_0[1]),.din(n4046));
	jspl jspl_w_n4048_0(.douta(w_n4048_0[0]),.doutb(w_n4048_0[1]),.din(n4048));
	jspl jspl_w_n4051_0(.douta(w_n4051_0[0]),.doutb(w_n4051_0[1]),.din(n4051));
	jspl jspl_w_n4052_0(.douta(w_n4052_0[0]),.doutb(w_n4052_0[1]),.din(n4052));
	jspl jspl_w_n4055_0(.douta(w_n4055_0[0]),.doutb(w_n4055_0[1]),.din(n4055));
	jspl jspl_w_n4059_0(.douta(w_n4059_0[0]),.doutb(w_n4059_0[1]),.din(n4059));
	jspl jspl_w_n4062_0(.douta(w_n4062_0[0]),.doutb(w_n4062_0[1]),.din(n4062));
	jspl jspl_w_n4063_0(.douta(w_n4063_0[0]),.doutb(w_n4063_0[1]),.din(n4063));
	jspl jspl_w_n4065_0(.douta(w_n4065_0[0]),.doutb(w_n4065_0[1]),.din(n4065));
	jspl jspl_w_n4066_0(.douta(w_n4066_0[0]),.doutb(w_n4066_0[1]),.din(n4066));
	jspl jspl_w_n4070_0(.douta(w_n4070_0[0]),.doutb(w_n4070_0[1]),.din(n4070));
	jspl jspl_w_n4071_0(.douta(w_n4071_0[0]),.doutb(w_n4071_0[1]),.din(n4071));
	jspl jspl_w_n4074_0(.douta(w_n4074_0[0]),.doutb(w_n4074_0[1]),.din(n4074));
	jspl jspl_w_n4076_0(.douta(w_n4076_0[0]),.doutb(w_n4076_0[1]),.din(n4076));
	jspl jspl_w_n4079_0(.douta(w_n4079_0[0]),.doutb(w_n4079_0[1]),.din(n4079));
	jspl jspl_w_n4080_0(.douta(w_n4080_0[0]),.doutb(w_n4080_0[1]),.din(n4080));
	jspl jspl_w_n4083_0(.douta(w_n4083_0[0]),.doutb(w_n4083_0[1]),.din(n4083));
	jspl jspl_w_n4087_0(.douta(w_n4087_0[0]),.doutb(w_n4087_0[1]),.din(n4087));
	jspl jspl_w_n4090_0(.douta(w_n4090_0[0]),.doutb(w_n4090_0[1]),.din(n4090));
	jspl jspl_w_n4091_0(.douta(w_n4091_0[0]),.doutb(w_n4091_0[1]),.din(n4091));
	jspl jspl_w_n4092_0(.douta(w_n4092_0[0]),.doutb(w_n4092_0[1]),.din(n4092));
	jspl jspl_w_n4096_0(.douta(w_n4096_0[0]),.doutb(w_n4096_0[1]),.din(n4096));
	jspl jspl_w_n4099_0(.douta(w_n4099_0[0]),.doutb(w_n4099_0[1]),.din(n4099));
	jspl jspl_w_n4101_0(.douta(w_n4101_0[0]),.doutb(w_n4101_0[1]),.din(n4101));
	jspl jspl_w_n4104_0(.douta(w_n4104_0[0]),.doutb(w_n4104_0[1]),.din(n4104));
	jspl jspl_w_n4108_0(.douta(w_n4108_0[0]),.doutb(w_n4108_0[1]),.din(n4108));
	jspl jspl_w_n4110_0(.douta(w_n4110_0[0]),.doutb(w_n4110_0[1]),.din(n4110));
	jspl jspl_w_n4114_0(.douta(w_n4114_0[0]),.doutb(w_n4114_0[1]),.din(n4114));
	jspl jspl_w_n4116_0(.douta(w_n4116_0[0]),.doutb(w_n4116_0[1]),.din(n4116));
	jspl jspl_w_n4125_0(.douta(w_n4125_0[0]),.doutb(w_n4125_0[1]),.din(n4125));
	jspl jspl_w_n4129_0(.douta(w_n4129_0[0]),.doutb(w_n4129_0[1]),.din(n4129));
	jspl jspl_w_n4133_0(.douta(w_n4133_0[0]),.doutb(w_n4133_0[1]),.din(n4133));
	jspl jspl_w_n4136_0(.douta(w_n4136_0[0]),.doutb(w_n4136_0[1]),.din(n4136));
	jspl jspl_w_n4138_0(.douta(w_n4138_0[0]),.doutb(w_n4138_0[1]),.din(n4138));
	jspl jspl_w_n4143_0(.douta(w_n4143_0[0]),.doutb(w_n4143_0[1]),.din(n4143));
	jspl jspl_w_n4145_0(.douta(w_n4145_0[0]),.doutb(w_n4145_0[1]),.din(n4145));
	jspl jspl_w_n4149_0(.douta(w_n4149_0[0]),.doutb(w_n4149_0[1]),.din(n4149));
	jspl jspl_w_n4153_0(.douta(w_n4153_0[0]),.doutb(w_n4153_0[1]),.din(n4153));
	jspl jspl_w_n4155_0(.douta(w_n4155_0[0]),.doutb(w_n4155_0[1]),.din(n4155));
	jspl jspl_w_n4158_0(.douta(w_n4158_0[0]),.doutb(w_n4158_0[1]),.din(n4158));
	jspl jspl_w_n4160_0(.douta(w_n4160_0[0]),.doutb(w_n4160_0[1]),.din(n4160));
	jspl jspl_w_n4162_0(.douta(w_n4162_0[0]),.doutb(w_n4162_0[1]),.din(n4162));
	jspl jspl_w_n4165_0(.douta(w_n4165_0[0]),.doutb(w_n4165_0[1]),.din(n4165));
	jspl jspl_w_n4167_0(.douta(w_n4167_0[0]),.doutb(w_n4167_0[1]),.din(n4167));
	jspl jspl_w_n4172_0(.douta(w_n4172_0[0]),.doutb(w_n4172_0[1]),.din(n4172));
	jspl jspl_w_n4173_0(.douta(w_n4173_0[0]),.doutb(w_n4173_0[1]),.din(n4173));
	jspl jspl_w_n4176_0(.douta(w_n4176_0[0]),.doutb(w_n4176_0[1]),.din(n4176));
	jspl jspl_w_n4181_0(.douta(w_n4181_0[0]),.doutb(w_n4181_0[1]),.din(n4181));
	jspl jspl_w_n4184_0(.douta(w_n4184_0[0]),.doutb(w_n4184_0[1]),.din(n4184));
	jspl jspl_w_n4185_0(.douta(w_n4185_0[0]),.doutb(w_n4185_0[1]),.din(n4185));
	jspl jspl_w_n4189_0(.douta(w_n4189_0[0]),.doutb(w_n4189_0[1]),.din(n4189));
	jspl jspl_w_n4190_0(.douta(w_n4190_0[0]),.doutb(w_n4190_0[1]),.din(n4190));
	jspl jspl_w_n4193_0(.douta(w_n4193_0[0]),.doutb(w_n4193_0[1]),.din(n4193));
	jspl jspl_w_n4196_0(.douta(w_n4196_0[0]),.doutb(w_n4196_0[1]),.din(n4196));
	jspl jspl_w_n4199_0(.douta(w_n4199_0[0]),.doutb(w_n4199_0[1]),.din(n4199));
	jspl jspl_w_n4202_0(.douta(w_n4202_0[0]),.doutb(w_n4202_0[1]),.din(n4202));
	jspl jspl_w_n4203_0(.douta(w_n4203_0[0]),.doutb(w_n4203_0[1]),.din(n4203));
	jspl jspl_w_n4205_0(.douta(w_n4205_0[0]),.doutb(w_n4205_0[1]),.din(n4205));
	jspl jspl_w_n4207_0(.douta(w_n4207_0[0]),.doutb(w_n4207_0[1]),.din(n4207));
	jspl jspl_w_n4210_0(.douta(w_n4210_0[0]),.doutb(w_n4210_0[1]),.din(n4210));
	jspl jspl_w_n4212_0(.douta(w_n4212_0[0]),.doutb(w_n4212_0[1]),.din(n4212));
	jspl jspl_w_n4214_0(.douta(w_n4214_0[0]),.doutb(w_n4214_0[1]),.din(n4214));
	jspl jspl_w_n4217_0(.douta(w_n4217_0[0]),.doutb(w_n4217_0[1]),.din(n4217));
	jspl jspl_w_n4222_0(.douta(w_n4222_0[0]),.doutb(w_n4222_0[1]),.din(n4222));
	jspl jspl_w_n4227_0(.douta(w_n4227_0[0]),.doutb(w_n4227_0[1]),.din(n4227));
	jspl jspl_w_n4229_0(.douta(w_n4229_0[0]),.doutb(w_n4229_0[1]),.din(n4229));
	jspl jspl_w_n4234_0(.douta(w_n4234_0[0]),.doutb(w_n4234_0[1]),.din(n4234));
	jspl jspl_w_n4236_0(.douta(w_n4236_0[0]),.doutb(w_n4236_0[1]),.din(n4236));
	jspl jspl_w_n4240_0(.douta(w_n4240_0[0]),.doutb(w_n4240_0[1]),.din(n4240));
	jspl jspl_w_n4245_0(.douta(w_n4245_0[0]),.doutb(w_n4245_0[1]),.din(n4245));
	jspl jspl_w_n4248_0(.douta(w_n4248_0[0]),.doutb(w_n4248_0[1]),.din(n4248));
	jspl jspl_w_n4251_0(.douta(w_n4251_0[0]),.doutb(w_n4251_0[1]),.din(n4251));
	jspl jspl_w_n4255_0(.douta(w_n4255_0[0]),.doutb(w_n4255_0[1]),.din(n4255));
	jspl jspl_w_n4259_0(.douta(w_n4259_0[0]),.doutb(w_n4259_0[1]),.din(n4259));
	jspl jspl_w_n4261_0(.douta(w_n4261_0[0]),.doutb(w_n4261_0[1]),.din(n4261));
	jspl jspl_w_n4266_0(.douta(w_n4266_0[0]),.doutb(w_n4266_0[1]),.din(n4266));
	jspl jspl_w_n4269_0(.douta(w_n4269_0[0]),.doutb(w_n4269_0[1]),.din(n4269));
	jspl jspl_w_n4272_0(.douta(w_n4272_0[0]),.doutb(w_n4272_0[1]),.din(n4272));
	jspl jspl_w_n4275_0(.douta(w_n4275_0[0]),.doutb(w_n4275_0[1]),.din(n4275));
	jspl jspl_w_n4280_0(.douta(w_n4280_0[0]),.doutb(w_n4280_0[1]),.din(n4280));
	jspl jspl_w_n4285_0(.douta(w_n4285_0[0]),.doutb(w_n4285_0[1]),.din(n4285));
	jspl jspl_w_n4287_0(.douta(w_n4287_0[0]),.doutb(w_n4287_0[1]),.din(n4287));
	jspl jspl_w_n4292_0(.douta(w_n4292_0[0]),.doutb(w_n4292_0[1]),.din(n4292));
	jspl jspl_w_n4294_0(.douta(w_n4294_0[0]),.doutb(w_n4294_0[1]),.din(n4294));
	jspl jspl_w_n4298_0(.douta(w_n4298_0[0]),.doutb(w_n4298_0[1]),.din(n4298));
	jspl jspl_w_n4302_0(.douta(w_n4302_0[0]),.doutb(w_n4302_0[1]),.din(n4302));
	jspl jspl_w_n4305_0(.douta(w_n4305_0[0]),.doutb(w_n4305_0[1]),.din(n4305));
	jspl jspl_w_n4308_0(.douta(w_n4308_0[0]),.doutb(w_n4308_0[1]),.din(n4308));
	jspl jspl_w_n4311_0(.douta(w_n4311_0[0]),.doutb(w_n4311_0[1]),.din(n4311));
	jspl jspl_w_n4316_0(.douta(w_n4316_0[0]),.doutb(w_n4316_0[1]),.din(n4316));
	jspl jspl_w_n4321_0(.douta(w_n4321_0[0]),.doutb(w_n4321_0[1]),.din(n4321));
	jspl jspl_w_n4323_0(.douta(w_n4323_0[0]),.doutb(w_n4323_0[1]),.din(n4323));
	jspl jspl_w_n4328_0(.douta(w_n4328_0[0]),.doutb(w_n4328_0[1]),.din(n4328));
	jspl jspl_w_n4330_0(.douta(w_n4330_0[0]),.doutb(w_n4330_0[1]),.din(n4330));
	jspl jspl_w_n4334_0(.douta(w_n4334_0[0]),.doutb(w_n4334_0[1]),.din(n4334));
	jspl jspl_w_n4338_0(.douta(w_n4338_0[0]),.doutb(w_n4338_0[1]),.din(n4338));
	jspl jspl_w_n4341_0(.douta(w_n4341_0[0]),.doutb(w_n4341_0[1]),.din(n4341));
	jspl jspl_w_n4344_0(.douta(w_n4344_0[0]),.doutb(w_n4344_0[1]),.din(n4344));
	jspl jspl_w_n4347_0(.douta(w_n4347_0[0]),.doutb(w_n4347_0[1]),.din(n4347));
	jspl jspl_w_n4352_0(.douta(w_n4352_0[0]),.doutb(w_n4352_0[1]),.din(n4352));
	jspl jspl_w_n4357_0(.douta(w_n4357_0[0]),.doutb(w_n4357_0[1]),.din(n4357));
	jspl jspl_w_n4359_0(.douta(w_n4359_0[0]),.doutb(w_n4359_0[1]),.din(n4359));
	jspl jspl_w_n4362_0(.douta(w_n4362_0[0]),.doutb(w_n4362_0[1]),.din(n4362));
	jspl jspl_w_n4368_0(.douta(w_n4368_0[0]),.doutb(w_n4368_0[1]),.din(n4368));
	jspl jspl_w_n4371_0(.douta(w_n4371_0[0]),.doutb(w_n4371_0[1]),.din(n4371));
	jspl jspl_w_n4372_0(.douta(w_n4372_0[0]),.doutb(w_n4372_0[1]),.din(n4372));
	jspl jspl_w_n4373_0(.douta(w_n4373_0[0]),.doutb(w_n4373_0[1]),.din(n4373));
	jspl jspl_w_n4374_0(.douta(w_n4374_0[0]),.doutb(w_n4374_0[1]),.din(n4374));
	jspl jspl_w_n4378_0(.douta(w_n4378_0[0]),.doutb(w_n4378_0[1]),.din(n4378));
	jspl jspl_w_n4379_0(.douta(w_n4379_0[0]),.doutb(w_n4379_0[1]),.din(n4379));
	jspl jspl_w_n4382_0(.douta(w_n4382_0[0]),.doutb(w_n4382_0[1]),.din(n4382));
	jspl jspl_w_n4384_0(.douta(w_n4384_0[0]),.doutb(w_n4384_0[1]),.din(n4384));
	jspl jspl_w_n4387_0(.douta(w_n4387_0[0]),.doutb(w_n4387_0[1]),.din(n4387));
	jspl jspl_w_n4388_0(.douta(w_n4388_0[0]),.doutb(w_n4388_0[1]),.din(n4388));
	jspl jspl_w_n4391_0(.douta(w_n4391_0[0]),.doutb(w_n4391_0[1]),.din(n4391));
	jspl jspl_w_n4394_0(.douta(w_n4394_0[0]),.doutb(w_n4394_0[1]),.din(n4394));
	jspl jspl_w_n4397_0(.douta(w_n4397_0[0]),.doutb(w_n4397_0[1]),.din(n4397));
	jspl jspl_w_n4400_0(.douta(w_n4400_0[0]),.doutb(w_n4400_0[1]),.din(n4400));
	jspl jspl_w_n4403_0(.douta(w_n4403_0[0]),.doutb(w_n4403_0[1]),.din(n4403));
	jspl jspl_w_n4407_0(.douta(w_n4407_0[0]),.doutb(w_n4407_0[1]),.din(n4407));
	jspl jspl_w_n4411_0(.douta(w_n4411_0[0]),.doutb(w_n4411_0[1]),.din(n4411));
	jspl jspl_w_n4413_0(.douta(w_n4413_0[0]),.doutb(w_n4413_0[1]),.din(n4413));
	jspl jspl_w_n4418_0(.douta(w_n4418_0[0]),.doutb(w_n4418_0[1]),.din(n4418));
	jspl jspl_w_n4419_0(.douta(w_n4419_0[0]),.doutb(w_n4419_0[1]),.din(n4419));
	jspl jspl_w_n4422_0(.douta(w_n4422_0[0]),.doutb(w_n4422_0[1]),.din(n4422));
	jspl jspl_w_n4427_0(.douta(w_n4427_0[0]),.doutb(w_n4427_0[1]),.din(n4427));
	jspl jspl_w_n4430_0(.douta(w_n4430_0[0]),.doutb(w_n4430_0[1]),.din(n4430));
	jspl jspl_w_n4431_0(.douta(w_n4431_0[0]),.doutb(w_n4431_0[1]),.din(n4431));
	jspl jspl_w_n4435_0(.douta(w_n4435_0[0]),.doutb(w_n4435_0[1]),.din(n4435));
	jspl jspl_w_n4436_0(.douta(w_n4436_0[0]),.doutb(w_n4436_0[1]),.din(n4436));
	jspl jspl_w_n4439_0(.douta(w_n4439_0[0]),.doutb(w_n4439_0[1]),.din(n4439));
	jspl jspl_w_n4442_0(.douta(w_n4442_0[0]),.doutb(w_n4442_0[1]),.din(n4442));
	jspl jspl_w_n4445_0(.douta(w_n4445_0[0]),.doutb(w_n4445_0[1]),.din(n4445));
	jspl jspl_w_n4448_0(.douta(w_n4448_0[0]),.doutb(w_n4448_0[1]),.din(n4448));
	jspl jspl_w_n4449_0(.douta(w_n4449_0[0]),.doutb(w_n4449_0[1]),.din(n4449));
	jspl jspl_w_n4451_0(.douta(w_n4451_0[0]),.doutb(w_n4451_0[1]),.din(n4451));
	jspl jspl_w_n4453_0(.douta(w_n4453_0[0]),.doutb(w_n4453_0[1]),.din(n4453));
	jspl jspl_w_n4456_0(.douta(w_n4456_0[0]),.doutb(w_n4456_0[1]),.din(n4456));
	jspl jspl_w_n4458_0(.douta(w_n4458_0[0]),.doutb(w_n4458_0[1]),.din(n4458));
	jspl jspl_w_n4460_0(.douta(w_n4460_0[0]),.doutb(w_n4460_0[1]),.din(n4460));
	jspl jspl_w_n4463_0(.douta(w_n4463_0[0]),.doutb(w_n4463_0[1]),.din(n4463));
	jspl jspl_w_n4468_0(.douta(w_n4468_0[0]),.doutb(w_n4468_0[1]),.din(n4468));
	jspl jspl_w_n4473_0(.douta(w_n4473_0[0]),.doutb(w_n4473_0[1]),.din(n4473));
	jspl jspl_w_n4503_0(.douta(w_n4503_0[0]),.doutb(w_n4503_0[1]),.din(n4503));
	jspl3 jspl3_w_n4506_0(.douta(w_n4506_0[0]),.doutb(w_n4506_0[1]),.doutc(w_n4506_0[2]),.din(n4506));
	jspl3 jspl3_w_n4515_0(.douta(w_n4515_0[0]),.doutb(w_n4515_0[1]),.doutc(w_n4515_0[2]),.din(n4515));
	jspl jspl_w_n4518_0(.douta(w_n4518_0[0]),.doutb(w_n4518_0[1]),.din(n4518));
	jspl jspl_w_n4526_0(.douta(w_n4526_0[0]),.doutb(w_n4526_0[1]),.din(n4526));
	jspl jspl_w_n4644_0(.douta(w_n4644_0[0]),.doutb(w_n4644_0[1]),.din(n4644));
	jspl3 jspl3_w_n4648_0(.douta(w_n4648_0[0]),.doutb(w_n4648_0[1]),.doutc(w_n4648_0[2]),.din(n4648));
	jspl3 jspl3_w_n4648_1(.douta(w_n4648_1[0]),.doutb(w_n4648_1[1]),.doutc(w_n4648_1[2]),.din(w_n4648_0[0]));
	jspl3 jspl3_w_n4648_2(.douta(w_n4648_2[0]),.doutb(w_n4648_2[1]),.doutc(w_n4648_2[2]),.din(w_n4648_0[1]));
	jspl3 jspl3_w_n4648_3(.douta(w_n4648_3[0]),.doutb(w_n4648_3[1]),.doutc(w_n4648_3[2]),.din(w_n4648_0[2]));
	jspl3 jspl3_w_n4648_4(.douta(w_n4648_4[0]),.doutb(w_n4648_4[1]),.doutc(w_n4648_4[2]),.din(w_n4648_1[0]));
	jspl3 jspl3_w_n4648_5(.douta(w_n4648_5[0]),.doutb(w_n4648_5[1]),.doutc(w_n4648_5[2]),.din(w_n4648_1[1]));
	jspl3 jspl3_w_n4648_6(.douta(w_n4648_6[0]),.doutb(w_n4648_6[1]),.doutc(w_n4648_6[2]),.din(w_n4648_1[2]));
	jspl3 jspl3_w_n4648_7(.douta(w_n4648_7[0]),.doutb(w_n4648_7[1]),.doutc(w_n4648_7[2]),.din(w_n4648_2[0]));
	jspl3 jspl3_w_n4648_8(.douta(w_n4648_8[0]),.doutb(w_n4648_8[1]),.doutc(w_n4648_8[2]),.din(w_n4648_2[1]));
	jspl3 jspl3_w_n4648_9(.douta(w_n4648_9[0]),.doutb(w_n4648_9[1]),.doutc(w_n4648_9[2]),.din(w_n4648_2[2]));
	jspl3 jspl3_w_n4648_10(.douta(w_n4648_10[0]),.doutb(w_n4648_10[1]),.doutc(w_n4648_10[2]),.din(w_n4648_3[0]));
	jspl3 jspl3_w_n4648_11(.douta(w_n4648_11[0]),.doutb(w_n4648_11[1]),.doutc(w_n4648_11[2]),.din(w_n4648_3[1]));
	jspl3 jspl3_w_n4648_12(.douta(w_n4648_12[0]),.doutb(w_n4648_12[1]),.doutc(w_n4648_12[2]),.din(w_n4648_3[2]));
	jspl3 jspl3_w_n4648_13(.douta(w_n4648_13[0]),.doutb(w_n4648_13[1]),.doutc(w_n4648_13[2]),.din(w_n4648_4[0]));
	jspl3 jspl3_w_n4648_14(.douta(w_n4648_14[0]),.doutb(w_n4648_14[1]),.doutc(w_n4648_14[2]),.din(w_n4648_4[1]));
	jspl3 jspl3_w_n4648_15(.douta(w_n4648_15[0]),.doutb(w_n4648_15[1]),.doutc(w_n4648_15[2]),.din(w_n4648_4[2]));
	jspl3 jspl3_w_n4648_16(.douta(w_n4648_16[0]),.doutb(w_n4648_16[1]),.doutc(w_n4648_16[2]),.din(w_n4648_5[0]));
	jspl3 jspl3_w_n4648_17(.douta(w_n4648_17[0]),.doutb(w_n4648_17[1]),.doutc(w_n4648_17[2]),.din(w_n4648_5[1]));
	jspl3 jspl3_w_n4648_18(.douta(w_n4648_18[0]),.doutb(w_n4648_18[1]),.doutc(w_n4648_18[2]),.din(w_n4648_5[2]));
	jspl3 jspl3_w_n4648_19(.douta(w_n4648_19[0]),.doutb(w_n4648_19[1]),.doutc(w_n4648_19[2]),.din(w_n4648_6[0]));
	jspl3 jspl3_w_n4648_20(.douta(w_n4648_20[0]),.doutb(w_n4648_20[1]),.doutc(w_n4648_20[2]),.din(w_n4648_6[1]));
	jspl3 jspl3_w_n4648_21(.douta(w_n4648_21[0]),.doutb(w_n4648_21[1]),.doutc(w_n4648_21[2]),.din(w_n4648_6[2]));
	jspl3 jspl3_w_n4648_22(.douta(w_n4648_22[0]),.doutb(w_n4648_22[1]),.doutc(w_n4648_22[2]),.din(w_n4648_7[0]));
	jspl3 jspl3_w_n4648_23(.douta(w_n4648_23[0]),.doutb(w_n4648_23[1]),.doutc(w_n4648_23[2]),.din(w_n4648_7[1]));
	jspl3 jspl3_w_n4648_24(.douta(w_n4648_24[0]),.doutb(w_n4648_24[1]),.doutc(w_n4648_24[2]),.din(w_n4648_7[2]));
	jspl3 jspl3_w_n4648_25(.douta(w_n4648_25[0]),.doutb(w_n4648_25[1]),.doutc(w_n4648_25[2]),.din(w_n4648_8[0]));
	jspl3 jspl3_w_n4648_26(.douta(w_n4648_26[0]),.doutb(w_n4648_26[1]),.doutc(w_n4648_26[2]),.din(w_n4648_8[1]));
	jspl3 jspl3_w_n4648_27(.douta(w_n4648_27[0]),.doutb(w_n4648_27[1]),.doutc(w_n4648_27[2]),.din(w_n4648_8[2]));
	jspl3 jspl3_w_n4648_28(.douta(w_n4648_28[0]),.doutb(w_n4648_28[1]),.doutc(w_n4648_28[2]),.din(w_n4648_9[0]));
	jspl3 jspl3_w_n4648_29(.douta(w_n4648_29[0]),.doutb(w_n4648_29[1]),.doutc(w_n4648_29[2]),.din(w_n4648_9[1]));
	jspl3 jspl3_w_n4648_30(.douta(w_n4648_30[0]),.doutb(w_n4648_30[1]),.doutc(w_n4648_30[2]),.din(w_n4648_9[2]));
	jspl3 jspl3_w_n4648_31(.douta(w_n4648_31[0]),.doutb(w_n4648_31[1]),.doutc(w_n4648_31[2]),.din(w_n4648_10[0]));
	jspl3 jspl3_w_n4648_32(.douta(w_n4648_32[0]),.doutb(w_n4648_32[1]),.doutc(w_n4648_32[2]),.din(w_n4648_10[1]));
	jspl3 jspl3_w_n4648_33(.douta(w_n4648_33[0]),.doutb(w_n4648_33[1]),.doutc(w_n4648_33[2]),.din(w_n4648_10[2]));
	jspl3 jspl3_w_n4648_34(.douta(w_n4648_34[0]),.doutb(w_n4648_34[1]),.doutc(w_n4648_34[2]),.din(w_n4648_11[0]));
	jspl3 jspl3_w_n4648_35(.douta(w_n4648_35[0]),.doutb(w_n4648_35[1]),.doutc(w_n4648_35[2]),.din(w_n4648_11[1]));
	jspl3 jspl3_w_n4648_36(.douta(w_n4648_36[0]),.doutb(w_n4648_36[1]),.doutc(w_n4648_36[2]),.din(w_n4648_11[2]));
	jspl3 jspl3_w_n4648_37(.douta(w_n4648_37[0]),.doutb(w_n4648_37[1]),.doutc(w_n4648_37[2]),.din(w_n4648_12[0]));
	jspl3 jspl3_w_n4648_38(.douta(w_n4648_38[0]),.doutb(w_n4648_38[1]),.doutc(w_n4648_38[2]),.din(w_n4648_12[1]));
	jspl3 jspl3_w_n4648_39(.douta(w_n4648_39[0]),.doutb(w_n4648_39[1]),.doutc(w_n4648_39[2]),.din(w_n4648_12[2]));
	jspl3 jspl3_w_n4648_40(.douta(w_n4648_40[0]),.doutb(w_n4648_40[1]),.doutc(w_n4648_40[2]),.din(w_n4648_13[0]));
	jspl3 jspl3_w_n4648_41(.douta(w_n4648_41[0]),.doutb(w_n4648_41[1]),.doutc(w_n4648_41[2]),.din(w_n4648_13[1]));
	jspl3 jspl3_w_n4648_42(.douta(w_n4648_42[0]),.doutb(w_n4648_42[1]),.doutc(w_n4648_42[2]),.din(w_n4648_13[2]));
	jspl3 jspl3_w_n4648_43(.douta(w_n4648_43[0]),.doutb(w_n4648_43[1]),.doutc(w_n4648_43[2]),.din(w_n4648_14[0]));
	jspl3 jspl3_w_n4648_44(.douta(w_n4648_44[0]),.doutb(w_n4648_44[1]),.doutc(w_n4648_44[2]),.din(w_n4648_14[1]));
	jspl3 jspl3_w_n4648_45(.douta(w_n4648_45[0]),.doutb(w_n4648_45[1]),.doutc(w_n4648_45[2]),.din(w_n4648_14[2]));
	jspl3 jspl3_w_n4648_46(.douta(w_n4648_46[0]),.doutb(w_n4648_46[1]),.doutc(w_n4648_46[2]),.din(w_n4648_15[0]));
	jspl3 jspl3_w_n4648_47(.douta(w_n4648_47[0]),.doutb(w_n4648_47[1]),.doutc(w_n4648_47[2]),.din(w_n4648_15[1]));
	jspl3 jspl3_w_n4648_48(.douta(w_n4648_48[0]),.doutb(w_n4648_48[1]),.doutc(w_n4648_48[2]),.din(w_n4648_15[2]));
	jspl3 jspl3_w_n4648_49(.douta(w_n4648_49[0]),.doutb(w_n4648_49[1]),.doutc(w_n4648_49[2]),.din(w_n4648_16[0]));
	jspl3 jspl3_w_n4648_50(.douta(w_n4648_50[0]),.doutb(w_n4648_50[1]),.doutc(w_n4648_50[2]),.din(w_n4648_16[1]));
	jspl3 jspl3_w_n4648_51(.douta(w_n4648_51[0]),.doutb(w_n4648_51[1]),.doutc(w_n4648_51[2]),.din(w_n4648_16[2]));
	jspl3 jspl3_w_n4648_52(.douta(w_n4648_52[0]),.doutb(w_n4648_52[1]),.doutc(w_n4648_52[2]),.din(w_n4648_17[0]));
	jspl3 jspl3_w_n4648_53(.douta(w_n4648_53[0]),.doutb(w_n4648_53[1]),.doutc(w_n4648_53[2]),.din(w_n4648_17[1]));
	jspl3 jspl3_w_n4648_54(.douta(w_n4648_54[0]),.doutb(w_n4648_54[1]),.doutc(w_n4648_54[2]),.din(w_n4648_17[2]));
	jspl3 jspl3_w_n4648_55(.douta(w_n4648_55[0]),.doutb(w_n4648_55[1]),.doutc(w_n4648_55[2]),.din(w_n4648_18[0]));
	jspl3 jspl3_w_n4648_56(.douta(w_n4648_56[0]),.doutb(w_n4648_56[1]),.doutc(w_n4648_56[2]),.din(w_n4648_18[1]));
	jspl3 jspl3_w_n4648_57(.douta(w_n4648_57[0]),.doutb(w_n4648_57[1]),.doutc(w_n4648_57[2]),.din(w_n4648_18[2]));
	jspl3 jspl3_w_n4648_58(.douta(w_n4648_58[0]),.doutb(w_n4648_58[1]),.doutc(w_n4648_58[2]),.din(w_n4648_19[0]));
	jspl3 jspl3_w_n4648_59(.douta(w_n4648_59[0]),.doutb(w_n4648_59[1]),.doutc(w_n4648_59[2]),.din(w_n4648_19[1]));
	jspl3 jspl3_w_n4648_60(.douta(w_n4648_60[0]),.doutb(w_n4648_60[1]),.doutc(w_n4648_60[2]),.din(w_n4648_19[2]));
	jspl3 jspl3_w_n4648_61(.douta(w_n4648_61[0]),.doutb(w_n4648_61[1]),.doutc(w_n4648_61[2]),.din(w_n4648_20[0]));
	jspl3 jspl3_w_n4648_62(.douta(w_n4648_62[0]),.doutb(w_n4648_62[1]),.doutc(w_n4648_62[2]),.din(w_n4648_20[1]));
	jspl jspl_w_n4648_63(.douta(w_n4648_63[0]),.doutb(w_n4648_63[1]),.din(w_n4648_20[2]));
	jdff dff_A_4jf92R4g9_2(.dout(w_dff_A_WvrfUvCs4_0),.din(w_dff_A_4jf92R4g9_2),.clk(gclk));
	jdff dff_A_WvrfUvCs4_0(.dout(w_dff_A_w2HmUyZ48_0),.din(w_dff_A_WvrfUvCs4_0),.clk(gclk));
	jdff dff_A_w2HmUyZ48_0(.dout(w_dff_A_cEcZOE7F6_0),.din(w_dff_A_w2HmUyZ48_0),.clk(gclk));
	jdff dff_A_cEcZOE7F6_0(.dout(w_dff_A_vRk2r0SD6_0),.din(w_dff_A_cEcZOE7F6_0),.clk(gclk));
	jdff dff_A_vRk2r0SD6_0(.dout(w_dff_A_qewfvzh80_0),.din(w_dff_A_vRk2r0SD6_0),.clk(gclk));
	jdff dff_A_qewfvzh80_0(.dout(w_dff_A_LulQbJwz3_0),.din(w_dff_A_qewfvzh80_0),.clk(gclk));
	jdff dff_A_LulQbJwz3_0(.dout(w_dff_A_cYvKdfOF7_0),.din(w_dff_A_LulQbJwz3_0),.clk(gclk));
	jdff dff_A_cYvKdfOF7_0(.dout(w_dff_A_9kGlvLfv2_0),.din(w_dff_A_cYvKdfOF7_0),.clk(gclk));
	jdff dff_A_9kGlvLfv2_0(.dout(w_dff_A_KiKbdZ2f2_0),.din(w_dff_A_9kGlvLfv2_0),.clk(gclk));
	jdff dff_A_KiKbdZ2f2_0(.dout(w_dff_A_Bb0zsgpd0_0),.din(w_dff_A_KiKbdZ2f2_0),.clk(gclk));
	jdff dff_A_Bb0zsgpd0_0(.dout(w_dff_A_NyxQ7mA05_0),.din(w_dff_A_Bb0zsgpd0_0),.clk(gclk));
	jdff dff_A_NyxQ7mA05_0(.dout(w_dff_A_X6eyEOAP9_0),.din(w_dff_A_NyxQ7mA05_0),.clk(gclk));
	jdff dff_A_X6eyEOAP9_0(.dout(w_dff_A_k0ryneHL6_0),.din(w_dff_A_X6eyEOAP9_0),.clk(gclk));
	jdff dff_A_k0ryneHL6_0(.dout(w_dff_A_AHlgEB6R8_0),.din(w_dff_A_k0ryneHL6_0),.clk(gclk));
	jdff dff_A_AHlgEB6R8_0(.dout(w_dff_A_nDuQPgox8_0),.din(w_dff_A_AHlgEB6R8_0),.clk(gclk));
	jdff dff_A_nDuQPgox8_0(.dout(w_dff_A_RkK6Y4jk9_0),.din(w_dff_A_nDuQPgox8_0),.clk(gclk));
	jdff dff_A_RkK6Y4jk9_0(.dout(w_dff_A_Mva2ZKpy1_0),.din(w_dff_A_RkK6Y4jk9_0),.clk(gclk));
	jdff dff_A_Mva2ZKpy1_0(.dout(w_dff_A_NM8nigdI3_0),.din(w_dff_A_Mva2ZKpy1_0),.clk(gclk));
	jdff dff_A_NM8nigdI3_0(.dout(w_dff_A_LSf5wbfi1_0),.din(w_dff_A_NM8nigdI3_0),.clk(gclk));
	jdff dff_A_LSf5wbfi1_0(.dout(w_dff_A_MlsONPWJ1_0),.din(w_dff_A_LSf5wbfi1_0),.clk(gclk));
	jdff dff_A_MlsONPWJ1_0(.dout(w_dff_A_7llmVHmU1_0),.din(w_dff_A_MlsONPWJ1_0),.clk(gclk));
	jdff dff_A_7llmVHmU1_0(.dout(w_dff_A_2EwzNxVk7_0),.din(w_dff_A_7llmVHmU1_0),.clk(gclk));
	jdff dff_A_2EwzNxVk7_0(.dout(w_dff_A_uyTbEu456_0),.din(w_dff_A_2EwzNxVk7_0),.clk(gclk));
	jdff dff_A_uyTbEu456_0(.dout(w_dff_A_73IGuFAb6_0),.din(w_dff_A_uyTbEu456_0),.clk(gclk));
	jdff dff_A_73IGuFAb6_0(.dout(w_dff_A_164mSSGv9_0),.din(w_dff_A_73IGuFAb6_0),.clk(gclk));
	jdff dff_A_164mSSGv9_0(.dout(w_dff_A_r8wBZGB90_0),.din(w_dff_A_164mSSGv9_0),.clk(gclk));
	jdff dff_A_r8wBZGB90_0(.dout(w_dff_A_zxTqd09L3_0),.din(w_dff_A_r8wBZGB90_0),.clk(gclk));
	jdff dff_A_zxTqd09L3_0(.dout(w_dff_A_ZfBg7EOm3_0),.din(w_dff_A_zxTqd09L3_0),.clk(gclk));
	jdff dff_A_ZfBg7EOm3_0(.dout(w_dff_A_eAoBdlQn5_0),.din(w_dff_A_ZfBg7EOm3_0),.clk(gclk));
	jdff dff_A_eAoBdlQn5_0(.dout(w_dff_A_UxAkDqS77_0),.din(w_dff_A_eAoBdlQn5_0),.clk(gclk));
	jdff dff_A_UxAkDqS77_0(.dout(w_dff_A_GUFhpf3f0_0),.din(w_dff_A_UxAkDqS77_0),.clk(gclk));
	jdff dff_A_GUFhpf3f0_0(.dout(w_dff_A_C2haGvds5_0),.din(w_dff_A_GUFhpf3f0_0),.clk(gclk));
	jdff dff_A_C2haGvds5_0(.dout(w_dff_A_iFd7aNBs5_0),.din(w_dff_A_C2haGvds5_0),.clk(gclk));
	jdff dff_A_iFd7aNBs5_0(.dout(w_dff_A_NUwyw1zB8_0),.din(w_dff_A_iFd7aNBs5_0),.clk(gclk));
	jdff dff_A_NUwyw1zB8_0(.dout(w_dff_A_oW4Z1SBK2_0),.din(w_dff_A_NUwyw1zB8_0),.clk(gclk));
	jdff dff_A_oW4Z1SBK2_0(.dout(w_dff_A_GkCBajpz2_0),.din(w_dff_A_oW4Z1SBK2_0),.clk(gclk));
	jdff dff_A_GkCBajpz2_0(.dout(w_dff_A_24eK7md31_0),.din(w_dff_A_GkCBajpz2_0),.clk(gclk));
	jdff dff_A_24eK7md31_0(.dout(w_dff_A_MQhPxitl4_0),.din(w_dff_A_24eK7md31_0),.clk(gclk));
	jdff dff_A_MQhPxitl4_0(.dout(w_dff_A_WemNEdjD0_0),.din(w_dff_A_MQhPxitl4_0),.clk(gclk));
	jdff dff_A_WemNEdjD0_0(.dout(w_dff_A_BjmyDr9S7_0),.din(w_dff_A_WemNEdjD0_0),.clk(gclk));
	jdff dff_A_BjmyDr9S7_0(.dout(w_dff_A_79a9Un1M3_0),.din(w_dff_A_BjmyDr9S7_0),.clk(gclk));
	jdff dff_A_79a9Un1M3_0(.dout(w_dff_A_ZgAAD1X23_0),.din(w_dff_A_79a9Un1M3_0),.clk(gclk));
	jdff dff_A_ZgAAD1X23_0(.dout(w_dff_A_W0hJcJng0_0),.din(w_dff_A_ZgAAD1X23_0),.clk(gclk));
	jdff dff_A_W0hJcJng0_0(.dout(w_dff_A_15VK5Byw3_0),.din(w_dff_A_W0hJcJng0_0),.clk(gclk));
	jdff dff_A_15VK5Byw3_0(.dout(w_dff_A_YXQp2haH1_0),.din(w_dff_A_15VK5Byw3_0),.clk(gclk));
	jdff dff_A_YXQp2haH1_0(.dout(w_dff_A_R013b8kh1_0),.din(w_dff_A_YXQp2haH1_0),.clk(gclk));
	jdff dff_A_R013b8kh1_0(.dout(w_dff_A_LcCBDxSe1_0),.din(w_dff_A_R013b8kh1_0),.clk(gclk));
	jdff dff_A_LcCBDxSe1_0(.dout(w_dff_A_5wIbKRAj5_0),.din(w_dff_A_LcCBDxSe1_0),.clk(gclk));
	jdff dff_A_5wIbKRAj5_0(.dout(w_dff_A_0QxsLgfB0_0),.din(w_dff_A_5wIbKRAj5_0),.clk(gclk));
	jdff dff_A_0QxsLgfB0_0(.dout(w_dff_A_3jFrOwCd1_0),.din(w_dff_A_0QxsLgfB0_0),.clk(gclk));
	jdff dff_A_3jFrOwCd1_0(.dout(w_dff_A_y9jp4VX77_0),.din(w_dff_A_3jFrOwCd1_0),.clk(gclk));
	jdff dff_A_y9jp4VX77_0(.dout(w_dff_A_4Qlnpg9M5_0),.din(w_dff_A_y9jp4VX77_0),.clk(gclk));
	jdff dff_A_4Qlnpg9M5_0(.dout(w_dff_A_uYaPzqZA3_0),.din(w_dff_A_4Qlnpg9M5_0),.clk(gclk));
	jdff dff_A_uYaPzqZA3_0(.dout(w_dff_A_kq1RummO1_0),.din(w_dff_A_uYaPzqZA3_0),.clk(gclk));
	jdff dff_A_kq1RummO1_0(.dout(w_dff_A_GfhJdHXK4_0),.din(w_dff_A_kq1RummO1_0),.clk(gclk));
	jdff dff_A_GfhJdHXK4_0(.dout(w_dff_A_vEYKv4WB4_0),.din(w_dff_A_GfhJdHXK4_0),.clk(gclk));
	jdff dff_A_vEYKv4WB4_0(.dout(w_dff_A_CDjyd4pp2_0),.din(w_dff_A_vEYKv4WB4_0),.clk(gclk));
	jdff dff_A_CDjyd4pp2_0(.dout(w_dff_A_jmRc3lFI4_0),.din(w_dff_A_CDjyd4pp2_0),.clk(gclk));
	jdff dff_A_jmRc3lFI4_0(.dout(w_dff_A_vw8shElw8_0),.din(w_dff_A_jmRc3lFI4_0),.clk(gclk));
	jdff dff_A_vw8shElw8_0(.dout(w_dff_A_y3Lzx6BD0_0),.din(w_dff_A_vw8shElw8_0),.clk(gclk));
	jdff dff_A_y3Lzx6BD0_0(.dout(w_dff_A_SP5SySG57_0),.din(w_dff_A_y3Lzx6BD0_0),.clk(gclk));
	jdff dff_A_SP5SySG57_0(.dout(w_dff_A_2moUPmxi5_0),.din(w_dff_A_SP5SySG57_0),.clk(gclk));
	jdff dff_A_2moUPmxi5_0(.dout(w_dff_A_X19Xa4qX4_0),.din(w_dff_A_2moUPmxi5_0),.clk(gclk));
	jdff dff_A_X19Xa4qX4_0(.dout(w_dff_A_DiDjfcNx9_0),.din(w_dff_A_X19Xa4qX4_0),.clk(gclk));
	jdff dff_A_DiDjfcNx9_0(.dout(w_dff_A_gJQ7MzSx4_0),.din(w_dff_A_DiDjfcNx9_0),.clk(gclk));
	jdff dff_A_gJQ7MzSx4_0(.dout(w_dff_A_frWp3oTl2_0),.din(w_dff_A_gJQ7MzSx4_0),.clk(gclk));
	jdff dff_A_frWp3oTl2_0(.dout(w_dff_A_zHUiaLRr5_0),.din(w_dff_A_frWp3oTl2_0),.clk(gclk));
	jdff dff_A_zHUiaLRr5_0(.dout(w_dff_A_EUKunzJq7_0),.din(w_dff_A_zHUiaLRr5_0),.clk(gclk));
	jdff dff_A_EUKunzJq7_0(.dout(w_dff_A_oQwMs0mW5_0),.din(w_dff_A_EUKunzJq7_0),.clk(gclk));
	jdff dff_A_oQwMs0mW5_0(.dout(w_dff_A_LSKIU1R72_0),.din(w_dff_A_oQwMs0mW5_0),.clk(gclk));
	jdff dff_A_LSKIU1R72_0(.dout(w_dff_A_YUFMEqV59_0),.din(w_dff_A_LSKIU1R72_0),.clk(gclk));
	jdff dff_A_YUFMEqV59_0(.dout(w_dff_A_T9pDQtWE9_0),.din(w_dff_A_YUFMEqV59_0),.clk(gclk));
	jdff dff_A_T9pDQtWE9_0(.dout(w_dff_A_t1ixKgFx5_0),.din(w_dff_A_T9pDQtWE9_0),.clk(gclk));
	jdff dff_A_t1ixKgFx5_0(.dout(w_dff_A_AGuJGsML4_0),.din(w_dff_A_t1ixKgFx5_0),.clk(gclk));
	jdff dff_A_AGuJGsML4_0(.dout(w_dff_A_Q2yISQDn5_0),.din(w_dff_A_AGuJGsML4_0),.clk(gclk));
	jdff dff_A_Q2yISQDn5_0(.dout(w_dff_A_6ukHgAXp8_0),.din(w_dff_A_Q2yISQDn5_0),.clk(gclk));
	jdff dff_A_6ukHgAXp8_0(.dout(w_dff_A_zxbKaZ869_0),.din(w_dff_A_6ukHgAXp8_0),.clk(gclk));
	jdff dff_A_zxbKaZ869_0(.dout(w_dff_A_24sfdZXr3_0),.din(w_dff_A_zxbKaZ869_0),.clk(gclk));
	jdff dff_A_24sfdZXr3_0(.dout(w_dff_A_GhuuM4nu2_0),.din(w_dff_A_24sfdZXr3_0),.clk(gclk));
	jdff dff_A_GhuuM4nu2_0(.dout(w_dff_A_vKtwxVRJ5_0),.din(w_dff_A_GhuuM4nu2_0),.clk(gclk));
	jdff dff_A_vKtwxVRJ5_0(.dout(w_dff_A_JXDjRnst9_0),.din(w_dff_A_vKtwxVRJ5_0),.clk(gclk));
	jdff dff_A_JXDjRnst9_0(.dout(w_dff_A_4TbC2bHw6_0),.din(w_dff_A_JXDjRnst9_0),.clk(gclk));
	jdff dff_A_4TbC2bHw6_0(.dout(w_dff_A_uYSMAWWk0_0),.din(w_dff_A_4TbC2bHw6_0),.clk(gclk));
	jdff dff_A_uYSMAWWk0_0(.dout(w_dff_A_SJgKgLkE7_0),.din(w_dff_A_uYSMAWWk0_0),.clk(gclk));
	jdff dff_A_SJgKgLkE7_0(.dout(w_dff_A_VTeFanvL9_0),.din(w_dff_A_SJgKgLkE7_0),.clk(gclk));
	jdff dff_A_VTeFanvL9_0(.dout(w_dff_A_sMHiCaPq4_0),.din(w_dff_A_VTeFanvL9_0),.clk(gclk));
	jdff dff_A_sMHiCaPq4_0(.dout(w_dff_A_6janH4c82_0),.din(w_dff_A_sMHiCaPq4_0),.clk(gclk));
	jdff dff_A_6janH4c82_0(.dout(w_dff_A_7jRGideT8_0),.din(w_dff_A_6janH4c82_0),.clk(gclk));
	jdff dff_A_7jRGideT8_0(.dout(w_dff_A_dO38tszJ1_0),.din(w_dff_A_7jRGideT8_0),.clk(gclk));
	jdff dff_A_dO38tszJ1_0(.dout(w_dff_A_ruoAbtlZ9_0),.din(w_dff_A_dO38tszJ1_0),.clk(gclk));
	jdff dff_A_ruoAbtlZ9_0(.dout(w_dff_A_4fiXhAXU2_0),.din(w_dff_A_ruoAbtlZ9_0),.clk(gclk));
	jdff dff_A_4fiXhAXU2_0(.dout(w_dff_A_egevUpLL9_0),.din(w_dff_A_4fiXhAXU2_0),.clk(gclk));
	jdff dff_A_egevUpLL9_0(.dout(w_dff_A_Nhdw7Kox2_0),.din(w_dff_A_egevUpLL9_0),.clk(gclk));
	jdff dff_A_Nhdw7Kox2_0(.dout(w_dff_A_rhyNALCV1_0),.din(w_dff_A_Nhdw7Kox2_0),.clk(gclk));
	jdff dff_A_rhyNALCV1_0(.dout(w_dff_A_E9BTpH219_0),.din(w_dff_A_rhyNALCV1_0),.clk(gclk));
	jdff dff_A_E9BTpH219_0(.dout(w_dff_A_vKsq5QJb0_0),.din(w_dff_A_E9BTpH219_0),.clk(gclk));
	jdff dff_A_vKsq5QJb0_0(.dout(w_dff_A_AgztGxiK8_0),.din(w_dff_A_vKsq5QJb0_0),.clk(gclk));
	jdff dff_A_AgztGxiK8_0(.dout(w_dff_A_t4IJCiJa6_0),.din(w_dff_A_AgztGxiK8_0),.clk(gclk));
	jdff dff_A_t4IJCiJa6_0(.dout(w_dff_A_N2ne8qw09_0),.din(w_dff_A_t4IJCiJa6_0),.clk(gclk));
	jdff dff_A_N2ne8qw09_0(.dout(w_dff_A_G7kqdhof8_0),.din(w_dff_A_N2ne8qw09_0),.clk(gclk));
	jdff dff_A_G7kqdhof8_0(.dout(w_dff_A_FBvnzSKB4_0),.din(w_dff_A_G7kqdhof8_0),.clk(gclk));
	jdff dff_A_FBvnzSKB4_0(.dout(w_dff_A_L0pTsOk01_0),.din(w_dff_A_FBvnzSKB4_0),.clk(gclk));
	jdff dff_A_L0pTsOk01_0(.dout(w_dff_A_i7MpsIXU1_0),.din(w_dff_A_L0pTsOk01_0),.clk(gclk));
	jdff dff_A_i7MpsIXU1_0(.dout(w_dff_A_Nx3X5url6_0),.din(w_dff_A_i7MpsIXU1_0),.clk(gclk));
	jdff dff_A_Nx3X5url6_0(.dout(w_dff_A_fUFtcc7W4_0),.din(w_dff_A_Nx3X5url6_0),.clk(gclk));
	jdff dff_A_fUFtcc7W4_0(.dout(w_dff_A_fKGTRAXk4_0),.din(w_dff_A_fUFtcc7W4_0),.clk(gclk));
	jdff dff_A_fKGTRAXk4_0(.dout(w_dff_A_TrFMigrB8_0),.din(w_dff_A_fKGTRAXk4_0),.clk(gclk));
	jdff dff_A_TrFMigrB8_0(.dout(w_dff_A_oY4d4AN77_0),.din(w_dff_A_TrFMigrB8_0),.clk(gclk));
	jdff dff_A_oY4d4AN77_0(.dout(w_dff_A_4rHXoMaq5_0),.din(w_dff_A_oY4d4AN77_0),.clk(gclk));
	jdff dff_A_4rHXoMaq5_0(.dout(w_dff_A_ne5OJtTS8_0),.din(w_dff_A_4rHXoMaq5_0),.clk(gclk));
	jdff dff_A_ne5OJtTS8_0(.dout(w_dff_A_TybogAPB0_0),.din(w_dff_A_ne5OJtTS8_0),.clk(gclk));
	jdff dff_A_TybogAPB0_0(.dout(w_dff_A_7an3FYwm6_0),.din(w_dff_A_TybogAPB0_0),.clk(gclk));
	jdff dff_A_7an3FYwm6_0(.dout(w_dff_A_KVbc8xCN0_0),.din(w_dff_A_7an3FYwm6_0),.clk(gclk));
	jdff dff_A_KVbc8xCN0_0(.dout(w_dff_A_LfXOHS0O4_0),.din(w_dff_A_KVbc8xCN0_0),.clk(gclk));
	jdff dff_A_LfXOHS0O4_0(.dout(w_dff_A_4NFpnNuN3_0),.din(w_dff_A_LfXOHS0O4_0),.clk(gclk));
	jdff dff_A_4NFpnNuN3_0(.dout(w_dff_A_y4WunLpr2_0),.din(w_dff_A_4NFpnNuN3_0),.clk(gclk));
	jdff dff_A_y4WunLpr2_0(.dout(w_dff_A_rkjJcYFu4_0),.din(w_dff_A_y4WunLpr2_0),.clk(gclk));
	jdff dff_A_rkjJcYFu4_0(.dout(w_dff_A_btioAenC8_0),.din(w_dff_A_rkjJcYFu4_0),.clk(gclk));
	jdff dff_A_btioAenC8_0(.dout(w_dff_A_zMWFq7u72_0),.din(w_dff_A_btioAenC8_0),.clk(gclk));
	jdff dff_A_zMWFq7u72_0(.dout(w_dff_A_5J0aoye44_0),.din(w_dff_A_zMWFq7u72_0),.clk(gclk));
	jdff dff_A_5J0aoye44_0(.dout(w_dff_A_JnTC9t918_0),.din(w_dff_A_5J0aoye44_0),.clk(gclk));
	jdff dff_A_JnTC9t918_0(.dout(w_dff_A_fuigrAIF3_0),.din(w_dff_A_JnTC9t918_0),.clk(gclk));
	jdff dff_A_fuigrAIF3_0(.dout(w_dff_A_k0vpDHaf5_0),.din(w_dff_A_fuigrAIF3_0),.clk(gclk));
	jdff dff_A_k0vpDHaf5_0(.dout(w_dff_A_n2Og61yG7_0),.din(w_dff_A_k0vpDHaf5_0),.clk(gclk));
	jdff dff_A_n2Og61yG7_0(.dout(w_dff_A_BwaUDQlb7_0),.din(w_dff_A_n2Og61yG7_0),.clk(gclk));
	jdff dff_A_BwaUDQlb7_0(.dout(w_dff_A_jvIRd8RD9_0),.din(w_dff_A_BwaUDQlb7_0),.clk(gclk));
	jdff dff_A_jvIRd8RD9_0(.dout(w_dff_A_t6DmL0hs4_0),.din(w_dff_A_jvIRd8RD9_0),.clk(gclk));
	jdff dff_A_t6DmL0hs4_0(.dout(w_dff_A_vKttdw0P8_0),.din(w_dff_A_t6DmL0hs4_0),.clk(gclk));
	jdff dff_A_vKttdw0P8_0(.dout(w_dff_A_zil5QNhd3_0),.din(w_dff_A_vKttdw0P8_0),.clk(gclk));
	jdff dff_A_zil5QNhd3_0(.dout(w_dff_A_eChi8Hp90_0),.din(w_dff_A_zil5QNhd3_0),.clk(gclk));
	jdff dff_A_eChi8Hp90_0(.dout(w_dff_A_h8NfFE6T9_0),.din(w_dff_A_eChi8Hp90_0),.clk(gclk));
	jdff dff_A_h8NfFE6T9_0(.dout(w_dff_A_WxOwicXM7_0),.din(w_dff_A_h8NfFE6T9_0),.clk(gclk));
	jdff dff_A_WxOwicXM7_0(.dout(w_dff_A_53ozTV0t8_0),.din(w_dff_A_WxOwicXM7_0),.clk(gclk));
	jdff dff_A_53ozTV0t8_0(.dout(w_dff_A_sHAhLXI65_0),.din(w_dff_A_53ozTV0t8_0),.clk(gclk));
	jdff dff_A_sHAhLXI65_0(.dout(w_dff_A_p6cK4d8e3_0),.din(w_dff_A_sHAhLXI65_0),.clk(gclk));
	jdff dff_A_p6cK4d8e3_0(.dout(w_dff_A_cNAUyyp40_0),.din(w_dff_A_p6cK4d8e3_0),.clk(gclk));
	jdff dff_A_cNAUyyp40_0(.dout(w_dff_A_B0ajDMg55_0),.din(w_dff_A_cNAUyyp40_0),.clk(gclk));
	jdff dff_A_B0ajDMg55_0(.dout(w_dff_A_bDDsIjFK5_0),.din(w_dff_A_B0ajDMg55_0),.clk(gclk));
	jdff dff_A_bDDsIjFK5_0(.dout(w_dff_A_zWmd4dhB0_0),.din(w_dff_A_bDDsIjFK5_0),.clk(gclk));
	jdff dff_A_zWmd4dhB0_0(.dout(w_dff_A_dFzYkT2w9_0),.din(w_dff_A_zWmd4dhB0_0),.clk(gclk));
	jdff dff_A_dFzYkT2w9_0(.dout(w_dff_A_WwnrpaUb3_0),.din(w_dff_A_dFzYkT2w9_0),.clk(gclk));
	jdff dff_A_WwnrpaUb3_0(.dout(w_dff_A_jCq1zhJR6_0),.din(w_dff_A_WwnrpaUb3_0),.clk(gclk));
	jdff dff_A_jCq1zhJR6_0(.dout(w_dff_A_3DB2Aomd0_0),.din(w_dff_A_jCq1zhJR6_0),.clk(gclk));
	jdff dff_A_3DB2Aomd0_0(.dout(w_dff_A_0MeMQ0W84_0),.din(w_dff_A_3DB2Aomd0_0),.clk(gclk));
	jdff dff_A_0MeMQ0W84_0(.dout(w_dff_A_rMxVGIVT7_0),.din(w_dff_A_0MeMQ0W84_0),.clk(gclk));
	jdff dff_A_rMxVGIVT7_0(.dout(w_dff_A_xWgZWwKi6_0),.din(w_dff_A_rMxVGIVT7_0),.clk(gclk));
	jdff dff_A_xWgZWwKi6_0(.dout(w_dff_A_OxDGxcuy0_0),.din(w_dff_A_xWgZWwKi6_0),.clk(gclk));
	jdff dff_A_OxDGxcuy0_0(.dout(w_dff_A_BAHS0BlU4_0),.din(w_dff_A_OxDGxcuy0_0),.clk(gclk));
	jdff dff_A_BAHS0BlU4_0(.dout(w_dff_A_1ur5BZkO0_0),.din(w_dff_A_BAHS0BlU4_0),.clk(gclk));
	jdff dff_A_1ur5BZkO0_0(.dout(w_dff_A_zU2Az30p3_0),.din(w_dff_A_1ur5BZkO0_0),.clk(gclk));
	jdff dff_A_zU2Az30p3_0(.dout(w_dff_A_pxdk0SaI5_0),.din(w_dff_A_zU2Az30p3_0),.clk(gclk));
	jdff dff_A_pxdk0SaI5_0(.dout(w_dff_A_IufjhC9z3_0),.din(w_dff_A_pxdk0SaI5_0),.clk(gclk));
	jdff dff_A_IufjhC9z3_0(.dout(w_dff_A_bUxsefr51_0),.din(w_dff_A_IufjhC9z3_0),.clk(gclk));
	jdff dff_A_bUxsefr51_0(.dout(w_dff_A_Nfv1pWz89_0),.din(w_dff_A_bUxsefr51_0),.clk(gclk));
	jdff dff_A_Nfv1pWz89_0(.dout(w_dff_A_Mi6vWPQd2_0),.din(w_dff_A_Nfv1pWz89_0),.clk(gclk));
	jdff dff_A_Mi6vWPQd2_0(.dout(w_dff_A_iZRgV53k8_0),.din(w_dff_A_Mi6vWPQd2_0),.clk(gclk));
	jdff dff_A_iZRgV53k8_0(.dout(w_dff_A_y9cqJ74O8_0),.din(w_dff_A_iZRgV53k8_0),.clk(gclk));
	jdff dff_A_y9cqJ74O8_0(.dout(w_dff_A_Yb7ypwXw3_0),.din(w_dff_A_y9cqJ74O8_0),.clk(gclk));
	jdff dff_A_Yb7ypwXw3_0(.dout(w_dff_A_ObOVeJRp9_0),.din(w_dff_A_Yb7ypwXw3_0),.clk(gclk));
	jdff dff_A_ObOVeJRp9_0(.dout(w_dff_A_KrQIAAHE3_0),.din(w_dff_A_ObOVeJRp9_0),.clk(gclk));
	jdff dff_A_KrQIAAHE3_0(.dout(w_dff_A_aoGDhvui2_0),.din(w_dff_A_KrQIAAHE3_0),.clk(gclk));
	jdff dff_A_aoGDhvui2_0(.dout(w_dff_A_KM4GCFim7_0),.din(w_dff_A_aoGDhvui2_0),.clk(gclk));
	jdff dff_A_KM4GCFim7_0(.dout(w_dff_A_kGuuD0dn6_0),.din(w_dff_A_KM4GCFim7_0),.clk(gclk));
	jdff dff_A_kGuuD0dn6_0(.dout(w_dff_A_TpFMWBtX0_0),.din(w_dff_A_kGuuD0dn6_0),.clk(gclk));
	jdff dff_A_TpFMWBtX0_0(.dout(w_dff_A_8ByzbrMU2_0),.din(w_dff_A_TpFMWBtX0_0),.clk(gclk));
	jdff dff_A_8ByzbrMU2_0(.dout(w_dff_A_AabcLQEi4_0),.din(w_dff_A_8ByzbrMU2_0),.clk(gclk));
	jdff dff_A_AabcLQEi4_0(.dout(w_dff_A_rTZdbN3s7_0),.din(w_dff_A_AabcLQEi4_0),.clk(gclk));
	jdff dff_A_rTZdbN3s7_0(.dout(w_dff_A_ck0PEhff7_0),.din(w_dff_A_rTZdbN3s7_0),.clk(gclk));
	jdff dff_A_ck0PEhff7_0(.dout(w_dff_A_cpY2kb4V7_0),.din(w_dff_A_ck0PEhff7_0),.clk(gclk));
	jdff dff_A_cpY2kb4V7_0(.dout(w_dff_A_p1PukFDF4_0),.din(w_dff_A_cpY2kb4V7_0),.clk(gclk));
	jdff dff_A_p1PukFDF4_0(.dout(w_dff_A_mVDadcX61_0),.din(w_dff_A_p1PukFDF4_0),.clk(gclk));
	jdff dff_A_mVDadcX61_0(.dout(w_dff_A_dy2I0UeI4_0),.din(w_dff_A_mVDadcX61_0),.clk(gclk));
	jdff dff_A_dy2I0UeI4_0(.dout(w_dff_A_cLy6gKfo5_0),.din(w_dff_A_dy2I0UeI4_0),.clk(gclk));
	jdff dff_A_cLy6gKfo5_0(.dout(w_dff_A_PRxsZe801_0),.din(w_dff_A_cLy6gKfo5_0),.clk(gclk));
	jdff dff_A_PRxsZe801_0(.dout(w_dff_A_sicOs0hc7_0),.din(w_dff_A_PRxsZe801_0),.clk(gclk));
	jdff dff_A_sicOs0hc7_0(.dout(w_dff_A_dSVYS6Sb0_0),.din(w_dff_A_sicOs0hc7_0),.clk(gclk));
	jdff dff_A_dSVYS6Sb0_0(.dout(w_dff_A_Y9MPNg2g7_0),.din(w_dff_A_dSVYS6Sb0_0),.clk(gclk));
	jdff dff_A_Y9MPNg2g7_0(.dout(w_dff_A_ENC5HKRE6_0),.din(w_dff_A_Y9MPNg2g7_0),.clk(gclk));
	jdff dff_A_ENC5HKRE6_0(.dout(w_dff_A_rTDKpKiJ5_0),.din(w_dff_A_ENC5HKRE6_0),.clk(gclk));
	jdff dff_A_rTDKpKiJ5_0(.dout(w_dff_A_n1KDeIFP5_0),.din(w_dff_A_rTDKpKiJ5_0),.clk(gclk));
	jdff dff_A_n1KDeIFP5_0(.dout(w_dff_A_QrykYaRi5_0),.din(w_dff_A_n1KDeIFP5_0),.clk(gclk));
	jdff dff_A_QrykYaRi5_0(.dout(w_dff_A_tX8FSWOw9_0),.din(w_dff_A_QrykYaRi5_0),.clk(gclk));
	jdff dff_A_tX8FSWOw9_0(.dout(w_dff_A_unj9VdsQ4_0),.din(w_dff_A_tX8FSWOw9_0),.clk(gclk));
	jdff dff_A_unj9VdsQ4_0(.dout(w_dff_A_y7AeHnxY2_0),.din(w_dff_A_unj9VdsQ4_0),.clk(gclk));
	jdff dff_A_y7AeHnxY2_0(.dout(w_dff_A_suiUbgLz3_0),.din(w_dff_A_y7AeHnxY2_0),.clk(gclk));
	jdff dff_A_suiUbgLz3_0(.dout(w_dff_A_Nt1BUMao2_0),.din(w_dff_A_suiUbgLz3_0),.clk(gclk));
	jdff dff_A_Nt1BUMao2_0(.dout(w_dff_A_E1qwy4311_0),.din(w_dff_A_Nt1BUMao2_0),.clk(gclk));
	jdff dff_A_E1qwy4311_0(.dout(w_dff_A_FEoc5rfZ4_0),.din(w_dff_A_E1qwy4311_0),.clk(gclk));
	jdff dff_A_FEoc5rfZ4_0(.dout(w_dff_A_zAIw19Ld1_0),.din(w_dff_A_FEoc5rfZ4_0),.clk(gclk));
	jdff dff_A_zAIw19Ld1_0(.dout(w_dff_A_gbW1I6Xw7_0),.din(w_dff_A_zAIw19Ld1_0),.clk(gclk));
	jdff dff_A_gbW1I6Xw7_0(.dout(w_dff_A_fjV7yB6Y1_0),.din(w_dff_A_gbW1I6Xw7_0),.clk(gclk));
	jdff dff_A_fjV7yB6Y1_0(.dout(w_dff_A_u9eCVOjx8_0),.din(w_dff_A_fjV7yB6Y1_0),.clk(gclk));
	jdff dff_A_u9eCVOjx8_0(.dout(w_dff_A_vxbIwSN15_0),.din(w_dff_A_u9eCVOjx8_0),.clk(gclk));
	jdff dff_A_vxbIwSN15_0(.dout(w_dff_A_habLXnNM8_0),.din(w_dff_A_vxbIwSN15_0),.clk(gclk));
	jdff dff_A_habLXnNM8_0(.dout(w_dff_A_HpcRdr2p2_0),.din(w_dff_A_habLXnNM8_0),.clk(gclk));
	jdff dff_A_HpcRdr2p2_0(.dout(w_dff_A_JpdZBD5e9_0),.din(w_dff_A_HpcRdr2p2_0),.clk(gclk));
	jdff dff_A_JpdZBD5e9_0(.dout(w_dff_A_CxWhO9FU8_0),.din(w_dff_A_JpdZBD5e9_0),.clk(gclk));
	jdff dff_A_CxWhO9FU8_0(.dout(w_dff_A_uZPd6kIb3_0),.din(w_dff_A_CxWhO9FU8_0),.clk(gclk));
	jdff dff_A_uZPd6kIb3_0(.dout(w_dff_A_mypM8eLS6_0),.din(w_dff_A_uZPd6kIb3_0),.clk(gclk));
	jdff dff_A_mypM8eLS6_0(.dout(w_dff_A_426B4d8m3_0),.din(w_dff_A_mypM8eLS6_0),.clk(gclk));
	jdff dff_A_426B4d8m3_0(.dout(w_dff_A_hYPFUOh12_0),.din(w_dff_A_426B4d8m3_0),.clk(gclk));
	jdff dff_A_hYPFUOh12_0(.dout(w_dff_A_jPWtj9QZ3_0),.din(w_dff_A_hYPFUOh12_0),.clk(gclk));
	jdff dff_A_jPWtj9QZ3_0(.dout(w_dff_A_pHcPiXMP2_0),.din(w_dff_A_jPWtj9QZ3_0),.clk(gclk));
	jdff dff_A_pHcPiXMP2_0(.dout(w_dff_A_0brnFmns3_0),.din(w_dff_A_pHcPiXMP2_0),.clk(gclk));
	jdff dff_A_0brnFmns3_0(.dout(w_dff_A_i4dkcnEv4_0),.din(w_dff_A_0brnFmns3_0),.clk(gclk));
	jdff dff_A_i4dkcnEv4_0(.dout(w_dff_A_1ZsJQvPo9_0),.din(w_dff_A_i4dkcnEv4_0),.clk(gclk));
	jdff dff_A_1ZsJQvPo9_0(.dout(w_dff_A_CfvqN9Yh0_0),.din(w_dff_A_1ZsJQvPo9_0),.clk(gclk));
	jdff dff_A_CfvqN9Yh0_0(.dout(w_dff_A_gVxwUDTJ2_0),.din(w_dff_A_CfvqN9Yh0_0),.clk(gclk));
	jdff dff_A_gVxwUDTJ2_0(.dout(w_dff_A_VSKG0pS21_0),.din(w_dff_A_gVxwUDTJ2_0),.clk(gclk));
	jdff dff_A_VSKG0pS21_0(.dout(w_dff_A_m6FTD2XC1_0),.din(w_dff_A_VSKG0pS21_0),.clk(gclk));
	jdff dff_A_m6FTD2XC1_0(.dout(w_dff_A_IUnjpRHq6_0),.din(w_dff_A_m6FTD2XC1_0),.clk(gclk));
	jdff dff_A_IUnjpRHq6_0(.dout(result127),.din(w_dff_A_IUnjpRHq6_0),.clk(gclk));
	jdff dff_A_J7blzP2R6_2(.dout(w_dff_A_PyOOYhAQ5_0),.din(w_dff_A_J7blzP2R6_2),.clk(gclk));
	jdff dff_A_PyOOYhAQ5_0(.dout(address1),.din(w_dff_A_PyOOYhAQ5_0),.clk(gclk));
endmodule

