/*

c5315:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jcb: 486
	jdff: 3236
	jand: 606

Summary:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jcb: 486
	jdff: 3236
	jand: 606
*/

module c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G4_0;
	wire [1:0] w_G11_0;
	wire [1:0] w_G14_0;
	wire [1:0] w_G17_0;
	wire [1:0] w_G20_0;
	wire [1:0] w_G37_0;
	wire [1:0] w_G40_0;
	wire [1:0] w_G43_0;
	wire [1:0] w_G46_0;
	wire [1:0] w_G49_0;
	wire [2:0] w_G54_0;
	wire [1:0] w_G61_0;
	wire [1:0] w_G64_0;
	wire [1:0] w_G67_0;
	wire [1:0] w_G70_0;
	wire [1:0] w_G73_0;
	wire [1:0] w_G76_0;
	wire [1:0] w_G91_0;
	wire [1:0] w_G100_0;
	wire [1:0] w_G103_0;
	wire [1:0] w_G106_0;
	wire [1:0] w_G109_0;
	wire [1:0] w_G123_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G137_2;
	wire [2:0] w_G137_3;
	wire [2:0] w_G137_4;
	wire [2:0] w_G137_5;
	wire [2:0] w_G137_6;
	wire [2:0] w_G137_7;
	wire [2:0] w_G137_8;
	wire [1:0] w_G137_9;
	wire [2:0] w_G141_0;
	wire [2:0] w_G141_1;
	wire [2:0] w_G141_2;
	wire [1:0] w_G146_0;
	wire [1:0] w_G149_0;
	wire [1:0] w_G152_0;
	wire [1:0] w_G155_0;
	wire [1:0] w_G158_0;
	wire [1:0] w_G161_0;
	wire [1:0] w_G164_0;
	wire [1:0] w_G167_0;
	wire [1:0] w_G170_0;
	wire [1:0] w_G173_0;
	wire [1:0] w_G182_0;
	wire [1:0] w_G185_0;
	wire [1:0] w_G188_0;
	wire [1:0] w_G191_0;
	wire [1:0] w_G194_0;
	wire [1:0] w_G197_0;
	wire [1:0] w_G200_0;
	wire [1:0] w_G203_0;
	wire [2:0] w_G206_0;
	wire [2:0] w_G206_1;
	wire [2:0] w_G210_0;
	wire [2:0] w_G210_1;
	wire [1:0] w_G210_2;
	wire [2:0] w_G218_0;
	wire [2:0] w_G218_1;
	wire [1:0] w_G218_2;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [1:0] w_G226_2;
	wire [2:0] w_G234_0;
	wire [2:0] w_G234_1;
	wire [1:0] w_G234_2;
	wire [2:0] w_G242_0;
	wire [1:0] w_G242_1;
	wire [1:0] w_G245_0;
	wire [2:0] w_G248_0;
	wire [2:0] w_G248_1;
	wire [2:0] w_G248_2;
	wire [2:0] w_G248_3;
	wire [2:0] w_G248_4;
	wire [2:0] w_G248_5;
	wire [2:0] w_G251_0;
	wire [2:0] w_G251_1;
	wire [2:0] w_G251_2;
	wire [2:0] w_G251_3;
	wire [2:0] w_G251_4;
	wire [1:0] w_G251_5;
	wire [2:0] w_G254_0;
	wire [1:0] w_G254_1;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [1:0] w_G257_2;
	wire [2:0] w_G265_0;
	wire [2:0] w_G265_1;
	wire [2:0] w_G273_0;
	wire [2:0] w_G273_1;
	wire [1:0] w_G273_2;
	wire [2:0] w_G281_0;
	wire [2:0] w_G281_1;
	wire [1:0] w_G281_2;
	wire [1:0] w_G289_0;
	wire [2:0] w_G293_0;
	wire [2:0] w_G299_0;
	wire [2:0] w_G302_0;
	wire [2:0] w_G308_0;
	wire [2:0] w_G308_1;
	wire [2:0] w_G316_0;
	wire [1:0] w_G316_1;
	wire [2:0] w_G324_0;
	wire [2:0] w_G324_1;
	wire [1:0] w_G331_0;
	wire [2:0] w_G332_0;
	wire [2:0] w_G332_1;
	wire [2:0] w_G332_2;
	wire [2:0] w_G332_3;
	wire [2:0] w_G335_0;
	wire [1:0] w_G338_0;
	wire [2:0] w_G341_0;
	wire [2:0] w_G341_1;
	wire [2:0] w_G341_2;
	wire [1:0] w_G348_0;
	wire [2:0] w_G351_0;
	wire [2:0] w_G351_1;
	wire [2:0] w_G351_2;
	wire [1:0] w_G358_0;
	wire [2:0] w_G361_0;
	wire [1:0] w_G361_1;
	wire [1:0] w_G366_0;
	wire [1:0] w_G369_0;
	wire [2:0] w_G374_0;
	wire [2:0] w_G374_1;
	wire [2:0] w_G389_0;
	wire [2:0] w_G389_1;
	wire [2:0] w_G400_0;
	wire [2:0] w_G400_1;
	wire [2:0] w_G411_0;
	wire [2:0] w_G411_1;
	wire [1:0] w_G411_2;
	wire [2:0] w_G422_0;
	wire [1:0] w_G422_1;
	wire [2:0] w_G435_0;
	wire [2:0] w_G435_1;
	wire [2:0] w_G446_0;
	wire [2:0] w_G446_1;
	wire [2:0] w_G457_0;
	wire [2:0] w_G457_1;
	wire [2:0] w_G468_0;
	wire [2:0] w_G468_1;
	wire [2:0] w_G479_0;
	wire [2:0] w_G490_0;
	wire [1:0] w_G490_1;
	wire [2:0] w_G503_0;
	wire [2:0] w_G503_1;
	wire [1:0] w_G503_2;
	wire [2:0] w_G514_0;
	wire [2:0] w_G514_1;
	wire [1:0] w_G514_2;
	wire [2:0] w_G523_0;
	wire [2:0] w_G523_1;
	wire [2:0] w_G534_0;
	wire [2:0] w_G534_1;
	wire [1:0] w_G534_2;
	wire [2:0] w_G545_0;
	wire [2:0] w_G549_0;
	wire [1:0] w_G552_0;
	wire [1:0] w_G559_0;
	wire [1:0] w_G562_0;
	wire [2:0] w_G1497_0;
	wire [2:0] w_G1689_0;
	wire [2:0] w_G1689_1;
	wire [2:0] w_G1689_2;
	wire [2:0] w_G1689_3;
	wire [2:0] w_G1689_4;
	wire [1:0] w_G1689_5;
	wire [2:0] w_G1690_0;
	wire [1:0] w_G1690_1;
	wire [2:0] w_G1691_0;
	wire [2:0] w_G1691_1;
	wire [2:0] w_G1691_2;
	wire [2:0] w_G1691_3;
	wire [2:0] w_G1691_4;
	wire [1:0] w_G1691_5;
	wire [2:0] w_G1694_0;
	wire [1:0] w_G1694_1;
	wire [2:0] w_G2174_0;
	wire [2:0] w_G2358_0;
	wire [2:0] w_G2358_1;
	wire [2:0] w_G2358_2;
	wire [1:0] w_G3173_0;
	wire [2:0] w_G3546_0;
	wire [2:0] w_G3546_1;
	wire [2:0] w_G3546_2;
	wire [2:0] w_G3546_3;
	wire [2:0] w_G3546_4;
	wire [1:0] w_G3546_5;
	wire [2:0] w_G3548_0;
	wire [2:0] w_G3548_1;
	wire [2:0] w_G3548_2;
	wire [2:0] w_G3548_3;
	wire [2:0] w_G3548_4;
	wire [1:0] w_G3552_0;
	wire [1:0] w_G3717_0;
	wire [2:0] w_G3724_0;
	wire [2:0] w_G4087_0;
	wire [2:0] w_G4087_1;
	wire [2:0] w_G4087_2;
	wire [2:0] w_G4087_3;
	wire [2:0] w_G4087_4;
	wire [2:0] w_G4088_0;
	wire [2:0] w_G4088_1;
	wire [2:0] w_G4088_2;
	wire [2:0] w_G4088_3;
	wire [2:0] w_G4088_4;
	wire [2:0] w_G4088_5;
	wire [2:0] w_G4088_6;
	wire [2:0] w_G4088_7;
	wire [2:0] w_G4088_8;
	wire [2:0] w_G4088_9;
	wire [2:0] w_G4089_0;
	wire [2:0] w_G4089_1;
	wire [2:0] w_G4089_2;
	wire [2:0] w_G4089_3;
	wire [2:0] w_G4089_4;
	wire [2:0] w_G4089_5;
	wire [2:0] w_G4089_6;
	wire [2:0] w_G4089_7;
	wire [2:0] w_G4089_8;
	wire [2:0] w_G4089_9;
	wire [2:0] w_G4090_0;
	wire [2:0] w_G4090_1;
	wire [2:0] w_G4090_2;
	wire [2:0] w_G4090_3;
	wire [2:0] w_G4090_4;
	wire [2:0] w_G4091_0;
	wire [2:0] w_G4091_1;
	wire [2:0] w_G4091_2;
	wire [2:0] w_G4091_3;
	wire [2:0] w_G4091_4;
	wire [2:0] w_G4091_5;
	wire [1:0] w_G4091_6;
	wire [2:0] w_G4092_0;
	wire [2:0] w_G4092_1;
	wire [2:0] w_G4092_2;
	wire [2:0] w_G4092_3;
	wire [2:0] w_G4092_4;
	wire [2:0] w_G4092_5;
	wire [2:0] w_G4092_6;
	wire [2:0] w_G4092_7;
	wire [2:0] w_G4092_8;
	wire [2:0] w_G4092_9;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire [2:0] w_G809_0;
	wire [2:0] w_G809_1;
	wire [2:0] w_G809_2;
	wire [1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G623_0;
	wire G623_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G998_0;
	wire G998_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G865_0;
	wire G865_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire [1:0] w_n316_0;
	wire [1:0] w_n318_0;
	wire [2:0] w_n326_0;
	wire [2:0] w_n326_1;
	wire [1:0] w_n326_2;
	wire [1:0] w_n333_0;
	wire [1:0] w_n336_0;
	wire [1:0] w_n361_0;
	wire [1:0] w_n365_0;
	wire [2:0] w_n366_0;
	wire [2:0] w_n366_1;
	wire [2:0] w_n369_0;
	wire [2:0] w_n369_1;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [2:0] w_n374_0;
	wire [1:0] w_n374_1;
	wire [2:0] w_n375_0;
	wire [2:0] w_n375_1;
	wire [2:0] w_n375_2;
	wire [2:0] w_n375_3;
	wire [2:0] w_n375_4;
	wire [2:0] w_n377_0;
	wire [1:0] w_n377_1;
	wire [2:0] w_n378_0;
	wire [2:0] w_n378_1;
	wire [2:0] w_n378_2;
	wire [2:0] w_n378_3;
	wire [2:0] w_n378_4;
	wire [1:0] w_n386_0;
	wire [2:0] w_n387_0;
	wire [1:0] w_n387_1;
	wire [2:0] w_n389_0;
	wire [1:0] w_n389_1;
	wire [1:0] w_n397_0;
	wire [1:0] w_n401_0;
	wire [2:0] w_n402_0;
	wire [2:0] w_n406_0;
	wire [2:0] w_n406_1;
	wire [2:0] w_n406_2;
	wire [2:0] w_n406_3;
	wire [2:0] w_n406_4;
	wire [1:0] w_n406_5;
	wire [2:0] w_n408_0;
	wire [2:0] w_n408_1;
	wire [2:0] w_n408_2;
	wire [2:0] w_n408_3;
	wire [2:0] w_n408_4;
	wire [2:0] w_n408_5;
	wire [2:0] w_n412_0;
	wire [1:0] w_n414_0;
	wire [1:0] w_n415_0;
	wire [2:0] w_n423_0;
	wire [2:0] w_n425_0;
	wire [2:0] w_n428_0;
	wire [1:0] w_n428_1;
	wire [1:0] w_n429_0;
	wire [2:0] w_n433_0;
	wire [2:0] w_n435_0;
	wire [2:0] w_n435_1;
	wire [1:0] w_n435_2;
	wire [1:0] w_n437_0;
	wire [1:0] w_n445_0;
	wire [2:0] w_n449_0;
	wire [2:0] w_n449_1;
	wire [2:0] w_n451_0;
	wire [1:0] w_n459_0;
	wire [2:0] w_n460_0;
	wire [2:0] w_n460_1;
	wire [2:0] w_n462_0;
	wire [1:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [2:0] w_n471_1;
	wire [2:0] w_n473_0;
	wire [1:0] w_n473_1;
	wire [1:0] w_n481_0;
	wire [2:0] w_n483_0;
	wire [2:0] w_n483_1;
	wire [1:0] w_n483_2;
	wire [2:0] w_n485_0;
	wire [1:0] w_n485_1;
	wire [1:0] w_n493_0;
	wire [2:0] w_n494_0;
	wire [2:0] w_n494_1;
	wire [2:0] w_n496_0;
	wire [1:0] w_n496_1;
	wire [1:0] w_n504_0;
	wire [2:0] w_n507_0;
	wire [2:0] w_n507_1;
	wire [2:0] w_n509_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n518_0;
	wire [2:0] w_n518_1;
	wire [2:0] w_n520_0;
	wire [1:0] w_n528_0;
	wire [2:0] w_n530_0;
	wire [2:0] w_n530_1;
	wire [2:0] w_n532_0;
	wire [1:0] w_n532_1;
	wire [1:0] w_n540_0;
	wire [1:0] w_n543_0;
	wire [2:0] w_n551_0;
	wire [2:0] w_n556_0;
	wire [2:0] w_n556_1;
	wire [2:0] w_n556_2;
	wire [2:0] w_n556_3;
	wire [2:0] w_n556_4;
	wire [2:0] w_n556_5;
	wire [2:0] w_n556_6;
	wire [2:0] w_n556_7;
	wire [1:0] w_n556_8;
	wire [1:0] w_n557_0;
	wire [1:0] w_n559_0;
	wire [2:0] w_n560_0;
	wire [2:0] w_n561_0;
	wire [1:0] w_n561_1;
	wire [1:0] w_n562_0;
	wire [1:0] w_n564_0;
	wire [2:0] w_n565_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n567_0;
	wire [1:0] w_n569_0;
	wire [1:0] w_n571_0;
	wire [2:0] w_n572_0;
	wire [2:0] w_n573_0;
	wire [2:0] w_n574_0;
	wire [2:0] w_n578_0;
	wire [1:0] w_n578_1;
	wire [2:0] w_n579_0;
	wire [1:0] w_n579_1;
	wire [1:0] w_n581_0;
	wire [2:0] w_n586_0;
	wire [1:0] w_n586_1;
	wire [1:0] w_n587_0;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [2:0] w_n591_0;
	wire [1:0] w_n591_1;
	wire [2:0] w_n592_0;
	wire [2:0] w_n596_0;
	wire [1:0] w_n596_1;
	wire [2:0] w_n597_0;
	wire [2:0] w_n601_0;
	wire [1:0] w_n601_1;
	wire [2:0] w_n602_0;
	wire [1:0] w_n603_0;
	wire [2:0] w_n607_0;
	wire [1:0] w_n607_1;
	wire [2:0] w_n608_0;
	wire [2:0] w_n609_0;
	wire [2:0] w_n611_0;
	wire [2:0] w_n613_0;
	wire [2:0] w_n613_1;
	wire [2:0] w_n613_2;
	wire [2:0] w_n613_3;
	wire [2:0] w_n613_4;
	wire [2:0] w_n613_5;
	wire [2:0] w_n617_0;
	wire [1:0] w_n617_1;
	wire [2:0] w_n618_0;
	wire [2:0] w_n619_0;
	wire [2:0] w_n619_1;
	wire [2:0] w_n620_0;
	wire [1:0] w_n620_1;
	wire [1:0] w_n621_0;
	wire [1:0] w_n623_0;
	wire [2:0] w_n624_0;
	wire [1:0] w_n625_0;
	wire [2:0] w_n627_0;
	wire [1:0] w_n627_1;
	wire [2:0] w_n628_0;
	wire [1:0] w_n631_0;
	wire [1:0] w_n632_0;
	wire [2:0] w_n635_0;
	wire [1:0] w_n635_1;
	wire [2:0] w_n636_0;
	wire [2:0] w_n637_0;
	wire [1:0] w_n638_0;
	wire [2:0] w_n639_0;
	wire [1:0] w_n640_0;
	wire [2:0] w_n641_0;
	wire [2:0] w_n641_1;
	wire [2:0] w_n644_0;
	wire [2:0] w_n648_0;
	wire [1:0] w_n648_1;
	wire [1:0] w_n649_0;
	wire [1:0] w_n650_0;
	wire [2:0] w_n653_0;
	wire [2:0] w_n654_0;
	wire [2:0] w_n654_1;
	wire [2:0] w_n654_2;
	wire [2:0] w_n658_0;
	wire [1:0] w_n658_1;
	wire [1:0] w_n659_0;
	wire [2:0] w_n660_0;
	wire [1:0] w_n660_1;
	wire [1:0] w_n661_0;
	wire [1:0] w_n670_0;
	wire [1:0] w_n680_0;
	wire [2:0] w_n682_0;
	wire [1:0] w_n684_0;
	wire [1:0] w_n685_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n690_0;
	wire [1:0] w_n692_0;
	wire [2:0] w_n694_0;
	wire [2:0] w_n695_0;
	wire [2:0] w_n699_0;
	wire [1:0] w_n701_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n710_0;
	wire [1:0] w_n711_0;
	wire [2:0] w_n713_0;
	wire [2:0] w_n715_0;
	wire [1:0] w_n717_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n720_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n722_0;
	wire [2:0] w_n725_0;
	wire [1:0] w_n726_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n733_0;
	wire [2:0] w_n735_0;
	wire [2:0] w_n737_0;
	wire [1:0] w_n737_1;
	wire [1:0] w_n738_0;
	wire [2:0] w_n742_0;
	wire [1:0] w_n745_0;
	wire [2:0] w_n746_0;
	wire [1:0] w_n747_0;
	wire [2:0] w_n749_0;
	wire [2:0] w_n749_1;
	wire [2:0] w_n749_2;
	wire [2:0] w_n749_3;
	wire [2:0] w_n749_4;
	wire [2:0] w_n749_5;
	wire [2:0] w_n749_6;
	wire [2:0] w_n749_7;
	wire [2:0] w_n749_8;
	wire [2:0] w_n749_9;
	wire [2:0] w_n749_10;
	wire [2:0] w_n749_11;
	wire [2:0] w_n749_12;
	wire [1:0] w_n749_13;
	wire [2:0] w_n750_0;
	wire [2:0] w_n750_1;
	wire [2:0] w_n750_2;
	wire [2:0] w_n750_3;
	wire [2:0] w_n750_4;
	wire [2:0] w_n750_5;
	wire [2:0] w_n750_6;
	wire [2:0] w_n750_7;
	wire [2:0] w_n750_8;
	wire [2:0] w_n753_0;
	wire [1:0] w_n753_1;
	wire [1:0] w_n755_0;
	wire [2:0] w_n763_0;
	wire [1:0] w_n767_0;
	wire [1:0] w_n779_0;
	wire [2:0] w_n786_0;
	wire [2:0] w_n788_0;
	wire [2:0] w_n790_0;
	wire [2:0] w_n792_0;
	wire [2:0] w_n795_0;
	wire [1:0] w_n795_1;
	wire [2:0] w_n797_0;
	wire [2:0] w_n797_1;
	wire [2:0] w_n797_2;
	wire [2:0] w_n797_3;
	wire [2:0] w_n797_4;
	wire [2:0] w_n797_5;
	wire [2:0] w_n797_6;
	wire [2:0] w_n797_7;
	wire [2:0] w_n797_8;
	wire [1:0] w_n797_9;
	wire [2:0] w_n798_0;
	wire [1:0] w_n798_1;
	wire [2:0] w_n800_0;
	wire [2:0] w_n800_1;
	wire [2:0] w_n800_2;
	wire [2:0] w_n800_3;
	wire [1:0] w_n800_4;
	wire [2:0] w_n801_0;
	wire [1:0] w_n801_1;
	wire [2:0] w_n814_0;
	wire [2:0] w_n819_0;
	wire [1:0] w_n821_0;
	wire [1:0] w_n824_0;
	wire [1:0] w_n827_0;
	wire [1:0] w_n836_0;
	wire [1:0] w_n847_0;
	wire [2:0] w_n852_0;
	wire [2:0] w_n852_1;
	wire [2:0] w_n852_2;
	wire [2:0] w_n852_3;
	wire [2:0] w_n852_4;
	wire [2:0] w_n852_5;
	wire [2:0] w_n852_6;
	wire [2:0] w_n852_7;
	wire [2:0] w_n852_8;
	wire [1:0] w_n852_9;
	wire [2:0] w_n854_0;
	wire [2:0] w_n854_1;
	wire [2:0] w_n854_2;
	wire [2:0] w_n854_3;
	wire [1:0] w_n854_4;
	wire [2:0] w_n865_0;
	wire [1:0] w_n867_0;
	wire [1:0] w_n868_0;
	wire [1:0] w_n870_0;
	wire [1:0] w_n871_0;
	wire [1:0] w_n880_0;
	wire [1:0] w_n890_0;
	wire [1:0] w_n901_0;
	wire [2:0] w_n923_0;
	wire [1:0] w_n935_0;
	wire [2:0] w_n938_0;
	wire [2:0] w_n940_0;
	wire [1:0] w_n940_1;
	wire [1:0] w_n944_0;
	wire [1:0] w_n949_0;
	wire [1:0] w_n953_0;
	wire [2:0] w_n954_0;
	wire [1:0] w_n957_0;
	wire [1:0] w_n962_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n969_0;
	wire [2:0] w_n977_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n986_0;
	wire [1:0] w_n989_0;
	wire [2:0] w_n993_0;
	wire [2:0] w_n993_1;
	wire [2:0] w_n993_2;
	wire [2:0] w_n993_3;
	wire [2:0] w_n993_4;
	wire [2:0] w_n994_0;
	wire [2:0] w_n994_1;
	wire [2:0] w_n994_2;
	wire [2:0] w_n994_3;
	wire [1:0] w_n994_4;
	wire [2:0] w_n996_0;
	wire [2:0] w_n996_1;
	wire [2:0] w_n996_2;
	wire [2:0] w_n996_3;
	wire [1:0] w_n996_4;
	wire [2:0] w_n999_0;
	wire [2:0] w_n999_1;
	wire [2:0] w_n999_2;
	wire [2:0] w_n999_3;
	wire [2:0] w_n1007_0;
	wire [2:0] w_n1007_1;
	wire [2:0] w_n1007_2;
	wire [2:0] w_n1007_3;
	wire [2:0] w_n1008_0;
	wire [2:0] w_n1008_1;
	wire [2:0] w_n1008_2;
	wire [2:0] w_n1008_3;
	wire [2:0] w_n1008_4;
	wire [2:0] w_n1012_0;
	wire [2:0] w_n1012_1;
	wire [2:0] w_n1012_2;
	wire [2:0] w_n1012_3;
	wire [1:0] w_n1012_4;
	wire [2:0] w_n1014_0;
	wire [2:0] w_n1014_1;
	wire [2:0] w_n1014_2;
	wire [2:0] w_n1014_3;
	wire [1:0] w_n1014_4;
	wire [2:0] w_n1019_0;
	wire [1:0] w_n1019_1;
	wire [2:0] w_n1021_0;
	wire [1:0] w_n1021_1;
	wire [2:0] w_n1030_0;
	wire [1:0] w_n1030_1;
	wire [2:0] w_n1032_0;
	wire [1:0] w_n1032_1;
	wire [2:0] w_n1041_0;
	wire [1:0] w_n1041_1;
	wire [2:0] w_n1043_0;
	wire [1:0] w_n1043_1;
	wire [2:0] w_n1052_0;
	wire [1:0] w_n1052_1;
	wire [2:0] w_n1054_0;
	wire [1:0] w_n1054_1;
	wire [1:0] w_n1177_0;
	wire [1:0] w_n1179_0;
	wire [2:0] w_n1196_0;
	wire [2:0] w_n1196_1;
	wire [2:0] w_n1201_0;
	wire [2:0] w_n1205_0;
	wire [2:0] w_n1205_1;
	wire [2:0] w_n1213_0;
	wire [2:0] w_n1213_1;
	wire [2:0] w_n1236_0;
	wire [2:0] w_n1236_1;
	wire [2:0] w_n1251_0;
	wire [2:0] w_n1251_1;
	wire [2:0] w_n1279_0;
	wire [1:0] w_n1279_1;
	wire [2:0] w_n1297_0;
	wire [1:0] w_n1297_1;
	wire [2:0] w_n1299_0;
	wire [1:0] w_n1299_1;
	wire [2:0] w_n1410_0;
	wire [2:0] w_n1412_0;
	wire [1:0] w_n1416_0;
	wire [1:0] w_n1422_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1428_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1451_0;
	wire [1:0] w_n1503_0;
	wire [1:0] w_n1504_0;
	wire [1:0] w_n1592_0;
	wire [1:0] w_n1593_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1599_0;
	wire [1:0] w_n1603_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1609_0;
	wire [2:0] w_n1611_0;
	wire [1:0] w_n1613_0;
	wire [1:0] w_n1615_0;
	wire [1:0] w_n1618_0;
	wire [1:0] w_n1633_0;
	wire [1:0] w_n1637_0;
	wire [1:0] w_n1643_0;
	wire [1:0] w_n1652_0;
	wire [1:0] w_n1665_0;
	wire [2:0] w_n1674_0;
	wire [1:0] w_n1675_0;
	wire [2:0] w_n1679_0;
	wire [1:0] w_n1680_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1695_0;
	wire [1:0] w_n1698_0;
	wire w_dff_B_1GtAzzyc1_1;
	wire w_dff_B_uqSiIOCB0_0;
	wire w_dff_A_9AfsaUq23_0;
	wire w_dff_B_kF86fxm53_0;
	wire w_dff_A_s5V3QPdz0_2;
	wire w_dff_B_vir5UhkS1_1;
	wire w_dff_B_80zcCL4t4_0;
	wire w_dff_B_iajVVK8S0_1;
	wire w_dff_A_ycvSEpNX4_0;
	wire w_dff_A_ntJFtxVS6_0;
	wire w_dff_A_zMFKEvft7_1;
	wire w_dff_A_V5xbFpuQ9_1;
	wire w_dff_B_WhznrxG92_0;
	wire w_dff_B_uKAsZBfU9_1;
	wire w_dff_B_6oA78GKR0_1;
	wire w_dff_B_i1OZVmBg6_1;
	wire w_dff_A_wBPBDoQH6_0;
	wire w_dff_A_kkDkeOtI7_1;
	wire w_dff_A_uOTPqfW57_0;
	wire w_dff_A_tBwK81W68_1;
	wire w_dff_A_URWs1D7U2_1;
	wire w_dff_A_KKMLDXxK0_2;
	wire w_dff_A_U92YXMBk7_2;
	wire w_dff_B_4OnXHcKF9_1;
	wire w_dff_B_n6bJKEiU7_1;
	wire w_dff_B_dIhJzJxG9_2;
	wire w_dff_B_yoaHrVYM0_2;
	wire w_dff_B_MadxbEbI1_2;
	wire w_dff_B_SXfYI3Is7_1;
	wire w_dff_B_RtgVay2W2_1;
	wire w_dff_B_D8iqVJ2Q6_1;
	wire w_dff_B_YAfW2rFd1_1;
	wire w_dff_B_F2MQMNNB6_1;
	wire w_dff_B_2I0qUByN0_1;
	wire w_dff_B_xx9DLbcD3_1;
	wire w_dff_B_9G05yIxf1_1;
	wire w_dff_B_SxrYm4o84_1;
	wire w_dff_B_9kpzX39X0_1;
	wire w_dff_B_waXr1BrN4_3;
	wire w_dff_B_xQTz6HIA3_3;
	wire w_dff_B_wgFKBdCJ0_1;
	wire w_dff_B_QS51zgDE7_1;
	wire w_dff_B_RuIzu3Mf8_2;
	wire w_dff_A_FlMFMgdf0_0;
	wire w_dff_B_6ySXAuP76_0;
	wire w_dff_B_KXacjP3V7_0;
	wire w_dff_B_eJVw89vJ1_0;
	wire w_dff_B_WuXnYcSF4_0;
	wire w_dff_B_J8ZGGgmS1_0;
	wire w_dff_B_HCKpntyI3_0;
	wire w_dff_B_kc2nmk4k9_0;
	wire w_dff_B_mUrQO9oR4_0;
	wire w_dff_B_UXsIwkmT9_0;
	wire w_dff_B_oP1k9NoK2_0;
	wire w_dff_B_lR45vIp78_0;
	wire w_dff_A_Yx7UmKv56_1;
	wire w_dff_A_Crq9RCt17_1;
	wire w_dff_A_9l0I1sTh6_1;
	wire w_dff_A_8X4C068P3_1;
	wire w_dff_A_UvY8o15y2_1;
	wire w_dff_A_jVnbCgHv4_1;
	wire w_dff_A_McIVgIT22_1;
	wire w_dff_A_eIOOudUf5_1;
	wire w_dff_A_J7RHUXOW9_1;
	wire w_dff_B_1tmFAwfe5_0;
	wire w_dff_B_hjy2jNaQ9_0;
	wire w_dff_B_YfZSxOQ37_0;
	wire w_dff_B_YXU6TZLL5_0;
	wire w_dff_B_Hn7n8Wbo9_0;
	wire w_dff_B_RDjAUUkT5_0;
	wire w_dff_B_4CJRazDM9_0;
	wire w_dff_B_Dj4j1axa2_0;
	wire w_dff_B_aSz2eNAo4_0;
	wire w_dff_B_nUPCiQug9_2;
	wire w_dff_B_WXh6wnPF1_0;
	wire w_dff_B_1lmb96HG0_0;
	wire w_dff_A_IqOfsAYC0_1;
	wire w_dff_A_v4pg8jNg8_1;
	wire w_dff_A_gRUaYSXs5_1;
	wire w_dff_A_tJBUgvJr6_1;
	wire w_dff_A_0cK7920E0_1;
	wire w_dff_A_Kxyba8K44_1;
	wire w_dff_A_zDdPMkYz0_1;
	wire w_dff_A_AGhSKuX16_1;
	wire w_dff_A_qM0F7uvM9_1;
	wire w_dff_B_D04IyGQz9_1;
	wire w_dff_B_B3ZV9v6v5_1;
	wire w_dff_B_Tdu0oli02_1;
	wire w_dff_B_jFyidKdb4_0;
	wire w_dff_B_LAnULZFI4_1;
	wire w_dff_B_1KWLkI3m7_1;
	wire w_dff_B_TfsNJWrF9_1;
	wire w_dff_B_aWhiiJLm3_1;
	wire w_dff_B_zdnkO2lt6_1;
	wire w_dff_B_CnJApNPj8_1;
	wire w_dff_B_XzphINxT3_1;
	wire w_dff_B_8ekjMiix1_1;
	wire w_dff_B_GHsEjHdk7_1;
	wire w_dff_B_VZZxT2BA5_1;
	wire w_dff_B_Ykn1hPsE6_1;
	wire w_dff_B_rNIQAiam6_1;
	wire w_dff_B_qEiUIF176_1;
	wire w_dff_B_BTRFv6GO1_1;
	wire w_dff_B_eHVGDM220_1;
	wire w_dff_B_MRVjuMTV2_1;
	wire w_dff_B_mQ31TKdw6_1;
	wire w_dff_B_VZpgtv9Y5_1;
	wire w_dff_B_KpDqVaos2_1;
	wire w_dff_B_PTVEC55W7_1;
	wire w_dff_B_0I1c4ZuX8_0;
	wire w_dff_B_WqgVAaty1_0;
	wire w_dff_B_FCWVVXmB8_0;
	wire w_dff_B_fEDGH8EZ6_0;
	wire w_dff_B_yb2JosEl9_0;
	wire w_dff_B_It7SPVGc1_0;
	wire w_dff_B_EnJDi84e9_0;
	wire w_dff_B_d6okdsGf8_0;
	wire w_dff_B_u0iXXtuK6_0;
	wire w_dff_B_lSXyQPV36_0;
	wire w_dff_B_QqXudnfC0_0;
	wire w_dff_B_VQGxCGCs8_1;
	wire w_dff_B_Lw4WQfms1_2;
	wire w_dff_B_esaDwXgw5_2;
	wire w_dff_B_menrNAlj4_2;
	wire w_dff_B_Q7gad6Bs4_1;
	wire w_dff_B_1XnVT89E6_1;
	wire w_dff_B_q6VYX1OR3_1;
	wire w_dff_B_ZB6kUhF76_1;
	wire w_dff_B_jPQLoBK69_1;
	wire w_dff_B_ANVSRo600_1;
	wire w_dff_B_5MbQrCJc8_1;
	wire w_dff_B_jgWblR193_1;
	wire w_dff_B_2hXGawTK9_0;
	wire w_dff_B_ZrCBIzZC1_0;
	wire w_dff_B_8HXx2yJO4_0;
	wire w_dff_B_QMQVtFwl1_0;
	wire w_dff_B_CQjF9HTI5_1;
	wire w_dff_A_rkyTETuQ0_0;
	wire w_dff_B_qq3VnTOQ7_1;
	wire w_dff_B_tsE0BllG0_1;
	wire w_dff_B_ttqqGnET9_1;
	wire w_dff_B_uoBLLF5g3_0;
	wire w_dff_A_3L5GuXNH8_0;
	wire w_dff_A_XwW2Wqu36_0;
	wire w_dff_A_BQh33GQT4_0;
	wire w_dff_A_Ju5TH4xT9_0;
	wire w_dff_A_m1c6lnTn3_0;
	wire w_dff_A_m9RpRpGy0_0;
	wire w_dff_A_cTMAdxYM3_0;
	wire w_dff_A_SiWftj9M9_0;
	wire w_dff_B_ZNVvaAH95_1;
	wire w_dff_B_RntSM2gG0_1;
	wire w_dff_A_vkfbRAzT5_0;
	wire w_dff_B_hVUzqmlY6_0;
	wire w_dff_B_p9rBhHSU0_0;
	wire w_dff_B_FJ70SmwN3_0;
	wire w_dff_B_cbjbzLry7_0;
	wire w_dff_B_VMPa116o2_0;
	wire w_dff_B_M5gKOCH17_0;
	wire w_dff_B_xQ7fOP5t3_0;
	wire w_dff_B_WfFlJPVz0_0;
	wire w_dff_B_HbDo0Dos1_0;
	wire w_dff_B_J1xabP3Y8_0;
	wire w_dff_B_5Af90yN23_0;
	wire w_dff_B_vGfTQHdt9_0;
	wire w_dff_A_fczZGPYb8_0;
	wire w_dff_A_HexWks2A7_0;
	wire w_dff_A_OPOV61q12_0;
	wire w_dff_A_fdTn3Grr8_0;
	wire w_dff_A_FoZjywm18_0;
	wire w_dff_B_in6b97hS3_0;
	wire w_dff_B_P8pCc4jI2_0;
	wire w_dff_B_Y8jhCHRY6_0;
	wire w_dff_B_DX72x1Dn3_0;
	wire w_dff_B_SpDAdqbM9_0;
	wire w_dff_B_L8oDlve46_0;
	wire w_dff_B_8IYxjELw4_0;
	wire w_dff_B_3xix8IXc8_0;
	wire w_dff_B_QABUrzbd0_0;
	wire w_dff_B_y2vmSPBM0_0;
	wire w_dff_B_i0Opn9fq0_0;
	wire w_dff_B_zNb3Rqgq0_0;
	wire w_dff_B_34QnpZ2M2_1;
	wire w_dff_A_ztp9UyxC4_0;
	wire w_dff_A_h9GlRIyz6_0;
	wire w_dff_A_ZBcZCkIP4_0;
	wire w_dff_A_jHY2LGTj7_0;
	wire w_dff_A_lYA67wRe7_0;
	wire w_dff_A_uTOJRq2Q8_0;
	wire w_dff_A_nLz6SNRi6_0;
	wire w_dff_A_furoJDwM6_0;
	wire w_dff_A_OPFZvC1U0_0;
	wire w_dff_A_HOZ7xEdp7_0;
	wire w_dff_A_P2qDmiei6_0;
	wire w_dff_A_ocmlcEj69_0;
	wire w_dff_A_CeCPHWaB6_2;
	wire w_dff_A_vyNwRoTY3_2;
	wire w_dff_A_jdFdgVQU4_2;
	wire w_dff_A_b2ctLjbA2_2;
	wire w_dff_A_ZeZAIU0i2_2;
	wire w_dff_A_gJiX4mCC6_2;
	wire w_dff_A_jVv2e0RD5_2;
	wire w_dff_A_3S53QUgj4_2;
	wire w_dff_A_QnGWxoCM5_2;
	wire w_dff_A_hWCudCpn0_2;
	wire w_dff_A_6ocjygVS8_2;
	wire w_dff_A_LiETSce14_2;
	wire w_dff_A_66blaznK0_0;
	wire w_dff_A_4FlJvVeE8_0;
	wire w_dff_A_O4QnsGew3_0;
	wire w_dff_A_yaUNVupM8_0;
	wire w_dff_A_Qbry0MNV0_0;
	wire w_dff_A_TAeVVpbe5_0;
	wire w_dff_A_Ffu6A3878_0;
	wire w_dff_A_fTZisUBx1_0;
	wire w_dff_A_A35UpjuI3_0;
	wire w_dff_A_X0uJt3xl3_0;
	wire w_dff_A_7CmtykPV7_0;
	wire w_dff_A_GZg8pH6M2_2;
	wire w_dff_A_cFPji26A3_2;
	wire w_dff_A_PyqQVyQN7_2;
	wire w_dff_A_hl3ZBUnU1_2;
	wire w_dff_A_xETbLDDh2_2;
	wire w_dff_A_xlG8cCWC5_2;
	wire w_dff_A_wOpDK0AH4_2;
	wire w_dff_A_kzUGrd8N4_2;
	wire w_dff_A_3AHbYvb48_2;
	wire w_dff_A_VhiWsFc44_2;
	wire w_dff_A_TsJubJMW8_2;
	wire w_dff_A_VNLjHoOq3_2;
	wire w_dff_B_THCpPPMj9_0;
	wire w_dff_B_yuabpuIt1_0;
	wire w_dff_B_G1tRvPUO4_0;
	wire w_dff_B_ToE7XJ3Z9_0;
	wire w_dff_B_7mWaczjN3_0;
	wire w_dff_B_chDO7ZiU7_0;
	wire w_dff_B_0JLmbahI5_0;
	wire w_dff_B_sKXTQ5WP4_0;
	wire w_dff_B_1vxwo5Pz7_0;
	wire w_dff_B_PDKL7CSO4_0;
	wire w_dff_B_Id00WzHI6_0;
	wire w_dff_B_j3L33nz34_1;
	wire w_dff_B_JuabviMb4_1;
	wire w_dff_B_l7ktTNTI3_1;
	wire w_dff_A_BfyTGzgp9_1;
	wire w_dff_A_PjX0Nso77_1;
	wire w_dff_A_gZxUrYBL8_1;
	wire w_dff_A_0eh4I4zt9_1;
	wire w_dff_A_CBI4nD3J7_1;
	wire w_dff_A_aBuZFZTV1_1;
	wire w_dff_A_VdyuK2dy6_1;
	wire w_dff_A_Jns33q6O2_1;
	wire w_dff_A_mhuAIWXF2_1;
	wire w_dff_A_8yAFZfdD0_1;
	wire w_dff_A_tK8GKuzK9_1;
	wire w_dff_A_wOOebpOE6_1;
	wire w_dff_A_LEvTjwJc2_1;
	wire w_dff_A_XHwHNi6B0_1;
	wire w_dff_A_b8chBR272_1;
	wire w_dff_A_ZnkAIT4d6_1;
	wire w_dff_A_HLLOjFs03_1;
	wire w_dff_A_wSRdn8vo9_1;
	wire w_dff_A_LFa27Mez9_1;
	wire w_dff_B_AKAmyV3f7_0;
	wire w_dff_B_0uXH1LMm7_0;
	wire w_dff_B_iQ8kPDyP1_0;
	wire w_dff_B_L4P7t1YE8_0;
	wire w_dff_B_PbuM9bPv0_0;
	wire w_dff_B_sh9XEXea2_0;
	wire w_dff_B_q45UdfyB3_0;
	wire w_dff_B_B6Fs37IB9_0;
	wire w_dff_B_5lTzlez44_0;
	wire w_dff_B_2fehSlEE1_0;
	wire w_dff_B_VUAjNiRH7_1;
	wire w_dff_A_CzjPq7vf6_1;
	wire w_dff_A_1RpyB4Tt6_2;
	wire w_dff_A_Lb63Q02A7_2;
	wire w_dff_B_bkMId1lU2_1;
	wire w_dff_B_B1mY836K8_1;
	wire w_dff_B_tdonufCY7_1;
	wire w_dff_B_7VECIvT16_1;
	wire w_dff_B_g9YK2ECl3_1;
	wire w_dff_B_66krYkky0_1;
	wire w_dff_B_CL5gt7K56_1;
	wire w_dff_B_YBHM59qu6_1;
	wire w_dff_B_cCAeGkO51_1;
	wire w_dff_B_kyj8czcF3_1;
	wire w_dff_B_afQvGX8Q3_1;
	wire w_dff_B_e1pr8F9p2_1;
	wire w_dff_B_8cMfT4eI0_1;
	wire w_dff_A_jxmC1sKZ1_0;
	wire w_dff_A_830J17vn4_0;
	wire w_dff_A_WKrrakNZ0_0;
	wire w_dff_A_L9wK2kU57_0;
	wire w_dff_A_Hk6TBfrL2_0;
	wire w_dff_A_paDHeFq52_0;
	wire w_dff_A_7k4NVCHH8_0;
	wire w_dff_B_cUkosmGA6_1;
	wire w_dff_B_jLkq5yPJ4_1;
	wire w_dff_B_ukQxG9DW5_2;
	wire w_dff_B_0hJPXdL73_1;
	wire w_dff_B_0w1RXKKs7_1;
	wire w_dff_B_T1A0bSTN8_1;
	wire w_dff_B_AOw2XQ8g8_1;
	wire w_dff_B_iXIiX3Fa9_1;
	wire w_dff_B_iw4G9YfW7_1;
	wire w_dff_B_lXQHtbLP6_1;
	wire w_dff_B_0p0r8dTy5_1;
	wire w_dff_B_HcPIsBDU7_1;
	wire w_dff_B_5E47tHTh1_1;
	wire w_dff_B_Znv1cIZd9_1;
	wire w_dff_B_5roB9hPP7_1;
	wire w_dff_B_ZC7hCloA9_1;
	wire w_dff_A_apcP3Tg10_1;
	wire w_dff_A_2uzeD8po6_1;
	wire w_dff_A_sbXKNuc64_1;
	wire w_dff_A_PUv7y5HW9_1;
	wire w_dff_A_v1eeMBvn0_1;
	wire w_dff_A_dX0ckGmA7_1;
	wire w_dff_A_uxSTdeKI9_1;
	wire w_dff_A_iMM9QvWc9_1;
	wire w_dff_A_H163rTMi4_1;
	wire w_dff_A_5VXQVjaE2_1;
	wire w_dff_A_v4yyboEx4_1;
	wire w_dff_A_e0eMipcg4_1;
	wire w_dff_B_im5dFBrE5_2;
	wire w_dff_A_xfvpJ84k2_1;
	wire w_dff_A_uAZ1J8Ip2_1;
	wire w_dff_A_bHC6A4543_1;
	wire w_dff_A_wW8clFLT8_1;
	wire w_dff_A_QWxAQkT58_1;
	wire w_dff_A_Nzr8a2qN5_1;
	wire w_dff_A_LAKDsYHP8_1;
	wire w_dff_A_RdLmMYTu7_1;
	wire w_dff_A_UBexyctJ2_1;
	wire w_dff_A_n5yHaSaD6_1;
	wire w_dff_A_NpbvhCOn5_1;
	wire w_dff_A_a3kVmaUn1_1;
	wire w_dff_B_e1qVRQzZ8_1;
	wire w_dff_B_22V7Vy6N1_1;
	wire w_dff_B_IzrZfD424_1;
	wire w_dff_B_u978ur932_1;
	wire w_dff_B_d535fkPZ6_1;
	wire w_dff_B_BpjImiYi7_1;
	wire w_dff_B_OGrMSw1B1_1;
	wire w_dff_B_xFBCjbib8_1;
	wire w_dff_B_rURzYWoP2_1;
	wire w_dff_B_9czpcr7Z2_1;
	wire w_dff_B_S6YzImyS1_0;
	wire w_dff_B_a5h5n6Vd2_0;
	wire w_dff_B_x9LEJhtA0_1;
	wire w_dff_B_JvDrFjIk7_1;
	wire w_dff_A_gC9GFFaA2_0;
	wire w_dff_A_H7CjY4PM5_0;
	wire w_dff_A_zlhhaP7h6_0;
	wire w_dff_A_6cHSBxia6_0;
	wire w_dff_A_4caa1qTa1_0;
	wire w_dff_A_09yBD5uR1_0;
	wire w_dff_A_0WovloHB4_0;
	wire w_dff_A_DxwT3zI21_0;
	wire w_dff_A_qBX3YmmR7_0;
	wire w_dff_A_AyIjvPMV7_0;
	wire w_dff_A_iYgs8HQM4_2;
	wire w_dff_A_tLZDn3Wx7_2;
	wire w_dff_A_iAP1tBFO5_2;
	wire w_dff_A_49aC9TyN1_2;
	wire w_dff_A_swNPezMS9_2;
	wire w_dff_A_XYFnRj8u9_2;
	wire w_dff_A_xmCOz98r2_2;
	wire w_dff_A_wdETEzoP6_2;
	wire w_dff_A_Z3oUY14E9_2;
	wire w_dff_A_VfOToTWh7_2;
	wire w_dff_A_D7jBCDW84_2;
	wire w_dff_B_sd2ZVu9e6_2;
	wire w_dff_A_pB4g1s7L5_0;
	wire w_dff_A_onfVLaOH9_0;
	wire w_dff_A_Eiwuvmvc4_0;
	wire w_dff_A_bO9pOKDo4_0;
	wire w_dff_A_BIeNcFBX7_0;
	wire w_dff_A_CUoMUWNW1_0;
	wire w_dff_A_Ih9IteqR9_0;
	wire w_dff_A_X2Qapz4v4_0;
	wire w_dff_A_y3Wiv0ee2_0;
	wire w_dff_A_qpN8pgB39_2;
	wire w_dff_A_NnKahwor1_2;
	wire w_dff_A_0VzkEIZ50_2;
	wire w_dff_A_z6xmCqAD5_2;
	wire w_dff_A_Ja8TycIr8_2;
	wire w_dff_A_NeB8eP9O1_2;
	wire w_dff_A_os5MzVpX6_2;
	wire w_dff_A_9NmrFACZ2_2;
	wire w_dff_A_YIpNymjH5_2;
	wire w_dff_A_7KEDcc1i1_2;
	wire w_dff_A_xeiLnNYM0_2;
	wire w_dff_A_Ydf7G1MN5_2;
	wire w_dff_B_lwxmTE3c0_0;
	wire w_dff_B_m2KtoGiw9_0;
	wire w_dff_B_gDfP0Q7f7_0;
	wire w_dff_B_77xP8QcO7_0;
	wire w_dff_B_ADUqRKjA4_0;
	wire w_dff_B_dSkavKle9_0;
	wire w_dff_B_rTgsmJ0K2_0;
	wire w_dff_B_Eu1dSeSi8_0;
	wire w_dff_B_Tit3b0uv4_0;
	wire w_dff_B_rOZqIJ489_0;
	wire w_dff_A_nEW9LA4a0_1;
	wire w_dff_A_POkQJsV80_2;
	wire w_dff_B_tQUug1ty3_2;
	wire w_dff_B_GtnUh3fp5_1;
	wire w_dff_A_vRa1EFPx1_1;
	wire w_dff_A_7V3vbrfp1_1;
	wire w_dff_A_7cLK4wxq1_2;
	wire w_dff_A_d4p14SI83_2;
	wire w_dff_A_wQvkC4ud0_2;
	wire w_dff_B_aGUeRP3L2_0;
	wire w_dff_B_tuBnLgZo4_0;
	wire w_dff_B_we40hQC63_0;
	wire w_dff_B_P0WeECj87_0;
	wire w_dff_B_OQZLYPfR4_0;
	wire w_dff_B_0bSE72zb7_0;
	wire w_dff_B_Sszl1lTC4_0;
	wire w_dff_B_Mg1CfUbk9_0;
	wire w_dff_B_DyFG6Q476_0;
	wire w_dff_B_2IaB2hQo2_0;
	wire w_dff_B_Z7X0DKjP1_0;
	wire w_dff_B_L0foX1gb2_0;
	wire w_dff_B_Zg1UhuNn4_0;
	wire w_dff_B_AbvrSSu94_1;
	wire w_dff_B_dHD2NsdS6_1;
	wire w_dff_B_BhCxatF42_0;
	wire w_dff_B_sjVkna3y0_0;
	wire w_dff_B_faJmfSlV7_0;
	wire w_dff_B_JmoLRkOZ1_0;
	wire w_dff_B_ujjSmdMT7_0;
	wire w_dff_B_dUuYIzS16_0;
	wire w_dff_B_LJrJXStQ8_0;
	wire w_dff_B_t34VBvls2_0;
	wire w_dff_B_4wdvpaih2_0;
	wire w_dff_B_OKBEGDpY5_0;
	wire w_dff_B_lLyMDWw12_1;
	wire w_dff_A_MDICiLQy1_0;
	wire w_dff_A_zPHzPfKF5_0;
	wire w_dff_A_nw6sdVGv8_0;
	wire w_dff_A_ejV6WJxp7_1;
	wire w_dff_A_aRx0CpwE4_1;
	wire w_dff_A_J7kLXnJZ0_1;
	wire w_dff_A_iXFLeoAz1_1;
	wire w_dff_A_auO0Ihs89_1;
	wire w_dff_A_V9tpnX0W9_1;
	wire w_dff_A_NcOedwtw7_0;
	wire w_dff_A_HQ4yem6X0_0;
	wire w_dff_A_wPirhIZM5_0;
	wire w_dff_A_x6QrGI4k9_1;
	wire w_dff_A_dO9R75Pk8_1;
	wire w_dff_A_YReokgF71_1;
	wire w_dff_A_kaPTMUid6_1;
	wire w_dff_A_hU8ufdTl1_1;
	wire w_dff_B_iITIKDNb5_0;
	wire w_dff_B_XH9LBuJk1_0;
	wire w_dff_B_Tpy8NYjg2_0;
	wire w_dff_B_mQxmRu629_0;
	wire w_dff_B_qdwiHKA33_0;
	wire w_dff_B_IcOzOlfV6_0;
	wire w_dff_B_afsLMNDS3_0;
	wire w_dff_B_2fcslUvf1_0;
	wire w_dff_B_K1KunLx38_0;
	wire w_dff_B_LuGLwxXH5_0;
	wire w_dff_B_OL3NLugM8_0;
	wire w_dff_B_201JWcL95_1;
	wire w_dff_B_mWlLAJF08_1;
	wire w_dff_B_4Z6Nypry4_1;
	wire w_dff_A_mbCLFJ1C0_0;
	wire w_dff_A_APz6jERG5_2;
	wire w_dff_A_rl5AWjRP2_2;
	wire w_dff_A_3m7ZcVHv3_2;
	wire w_dff_B_bjQmrv3o6_0;
	wire w_dff_B_9PWobMtC4_0;
	wire w_dff_B_cMl2pxRp0_0;
	wire w_dff_B_jKGfgZXT8_0;
	wire w_dff_B_bi8BQgi44_0;
	wire w_dff_B_LZM14I1d0_0;
	wire w_dff_B_XrJbQawW4_0;
	wire w_dff_B_eP20ZFRJ2_0;
	wire w_dff_B_RF74xTuM8_0;
	wire w_dff_B_g3a2nV270_0;
	wire w_dff_B_mzqMQWYO7_0;
	wire w_dff_B_TRI8VtAe1_0;
	wire w_dff_B_rNLC0A6b9_1;
	wire w_dff_A_I7cFGMOk0_0;
	wire w_dff_A_5zgclu6e2_0;
	wire w_dff_A_WrwQKUNH7_1;
	wire w_dff_B_QNE4u8UD2_1;
	wire w_dff_B_2OibqZSg5_1;
	wire w_dff_B_cmJ4Sanv8_1;
	wire w_dff_B_GZNcX2g00_1;
	wire w_dff_B_ZcOcE4TC4_1;
	wire w_dff_B_DqEEM4R79_1;
	wire w_dff_B_EmpDHZlQ2_1;
	wire w_dff_B_OQ8RAhaU2_1;
	wire w_dff_B_QW1gJaCr4_1;
	wire w_dff_B_cZtruJZp8_1;
	wire w_dff_B_9dKtiNDO5_1;
	wire w_dff_B_O8UO2SZW0_1;
	wire w_dff_B_fOThIB7Q0_1;
	wire w_dff_B_vdVXqaMK2_1;
	wire w_dff_B_hxRqJRzm1_1;
	wire w_dff_B_kaGws2ym7_1;
	wire w_dff_B_6EJG7CkC3_1;
	wire w_dff_B_lvafxM903_1;
	wire w_dff_B_aJ4zOciI9_1;
	wire w_dff_B_8CPFJZ6j1_1;
	wire w_dff_B_0SJciPGz8_1;
	wire w_dff_B_IcIzwzrP5_1;
	wire w_dff_B_aUAbdcNR7_1;
	wire w_dff_B_6ZKop9ww7_1;
	wire w_dff_B_039QYSRB1_1;
	wire w_dff_B_beWqPsAs9_0;
	wire w_dff_B_SCNZweY59_1;
	wire w_dff_B_VnrBFmea0_1;
	wire w_dff_B_WwWbbkQL5_1;
	wire w_dff_B_6tLdqHvS2_1;
	wire w_dff_B_y8BTqAfv6_1;
	wire w_dff_B_9RWlcmWY9_1;
	wire w_dff_B_DoV4iL8k7_0;
	wire w_dff_B_48oF9AZD9_0;
	wire w_dff_B_6v9iZpdS7_0;
	wire w_dff_B_YOF0tylv7_0;
	wire w_dff_B_TIa6Cguv5_0;
	wire w_dff_B_sL7vJs5x6_0;
	wire w_dff_A_s0mWYLZx6_1;
	wire w_dff_B_F9EoP2rl4_1;
	wire w_dff_B_MTFsqagk5_1;
	wire w_dff_B_z3Nd8qxk9_1;
	wire w_dff_B_LjCjvAaW5_1;
	wire w_dff_B_sedO53ka2_1;
	wire w_dff_B_c2WqjHWj4_1;
	wire w_dff_B_JwiEoX8s2_1;
	wire w_dff_B_Tala5Q3g3_1;
	wire w_dff_B_QZpvcZaB4_1;
	wire w_dff_B_TyevNExH3_1;
	wire w_dff_B_laLYCMTy3_1;
	wire w_dff_B_NvWPEA940_1;
	wire w_dff_B_GfAwnbcw4_1;
	wire w_dff_B_ZsiKmdKd1_1;
	wire w_dff_B_GtDlaz1j4_0;
	wire w_dff_B_0z7eOQJI9_0;
	wire w_dff_B_dyc5tWD73_0;
	wire w_dff_B_FU3Szuor4_0;
	wire w_dff_B_sIoewJFH8_0;
	wire w_dff_B_TK1m8UMz9_0;
	wire w_dff_B_myhdTuYj6_0;
	wire w_dff_B_1JyXEtsm3_1;
	wire w_dff_B_SauEUFGf6_1;
	wire w_dff_B_c5kHQJeJ9_1;
	wire w_dff_B_fJjEArNj5_2;
	wire w_dff_B_FU2GyNtp4_2;
	wire w_dff_B_P7lro8k06_2;
	wire w_dff_B_kRSMxXCm1_0;
	wire w_dff_B_M1dIrjKe6_0;
	wire w_dff_B_wrTZK3aY2_0;
	wire w_dff_B_X8HOIuIg7_0;
	wire w_dff_B_cOEWvLM80_0;
	wire w_dff_B_C2RHxMHD5_0;
	wire w_dff_B_nYyjJrNm4_0;
	wire w_dff_B_uERNU9TH2_0;
	wire w_dff_B_7VhNgJT62_0;
	wire w_dff_B_Nxu03oUQ0_0;
	wire w_dff_B_Qku3HVSq6_2;
	wire w_dff_B_F43lJ4044_2;
	wire w_dff_B_fBz5XXFX2_2;
	wire w_dff_B_6d5lY3U59_1;
	wire w_dff_B_aJo1nRbC1_1;
	wire w_dff_B_bgvZjZNJ3_1;
	wire w_dff_B_73awkLfH9_1;
	wire w_dff_B_aqObUz5T9_1;
	wire w_dff_B_MKcm9QhE1_0;
	wire w_dff_B_uYkATdKd6_0;
	wire w_dff_B_vNOiyNA02_0;
	wire w_dff_B_D2gjCNcq2_0;
	wire w_dff_B_aMvWkg9f4_1;
	wire w_dff_A_dBRegjB43_0;
	wire w_dff_A_F6Ryisq53_0;
	wire w_dff_B_zW1FaUDe4_1;
	wire w_dff_B_uc5mNuws3_1;
	wire w_dff_A_mnVniqVR9_1;
	wire w_dff_A_U9FwaGHB7_1;
	wire w_dff_A_hp6tJ3RD6_1;
	wire w_dff_A_ARkK3bjp4_1;
	wire w_dff_B_YpfmQm0m0_1;
	wire w_dff_B_lNitwqbK2_1;
	wire w_dff_B_qdjYAWkp4_1;
	wire w_dff_B_WKaXesSI6_1;
	wire w_dff_B_KfCYvZFK0_0;
	wire w_dff_B_fyau8eTK4_0;
	wire w_dff_B_bccpTALs6_0;
	wire w_dff_B_xvh3OphK0_0;
	wire w_dff_B_nek1dyeV9_1;
	wire w_dff_B_BWMxTbrC1_0;
	wire w_dff_B_PKKUPnJQ6_0;
	wire w_dff_B_bvUdY8NE0_0;
	wire w_dff_A_syCrgftP0_0;
	wire w_dff_A_819bBhEI4_0;
	wire w_dff_A_wdVqBrym4_0;
	wire w_dff_A_hurffN830_0;
	wire w_dff_A_5qpZxzkn1_0;
	wire w_dff_A_GAPszGMA6_0;
	wire w_dff_B_V4cX5wPa7_1;
	wire w_dff_B_EDicO3ac1_1;
	wire w_dff_A_qPIwHP0t4_1;
	wire w_dff_A_nyqAEYAd7_1;
	wire w_dff_A_ZkMZMwwK5_1;
	wire w_dff_A_w6xNupWn1_2;
	wire w_dff_A_LHfbv8a61_2;
	wire w_dff_A_nslVg6tw9_0;
	wire w_dff_A_qWjcXWzl4_1;
	wire w_dff_B_84nPq5fe2_0;
	wire w_dff_B_BSRtKwJs3_0;
	wire w_dff_B_8tJOCkGq1_0;
	wire w_dff_B_CpK3WHEH9_0;
	wire w_dff_B_WOn2ylnQ3_0;
	wire w_dff_B_HL7G0cZb0_0;
	wire w_dff_B_iGPXOkeR0_0;
	wire w_dff_B_yWfnQGqC1_0;
	wire w_dff_B_GN5pjDSK5_0;
	wire w_dff_B_tb7gYmZ10_0;
	wire w_dff_B_oc0B1lNu8_0;
	wire w_dff_B_QRfzaI208_2;
	wire w_dff_B_EkoNtpq80_2;
	wire w_dff_B_BpTF5GQy4_2;
	wire w_dff_B_aSaFLFPL9_1;
	wire w_dff_B_Fv6no2Ey8_1;
	wire w_dff_B_knRvT7tP7_1;
	wire w_dff_B_9TVfkL8R6_1;
	wire w_dff_B_F1guUStm2_1;
	wire w_dff_B_NKLB37uY2_1;
	wire w_dff_B_MZgEDszm3_1;
	wire w_dff_B_3QS9wXdt8_1;
	wire w_dff_B_qUJx8LBb8_0;
	wire w_dff_B_bsfaDhKk9_0;
	wire w_dff_B_xxqTxMre1_0;
	wire w_dff_B_bTvv8oSU1_0;
	wire w_dff_B_dLxIWmEe6_0;
	wire w_dff_B_Tgn2H91z5_1;
	wire w_dff_B_z1Eielot2_0;
	wire w_dff_B_vFwuNlNw2_1;
	wire w_dff_B_Hp7PbKvj2_1;
	wire w_dff_B_rNs4GD8K8_1;
	wire w_dff_B_NLM2AQr62_1;
	wire w_dff_B_trAlkVrw5_1;
	wire w_dff_B_zzFaTFQg8_1;
	wire w_dff_B_lghMQ7Yz0_1;
	wire w_dff_B_7n3YPTJS0_1;
	wire w_dff_A_30dIqxAf0_0;
	wire w_dff_A_qOxMpK4H6_0;
	wire w_dff_A_ae4ddyxY3_0;
	wire w_dff_A_ww4RAWBC9_0;
	wire w_dff_B_SWNB9SoI5_1;
	wire w_dff_B_8gFBKhv31_1;
	wire w_dff_B_qVeNaaDJ7_1;
	wire w_dff_B_026NcNg70_0;
	wire w_dff_B_pFSwHHtb2_0;
	wire w_dff_B_jkWuy1ni8_0;
	wire w_dff_B_JXbAYvgO8_0;
	wire w_dff_B_jMxPL8SS5_0;
	wire w_dff_B_LCkv9DTj6_0;
	wire w_dff_B_qGXRgWgy9_0;
	wire w_dff_B_ZUjZvtYv0_0;
	wire w_dff_B_tHPhL2Gm9_0;
	wire w_dff_B_2zxle7Eu4_0;
	wire w_dff_B_coJcKL1t1_0;
	wire w_dff_B_8jjA69mY4_0;
	wire w_dff_B_CUdKH9X76_2;
	wire w_dff_B_r0QTEMSG2_2;
	wire w_dff_B_Vtj1ABIZ9_2;
	wire w_dff_B_wnl81Iyh3_1;
	wire w_dff_B_9whXdIIs9_1;
	wire w_dff_B_Q1rEGta80_1;
	wire w_dff_B_eOBOxAxZ8_1;
	wire w_dff_B_uM8Jl3zU7_1;
	wire w_dff_B_sSNvPANC4_1;
	wire w_dff_B_ODrs3Hv98_1;
	wire w_dff_B_8hVuXK618_0;
	wire w_dff_B_i7CxdktL4_0;
	wire w_dff_B_q9OM7uZS4_0;
	wire w_dff_B_dqrFfrfa0_0;
	wire w_dff_B_5huyXDVK3_0;
	wire w_dff_B_Gip1KnOr8_0;
	wire w_dff_B_ns3mmr1l6_1;
	wire w_dff_A_AuhDZwQi4_2;
	wire w_dff_A_HB1k4VTa7_2;
	wire w_dff_A_sVMre9Ik6_2;
	wire w_dff_A_MV8w9BWA8_0;
	wire w_dff_A_qQK4ptO99_0;
	wire w_dff_A_9GCQO9zD4_0;
	wire w_dff_A_9gC8U8aS1_1;
	wire w_dff_A_clEifxhA9_2;
	wire w_dff_A_VBoCBJqN8_2;
	wire w_dff_B_lXrQxOTa6_1;
	wire w_dff_B_bMPd2nWQ2_1;
	wire w_dff_A_CJHvcAcc3_0;
	wire w_dff_A_BaOSPFsm5_0;
	wire w_dff_A_rDg5QNjv5_1;
	wire w_dff_B_SyrpvCGw4_1;
	wire w_dff_B_cF1kL6Ir0_1;
	wire w_dff_B_n5R4Zt7E6_1;
	wire w_dff_B_6QAueIRe5_1;
	wire w_dff_B_6AfSqez20_1;
	wire w_dff_B_ETrn17uu3_1;
	wire w_dff_B_aHYp6zQn1_0;
	wire w_dff_B_7XkRhDja7_0;
	wire w_dff_B_p9Yvvedh9_0;
	wire w_dff_B_McGf1tEs0_0;
	wire w_dff_B_6LzYTQeG1_0;
	wire w_dff_B_6H8o4d9y1_0;
	wire w_dff_B_de19BWZc6_1;
	wire w_dff_A_WqWAB9at4_0;
	wire w_dff_A_DwUkGJs80_0;
	wire w_dff_A_L8dLDJ6w5_0;
	wire w_dff_A_5bRvF0Nh4_0;
	wire w_dff_A_FIlawX3a4_1;
	wire w_dff_A_aQ50xBuz5_1;
	wire w_dff_A_3bDdvGbk4_2;
	wire w_dff_A_2WmamI4n2_2;
	wire w_dff_A_beQmwRy67_2;
	wire w_dff_A_ks8FVTFN3_2;
	wire w_dff_A_4WBJbeab2_2;
	wire w_dff_B_t1FXFAaZ7_3;
	wire w_dff_A_DHNOFN4p6_0;
	wire w_dff_A_WGV5FVai3_0;
	wire w_dff_A_AdnlTC4Y5_0;
	wire w_dff_A_smjPFL1o7_0;
	wire w_dff_A_EWBqzcHE4_2;
	wire w_dff_A_Jyys0oDK4_2;
	wire w_dff_A_rbirpuik2_2;
	wire w_dff_B_bLfx55vc8_1;
	wire w_dff_B_9OEG3cWT9_1;
	wire w_dff_B_tO0mzwg96_1;
	wire w_dff_B_lhRGlw9K9_1;
	wire w_dff_B_FQQWkwii8_1;
	wire w_dff_B_wn5iN9zw9_1;
	wire w_dff_B_SjU1yt2V7_1;
	wire w_dff_B_unZKnTdD0_1;
	wire w_dff_B_70wxUfHc4_1;
	wire w_dff_B_B7UMTwev4_1;
	wire w_dff_B_FlQNaKcG7_1;
	wire w_dff_B_eQteUKjZ2_1;
	wire w_dff_B_XLSHq1Th9_1;
	wire w_dff_B_2u0ShZUG1_1;
	wire w_dff_B_NGnx5LnA9_1;
	wire w_dff_B_198XHMzy8_1;
	wire w_dff_B_PSrErrhy7_1;
	wire w_dff_B_qynal3SP1_1;
	wire w_dff_B_QekT2fM28_1;
	wire w_dff_B_Xt9Y9EYs6_1;
	wire w_dff_B_QyHALjbl8_0;
	wire w_dff_B_8p7F8Wpz3_0;
	wire w_dff_B_D4sCE0H09_0;
	wire w_dff_B_KmYStiCn2_0;
	wire w_dff_B_vhdNbXMJ9_0;
	wire w_dff_B_BqG7FfWw6_0;
	wire w_dff_B_owT8PVMb3_0;
	wire w_dff_B_VTJlbBN22_0;
	wire w_dff_B_Vl5L1zmB2_0;
	wire w_dff_B_7lHRc8zN2_0;
	wire w_dff_B_KnwnaKGM1_0;
	wire w_dff_B_ITFQcYXI8_1;
	wire w_dff_B_0qpq5DAt7_1;
	wire w_dff_B_KgvbjEim3_1;
	wire w_dff_B_fPVcmVYO6_1;
	wire w_dff_B_ajBqM8tc6_1;
	wire w_dff_B_CQpxvma20_1;
	wire w_dff_B_P0bI9bgD6_1;
	wire w_dff_A_szaHesc36_0;
	wire w_dff_A_vXyBZDLX0_0;
	wire w_dff_A_WfZzG6FB3_0;
	wire w_dff_A_bln2jIrX8_0;
	wire w_dff_A_SVYpcLbw9_0;
	wire w_dff_A_C1IDkzsS0_0;
	wire w_dff_A_i4bemp5d7_0;
	wire w_dff_B_o9gmxaQ76_2;
	wire w_dff_B_UCILfZAn5_2;
	wire w_dff_B_RSIx4bsn9_2;
	wire w_dff_B_cMRgaMlm1_2;
	wire w_dff_A_pZ8QkzW89_1;
	wire w_dff_A_UrsF4Apy8_2;
	wire w_dff_A_c54t0iqu8_2;
	wire w_dff_A_wwcE1kRT2_2;
	wire w_dff_A_3iQpeY224_0;
	wire w_dff_A_o5mE3gb71_0;
	wire w_dff_A_VN0ZYhaT8_0;
	wire w_dff_A_quFaGz0f9_0;
	wire w_dff_A_lDlSrtFN3_0;
	wire w_dff_A_Gplb7tj13_0;
	wire w_dff_A_euOf8vAs0_0;
	wire w_dff_B_EdChOtUI6_1;
	wire w_dff_B_IgrB5vSH2_1;
	wire w_dff_B_K6VgBYY54_1;
	wire w_dff_B_oRispRRq4_1;
	wire w_dff_B_KZEWDumJ5_0;
	wire w_dff_B_3nXIKtGi0_0;
	wire w_dff_B_LDROBFzc7_0;
	wire w_dff_B_kmLJ1tZm4_0;
	wire w_dff_B_CqnFOVbl3_0;
	wire w_dff_A_voFT6FAY7_0;
	wire w_dff_A_5dlESbO32_0;
	wire w_dff_B_8m802Xw05_0;
	wire w_dff_B_HrWB5H7K4_1;
	wire w_dff_B_ieA4H7A44_1;
	wire w_dff_B_oLh5Lp4R4_1;
	wire w_dff_B_uBK8rf9p3_1;
	wire w_dff_B_6hPxrTld8_1;
	wire w_dff_B_ZQaKcf964_0;
	wire w_dff_B_ubAaVd4l6_1;
	wire w_dff_B_jCDCYhlj0_0;
	wire w_dff_B_5GvTtmRH5_0;
	wire w_dff_B_i8kUr1e56_1;
	wire w_dff_B_lprhXOTy9_1;
	wire w_dff_B_nmbHJMig4_1;
	wire w_dff_B_YidhlQNS8_0;
	wire w_dff_B_AjBRgu6e9_0;
	wire w_dff_B_yQZ9oo2Z6_0;
	wire w_dff_B_UkrEuE9s7_0;
	wire w_dff_B_VDU12DIm5_1;
	wire w_dff_A_cIv5IQkG3_0;
	wire w_dff_A_xRo5UZdV2_0;
	wire w_dff_A_BsGQ8ETt0_0;
	wire w_dff_A_G9Pwthw85_0;
	wire w_dff_B_M65zM5Hf2_1;
	wire w_dff_B_zeRRCORY7_1;
	wire w_dff_B_pZDJJ7u89_1;
	wire w_dff_B_SayaEkvV4_1;
	wire w_dff_B_gagvMuUz4_1;
	wire w_dff_B_miCOhRWA2_1;
	wire w_dff_B_8zVrpvmF9_1;
	wire w_dff_B_7Aumt0np9_1;
	wire w_dff_B_R3GMazw41_1;
	wire w_dff_B_CcFBvzJs4_1;
	wire w_dff_B_6rxe9iZv5_1;
	wire w_dff_B_6ai4waMO7_1;
	wire w_dff_B_jyX6kh7H4_1;
	wire w_dff_B_HpivnRXk6_1;
	wire w_dff_B_kjUlIwkl0_1;
	wire w_dff_B_1r5N1f4X6_1;
	wire w_dff_B_7Gg8tduh0_1;
	wire w_dff_B_y4GRpozF4_1;
	wire w_dff_B_UpTPaB8V4_1;
	wire w_dff_B_l5liVw6T3_0;
	wire w_dff_B_x1Sxh1Kz0_1;
	wire w_dff_B_oIzlAM068_1;
	wire w_dff_A_4RjYFG4K9_2;
	wire w_dff_A_ZLMebdVg6_2;
	wire w_dff_A_rCyVFMDg6_2;
	wire w_dff_A_wHMLXklS3_2;
	wire w_dff_A_DsOyQXxt6_2;
	wire w_dff_A_ob3Uspce6_2;
	wire w_dff_A_X1HmajJw6_2;
	wire w_dff_A_NvnRKjZL9_2;
	wire w_dff_A_9x3Yo8EN9_2;
	wire w_dff_A_8JGtiVNQ6_2;
	wire w_dff_A_LMOioVDJ3_2;
	wire w_dff_A_eJYbyVf70_2;
	wire w_dff_A_GEgtIHgQ6_2;
	wire w_dff_A_CAXsjpkX6_2;
	wire w_dff_A_PNDRObHB4_2;
	wire w_dff_A_Z519ggSy1_2;
	wire w_dff_A_d22uQCar0_2;
	wire w_dff_A_JDItCrtt2_2;
	wire w_dff_A_YrEGUGTu5_2;
	wire w_dff_B_HSLOQpXc2_0;
	wire w_dff_B_lgbymOOJ9_0;
	wire w_dff_B_N9vB34J35_0;
	wire w_dff_B_XSoYDXjI0_0;
	wire w_dff_B_K9jChpCQ0_0;
	wire w_dff_B_sjwgHYEH6_0;
	wire w_dff_B_pUomxi3t2_0;
	wire w_dff_B_3fI1vQaf1_0;
	wire w_dff_B_AL122XYB9_0;
	wire w_dff_B_LWtPXt185_0;
	wire w_dff_B_GLeeVZ5K7_0;
	wire w_dff_B_QZjZ94RC1_0;
	wire w_dff_B_ciHm6jhR3_0;
	wire w_dff_B_8CktlJcR5_0;
	wire w_dff_B_cP2vFUK47_0;
	wire w_dff_B_Ys6cIc8n8_2;
	wire w_dff_B_X6mec9Ar6_1;
	wire w_dff_B_tII93kEQ5_1;
	wire w_dff_B_beRkpLEE2_1;
	wire w_dff_A_EIhygtvp0_0;
	wire w_dff_A_0xH5TIIg0_0;
	wire w_dff_A_mfQpytnV1_0;
	wire w_dff_A_WKC49Meu0_0;
	wire w_dff_A_1gxq7JWy7_0;
	wire w_dff_A_bevwvuwM9_0;
	wire w_dff_A_ZxnVxvec0_0;
	wire w_dff_A_fPSPLAGd1_0;
	wire w_dff_A_d0MrzTYe8_0;
	wire w_dff_A_ShtoPeI53_0;
	wire w_dff_A_wRUR3CdM8_0;
	wire w_dff_A_Z5xKLcse1_0;
	wire w_dff_A_7paWf7me8_0;
	wire w_dff_A_i7vIy5nd8_0;
	wire w_dff_A_l07kGdf07_2;
	wire w_dff_A_QALrA6Ug2_2;
	wire w_dff_A_3ov9t8sz4_2;
	wire w_dff_A_Cr28jNBd5_2;
	wire w_dff_A_tShaQ5nr3_2;
	wire w_dff_A_OAWtnM404_2;
	wire w_dff_A_qdqH9rKd4_2;
	wire w_dff_A_blZP9Hfz6_2;
	wire w_dff_A_w1EBiFrA3_2;
	wire w_dff_A_8X7AsI6h6_0;
	wire w_dff_A_ZVZPeOv60_0;
	wire w_dff_A_Kz9vVoEa0_0;
	wire w_dff_A_dpSplsPl5_0;
	wire w_dff_A_GgguOPOl9_0;
	wire w_dff_A_WLwsBMxg3_0;
	wire w_dff_A_vBD5oPDR3_0;
	wire w_dff_A_Jf6CIFIy8_0;
	wire w_dff_A_ggBehG243_0;
	wire w_dff_A_AMZqHj9V9_0;
	wire w_dff_A_ogHOGOfJ8_0;
	wire w_dff_A_qH8pCZaJ4_0;
	wire w_dff_A_wmvximqy1_0;
	wire w_dff_A_LeDPvtRG1_2;
	wire w_dff_A_Uyg8AFmx8_2;
	wire w_dff_A_Fj7z8uzD1_2;
	wire w_dff_A_Vd5jpfGX2_2;
	wire w_dff_A_N8utaI5B1_2;
	wire w_dff_A_KZnepCYa3_2;
	wire w_dff_A_T1rtKHIl4_2;
	wire w_dff_A_6NJ7VYnd6_2;
	wire w_dff_A_R7j4hwe17_2;
	wire w_dff_A_aO7SEFju5_2;
	wire w_dff_B_4bNGrXUQ9_0;
	wire w_dff_B_07wly5Ol4_0;
	wire w_dff_B_56WsX3sS6_0;
	wire w_dff_B_dbuNXJN80_0;
	wire w_dff_B_DuhFN4vE0_0;
	wire w_dff_B_HlmbQFyF2_0;
	wire w_dff_B_9IIJg3y20_0;
	wire w_dff_B_P0P025ms5_0;
	wire w_dff_B_MqEipejA5_0;
	wire w_dff_B_Fp31TEwl9_0;
	wire w_dff_B_7nnYvt1J9_0;
	wire w_dff_B_qAfv0Rnk6_0;
	wire w_dff_B_pguaHEhJ4_0;
	wire w_dff_B_CyOCDMME2_0;
	wire w_dff_B_fbzNMePi9_0;
	wire w_dff_B_ozTQxUHt5_1;
	wire w_dff_B_M8TbZGfO8_1;
	wire w_dff_B_VvxiDDw61_1;
	wire w_dff_A_61hyrzFl7_1;
	wire w_dff_A_YosYbhOc1_1;
	wire w_dff_A_fifs4hFG3_1;
	wire w_dff_A_XebadTqn6_1;
	wire w_dff_A_m5QyaTK99_1;
	wire w_dff_A_awIwdeP06_1;
	wire w_dff_A_I3aCi0CK7_1;
	wire w_dff_A_mkestAyB1_1;
	wire w_dff_A_FnL4gZXA3_1;
	wire w_dff_A_5MYECC5F6_1;
	wire w_dff_A_QKLOlKfY0_1;
	wire w_dff_A_QaMlli2f3_1;
	wire w_dff_A_gRAkpv5i7_1;
	wire w_dff_A_83cHrO3Z0_1;
	wire w_dff_A_tUFwpcmo8_1;
	wire w_dff_A_MFEXzr504_1;
	wire w_dff_A_6RRPLTSU8_1;
	wire w_dff_A_HLeZWtBx3_1;
	wire w_dff_A_J21HaI1L7_1;
	wire w_dff_A_KzwLaXnn5_1;
	wire w_dff_A_raXqmRL08_1;
	wire w_dff_A_2LiweVeY7_1;
	wire w_dff_A_lwEotw011_1;
	wire w_dff_A_AH3fLX0w5_1;
	wire w_dff_A_ETld6wek7_1;
	wire w_dff_A_sjYm9l1t9_1;
	wire w_dff_A_aBzkJTVZ8_1;
	wire w_dff_B_RVRPJh1j7_0;
	wire w_dff_B_rqBZ1JQI3_0;
	wire w_dff_B_LwpIlTuo8_0;
	wire w_dff_B_5HhsiZ1R5_0;
	wire w_dff_B_aRBGPgfP2_0;
	wire w_dff_B_zYZ7TxIn0_0;
	wire w_dff_B_LskRZRaP1_0;
	wire w_dff_B_dqXOf1pv5_0;
	wire w_dff_B_0Ej2agMG2_0;
	wire w_dff_B_2nWOtnAg5_0;
	wire w_dff_B_JodKFaiP1_0;
	wire w_dff_B_iR0DYSKz7_0;
	wire w_dff_B_8JZi2Twq7_0;
	wire w_dff_B_3RpqSXkc4_0;
	wire w_dff_B_JomtzdNK1_1;
	wire w_dff_B_CkXm9KeI4_1;
	wire w_dff_B_CFSdghtJ8_1;
	wire w_dff_A_VSsgog7F1_1;
	wire w_dff_A_PnFovOBO9_2;
	wire w_dff_B_2daa77Bo1_0;
	wire w_dff_B_y3IsT7Ic0_0;
	wire w_dff_B_mxCDFJq14_0;
	wire w_dff_B_iWbjM1nD3_0;
	wire w_dff_B_A3D80apv4_0;
	wire w_dff_B_vGlipJHY2_0;
	wire w_dff_B_3fVfgQg17_0;
	wire w_dff_B_hUH6JMAN9_0;
	wire w_dff_B_UkIEKpXw8_0;
	wire w_dff_B_aZyKo8Bx4_0;
	wire w_dff_B_hju0W5HN8_0;
	wire w_dff_B_51FasEN76_0;
	wire w_dff_B_kZpqylnS4_0;
	wire w_dff_B_dxwp7vRm7_0;
	wire w_dff_B_xeFe8tDL3_0;
	wire w_dff_B_R6k2vql07_1;
	wire w_dff_B_KgK6Eytl0_1;
	wire w_dff_B_DCa37vzH1_1;
	wire w_dff_A_3dhf2zH69_0;
	wire w_dff_A_PKD4sYhK0_0;
	wire w_dff_A_X5907bwN2_0;
	wire w_dff_A_ftdpoaOF7_0;
	wire w_dff_A_gfXIgObn6_0;
	wire w_dff_A_aGWmHD8e7_0;
	wire w_dff_A_zRzgAmkL3_0;
	wire w_dff_A_duxIveYA0_0;
	wire w_dff_A_ulhTxpCP3_0;
	wire w_dff_A_O0yG5oUA9_0;
	wire w_dff_A_mEXwCAXT9_0;
	wire w_dff_A_ErQlNHns9_0;
	wire w_dff_A_z9bYcK5w1_0;
	wire w_dff_A_drLVlnn43_0;
	wire w_dff_A_le1zyTkC4_2;
	wire w_dff_A_PqxpfCk62_2;
	wire w_dff_A_aTmrLBR34_2;
	wire w_dff_A_Pq8d67pW6_2;
	wire w_dff_A_PAzRvVhk5_2;
	wire w_dff_A_mhv7YP2y6_2;
	wire w_dff_A_YcDjhT8T3_2;
	wire w_dff_A_9tAP6bGr6_2;
	wire w_dff_A_ssWpAkUp1_2;
	wire w_dff_A_XgDTtMqh7_2;
	wire w_dff_A_BgfEetLh3_2;
	wire w_dff_A_OsqZJsAF7_2;
	wire w_dff_A_Jk8JySbY0_2;
	wire w_dff_A_9qaF3s5p9_0;
	wire w_dff_A_7fm7OJu09_0;
	wire w_dff_A_jyxjwfih5_0;
	wire w_dff_A_2S7sEQvu7_0;
	wire w_dff_A_MSD0T39I1_0;
	wire w_dff_A_7Zw8XIoB1_0;
	wire w_dff_A_0HY2OVzG1_0;
	wire w_dff_A_62iO4Jzp4_0;
	wire w_dff_A_CT3P7VP80_0;
	wire w_dff_A_iy7aQw1i7_0;
	wire w_dff_A_KdpGOKs31_0;
	wire w_dff_A_DeriYlGF3_0;
	wire w_dff_A_GtycS8g76_0;
	wire w_dff_A_FMu5tN8o6_2;
	wire w_dff_A_9sHGJc3t5_2;
	wire w_dff_A_NXiR1U0V0_2;
	wire w_dff_A_2sNnIkIh8_2;
	wire w_dff_A_xmUYwhiP2_2;
	wire w_dff_A_O1X7TDLI6_2;
	wire w_dff_A_5SehsGnv5_2;
	wire w_dff_A_yB35zGkT9_2;
	wire w_dff_A_BLaCUOQs4_2;
	wire w_dff_A_ygAWogll4_2;
	wire w_dff_A_KE703snk8_2;
	wire w_dff_A_UR13TOBk4_2;
	wire w_dff_B_TPOkjn7r9_0;
	wire w_dff_B_p8ObpuHO3_0;
	wire w_dff_B_RfTKynf52_0;
	wire w_dff_B_63rkuWgi5_0;
	wire w_dff_B_QEICD4B38_0;
	wire w_dff_B_GMDvtPfY9_0;
	wire w_dff_B_7dm3CGsX4_0;
	wire w_dff_B_sIaBciIM1_0;
	wire w_dff_B_aRrUP5Cf8_0;
	wire w_dff_B_FxrUoyKA7_0;
	wire w_dff_B_h57xBb8Q8_0;
	wire w_dff_B_KGCyfljf0_0;
	wire w_dff_B_byXYpk5q8_0;
	wire w_dff_B_32PVOr4o8_0;
	wire w_dff_B_IBbsAM0P4_0;
	wire w_dff_B_FAo4GoRd6_2;
	wire w_dff_B_hnCBB4eR5_1;
	wire w_dff_B_DyAbswhy2_1;
	wire w_dff_B_jxdHE5yx0_1;
	wire w_dff_A_6aP60U6S4_1;
	wire w_dff_A_fgkpfRl94_1;
	wire w_dff_A_QfBA7mrf1_1;
	wire w_dff_A_OvoeYs2x9_1;
	wire w_dff_A_FBcZg9x53_1;
	wire w_dff_A_Holf9ScS6_1;
	wire w_dff_A_7l85le1F3_1;
	wire w_dff_A_wpAQBJA69_1;
	wire w_dff_A_2AfTwmzk5_1;
	wire w_dff_A_N0ozBPZ51_1;
	wire w_dff_A_66Jggwrk1_1;
	wire w_dff_A_QaoKRL2z1_1;
	wire w_dff_A_JC9hUCkI0_1;
	wire w_dff_A_0wRL0BA83_1;
	wire w_dff_A_wtQfZ54e8_2;
	wire w_dff_A_3s2nxqKQ7_2;
	wire w_dff_A_GWVoku2z4_2;
	wire w_dff_A_8FAIC1IA6_2;
	wire w_dff_A_UNXSZwcO3_2;
	wire w_dff_A_nUGKIQoW7_2;
	wire w_dff_A_OL45Dp2D4_2;
	wire w_dff_A_EIgBiJQD5_2;
	wire w_dff_A_iqcoUGm54_2;
	wire w_dff_A_VAGYgt9E0_2;
	wire w_dff_A_3UeJjg4D4_2;
	wire w_dff_A_VwWoXtQT7_2;
	wire w_dff_A_lVk8emyb5_2;
	wire w_dff_A_2rHcka5g9_2;
	wire w_dff_A_pNqj457g1_1;
	wire w_dff_A_iNC929Ew3_1;
	wire w_dff_A_v0z2JNA78_1;
	wire w_dff_A_ynkmJDs31_1;
	wire w_dff_A_O0fpEPtx0_1;
	wire w_dff_A_WNltdT4J2_1;
	wire w_dff_A_I74UbD4Q0_1;
	wire w_dff_A_AOLGFEfp6_1;
	wire w_dff_A_xnZJRa9L2_1;
	wire w_dff_A_fslFyC5k4_1;
	wire w_dff_A_SpFxxcgd2_1;
	wire w_dff_A_dRVvHzKp6_1;
	wire w_dff_A_QQ3cgWxW8_1;
	wire w_dff_A_PIfmCQ6N7_2;
	wire w_dff_A_xwa0luW98_2;
	wire w_dff_A_tp3c67SQ3_2;
	wire w_dff_A_tE3ebmNO9_2;
	wire w_dff_A_mfoznz4J2_2;
	wire w_dff_A_a7hfHu3R2_2;
	wire w_dff_A_hT1yPn2v2_2;
	wire w_dff_A_Pie7opTS9_2;
	wire w_dff_A_o0Bu0caV0_2;
	wire w_dff_A_g0xY0OlP5_2;
	wire w_dff_A_nTcqnpTW6_2;
	wire w_dff_A_GOdr2Bnl9_2;
	wire w_dff_A_7jshLYJC7_2;
	wire w_dff_B_Sg1nqh8g2_0;
	wire w_dff_B_8itE12jJ8_0;
	wire w_dff_B_2bqiqs3G1_0;
	wire w_dff_B_66y0M8Z94_0;
	wire w_dff_B_oVOUaFwl9_0;
	wire w_dff_B_SNIr9ggv9_0;
	wire w_dff_B_JfUnKVtE0_0;
	wire w_dff_B_z6QokRgv8_0;
	wire w_dff_B_PIOSjjUD6_0;
	wire w_dff_B_ZsuFXeVN4_0;
	wire w_dff_B_zVEyLM8N0_0;
	wire w_dff_B_JDCBK7gm0_0;
	wire w_dff_B_teWfjeAf5_0;
	wire w_dff_B_rfKSEMge0_0;
	wire w_dff_A_tSDqlSZB3_2;
	wire w_dff_B_HxTIoVvv0_2;
	wire w_dff_B_s8OaSu7E6_1;
	wire w_dff_B_6zEZas013_1;
	wire w_dff_B_vOeuLJoV2_1;
	wire w_dff_A_uPx2Fj0u1_0;
	wire w_dff_A_uFQUb5RD5_1;
	wire w_dff_A_Yb84MPbL5_1;
	wire w_dff_B_I9jx0YZ58_0;
	wire w_dff_B_tOBh2K0e2_0;
	wire w_dff_B_FQjJiZYQ9_0;
	wire w_dff_B_GensyDvK0_0;
	wire w_dff_B_cptc2s1c5_0;
	wire w_dff_B_xj22PHBG8_0;
	wire w_dff_B_vPmcNdxc6_0;
	wire w_dff_B_eRivflNn0_0;
	wire w_dff_B_RH4Zyh2w2_0;
	wire w_dff_B_CP3Zu8BA1_0;
	wire w_dff_B_IQNqM0gy0_0;
	wire w_dff_B_Lkey5Jve4_0;
	wire w_dff_B_zFvtv3yL9_0;
	wire w_dff_B_FYUnYL8X0_0;
	wire w_dff_B_1e1NwGhf7_0;
	wire w_dff_B_wGJVb2R39_2;
	wire w_dff_B_kbhrdEkE0_1;
	wire w_dff_B_Ywmvo4SI5_1;
	wire w_dff_B_vCC4io5f0_1;
	wire w_dff_A_GY5BZJ6C9_0;
	wire w_dff_A_W01AA77Q2_0;
	wire w_dff_A_lmW0h3uF2_0;
	wire w_dff_A_YX9lb0hU1_0;
	wire w_dff_A_kZBXivu82_0;
	wire w_dff_A_7m510Wrv0_0;
	wire w_dff_A_Hs43XAUq3_0;
	wire w_dff_A_pFnoTz3C2_0;
	wire w_dff_A_IBbXRGp16_0;
	wire w_dff_A_JJHqbZGP9_0;
	wire w_dff_A_6Y3XtMLv4_0;
	wire w_dff_A_YrhwLuMm5_0;
	wire w_dff_A_IGaPKrFy8_0;
	wire w_dff_A_cCkSWa6R3_0;
	wire w_dff_A_VuEfhJ3T6_2;
	wire w_dff_A_MG3D1TRD1_2;
	wire w_dff_A_Ud2VEXUf0_2;
	wire w_dff_A_6IZqZPyg9_2;
	wire w_dff_A_FGlp4Xtm2_2;
	wire w_dff_A_6GbMvlJj3_2;
	wire w_dff_A_PPwvwhUc5_2;
	wire w_dff_A_aLQqy7yi0_2;
	wire w_dff_A_fbDVu2WR5_2;
	wire w_dff_A_UzVHen974_2;
	wire w_dff_A_wMPb9Ryy0_2;
	wire w_dff_A_TA0Xv2M69_2;
	wire w_dff_A_0BqAqfk73_2;
	wire w_dff_A_MpiDd9nl5_0;
	wire w_dff_A_qdjRQbK42_0;
	wire w_dff_A_DD26uquh0_0;
	wire w_dff_A_Gdm1Zirz0_0;
	wire w_dff_A_cRnDkwLg0_0;
	wire w_dff_A_h01dXzPP6_0;
	wire w_dff_A_toTduXpH7_0;
	wire w_dff_A_j0LIvh7i8_0;
	wire w_dff_A_ukqEtCJK1_0;
	wire w_dff_A_mqLH5R708_0;
	wire w_dff_A_9WNOy34A7_0;
	wire w_dff_A_ZiFLynTk1_0;
	wire w_dff_A_3Q17h9HF4_0;
	wire w_dff_A_u5e2CJke9_2;
	wire w_dff_A_VXp3BJCA6_2;
	wire w_dff_A_6ZMsb2EU6_2;
	wire w_dff_A_a0PoRZX68_2;
	wire w_dff_A_6gUPEj5n4_2;
	wire w_dff_A_J32Kr23S0_2;
	wire w_dff_A_x8InVjLI7_2;
	wire w_dff_A_5u2vZdMK1_2;
	wire w_dff_A_1VsaclCc0_2;
	wire w_dff_A_EgZuTeVk5_2;
	wire w_dff_A_kBEpjhWt0_2;
	wire w_dff_A_KC6qS1y01_2;
	wire w_dff_B_I5TLcTiR9_0;
	wire w_dff_B_6fTDir3V2_0;
	wire w_dff_B_Jwz1yg6a4_0;
	wire w_dff_B_QHHtFVdr8_0;
	wire w_dff_B_u2amd3L69_0;
	wire w_dff_B_QP1psu2c3_0;
	wire w_dff_B_PrVnu9W26_0;
	wire w_dff_B_RLgeHdSq9_0;
	wire w_dff_B_3Pk5V8qq8_0;
	wire w_dff_B_YrQQ7jc00_0;
	wire w_dff_B_3iFp6ebg9_0;
	wire w_dff_B_mzHjuo2t5_0;
	wire w_dff_B_hnIG4mRO0_0;
	wire w_dff_B_qyRUhJ1b1_0;
	wire w_dff_B_y8RlDIqL2_0;
	wire w_dff_B_pFa5jgYj1_1;
	wire w_dff_B_Wz45cKCp9_1;
	wire w_dff_B_TvoVTqyh9_1;
	wire w_dff_A_UMCHUZ8v0_0;
	wire w_dff_A_Pizrzpdm6_0;
	wire w_dff_A_jmdxMLRo3_0;
	wire w_dff_A_w5yFxTCv2_0;
	wire w_dff_A_Nfz1J6KG2_1;
	wire w_dff_A_0sNIWVYG8_0;
	wire w_dff_A_rYzoHzx23_0;
	wire w_dff_A_DN4yzRBO6_0;
	wire w_dff_A_ub3jo0QX4_0;
	wire w_dff_A_wIeQAxNX2_1;
	wire w_dff_A_9otecso84_1;
	wire w_dff_A_Z3m41yRD3_1;
	wire w_dff_A_S2j9JxC38_0;
	wire w_dff_A_P2Xr5Aeo9_0;
	wire w_dff_A_6gFxThkW6_0;
	wire w_dff_A_rdQSBNhP1_0;
	wire w_dff_A_ZlA3nojh2_1;
	wire w_dff_B_5LUGeVFv0_0;
	wire w_dff_B_R5y6A9X89_0;
	wire w_dff_B_kF0Wv8Js3_0;
	wire w_dff_B_NCBxH3Uw1_0;
	wire w_dff_B_BF6TFLkP3_0;
	wire w_dff_B_Mrz1JR5b7_0;
	wire w_dff_B_AVqrgRJA5_0;
	wire w_dff_B_qf99JQde5_0;
	wire w_dff_B_9GZWId6o1_0;
	wire w_dff_B_57bqmZdz0_0;
	wire w_dff_B_8HX3QIPU8_0;
	wire w_dff_B_ZNHaclVH4_0;
	wire w_dff_B_CvCeRqJO4_0;
	wire w_dff_B_cc0SnLEB2_0;
	wire w_dff_B_0GoxrDj70_1;
	wire w_dff_B_4r1oWU3g5_1;
	wire w_dff_B_eHmNBG1g9_1;
	wire w_dff_B_YW2B18rA1_1;
	wire w_dff_B_kVckMQ4n5_1;
	wire w_dff_B_vaRZSY4B9_1;
	wire w_dff_B_tp1CVz8i4_1;
	wire w_dff_B_QJQuMFGs9_1;
	wire w_dff_B_4LTrpdAO9_1;
	wire w_dff_B_OElp9HZj9_1;
	wire w_dff_B_a1wItpK42_1;
	wire w_dff_B_85cD58965_1;
	wire w_dff_B_DDK25lXU2_1;
	wire w_dff_B_UIxyaktK2_1;
	wire w_dff_B_Sxo3aIoO6_1;
	wire w_dff_B_8BAIfOQ66_1;
	wire w_dff_A_eu48OquP3_0;
	wire w_dff_A_t4Fis4ED6_2;
	wire w_dff_B_pLg1x5Uh2_0;
	wire w_dff_B_6Q7NCzT81_1;
	wire w_dff_B_rmn2sUrR2_1;
	wire w_dff_B_iR3KjVcr2_1;
	wire w_dff_B_mp5hQn448_1;
	wire w_dff_B_d8NuR7cB6_1;
	wire w_dff_B_RGYJOLm64_1;
	wire w_dff_B_keGQCtis8_1;
	wire w_dff_B_mOX6zrRQ9_1;
	wire w_dff_B_RlCYQF7t8_1;
	wire w_dff_B_3V60uW6S5_1;
	wire w_dff_B_cF2rsD8Y6_1;
	wire w_dff_B_XlM9oqnq7_1;
	wire w_dff_B_imWam3ti3_1;
	wire w_dff_B_ISUm5JJD8_1;
	wire w_dff_B_lX5igOiU7_1;
	wire w_dff_B_zlpaa5gV7_1;
	wire w_dff_A_dbL7HgUb5_0;
	wire w_dff_A_5gv99wKp5_1;
	wire w_dff_A_Fj9jsS5V1_0;
	wire w_dff_A_JrqsoFpp4_0;
	wire w_dff_A_zlOU3PFR9_0;
	wire w_dff_A_YtguDoaI5_0;
	wire w_dff_A_Pb6fzhMu8_1;
	wire w_dff_A_SnaBn54J6_1;
	wire w_dff_A_ytPiS0pz5_1;
	wire w_dff_A_OSrG8lVv8_1;
	wire w_dff_A_KkYYGaHB2_0;
	wire w_dff_A_lAfnskW83_0;
	wire w_dff_A_SAJoHOUv1_0;
	wire w_dff_A_fjTSXSRj5_0;
	wire w_dff_A_nJlTbF2Y5_0;
	wire w_dff_A_0wWwtRaZ5_1;
	wire w_dff_A_pVYye2o71_1;
	wire w_dff_A_R3I00uET6_1;
	wire w_dff_A_jDTP8mhR3_1;
	wire w_dff_B_RJjV95fk3_3;
	wire w_dff_B_YB1lEoVq0_3;
	wire w_dff_B_vWiWSM1t5_3;
	wire w_dff_B_Y3drOONr1_3;
	wire w_dff_B_LH9e32Fv6_3;
	wire w_dff_B_YUHuGYOJ2_3;
	wire w_dff_B_3wmX0kaV8_0;
	wire w_dff_A_fPXvYNu72_0;
	wire w_dff_A_nbfowXPv7_0;
	wire w_dff_A_dQQ7lR6d4_1;
	wire w_dff_A_Gr1OsUZM4_1;
	wire w_dff_B_SYDnRnlS3_0;
	wire w_dff_B_uOa2Om2A3_0;
	wire w_dff_B_KhXMwgVZ5_0;
	wire w_dff_B_qRoGwaHe0_0;
	wire w_dff_B_Sdsdwj048_0;
	wire w_dff_B_2p7wOymw9_0;
	wire w_dff_B_Axfwu7PD6_0;
	wire w_dff_B_IqrRWfvF6_0;
	wire w_dff_B_aWplygT04_0;
	wire w_dff_B_D0x8W2UY0_0;
	wire w_dff_B_L8RbnZAH0_0;
	wire w_dff_B_z56sPEOa1_0;
	wire w_dff_B_OfaiaSDA2_0;
	wire w_dff_B_DhhOIGEd6_0;
	wire w_dff_B_HmpjpagX4_0;
	wire w_dff_B_kl9TYwy45_2;
	wire w_dff_B_9JfofeCC7_2;
	wire w_dff_B_a6wgwdlZ7_2;
	wire w_dff_B_3OT5K5BX1_1;
	wire w_dff_B_FUvMHAoG8_1;
	wire w_dff_B_Maw3qAoo6_1;
	wire w_dff_B_ZixKtjTy0_1;
	wire w_dff_B_omGMbmO87_1;
	wire w_dff_B_Sb5K7Lkr7_1;
	wire w_dff_B_cXYwp4QC8_1;
	wire w_dff_B_MhK4R2VP5_1;
	wire w_dff_B_lnV2xwj59_1;
	wire w_dff_B_JTVD6QjC1_1;
	wire w_dff_B_0dqQCNPE0_1;
	wire w_dff_B_3KgK7ttF1_1;
	wire w_dff_B_FUlOgvlE4_0;
	wire w_dff_B_sXdgtlN89_0;
	wire w_dff_B_IzmcUFDw6_0;
	wire w_dff_B_NZvyk9B59_0;
	wire w_dff_B_giUEsZHo8_0;
	wire w_dff_B_xbwqmf6Y6_0;
	wire w_dff_B_LaNUnhTa0_0;
	wire w_dff_B_aT3NvJZB9_0;
	wire w_dff_B_doZsvJYt5_0;
	wire w_dff_B_uRSWtzdc4_1;
	wire w_dff_B_2ghFBc636_1;
	wire w_dff_B_mQPe3CN02_1;
	wire w_dff_A_KfgNAJJQ1_0;
	wire w_dff_A_8emau9tp9_0;
	wire w_dff_A_rt8DgwgD2_0;
	wire w_dff_A_94cTNurI0_0;
	wire w_dff_A_mcsujQa73_1;
	wire w_dff_B_eH6XZ9HE6_1;
	wire w_dff_B_99Jp3u7C1_1;
	wire w_dff_B_d1vcH2rp8_1;
	wire w_dff_B_kTa99tev8_1;
	wire w_dff_B_tW1fGQ8W6_1;
	wire w_dff_B_bfYeBHZJ5_1;
	wire w_dff_B_tQhKUQkb1_1;
	wire w_dff_B_qsP9iLyS2_0;
	wire w_dff_B_P0VoA2qX3_0;
	wire w_dff_B_U4764NVg8_0;
	wire w_dff_B_X4qyWCUQ9_0;
	wire w_dff_B_BXVMmKux4_0;
	wire w_dff_B_8miCOP7x2_0;
	wire w_dff_B_xnScEtc77_0;
	wire w_dff_A_GTSqUhit9_1;
	wire w_dff_A_VvpmMaxw4_1;
	wire w_dff_B_XgWeIoQq1_1;
	wire w_dff_B_8itSGbJL9_1;
	wire w_dff_B_zz6sdQL49_1;
	wire w_dff_B_9Jufj2dn4_1;
	wire w_dff_B_WdEBxlLx2_1;
	wire w_dff_A_CsIMUsMA1_0;
	wire w_dff_A_YhaeeRwc3_0;
	wire w_dff_A_fvuRWb520_0;
	wire w_dff_A_PoXbhRtG3_0;
	wire w_dff_A_OZrfM07g6_1;
	wire w_dff_A_MVJX8e971_1;
	wire w_dff_A_jsFtZQH11_1;
	wire w_dff_B_jRkXEa4G8_1;
	wire w_dff_B_hIpkgZVf9_1;
	wire w_dff_B_KprD1YzT0_1;
	wire w_dff_B_LSMEqjdP5_1;
	wire w_dff_B_wyrr0KVs3_1;
	wire w_dff_B_QmSWv1xo5_1;
	wire w_dff_B_q2ZlH6GD6_1;
	wire w_dff_B_UUnfP5AT5_1;
	wire w_dff_B_EvaoAqRi2_1;
	wire w_dff_B_NKhI9E6Q0_1;
	wire w_dff_B_X73lLezi7_1;
	wire w_dff_B_CKPptlEW0_1;
	wire w_dff_B_Ne8oZc1E3_1;
	wire w_dff_B_uPXEjoAm5_1;
	wire w_dff_B_AyFQlIRn2_1;
	wire w_dff_B_geOM1XqB1_1;
	wire w_dff_B_ilvktEQ82_1;
	wire w_dff_B_ueYmJDVK8_1;
	wire w_dff_B_D3cU6MAc4_1;
	wire w_dff_B_pKtBL8wo0_1;
	wire w_dff_B_pPEyHNkF5_1;
	wire w_dff_B_cqMlWShW7_1;
	wire w_dff_B_e7voZlXf7_1;
	wire w_dff_B_JLq5iGFx1_1;
	wire w_dff_B_bF1nBn231_1;
	wire w_dff_B_8v49LUSi5_1;
	wire w_dff_B_mVCr4D5P8_1;
	wire w_dff_B_Muchwt741_1;
	wire w_dff_B_WsIOQDBW7_1;
	wire w_dff_B_ZBHpFyMZ4_1;
	wire w_dff_B_8se2icQt3_1;
	wire w_dff_B_SQcqYZmX4_1;
	wire w_dff_B_Cl0PRBtX8_1;
	wire w_dff_B_F2YdCrcQ2_1;
	wire w_dff_B_iZbEqrwL4_1;
	wire w_dff_B_L7mduJ635_1;
	wire w_dff_B_p8HR99bd4_1;
	wire w_dff_B_20fjxLOe7_1;
	wire w_dff_B_8kpeJ6dk8_1;
	wire w_dff_B_cUsp9VPF8_1;
	wire w_dff_B_HKwz4r8D7_1;
	wire w_dff_B_fyVm4Obu7_1;
	wire w_dff_B_Sf6XW2lO0_1;
	wire w_dff_B_m6C7XxgQ5_1;
	wire w_dff_B_tSjut3WQ4_1;
	wire w_dff_B_GPrc29YB8_1;
	wire w_dff_B_WsOgnKMC5_1;
	wire w_dff_B_qiqA1Udo2_1;
	wire w_dff_B_73X1Uyel6_1;
	wire w_dff_B_IMkZVaau5_1;
	wire w_dff_B_l0lvpBRH7_1;
	wire w_dff_B_GyhXUum03_0;
	wire w_dff_B_mgJ7Dxo54_0;
	wire w_dff_B_4JmHfGlC0_0;
	wire w_dff_B_prtKVrCG4_0;
	wire w_dff_B_uCDM9g1o6_0;
	wire w_dff_B_9LvvXecj4_0;
	wire w_dff_B_7R0hRiq00_1;
	wire w_dff_B_WuaJGEol0_1;
	wire w_dff_B_oANVJYZs4_1;
	wire w_dff_B_DyVAr6xK6_1;
	wire w_dff_B_la9Hy5cp1_1;
	wire w_dff_B_rrZli3ql8_1;
	wire w_dff_B_BF6jpSG08_1;
	wire w_dff_B_nDHupgS93_1;
	wire w_dff_B_bxnokhrt3_1;
	wire w_dff_B_rEPQrDHN1_0;
	wire w_dff_B_xzRqBeyM5_2;
	wire w_dff_B_2NcDcZ4t1_2;
	wire w_dff_B_LbQbXpqE0_2;
	wire w_dff_B_G0TdlR5Q6_0;
	wire w_dff_B_ulbvS3w21_0;
	wire w_dff_B_rxCsvLWZ1_0;
	wire w_dff_B_xb12rojj6_0;
	wire w_dff_B_p7XqTf1S1_0;
	wire w_dff_B_7E62Ck327_0;
	wire w_dff_B_uYJPnmsC3_0;
	wire w_dff_B_6FbSOT536_0;
	wire w_dff_B_OXbUoqo60_0;
	wire w_dff_B_upJEYTwM5_0;
	wire w_dff_B_U7QwuuLY5_0;
	wire w_dff_B_IEVt0auh7_0;
	wire w_dff_B_eG8Y03wf1_0;
	wire w_dff_B_z6GN4o6J4_0;
	wire w_dff_B_bTO4pNdS5_0;
	wire w_dff_B_Z4HedfuY6_2;
	wire w_dff_B_QCywYnxs3_2;
	wire w_dff_B_0c6JP3fR4_2;
	wire w_dff_B_Z3R43VgP3_1;
	wire w_dff_B_qT4UQQcZ1_1;
	wire w_dff_B_5vZSiFMv0_1;
	wire w_dff_B_EKRjpc7W1_1;
	wire w_dff_B_ZT7uiZGu0_1;
	wire w_dff_B_JpGydxwo8_1;
	wire w_dff_B_Xp0iKvHv0_1;
	wire w_dff_B_pGwEHb6S2_1;
	wire w_dff_B_dQ7mUAgC6_1;
	wire w_dff_B_svvvIDDB7_1;
	wire w_dff_B_loHEoTp43_1;
	wire w_dff_B_8k09gzto0_1;
	wire w_dff_B_GPvXg0MZ2_0;
	wire w_dff_B_wLqZL7Tu7_0;
	wire w_dff_B_QwjycpWc7_0;
	wire w_dff_B_i2kKjPjL7_0;
	wire w_dff_B_3vRC0caK2_0;
	wire w_dff_B_KUmo848l3_0;
	wire w_dff_B_N1FDV6gt3_0;
	wire w_dff_B_1mlDaVVb1_0;
	wire w_dff_B_EDvBLAjE8_0;
	wire w_dff_A_aQPlSkov2_1;
	wire w_dff_A_ogj2uxWd9_1;
	wire w_dff_A_2QrO1eFJ5_1;
	wire w_dff_B_ls9Jbc5m9_1;
	wire w_dff_B_dTX8841M8_3;
	wire w_dff_A_ayZfTGbW7_0;
	wire w_dff_A_hKrFVRUb9_0;
	wire w_dff_A_FRRHhxFu1_0;
	wire w_dff_A_q1GhjYhb4_0;
	wire w_dff_A_1iDa6NEo0_0;
	wire w_dff_A_71HeBFXT1_0;
	wire w_dff_A_mjUWrnhX0_0;
	wire w_dff_A_61pbxiN61_0;
	wire w_dff_A_XkHPpHga1_0;
	wire w_dff_A_heEpW0bd2_1;
	wire w_dff_A_prQ93bQ73_1;
	wire w_dff_B_AbTt4sVP2_1;
	wire w_dff_B_STdf4kd25_1;
	wire w_dff_B_k9d95q3R6_1;
	wire w_dff_B_u6wb1a4G8_1;
	wire w_dff_A_5uB1OBD08_0;
	wire w_dff_A_X20EqEFP2_0;
	wire w_dff_A_7210V7iL2_1;
	wire w_dff_A_WX1kDifk3_1;
	wire w_dff_B_8TlBesEM9_1;
	wire w_dff_B_mtf1kKtJ0_1;
	wire w_dff_A_hmk7Jl116_0;
	wire w_dff_A_Jdvyeqj88_2;
	wire w_dff_B_qbT2jZtg7_1;
	wire w_dff_B_2mGFCHHN0_1;
	wire w_dff_B_fYJgsvkO4_1;
	wire w_dff_B_fQU27Otu8_1;
	wire w_dff_B_fvCy5GTE6_1;
	wire w_dff_B_VkPjJjyO6_1;
	wire w_dff_B_KOcVQ9zg7_1;
	wire w_dff_B_rWjubk8T0_1;
	wire w_dff_B_klFXr6gf2_1;
	wire w_dff_B_sZyG1Hue7_1;
	wire w_dff_B_Zwbz9OBi8_1;
	wire w_dff_B_AspQvzbM2_1;
	wire w_dff_B_Gz3wjFV38_1;
	wire w_dff_B_wOBoi8IA9_1;
	wire w_dff_B_fLhK1Rzp7_1;
	wire w_dff_B_3KVuhrsb7_1;
	wire w_dff_B_JPiiHemD4_1;
	wire w_dff_A_gzuh0Vkx4_0;
	wire w_dff_A_aYiZxmTq2_0;
	wire w_dff_A_ktkeExIF9_0;
	wire w_dff_A_sfX1liGi1_0;
	wire w_dff_A_UkKsjaYi3_0;
	wire w_dff_A_IPzIfzM83_1;
	wire w_dff_A_MrX19JTA6_1;
	wire w_dff_A_TfoO0VLG6_1;
	wire w_dff_A_4CBp8hWE2_1;
	wire w_dff_A_TokjpKAi3_1;
	wire w_dff_A_4Xb8R5PN6_1;
	wire w_dff_A_KSXKHMFr5_1;
	wire w_dff_A_va9v80OY8_1;
	wire w_dff_A_xvASDEsW2_2;
	wire w_dff_A_5aatTcDn9_2;
	wire w_dff_A_EOLXLQar4_2;
	wire w_dff_A_8BBXttcs1_2;
	wire w_dff_A_v26VStLg6_2;
	wire w_dff_A_NqJ4XrW94_2;
	wire w_dff_A_gYIti0uh0_2;
	wire w_dff_A_vPH2o0Fx6_2;
	wire w_dff_B_VLxEDSOP3_1;
	wire w_dff_B_WmGzb8lC6_1;
	wire w_dff_A_LgkekKzh6_0;
	wire w_dff_A_EMhafzSt0_2;
	wire w_dff_A_1GrhbAQ60_0;
	wire w_dff_A_FbGtgUkM4_0;
	wire w_dff_A_uT9IiILD1_0;
	wire w_dff_A_2Vlbq6zP4_1;
	wire w_dff_A_aLRzdaaN3_1;
	wire w_dff_B_l5H6hofB7_0;
	wire w_dff_B_hM19lVyP3_0;
	wire w_dff_B_gkyLdtlt2_0;
	wire w_dff_B_1QXHFnVa1_0;
	wire w_dff_B_6TUkHkPM8_0;
	wire w_dff_B_IjZOVqmv6_0;
	wire w_dff_B_VaQRqlkY2_0;
	wire w_dff_B_79tvpKwJ8_0;
	wire w_dff_B_pJdWxdzJ7_0;
	wire w_dff_B_YQnm9lIU5_0;
	wire w_dff_B_lyyle7KZ7_0;
	wire w_dff_B_LdgVtUsB5_0;
	wire w_dff_B_CLCqBe9Z7_0;
	wire w_dff_B_qJoWdEf78_0;
	wire w_dff_B_ILB9o4r96_2;
	wire w_dff_B_xbca8g1s8_2;
	wire w_dff_B_Yf51D3so8_2;
	wire w_dff_B_19CUk0R73_0;
	wire w_dff_B_mUxvoqsy5_1;
	wire w_dff_B_i1CuZtu87_1;
	wire w_dff_B_s5tZkZh78_1;
	wire w_dff_B_EDHVQyou6_1;
	wire w_dff_B_3vonscR97_1;
	wire w_dff_B_9YS5VVDT3_1;
	wire w_dff_B_X6IwygaY6_1;
	wire w_dff_B_fGuWyEnw0_1;
	wire w_dff_B_6m1TaVSt3_1;
	wire w_dff_B_QRrdICxI0_1;
	wire w_dff_B_7hQKRca92_0;
	wire w_dff_B_j5Vcf3KU3_0;
	wire w_dff_B_ZmKB1oqU3_0;
	wire w_dff_B_hMJL2LoC0_0;
	wire w_dff_B_iZowr3dP7_0;
	wire w_dff_B_AYsJGttp0_0;
	wire w_dff_B_yWAWEi9S4_0;
	wire w_dff_B_0ppLAxZZ8_0;
	wire w_dff_A_HIvEGoOw6_1;
	wire w_dff_A_gsEPuZkl3_2;
	wire w_dff_B_1HfbonEU1_0;
	wire w_dff_A_zZPHMM180_0;
	wire w_dff_A_U5gn7ozT5_0;
	wire w_dff_A_mUiANa5l0_0;
	wire w_dff_A_GH6Ko2pe0_0;
	wire w_dff_A_xJ27gl944_0;
	wire w_dff_A_3NAf5tD94_0;
	wire w_dff_A_YoXMoOQg9_0;
	wire w_dff_A_YzfQGdLU0_0;
	wire w_dff_A_Kz347l3Y3_1;
	wire w_dff_A_ZRRNMtCC4_1;
	wire w_dff_A_PcRgOJNS6_1;
	wire w_dff_A_Qmr2zLjk1_0;
	wire w_dff_A_pFcrzKxj4_0;
	wire w_dff_A_epYM8dkX3_0;
	wire w_dff_A_ZpYjSdeL0_2;
	wire w_dff_A_pd2Fzd3t8_2;
	wire w_dff_A_tfnyL9Sh2_2;
	wire w_dff_A_AFUj7jRN3_2;
	wire w_dff_A_ivQD28eW9_2;
	wire w_dff_A_OAgB92s37_2;
	wire w_dff_A_jfWpfTDY8_2;
	wire w_dff_A_vIa3IA8D7_2;
	wire w_dff_A_O9JtnTrn7_2;
	wire w_dff_A_LPew5BSL7_2;
	wire w_dff_A_aaTwBJgH3_0;
	wire w_dff_A_ySZyEEnd2_0;
	wire w_dff_A_AgVAjbLj8_0;
	wire w_dff_A_I9Uio7DV6_1;
	wire w_dff_A_OVor5WGP0_1;
	wire w_dff_A_rWnb6qNO3_1;
	wire w_dff_A_DJ51JjTe3_2;
	wire w_dff_A_LNXDQdP04_2;
	wire w_dff_A_wCJR7GEK4_0;
	wire w_dff_A_MZ0SB1Ps2_0;
	wire w_dff_A_7Vx558mB1_0;
	wire w_dff_A_KdQ8m5yz3_1;
	wire w_dff_B_dq8pL2kY4_3;
	wire w_dff_B_OJWZcLhd3_3;
	wire w_dff_B_7s44NM8a3_3;
	wire w_dff_B_olm5LHQs1_3;
	wire w_dff_B_hcZfaSak9_3;
	wire w_dff_B_eGRdpZ4f2_3;
	wire w_dff_B_GOYTWufs0_3;
	wire w_dff_B_aZlbDHqr4_3;
	wire w_dff_B_sxP123rE8_3;
	wire w_dff_B_aj7JN7wK2_1;
	wire w_dff_B_n8aV7hLb3_1;
	wire w_dff_B_jHBprmgF4_1;
	wire w_dff_B_ww1Bb9T24_1;
	wire w_dff_B_NMJHJAad8_1;
	wire w_dff_B_vzvGqzOA3_1;
	wire w_dff_B_74pk0Hhd3_1;
	wire w_dff_B_A20ilHKs1_1;
	wire w_dff_B_7wfDf1vh2_1;
	wire w_dff_B_VabMyFf63_1;
	wire w_dff_B_w4R4vMFd2_1;
	wire w_dff_B_Z5W0Ta4I1_1;
	wire w_dff_B_Q3TlPJxP2_1;
	wire w_dff_B_h2nWPywg7_1;
	wire w_dff_B_4yEh5cb65_1;
	wire w_dff_B_5gXxx9iH9_1;
	wire w_dff_B_oPnMMCzm4_1;
	wire w_dff_B_bbVZubYC8_1;
	wire w_dff_B_tL06usoO3_1;
	wire w_dff_B_4qdcCPL31_1;
	wire w_dff_B_lViDy4wq4_1;
	wire w_dff_B_DQ2VEUdN9_1;
	wire w_dff_B_uLRIozM67_1;
	wire w_dff_B_Uv48ZgDn4_1;
	wire w_dff_B_ntnPPHuU4_1;
	wire w_dff_B_GtS36WCP5_1;
	wire w_dff_B_twIV5z9g9_1;
	wire w_dff_B_XK3P6TBA8_1;
	wire w_dff_B_vttHX3IB0_1;
	wire w_dff_B_acIVQIkn5_1;
	wire w_dff_B_fqtln7K09_1;
	wire w_dff_A_FvxgaWv24_1;
	wire w_dff_B_cg5oOrxl3_3;
	wire w_dff_B_fTYU1qt46_3;
	wire w_dff_B_FgEDfhrY8_3;
	wire w_dff_B_snmdC2Cj1_3;
	wire w_dff_B_DAGiszlx7_3;
	wire w_dff_A_Z9NEU7h14_0;
	wire w_dff_A_fRRVBTaS4_1;
	wire w_dff_A_1DbhtSJM9_1;
	wire w_dff_B_bC0IgXju0_3;
	wire w_dff_B_sjm3CCUl6_3;
	wire w_dff_B_3uFfUMeF0_3;
	wire w_dff_B_bYGZBYfd5_3;
	wire w_dff_B_rohqyra99_3;
	wire w_dff_B_ektyliWy8_3;
	wire w_dff_B_FOcgl5Ig0_3;
	wire w_dff_B_HqbpNqwJ4_3;
	wire w_dff_B_K8qLVtPj7_3;
	wire w_dff_B_sWMDizUz3_3;
	wire w_dff_A_2uR8uR269_0;
	wire w_dff_A_Z2gtRlb27_0;
	wire w_dff_A_gyfPRPyR1_0;
	wire w_dff_A_gJuftH4B6_0;
	wire w_dff_A_htGz29MJ5_1;
	wire w_dff_A_BdUeDT9A7_1;
	wire w_dff_A_ocZONREd9_1;
	wire w_dff_A_OdaYqszP2_1;
	wire w_dff_A_ndj4ZMr78_0;
	wire w_dff_A_0va8SZaj1_0;
	wire w_dff_A_fGBivi058_0;
	wire w_dff_A_m8v6DEEs9_0;
	wire w_dff_A_HCwU8CDC3_0;
	wire w_dff_A_OePnhah88_0;
	wire w_dff_A_reBb0rZg7_0;
	wire w_dff_A_Og6BaQ0q0_0;
	wire w_dff_A_DCplg5J53_0;
	wire w_dff_A_9g7kbvuQ0_0;
	wire w_dff_A_kmiPpjBM6_0;
	wire w_dff_A_GaxJsdja4_1;
	wire w_dff_B_6DIDidrH7_1;
	wire w_dff_B_DhEh2tGG5_1;
	wire w_dff_B_5MmuVgut9_0;
	wire w_dff_B_HevVietn9_0;
	wire w_dff_B_lGoLgcqN5_0;
	wire w_dff_B_cmkLnFvo7_0;
	wire w_dff_B_c3VDItoR1_0;
	wire w_dff_B_FHZJGFsU5_0;
	wire w_dff_B_fXYcpbP90_0;
	wire w_dff_B_p40PdWak6_0;
	wire w_dff_B_1j1dvsn16_0;
	wire w_dff_B_ZFHAwiAm3_0;
	wire w_dff_B_KxcdlZft6_0;
	wire w_dff_B_65cWIXBY4_0;
	wire w_dff_B_hUtUCUUQ1_0;
	wire w_dff_B_O2wXCame6_0;
	wire w_dff_B_O0bUaAGo0_1;
	wire w_dff_B_RgUjy1Im3_1;
	wire w_dff_B_azXsQYim8_1;
	wire w_dff_B_M85N0d3R5_0;
	wire w_dff_B_aS2Vih3x8_0;
	wire w_dff_B_3vhFUZGe2_0;
	wire w_dff_B_3Czds3JZ4_0;
	wire w_dff_B_8VeSpgzn0_0;
	wire w_dff_B_EjvNbbix8_0;
	wire w_dff_B_NZ8cTK9S6_0;
	wire w_dff_B_hAQsKl8j3_0;
	wire w_dff_B_mmXdeAtT8_0;
	wire w_dff_B_dxH2p7S05_0;
	wire w_dff_B_MORgfw408_0;
	wire w_dff_B_aPJmDf3D1_0;
	wire w_dff_B_SBDAbhRx1_1;
	wire w_dff_B_zjSNR6RA8_1;
	wire w_dff_B_3I40ZzvN4_1;
	wire w_dff_A_vZjRr1JT6_0;
	wire w_dff_A_fZCZTDzz3_0;
	wire w_dff_A_LlDY6nhZ3_0;
	wire w_dff_A_YcAksiy49_1;
	wire w_dff_A_qcE08D9l5_1;
	wire w_dff_A_gmf8R17O2_1;
	wire w_dff_A_nWhYw17j6_0;
	wire w_dff_A_OXZn5mpO3_0;
	wire w_dff_A_J7Y9NuWP2_0;
	wire w_dff_A_UmKEUOuR3_1;
	wire w_dff_A_VhiGAHnE3_1;
	wire w_dff_A_RqxKpO2m6_1;
	wire w_dff_A_BXfgeJqU2_0;
	wire w_dff_A_CyS8Dk7A7_0;
	wire w_dff_B_XtHccHky7_1;
	wire w_dff_B_aMDTVFoh8_1;
	wire w_dff_B_GBfP93RP8_1;
	wire w_dff_B_zWMPtATj4_1;
	wire w_dff_B_XgLeXI1C6_1;
	wire w_dff_B_cWHhm0ZB5_1;
	wire w_dff_B_2QlkjtgU7_1;
	wire w_dff_B_Av4cuTYC5_1;
	wire w_dff_B_YHHqLzvp5_1;
	wire w_dff_B_SdTOLAfJ3_1;
	wire w_dff_B_Lo0ttyBg6_1;
	wire w_dff_B_hyJSHAJk7_1;
	wire w_dff_B_ldIlUEcz3_1;
	wire w_dff_B_g5hIqvbP5_1;
	wire w_dff_B_hCzt0KMs8_1;
	wire w_dff_B_bWI8XA087_1;
	wire w_dff_B_YpajO6WT8_1;
	wire w_dff_B_WSmL8jgO8_1;
	wire w_dff_B_fknJvqcH6_1;
	wire w_dff_B_eVwt8nyF3_1;
	wire w_dff_B_eFyZ6tLA9_1;
	wire w_dff_A_nYSjvWRp9_1;
	wire w_dff_A_gJMNuNEo9_1;
	wire w_dff_A_Vov5Eqjr7_1;
	wire w_dff_A_9oO42x6x2_1;
	wire w_dff_A_SAZg6pwQ3_1;
	wire w_dff_A_FZATdq0d0_1;
	wire w_dff_A_nhAMpXcO2_1;
	wire w_dff_A_XpWiRjSv1_1;
	wire w_dff_A_H4koN1yK6_1;
	wire w_dff_A_aIyR34lZ1_1;
	wire w_dff_A_UAkVqxtG8_1;
	wire w_dff_A_Ox8FuV760_1;
	wire w_dff_A_brTgIcGo0_2;
	wire w_dff_A_BfrDUMvr9_2;
	wire w_dff_A_3y2Y8qjJ8_2;
	wire w_dff_A_7pV8ofrA4_2;
	wire w_dff_A_mZ2chaRB9_2;
	wire w_dff_A_hlHgs7Jf6_2;
	wire w_dff_A_hXs8wCCM1_2;
	wire w_dff_A_DSftXgBI3_2;
	wire w_dff_A_3WfPR8XK6_1;
	wire w_dff_A_5Yf3umdy3_1;
	wire w_dff_A_EWRqoXPE5_1;
	wire w_dff_A_1Vrka3nn3_1;
	wire w_dff_A_0gF9QG569_1;
	wire w_dff_A_wpr6RYoH4_1;
	wire w_dff_A_3NmwBAyE8_1;
	wire w_dff_A_mPQrTci48_2;
	wire w_dff_A_hUqzAPow8_2;
	wire w_dff_A_hOX6vQYZ3_2;
	wire w_dff_B_SunLTDhH8_3;
	wire w_dff_B_NDU8Wrav9_3;
	wire w_dff_B_CFEXWSiw5_3;
	wire w_dff_B_ifJc5Jiq5_3;
	wire w_dff_B_GimFYhXu0_3;
	wire w_dff_B_w6LEIGgm5_3;
	wire w_dff_B_qceph8Jg1_1;
	wire w_dff_B_gqy9HQBB1_1;
	wire w_dff_A_Ny8CW9t27_0;
	wire w_dff_A_I6xnkGRK0_0;
	wire w_dff_A_HOiwcsfq9_0;
	wire w_dff_A_Sy0nyQxk0_0;
	wire w_dff_A_n3XMWM151_0;
	wire w_dff_A_ceGG89cq8_0;
	wire w_dff_A_uv1pBWGx9_0;
	wire w_dff_A_Fnx7eK0y1_0;
	wire w_dff_A_I3jfBtvS7_0;
	wire w_dff_A_sqbawJ0Y8_0;
	wire w_dff_A_ci3ckk8m1_0;
	wire w_dff_A_lQLNx10j0_0;
	wire w_dff_A_taRnpM5n2_0;
	wire w_dff_A_81OM5YjI4_0;
	wire w_dff_A_m3HysKyj2_0;
	wire w_dff_A_rkrxYc2d2_0;
	wire w_dff_A_AQxbrSVC9_1;
	wire w_dff_A_onMi9TXx1_1;
	wire w_dff_A_EpAJ3cIs1_1;
	wire w_dff_A_3i54SPcU4_1;
	wire w_dff_A_9N6E4uSX1_1;
	wire w_dff_A_nxj1Y6cT6_1;
	wire w_dff_A_uA12pxJ92_1;
	wire w_dff_A_ZY4mbvov9_1;
	wire w_dff_A_46c1UTu87_0;
	wire w_dff_A_l57HmlmH3_0;
	wire w_dff_A_5POZ5v0y5_0;
	wire w_dff_A_m7LijZU08_0;
	wire w_dff_A_KhHYVNol9_0;
	wire w_dff_A_nHotHTxJ2_0;
	wire w_dff_A_urAmzmBm2_0;
	wire w_dff_A_w52yENHX9_0;
	wire w_dff_A_yodGdyjF1_0;
	wire w_dff_A_JgmYUvvq4_0;
	wire w_dff_A_IjWZ0cjW0_0;
	wire w_dff_A_G5IAFQDd9_0;
	wire w_dff_A_pZgEnPBt3_0;
	wire w_dff_A_PdO99CxA0_0;
	wire w_dff_A_BOkVioFP1_0;
	wire w_dff_A_P6qfhyQ55_0;
	wire w_dff_A_g64oOjpf2_0;
	wire w_dff_A_PlrVWtov6_0;
	wire w_dff_A_iPVAgh5r5_0;
	wire w_dff_B_b2rcfOAo5_1;
	wire w_dff_B_iJpBJpJC6_1;
	wire w_dff_B_umm4bBqh9_1;
	wire w_dff_B_EuiMQ7PN3_1;
	wire w_dff_B_ob3ULvyY1_1;
	wire w_dff_B_oaXQrTyF6_1;
	wire w_dff_B_zA3ZIGSj0_1;
	wire w_dff_B_PXIRLwyN1_1;
	wire w_dff_B_lXZpWuCN0_1;
	wire w_dff_B_TO98OCIr0_1;
	wire w_dff_B_L3SOA6hu7_1;
	wire w_dff_B_HUfmvg2j8_1;
	wire w_dff_B_zEHCLY6G9_1;
	wire w_dff_B_Dn1zFS835_1;
	wire w_dff_B_za3APN9P7_1;
	wire w_dff_B_tUVxwxxA9_1;
	wire w_dff_B_aBbydeJj2_1;
	wire w_dff_B_bGSCQJIQ0_1;
	wire w_dff_B_mDpCqA5d6_1;
	wire w_dff_B_nj8by4FA8_1;
	wire w_dff_B_0X0GAI739_1;
	wire w_dff_A_JmxG3i3X7_1;
	wire w_dff_A_OpYYQD5b6_1;
	wire w_dff_A_aRJxquyA2_1;
	wire w_dff_A_52sKUUFg7_1;
	wire w_dff_A_7hBvdyLN6_1;
	wire w_dff_A_s0qnuZSx5_1;
	wire w_dff_A_Lu97yoc89_1;
	wire w_dff_A_Lfa3XIpl8_1;
	wire w_dff_A_OzKf7yLM5_1;
	wire w_dff_A_ZR5gk7BB6_1;
	wire w_dff_A_SJBnhBHh9_1;
	wire w_dff_A_TUOlpUU97_1;
	wire w_dff_A_EaFBdXsk9_2;
	wire w_dff_A_mkt2cZNu2_2;
	wire w_dff_A_kzgIon3V5_2;
	wire w_dff_A_7c826gqM9_2;
	wire w_dff_A_v26QQYFn9_2;
	wire w_dff_A_w7FbCt0k0_2;
	wire w_dff_A_rzEmcvym0_2;
	wire w_dff_A_AU70l0BR0_2;
	wire w_dff_A_i0pT8b6p8_1;
	wire w_dff_A_BNdz5W6v2_1;
	wire w_dff_A_K4876BO89_1;
	wire w_dff_A_jZci6xpn7_1;
	wire w_dff_A_fYsXlsdV7_1;
	wire w_dff_A_HyE5cwxc9_1;
	wire w_dff_A_FyeoVdrP6_2;
	wire w_dff_A_iXrQXtt85_2;
	wire w_dff_A_VhhiEz3N5_2;
	wire w_dff_B_zaDwqqmF6_3;
	wire w_dff_B_wOClTlYS3_3;
	wire w_dff_B_24cfXtf52_3;
	wire w_dff_B_waseNjwI4_3;
	wire w_dff_B_DBVmso4B8_3;
	wire w_dff_B_ywEgtm6v0_3;
	wire w_dff_A_WrtBaxLL7_0;
	wire w_dff_B_u5pwc04z4_1;
	wire w_dff_B_pkcCmuYD8_1;
	wire w_dff_A_udlUBLP06_0;
	wire w_dff_A_vzChoUuX1_0;
	wire w_dff_A_PcFUTzKt3_0;
	wire w_dff_A_ow5hqszk7_0;
	wire w_dff_A_kS82MclJ4_0;
	wire w_dff_A_7Dny0Fmu2_0;
	wire w_dff_A_pUE2wtYt5_0;
	wire w_dff_A_MrGUDlWU7_0;
	wire w_dff_A_RXNtSKFm3_0;
	wire w_dff_A_bpOFpYJ53_0;
	wire w_dff_A_i6zAf3cG0_0;
	wire w_dff_A_yKf2mi5S0_0;
	wire w_dff_A_bJUARkVp5_0;
	wire w_dff_A_mEVVDa5N0_0;
	wire w_dff_A_uJPWIQjh3_0;
	wire w_dff_A_aOhPuqhi6_0;
	wire w_dff_A_dpglei4F4_1;
	wire w_dff_A_t0m4ID4x1_1;
	wire w_dff_A_2KOzwYRg4_1;
	wire w_dff_A_IZQsoj7U4_1;
	wire w_dff_A_p2ubC7BX0_1;
	wire w_dff_A_VaIEA5X51_1;
	wire w_dff_A_HgcJxiAs8_1;
	wire w_dff_B_FLJVpyGZ3_2;
	wire w_dff_A_vnoqIWWT6_1;
	wire w_dff_A_pdrTJy1i8_0;
	wire w_dff_A_pRDjoIEm6_0;
	wire w_dff_A_8H1KD62R8_0;
	wire w_dff_A_agSwbR1e5_0;
	wire w_dff_A_4sJq9ubV8_0;
	wire w_dff_A_3kKFd0Ze5_0;
	wire w_dff_A_n6YfRw1H9_0;
	wire w_dff_A_fvRLohg12_0;
	wire w_dff_A_ptnRsuft4_0;
	wire w_dff_A_8NSOpAOV3_0;
	wire w_dff_A_wWmCWJnk6_0;
	wire w_dff_A_i1t2QG4h2_0;
	wire w_dff_A_WCnWyzAE5_0;
	wire w_dff_A_o44IDXQl3_0;
	wire w_dff_A_AkHnZjDH1_0;
	wire w_dff_A_2atQeOyk4_0;
	wire w_dff_A_sdYBnwaJ0_0;
	wire w_dff_A_DjEUFzkF4_0;
	wire w_dff_A_WJPfpayy3_0;
	wire w_dff_B_pJffjcOQ2_1;
	wire w_dff_B_xXhgzhoq6_1;
	wire w_dff_B_Poi6ZA9Y7_1;
	wire w_dff_B_hXHJsLcI2_1;
	wire w_dff_B_TsTuR1uN9_1;
	wire w_dff_B_SuyYcSTo5_1;
	wire w_dff_B_j5GPUGIl5_1;
	wire w_dff_B_Q8jC2qi76_1;
	wire w_dff_B_ABaEJwPX7_1;
	wire w_dff_B_MODYTMI39_1;
	wire w_dff_B_wmFzOJ4K7_1;
	wire w_dff_B_ulVjxbAe7_1;
	wire w_dff_B_PbDOvcpb8_1;
	wire w_dff_B_fi1EYCqG0_1;
	wire w_dff_B_TW288oSk7_1;
	wire w_dff_B_AaXn2NDy6_1;
	wire w_dff_B_mKkKryGu0_1;
	wire w_dff_B_qEMVhYvC0_1;
	wire w_dff_B_lF41FNti2_1;
	wire w_dff_B_KCYizpgs9_1;
	wire w_dff_B_Gnpx6ZxS1_1;
	wire w_dff_B_WoAadTlh5_1;
	wire w_dff_B_tO25t6dS4_1;
	wire w_dff_B_Ar6ZUzHm5_1;
	wire w_dff_B_H7DX6pVw0_1;
	wire w_dff_B_YfBEjTHl2_1;
	wire w_dff_B_d66XZqqJ8_1;
	wire w_dff_B_ppgMSckT3_1;
	wire w_dff_B_4n2AyCD48_1;
	wire w_dff_B_3hb8bEZZ3_1;
	wire w_dff_B_YBuJYGdY9_1;
	wire w_dff_B_w0CSvFMJ9_1;
	wire w_dff_B_PrC8srmz1_1;
	wire w_dff_B_nvqN5uz61_1;
	wire w_dff_B_2ioENHB65_1;
	wire w_dff_B_EMUBajAW9_1;
	wire w_dff_A_8xK8VXFh7_0;
	wire w_dff_A_1aatv5mw9_0;
	wire w_dff_A_puEjy21F4_0;
	wire w_dff_A_UqERjw0i5_0;
	wire w_dff_A_Q6NcDjzu2_0;
	wire w_dff_A_oQrl6rLs7_0;
	wire w_dff_A_iULWfgfT4_0;
	wire w_dff_A_gcXW73iw7_0;
	wire w_dff_A_XUX3r3iv1_0;
	wire w_dff_A_VtkPEHmx9_0;
	wire w_dff_A_k9hWg1wo0_0;
	wire w_dff_A_YwEznwgY8_0;
	wire w_dff_A_cRUsgrtb4_1;
	wire w_dff_A_BuoCDXTF6_1;
	wire w_dff_A_oheE48JG9_1;
	wire w_dff_A_Oy5oOTlU2_1;
	wire w_dff_A_1pa8uRPx7_1;
	wire w_dff_A_hh5YWipl6_1;
	wire w_dff_A_GOfz4csY9_1;
	wire w_dff_A_jMuMy8Wk7_1;
	wire w_dff_A_hmqJmvhe9_1;
	wire w_dff_A_bxFPa8u93_1;
	wire w_dff_A_WfuOkAOV8_1;
	wire w_dff_A_iIvhlGgr9_1;
	wire w_dff_A_6QchqKpk5_1;
	wire w_dff_A_dC3enEGa0_1;
	wire w_dff_A_HqZ9htgT0_1;
	wire w_dff_A_CfthQPG70_1;
	wire w_dff_A_cObrOEkK4_1;
	wire w_dff_A_09DbJUja3_1;
	wire w_dff_A_4dLxQPcd1_1;
	wire w_dff_A_DUsB57ym2_1;
	wire w_dff_A_GYmrlpJv3_1;
	wire w_dff_A_fffNOiRE9_1;
	wire w_dff_A_egOg8bec8_1;
	wire w_dff_A_OM7OUMoI5_1;
	wire w_dff_A_qUsJx8Qp0_1;
	wire w_dff_A_sIofJAnO1_1;
	wire w_dff_A_bMj26oXv2_2;
	wire w_dff_A_gfaXRvDY4_2;
	wire w_dff_A_d5ywrFJG8_2;
	wire w_dff_A_aKHTaF592_2;
	wire w_dff_A_2HjCF51g9_2;
	wire w_dff_A_ADMGUHmx8_2;
	wire w_dff_A_cnw3HkUX6_2;
	wire w_dff_A_TcitEqyr9_2;
	wire w_dff_A_wxwLr7ba7_2;
	wire w_dff_A_VpcbP0Cs6_2;
	wire w_dff_A_4vJo3Nhw6_2;
	wire w_dff_A_6sIYz1BS8_2;
	wire w_dff_A_xU9ffot83_2;
	wire w_dff_A_iJo7wsB24_2;
	wire w_dff_A_qnFqvISH0_1;
	wire w_dff_A_74tlJx2G5_1;
	wire w_dff_A_Q37oWraE4_1;
	wire w_dff_A_3mmU56vm8_1;
	wire w_dff_A_LITqAKQa6_1;
	wire w_dff_A_h44018j13_1;
	wire w_dff_A_KOXHWqVg0_1;
	wire w_dff_A_TXcFZWv89_1;
	wire w_dff_A_KU4MEAzF4_1;
	wire w_dff_A_94TvaCZy6_1;
	wire w_dff_A_UTp8sruD6_1;
	wire w_dff_A_qPTMqRIg5_1;
	wire w_dff_A_IAF5Qtnl9_1;
	wire w_dff_A_Ocg1H20t9_2;
	wire w_dff_A_GLKjOtYb7_2;
	wire w_dff_A_n81TeKAl8_2;
	wire w_dff_A_ViFLau3t7_2;
	wire w_dff_A_2I9S8XQp6_2;
	wire w_dff_A_C3OqboqI7_2;
	wire w_dff_A_VvoNm4nn9_2;
	wire w_dff_A_0O2kpQdZ4_2;
	wire w_dff_A_8376GmCA9_2;
	wire w_dff_A_XlDx9OSS6_1;
	wire w_dff_A_xkrDxope0_1;
	wire w_dff_A_nGqoYRDg4_1;
	wire w_dff_A_YgZ58kRh5_1;
	wire w_dff_A_7LyVNPUy3_1;
	wire w_dff_A_jECS5YH59_1;
	wire w_dff_A_LnrAmqGP8_1;
	wire w_dff_A_dzJXTCCT9_1;
	wire w_dff_A_f0rXsL5M1_1;
	wire w_dff_A_a728PDv13_1;
	wire w_dff_A_ttFflHNJ8_1;
	wire w_dff_A_n4lnK1VF4_1;
	wire w_dff_A_x75IVeFP2_1;
	wire w_dff_A_9kvR0RHU7_1;
	wire w_dff_A_Ub4t46gV0_1;
	wire w_dff_A_G8NnnIVa3_1;
	wire w_dff_A_JptWlgdZ2_1;
	wire w_dff_A_OZ4fZ4xv6_1;
	wire w_dff_A_5eaAx21E9_1;
	wire w_dff_A_f405pS0G7_1;
	wire w_dff_A_7h0amuuZ1_0;
	wire w_dff_A_o5wOCgQ61_0;
	wire w_dff_A_8ybaW9IF6_0;
	wire w_dff_A_0ChQ87o71_0;
	wire w_dff_A_LbZ03N6A8_0;
	wire w_dff_A_vbvg9F0Z0_0;
	wire w_dff_A_yn9tlmaF7_0;
	wire w_dff_A_H5kKxkqm6_2;
	wire w_dff_A_vItqtTeF6_2;
	wire w_dff_A_Vbwb1EMG9_2;
	wire w_dff_A_w9MX6vb47_2;
	wire w_dff_A_Od3aWPll0_2;
	wire w_dff_A_xvTRKp3k9_2;
	wire w_dff_A_XJgAsCsE9_2;
	wire w_dff_A_5R0xYeGe7_2;
	wire w_dff_A_J62SNFk35_2;
	wire w_dff_A_Eh8SxKZM5_2;
	wire w_dff_A_ySTgQNO37_2;
	wire w_dff_A_KK8seJc28_2;
	wire w_dff_A_9Y6mym4t4_2;
	wire w_dff_A_V4SPeXWY4_2;
	wire w_dff_A_eKCvZG224_2;
	wire w_dff_A_ZGEwQbOp8_2;
	wire w_dff_A_YjWwCsyN2_1;
	wire w_dff_A_amHV6v8B9_1;
	wire w_dff_A_avyApZ9t5_1;
	wire w_dff_A_uzOaPsZv1_1;
	wire w_dff_A_qKu5EPsF5_1;
	wire w_dff_A_wNrZFBS95_1;
	wire w_dff_A_XVpHqNjm7_1;
	wire w_dff_A_Fy9rEV3l5_1;
	wire w_dff_A_wjoPMRhT6_1;
	wire w_dff_A_nLoa28D20_1;
	wire w_dff_A_KhwDJsyE7_1;
	wire w_dff_A_QXu7rwtx6_1;
	wire w_dff_A_Cg8fNTzH5_2;
	wire w_dff_A_duePGjtb9_2;
	wire w_dff_A_BoSfbFG50_2;
	wire w_dff_A_yxkdMpGz0_2;
	wire w_dff_A_FzKve4SU4_2;
	wire w_dff_A_Px1p9vNX5_2;
	wire w_dff_A_77eWdI954_2;
	wire w_dff_A_HYv2veyb9_2;
	wire w_dff_A_vbkxWPKJ6_2;
	wire w_dff_B_g1NZdqsi7_1;
	wire w_dff_B_T4yHuf3p1_1;
	wire w_dff_B_B4sIOW8K3_1;
	wire w_dff_B_TTFgYehI2_1;
	wire w_dff_B_rcFwh1Hh7_1;
	wire w_dff_B_RS0J7QR09_1;
	wire w_dff_B_JslYyxcs4_1;
	wire w_dff_B_YOdUTLAu9_1;
	wire w_dff_B_vxD1Olrk3_1;
	wire w_dff_B_kCsAirVz0_1;
	wire w_dff_B_zY7v3CCW5_1;
	wire w_dff_B_wHJSwFaZ5_1;
	wire w_dff_B_CAgiRPfG3_1;
	wire w_dff_B_LhugXMuJ7_1;
	wire w_dff_B_PJTbO05R6_1;
	wire w_dff_B_POLCdHC48_1;
	wire w_dff_B_yM3NqG9g3_1;
	wire w_dff_B_O7Z1AKZ68_1;
	wire w_dff_B_lb5dKOg98_1;
	wire w_dff_B_O5E94j3c4_1;
	wire w_dff_B_jXMyg2c55_1;
	wire w_dff_B_R1Wkhd6v8_1;
	wire w_dff_B_1X07Wmza9_1;
	wire w_dff_B_hlgieTYN3_1;
	wire w_dff_B_buQdeXio7_1;
	wire w_dff_B_y5vdR8xS0_1;
	wire w_dff_B_uz9elGk93_1;
	wire w_dff_B_sOcVv01b4_1;
	wire w_dff_B_uCZ8kTj63_1;
	wire w_dff_B_7o671Esm1_1;
	wire w_dff_B_ofgYCHXe7_1;
	wire w_dff_B_pdIoJ7S96_1;
	wire w_dff_B_7MPljmG90_1;
	wire w_dff_B_u18zMVPH2_1;
	wire w_dff_B_0598kKp94_1;
	wire w_dff_B_hGr6wSUJ7_1;
	wire w_dff_B_fPissgFc5_0;
	wire w_dff_B_TFlZORKh3_0;
	wire w_dff_B_RY666wF85_0;
	wire w_dff_B_7dnT8Qwg9_0;
	wire w_dff_B_g6AtUCyW1_0;
	wire w_dff_B_cloTSarb4_0;
	wire w_dff_B_r29TzAEK4_0;
	wire w_dff_B_YvNukTC68_0;
	wire w_dff_B_0dkMnsUl1_0;
	wire w_dff_B_RHNi9xVM6_0;
	wire w_dff_B_xPLCufXR0_0;
	wire w_dff_B_eSl6CPWI9_0;
	wire w_dff_B_gk2FnGnp0_0;
	wire w_dff_B_vNEaLbEW9_0;
	wire w_dff_B_LR7OJ1I74_0;
	wire w_dff_B_DjlpOAtG3_0;
	wire w_dff_B_hV5agPxn8_0;
	wire w_dff_B_QZw4TMhB7_0;
	wire w_dff_B_VkeaUpgj9_0;
	wire w_dff_B_shnPEXPY1_0;
	wire w_dff_B_px5ZdUIe7_0;
	wire w_dff_B_0Nr7RXnD4_0;
	wire w_dff_B_Rqgp33VM1_0;
	wire w_dff_B_iv4zvYdQ6_1;
	wire w_dff_A_K26thiWr8_0;
	wire w_dff_B_pOQmJj3U1_1;
	wire w_dff_A_qS9klzNj2_1;
	wire w_dff_A_k3JB3iCB9_0;
	wire w_dff_B_UnBdhMhv8_1;
	wire w_dff_B_TTFTocGu1_2;
	wire w_dff_A_GApiUB9Q9_0;
	wire w_dff_A_WA0s8Mnc6_0;
	wire w_dff_B_ojyNWK7c7_1;
	wire w_dff_B_eZqKCXTv8_1;
	wire w_dff_A_xQfn7MGY8_1;
	wire w_dff_B_rGnss2399_1;
	wire w_dff_A_3YLb6Y9c1_1;
	wire w_dff_B_F8AqNKUb9_0;
	wire w_dff_B_a3QL1NSg6_0;
	wire w_dff_B_VjOJsnXf6_0;
	wire w_dff_B_rk4d4Bjk7_0;
	wire w_dff_B_OzS5BOtS0_0;
	wire w_dff_A_ltpBvl6H1_0;
	wire w_dff_A_cB9ztAZT6_0;
	wire w_dff_A_2JdLEy3j5_0;
	wire w_dff_A_HpiOvwHi4_1;
	wire w_dff_A_rgcPklOv7_1;
	wire w_dff_A_9FMqmy381_1;
	wire w_dff_A_OWQkBT059_1;
	wire w_dff_A_FhEXZ4ZW6_1;
	wire w_dff_A_38JcmSs84_1;
	wire w_dff_A_wCRS4pXC5_1;
	wire w_dff_A_tVNUeOV68_1;
	wire w_dff_A_HhRntZwZ4_1;
	wire w_dff_A_bZyt1uXS4_1;
	wire w_dff_A_WV7wOBFw4_1;
	wire w_dff_B_Snf1LqFt0_0;
	wire w_dff_B_jMQYmiD85_0;
	wire w_dff_B_cw8LeY8W6_0;
	wire w_dff_B_Jh3TekGu0_0;
	wire w_dff_A_HyanecyJ0_0;
	wire w_dff_A_53lSuFD73_0;
	wire w_dff_A_8IqcREHf8_0;
	wire w_dff_B_V58b9dXk3_0;
	wire w_dff_B_pVM2lMhF9_1;
	wire w_dff_A_SF2gKTs29_0;
	wire w_dff_A_hCMtiU4E1_0;
	wire w_dff_A_SehYSrqj3_0;
	wire w_dff_A_foB81kUL3_0;
	wire w_dff_A_jHvo7Xlk4_0;
	wire w_dff_A_PwUBuEfH9_0;
	wire w_dff_B_T3sxnq1M5_1;
	wire w_dff_B_qYaK45dp7_1;
	wire w_dff_B_ZUAYicvz0_1;
	wire w_dff_B_5mPxYXIv3_0;
	wire w_dff_B_fdGNECGl8_0;
	wire w_dff_B_8e85yDFP6_0;
	wire w_dff_B_d3LsgjpI8_1;
	wire w_dff_A_WwVYqvUf4_0;
	wire w_dff_A_5dDgk8ii0_0;
	wire w_dff_B_uNP6423W8_2;
	wire w_dff_A_Q8QOtOSR2_0;
	wire w_dff_B_b6pFW9900_3;
	wire w_dff_B_1QNdUh026_3;
	wire w_dff_A_Fwgg2QO98_1;
	wire w_dff_A_5nqX0Onf0_1;
	wire w_dff_A_9Oj3ozNS6_1;
	wire w_dff_A_FaTiuKzn8_1;
	wire w_dff_A_QrF8qCpc9_1;
	wire w_dff_A_tLWPBBaU6_1;
	wire w_dff_A_QTSfA3wV0_1;
	wire w_dff_A_7xNlXekK5_2;
	wire w_dff_A_WXrc9FmN1_2;
	wire w_dff_A_ypQB3onv6_2;
	wire w_dff_A_Kfw9dmFK2_2;
	wire w_dff_A_pvFXFeQb3_2;
	wire w_dff_A_ILyOpGBO9_2;
	wire w_dff_A_JjMk9zlO8_1;
	wire w_dff_A_0H4spKl57_1;
	wire w_dff_A_dEErKEAa2_1;
	wire w_dff_A_raMBdhc38_2;
	wire w_dff_A_5GC5YbDb3_2;
	wire w_dff_B_xUii6bHv2_1;
	wire w_dff_B_9bgltcn55_1;
	wire w_dff_B_VZZTiSp49_1;
	wire w_dff_B_eNGpBWf86_1;
	wire w_dff_B_fRw42wEj5_1;
	wire w_dff_B_zsdy9Zl82_1;
	wire w_dff_A_50hmwSDu7_2;
	wire w_dff_A_9kVgspdK1_2;
	wire w_dff_A_vhzWELfx7_2;
	wire w_dff_A_e4X0ADm52_2;
	wire w_dff_A_OXBJvEML1_2;
	wire w_dff_A_tg4nSsv12_2;
	wire w_dff_A_ZmXU0taD4_2;
	wire w_dff_A_O57uuZ4N1_2;
	wire w_dff_A_yb7Rrzvm3_1;
	wire w_dff_A_l9btvlHH5_1;
	wire w_dff_A_YtBF5r7W8_1;
	wire w_dff_A_tFxOJqQM1_1;
	wire w_dff_A_tLdKHldY0_1;
	wire w_dff_A_hIUaBKai6_1;
	wire w_dff_A_xjVBSbwO5_1;
	wire w_dff_A_GNJrBlpy1_2;
	wire w_dff_A_NkL8CpXt2_1;
	wire w_dff_A_pYkteeSe7_1;
	wire w_dff_B_WYHw19yU4_2;
	wire w_dff_B_bSGZwCqE4_2;
	wire w_dff_B_X0R6Lci53_0;
	wire w_dff_A_75SbOFsv8_1;
	wire w_dff_A_ZdDOikhV5_1;
	wire w_dff_B_c2vrybp85_1;
	wire w_dff_B_Tw5JmFPd0_1;
	wire w_dff_B_e2WDhi7A7_1;
	wire w_dff_B_UO8pbqDg9_1;
	wire w_dff_A_QpH1FV798_1;
	wire w_dff_A_jTs244OI7_1;
	wire w_dff_A_xhbIWgCU4_1;
	wire w_dff_A_SXc5389j0_1;
	wire w_dff_A_hPXqXdMT6_0;
	wire w_dff_A_IPnPPsxj1_0;
	wire w_dff_A_PNJXGsJi1_1;
	wire w_dff_A_4L6nhCvO8_1;
	wire w_dff_B_aWKtNM9w2_1;
	wire w_dff_B_V7Kax62f0_3;
	wire w_dff_A_yyZ7EeFx5_0;
	wire w_dff_A_IFGDUsUK7_0;
	wire w_dff_A_3hgCUxs04_1;
	wire w_dff_A_AOtu1sjH4_1;
	wire w_dff_A_HCs8vNtd3_1;
	wire w_dff_A_DiOjrdAz9_1;
	wire w_dff_A_jvyrUwuN8_1;
	wire w_dff_A_Xpu7Qeg40_2;
	wire w_dff_A_XbTzPN4r2_2;
	wire w_dff_A_EE610UcN3_2;
	wire w_dff_B_0moUcKQS9_3;
	wire w_dff_B_0gyQMMzy0_3;
	wire w_dff_B_wgle9SfE6_3;
	wire w_dff_B_gmsZvxHJ0_3;
	wire w_dff_B_YUyPreZ66_3;
	wire w_dff_B_kshmEO0R7_3;
	wire w_dff_B_33bhuAvl8_3;
	wire w_dff_A_q4NEHzuz9_0;
	wire w_dff_A_tT6hAK6U7_0;
	wire w_dff_A_BrgZqVO46_0;
	wire w_dff_A_4UhCQXfS6_0;
	wire w_dff_A_aujhon4S8_0;
	wire w_dff_A_OThn2ABh0_0;
	wire w_dff_A_blw3zNgs9_0;
	wire w_dff_A_WWV3D3Pb2_0;
	wire w_dff_A_5oUjxY3r0_0;
	wire w_dff_A_lsRdNO4i9_0;
	wire w_dff_A_HftPVBkU4_0;
	wire w_dff_A_aXXG4IeB4_1;
	wire w_dff_A_CjNDb0Us0_1;
	wire w_dff_A_vgwD9PvH1_1;
	wire w_dff_A_HSb0cIJS1_1;
	wire w_dff_A_z1hpwgbH6_1;
	wire w_dff_A_AKymWHSA7_1;
	wire w_dff_A_dEf9Dms78_1;
	wire w_dff_B_OpOkjfm44_0;
	wire w_dff_B_1pkzOlgn8_0;
	wire w_dff_A_5VmbqH5C2_0;
	wire w_dff_A_HHssrEh99_0;
	wire w_dff_A_BCuU1Rr21_0;
	wire w_dff_B_znryO9ie9_2;
	wire w_dff_A_67QwtZ6x4_0;
	wire w_dff_A_VgQhHTKt5_0;
	wire w_dff_A_GewbPXuV0_1;
	wire w_dff_A_iBUMR8Ew2_1;
	wire w_dff_A_HNSQBfCa2_1;
	wire w_dff_A_BTCzLtU25_1;
	wire w_dff_A_Gv755MUa6_0;
	wire w_dff_A_sCyLSq6K7_0;
	wire w_dff_A_nUcGYgwi3_0;
	wire w_dff_A_VtPrfV8H4_0;
	wire w_dff_A_QzxyHL7W6_0;
	wire w_dff_A_pfeWfZUr8_2;
	wire w_dff_A_67GSnaxY0_2;
	wire w_dff_A_SokhPaHg7_2;
	wire w_dff_A_8pzO0rXC3_1;
	wire w_dff_A_bow1sMlW8_1;
	wire w_dff_B_TRF4NlcU8_1;
	wire w_dff_B_MF1kEDRA6_1;
	wire w_dff_B_67dmE65F9_1;
	wire w_dff_B_hbgrprrW0_1;
	wire w_dff_A_BFctmDTz3_1;
	wire w_dff_A_zNwLQdnp5_1;
	wire w_dff_A_4osPnoRv1_1;
	wire w_dff_A_ttlHbz9T1_1;
	wire w_dff_B_TBImO6FS6_0;
	wire w_dff_B_OF3KwrDd9_0;
	wire w_dff_B_aVgFD1dL9_1;
	wire w_dff_A_h3z2YUrv4_2;
	wire w_dff_A_IUNEtqDF8_1;
	wire w_dff_A_FUCJ8oFp2_1;
	wire w_dff_A_1B2tUJY09_1;
	wire w_dff_A_1btaIGhu2_1;
	wire w_dff_A_TJSNIQ1X7_2;
	wire w_dff_A_z9A9yAvg2_2;
	wire w_dff_A_x1trZjX05_2;
	wire w_dff_A_OezKpDzA1_2;
	wire w_dff_A_r31cBjW88_0;
	wire w_dff_A_JWWby9fX1_0;
	wire w_dff_B_VydjEBBC5_3;
	wire w_dff_B_Xxy0llxD2_3;
	wire w_dff_A_kNM03czV2_0;
	wire w_dff_A_CC5zD9ys5_0;
	wire w_dff_B_iO5cs4jZ7_1;
	wire w_dff_B_McNbNlnj5_1;
	wire w_dff_A_rJlRsTwe4_0;
	wire w_dff_B_7V7pwQqq8_2;
	wire w_dff_A_HP5uExgC5_0;
	wire w_dff_A_DybV0qOA6_0;
	wire w_dff_A_9u4yvsA51_1;
	wire w_dff_A_klxydncY7_1;
	wire w_dff_A_gI5B2grv5_1;
	wire w_dff_A_faQzdlrd2_1;
	wire w_dff_A_M7bze1R01_1;
	wire w_dff_A_0voaKU4p9_1;
	wire w_dff_A_oXvTveG19_2;
	wire w_dff_A_dflQyUH87_2;
	wire w_dff_A_nGeZXjpX6_2;
	wire w_dff_A_0VnuRAWd0_2;
	wire w_dff_A_mQMoIth09_2;
	wire w_dff_B_QlA5UopO3_0;
	wire w_dff_B_r1zOMHRi2_0;
	wire w_dff_B_fshypG5j3_1;
	wire w_dff_A_Q6s4J0Ok9_0;
	wire w_dff_A_NemSBIxA4_1;
	wire w_dff_A_UwMNUtlo7_1;
	wire w_dff_A_h7wfmPoq5_2;
	wire w_dff_A_cMvc9Qws4_2;
	wire w_dff_A_HIWORh2d2_2;
	wire w_dff_A_k3vSyhWN3_2;
	wire w_dff_A_sgODAPR95_0;
	wire w_dff_B_tS6mCmRe0_0;
	wire w_dff_A_AuRtYqI56_0;
	wire w_dff_A_eAEeDcZA9_1;
	wire w_dff_A_hNwrlskJ5_1;
	wire w_dff_B_of19NiuT7_1;
	wire w_dff_A_tUR2AhzW3_0;
	wire w_dff_A_AJsusLjk2_0;
	wire w_dff_A_xm5kZ9st4_2;
	wire w_dff_A_LnjJ634u3_0;
	wire w_dff_A_00MTdIt77_0;
	wire w_dff_A_LwvZZmhx1_2;
	wire w_dff_A_z1gmnbMd3_2;
	wire w_dff_A_CLGdv8Ko1_0;
	wire w_dff_A_tG7bxNfY2_1;
	wire w_dff_A_PsHvd5hW2_2;
	wire w_dff_A_tWNU14720_0;
	wire w_dff_A_mDu6K7KB9_0;
	wire w_dff_A_0VsX9gSj1_2;
	wire w_dff_A_22TePM3N9_2;
	wire w_dff_A_K3Qbqy7G6_0;
	wire w_dff_B_Y6uJcumH7_1;
	wire w_dff_A_d0mXA9PV1_0;
	wire w_dff_A_oJvT7yWN6_1;
	wire w_dff_A_FW533wll0_1;
	wire w_dff_A_ppkAAw5J0_2;
	wire w_dff_B_heec8Ysv9_3;
	wire w_dff_A_ynpSuS5k6_0;
	wire w_dff_A_sHe4h7fx4_0;
	wire w_dff_A_pxelVl3Z0_1;
	wire w_dff_A_RZ5VYcc30_1;
	wire w_dff_A_236AP8nm2_1;
	wire w_dff_A_tWoPz4ME8_1;
	wire w_dff_A_zrSjxQI90_2;
	wire w_dff_A_mckreH0L8_2;
	wire w_dff_A_gRoyY9iG4_1;
	wire w_dff_A_n3Pl6qdE0_1;
	wire w_dff_A_x5eB3vcn8_1;
	wire w_dff_A_ELEi7V7m7_1;
	wire w_dff_A_k5dAjeXQ4_1;
	wire w_dff_A_11KyuPkZ3_1;
	wire w_dff_A_N68OXoit7_1;
	wire w_dff_A_qYgJoz2A4_1;
	wire w_dff_A_sUq2AmRE2_1;
	wire w_dff_A_kvH05xRp7_1;
	wire w_dff_A_LtwD0vNX5_0;
	wire w_dff_A_GEsH3DP62_0;
	wire w_dff_A_p7EyMcTN4_2;
	wire w_dff_A_jvNcSafF1_1;
	wire w_dff_A_Udpa4Dlm8_1;
	wire w_dff_A_LSWA4SK34_1;
	wire w_dff_A_iYbMZzK97_1;
	wire w_dff_B_EV41gs3b0_0;
	wire w_dff_B_dCZwKOI10_0;
	wire w_dff_A_Oz1kqe4N9_1;
	wire w_dff_A_jOXfclfh5_1;
	wire w_dff_A_PD6kO0Ym0_2;
	wire w_dff_A_x0IUNIDN8_0;
	wire w_dff_A_K44uDDF16_0;
	wire w_dff_A_DvWIhjLR1_0;
	wire w_dff_A_JxeyMOSj2_0;
	wire w_dff_A_T7tHFmi49_2;
	wire w_dff_A_WcQnB2JF9_0;
	wire w_dff_A_nRuNkL557_0;
	wire w_dff_A_PFfUAP3b8_0;
	wire w_dff_A_CVj66qHQ4_0;
	wire w_dff_A_pula1oiE2_0;
	wire w_dff_A_osDBOpXY5_0;
	wire w_dff_A_Q6r4r7rb3_0;
	wire w_dff_A_umhkggfb1_0;
	wire w_dff_A_jTzFy5wh3_0;
	wire w_dff_A_yCuGPY7Q1_0;
	wire w_dff_A_CzWOorUO5_0;
	wire w_dff_A_mmVvdwBw5_0;
	wire w_dff_A_bOzkJjjs5_0;
	wire w_dff_A_hj3Pxhih1_0;
	wire w_dff_A_Ft5dKWl73_0;
	wire w_dff_A_u5ptFPJO7_0;
	wire w_dff_A_0c2haayH0_0;
	wire w_dff_A_PsXMDqsn9_2;
	wire w_dff_A_8Iwc0BAH6_2;
	wire w_dff_A_2xvx20Dz2_2;
	wire w_dff_B_B180yI9l9_0;
	wire w_dff_B_wa4N5EPW1_0;
	wire w_dff_B_I6Vmu5Qf7_0;
	wire w_dff_B_EmxxxWDC5_0;
	wire w_dff_B_VH6yGqaa3_0;
	wire w_dff_B_AUeL5z2w3_0;
	wire w_dff_B_lZPwmdJr5_0;
	wire w_dff_B_m0LBZ8ps8_0;
	wire w_dff_B_H7y67g0v5_0;
	wire w_dff_B_V825YOW41_0;
	wire w_dff_B_nwpjwDy64_0;
	wire w_dff_B_wanWD0270_0;
	wire w_dff_B_ytyy4KYs9_0;
	wire w_dff_B_bkjl5Xja4_1;
	wire w_dff_B_G2zMsgd27_1;
	wire w_dff_B_XrdMZr1n8_1;
	wire w_dff_B_tVYseWYk3_1;
	wire w_dff_B_o5Sivf2n5_1;
	wire w_dff_B_PYbTzFi39_1;
	wire w_dff_B_1WUmjhl90_0;
	wire w_dff_B_umz6snDn7_0;
	wire w_dff_B_ptrbJwoT9_1;
	wire w_dff_B_klZCwMge2_1;
	wire w_dff_B_KVxKDGVU1_1;
	wire w_dff_B_L5oVnzO48_1;
	wire w_dff_B_pk3vYg6W7_0;
	wire w_dff_A_duw3mAMP8_0;
	wire w_dff_A_RIzvgUbT6_1;
	wire w_dff_A_fbotVb362_1;
	wire w_dff_A_9V0wUiED8_1;
	wire w_dff_A_BFAkwIrk5_1;
	wire w_dff_A_hHwEEgIP3_1;
	wire w_dff_A_hpqvISpo6_1;
	wire w_dff_A_jBj7RvZ02_1;
	wire w_dff_A_jwKbbin55_1;
	wire w_dff_A_USAtdbCA6_1;
	wire w_dff_A_MOvyumZz3_1;
	wire w_dff_A_ZGWavH5e8_2;
	wire w_dff_A_LrKwF3DL8_2;
	wire w_dff_A_vmsZkfZI1_2;
	wire w_dff_B_RCuyKb0I8_1;
	wire w_dff_B_LFGWI0nG2_1;
	wire w_dff_B_LKZCUakw4_1;
	wire w_dff_B_GCIUjCEb3_1;
	wire w_dff_A_z9nyDZ5I5_0;
	wire w_dff_A_tvJ5pTrB9_1;
	wire w_dff_A_02E25KrJ1_1;
	wire w_dff_A_YdvRnKQC1_1;
	wire w_dff_A_MbcZdtJF0_1;
	wire w_dff_A_77v8mn7W1_1;
	wire w_dff_A_B77uRN4V4_0;
	wire w_dff_A_1xSnFRRZ7_0;
	wire w_dff_A_UUoHSVdh5_0;
	wire w_dff_A_gndSIIHq5_0;
	wire w_dff_A_DaFQTWao4_0;
	wire w_dff_A_SVP84Jxj8_0;
	wire w_dff_A_ybkX4O3d6_0;
	wire w_dff_A_c8BxFHsH8_0;
	wire w_dff_A_RfEBFwxt1_0;
	wire w_dff_A_uFn72zPK9_0;
	wire w_dff_A_a3aub9DV0_0;
	wire w_dff_B_yPMzt06f5_2;
	wire w_dff_A_eQKtaybn8_1;
	wire w_dff_A_0l2Sv8Ge0_1;
	wire w_dff_A_SsqQ17Nc6_1;
	wire w_dff_A_QbxZYPDn2_1;
	wire w_dff_A_hH69EzeS0_1;
	wire w_dff_A_L4AHDBsg0_1;
	wire w_dff_B_KTcfb66q6_0;
	wire w_dff_B_sb7ax8Z62_0;
	wire w_dff_B_6l8Es9rU3_1;
	wire w_dff_A_rPMYSFAn3_0;
	wire w_dff_A_uX3tdavN5_0;
	wire w_dff_A_6uAxBoPZ0_2;
	wire w_dff_A_vpZNlNcy9_2;
	wire w_dff_A_cCq4LzdO9_2;
	wire w_dff_B_YBkNYZOG6_1;
	wire w_dff_B_VWEEJY1S1_1;
	wire w_dff_A_5gwSCMZM8_0;
	wire w_dff_A_4wNAwRAf9_0;
	wire w_dff_A_tVHTqF3h4_0;
	wire w_dff_B_rEpscLp15_2;
	wire w_dff_A_OdkKpBji1_2;
	wire w_dff_A_XqoSx2Ot9_2;
	wire w_dff_A_bluO7SOM9_2;
	wire w_dff_B_Ol8i2kYi7_2;
	wire w_dff_A_k86KeRhH0_1;
	wire w_dff_B_ez15tSP66_0;
	wire w_dff_B_Rvnwe1wD7_0;
	wire w_dff_B_Bfz9YGEj0_1;
	wire w_dff_B_qSDASetN6_0;
	wire w_dff_B_vi8uLsP27_0;
	wire w_dff_B_JUCzJ7sa9_1;
	wire w_dff_A_TrHiYAnk6_1;
	wire w_dff_A_L2wK5FBO0_0;
	wire w_dff_A_T52GB4Ep1_0;
	wire w_dff_B_CoCtGuNQ8_2;
	wire w_dff_A_PL9bxoyz9_0;
	wire w_dff_A_E2bAMQPb5_1;
	wire w_dff_A_plI47xaI9_1;
	wire w_dff_A_OdD1Xs1X1_1;
	wire w_dff_A_hoaHWpBQ4_1;
	wire w_dff_A_Vg9ppsk36_2;
	wire w_dff_A_HmoeU2K61_2;
	wire w_dff_A_JHbzWgM82_2;
	wire w_dff_A_JSKQu7Ck0_2;
	wire w_dff_B_6sMTLta98_0;
	wire w_dff_B_wzqnqoXo6_0;
	wire w_dff_B_2rOS53rP8_0;
	wire w_dff_B_EZuZnK921_0;
	wire w_dff_B_MIfKNEgW7_0;
	wire w_dff_B_Bci5bNEN8_0;
	wire w_dff_B_0cOJAhcX5_0;
	wire w_dff_B_o79XuoKI2_1;
	wire w_dff_B_R6T6ydsP1_0;
	wire w_dff_B_kyzhpD2z1_0;
	wire w_dff_B_as1BGSdU2_0;
	wire w_dff_B_a5rfNWOn7_0;
	wire w_dff_A_x9GwPzIU3_0;
	wire w_dff_A_JE3qdwRv2_0;
	wire w_dff_B_eaoXcS7P6_2;
	wire w_dff_B_J3UtZMY82_2;
	wire w_dff_B_p9whTygG0_2;
	wire w_dff_B_UaKwaDPw5_2;
	wire w_dff_B_sMBNa4lp7_2;
	wire w_dff_B_u1wcZca27_2;
	wire w_dff_B_Nl6AlKv06_2;
	wire w_dff_B_4p4PURqQ7_2;
	wire w_dff_B_2Wbpd6sD9_2;
	wire w_dff_A_7bwjDdvK2_0;
	wire w_dff_A_7qPjqhdK9_0;
	wire w_dff_A_jczKTll98_0;
	wire w_dff_A_Aok4hIju0_0;
	wire w_dff_A_btxep7797_0;
	wire w_dff_A_qZJYF48m2_0;
	wire w_dff_A_O2MWxzCe1_0;
	wire w_dff_A_Cp2LwsjL6_0;
	wire w_dff_A_Sbe6xNlx1_0;
	wire w_dff_A_ZjZ2DZ7l8_0;
	wire w_dff_A_K1zS4y1F5_0;
	wire w_dff_A_Zt4aQlix2_1;
	wire w_dff_A_I00WpwUb5_1;
	wire w_dff_A_g1Svti6l9_1;
	wire w_dff_A_DrpQAFGN2_1;
	wire w_dff_A_7Mj91jPD4_1;
	wire w_dff_A_lI3RzP6B5_1;
	wire w_dff_A_PODq0vZL2_1;
	wire w_dff_A_V13W4NhE3_1;
	wire w_dff_A_ODvgMo6Y2_1;
	wire w_dff_B_sOIUIeEh4_1;
	wire w_dff_B_rXtbchKY7_0;
	wire w_dff_A_xh1MlD5z4_0;
	wire w_dff_A_x94Gyz5M4_2;
	wire w_dff_A_rhu1SLX75_2;
	wire w_dff_A_VMAvBlKx6_2;
	wire w_dff_A_otpvEPg61_1;
	wire w_dff_A_VmCc0SdF6_1;
	wire w_dff_A_gspL3bJU9_1;
	wire w_dff_B_JGqTnb7k3_0;
	wire w_dff_B_xbfNDrb60_0;
	wire w_dff_B_s1Lg2lHD0_1;
	wire w_dff_B_U8dG6jcS2_0;
	wire w_dff_A_usuy5aFg9_0;
	wire w_dff_B_HQmzkpsW9_2;
	wire w_dff_A_AyQKETKV8_1;
	wire w_dff_A_End4mDRM1_1;
	wire w_dff_A_a0Lwgxvx6_1;
	wire w_dff_A_khTp7iO64_1;
	wire w_dff_A_mdmMYsyg7_1;
	wire w_dff_A_633fGYG73_1;
	wire w_dff_A_DfkzCR1E7_1;
	wire w_dff_B_weWeD51m0_0;
	wire w_dff_A_n64hHnDN6_1;
	wire w_dff_A_KwzCzioj9_1;
	wire w_dff_A_JZ5umaZO8_2;
	wire w_dff_A_gGE1DTIe7_2;
	wire w_dff_A_8m8VzK7g3_2;
	wire w_dff_B_75ERfvS76_0;
	wire w_dff_B_RJyCFA7L9_0;
	wire w_dff_B_Z0FhR6SO8_1;
	wire w_dff_A_AbPZAwis7_1;
	wire w_dff_A_TtdV9xNS0_0;
	wire w_dff_B_SVP5Y5N34_0;
	wire w_dff_B_CkHicxHn5_0;
	wire w_dff_B_P5UkVFyp5_0;
	wire w_dff_A_DZ4rb1pn2_2;
	wire w_dff_A_RqEWupQx7_2;
	wire w_dff_B_uCsSlT233_1;
	wire w_dff_A_KiCxKFaz6_0;
	wire w_dff_A_AoskPmD63_1;
	wire w_dff_A_6zW5vQiK3_1;
	wire w_dff_A_m3dvtZfp2_1;
	wire w_dff_B_5UMaX4ZM0_1;
	wire w_dff_B_Rd6uJHVp0_1;
	wire w_dff_B_dEl6L4no0_0;
	wire w_dff_A_92TCUL8i1_1;
	wire w_dff_B_WqTalyok5_0;
	wire w_dff_A_1iQtT2Lb3_1;
	wire w_dff_A_wZAo4vm67_1;
	wire w_dff_B_H8GXBcUn2_1;
	wire w_dff_A_lQRMyj9D2_0;
	wire w_dff_A_gGnrurns2_1;
	wire w_dff_A_SRqVufOq5_1;
	wire w_dff_B_N5KTHUmM9_1;
	wire w_dff_A_F8hozB7X3_0;
	wire w_dff_A_QCsdzEps4_1;
	wire w_dff_A_VCHzWWBO2_1;
	wire w_dff_B_xvI34cRN7_1;
	wire w_dff_B_OaFX81gL2_0;
	wire w_dff_B_8xCPJpTY7_1;
	wire w_dff_A_XZylqcdf9_0;
	wire w_dff_A_zngNaiEX2_1;
	wire w_dff_A_SrzM1ZCC3_1;
	wire w_dff_B_glHv4Be06_3;
	wire w_dff_A_0e8Tz4Da4_0;
	wire w_dff_A_Nen14reh1_0;
	wire w_dff_A_SLOptLUN8_0;
	wire w_dff_A_29KEvHpM3_0;
	wire w_dff_A_1AcOq1Na9_1;
	wire w_dff_A_dVbwrVjr4_1;
	wire w_dff_A_m5XaaJW91_1;
	wire w_dff_A_UpmAJVRc9_1;
	wire w_dff_A_s37Gi0y91_2;
	wire w_dff_A_stElDjSk7_2;
	wire w_dff_A_btWbsP4p8_2;
	wire w_dff_A_wCHQqrQ66_2;
	wire w_dff_A_eCxoAzf34_2;
	wire w_dff_B_RYzTC9Qw3_1;
	wire w_dff_A_k924Gbdg9_1;
	wire w_dff_A_ynWu1gvJ3_1;
	wire w_dff_B_Jd8Y8iK58_3;
	wire w_dff_A_ENpVegIb2_0;
	wire w_dff_A_BPiz1hj92_0;
	wire w_dff_A_6oM2yfUC7_0;
	wire w_dff_A_ewlGzfSJ4_0;
	wire w_dff_A_hiaybn1G9_1;
	wire w_dff_A_SE6sVdrN9_1;
	wire w_dff_B_9sfsuSSR1_1;
	wire w_dff_A_8zdwvfop7_0;
	wire w_dff_A_HOf4kQdV8_1;
	wire w_dff_A_cQUCsWo01_2;
	wire w_dff_A_LM8TSfZa7_2;
	wire w_dff_A_Zhpq7rLM0_2;
	wire w_dff_A_penQLU6r8_2;
	wire w_dff_A_ayZZV8Mh8_0;
	wire w_dff_B_DrhtTbPM2_1;
	wire w_dff_A_hSJTcLhb5_0;
	wire w_dff_A_A5K82NNl8_2;
	wire w_dff_A_IGkRkcEo3_2;
	wire w_dff_A_21qrzfBF6_2;
	wire w_dff_B_2Ugq5SDK0_3;
	wire w_dff_A_4en0RrWo9_0;
	wire w_dff_A_UaZNyiSJ8_0;
	wire w_dff_A_9eAdTEaV6_1;
	wire w_dff_A_6QueWslw8_1;
	wire w_dff_A_lnyqTAaI3_2;
	wire w_dff_A_0u4JD2Gl6_2;
	wire w_dff_A_2yAw5N0q6_2;
	wire w_dff_A_OW3w21rU4_2;
	wire w_dff_A_Hk7IFeeq8_2;
	wire w_dff_B_OQMF5acT7_1;
	wire w_dff_B_2EtDnD859_1;
	wire w_dff_A_cjOigGYo4_0;
	wire w_dff_A_PUPbGg4F4_0;
	wire w_dff_A_pWTYFmGH7_1;
	wire w_dff_A_tBxglOLO9_1;
	wire w_dff_A_MZY9Vevh7_1;
	wire w_dff_A_0GvYtfUI6_1;
	wire w_dff_A_t3r0Xzeu5_2;
	wire w_dff_A_8HkfzeEk4_2;
	wire w_dff_A_NIY42FNy3_0;
	wire w_dff_B_Cp9r5I7Y0_1;
	wire w_dff_B_DtwF8QNr1_1;
	wire w_dff_B_HSff3Y947_1;
	wire w_dff_A_LHGc20gx9_0;
	wire w_dff_A_B6Hz6mmi1_1;
	wire w_dff_A_PNelFTlN8_1;
	wire w_dff_A_xoOMif9N4_1;
	wire w_dff_B_JkwMTCpa0_3;
	wire w_dff_A_YWRSlTvL2_0;
	wire w_dff_A_dYJCZRIB4_0;
	wire w_dff_A_OrtdOlk18_0;
	wire w_dff_A_zI9PDHAN4_0;
	wire w_dff_A_nYRQNxeO5_1;
	wire w_dff_A_Vy5T5x4G7_1;
	wire w_dff_A_285xZoKg6_1;
	wire w_dff_A_sleKAM1H8_1;
	wire w_dff_A_skKD6xIe2_2;
	wire w_dff_A_oViVnr2g9_2;
	wire w_dff_A_OGIteHFE9_2;
	wire w_dff_A_Z4jqWwkk4_2;
	wire w_dff_A_ufYN7Zob3_2;
	wire w_dff_B_A039z5SO3_1;
	wire w_dff_A_bjpd9y5w2_0;
	wire w_dff_A_CMqjyJc04_1;
	wire w_dff_A_FrwNMP6u2_1;
	wire w_dff_B_jUzy2tsp4_3;
	wire w_dff_A_PxqJO5hw7_0;
	wire w_dff_A_qfppex116_0;
	wire w_dff_A_jZfgkex86_0;
	wire w_dff_A_Sgh0BycS8_0;
	wire w_dff_A_O7RXdq8e7_1;
	wire w_dff_A_6XZQcvXs7_1;
	wire w_dff_A_mwTnOLeO1_1;
	wire w_dff_A_KMlWaPwz4_1;
	wire w_dff_A_r9tMHijF2_2;
	wire w_dff_A_nUbNzVq17_2;
	wire w_dff_A_dWNlxkLb4_2;
	wire w_dff_A_04DJAaSG2_2;
	wire w_dff_A_nUkqtVwk2_2;
	wire w_dff_B_07KldbNH7_1;
	wire w_dff_B_dULN66I59_3;
	wire w_dff_A_9tFWFHYi0_0;
	wire w_dff_A_sRjpLi1M0_0;
	wire w_dff_A_TYVHvv0x4_0;
	wire w_dff_A_ddJZg2O26_0;
	wire w_dff_A_c8Uegmih4_1;
	wire w_dff_A_6PT9UaPV7_1;
	wire w_dff_B_m86AmQ6o9_1;
	wire w_dff_A_igLneryp8_0;
	wire w_dff_A_pKnYCdRQ0_0;
	wire w_dff_A_hnZVdOah8_2;
	wire w_dff_A_2ZG2lwal3_1;
	wire w_dff_A_aPfAbq2E5_2;
	wire w_dff_A_4uQpMDMp0_2;
	wire w_dff_A_aV5iv32c8_2;
	wire w_dff_A_F0aoAc7Z5_2;
	wire w_dff_A_p5KaWxUz0_1;
	wire w_dff_A_28hBAJIf9_2;
	wire w_dff_B_RfWK9qRM9_1;
	wire w_dff_A_tmfqrQf33_0;
	wire w_dff_B_dbez48296_3;
	wire w_dff_A_Qa2dTJtU4_0;
	wire w_dff_A_tSSnMQyO4_0;
	wire w_dff_A_UvCznFnx1_0;
	wire w_dff_A_iT0XC6JC1_0;
	wire w_dff_A_icIKl32y3_1;
	wire w_dff_A_AYOFg4f10_1;
	wire w_dff_A_lSwGBZ3P3_1;
	wire w_dff_A_N7rosL8O5_1;
	wire w_dff_A_zOUCRTkq8_2;
	wire w_dff_A_yE0fdLE20_2;
	wire w_dff_A_OpVGVuUx8_2;
	wire w_dff_A_xG4huGW33_2;
	wire w_dff_A_35IMdrIP4_2;
	wire w_dff_A_d4OfE2S05_0;
	wire w_dff_A_eePLoI0R8_1;
	wire w_dff_A_yHUCZuC37_2;
	wire w_dff_B_IfxoEAop5_1;
	wire w_dff_A_JXrCIJvl2_0;
	wire w_dff_A_6pD16Eak7_1;
	wire w_dff_A_TGig5Ra66_2;
	wire w_dff_B_y2eLDWYg9_3;
	wire w_dff_A_M0w1qVb91_0;
	wire w_dff_A_H2IaVxAx0_0;
	wire w_dff_A_q5diUuo23_0;
	wire w_dff_A_YTcr934E7_0;
	wire w_dff_A_nuWETZuz2_0;
	wire w_dff_A_cQUuhADp8_0;
	wire w_dff_A_LmPcdkiY6_2;
	wire w_dff_A_pMF7ZgcW6_2;
	wire w_dff_A_6FuuZyO67_1;
	wire w_dff_A_x7sGiAdx3_2;
	wire w_dff_A_8w6nNEqq5_2;
	wire w_dff_A_rxPgrNyV1_1;
	wire w_dff_A_cNoIiuvb4_1;
	wire w_dff_A_1jd7x19Q3_1;
	wire w_dff_A_6o6y199y8_1;
	wire w_dff_A_cwmGlU5W8_1;
	wire w_dff_A_41ACyzYg9_1;
	wire w_dff_A_A3zQ4tk19_1;
	wire w_dff_A_ZrgidNM39_1;
	wire w_dff_A_qlGK1zUc2_1;
	wire w_dff_A_A5S280Jx3_1;
	wire w_dff_A_Fgb2w0BH6_1;
	wire w_dff_A_q5RmSlfg8_1;
	wire w_dff_A_dw7vFQVK4_1;
	wire w_dff_A_A35gOGjj3_2;
	wire w_dff_A_fnaYPgvu8_2;
	wire w_dff_A_88nBEgWt0_2;
	wire w_dff_A_S5mqmuTU2_2;
	wire w_dff_A_megjtH8p1_2;
	wire w_dff_A_jKQg6Bzu4_2;
	wire w_dff_A_M17gvMOR8_1;
	wire w_dff_A_8MyeU4p57_1;
	wire w_dff_A_RwmHz5dF8_2;
	wire w_dff_A_knUKgd3s9_2;
	wire w_dff_A_ldal8IrY6_1;
	wire w_dff_A_gPehqFNi3_2;
	wire w_dff_A_D9J3qCLC2_2;
	wire w_dff_A_eqHfnncg7_0;
	wire w_dff_A_RVF50Q914_0;
	wire w_dff_A_b4pEDyG90_0;
	wire w_dff_A_jgyoAhAo8_0;
	wire w_dff_A_ki72DMDT7_0;
	wire w_dff_A_EhPNGhGT5_0;
	wire w_dff_A_PwyVWGro2_0;
	wire w_dff_A_zLfcPr794_0;
	wire w_dff_A_gTTEjKUO8_0;
	wire w_dff_A_RKSBBxJA8_0;
	wire w_dff_A_JNsW3kQF0_1;
	wire w_dff_A_6XeykArG8_1;
	wire w_dff_A_eTnnq1VJ1_1;
	wire w_dff_A_K662OT5o9_1;
	wire w_dff_A_5juf2MdT5_1;
	wire w_dff_A_XXhFatY62_1;
	wire w_dff_A_k5UnAS1S9_1;
	wire w_dff_A_snpIkSUm6_1;
	wire w_dff_A_5g0c3fXV9_1;
	wire w_dff_A_NwjZZOGG4_1;
	wire w_dff_A_AejevhVk9_1;
	wire w_dff_A_OrmFKQiS4_1;
	wire w_dff_A_6RrIfPak4_1;
	wire w_dff_A_g7QYx8QW5_1;
	wire w_dff_A_bnX6o2SG7_1;
	wire w_dff_A_sS9p3uYW1_1;
	wire w_dff_A_mRgHOw5y3_1;
	wire w_dff_A_8XNAnQuR4_2;
	wire w_dff_A_qZxqNWs10_2;
	wire w_dff_A_bmhauP1P5_2;
	wire w_dff_A_AkGAOCEU5_2;
	wire w_dff_A_bQgOdBIg8_2;
	wire w_dff_A_CnavchMN2_2;
	wire w_dff_A_uyKqCI4e6_2;
	wire w_dff_A_DCvm9Jp54_2;
	wire w_dff_A_9YFfn4a95_2;
	wire w_dff_A_8xMWlhgR6_2;
	wire w_dff_A_LQ8hzgDA8_2;
	wire w_dff_A_9YRwvugD1_2;
	wire w_dff_A_VzLreYgr4_2;
	wire w_dff_A_xNoEALuA2_2;
	wire w_dff_A_UbJTOfwr6_2;
	wire w_dff_A_6FTyiP646_2;
	wire w_dff_A_UIjB0zyY5_2;
	wire w_dff_A_bOJsdiR19_2;
	wire w_dff_A_UBaovMR50_2;
	wire w_dff_A_S5ECTJ9d4_2;
	wire w_dff_A_SDm1thEd8_2;
	wire w_dff_A_CiHQhXAV7_2;
	wire w_dff_A_lcXMExnl1_1;
	wire w_dff_A_F65Acl362_0;
	wire w_dff_A_i0oV3XBq1_0;
	wire w_dff_A_snNBHj0t4_0;
	wire w_dff_A_kEfVqUx53_0;
	wire w_dff_A_JEwSdVin5_0;
	wire w_dff_A_TQvhzHIO7_0;
	wire w_dff_A_zrzRwFII8_0;
	wire w_dff_A_AuMGgbfJ1_0;
	wire w_dff_A_KYRcokFw2_0;
	wire w_dff_A_LcG0xPmX8_0;
	wire w_dff_A_mX3aNj423_0;
	wire w_dff_A_9ZG8s6Sg5_0;
	wire w_dff_A_QukYTuNX7_2;
	wire w_dff_A_SPBSTZgc6_2;
	wire w_dff_A_0bta0lHL3_2;
	wire w_dff_A_4QQCIver8_2;
	wire w_dff_A_kUq32hEe8_2;
	wire w_dff_A_KPvFGWBZ2_2;
	wire w_dff_A_EJ0zEH3n7_2;
	wire w_dff_A_B06BWju75_2;
	wire w_dff_A_LO8UWQR42_2;
	wire w_dff_A_8zre90L10_1;
	wire w_dff_A_7ydOL1c61_1;
	wire w_dff_A_q0t9VMXc4_1;
	wire w_dff_A_ksNc1iY76_1;
	wire w_dff_A_wffFOdSi9_1;
	wire w_dff_A_YaGHig3H8_1;
	wire w_dff_A_u3D6O5KS0_1;
	wire w_dff_A_GU6ZFazo1_1;
	wire w_dff_A_2D7vCtPn4_1;
	wire w_dff_A_R3482hnf5_1;
	wire w_dff_A_NPysg0Ys9_1;
	wire w_dff_A_Nv2vdjzc6_1;
	wire w_dff_A_QjwkVGAL1_1;
	wire w_dff_A_YIwVEM0L8_1;
	wire w_dff_A_cIZq431Z6_1;
	wire w_dff_A_DR3U9k6v4_1;
	wire w_dff_A_HlNI22Kk6_1;
	wire w_dff_A_H6j9jbvz4_2;
	wire w_dff_A_O6IDgJcS2_2;
	wire w_dff_A_1TCpeAM55_2;
	wire w_dff_A_isMvM8cf3_2;
	wire w_dff_A_vrhIlXCD6_2;
	wire w_dff_A_3bxwuoaJ1_2;
	wire w_dff_A_cs4Q6h1Q4_2;
	wire w_dff_A_zA4o0ooZ6_2;
	wire w_dff_A_GA2HNsza2_2;
	wire w_dff_A_7m5TB6Hu8_2;
	wire w_dff_A_wUErHdW35_2;
	wire w_dff_A_txNEyoiR7_2;
	wire w_dff_A_IPMSuDzf2_2;
	wire w_dff_A_smbwUTM68_2;
	wire w_dff_A_i63KIdhp9_1;
	wire w_dff_A_EWHvyPZ43_1;
	wire w_dff_A_R62Qy0032_1;
	wire w_dff_A_1MyqPzEA3_1;
	wire w_dff_A_HUcL8UEe1_1;
	wire w_dff_A_iKs1Z2Sm7_1;
	wire w_dff_A_XZvDag2a6_1;
	wire w_dff_A_jlxOl8lR9_1;
	wire w_dff_A_qtHWGnv13_1;
	wire w_dff_A_wSTKM3NH4_1;
	wire w_dff_A_ggyk9r9m9_1;
	wire w_dff_A_6SweCnPu6_1;
	wire w_dff_A_BDIoTfWJ6_1;
	wire w_dff_A_bXRX2Atc4_2;
	wire w_dff_A_R7p5KH6R4_2;
	wire w_dff_A_6qA5t5FI6_2;
	wire w_dff_A_Z2wR5NnP2_2;
	wire w_dff_A_dj7r3Jwf1_2;
	wire w_dff_A_TowleIEi1_2;
	wire w_dff_A_uzoQmpYe7_2;
	wire w_dff_A_k7brtZ6F5_2;
	wire w_dff_A_ctauFzo35_2;
	wire w_dff_A_IlVo0zOt8_1;
	wire w_dff_A_o45xLZWt3_1;
	wire w_dff_A_3DUBTaA16_1;
	wire w_dff_A_C2zHLIrd9_1;
	wire w_dff_A_3HhAzPlm5_1;
	wire w_dff_A_buTNbRHs9_1;
	wire w_dff_A_o4grvfCh0_1;
	wire w_dff_B_L5yK2An24_2;
	wire w_dff_B_NlFn00mt7_2;
	wire w_dff_A_pW95h57B1_1;
	wire w_dff_A_rLR0GM5D0_1;
	wire w_dff_A_X2vG03Rq7_1;
	wire w_dff_A_rVCZxvPw7_1;
	wire w_dff_A_ArLHnBfi5_1;
	wire w_dff_A_CuZygEpU4_1;
	wire w_dff_A_xYijioYp3_1;
	wire w_dff_A_i4VqygTe9_1;
	wire w_dff_A_tm973Edl8_1;
	wire w_dff_A_d6J6DxjB6_1;
	wire w_dff_A_C3D2yfgo8_1;
	wire w_dff_A_M9Qz2cnI1_1;
	wire w_dff_A_5U9Gkiec9_1;
	wire w_dff_A_g4KbrXBc9_1;
	wire w_dff_A_TS2FEWC16_1;
	wire w_dff_A_ffOTLJoC2_1;
	wire w_dff_A_BKUf7AhY0_1;
	wire w_dff_A_1f13skSO0_1;
	wire w_dff_A_aQCxkdfb3_1;
	wire w_dff_A_gU3g5sc85_2;
	wire w_dff_A_SA0aRm868_0;
	wire w_dff_A_hlsP0tkn5_0;
	wire w_dff_A_yEN9h9Ia0_0;
	wire w_dff_A_xC4n3mcC6_0;
	wire w_dff_A_iIBkXhEP4_0;
	wire w_dff_A_q4Cjv6fi9_0;
	wire w_dff_A_phz25t3F0_0;
	wire w_dff_A_gi3NMY6U2_0;
	wire w_dff_A_ZWXnm81p5_0;
	wire w_dff_A_WEuSM3HY6_0;
	wire w_dff_A_x5nFVwmE1_1;
	wire w_dff_A_KykJahah3_1;
	wire w_dff_A_l3SNMPq15_1;
	wire w_dff_A_iNnfzujs5_1;
	wire w_dff_A_wEyEDtv12_1;
	wire w_dff_A_KQEVPLUt0_1;
	wire w_dff_A_ZY0JdPxh1_1;
	wire w_dff_A_nUQmyL3F4_1;
	wire w_dff_A_FelI4awa8_1;
	wire w_dff_A_9W1IDtR54_1;
	wire w_dff_A_xymTSAXO9_1;
	wire w_dff_A_5oOWpqjS6_1;
	wire w_dff_A_9LYk3EoK9_2;
	wire w_dff_A_qf8uLdAk2_2;
	wire w_dff_A_1MQCro9E7_2;
	wire w_dff_A_1nU3WNDh3_2;
	wire w_dff_A_2rmSXgSW0_2;
	wire w_dff_A_mM8ZiayI8_2;
	wire w_dff_A_QNQfnR0t9_2;
	wire w_dff_A_zm4VkXNN3_2;
	wire w_dff_A_cQyQM5eZ8_2;
	wire w_dff_A_6kqBPqRu1_2;
	wire w_dff_A_tJva2PYj6_2;
	wire w_dff_A_XeKFCu0r5_2;
	wire w_dff_A_d3R4En5E1_2;
	wire w_dff_A_EwsDexbo7_2;
	wire w_dff_A_BbMNcHjw6_2;
	wire w_dff_A_iZXm6Txu5_2;
	wire w_dff_A_4hGzf6Sl6_1;
	wire w_dff_A_Mu3YnyXy6_1;
	wire w_dff_A_AP9auKRN9_1;
	wire w_dff_A_rKbTQJGZ6_1;
	wire w_dff_A_BET9gSeQ8_1;
	wire w_dff_A_oR4Wcep23_1;
	wire w_dff_A_whE6azjg4_1;
	wire w_dff_A_1ME0lkkO0_1;
	wire w_dff_A_FVri9oHp2_1;
	wire w_dff_A_wAZfXtje8_1;
	wire w_dff_A_rpLuG0iX9_1;
	wire w_dff_A_RulbiuaA4_1;
	wire w_dff_A_Dyg1rBGL7_2;
	wire w_dff_A_nOtk7jjB4_2;
	wire w_dff_A_zLp1h93Q8_2;
	wire w_dff_A_hG2bJ7Ph4_2;
	wire w_dff_A_m6syC80A3_2;
	wire w_dff_A_6jFDG3866_2;
	wire w_dff_A_HVvWM4KM0_2;
	wire w_dff_A_riK0dFw99_2;
	wire w_dff_A_4Py8OvaH9_2;
	wire w_dff_B_Jzd9k4Fx3_2;
	wire w_dff_B_6m41WtIX8_2;
	wire w_dff_B_Xt0mqTLH7_2;
	wire w_dff_B_uYZGv2q40_2;
	wire w_dff_B_GU1dWDT25_2;
	wire w_dff_B_RYSmBXTS4_2;
	wire w_dff_B_tn5PMLcw8_2;
	wire w_dff_B_1yTd4z8I9_2;
	wire w_dff_B_xQZbUEyq2_2;
	wire w_dff_B_0U5GZGzw6_2;
	wire w_dff_B_RHe6sdbS3_2;
	wire w_dff_B_qWPlpAAc5_2;
	wire w_dff_B_6z3xrdX69_2;
	wire w_dff_B_zcZ4tKoi5_2;
	wire w_dff_B_pWMBnui65_2;
	wire w_dff_B_4FAhZVik4_2;
	wire w_dff_B_R8zUJDv94_2;
	wire w_dff_B_GpoS2ciP9_2;
	wire w_dff_B_Gx5RMmQk2_2;
	wire w_dff_B_ho6CeItt7_2;
	wire w_dff_B_CBr7vovW7_2;
	wire w_dff_A_2tJH9mlD7_2;
	wire w_dff_A_6HyZwmq06_2;
	wire w_dff_A_LDkkK9UI8_2;
	wire w_dff_A_ocoDvnBD0_2;
	wire w_dff_A_Iz8hZefj9_2;
	wire w_dff_A_GPgtXtqb4_2;
	wire w_dff_A_KydmmE2h0_2;
	wire w_dff_A_hEM6JJns1_2;
	wire w_dff_A_3tgqsPRM3_2;
	wire w_dff_A_Xe41X6qo2_2;
	wire w_dff_A_IbsehqEZ1_2;
	wire w_dff_A_z8dv6Cyc3_2;
	wire w_dff_A_0cc3bsGT0_2;
	wire w_dff_A_nRmQI1pI1_2;
	wire w_dff_A_nuPWCobX3_2;
	wire w_dff_A_ODBhPCbc7_2;
	wire w_dff_A_Ze6XHiJr6_0;
	wire w_dff_A_XKMUUbtb7_0;
	wire w_dff_A_eaEClgUN7_0;
	wire w_dff_A_HSS8BUx25_0;
	wire w_dff_A_vPjYaV1C4_0;
	wire w_dff_A_9nIqZS5z3_0;
	wire w_dff_A_NiUr84898_0;
	wire w_dff_A_jP0WDR4F1_0;
	wire w_dff_A_USwOKz9E2_0;
	wire w_dff_A_3rCqbU0j3_0;
	wire w_dff_A_w5Oe1Zku4_0;
	wire w_dff_A_ijZOQv6z9_0;
	wire w_dff_A_QLuiCQ632_0;
	wire w_dff_A_EQzlzmTc5_1;
	wire w_dff_A_rWTdhc5P9_1;
	wire w_dff_A_HvH6bxXn1_1;
	wire w_dff_A_lMyJxd4G7_1;
	wire w_dff_A_jW4Q9AXx7_1;
	wire w_dff_A_9vBTLN8Z5_1;
	wire w_dff_A_I3nsEFKs9_1;
	wire w_dff_A_OEVyauOl2_1;
	wire w_dff_A_0xYZ7qo33_1;
	wire w_dff_A_QBXP7ueY5_1;
	wire w_dff_A_eQi5s9X70_1;
	jnot g0000(.din(w_G545_0[2]),.dout(G594),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(w_G366_0[1]),.dout(G600),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(G602),.clk(gclk));
	jnot g0005(.din(w_G338_0[1]),.dout(G611),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(G810),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(G848),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(G849),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(G850),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(G851),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(G634),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_1GtAzzyc1_1),.dout(G815),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jcb g0016(.dina(w_dff_B_uqSiIOCB0_0),.dinb(w_n316_0[1]),.dout(G845));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(G847),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jcb g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_));
	jcb g0022(.dina(w_G809_3[1]),.dinb(n320),.dout(G656));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jcb g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330));
	jcb g0030(.dina(n330),.dinb(n327),.dout(G636));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jcb g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336));
	jcb g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(G704));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jcb g0038(.dina(w_G809_2[1]),.dinb(n338),.dout(G820));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_vir5UhkS1_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jcb g0041(.dina(n341),.dinb(w_G809_2[0]),.dout(n342));
	jcb g0042(.dina(w_dff_B_kF86fxm53_0),.dinb(n340),.dout(n343));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(G639),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_iajVVK8S0_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jcb g0046(.dina(n346),.dinb(w_G809_1[2]),.dout(n347));
	jcb g0047(.dina(w_dff_B_80zcCL4t4_0),.dinb(n345),.dout(n348));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(G673),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_uKAsZBfU9_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jcb g0051(.dina(n351),.dinb(w_G809_1[1]),.dout(n352));
	jcb g0052(.dina(w_dff_B_WhznrxG92_0),.dinb(n350),.dout(n353));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(G707),.clk(gclk));
	jand g0054(.dina(w_G2358_0[2]),.dinb(G80),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_n326_0[2]),.dinb(w_dff_B_i1OZVmBg6_1),.dout(n356),.clk(gclk));
	jcb g0056(.dina(n356),.dinb(w_G809_1[0]),.dout(n357));
	jcb g0057(.dina(n357),.dinb(w_dff_B_6oA78GKR0_1),.dout(n358));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(G715),.clk(gclk));
	jand g0059(.dina(w_G3552_0[1]),.dinb(w_G514_2[1]),.dout(n360),.clk(gclk));
	jnot g0060(.din(w_G514_2[0]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G3546_5[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(n362),.dinb(w_n361_0[1]),.dout(n363),.clk(gclk));
	jcb g0063(.dina(n363),.dinb(w_dff_B_de19BWZc6_1),.dout(n364));
	jnot g0064(.din(n364),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G251_5[1]),.dout(n366),.clk(gclk));
	jnot g0066(.din(w_G361_1[1]),.dout(n367),.clk(gclk));
	jand g0067(.dina(n367),.dinb(w_n366_1[2]),.dout(n368),.clk(gclk));
	jnot g0068(.din(w_G248_5[2]),.dout(n369),.clk(gclk));
	jand g0069(.dina(w_G361_1[0]),.dinb(w_n369_1[2]),.dout(n370),.clk(gclk));
	jcb g0070(.dina(n370),.dinb(n368),.dout(n371));
	jnot g0071(.din(w_n371_0[1]),.dout(n372),.clk(gclk));
	jand g0072(.dina(w_n372_0[1]),.dinb(w_n365_0[1]),.dout(n373),.clk(gclk));
	jnot g0073(.din(w_G351_2[2]),.dout(n374),.clk(gclk));
	jnot g0074(.din(G3550),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_n375_4[2]),.dinb(w_n374_1[1]),.dout(n376),.clk(gclk));
	jnot g0076(.din(w_G534_2[1]),.dout(n377),.clk(gclk));
	jnot g0077(.din(w_G3552_0[0]),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n378_4[2]),.dinb(w_G351_2[1]),.dout(n379),.clk(gclk));
	jcb g0079(.dina(n379),.dinb(w_n377_1[1]),.dout(n380));
	jcb g0080(.dina(n380),.dinb(n376),.dout(n381));
	jand g0081(.dina(w_G3546_5[0]),.dinb(w_G351_2[0]),.dout(n382),.clk(gclk));
	jand g0082(.dina(w_G3548_4[2]),.dinb(w_n374_1[0]),.dout(n383),.clk(gclk));
	jcb g0083(.dina(n383),.dinb(w_dff_B_nek1dyeV9_1),.dout(n384));
	jcb g0084(.dina(n384),.dinb(w_G534_2[0]),.dout(n385));
	jand g0085(.dina(n385),.dinb(n381),.dout(n386),.clk(gclk));
	jnot g0086(.din(w_G341_2[2]),.dout(n387),.clk(gclk));
	jand g0087(.dina(w_n375_4[1]),.dinb(w_n387_1[1]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G523_1[2]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n378_4[1]),.dinb(w_G341_2[1]),.dout(n390),.clk(gclk));
	jcb g0090(.dina(n390),.dinb(w_n389_1[1]),.dout(n391));
	jcb g0091(.dina(n391),.dinb(n388),.dout(n392));
	jand g0092(.dina(w_G3546_4[2]),.dinb(w_G341_2[0]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3548_4[1]),.dinb(w_n387_1[0]),.dout(n394),.clk(gclk));
	jcb g0094(.dina(n394),.dinb(w_dff_B_SWNB9SoI5_1),.dout(n395));
	jcb g0095(.dina(n395),.dinb(w_G523_1[1]),.dout(n396));
	jand g0096(.dina(n396),.dinb(n392),.dout(n397),.clk(gclk));
	jand g0097(.dina(w_n397_0[1]),.dinb(w_n386_0[1]),.dout(n398),.clk(gclk));
	jand g0098(.dina(n398),.dinb(n373),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G316_1[1]),.dinb(w_G248_5[1]),.dout(n400),.clk(gclk));
	jnot g0100(.din(w_G490_1[1]),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G316_1[0]),.dout(n402),.clk(gclk));
	jand g0102(.dina(w_n402_0[2]),.dinb(w_G251_5[0]),.dout(n403),.clk(gclk));
	jcb g0103(.dina(n403),.dinb(w_n401_0[1]),.dout(n404));
	jcb g0104(.dina(n404),.dinb(w_dff_B_pOQmJj3U1_1),.dout(n405));
	jnot g0105(.din(w_G254_1[1]),.dout(n406),.clk(gclk));
	jand g0106(.dina(w_n402_0[1]),.dinb(w_n406_5[1]),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_G242_1[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_G316_0[2]),.dinb(w_n408_5[2]),.dout(n409),.clk(gclk));
	jcb g0109(.dina(n409),.dinb(n407),.dout(n410));
	jcb g0110(.dina(n410),.dinb(w_G490_1[0]),.dout(n411));
	jand g0111(.dina(n411),.dinb(n405),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G308_1[2]),.dinb(w_G248_5[0]),.dout(n413),.clk(gclk));
	jnot g0113(.din(w_G479_0[2]),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_G308_1[1]),.dout(n415),.clk(gclk));
	jand g0115(.dina(w_n415_0[1]),.dinb(w_G251_4[2]),.dout(n416),.clk(gclk));
	jcb g0116(.dina(n416),.dinb(w_n414_0[1]),.dout(n417));
	jcb g0117(.dina(n417),.dinb(w_dff_B_iv4zvYdQ6_1),.dout(n418));
	jand g0118(.dina(w_n415_0[0]),.dinb(w_n406_5[0]),.dout(n419),.clk(gclk));
	jand g0119(.dina(w_G308_1[0]),.dinb(w_n408_5[1]),.dout(n420),.clk(gclk));
	jcb g0120(.dina(n420),.dinb(n419),.dout(n421));
	jcb g0121(.dina(n421),.dinb(w_G479_0[1]),.dout(n422));
	jand g0122(.dina(n422),.dinb(n418),.dout(n423),.clk(gclk));
	jand g0123(.dina(w_n423_0[2]),.dinb(w_n412_0[2]),.dout(n424),.clk(gclk));
	jnot g0124(.din(w_G293_0[2]),.dout(n425),.clk(gclk));
	jand g0125(.dina(w_n425_0[2]),.dinb(w_n406_4[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_G293_0[1]),.dinb(w_n408_5[0]),.dout(n427),.clk(gclk));
	jcb g0127(.dina(n427),.dinb(n426),.dout(n428));
	jnot g0128(.din(w_G302_0[2]),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_n429_0[1]),.dinb(w_n366_1[1]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G302_0[1]),.dinb(w_n369_1[1]),.dout(n431),.clk(gclk));
	jcb g0131(.dina(n431),.dinb(n430),.dout(n432));
	jnot g0132(.din(n432),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_n433_0[2]),.dinb(w_n428_1[1]),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G324_1[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n375_4[0]),.dinb(w_n435_2[1]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G503_2[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n378_4[0]),.dinb(w_G324_1[1]),.dout(n438),.clk(gclk));
	jcb g0138(.dina(n438),.dinb(w_n437_0[1]),.dout(n439));
	jcb g0139(.dina(n439),.dinb(n436),.dout(n440));
	jand g0140(.dina(w_G3546_4[1]),.dinb(w_G324_1[0]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3548_4[0]),.dinb(w_n435_2[0]),.dout(n442),.clk(gclk));
	jcb g0142(.dina(n442),.dinb(w_dff_B_F9EoP2rl4_1),.dout(n443));
	jcb g0143(.dina(n443),.dinb(w_G503_2[0]),.dout(n444));
	jand g0144(.dina(n444),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(n434),.dout(n446),.clk(gclk));
	jand g0146(.dina(n446),.dinb(w_dff_B_n6bJKEiU7_1),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(w_dff_B_4OnXHcKF9_1),.dout(G598),.clk(gclk));
	jnot g0148(.din(w_G210_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n375_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G457_1[2]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n378_3[2]),.dinb(w_G210_2[0]),.dout(n452),.clk(gclk));
	jcb g0152(.dina(n452),.dinb(w_n451_0[2]),.dout(n453));
	jcb g0153(.dina(n453),.dinb(n450),.dout(n454));
	jand g0154(.dina(w_G3546_4[0]),.dinb(w_G210_1[2]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n456),.clk(gclk));
	jcb g0156(.dina(n456),.dinb(w_dff_B_ls9Jbc5m9_1),.dout(n457));
	jcb g0157(.dina(n457),.dinb(w_G457_1[1]),.dout(n458));
	jand g0158(.dina(n458),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n375_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n378_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jcb g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464));
	jcb g0164(.dina(n464),.dinb(n461),.dout(n465));
	jand g0165(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n467),.clk(gclk));
	jcb g0167(.dina(n467),.dinb(w_dff_B_1JyXEtsm3_1),.dout(n468));
	jcb g0168(.dina(n468),.dinb(w_G435_1[1]),.dout(n469));
	jand g0169(.dina(n469),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G273_2[1]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n375_3[0]),.dinb(w_n471_1[2]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G411_2[1]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n378_3[0]),.dinb(w_G273_2[0]),.dout(n474),.clk(gclk));
	jcb g0174(.dina(n474),.dinb(w_n473_1[1]),.dout(n475));
	jcb g0175(.dina(n475),.dinb(n472),.dout(n476));
	jand g0176(.dina(w_G3546_3[1]),.dinb(w_G273_1[2]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3548_3[0]),.dinb(w_n471_1[1]),.dout(n478),.clk(gclk));
	jcb g0178(.dina(n478),.dinb(w_dff_B_aMvWkg9f4_1),.dout(n479));
	jcb g0179(.dina(n479),.dinb(w_G411_2[0]),.dout(n480));
	jand g0180(.dina(n480),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jnot g0182(.din(w_G265_1[2]),.dout(n483),.clk(gclk));
	jand g0183(.dina(w_n375_2[2]),.dinb(w_n483_2[1]),.dout(n484),.clk(gclk));
	jnot g0184(.din(w_G400_1[2]),.dout(n485),.clk(gclk));
	jand g0185(.dina(w_n378_2[2]),.dinb(w_G265_1[1]),.dout(n486),.clk(gclk));
	jcb g0186(.dina(n486),.dinb(w_n485_1[1]),.dout(n487));
	jcb g0187(.dina(n487),.dinb(n484),.dout(n488));
	jand g0188(.dina(w_G3546_3[0]),.dinb(w_G265_1[0]),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n483_2[0]),.dout(n490),.clk(gclk));
	jcb g0190(.dina(n490),.dinb(w_dff_B_Tgn2H91z5_1),.dout(n491));
	jcb g0191(.dina(n491),.dinb(w_G400_1[1]),.dout(n492));
	jand g0192(.dina(n492),.dinb(n488),.dout(n493),.clk(gclk));
	jnot g0193(.din(w_G226_2[1]),.dout(n494),.clk(gclk));
	jand g0194(.dina(w_n375_2[1]),.dinb(w_n494_1[2]),.dout(n495),.clk(gclk));
	jnot g0195(.din(w_G422_1[1]),.dout(n496),.clk(gclk));
	jand g0196(.dina(w_n378_2[1]),.dinb(w_G226_2[0]),.dout(n497),.clk(gclk));
	jcb g0197(.dina(n497),.dinb(w_n496_1[1]),.dout(n498));
	jcb g0198(.dina(n498),.dinb(n495),.dout(n499));
	jand g0199(.dina(w_G3546_2[2]),.dinb(w_G226_1[2]),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n494_1[1]),.dout(n501),.clk(gclk));
	jcb g0201(.dina(n501),.dinb(w_dff_B_uRSWtzdc4_1),.dout(n502));
	jcb g0202(.dina(n502),.dinb(w_G422_1[0]),.dout(n503));
	jand g0203(.dina(n503),.dinb(n499),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_n504_0[1]),.dinb(w_n493_0[1]),.dout(n505),.clk(gclk));
	jand g0205(.dina(n505),.dinb(n482),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[1]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n375_2[0]),.dinb(w_n507_1[2]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n378_2[0]),.dinb(w_G218_2[0]),.dout(n510),.clk(gclk));
	jcb g0210(.dina(n510),.dinb(w_n509_0[2]),.dout(n511));
	jcb g0211(.dina(n511),.dinb(n508),.dout(n512));
	jand g0212(.dina(w_G3546_2[1]),.dinb(w_G218_1[2]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3548_2[0]),.dinb(w_n507_1[1]),.dout(n514),.clk(gclk));
	jcb g0214(.dina(n514),.dinb(w_dff_B_cUsp9VPF8_1),.dout(n515));
	jcb g0215(.dina(n515),.dinb(w_G468_1[1]),.dout(n516));
	jand g0216(.dina(n516),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G257_2[1]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_n375_1[2]),.dinb(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G389_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_n378_1[2]),.dinb(w_G257_2[0]),.dout(n521),.clk(gclk));
	jcb g0221(.dina(n521),.dinb(w_n520_0[2]),.dout(n522));
	jcb g0222(.dina(n522),.dinb(n519),.dout(n523));
	jand g0223(.dina(w_G3546_2[0]),.dinb(w_G257_1[2]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_G3548_1[2]),.dinb(w_n518_1[1]),.dout(n525),.clk(gclk));
	jcb g0225(.dina(n525),.dinb(w_dff_B_ns3mmr1l6_1),.dout(n526));
	jcb g0226(.dina(n526),.dinb(w_G389_1[1]),.dout(n527));
	jand g0227(.dina(n527),.dinb(n523),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[1]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G281_2[1]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n375_1[1]),.dinb(w_n530_1[2]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G374_1[2]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n378_1[1]),.dinb(w_G281_2[0]),.dout(n533),.clk(gclk));
	jcb g0233(.dina(n533),.dinb(w_n532_1[1]),.dout(n534));
	jcb g0234(.dina(n534),.dinb(n531),.dout(n535));
	jand g0235(.dina(w_G3546_1[2]),.dinb(w_G281_1[2]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3548_1[1]),.dinb(w_n530_1[1]),.dout(n537),.clk(gclk));
	jcb g0237(.dina(n537),.dinb(w_dff_B_CQjF9HTI5_1),.dout(n538));
	jcb g0238(.dina(n538),.dinb(w_G374_1[1]),.dout(n539));
	jand g0239(.dina(n539),.dinb(n535),.dout(n540),.clk(gclk));
	jand g0240(.dina(w_G248_4[2]),.dinb(w_G206_1[2]),.dout(n541),.clk(gclk));
	jnot g0241(.din(w_G446_1[2]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G206_1[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_G251_4[1]),.dinb(w_n543_0[1]),.dout(n544),.clk(gclk));
	jcb g0244(.dina(n544),.dinb(w_dff_B_2EtDnD859_1),.dout(n545));
	jcb g0245(.dina(n545),.dinb(w_dff_B_OQMF5acT7_1),.dout(n546));
	jand g0246(.dina(w_n406_4[1]),.dinb(w_n543_0[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_n408_4[2]),.dinb(w_G206_1[0]),.dout(n548),.clk(gclk));
	jcb g0248(.dina(n548),.dinb(n547),.dout(n549));
	jcb g0249(.dina(n549),.dinb(w_G446_1[1]),.dout(n550));
	jand g0250(.dina(n550),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[2]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(n506),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_n459_0[1]),.dout(G610),.clk(gclk));
	jnot g0255(.din(w_G335_0[2]),.dout(n556),.clk(gclk));
	jand g0256(.dina(w_n556_8[1]),.dinb(w_n530_1[0]),.dout(n557),.clk(gclk));
	jnot g0257(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jcb g0258(.dina(w_n556_8[0]),.dinb(w_dff_B_N5KTHUmM9_1),.dout(n559));
	jand g0259(.dina(w_n559_0[1]),.dinb(n558),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_0[2]),.dinb(w_G374_1[0]),.dout(n561),.clk(gclk));
	jand g0261(.dina(w_n556_7[2]),.dinb(w_n471_1[0]),.dout(n562),.clk(gclk));
	jnot g0262(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jcb g0263(.dina(w_n556_7[1]),.dinb(w_dff_B_H8GXBcUn2_1),.dout(n564));
	jand g0264(.dina(w_n564_0[1]),.dinb(n563),.dout(n565),.clk(gclk));
	jxor g0265(.dina(w_n565_0[2]),.dinb(w_G411_1[2]),.dout(n566),.clk(gclk));
	jand g0266(.dina(w_n566_0[2]),.dinb(w_n561_1[1]),.dout(n567),.clk(gclk));
	jnot g0267(.din(w_n567_0[2]),.dout(n568),.clk(gclk));
	jand g0268(.dina(w_n556_7[0]),.dinb(w_n483_1[2]),.dout(n569),.clk(gclk));
	jnot g0269(.din(w_n569_0[1]),.dout(n570),.clk(gclk));
	jcb g0270(.dina(w_n556_6[2]),.dinb(w_dff_B_xvI34cRN7_1),.dout(n571));
	jand g0271(.dina(w_n571_0[1]),.dinb(n570),.dout(n572),.clk(gclk));
	jxor g0272(.dina(w_n572_0[2]),.dinb(w_G400_1[0]),.dout(n573),.clk(gclk));
	jnot g0273(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jand g0274(.dina(w_n556_6[1]),.dinb(w_n518_1[0]),.dout(n575),.clk(gclk));
	jnot g0275(.din(n575),.dout(n576),.clk(gclk));
	jcb g0276(.dina(w_n556_6[0]),.dinb(w_dff_B_Z0FhR6SO8_1),.dout(n577));
	jand g0277(.dina(w_dff_B_RJyCFA7L9_0),.dinb(n576),.dout(n578),.clk(gclk));
	jxor g0278(.dina(w_n578_1[1]),.dinb(w_n520_0[1]),.dout(n579),.clk(gclk));
	jcb g0279(.dina(w_n579_1[1]),.dinb(w_n574_0[2]),.dout(n580));
	jcb g0280(.dina(w_dff_B_weWeD51m0_0),.dinb(n568),.dout(n581));
	jnot g0281(.din(w_n581_0[1]),.dout(n582),.clk(gclk));
	jand g0282(.dina(w_n556_5[2]),.dinb(w_n460_1[0]),.dout(n583),.clk(gclk));
	jnot g0283(.din(n583),.dout(n584),.clk(gclk));
	jcb g0284(.dina(w_n556_5[1]),.dinb(w_dff_B_s1Lg2lHD0_1),.dout(n585));
	jand g0285(.dina(w_dff_B_xbfNDrb60_0),.dinb(n584),.dout(n586),.clk(gclk));
	jxor g0286(.dina(w_n586_1[1]),.dinb(w_G435_1[0]),.dout(n587),.clk(gclk));
	jand g0287(.dina(w_n587_0[1]),.dinb(n582),.dout(n588),.clk(gclk));
	jcb g0288(.dina(w_G335_0[1]),.dinb(w_G206_0[2]),.dout(n589));
	jcb g0289(.dina(w_n556_5[0]),.dinb(w_dff_B_VWEEJY1S1_1),.dout(n590));
	jand g0290(.dina(n590),.dinb(w_dff_B_YBkNYZOG6_1),.dout(n591),.clk(gclk));
	jxor g0291(.dina(w_n591_1[1]),.dinb(w_G446_1[0]),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_4[2]),.dinb(w_n494_1[0]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jcb g0294(.dina(w_n556_4[1]),.dinb(w_dff_B_JUCzJ7sa9_1),.dout(n595));
	jand g0295(.dina(w_dff_B_vi8uLsP27_0),.dinb(n594),.dout(n596),.clk(gclk));
	jxor g0296(.dina(w_n596_1[1]),.dinb(w_n496_1[0]),.dout(n597),.clk(gclk));
	jand g0297(.dina(w_n556_4[0]),.dinb(w_n507_1[0]),.dout(n598),.clk(gclk));
	jnot g0298(.din(n598),.dout(n599),.clk(gclk));
	jcb g0299(.dina(w_n556_3[2]),.dinb(w_dff_B_Bfz9YGEj0_1),.dout(n600));
	jand g0300(.dina(w_dff_B_Rvnwe1wD7_0),.dinb(n599),.dout(n601),.clk(gclk));
	jxor g0301(.dina(w_n601_1[1]),.dinb(w_n509_0[1]),.dout(n602),.clk(gclk));
	jcb g0302(.dina(w_n602_0[2]),.dinb(w_n597_0[2]),.dout(n603));
	jand g0303(.dina(w_n556_3[1]),.dinb(w_n449_1[0]),.dout(n604),.clk(gclk));
	jnot g0304(.din(n604),.dout(n605),.clk(gclk));
	jcb g0305(.dina(w_n556_3[0]),.dinb(w_dff_B_6l8Es9rU3_1),.dout(n606));
	jand g0306(.dina(w_dff_B_sb7ax8Z62_0),.dinb(n605),.dout(n607),.clk(gclk));
	jxor g0307(.dina(w_n607_1[1]),.dinb(w_n451_0[1]),.dout(n608),.clk(gclk));
	jcb g0308(.dina(w_n608_0[2]),.dinb(w_n603_0[1]),.dout(n609));
	jnot g0309(.din(w_n609_0[2]),.dout(n610),.clk(gclk));
	jand g0310(.dina(n610),.dinb(w_n592_0[2]),.dout(n611),.clk(gclk));
	jand g0311(.dina(w_n611_0[2]),.dinb(w_n588_1[1]),.dout(G588),.clk(gclk));
	jnot g0312(.din(w_G332_3[2]),.dout(n613),.clk(gclk));
	jand g0313(.dina(w_n613_5[2]),.dinb(w_n435_1[2]),.dout(n614),.clk(gclk));
	jnot g0314(.din(n614),.dout(n615),.clk(gclk));
	jcb g0315(.dina(w_n613_5[1]),.dinb(w_G331_0[1]),.dout(n616));
	jand g0316(.dina(w_dff_B_dCZwKOI10_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_G503_1[2]),.dout(n618),.clk(gclk));
	jcb g0318(.dina(w_G338_0[0]),.dinb(w_n613_5[0]),.dout(n619));
	jxor g0319(.dina(w_n619_1[2]),.dinb(w_G514_1[2]),.dout(n620),.clk(gclk));
	jcb g0320(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n621));
	jcb g0321(.dina(w_G348_0[0]),.dinb(w_n613_4[2]),.dout(n622));
	jand g0322(.dina(n622),.dinb(w_n621_0[1]),.dout(n623),.clk(gclk));
	jxor g0323(.dina(w_n623_0[1]),.dinb(w_G523_1[0]),.dout(n624),.clk(gclk));
	jcb g0324(.dina(w_G351_1[2]),.dinb(w_G332_3[0]),.dout(n625));
	jcb g0325(.dina(w_G358_0[0]),.dinb(w_n613_4[1]),.dout(n626));
	jand g0326(.dina(n626),.dinb(w_n625_0[1]),.dout(n627),.clk(gclk));
	jcb g0327(.dina(w_n627_1[1]),.dinb(w_G534_1[2]),.dout(n628));
	jnot g0328(.din(w_n625_0[0]),.dout(n629),.clk(gclk));
	jand g0329(.dina(w_G612_0),.dinb(w_G332_2[2]),.dout(n630),.clk(gclk));
	jcb g0330(.dina(n630),.dinb(w_dff_B_aWKtNM9w2_1),.dout(n631));
	jcb g0331(.dina(w_n631_0[1]),.dinb(w_n377_1[0]),.dout(n632));
	jcb g0332(.dina(w_G361_0[2]),.dinb(w_G332_2[1]),.dout(n633));
	jcb g0333(.dina(w_G366_0[0]),.dinb(w_n613_4[0]),.dout(n634));
	jand g0334(.dina(n634),.dinb(w_dff_B_of19NiuT7_1),.dout(n635),.clk(gclk));
	jnot g0335(.din(w_n635_1[1]),.dout(n636),.clk(gclk));
	jand g0336(.dina(w_n636_0[2]),.dinb(w_n632_0[1]),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n637_0[2]),.dinb(w_n628_0[2]),.dout(n638),.clk(gclk));
	jand g0338(.dina(w_n638_0[1]),.dinb(w_n624_0[2]),.dout(n639),.clk(gclk));
	jand g0339(.dina(w_n639_0[2]),.dinb(w_n620_1[1]),.dout(n640),.clk(gclk));
	jand g0340(.dina(w_n640_0[1]),.dinb(w_n618_0[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n613_3[2]),.dinb(w_n425_0[1]),.dout(n642),.clk(gclk));
	jand g0342(.dina(w_G332_2[0]),.dinb(w_G593_0),.dout(n643),.clk(gclk));
	jcb g0343(.dina(n643),.dinb(n642),.dout(n644));
	jand g0344(.dina(w_n613_3[1]),.dinb(w_n429_0[0]),.dout(n645),.clk(gclk));
	jnot g0345(.din(n645),.dout(n646),.clk(gclk));
	jcb g0346(.dina(w_n613_3[0]),.dinb(w_dff_B_fshypG5j3_1),.dout(n647));
	jand g0347(.dina(w_dff_B_r1zOMHRi2_0),.dinb(n646),.dout(n648),.clk(gclk));
	jnot g0348(.din(w_n648_1[1]),.dout(n649),.clk(gclk));
	jand g0349(.dina(w_n649_0[1]),.dinb(w_n644_0[2]),.dout(n650),.clk(gclk));
	jcb g0350(.dina(w_G332_1[2]),.dinb(w_G308_0[2]),.dout(n651));
	jcb g0351(.dina(w_n613_2[2]),.dinb(w_dff_B_McNbNlnj5_1),.dout(n652));
	jand g0352(.dina(n652),.dinb(w_dff_B_iO5cs4jZ7_1),.dout(n653),.clk(gclk));
	jxor g0353(.dina(w_n653_0[2]),.dinb(w_G479_0[0]),.dout(n654),.clk(gclk));
	jand g0354(.dina(w_n613_2[1]),.dinb(w_n402_0[0]),.dout(n655),.clk(gclk));
	jnot g0355(.din(n655),.dout(n656),.clk(gclk));
	jcb g0356(.dina(w_n613_2[0]),.dinb(w_dff_B_aVgFD1dL9_1),.dout(n657));
	jand g0357(.dina(w_dff_B_OF3KwrDd9_0),.dinb(n656),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_n658_1[1]),.dinb(w_G490_0[2]),.dout(n659),.clk(gclk));
	jand g0359(.dina(w_n659_0[1]),.dinb(w_n654_2[2]),.dout(n660),.clk(gclk));
	jand g0360(.dina(w_n660_1[1]),.dinb(w_n650_0[1]),.dout(n661),.clk(gclk));
	jand g0361(.dina(w_n661_0[1]),.dinb(w_n641_1[2]),.dout(G615),.clk(gclk));
	jxor g0362(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G302_0[0]),.dinb(w_n425_0[0]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(w_dff_B_HrWB5H7K4_1),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G369_0[1]),.dinb(w_G361_0[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(n666),.dinb(w_n435_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_dff_B_8m802Xw05_0),.dinb(n667),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n665),.dout(n670),.clk(gclk));
	jnot g0370(.din(w_n670_0[1]),.dout(G1002),.clk(gclk));
	jxor g0371(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n672),.clk(gclk));
	jxor g0372(.dina(w_G273_1[1]),.dinb(w_n483_1[1]),.dout(n673),.clk(gclk));
	jxor g0373(.dina(n673),.dinb(w_dff_B_VDU12DIm5_1),.dout(n674),.clk(gclk));
	jxor g0374(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n675),.clk(gclk));
	jxor g0375(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n676),.clk(gclk));
	jxor g0376(.dina(n676),.dinb(n675),.dout(n677),.clk(gclk));
	jxor g0377(.dina(w_G210_1[1]),.dinb(w_G206_0[1]),.dout(n678),.clk(gclk));
	jxor g0378(.dina(w_dff_B_UkrEuE9s7_0),.dinb(n677),.dout(n679),.clk(gclk));
	jxor g0379(.dina(n679),.dinb(n674),.dout(n680),.clk(gclk));
	jnot g0380(.din(w_n680_0[1]),.dout(G1004),.clk(gclk));
	jand g0381(.dina(w_n586_1[0]),.dinb(w_G435_0[2]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_n586_0[2]),.dout(n683),.clk(gclk));
	jand g0383(.dina(n683),.dinb(w_n462_0[1]),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n684_0[1]),.dout(n685),.clk(gclk));
	jand g0385(.dina(w_n578_1[0]),.dinb(w_G389_1[0]),.dout(n686),.clk(gclk));
	jcb g0386(.dina(w_n578_0[2]),.dinb(w_G389_0[2]),.dout(n687));
	jnot g0387(.din(w_n571_0[0]),.dout(n688),.clk(gclk));
	jcb g0388(.dina(n688),.dinb(w_n569_0[0]),.dout(n689));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n485_1[0]),.dout(n690),.clk(gclk));
	jnot g0390(.din(w_n690_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n560_0[1]),.dinb(w_G374_0[2]),.dout(n692),.clk(gclk));
	jcb g0392(.dina(w_n565_0[1]),.dinb(w_G411_1[1]),.dout(n693));
	jand g0393(.dina(w_dff_B_WqTalyok5_0),.dinb(w_n692_0[1]),.dout(n694),.clk(gclk));
	jand g0394(.dina(w_n565_0[0]),.dinb(w_G411_1[0]),.dout(n695),.clk(gclk));
	jand g0395(.dina(w_n572_0[1]),.dinb(w_G400_0[2]),.dout(n696),.clk(gclk));
	jcb g0396(.dina(n696),.dinb(w_n695_0[2]),.dout(n697));
	jcb g0397(.dina(w_dff_B_dEl6L4no0_0),.dinb(w_n694_0[2]),.dout(n698));
	jand g0398(.dina(n698),.dinb(w_dff_B_Rd6uJHVp0_1),.dout(n699),.clk(gclk));
	jand g0399(.dina(w_n699_0[2]),.dinb(w_n687_0[1]),.dout(n700),.clk(gclk));
	jcb g0400(.dina(n700),.dinb(w_n686_0[1]),.dout(n701));
	jand g0401(.dina(w_n701_0[1]),.dinb(w_n685_0[1]),.dout(n702),.clk(gclk));
	jcb g0402(.dina(n702),.dinb(w_n682_0[2]),.dout(n703));
	jand g0403(.dina(w_n703_0[2]),.dinb(w_n611_0[1]),.dout(n704),.clk(gclk));
	jand g0404(.dina(w_n591_1[0]),.dinb(w_G446_0[2]),.dout(n705),.clk(gclk));
	jcb g0405(.dina(w_n591_0[2]),.dinb(w_G446_0[1]),.dout(n706));
	jand g0406(.dina(w_n607_1[0]),.dinb(w_G457_1[0]),.dout(n707),.clk(gclk));
	jcb g0407(.dina(w_n607_0[2]),.dinb(w_G457_0[2]),.dout(n708));
	jand g0408(.dina(w_n601_1[0]),.dinb(w_G468_1[0]),.dout(n709),.clk(gclk));
	jand g0409(.dina(w_n596_1[0]),.dinb(w_G422_0[2]),.dout(n710),.clk(gclk));
	jcb g0410(.dina(w_n601_0[2]),.dinb(w_G468_0[2]),.dout(n711));
	jand g0411(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jcb g0412(.dina(n712),.dinb(w_n709_0[1]),.dout(n713));
	jand g0413(.dina(w_n713_0[2]),.dinb(w_dff_B_GCIUjCEb3_1),.dout(n714),.clk(gclk));
	jcb g0414(.dina(n714),.dinb(w_dff_B_LFGWI0nG2_1),.dout(n715));
	jand g0415(.dina(w_n715_0[2]),.dinb(w_dff_B_9kpzX39X0_1),.dout(n716),.clk(gclk));
	jcb g0416(.dina(n716),.dinb(w_dff_B_F2MQMNNB6_1),.dout(n717));
	jcb g0417(.dina(w_n717_0[1]),.dinb(w_n704_0[1]),.dout(G591));
	jand g0418(.dina(w_n617_1[0]),.dinb(w_G503_1[1]),.dout(n719),.clk(gclk));
	jcb g0419(.dina(w_n617_0[2]),.dinb(w_G503_1[0]),.dout(n720));
	jcb g0420(.dina(w_n619_1[1]),.dinb(w_G514_1[1]),.dout(n721));
	jand g0421(.dina(w_n619_1[0]),.dinb(w_G514_1[0]),.dout(n722),.clk(gclk));
	jnot g0422(.din(w_n621_0[0]),.dout(n723),.clk(gclk));
	jand g0423(.dina(w_G599_0),.dinb(w_G332_1[1]),.dout(n724),.clk(gclk));
	jcb g0424(.dina(n724),.dinb(w_dff_B_Y6uJcumH7_1),.dout(n725));
	jand g0425(.dina(w_n725_0[2]),.dinb(w_n389_1[0]),.dout(n726),.clk(gclk));
	jnot g0426(.din(w_n726_0[1]),.dout(n727),.clk(gclk));
	jand g0427(.dina(w_n635_1[0]),.dinb(w_n628_0[1]),.dout(n728),.clk(gclk));
	jand g0428(.dina(w_n623_0[0]),.dinb(w_G523_0[2]),.dout(n729),.clk(gclk));
	jand g0429(.dina(w_n627_1[0]),.dinb(w_G534_1[1]),.dout(n730),.clk(gclk));
	jcb g0430(.dina(n730),.dinb(n729),.dout(n731));
	jcb g0431(.dina(n731),.dinb(w_n728_0[1]),.dout(n732));
	jand g0432(.dina(w_dff_B_tS6mCmRe0_0),.dinb(n727),.dout(n733),.clk(gclk));
	jcb g0433(.dina(w_n733_0[2]),.dinb(w_n722_0[1]),.dout(n734));
	jand g0434(.dina(n734),.dinb(w_n721_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[2]),.dinb(w_n720_0[1]),.dout(n736),.clk(gclk));
	jcb g0436(.dina(n736),.dinb(w_n719_0[1]),.dout(n737));
	jand g0437(.dina(w_n737_1[1]),.dinb(w_n660_1[0]),.dout(n738),.clk(gclk));
	jnot g0438(.din(w_n650_0[0]),.dout(n739),.clk(gclk));
	jnot g0439(.din(w_n653_0[1]),.dout(n740),.clk(gclk));
	jcb g0440(.dina(n740),.dinb(w_n414_0[0]),.dout(n741));
	jand g0441(.dina(w_n658_1[0]),.dinb(w_G490_0[1]),.dout(n742),.clk(gclk));
	jand g0442(.dina(w_n742_0[2]),.dinb(w_n654_2[1]),.dout(n743),.clk(gclk));
	jnot g0443(.din(n743),.dout(n744),.clk(gclk));
	jand g0444(.dina(n744),.dinb(w_dff_B_hbgrprrW0_1),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_n745_0[1]),.dout(n746),.clk(gclk));
	jcb g0446(.dina(w_n746_0[2]),.dinb(w_dff_B_QS51zgDE7_1),.dout(n747));
	jcb g0447(.dina(w_n747_0[1]),.dinb(w_n738_0[1]),.dout(G618));
	jnot g0448(.din(w_G4091_6[1]),.dout(n749),.clk(gclk));
	jand g0449(.dina(w_G4092_9[2]),.dinb(w_n749_13[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n750_8[2]),.dinb(w_dff_B_RntSM2gG0_1),.dout(n751),.clk(gclk));
	jnot g0451(.din(n751),.dout(n752),.clk(gclk));
	jnot g0452(.din(w_G54_0[2]),.dout(n753),.clk(gclk));
	jxor g0453(.dina(w_n635_0[2]),.dinb(w_n753_1[1]),.dout(n754),.clk(gclk));
	jnot g0454(.din(n754),.dout(n755),.clk(gclk));
	jand g0455(.dina(w_n755_0[1]),.dinb(w_G4091_6[0]),.dout(n756),.clk(gclk));
	jand g0456(.dina(w_n372_0[0]),.dinb(w_n749_13[0]),.dout(n757),.clk(gclk));
	jcb g0457(.dina(n757),.dinb(w_G4092_9[1]),.dout(n758));
	jcb g0458(.dina(w_dff_B_uoBLLF5g3_0),.dinb(n756),.dout(n759));
	jand g0459(.dina(n759),.dinb(w_dff_B_ttqqGnET9_1),.dout(G822_fa_),.clk(gclk));
	jand g0460(.dina(w_n750_8[1]),.dinb(w_dff_B_EDicO3ac1_1),.dout(n761),.clk(gclk));
	jnot g0461(.din(n761),.dout(n762),.clk(gclk));
	jxor g0462(.dina(w_n627_0[2]),.dinb(w_G534_1[0]),.dout(n763),.clk(gclk));
	jnot g0463(.din(w_n763_0[2]),.dout(n764),.clk(gclk));
	jand g0464(.dina(n764),.dinb(w_n635_0[1]),.dout(n765),.clk(gclk));
	jcb g0465(.dina(n765),.dinb(w_n638_0[0]),.dout(n766));
	jnot g0466(.din(n766),.dout(n767),.clk(gclk));
	jand g0467(.dina(w_n767_0[1]),.dinb(w_n753_1[0]),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_n763_0[1]),.dinb(w_G54_0[1]),.dout(n769),.clk(gclk));
	jcb g0469(.dina(w_dff_B_bvUdY8NE0_0),.dinb(n768),.dout(n770));
	jand g0470(.dina(n770),.dinb(w_G4091_5[2]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n386_0[0]),.dinb(w_n749_12[2]),.dout(n772),.clk(gclk));
	jcb g0472(.dina(n772),.dinb(w_G4092_9[0]),.dout(n773));
	jcb g0473(.dina(w_dff_B_xvh3OphK0_0),.dinb(n771),.dout(n774));
	jand g0474(.dina(n774),.dinb(w_dff_B_WKaXesSI6_1),.dout(G838_fa_),.clk(gclk));
	jand g0475(.dina(w_n750_8[0]),.dinb(w_dff_B_tsE0BllG0_1),.dout(n776),.clk(gclk));
	jnot g0476(.din(n776),.dout(n777),.clk(gclk));
	jxor g0477(.dina(w_n561_1[0]),.dinb(w_G4_0[2]),.dout(n778),.clk(gclk));
	jnot g0478(.din(n778),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n779_0[1]),.dinb(w_G4091_5[1]),.dout(n780),.clk(gclk));
	jand g0480(.dina(w_n540_0[0]),.dinb(w_n749_12[1]),.dout(n781),.clk(gclk));
	jcb g0481(.dina(n781),.dinb(w_G4092_8[2]),.dout(n782));
	jcb g0482(.dina(w_dff_B_QMQVtFwl1_0),.dinb(n780),.dout(n783));
	jand g0483(.dina(n783),.dinb(w_dff_B_jgWblR193_1),.dout(G861_fa_),.clk(gclk));
	jand g0484(.dina(w_n641_1[1]),.dinb(w_G54_0[0]),.dout(n785),.clk(gclk));
	jcb g0485(.dina(n785),.dinb(w_n737_1[0]),.dout(n786));
	jand g0486(.dina(w_n786_0[2]),.dinb(w_n660_0[2]),.dout(n787),.clk(gclk));
	jcb g0487(.dina(n787),.dinb(w_n746_0[1]),.dout(n788));
	jnot g0488(.din(w_n788_0[2]),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n644_0[1]),.dout(n790),.clk(gclk));
	jxor g0490(.dina(w_n648_1[0]),.dinb(w_n790_0[2]),.dout(n791),.clk(gclk));
	jnot g0491(.din(n791),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_n792_0[2]),.dinb(n789),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n788_0[1]),.dinb(w_n790_0[1]),.dout(n794),.clk(gclk));
	jcb g0494(.dina(w_dff_B_1HfbonEU1_0),.dinb(n793),.dout(n795));
	jnot g0495(.din(w_n795_1[1]),.dout(G623_fa_),.clk(gclk));
	jnot g0496(.din(w_G4088_9[2]),.dout(n797),.clk(gclk));
	jnot g0497(.din(w_G861_0),.dout(n798),.clk(gclk));
	jcb g0498(.dina(w_n798_1[1]),.dinb(w_n797_9[1]),.dout(n799));
	jnot g0499(.din(w_G4087_4[2]),.dout(n800),.clk(gclk));
	jnot g0500(.din(w_G822_0),.dout(n801),.clk(gclk));
	jcb g0501(.dina(w_n801_1[1]),.dinb(w_G4088_9[1]),.dout(n802));
	jand g0502(.dina(n802),.dinb(w_n800_4[1]),.dout(n803),.clk(gclk));
	jand g0503(.dina(w_dff_B_lR45vIp78_0),.dinb(n799),.dout(n804),.clk(gclk));
	jcb g0504(.dina(w_n797_9[0]),.dinb(w_G61_0[1]),.dout(n805));
	jcb g0505(.dina(w_G4088_9[0]),.dinb(w_G11_0[1]),.dout(n806));
	jand g0506(.dina(n806),.dinb(w_G4087_4[1]),.dout(n807),.clk(gclk));
	jand g0507(.dina(n807),.dinb(n805),.dout(n808),.clk(gclk));
	jcb g0508(.dina(w_dff_B_UXsIwkmT9_0),.dinb(n804),.dout(G722));
	jand g0509(.dina(w_n750_7[2]),.dinb(w_dff_B_JwiEoX8s2_1),.dout(n810),.clk(gclk));
	jnot g0510(.din(n810),.dout(n811),.clk(gclk));
	jnot g0511(.din(w_n721_0[0]),.dout(n812),.clk(gclk));
	jnot g0512(.din(w_n722_0[0]),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_n631_0[0]),.dinb(w_n377_0[2]),.dout(n814),.clk(gclk));
	jcb g0514(.dina(w_n636_0[1]),.dinb(w_n814_0[2]),.dout(n815));
	jcb g0515(.dina(w_n725_0[1]),.dinb(w_n389_0[2]),.dout(n816));
	jand g0516(.dina(w_n632_0[0]),.dinb(n816),.dout(n817),.clk(gclk));
	jand g0517(.dina(n817),.dinb(n815),.dout(n818),.clk(gclk));
	jcb g0518(.dina(n818),.dinb(w_n726_0[0]),.dout(n819));
	jand g0519(.dina(w_n819_0[2]),.dinb(w_dff_B_UO8pbqDg9_1),.dout(n820),.clk(gclk));
	jcb g0520(.dina(n820),.dinb(w_dff_B_e2WDhi7A7_1),.dout(n821));
	jnot g0521(.din(w_n620_1[0]),.dout(n822),.clk(gclk));
	jnot g0522(.din(w_n639_0[1]),.dout(n823),.clk(gclk));
	jcb g0523(.dina(n823),.dinb(w_n753_0[2]),.dout(n824));
	jcb g0524(.dina(w_n824_0[1]),.dinb(w_dff_B_sedO53ka2_1),.dout(n825));
	jand g0525(.dina(n825),.dinb(w_n821_0[1]),.dout(n826),.clk(gclk));
	jxor g0526(.dina(n826),.dinb(w_n618_0[1]),.dout(n827),.clk(gclk));
	jand g0527(.dina(w_n827_0[1]),.dinb(w_G4091_5[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n445_0[0]),.dinb(w_n749_12[0]),.dout(n829),.clk(gclk));
	jcb g0529(.dina(n829),.dinb(w_G4092_8[1]),.dout(n830));
	jcb g0530(.dina(w_dff_B_sL7vJs5x6_0),.dinb(n828),.dout(n831));
	jand g0531(.dina(n831),.dinb(w_dff_B_9RWlcmWY9_1),.dout(G832_fa_),.clk(gclk));
	jand g0532(.dina(w_n750_7[1]),.dinb(w_dff_B_9OEG3cWT9_1),.dout(n833),.clk(gclk));
	jnot g0533(.din(n833),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n824_0[0]),.dinb(w_n819_0[1]),.dout(n835),.clk(gclk));
	jxor g0535(.dina(n835),.dinb(w_n620_0[2]),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_n836_0[1]),.dinb(w_G4091_4[2]),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_n365_0[0]),.dinb(w_n749_11[2]),.dout(n838),.clk(gclk));
	jcb g0538(.dina(n838),.dinb(w_G4092_8[0]),.dout(n839));
	jcb g0539(.dina(w_dff_B_6H8o4d9y1_0),.dinb(n837),.dout(n840));
	jand g0540(.dina(n840),.dinb(w_dff_B_ETrn17uu3_1),.dout(G834_fa_),.clk(gclk));
	jand g0541(.dina(w_n750_7[0]),.dinb(w_dff_B_qVeNaaDJ7_1),.dout(n842),.clk(gclk));
	jnot g0542(.din(n842),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n397_0[0]),.dinb(w_n749_11[1]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_n637_0[1]),.dinb(w_n753_0[1]),.dout(n845),.clk(gclk));
	jcb g0545(.dina(n845),.dinb(w_n814_0[1]),.dout(n846));
	jxor g0546(.dina(n846),.dinb(w_n624_0[1]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_0[1]),.dinb(w_G4091_4[1]),.dout(n848),.clk(gclk));
	jcb g0548(.dina(n848),.dinb(w_G4092_7[2]),.dout(n849));
	jcb g0549(.dina(n849),.dinb(w_dff_B_7n3YPTJS0_1),.dout(n850));
	jand g0550(.dina(n850),.dinb(w_dff_B_trAlkVrw5_1),.dout(G836_fa_),.clk(gclk));
	jnot g0551(.din(w_G4089_9[2]),.dout(n852),.clk(gclk));
	jcb g0552(.dina(w_n798_1[0]),.dinb(w_n852_9[1]),.dout(n853));
	jnot g0553(.din(w_G4090_4[2]),.dout(n854),.clk(gclk));
	jcb g0554(.dina(w_n801_1[0]),.dinb(w_G4089_9[1]),.dout(n855));
	jand g0555(.dina(n855),.dinb(w_n854_4[1]),.dout(n856),.clk(gclk));
	jand g0556(.dina(w_dff_B_1lmb96HG0_0),.dinb(n853),.dout(n857),.clk(gclk));
	jcb g0557(.dina(w_n852_9[0]),.dinb(w_G61_0[0]),.dout(n858));
	jcb g0558(.dina(w_G4089_9[0]),.dinb(w_G11_0[0]),.dout(n859));
	jand g0559(.dina(n859),.dinb(w_G4090_4[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(n858),.dout(n861),.clk(gclk));
	jcb g0561(.dina(w_dff_B_aSz2eNAo4_0),.dinb(n857),.dout(G859));
	jand g0562(.dina(w_n750_6[2]),.dinb(w_dff_B_c5kHQJeJ9_1),.dout(n863),.clk(gclk));
	jnot g0563(.din(n863),.dout(n864),.clk(gclk));
	jnot g0564(.din(w_n587_0[0]),.dout(n865),.clk(gclk));
	jnot g0565(.din(w_n579_1[0]),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_n567_0[1]),.dinb(w_G4_0[1]),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_n867_0[1]),.dinb(w_n573_0[1]),.dout(n868),.clk(gclk));
	jand g0568(.dina(w_n868_0[1]),.dinb(w_dff_B_fqtln7K09_1),.dout(n869),.clk(gclk));
	jcb g0569(.dina(n869),.dinb(w_n701_0[0]),.dout(n870));
	jxor g0570(.dina(w_n870_0[1]),.dinb(w_n865_0[2]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n871_0[1]),.dinb(w_G4091_4[0]),.dout(n872),.clk(gclk));
	jand g0572(.dina(w_n470_0[0]),.dinb(w_n749_11[0]),.dout(n873),.clk(gclk));
	jcb g0573(.dina(n873),.dinb(w_G4092_7[1]),.dout(n874));
	jcb g0574(.dina(w_dff_B_myhdTuYj6_0),.dinb(n872),.dout(n875));
	jand g0575(.dina(n875),.dinb(w_dff_B_ZsiKmdKd1_1),.dout(G871_fa_),.clk(gclk));
	jand g0576(.dina(w_n750_6[1]),.dinb(w_dff_B_bMPd2nWQ2_1),.dout(n877),.clk(gclk));
	jnot g0577(.din(n877),.dout(n878),.clk(gclk));
	jcb g0578(.dina(w_n868_0[0]),.dinb(w_n699_0[1]),.dout(n879));
	jxor g0579(.dina(n879),.dinb(w_n579_0[2]),.dout(n880),.clk(gclk));
	jand g0580(.dina(w_n880_0[1]),.dinb(w_G4091_3[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n528_0[0]),.dinb(w_n749_10[2]),.dout(n882),.clk(gclk));
	jcb g0582(.dina(n882),.dinb(w_G4092_7[0]),.dout(n883));
	jcb g0583(.dina(w_dff_B_Gip1KnOr8_0),.dinb(n881),.dout(n884));
	jand g0584(.dina(n884),.dinb(w_dff_B_ODrs3Hv98_1),.dout(G873_fa_),.clk(gclk));
	jand g0585(.dina(w_n750_6[0]),.dinb(w_dff_B_Hp7PbKvj2_1),.dout(n886),.clk(gclk));
	jnot g0586(.din(n886),.dout(n887),.clk(gclk));
	jcb g0587(.dina(w_n694_0[1]),.dinb(w_n695_0[1]),.dout(n888));
	jcb g0588(.dina(w_dff_B_z1Eielot2_0),.dinb(w_n867_0[0]),.dout(n889));
	jxor g0589(.dina(n889),.dinb(w_n574_0[1]),.dout(n890),.clk(gclk));
	jand g0590(.dina(w_n890_0[1]),.dinb(w_G4091_3[1]),.dout(n891),.clk(gclk));
	jand g0591(.dina(w_n493_0[0]),.dinb(w_n749_10[1]),.dout(n892),.clk(gclk));
	jcb g0592(.dina(n892),.dinb(w_G4092_6[2]),.dout(n893));
	jcb g0593(.dina(w_dff_B_dLxIWmEe6_0),.dinb(n891),.dout(n894));
	jand g0594(.dina(n894),.dinb(w_dff_B_3QS9wXdt8_1),.dout(G875_fa_),.clk(gclk));
	jand g0595(.dina(w_n750_5[2]),.dinb(w_dff_B_uc5mNuws3_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jnot g0597(.din(w_n566_0[1]),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_n561_0[2]),.dinb(w_G4_0[0]),.dout(n899),.clk(gclk));
	jcb g0599(.dina(n899),.dinb(w_n692_0[0]),.dout(n900));
	jxor g0600(.dina(n900),.dinb(n898),.dout(n901),.clk(gclk));
	jand g0601(.dina(w_n901_0[1]),.dinb(w_G4091_3[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_n481_0[0]),.dinb(w_n749_10[0]),.dout(n903),.clk(gclk));
	jcb g0603(.dina(n903),.dinb(w_G4092_6[1]),.dout(n904));
	jcb g0604(.dina(w_dff_B_D2gjCNcq2_0),.dinb(n902),.dout(n905));
	jand g0605(.dina(n905),.dinb(w_dff_B_aqObUz5T9_1),.dout(G877_fa_),.clk(gclk));
	jnot g0606(.din(w_G331_0[0]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_n619_0[2]),.dout(n908),.clk(gclk));
	jand g0608(.dina(n908),.dinb(w_dff_B_nmbHJMig4_1),.dout(n909),.clk(gclk));
	jand g0609(.dina(w_n619_0[1]),.dinb(w_n617_0[1]),.dout(n910),.clk(gclk));
	jcb g0610(.dina(n910),.dinb(w_dff_B_lprhXOTy9_1),.dout(n911));
	jxor g0611(.dina(w_dff_B_5GvTtmRH5_0),.dinb(w_n792_0[1]),.dout(n912),.clk(gclk));
	jcb g0612(.dina(w_G369_0[0]),.dinb(w_G332_1[0]),.dout(n913));
	jcb g0613(.dina(w_dff_B_jCDCYhlj0_0),.dinb(w_n613_1[2]),.dout(n914));
	jand g0614(.dina(n914),.dinb(w_dff_B_ubAaVd4l6_1),.dout(n915),.clk(gclk));
	jxor g0615(.dina(w_dff_B_ZQaKcf964_0),.dinb(w_n636_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n627_0[1]),.dinb(w_n725_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(w_n658_0[2]),.dinb(w_n653_0[0]),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_dff_B_6hPxrTld8_1),.dout(n919),.clk(gclk));
	jxor g0619(.dina(n919),.dinb(w_dff_B_oLh5Lp4R4_1),.dout(n920),.clk(gclk));
	jxor g0620(.dina(n920),.dinb(n912),.dout(G998_fa_),.clk(gclk));
	jnot g0621(.din(w_n564_0[0]),.dout(n922),.clk(gclk));
	jcb g0622(.dina(n922),.dinb(w_n562_0[0]),.dout(n923));
	jxor g0623(.dina(w_n578_0[1]),.dinb(w_n923_0[2]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n572_0[0]),.dinb(w_n560_0[0]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jcb g0626(.dina(w_G335_0[0]),.dinb(w_G289_0[0]),.dout(n927));
	jcb g0627(.dina(w_n556_2[2]),.dinb(w_dff_B_miCOhRWA2_1),.dout(n928));
	jand g0628(.dina(n928),.dinb(w_dff_B_gagvMuUz4_1),.dout(n929),.clk(gclk));
	jxor g0629(.dina(n929),.dinb(w_n591_0[1]),.dout(n930),.clk(gclk));
	jxor g0630(.dina(w_n596_0[2]),.dinb(w_n586_0[1]),.dout(n931),.clk(gclk));
	jxor g0631(.dina(w_n607_0[1]),.dinb(w_n601_0[1]),.dout(n932),.clk(gclk));
	jxor g0632(.dina(n932),.dinb(n931),.dout(n933),.clk(gclk));
	jxor g0633(.dina(n933),.dinb(w_dff_B_SayaEkvV4_1),.dout(n934),.clk(gclk));
	jxor g0634(.dina(n934),.dinb(w_dff_B_M65zM5Hf2_1),.dout(n935),.clk(gclk));
	jnot g0635(.din(w_n935_0[1]),.dout(G1000),.clk(gclk));
	jnot g0636(.din(w_n592_0[1]),.dout(n937),.clk(gclk));
	jnot g0637(.din(w_n715_0[1]),.dout(n938),.clk(gclk));
	jcb g0638(.dina(w_n870_0[0]),.dinb(w_n682_0[1]),.dout(n939));
	jand g0639(.dina(n939),.dinb(w_n685_0[0]),.dout(n940),.clk(gclk));
	jnot g0640(.din(w_n940_1[1]),.dout(n941),.clk(gclk));
	jcb g0641(.dina(n941),.dinb(w_n609_0[1]),.dout(n942));
	jand g0642(.dina(n942),.dinb(w_n938_0[2]),.dout(n943),.clk(gclk));
	jxor g0643(.dina(n943),.dinb(w_dff_B_vttHX3IB0_1),.dout(n944),.clk(gclk));
	jnot g0644(.din(w_n944_0[1]),.dout(n945),.clk(gclk));
	jnot g0645(.din(w_n603_0[0]),.dout(n946),.clk(gclk));
	jand g0646(.dina(w_n940_1[0]),.dinb(w_dff_B_u6wb1a4G8_1),.dout(n947),.clk(gclk));
	jcb g0647(.dina(n947),.dinb(w_n713_0[1]),.dout(n948));
	jxor g0648(.dina(n948),.dinb(w_n608_0[1]),.dout(n949),.clk(gclk));
	jand g0649(.dina(w_n949_0[1]),.dinb(n945),.dout(n950),.clk(gclk));
	jnot g0650(.din(w_n602_0[1]),.dout(n951),.clk(gclk));
	jnot g0651(.din(w_n596_0[1]),.dout(n952),.clk(gclk));
	jand g0652(.dina(n952),.dinb(w_n496_0[2]),.dout(n953),.clk(gclk));
	jnot g0653(.din(w_n953_0[1]),.dout(n954),.clk(gclk));
	jcb g0654(.dina(w_n940_0[2]),.dinb(w_n710_0[0]),.dout(n955));
	jand g0655(.dina(n955),.dinb(w_n954_0[2]),.dout(n956),.clk(gclk));
	jxor g0656(.dina(n956),.dinb(w_dff_B_8kpeJ6dk8_1),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n957_0[1]),.dout(n958),.clk(gclk));
	jand g0658(.dina(w_n890_0[0]),.dinb(w_n779_0[0]),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(w_n901_0[0]),.dout(n960),.clk(gclk));
	jand g0660(.dina(n960),.dinb(w_n871_0[0]),.dout(n961),.clk(gclk));
	jnot g0661(.din(w_n597_0[1]),.dout(n962),.clk(gclk));
	jxor g0662(.dina(w_n940_0[1]),.dinb(w_n962_0[1]),.dout(n963),.clk(gclk));
	jnot g0663(.din(n963),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_n964_0[1]),.dinb(w_n880_0[0]),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(w_dff_B_Tdu0oli02_1),.dout(n966),.clk(gclk));
	jand g0666(.dina(n966),.dinb(w_dff_B_D04IyGQz9_1),.dout(n967),.clk(gclk));
	jand g0667(.dina(n967),.dinb(n950),.dout(G575),.clk(gclk));
	jxor g0668(.dina(w_n788_0[0]),.dinb(w_n649_0[0]),.dout(n969),.clk(gclk));
	jnot g0669(.din(w_n969_0[1]),.dout(n970),.clk(gclk));
	jand g0670(.dina(n970),.dinb(w_n755_0[0]),.dout(n971),.clk(gclk));
	jand g0671(.dina(w_n836_0[0]),.dinb(w_G623_0),.dout(n972),.clk(gclk));
	jand g0672(.dina(n972),.dinb(w_dff_B_TfsNJWrF9_1),.dout(n973),.clk(gclk));
	jand g0673(.dina(w_n827_0[0]),.dinb(w_n763_0[0]),.dout(n974),.clk(gclk));
	jand g0674(.dina(n974),.dinb(w_n847_0[0]),.dout(n975),.clk(gclk));
	jnot g0675(.din(w_n658_0[1]),.dout(n976),.clk(gclk));
	jand g0676(.dina(n976),.dinb(w_n401_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_n977_0[2]),.dinb(w_n654_2[0]),.dout(n978),.clk(gclk));
	jcb g0678(.dina(w_n977_0[1]),.dinb(w_n654_1[2]),.dout(n979));
	jnot g0679(.din(n979),.dout(n980),.clk(gclk));
	jcb g0680(.dina(w_n786_0[1]),.dinb(w_n742_0[1]),.dout(n981));
	jand g0681(.dina(w_n981_0[1]),.dinb(w_dff_B_BF6jpSG08_1),.dout(n982),.clk(gclk));
	jnot g0682(.din(w_n981_0[0]),.dout(n983),.clk(gclk));
	jand g0683(.dina(n983),.dinb(w_n654_1[1]),.dout(n984),.clk(gclk));
	jcb g0684(.dina(n984),.dinb(w_dff_B_la9Hy5cp1_1),.dout(n985));
	jcb g0685(.dina(n985),.dinb(w_dff_B_DyVAr6xK6_1),.dout(n986));
	jnot g0686(.din(w_n986_0[1]),.dout(n987),.clk(gclk));
	jnot g0687(.din(w_n659_0[0]),.dout(n988),.clk(gclk));
	jxor g0688(.dina(w_n786_0[0]),.dinb(w_dff_B_zz6sdQL49_1),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_n989_0[1]),.dinb(n987),.dout(n990),.clk(gclk));
	jand g0690(.dina(n990),.dinb(w_dff_B_1KWLkI3m7_1),.dout(n991),.clk(gclk));
	jand g0691(.dina(w_dff_B_jFyidKdb4_0),.dinb(n973),.dout(G585),.clk(gclk));
	jnot g0692(.din(w_G1689_5[1]),.dout(n993),.clk(gclk));
	jand g0693(.dina(w_G1690_1[1]),.dinb(w_n993_4[2]),.dout(n994),.clk(gclk));
	jand g0694(.dina(w_n994_4[1]),.dinb(w_G182_0[1]),.dout(n995),.clk(gclk));
	jand g0695(.dina(w_G1690_1[0]),.dinb(w_G1689_5[0]),.dout(n996),.clk(gclk));
	jand g0696(.dina(w_n996_4[1]),.dinb(w_G185_0[1]),.dout(n997),.clk(gclk));
	jcb g0697(.dina(w_n798_0[2]),.dinb(w_n993_4[1]),.dout(n998));
	jnot g0698(.din(w_G1690_0[2]),.dout(n999),.clk(gclk));
	jcb g0699(.dina(w_n801_0[2]),.dinb(w_G1689_4[2]),.dout(n1000));
	jand g0700(.dina(n1000),.dinb(w_n999_3[2]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_dff_B_WqgVAaty1_0),.dinb(n998),.dout(n1002),.clk(gclk));
	jcb g0702(.dina(n1002),.dinb(w_dff_B_PTVEC55W7_1),.dout(n1003));
	jcb g0703(.dina(n1003),.dinb(w_dff_B_Ykn1hPsE6_1),.dout(n1004));
	jand g0704(.dina(n1004),.dinb(w_G137_9[1]),.dout(G661),.clk(gclk));
	jcb g0705(.dina(w_n801_0[1]),.dinb(w_G1691_5[1]),.dout(n1006));
	jnot g0706(.din(w_G1694_1[1]),.dout(n1007),.clk(gclk));
	jnot g0707(.din(w_G1691_5[0]),.dout(n1008),.clk(gclk));
	jcb g0708(.dina(w_n798_0[1]),.dinb(w_n1008_4[2]),.dout(n1009));
	jand g0709(.dina(n1009),.dinb(w_n1007_3[2]),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_dff_B_ZB6kUhF76_1),.dout(n1011),.clk(gclk));
	jand g0711(.dina(w_G1694_1[0]),.dinb(w_G1691_4[2]),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_4[1]),.dinb(w_G185_0[0]),.dout(n1013),.clk(gclk));
	jand g0713(.dina(w_G1694_0[2]),.dinb(w_n1008_4[1]),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_4[1]),.dinb(w_G182_0[0]),.dout(n1015),.clk(gclk));
	jcb g0715(.dina(n1015),.dinb(w_dff_B_VQGxCGCs8_1),.dout(n1016));
	jcb g0716(.dina(w_dff_B_QqXudnfC0_0),.dinb(n1011),.dout(n1017));
	jand g0717(.dina(n1017),.dinb(w_G137_9[0]),.dout(G693),.clk(gclk));
	jnot g0718(.din(w_G871_0),.dout(n1019),.clk(gclk));
	jcb g0719(.dina(w_n1019_1[1]),.dinb(w_n797_8[2]),.dout(n1020));
	jnot g0720(.din(w_G832_0),.dout(n1021),.clk(gclk));
	jcb g0721(.dina(w_n1021_1[1]),.dinb(w_G4088_8[2]),.dout(n1022));
	jand g0722(.dina(n1022),.dinb(w_n800_4[0]),.dout(n1023),.clk(gclk));
	jand g0723(.dina(n1023),.dinb(n1020),.dout(n1024),.clk(gclk));
	jcb g0724(.dina(w_n797_8[1]),.dinb(w_G37_0[1]),.dout(n1025));
	jcb g0725(.dina(w_G4088_8[1]),.dinb(w_G43_0[1]),.dout(n1026));
	jand g0726(.dina(n1026),.dinb(w_G4087_4[0]),.dout(n1027),.clk(gclk));
	jand g0727(.dina(n1027),.dinb(n1025),.dout(n1028),.clk(gclk));
	jcb g0728(.dina(w_dff_B_vGfTQHdt9_0),.dinb(n1024),.dout(G747));
	jnot g0729(.din(w_G873_0),.dout(n1030),.clk(gclk));
	jcb g0730(.dina(w_n1030_1[1]),.dinb(w_n797_8[0]),.dout(n1031));
	jnot g0731(.din(w_G834_0),.dout(n1032),.clk(gclk));
	jcb g0732(.dina(w_n1032_1[1]),.dinb(w_G4088_8[0]),.dout(n1033));
	jand g0733(.dina(n1033),.dinb(w_n800_3[2]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(n1034),.dinb(w_dff_B_34QnpZ2M2_1),.dout(n1035),.clk(gclk));
	jcb g0735(.dina(w_n797_7[2]),.dinb(w_G20_0[1]),.dout(n1036));
	jcb g0736(.dina(w_G4088_7[2]),.dinb(w_G76_0[1]),.dout(n1037));
	jand g0737(.dina(n1037),.dinb(w_G4087_3[2]),.dout(n1038),.clk(gclk));
	jand g0738(.dina(n1038),.dinb(n1036),.dout(n1039),.clk(gclk));
	jcb g0739(.dina(w_dff_B_zNb3Rqgq0_0),.dinb(n1035),.dout(G752));
	jnot g0740(.din(w_G836_0),.dout(n1041),.clk(gclk));
	jcb g0741(.dina(w_n1041_1[1]),.dinb(w_G4088_7[1]),.dout(n1042));
	jnot g0742(.din(w_G875_0),.dout(n1043),.clk(gclk));
	jcb g0743(.dina(w_n1043_1[1]),.dinb(w_n797_7[1]),.dout(n1044));
	jand g0744(.dina(n1044),.dinb(w_n800_3[1]),.dout(n1045),.clk(gclk));
	jand g0745(.dina(n1045),.dinb(w_dff_B_l7ktTNTI3_1),.dout(n1046),.clk(gclk));
	jcb g0746(.dina(w_n797_7[0]),.dinb(w_G17_0[1]),.dout(n1047));
	jcb g0747(.dina(w_G4088_7[0]),.dinb(w_G73_0[1]),.dout(n1048));
	jand g0748(.dina(n1048),.dinb(w_G4087_3[1]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(n1049),.dinb(n1047),.dout(n1050),.clk(gclk));
	jcb g0750(.dina(w_dff_B_Id00WzHI6_0),.dinb(n1046),.dout(G757));
	jnot g0751(.din(w_G877_0),.dout(n1052),.clk(gclk));
	jcb g0752(.dina(w_n1052_1[1]),.dinb(w_n797_6[2]),.dout(n1053));
	jnot g0753(.din(w_G838_0),.dout(n1054),.clk(gclk));
	jcb g0754(.dina(w_n1054_1[1]),.dinb(w_G4088_6[2]),.dout(n1055));
	jand g0755(.dina(n1055),.dinb(w_n800_3[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(n1056),.dinb(w_dff_B_VUAjNiRH7_1),.dout(n1057),.clk(gclk));
	jcb g0757(.dina(w_n797_6[1]),.dinb(w_G70_0[1]),.dout(n1058));
	jcb g0758(.dina(w_G4088_6[1]),.dinb(w_G67_0[1]),.dout(n1059));
	jand g0759(.dina(n1059),.dinb(w_G4087_3[0]),.dout(n1060),.clk(gclk));
	jand g0760(.dina(n1060),.dinb(n1058),.dout(n1061),.clk(gclk));
	jcb g0761(.dina(w_dff_B_2fehSlEE1_0),.dinb(n1057),.dout(G762));
	jcb g0762(.dina(w_G4089_8[2]),.dinb(w_G43_0[0]),.dout(n1063));
	jcb g0763(.dina(w_n852_8[2]),.dinb(w_G37_0[0]),.dout(n1064));
	jand g0764(.dina(n1064),.dinb(w_G4090_4[0]),.dout(n1065),.clk(gclk));
	jand g0765(.dina(n1065),.dinb(w_dff_B_jLkq5yPJ4_1),.dout(n1066),.clk(gclk));
	jcb g0766(.dina(w_n1021_1[0]),.dinb(w_G4089_8[1]),.dout(n1067));
	jcb g0767(.dina(w_n1019_1[0]),.dinb(w_n852_8[1]),.dout(n1068));
	jand g0768(.dina(n1068),.dinb(w_dff_B_8cMfT4eI0_1),.dout(n1069),.clk(gclk));
	jand g0769(.dina(n1069),.dinb(w_n854_4[0]),.dout(n1070),.clk(gclk));
	jcb g0770(.dina(n1070),.dinb(w_dff_B_e1pr8F9p2_1),.dout(G787));
	jcb g0771(.dina(w_G4089_8[0]),.dinb(w_G76_0[0]),.dout(n1072));
	jcb g0772(.dina(w_n852_8[0]),.dinb(w_G20_0[0]),.dout(n1073));
	jand g0773(.dina(n1073),.dinb(w_G4090_3[2]),.dout(n1074),.clk(gclk));
	jand g0774(.dina(n1074),.dinb(w_dff_B_ZC7hCloA9_1),.dout(n1075),.clk(gclk));
	jcb g0775(.dina(w_n1032_1[0]),.dinb(w_G4089_7[2]),.dout(n1076));
	jcb g0776(.dina(w_n1030_1[0]),.dinb(w_n852_7[2]),.dout(n1077));
	jand g0777(.dina(n1077),.dinb(n1076),.dout(n1078),.clk(gclk));
	jand g0778(.dina(n1078),.dinb(w_n854_3[2]),.dout(n1079),.clk(gclk));
	jcb g0779(.dina(n1079),.dinb(w_dff_B_Znv1cIZd9_1),.dout(G792));
	jcb g0780(.dina(w_G4089_7[1]),.dinb(w_G73_0[0]),.dout(n1081));
	jcb g0781(.dina(w_n852_7[1]),.dinb(w_G17_0[0]),.dout(n1082));
	jand g0782(.dina(n1082),.dinb(w_G4090_3[1]),.dout(n1083),.clk(gclk));
	jand g0783(.dina(n1083),.dinb(w_dff_B_JvDrFjIk7_1),.dout(n1084),.clk(gclk));
	jcb g0784(.dina(w_n1043_1[0]),.dinb(w_n852_7[0]),.dout(n1085));
	jcb g0785(.dina(w_n1041_1[0]),.dinb(w_G4089_7[0]),.dout(n1086));
	jand g0786(.dina(w_dff_B_a5h5n6Vd2_0),.dinb(n1085),.dout(n1087),.clk(gclk));
	jand g0787(.dina(n1087),.dinb(w_n854_3[1]),.dout(n1088),.clk(gclk));
	jcb g0788(.dina(n1088),.dinb(w_dff_B_9czpcr7Z2_1),.dout(G797));
	jcb g0789(.dina(w_n1052_1[0]),.dinb(w_n852_6[2]),.dout(n1090));
	jcb g0790(.dina(w_n1054_1[0]),.dinb(w_G4089_6[2]),.dout(n1091));
	jand g0791(.dina(n1091),.dinb(w_n854_3[0]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(n1092),.dinb(w_dff_B_GtnUh3fp5_1),.dout(n1093),.clk(gclk));
	jcb g0793(.dina(w_n852_6[1]),.dinb(w_G70_0[0]),.dout(n1094));
	jcb g0794(.dina(w_G4089_6[1]),.dinb(w_G67_0[0]),.dout(n1095));
	jand g0795(.dina(n1095),.dinb(w_G4090_3[0]),.dout(n1096),.clk(gclk));
	jand g0796(.dina(n1096),.dinb(n1094),.dout(n1097),.clk(gclk));
	jcb g0797(.dina(w_dff_B_rOZqIJ489_0),.dinb(n1093),.dout(G802));
	jcb g0798(.dina(w_n1021_0[2]),.dinb(w_G1689_4[1]),.dout(n1099));
	jcb g0799(.dina(w_n1019_0[2]),.dinb(w_n993_4[0]),.dout(n1100));
	jand g0800(.dina(n1100),.dinb(w_n999_3[1]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(n1101),.dinb(w_dff_B_dHD2NsdS6_1),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n994_4[0]),.dinb(w_G200_0[1]),.dout(n1103),.clk(gclk));
	jand g0803(.dina(w_n996_4[0]),.dinb(w_G170_0[1]),.dout(n1104),.clk(gclk));
	jcb g0804(.dina(w_dff_B_Zg1UhuNn4_0),.dinb(n1103),.dout(n1105));
	jcb g0805(.dina(w_dff_B_L0foX1gb2_0),.dinb(n1102),.dout(n1106));
	jand g0806(.dina(n1106),.dinb(w_G137_8[2]),.dout(G642),.clk(gclk));
	jcb g0807(.dina(w_n1054_0[2]),.dinb(w_G1689_4[0]),.dout(n1108));
	jcb g0808(.dina(w_n1052_0[2]),.dinb(w_n993_3[2]),.dout(n1109));
	jand g0809(.dina(n1109),.dinb(w_n999_3[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(n1110),.dinb(w_dff_B_lLyMDWw12_1),.dout(n1111),.clk(gclk));
	jand g0811(.dina(w_n994_3[2]),.dinb(w_G188_0[1]),.dout(n1112),.clk(gclk));
	jand g0812(.dina(w_n996_3[2]),.dinb(w_G158_0[1]),.dout(n1113),.clk(gclk));
	jcb g0813(.dina(w_dff_B_OKBEGDpY5_0),.dinb(n1112),.dout(n1114));
	jcb g0814(.dina(w_dff_B_4wdvpaih2_0),.dinb(n1111),.dout(n1115));
	jand g0815(.dina(n1115),.dinb(w_G137_8[1]),.dout(G664),.clk(gclk));
	jcb g0816(.dina(w_n1041_0[2]),.dinb(w_G1689_3[2]),.dout(n1117));
	jcb g0817(.dina(w_n1043_0[2]),.dinb(w_n993_3[1]),.dout(n1118));
	jand g0818(.dina(n1118),.dinb(w_n999_2[2]),.dout(n1119),.clk(gclk));
	jand g0819(.dina(n1119),.dinb(w_dff_B_4Z6Nypry4_1),.dout(n1120),.clk(gclk));
	jand g0820(.dina(w_n994_3[1]),.dinb(w_G155_0[1]),.dout(n1121),.clk(gclk));
	jand g0821(.dina(w_n996_3[1]),.dinb(w_G152_0[1]),.dout(n1122),.clk(gclk));
	jcb g0822(.dina(w_dff_B_OL3NLugM8_0),.dinb(n1121),.dout(n1123));
	jcb g0823(.dina(w_dff_B_LuGLwxXH5_0),.dinb(n1120),.dout(n1124));
	jand g0824(.dina(n1124),.dinb(w_G137_8[0]),.dout(G667),.clk(gclk));
	jcb g0825(.dina(w_n1032_0[2]),.dinb(w_G1689_3[1]),.dout(n1126));
	jcb g0826(.dina(w_n1030_0[2]),.dinb(w_n993_3[0]),.dout(n1127));
	jand g0827(.dina(n1127),.dinb(w_n999_2[1]),.dout(n1128),.clk(gclk));
	jand g0828(.dina(n1128),.dinb(w_dff_B_rNLC0A6b9_1),.dout(n1129),.clk(gclk));
	jand g0829(.dina(w_n994_3[0]),.dinb(w_G149_0[1]),.dout(n1130),.clk(gclk));
	jand g0830(.dina(w_n996_3[0]),.dinb(w_G146_0[1]),.dout(n1131),.clk(gclk));
	jcb g0831(.dina(w_dff_B_TRI8VtAe1_0),.dinb(n1130),.dout(n1132));
	jcb g0832(.dina(w_dff_B_mzqMQWYO7_0),.dinb(n1129),.dout(n1133));
	jand g0833(.dina(n1133),.dinb(w_G137_7[2]),.dout(G670),.clk(gclk));
	jand g0834(.dina(w_n1014_4[0]),.dinb(w_G200_0[0]),.dout(n1135),.clk(gclk));
	jand g0835(.dina(w_n1012_4[0]),.dinb(w_G170_0[0]),.dout(n1136),.clk(gclk));
	jcb g0836(.dina(w_n1019_0[1]),.dinb(w_n1008_4[0]),.dout(n1137));
	jcb g0837(.dina(w_n1021_0[1]),.dinb(w_G1691_4[1]),.dout(n1138));
	jand g0838(.dina(w_dff_B_beWqPsAs9_0),.dinb(n1137),.dout(n1139),.clk(gclk));
	jand g0839(.dina(n1139),.dinb(w_n1007_3[1]),.dout(n1140),.clk(gclk));
	jcb g0840(.dina(n1140),.dinb(w_dff_B_039QYSRB1_1),.dout(n1141));
	jcb g0841(.dina(n1141),.dinb(w_dff_B_O8UO2SZW0_1),.dout(n1142));
	jand g0842(.dina(n1142),.dinb(w_G137_7[1]),.dout(G676),.clk(gclk));
	jcb g0843(.dina(w_n1054_0[1]),.dinb(w_G1691_4[0]),.dout(n1144));
	jcb g0844(.dina(w_n1052_0[1]),.dinb(w_n1008_3[2]),.dout(n1145));
	jand g0845(.dina(n1145),.dinb(w_n1007_3[0]),.dout(n1146),.clk(gclk));
	jand g0846(.dina(n1146),.dinb(w_dff_B_6d5lY3U59_1),.dout(n1147),.clk(gclk));
	jand g0847(.dina(w_n1014_3[2]),.dinb(w_G188_0[0]),.dout(n1148),.clk(gclk));
	jand g0848(.dina(w_n1012_3[2]),.dinb(w_G158_0[0]),.dout(n1149),.clk(gclk));
	jcb g0849(.dina(w_dff_B_Nxu03oUQ0_0),.dinb(n1148),.dout(n1150));
	jcb g0850(.dina(w_dff_B_7VhNgJT62_0),.dinb(n1147),.dout(n1151));
	jand g0851(.dina(n1151),.dinb(w_G137_7[0]),.dout(G696),.clk(gclk));
	jcb g0852(.dina(w_n1041_0[1]),.dinb(w_G1691_3[2]),.dout(n1153));
	jcb g0853(.dina(w_n1043_0[1]),.dinb(w_n1008_3[1]),.dout(n1154));
	jand g0854(.dina(n1154),.dinb(w_n1007_2[2]),.dout(n1155),.clk(gclk));
	jand g0855(.dina(n1155),.dinb(w_dff_B_knRvT7tP7_1),.dout(n1156),.clk(gclk));
	jand g0856(.dina(w_n1014_3[1]),.dinb(w_G155_0[0]),.dout(n1157),.clk(gclk));
	jand g0857(.dina(w_n1012_3[1]),.dinb(w_G152_0[0]),.dout(n1158),.clk(gclk));
	jcb g0858(.dina(w_dff_B_oc0B1lNu8_0),.dinb(n1157),.dout(n1159));
	jcb g0859(.dina(w_dff_B_tb7gYmZ10_0),.dinb(n1156),.dout(n1160));
	jand g0860(.dina(n1160),.dinb(w_G137_6[2]),.dout(G699),.clk(gclk));
	jcb g0861(.dina(w_n1032_0[1]),.dinb(w_G1691_3[1]),.dout(n1162));
	jcb g0862(.dina(w_n1030_0[1]),.dinb(w_n1008_3[0]),.dout(n1163));
	jand g0863(.dina(n1163),.dinb(w_n1007_2[1]),.dout(n1164),.clk(gclk));
	jand g0864(.dina(n1164),.dinb(w_dff_B_wnl81Iyh3_1),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n1014_3[0]),.dinb(w_G149_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n1012_3[0]),.dinb(w_G146_0[0]),.dout(n1167),.clk(gclk));
	jcb g0867(.dina(w_dff_B_8jjA69mY4_0),.dinb(n1166),.dout(n1168));
	jcb g0868(.dina(w_dff_B_coJcKL1t1_0),.dinb(n1165),.dout(n1169));
	jand g0869(.dina(n1169),.dinb(w_G137_6[1]),.dout(G702),.clk(gclk));
	jnot g0870(.din(G135),.dout(n1171),.clk(gclk));
	jnot g0871(.din(G4115),.dout(n1172),.clk(gclk));
	jcb g0872(.dina(n1172),.dinb(n1171),.dout(n1173));
	jnot g0873(.din(w_n428_1[0]),.dout(n1174),.clk(gclk));
	jcb g0874(.dina(n1174),.dinb(w_G3724_0[2]),.dout(n1175));
	jnot g0875(.din(w_G3717_0[1]),.dout(n1176),.clk(gclk));
	jnot g0876(.din(w_G3724_0[1]),.dout(n1177),.clk(gclk));
	jxor g0877(.dina(w_n790_0[0]),.dinb(w_dff_B_K6VgBYY54_1),.dout(n1178),.clk(gclk));
	jnot g0878(.din(n1178),.dout(n1179),.clk(gclk));
	jcb g0879(.dina(w_n1179_0[1]),.dinb(w_n1177_0[1]),.dout(n1180));
	jand g0880(.dina(n1180),.dinb(w_dff_B_P0bI9bgD6_1),.dout(n1181),.clk(gclk));
	jand g0881(.dina(n1181),.dinb(w_dff_B_KgvbjEim3_1),.dout(n1182),.clk(gclk));
	jcb g0882(.dina(w_n795_1[0]),.dinb(w_n1177_0[0]),.dout(n1183));
	jcb g0883(.dina(w_G3724_0[0]),.dinb(w_G123_0[1]),.dout(n1184));
	jand g0884(.dina(n1184),.dinb(w_G3717_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(w_dff_B_KnwnaKGM1_0),.dinb(n1183),.dout(n1186),.clk(gclk));
	jcb g0886(.dina(n1186),.dinb(w_dff_B_Xt9Y9EYs6_1),.dout(n1187));
	jand g0887(.dina(n1187),.dinb(w_dff_B_2u0ShZUG1_1),.dout(G818),.clk(gclk));
	jxor g0888(.dina(w_n1179_0[0]),.dinb(w_n795_0[2]),.dout(G813),.clk(gclk));
	jand g0889(.dina(w_n750_5[1]),.dinb(w_G123_0[0]),.dout(n1190),.clk(gclk));
	jcb g0890(.dina(w_n795_0[1]),.dinb(w_n749_9[2]),.dout(n1191));
	jand g0891(.dina(w_n428_0[2]),.dinb(w_n749_9[1]),.dout(n1192),.clk(gclk));
	jcb g0892(.dina(n1192),.dinb(w_G4092_6[0]),.dout(n1193));
	jnot g0893(.din(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_dff_B_0ppLAxZZ8_0),.dinb(n1191),.dout(n1195),.clk(gclk));
	jcb g0895(.dina(n1195),.dinb(w_dff_B_QRrdICxI0_1),.dout(n1196));
	jnot g0896(.din(w_n1196_1[2]),.dout(G824),.clk(gclk));
	jand g0897(.dina(w_n750_5[0]),.dinb(w_dff_B_WmGzb8lC6_1),.dout(n1198),.clk(gclk));
	jand g0898(.dina(w_n433_0[1]),.dinb(w_n749_9[0]),.dout(n1199),.clk(gclk));
	jnot g0899(.din(n1199),.dout(n1200),.clk(gclk));
	jnot g0900(.din(w_G4092_5[2]),.dout(n1201),.clk(gclk));
	jcb g0901(.dina(w_n969_0[0]),.dinb(w_n749_8[2]),.dout(n1202));
	jand g0902(.dina(n1202),.dinb(w_n1201_0[2]),.dout(n1203),.clk(gclk));
	jand g0903(.dina(n1203),.dinb(w_dff_B_JPiiHemD4_1),.dout(n1204),.clk(gclk));
	jcb g0904(.dina(n1204),.dinb(w_dff_B_sZyG1Hue7_1),.dout(n1205));
	jnot g0905(.din(w_n1205_1[2]),.dout(G826),.clk(gclk));
	jand g0906(.dina(w_n750_4[2]),.dinb(w_dff_B_bxnokhrt3_1),.dout(n1207),.clk(gclk));
	jcb g0907(.dina(w_n986_0[0]),.dinb(w_n749_8[1]),.dout(n1208));
	jand g0908(.dina(w_n423_0[1]),.dinb(w_n749_8[0]),.dout(n1209),.clk(gclk));
	jcb g0909(.dina(n1209),.dinb(w_G4092_5[1]),.dout(n1210));
	jnot g0910(.din(n1210),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_9LvvXecj4_0),.dinb(n1208),.dout(n1212),.clk(gclk));
	jcb g0912(.dina(n1212),.dinb(w_dff_B_l0lvpBRH7_1),.dout(n1213));
	jnot g0913(.din(w_n1213_1[2]),.dout(G828),.clk(gclk));
	jand g0914(.dina(w_n750_4[1]),.dinb(w_dff_B_WdEBxlLx2_1),.dout(n1215),.clk(gclk));
	jnot g0915(.din(n1215),.dout(n1216),.clk(gclk));
	jand g0916(.dina(w_n989_0[0]),.dinb(w_G4091_2[2]),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_n412_0[1]),.dinb(w_n749_7[2]),.dout(n1218),.clk(gclk));
	jcb g0918(.dina(n1218),.dinb(w_G4092_5[0]),.dout(n1219));
	jcb g0919(.dina(w_dff_B_xnScEtc77_0),.dinb(n1217),.dout(n1220));
	jand g0920(.dina(n1220),.dinb(w_dff_B_tQhKUQkb1_1),.dout(G830_fa_),.clk(gclk));
	jand g0921(.dina(w_n680_0[0]),.dinb(w_G245_0[0]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_dff_B_yQZ9oo2Z6_0),.dinb(w_n935_0[0]),.dout(n1223),.clk(gclk));
	jnot g0923(.din(w_G998_0),.dout(n1224),.clk(gclk));
	jand g0924(.dina(w_n318_0[0]),.dinb(w_G601_0),.dout(n1225),.clk(gclk));
	jand g0925(.dina(n1225),.dinb(w_G559_0[0]),.dout(n1226),.clk(gclk));
	jand g0926(.dina(w_dff_B_CqnFOVbl3_0),.dinb(w_n670_0[0]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_dff_B_kmLJ1tZm4_0),.dinb(n1224),.dout(n1228),.clk(gclk));
	jand g0928(.dina(n1228),.dinb(w_dff_B_oRispRRq4_1),.dout(G854),.clk(gclk));
	jand g0929(.dina(w_n750_4[0]),.dinb(w_dff_B_DhEh2tGG5_1),.dout(n1230),.clk(gclk));
	jand g0930(.dina(w_n551_0[1]),.dinb(w_n749_7[1]),.dout(n1231),.clk(gclk));
	jnot g0931(.din(n1231),.dout(n1232),.clk(gclk));
	jcb g0932(.dina(w_n944_0[0]),.dinb(w_n749_7[0]),.dout(n1233));
	jand g0933(.dina(n1233),.dinb(w_n1201_0[1]),.dout(n1234),.clk(gclk));
	jand g0934(.dina(n1234),.dinb(w_dff_B_lViDy4wq4_1),.dout(n1235),.clk(gclk));
	jcb g0935(.dina(n1235),.dinb(w_dff_B_Z5W0Ta4I1_1),.dout(n1236));
	jnot g0936(.din(w_n1236_1[2]),.dout(G863),.clk(gclk));
	jand g0937(.dina(w_n750_3[2]),.dinb(w_dff_B_mtf1kKtJ0_1),.dout(n1238),.clk(gclk));
	jnot g0938(.din(n1238),.dout(n1239),.clk(gclk));
	jand g0939(.dina(w_n949_0[0]),.dinb(w_G4091_2[1]),.dout(n1240),.clk(gclk));
	jand g0940(.dina(w_n459_0[0]),.dinb(w_n749_6[2]),.dout(n1241),.clk(gclk));
	jcb g0941(.dina(n1241),.dinb(w_G4092_4[2]),.dout(n1242));
	jcb g0942(.dina(w_dff_B_EDvBLAjE8_0),.dinb(n1240),.dout(n1243));
	jand g0943(.dina(n1243),.dinb(w_dff_B_8k09gzto0_1),.dout(G865_fa_),.clk(gclk));
	jand g0944(.dina(w_n750_3[1]),.dinb(w_dff_B_fyVm4Obu7_1),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n517_0[0]),.dinb(w_n749_6[1]),.dout(n1246),.clk(gclk));
	jnot g0946(.din(n1246),.dout(n1247),.clk(gclk));
	jcb g0947(.dina(w_n957_0[0]),.dinb(w_n749_6[0]),.dout(n1248));
	jand g0948(.dina(n1248),.dinb(w_n1201_0[0]),.dout(n1249),.clk(gclk));
	jand g0949(.dina(n1249),.dinb(w_dff_B_F2YdCrcQ2_1),.dout(n1250),.clk(gclk));
	jcb g0950(.dina(n1250),.dinb(w_dff_B_8v49LUSi5_1),.dout(n1251));
	jnot g0951(.din(w_n1251_1[2]),.dout(G867),.clk(gclk));
	jand g0952(.dina(w_n750_3[0]),.dinb(w_dff_B_mQPe3CN02_1),.dout(n1253),.clk(gclk));
	jnot g0953(.din(n1253),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n964_0[0]),.dinb(w_G4091_2[0]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n504_0[0]),.dinb(w_n749_5[2]),.dout(n1256),.clk(gclk));
	jcb g0956(.dina(n1256),.dinb(w_G4092_4[1]),.dout(n1257));
	jcb g0957(.dina(w_dff_B_doZsvJYt5_0),.dinb(n1255),.dout(n1258));
	jand g0958(.dina(n1258),.dinb(w_dff_B_3KgK7ttF1_1),.dout(G869_fa_),.clk(gclk));
	jcb g0959(.dina(w_G4089_6[0]),.dinb(w_G109_0[1]),.dout(n1260));
	jcb g0960(.dina(w_n852_6[0]),.dinb(w_G106_0[1]),.dout(n1261));
	jand g0961(.dina(n1261),.dinb(w_G4090_2[2]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(n1262),.dinb(w_dff_B_oIzlAM068_1),.dout(n1263),.clk(gclk));
	jcb g0963(.dina(w_n1236_1[1]),.dinb(w_n852_5[2]),.dout(n1264));
	jcb g0964(.dina(w_n1196_1[1]),.dinb(w_G4089_5[2]),.dout(n1265));
	jand g0965(.dina(n1265),.dinb(w_n854_2[2]),.dout(n1266),.clk(gclk));
	jand g0966(.dina(w_dff_B_l5liVw6T3_0),.dinb(n1264),.dout(n1267),.clk(gclk));
	jcb g0967(.dina(n1267),.dinb(w_dff_B_UpTPaB8V4_1),.dout(G712));
	jcb g0968(.dina(w_n1196_1[0]),.dinb(w_G4088_6[0]),.dout(n1269));
	jcb g0969(.dina(w_n1236_1[0]),.dinb(w_n797_6[0]),.dout(n1270));
	jand g0970(.dina(n1270),.dinb(w_n800_2[2]),.dout(n1271),.clk(gclk));
	jand g0971(.dina(n1271),.dinb(w_dff_B_beRkpLEE2_1),.dout(n1272),.clk(gclk));
	jcb g0972(.dina(w_n797_5[2]),.dinb(w_G106_0[0]),.dout(n1273));
	jcb g0973(.dina(w_G4088_5[2]),.dinb(w_G109_0[0]),.dout(n1274));
	jand g0974(.dina(n1274),.dinb(w_G4087_2[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(n1275),.dinb(n1273),.dout(n1276),.clk(gclk));
	jcb g0976(.dina(w_dff_B_cP2vFUK47_0),.dinb(n1272),.dout(G727));
	jcb g0977(.dina(w_n1205_1[1]),.dinb(w_G4088_5[1]),.dout(n1278));
	jnot g0978(.din(w_G865_0),.dout(n1279),.clk(gclk));
	jcb g0979(.dina(w_n1279_1[1]),.dinb(w_n797_5[1]),.dout(n1280));
	jand g0980(.dina(n1280),.dinb(w_n800_2[1]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(n1281),.dinb(w_dff_B_VvxiDDw61_1),.dout(n1282),.clk(gclk));
	jcb g0982(.dina(w_n797_5[0]),.dinb(w_G49_0[1]),.dout(n1283));
	jcb g0983(.dina(w_G4088_5[0]),.dinb(w_G46_0[1]),.dout(n1284));
	jand g0984(.dina(n1284),.dinb(w_G4087_2[1]),.dout(n1285),.clk(gclk));
	jand g0985(.dina(n1285),.dinb(n1283),.dout(n1286),.clk(gclk));
	jcb g0986(.dina(w_dff_B_fbzNMePi9_0),.dinb(n1282),.dout(G732));
	jcb g0987(.dina(w_n1213_1[1]),.dinb(w_G4088_4[2]),.dout(n1288));
	jcb g0988(.dina(w_n1251_1[1]),.dinb(w_n797_4[2]),.dout(n1289));
	jand g0989(.dina(n1289),.dinb(w_n800_2[0]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(n1290),.dinb(w_dff_B_CFSdghtJ8_1),.dout(n1291),.clk(gclk));
	jcb g0991(.dina(w_n797_4[1]),.dinb(w_G103_0[1]),.dout(n1292));
	jcb g0992(.dina(w_G4088_4[1]),.dinb(w_G100_0[1]),.dout(n1293));
	jand g0993(.dina(n1293),.dinb(w_G4087_2[0]),.dout(n1294),.clk(gclk));
	jand g0994(.dina(n1294),.dinb(n1292),.dout(n1295),.clk(gclk));
	jcb g0995(.dina(w_dff_B_3RpqSXkc4_0),.dinb(n1291),.dout(G737));
	jnot g0996(.din(w_G830_0),.dout(n1297),.clk(gclk));
	jcb g0997(.dina(w_n1297_1[1]),.dinb(w_G4088_4[0]),.dout(n1298));
	jnot g0998(.din(w_G869_0),.dout(n1299),.clk(gclk));
	jcb g0999(.dina(w_n1299_1[1]),.dinb(w_n797_4[0]),.dout(n1300));
	jand g1000(.dina(n1300),.dinb(w_n800_1[2]),.dout(n1301),.clk(gclk));
	jand g1001(.dina(n1301),.dinb(w_dff_B_DCa37vzH1_1),.dout(n1302),.clk(gclk));
	jcb g1002(.dina(w_n797_3[2]),.dinb(w_G40_0[1]),.dout(n1303));
	jcb g1003(.dina(w_G4088_3[2]),.dinb(w_G91_0[1]),.dout(n1304));
	jand g1004(.dina(n1304),.dinb(w_G4087_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(n1305),.dinb(n1303),.dout(n1306),.clk(gclk));
	jcb g1006(.dina(w_dff_B_xeFe8tDL3_0),.dinb(n1302),.dout(G742));
	jcb g1007(.dina(w_n1205_1[0]),.dinb(w_G4089_5[1]),.dout(n1308));
	jcb g1008(.dina(w_n1279_1[0]),.dinb(w_n852_5[1]),.dout(n1309));
	jand g1009(.dina(n1309),.dinb(w_n854_2[1]),.dout(n1310),.clk(gclk));
	jand g1010(.dina(n1310),.dinb(w_dff_B_jxdHE5yx0_1),.dout(n1311),.clk(gclk));
	jcb g1011(.dina(w_n852_5[0]),.dinb(w_G49_0[0]),.dout(n1312));
	jcb g1012(.dina(w_G4089_5[0]),.dinb(w_G46_0[0]),.dout(n1313));
	jand g1013(.dina(n1313),.dinb(w_G4090_2[1]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(n1314),.dinb(n1312),.dout(n1315),.clk(gclk));
	jcb g1015(.dina(w_dff_B_IBbsAM0P4_0),.dinb(n1311),.dout(G772));
	jcb g1016(.dina(w_n1213_1[0]),.dinb(w_G4089_4[2]),.dout(n1317));
	jcb g1017(.dina(w_n1251_1[0]),.dinb(w_n852_4[2]),.dout(n1318));
	jand g1018(.dina(n1318),.dinb(w_n854_2[0]),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_dff_B_vOeuLJoV2_1),.dout(n1320),.clk(gclk));
	jcb g1020(.dina(w_n852_4[1]),.dinb(w_G103_0[0]),.dout(n1321));
	jcb g1021(.dina(w_G4089_4[1]),.dinb(w_G100_0[0]),.dout(n1322));
	jand g1022(.dina(n1322),.dinb(w_G4090_2[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(n1323),.dinb(n1321),.dout(n1324),.clk(gclk));
	jcb g1024(.dina(w_dff_B_rfKSEMge0_0),.dinb(n1320),.dout(G777));
	jcb g1025(.dina(w_n1297_1[0]),.dinb(w_G4089_4[0]),.dout(n1326));
	jcb g1026(.dina(w_n1299_1[0]),.dinb(w_n852_4[0]),.dout(n1327));
	jand g1027(.dina(n1327),.dinb(w_n854_1[2]),.dout(n1328),.clk(gclk));
	jand g1028(.dina(n1328),.dinb(w_dff_B_vCC4io5f0_1),.dout(n1329),.clk(gclk));
	jcb g1029(.dina(w_n852_3[2]),.dinb(w_G40_0[0]),.dout(n1330));
	jcb g1030(.dina(w_G4089_3[2]),.dinb(w_G91_0[0]),.dout(n1331));
	jand g1031(.dina(n1331),.dinb(w_G4090_1[2]),.dout(n1332),.clk(gclk));
	jand g1032(.dina(n1332),.dinb(n1330),.dout(n1333),.clk(gclk));
	jcb g1033(.dina(w_dff_B_1e1NwGhf7_0),.dinb(n1329),.dout(G782));
	jcb g1034(.dina(w_n1297_0[2]),.dinb(w_G1689_3[0]),.dout(n1335));
	jcb g1035(.dina(w_n1299_0[2]),.dinb(w_n993_2[2]),.dout(n1336));
	jand g1036(.dina(n1336),.dinb(w_n999_2[0]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(n1337),.dinb(w_dff_B_TvoVTqyh9_1),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n994_2[2]),.dinb(w_G203_0[1]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n996_2[2]),.dinb(w_G173_0[1]),.dout(n1340),.clk(gclk));
	jcb g1040(.dina(w_dff_B_y8RlDIqL2_0),.dinb(n1339),.dout(n1341));
	jcb g1041(.dina(w_dff_B_qyRUhJ1b1_0),.dinb(n1338),.dout(n1342));
	jand g1042(.dina(n1342),.dinb(w_G137_6[0]),.dout(G645),.clk(gclk));
	jcb g1043(.dina(w_n1251_0[2]),.dinb(w_n993_2[1]),.dout(n1344));
	jcb g1044(.dina(w_n1213_0[2]),.dinb(w_G1689_2[2]),.dout(n1345));
	jand g1045(.dina(n1345),.dinb(w_n999_1[2]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(w_dff_B_cc0SnLEB2_0),.dinb(n1344),.dout(n1347),.clk(gclk));
	jand g1047(.dina(w_n994_2[1]),.dinb(w_G197_0[1]),.dout(n1348),.clk(gclk));
	jand g1048(.dina(w_n996_2[1]),.dinb(w_G167_0[1]),.dout(n1349),.clk(gclk));
	jcb g1049(.dina(w_dff_B_CvCeRqJO4_0),.dinb(n1348),.dout(n1350));
	jcb g1050(.dina(w_dff_B_ZNHaclVH4_0),.dinb(n1347),.dout(n1351));
	jand g1051(.dina(n1351),.dinb(w_G137_5[2]),.dout(G648),.clk(gclk));
	jand g1052(.dina(w_n994_2[0]),.dinb(w_G194_0[1]),.dout(n1353),.clk(gclk));
	jand g1053(.dina(w_n996_2[0]),.dinb(w_G164_0[1]),.dout(n1354),.clk(gclk));
	jcb g1054(.dina(w_dff_B_pLg1x5Uh2_0),.dinb(n1353),.dout(n1355));
	jcb g1055(.dina(w_n1205_0[2]),.dinb(w_G1689_2[1]),.dout(n1356));
	jcb g1056(.dina(w_n1279_0[2]),.dinb(w_n993_2[0]),.dout(n1357));
	jand g1057(.dina(n1357),.dinb(w_dff_B_8BAIfOQ66_1),.dout(n1358),.clk(gclk));
	jand g1058(.dina(n1358),.dinb(w_n999_1[1]),.dout(n1359),.clk(gclk));
	jcb g1059(.dina(n1359),.dinb(w_dff_B_UIxyaktK2_1),.dout(n1360));
	jand g1060(.dina(n1360),.dinb(w_G137_5[1]),.dout(G651),.clk(gclk));
	jand g1061(.dina(w_n994_1[2]),.dinb(w_G191_0[1]),.dout(n1362),.clk(gclk));
	jand g1062(.dina(w_n996_1[2]),.dinb(w_G161_0[1]),.dout(n1363),.clk(gclk));
	jcb g1063(.dina(w_dff_B_3wmX0kaV8_0),.dinb(n1362),.dout(n1364));
	jcb g1064(.dina(w_n1196_0[2]),.dinb(w_G1689_2[0]),.dout(n1365));
	jcb g1065(.dina(w_n1236_0[2]),.dinb(w_n993_1[2]),.dout(n1366));
	jand g1066(.dina(n1366),.dinb(w_dff_B_zlpaa5gV7_1),.dout(n1367),.clk(gclk));
	jand g1067(.dina(n1367),.dinb(w_n999_1[0]),.dout(n1368),.clk(gclk));
	jcb g1068(.dina(n1368),.dinb(w_dff_B_ISUm5JJD8_1),.dout(n1369));
	jand g1069(.dina(n1369),.dinb(w_G137_5[0]),.dout(G654),.clk(gclk));
	jcb g1070(.dina(w_n1297_0[1]),.dinb(w_G1691_3[0]),.dout(n1371));
	jcb g1071(.dina(w_n1299_0[1]),.dinb(w_n1008_2[2]),.dout(n1372));
	jand g1072(.dina(n1372),.dinb(w_n1007_2[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(n1373),.dinb(w_dff_B_Maw3qAoo6_1),.dout(n1374),.clk(gclk));
	jand g1074(.dina(w_n1014_2[2]),.dinb(w_G203_0[0]),.dout(n1375),.clk(gclk));
	jand g1075(.dina(w_n1012_2[2]),.dinb(w_G173_0[0]),.dout(n1376),.clk(gclk));
	jcb g1076(.dina(w_dff_B_HmpjpagX4_0),.dinb(n1375),.dout(n1377));
	jcb g1077(.dina(w_dff_B_DhhOIGEd6_0),.dinb(n1374),.dout(n1378));
	jand g1078(.dina(n1378),.dinb(w_G137_4[2]),.dout(G679),.clk(gclk));
	jand g1079(.dina(w_n1014_2[1]),.dinb(w_G197_0[0]),.dout(n1380),.clk(gclk));
	jand g1080(.dina(w_n1012_2[1]),.dinb(w_G167_0[0]),.dout(n1381),.clk(gclk));
	jcb g1081(.dina(w_dff_B_rEPQrDHN1_0),.dinb(n1380),.dout(n1382));
	jcb g1082(.dina(w_n1213_0[1]),.dinb(w_G1691_2[2]),.dout(n1383));
	jcb g1083(.dina(w_n1251_0[1]),.dinb(w_n1008_2[1]),.dout(n1384));
	jand g1084(.dina(n1384),.dinb(w_dff_B_AyFQlIRn2_1),.dout(n1385),.clk(gclk));
	jand g1085(.dina(n1385),.dinb(w_n1007_1[2]),.dout(n1386),.clk(gclk));
	jcb g1086(.dina(n1386),.dinb(w_dff_B_Ne8oZc1E3_1),.dout(n1387));
	jand g1087(.dina(n1387),.dinb(w_G137_4[1]),.dout(G682),.clk(gclk));
	jcb g1088(.dina(w_n1205_0[1]),.dinb(w_G1691_2[1]),.dout(n1389));
	jcb g1089(.dina(w_n1279_0[1]),.dinb(w_n1008_2[0]),.dout(n1390));
	jand g1090(.dina(n1390),.dinb(w_n1007_1[1]),.dout(n1391),.clk(gclk));
	jand g1091(.dina(n1391),.dinb(w_dff_B_5vZSiFMv0_1),.dout(n1392),.clk(gclk));
	jand g1092(.dina(w_n1014_2[0]),.dinb(w_G194_0[0]),.dout(n1393),.clk(gclk));
	jand g1093(.dina(w_n1012_2[0]),.dinb(w_G164_0[0]),.dout(n1394),.clk(gclk));
	jcb g1094(.dina(w_dff_B_bTO4pNdS5_0),.dinb(n1393),.dout(n1395));
	jcb g1095(.dina(w_dff_B_z6GN4o6J4_0),.dinb(n1392),.dout(n1396));
	jand g1096(.dina(n1396),.dinb(w_G137_4[0]),.dout(G685),.clk(gclk));
	jcb g1097(.dina(w_n1236_0[1]),.dinb(w_n1008_1[2]),.dout(n1398));
	jcb g1098(.dina(w_n1196_0[1]),.dinb(w_G1691_2[0]),.dout(n1399));
	jand g1099(.dina(n1399),.dinb(w_n1007_1[0]),.dout(n1400),.clk(gclk));
	jand g1100(.dina(w_dff_B_19CUk0R73_0),.dinb(n1398),.dout(n1401),.clk(gclk));
	jand g1101(.dina(w_n1014_1[2]),.dinb(w_G191_0[0]),.dout(n1402),.clk(gclk));
	jand g1102(.dina(w_n1012_1[2]),.dinb(w_G161_0[0]),.dout(n1403),.clk(gclk));
	jcb g1103(.dina(w_dff_B_qJoWdEf78_0),.dinb(n1402),.dout(n1404));
	jcb g1104(.dina(w_dff_B_CLCqBe9Z7_0),.dinb(n1401),.dout(n1405));
	jand g1105(.dina(n1405),.dinb(w_G137_3[2]),.dout(G688),.clk(gclk));
	jand g1106(.dina(w_n746_0[0]),.dinb(w_n648_0[2]),.dout(n1407),.clk(gclk));
	jxor g1107(.dina(w_n977_0[0]),.dinb(w_n654_1[0]),.dout(n1408),.clk(gclk));
	jxor g1108(.dina(n1408),.dinb(w_n644_0[0]),.dout(n1409),.clk(gclk));
	jxor g1109(.dina(w_dff_B_1pkzOlgn8_0),.dinb(n1407),.dout(n1410),.clk(gclk));
	jcb g1110(.dina(w_n1410_0[2]),.dinb(w_n737_0[2]),.dout(n1411));
	jnot g1111(.din(w_G2174_0[2]),.dout(n1412),.clk(gclk));
	jnot g1112(.din(w_n719_0[0]),.dout(n1413),.clk(gclk));
	jnot g1113(.din(w_n720_0[0]),.dout(n1414),.clk(gclk));
	jcb g1114(.dina(w_n821_0[0]),.dinb(n1414),.dout(n1415));
	jand g1115(.dina(w_dff_B_X0R6Lci53_0),.dinb(n1413),.dout(n1416),.clk(gclk));
	jxor g1116(.dina(w_n742_0[0]),.dinb(w_n654_0[2]),.dout(n1417),.clk(gclk));
	jxor g1117(.dina(n1417),.dinb(w_n792_0[0]),.dout(n1418),.clk(gclk));
	jnot g1118(.din(w_n660_0[1]),.dout(n1419),.clk(gclk));
	jand g1119(.dina(w_n745_0[0]),.dinb(w_n648_0[1]),.dout(n1420),.clk(gclk));
	jand g1120(.dina(n1420),.dinb(w_dff_B_zsdy9Zl82_1),.dout(n1421),.clk(gclk));
	jxor g1121(.dina(n1421),.dinb(w_dff_B_eNGpBWf86_1),.dout(n1422),.clk(gclk));
	jcb g1122(.dina(w_n1422_0[1]),.dinb(w_n1416_0[1]),.dout(n1423));
	jand g1123(.dina(n1423),.dinb(w_n1412_0[2]),.dout(n1424),.clk(gclk));
	jand g1124(.dina(n1424),.dinb(w_dff_B_xUii6bHv2_1),.dout(n1425),.clk(gclk));
	jnot g1125(.din(w_n1425_0[1]),.dout(n1426),.clk(gclk));
	jnot g1126(.din(w_n641_1[0]),.dout(n1427),.clk(gclk));
	jand g1127(.dina(w_n1416_0[0]),.dinb(n1427),.dout(n1428),.clk(gclk));
	jcb g1128(.dina(w_n1428_0[1]),.dinb(w_n1422_0[0]),.dout(n1429));
	jnot g1129(.din(w_n1429_0[1]),.dout(n1430),.clk(gclk));
	jnot g1130(.din(w_n1410_0[1]),.dout(n1431),.clk(gclk));
	jand g1131(.dina(w_n1428_0[0]),.dinb(n1431),.dout(n1432),.clk(gclk));
	jcb g1132(.dina(n1432),.dinb(w_n1412_0[1]),.dout(n1433));
	jcb g1133(.dina(n1433),.dinb(w_dff_B_d3LsgjpI8_1),.dout(n1434));
	jand g1134(.dina(w_dff_B_8e85yDFP6_0),.dinb(n1426),.dout(n1435),.clk(gclk));
	jcb g1135(.dina(w_n728_0[0]),.dinb(w_n637_0[0]),.dout(n1436));
	jxor g1136(.dina(w_dff_B_fdGNECGl8_0),.dinb(w_n733_0[1]),.dout(n1437),.clk(gclk));
	jxor g1137(.dina(n1437),.dinb(w_n735_0[1]),.dout(n1438),.clk(gclk));
	jcb g1138(.dina(n1438),.dinb(w_G2174_0[1]),.dout(n1439));
	jcb g1139(.dina(w_n735_0[0]),.dinb(w_n640_0[0]),.dout(n1440));
	jcb g1140(.dina(w_n819_0[0]),.dinb(w_n628_0[0]),.dout(n1441));
	jcb g1141(.dina(w_n733_0[0]),.dinb(w_n814_0[0]),.dout(n1442));
	jcb g1142(.dina(w_dff_B_5mPxYXIv3_0),.dinb(w_n639_0[0]),.dout(n1443));
	jand g1143(.dina(n1443),.dinb(w_dff_B_ZUAYicvz0_1),.dout(n1444),.clk(gclk));
	jxor g1144(.dina(n1444),.dinb(n1440),.dout(n1445),.clk(gclk));
	jcb g1145(.dina(n1445),.dinb(w_n1412_0[0]),.dout(n1446));
	jand g1146(.dina(n1446),.dinb(w_dff_B_T3sxnq1M5_1),.dout(n1447),.clk(gclk));
	jxor g1147(.dina(w_n620_0[1]),.dinb(w_n618_0[0]),.dout(n1448),.clk(gclk));
	jxor g1148(.dina(w_n767_0[0]),.dinb(w_n624_0[0]),.dout(n1449),.clk(gclk));
	jxor g1149(.dina(n1449),.dinb(w_dff_B_pVM2lMhF9_1),.dout(n1450),.clk(gclk));
	jxor g1150(.dina(w_dff_B_V58b9dXk3_0),.dinb(n1447),.dout(n1451),.clk(gclk));
	jnot g1151(.din(w_n1451_0[1]),.dout(n1452),.clk(gclk));
	jand g1152(.dina(w_dff_B_Jh3TekGu0_0),.dinb(n1435),.dout(n1453),.clk(gclk));
	jcb g1153(.dina(w_n737_0[1]),.dinb(w_n641_0[2]),.dout(n1454));
	jcb g1154(.dina(w_dff_B_OzS5BOtS0_0),.dinb(w_n1410_0[0]),.dout(n1455));
	jand g1155(.dina(n1455),.dinb(w_G2174_0[0]),.dout(n1456),.clk(gclk));
	jand g1156(.dina(n1456),.dinb(w_n1429_0[0]),.dout(n1457),.clk(gclk));
	jcb g1157(.dina(n1457),.dinb(w_n1425_0[0]),.dout(n1458));
	jand g1158(.dina(w_n1451_0[0]),.dinb(n1458),.dout(n1459),.clk(gclk));
	jcb g1159(.dina(n1459),.dinb(w_n749_5[1]),.dout(n1460));
	jcb g1160(.dina(w_dff_B_a3QL1NSg6_0),.dinb(n1453),.dout(n1461));
	jand g1161(.dina(w_G351_1[0]),.dinb(w_G248_4[1]),.dout(n1462),.clk(gclk));
	jand g1162(.dina(w_n374_0[2]),.dinb(w_G251_4[0]),.dout(n1463),.clk(gclk));
	jcb g1163(.dina(n1463),.dinb(w_n377_0[1]),.dout(n1464));
	jcb g1164(.dina(n1464),.dinb(w_dff_B_rGnss2399_1),.dout(n1465));
	jand g1165(.dina(w_n374_0[1]),.dinb(w_n406_4[0]),.dout(n1466),.clk(gclk));
	jand g1166(.dina(w_G351_0[2]),.dinb(w_n408_4[1]),.dout(n1467),.clk(gclk));
	jcb g1167(.dina(n1467),.dinb(n1466),.dout(n1468));
	jcb g1168(.dina(n1468),.dinb(w_G534_0[2]),.dout(n1469));
	jand g1169(.dina(n1469),.dinb(n1465),.dout(n1470),.clk(gclk));
	jand g1170(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1471),.clk(gclk));
	jand g1171(.dina(w_n387_0[2]),.dinb(w_G251_3[2]),.dout(n1472),.clk(gclk));
	jcb g1172(.dina(n1472),.dinb(w_n389_0[1]),.dout(n1473));
	jcb g1173(.dina(n1473),.dinb(w_dff_B_eZqKCXTv8_1),.dout(n1474));
	jand g1174(.dina(w_n387_0[1]),.dinb(w_n406_3[2]),.dout(n1475),.clk(gclk));
	jand g1175(.dina(w_G341_0[2]),.dinb(w_n408_4[0]),.dout(n1476),.clk(gclk));
	jcb g1176(.dina(n1476),.dinb(n1475),.dout(n1477));
	jcb g1177(.dina(n1477),.dinb(w_G523_0[1]),.dout(n1478));
	jand g1178(.dina(n1478),.dinb(n1474),.dout(n1479),.clk(gclk));
	jxor g1179(.dina(n1479),.dinb(n1470),.dout(n1480),.clk(gclk));
	jcb g1180(.dina(w_n435_1[0]),.dinb(w_n369_1[0]),.dout(n1481));
	jcb g1181(.dina(w_G324_0[2]),.dinb(w_n366_1[0]),.dout(n1482));
	jand g1182(.dina(n1482),.dinb(w_G503_0[2]),.dout(n1483),.clk(gclk));
	jand g1183(.dina(n1483),.dinb(w_dff_B_ojyNWK7c7_1),.dout(n1484),.clk(gclk));
	jcb g1184(.dina(w_G324_0[1]),.dinb(w_G254_1[0]),.dout(n1485));
	jcb g1185(.dina(w_n435_0[2]),.dinb(w_G242_1[0]),.dout(n1486));
	jand g1186(.dina(n1486),.dinb(w_dff_B_UnBdhMhv8_1),.dout(n1487),.clk(gclk));
	jand g1187(.dina(n1487),.dinb(w_n437_0[0]),.dout(n1488),.clk(gclk));
	jcb g1188(.dina(n1488),.dinb(n1484),.dout(n1489));
	jcb g1189(.dina(w_G514_0[2]),.dinb(w_n408_3[2]),.dout(n1490));
	jcb g1190(.dina(w_n361_0[0]),.dinb(w_G248_3[2]),.dout(n1491));
	jand g1191(.dina(n1491),.dinb(n1490),.dout(n1492),.clk(gclk));
	jxor g1192(.dina(n1492),.dinb(w_n371_0[0]),.dout(n1493),.clk(gclk));
	jxor g1193(.dina(n1493),.dinb(n1489),.dout(n1494),.clk(gclk));
	jxor g1194(.dina(n1494),.dinb(n1480),.dout(n1495),.clk(gclk));
	jxor g1195(.dina(w_n433_0[0]),.dinb(w_n428_0[1]),.dout(n1496),.clk(gclk));
	jxor g1196(.dina(w_n423_0[0]),.dinb(w_n412_0[0]),.dout(n1497),.clk(gclk));
	jxor g1197(.dina(n1497),.dinb(n1496),.dout(n1498),.clk(gclk));
	jxor g1198(.dina(n1498),.dinb(n1495),.dout(n1499),.clk(gclk));
	jand g1199(.dina(n1499),.dinb(w_n749_5[0]),.dout(n1500),.clk(gclk));
	jnot g1200(.din(n1500),.dout(n1501),.clk(gclk));
	jand g1201(.dina(w_dff_B_Rqgp33VM1_0),.dinb(n1461),.dout(n1502),.clk(gclk));
	jcb g1202(.dina(n1502),.dinb(w_G4092_4[0]),.dout(n1503));
	jnot g1203(.din(w_n750_2[2]),.dout(n1504),.clk(gclk));
	jcb g1204(.dina(w_n1504_0[1]),.dinb(w_dff_B_azXsQYim8_1),.dout(n1505));
	jand g1205(.dina(w_dff_B_O2wXCame6_0),.dinb(w_n1503_0[1]),.dout(G843),.clk(gclk));
	jand g1206(.dina(w_G273_1[0]),.dinb(w_G248_3[1]),.dout(n1507),.clk(gclk));
	jand g1207(.dina(w_n471_0[2]),.dinb(w_G251_3[1]),.dout(n1508),.clk(gclk));
	jcb g1208(.dina(n1508),.dinb(w_n473_1[0]),.dout(n1509));
	jcb g1209(.dina(n1509),.dinb(w_dff_B_IfxoEAop5_1),.dout(n1510));
	jand g1210(.dina(w_n471_0[1]),.dinb(w_n406_3[1]),.dout(n1511),.clk(gclk));
	jand g1211(.dina(w_G273_0[2]),.dinb(w_n408_3[1]),.dout(n1512),.clk(gclk));
	jcb g1212(.dina(n1512),.dinb(n1511),.dout(n1513));
	jcb g1213(.dina(n1513),.dinb(w_G411_0[2]),.dout(n1514));
	jand g1214(.dina(n1514),.dinb(n1510),.dout(n1515),.clk(gclk));
	jand g1215(.dina(w_G281_1[0]),.dinb(w_G248_3[0]),.dout(n1516),.clk(gclk));
	jand g1216(.dina(w_n530_0[2]),.dinb(w_G251_3[0]),.dout(n1517),.clk(gclk));
	jcb g1217(.dina(n1517),.dinb(w_n532_1[0]),.dout(n1518));
	jcb g1218(.dina(n1518),.dinb(w_dff_B_RfWK9qRM9_1),.dout(n1519));
	jand g1219(.dina(w_n530_0[1]),.dinb(w_n406_3[0]),.dout(n1520),.clk(gclk));
	jand g1220(.dina(w_G281_0[2]),.dinb(w_n408_3[0]),.dout(n1521),.clk(gclk));
	jcb g1221(.dina(n1521),.dinb(n1520),.dout(n1522));
	jcb g1222(.dina(n1522),.dinb(w_G374_0[1]),.dout(n1523));
	jand g1223(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jxor g1224(.dina(n1524),.dinb(n1515),.dout(n1525),.clk(gclk));
	jcb g1225(.dina(w_n483_1[0]),.dinb(w_n369_0[2]),.dout(n1526));
	jcb g1226(.dina(w_G265_0[2]),.dinb(w_n366_0[2]),.dout(n1527));
	jand g1227(.dina(n1527),.dinb(w_G400_0[1]),.dout(n1528),.clk(gclk));
	jand g1228(.dina(n1528),.dinb(w_dff_B_m86AmQ6o9_1),.dout(n1529),.clk(gclk));
	jcb g1229(.dina(w_G265_0[1]),.dinb(w_G254_0[2]),.dout(n1530));
	jcb g1230(.dina(w_n483_0[2]),.dinb(w_G242_0[2]),.dout(n1531));
	jand g1231(.dina(n1531),.dinb(w_dff_B_07KldbNH7_1),.dout(n1532),.clk(gclk));
	jand g1232(.dina(n1532),.dinb(w_n485_0[2]),.dout(n1533),.clk(gclk));
	jcb g1233(.dina(n1533),.dinb(n1529),.dout(n1534));
	jand g1234(.dina(w_G257_1[0]),.dinb(w_G248_2[2]),.dout(n1535),.clk(gclk));
	jand g1235(.dina(w_n518_0[2]),.dinb(w_G251_2[2]),.dout(n1536),.clk(gclk));
	jcb g1236(.dina(n1536),.dinb(w_n520_0[0]),.dout(n1537));
	jcb g1237(.dina(n1537),.dinb(w_dff_B_A039z5SO3_1),.dout(n1538));
	jand g1238(.dina(w_n518_0[1]),.dinb(w_n406_2[2]),.dout(n1539),.clk(gclk));
	jand g1239(.dina(w_G257_0[2]),.dinb(w_n408_2[2]),.dout(n1540),.clk(gclk));
	jcb g1240(.dina(n1540),.dinb(n1539),.dout(n1541));
	jcb g1241(.dina(n1541),.dinb(w_G389_0[1]),.dout(n1542));
	jand g1242(.dina(n1542),.dinb(n1538),.dout(n1543),.clk(gclk));
	jand g1243(.dina(w_G248_2[1]),.dinb(w_G234_1[0]),.dout(n1544),.clk(gclk));
	jand g1244(.dina(w_G251_2[1]),.dinb(w_n460_0[2]),.dout(n1545),.clk(gclk));
	jcb g1245(.dina(n1545),.dinb(w_n462_0[0]),.dout(n1546));
	jcb g1246(.dina(n1546),.dinb(w_dff_B_HSff3Y947_1),.dout(n1547));
	jand g1247(.dina(w_n406_2[1]),.dinb(w_n460_0[1]),.dout(n1548),.clk(gclk));
	jand g1248(.dina(w_n408_2[1]),.dinb(w_G234_0[2]),.dout(n1549),.clk(gclk));
	jcb g1249(.dina(n1549),.dinb(n1548),.dout(n1550));
	jcb g1250(.dina(n1550),.dinb(w_G435_0[1]),.dout(n1551));
	jand g1251(.dina(n1551),.dinb(n1547),.dout(n1552),.clk(gclk));
	jxor g1252(.dina(n1552),.dinb(n1543),.dout(n1553),.clk(gclk));
	jxor g1253(.dina(n1553),.dinb(w_dff_B_DtwF8QNr1_1),.dout(n1554),.clk(gclk));
	jxor g1254(.dina(n1554),.dinb(w_dff_B_Cp9r5I7Y0_1),.dout(n1555),.clk(gclk));
	jand g1255(.dina(w_G248_2[0]),.dinb(w_G226_1[0]),.dout(n1556),.clk(gclk));
	jand g1256(.dina(w_G251_2[0]),.dinb(w_n494_0[2]),.dout(n1557),.clk(gclk));
	jcb g1257(.dina(n1557),.dinb(w_n496_0[1]),.dout(n1558));
	jcb g1258(.dina(n1558),.dinb(w_dff_B_DrhtTbPM2_1),.dout(n1559));
	jand g1259(.dina(w_n406_2[0]),.dinb(w_n494_0[1]),.dout(n1560),.clk(gclk));
	jand g1260(.dina(w_n408_2[0]),.dinb(w_G226_0[2]),.dout(n1561),.clk(gclk));
	jcb g1261(.dina(n1561),.dinb(n1560),.dout(n1562));
	jcb g1262(.dina(n1562),.dinb(w_G422_0[1]),.dout(n1563));
	jand g1263(.dina(n1563),.dinb(n1559),.dout(n1564),.clk(gclk));
	jxor g1264(.dina(n1564),.dinb(w_n551_0[0]),.dout(n1565),.clk(gclk));
	jcb g1265(.dina(w_n369_0[1]),.dinb(w_n507_0[2]),.dout(n1566));
	jcb g1266(.dina(w_n366_0[1]),.dinb(w_G218_1[0]),.dout(n1567));
	jand g1267(.dina(n1567),.dinb(w_G468_0[1]),.dout(n1568),.clk(gclk));
	jand g1268(.dina(n1568),.dinb(w_dff_B_9sfsuSSR1_1),.dout(n1569),.clk(gclk));
	jcb g1269(.dina(w_G254_0[1]),.dinb(w_G218_0[2]),.dout(n1570));
	jcb g1270(.dina(w_G242_0[1]),.dinb(w_n507_0[1]),.dout(n1571));
	jand g1271(.dina(n1571),.dinb(w_dff_B_RYzTC9Qw3_1),.dout(n1572),.clk(gclk));
	jand g1272(.dina(n1572),.dinb(w_n509_0[0]),.dout(n1573),.clk(gclk));
	jcb g1273(.dina(n1573),.dinb(n1569),.dout(n1574));
	jand g1274(.dina(w_G248_1[2]),.dinb(w_G210_1[0]),.dout(n1575),.clk(gclk));
	jand g1275(.dina(w_G251_1[2]),.dinb(w_n449_0[2]),.dout(n1576),.clk(gclk));
	jcb g1276(.dina(n1576),.dinb(w_n451_0[0]),.dout(n1577));
	jcb g1277(.dina(n1577),.dinb(w_dff_B_8xCPJpTY7_1),.dout(n1578));
	jand g1278(.dina(w_n406_1[2]),.dinb(w_n449_0[1]),.dout(n1579),.clk(gclk));
	jand g1279(.dina(w_n408_1[2]),.dinb(w_G210_0[2]),.dout(n1580),.clk(gclk));
	jcb g1280(.dina(n1580),.dinb(n1579),.dout(n1581));
	jcb g1281(.dina(n1581),.dinb(w_G457_0[1]),.dout(n1582));
	jand g1282(.dina(n1582),.dinb(n1578),.dout(n1583),.clk(gclk));
	jxor g1283(.dina(n1583),.dinb(n1574),.dout(n1584),.clk(gclk));
	jxor g1284(.dina(n1584),.dinb(n1565),.dout(n1585),.clk(gclk));
	jxor g1285(.dina(w_dff_B_OaFX81gL2_0),.dinb(n1555),.dout(n1586),.clk(gclk));
	jand g1286(.dina(n1586),.dinb(w_n749_4[2]),.dout(n1587),.clk(gclk));
	jnot g1287(.din(n1587),.dout(n1588),.clk(gclk));
	jand g1288(.dina(w_n573_0[0]),.dinb(w_n567_0[0]),.dout(n1589),.clk(gclk));
	jcb g1289(.dina(n1589),.dinb(w_n699_0[0]),.dout(n1590));
	jnot g1290(.din(w_n559_0[0]),.dout(n1591),.clk(gclk));
	jcb g1291(.dina(n1591),.dinb(w_n557_0[0]),.dout(n1592));
	jand g1292(.dina(w_n1592_0[1]),.dinb(w_n532_0[2]),.dout(n1593),.clk(gclk));
	jnot g1293(.din(w_n1593_0[1]),.dout(n1594),.clk(gclk));
	jcb g1294(.dina(w_n695_0[0]),.dinb(w_dff_B_uCsSlT233_1),.dout(n1595));
	jand g1295(.dina(w_n923_0[1]),.dinb(w_n473_0[2]),.dout(n1596),.clk(gclk));
	jcb g1296(.dina(w_n1596_0[1]),.dinb(w_n1593_0[0]),.dout(n1597));
	jand g1297(.dina(w_dff_B_P5UkVFyp5_0),.dinb(n1595),.dout(n1598),.clk(gclk));
	jxor g1298(.dina(w_dff_B_SVP5Y5N34_0),.dinb(n1590),.dout(n1599),.clk(gclk));
	jnot g1299(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jnot g1300(.din(w_n686_0[0]),.dout(n1601),.clk(gclk));
	jnot g1301(.din(w_n687_0[0]),.dout(n1602),.clk(gclk));
	jcb g1302(.dina(w_n1592_0[0]),.dinb(w_n532_0[1]),.dout(n1603));
	jcb g1303(.dina(w_n1596_0[0]),.dinb(w_n1603_0[1]),.dout(n1604));
	jcb g1304(.dina(w_n923_0[0]),.dinb(w_n473_0[1]),.dout(n1605));
	jcb g1305(.dina(w_n689_0[0]),.dinb(w_n485_0[1]),.dout(n1606));
	jand g1306(.dina(n1606),.dinb(w_n1605_0[1]),.dout(n1607),.clk(gclk));
	jand g1307(.dina(n1607),.dinb(n1604),.dout(n1608),.clk(gclk));
	jcb g1308(.dina(n1608),.dinb(w_n690_0[0]),.dout(n1609));
	jcb g1309(.dina(w_n1609_0[1]),.dinb(n1602),.dout(n1610));
	jand g1310(.dina(w_dff_B_U8dG6jcS2_0),.dinb(n1601),.dout(n1611),.clk(gclk));
	jand g1311(.dina(w_n1611_0[2]),.dinb(w_n581_0[0]),.dout(n1612),.clk(gclk));
	jxor g1312(.dina(w_n566_0[0]),.dinb(w_n561_0[1]),.dout(n1613),.clk(gclk));
	jxor g1313(.dina(w_n1613_0[1]),.dinb(w_n865_0[1]),.dout(n1614),.clk(gclk));
	jxor g1314(.dina(w_dff_B_rXtbchKY7_0),.dinb(n1612),.dout(n1615),.clk(gclk));
	jnot g1315(.din(w_n1615_0[1]),.dout(n1616),.clk(gclk));
	jand g1316(.dina(n1616),.dinb(w_dff_B_sOIUIeEh4_1),.dout(n1617),.clk(gclk));
	jnot g1317(.din(w_G1497_0[2]),.dout(n1618),.clk(gclk));
	jand g1318(.dina(w_n1615_0[0]),.dinb(w_n1599_0[0]),.dout(n1619),.clk(gclk));
	jcb g1319(.dina(n1619),.dinb(w_n1618_0[1]),.dout(n1620));
	jcb g1320(.dina(w_dff_B_a5rfNWOn7_0),.dinb(n1617),.dout(n1621));
	jand g1321(.dina(w_n1605_0[0]),.dinb(w_n1603_0[0]),.dout(n1622),.clk(gclk));
	jcb g1322(.dina(w_dff_B_as1BGSdU2_0),.dinb(w_n694_0[0]),.dout(n1623));
	jxor g1323(.dina(w_n1613_0[0]),.dinb(w_n1609_0[0]),.dout(n1624),.clk(gclk));
	jxor g1324(.dina(n1624),.dinb(w_dff_B_o79XuoKI2_1),.dout(n1625),.clk(gclk));
	jxor g1325(.dina(w_n1611_0[1]),.dinb(w_n865_0[0]),.dout(n1626),.clk(gclk));
	jxor g1326(.dina(n1626),.dinb(n1625),.dout(n1627),.clk(gclk));
	jcb g1327(.dina(n1627),.dinb(w_G1497_0[1]),.dout(n1628));
	jand g1328(.dina(w_dff_B_0cOJAhcX5_0),.dinb(n1621),.dout(n1629),.clk(gclk));
	jxor g1329(.dina(w_n579_0[1]),.dinb(w_n574_0[0]),.dout(n1630),.clk(gclk));
	jxor g1330(.dina(w_dff_B_MIfKNEgW7_0),.dinb(n1629),.dout(n1631),.clk(gclk));
	jnot g1331(.din(w_n709_0[0]),.dout(n1632),.clk(gclk));
	jand g1332(.dina(n1632),.dinb(w_n953_0[0]),.dout(n1633),.clk(gclk));
	jand g1333(.dina(w_n711_0[0]),.dinb(w_n954_0[1]),.dout(n1634),.clk(gclk));
	jcb g1334(.dina(n1634),.dinb(w_n1633_0[1]),.dout(n1635));
	jxor g1335(.dina(w_n608_0[0]),.dinb(w_n592_0[0]),.dout(n1636),.clk(gclk));
	jxor g1336(.dina(n1636),.dinb(w_n602_0[0]),.dout(n1637),.clk(gclk));
	jxor g1337(.dina(w_n1637_0[1]),.dinb(n1635),.dout(n1638),.clk(gclk));
	jcb g1338(.dina(w_n938_0[1]),.dinb(w_n597_0[0]),.dout(n1639));
	jand g1339(.dina(w_n609_0[0]),.dinb(w_n962_0[0]),.dout(n1640),.clk(gclk));
	jcb g1340(.dina(n1640),.dinb(w_n715_0[0]),.dout(n1641));
	jand g1341(.dina(w_dff_B_pk3vYg6W7_0),.dinb(n1639),.dout(n1642),.clk(gclk));
	jxor g1342(.dina(n1642),.dinb(n1638),.dout(n1643),.clk(gclk));
	jand g1343(.dina(w_n1643_0[1]),.dinb(w_n703_0[1]),.dout(n1644),.clk(gclk));
	jnot g1344(.din(w_n682_0[0]),.dout(n1645),.clk(gclk));
	jcb g1345(.dina(w_n1611_0[0]),.dinb(w_n684_0[0]),.dout(n1646));
	jand g1346(.dina(n1646),.dinb(w_dff_B_L5oVnzO48_1),.dout(n1647),.clk(gclk));
	jand g1347(.dina(w_n713_0[0]),.dinb(w_n954_0[0]),.dout(n1648),.clk(gclk));
	jcb g1348(.dina(n1648),.dinb(w_n1633_0[0]),.dout(n1649));
	jxor g1349(.dina(n1649),.dinb(w_n938_0[0]),.dout(n1650),.clk(gclk));
	jxor g1350(.dina(n1650),.dinb(w_n1637_0[0]),.dout(n1651),.clk(gclk));
	jand g1351(.dina(n1651),.dinb(w_dff_B_KVxKDGVU1_1),.dout(n1652),.clk(gclk));
	jcb g1352(.dina(w_n1652_0[1]),.dinb(n1644),.dout(n1653));
	jcb g1353(.dina(n1653),.dinb(w_G1497_0[0]),.dout(n1654));
	jnot g1354(.din(w_n588_1[0]),.dout(n1655),.clk(gclk));
	jand g1355(.dina(w_n1652_0[0]),.dinb(w_dff_B_ptrbJwoT9_1),.dout(n1656),.clk(gclk));
	jcb g1356(.dina(w_n703_0[0]),.dinb(w_n588_0[2]),.dout(n1657));
	jand g1357(.dina(w_dff_B_umz6snDn7_0),.dinb(w_n1643_0[0]),.dout(n1658),.clk(gclk));
	jcb g1358(.dina(w_dff_B_1WUmjhl90_0),.dinb(n1656),.dout(n1659));
	jcb g1359(.dina(n1659),.dinb(w_n1618_0[0]),.dout(n1660));
	jand g1360(.dina(n1660),.dinb(w_dff_B_PYbTzFi39_1),.dout(n1661),.clk(gclk));
	jxor g1361(.dina(n1661),.dinb(n1631),.dout(n1662),.clk(gclk));
	jcb g1362(.dina(n1662),.dinb(w_n749_4[1]),.dout(n1663));
	jand g1363(.dina(n1663),.dinb(w_dff_B_o5Sivf2n5_1),.dout(n1664),.clk(gclk));
	jcb g1364(.dina(n1664),.dinb(w_G4092_3[2]),.dout(n1665));
	jcb g1365(.dina(w_n1504_0[0]),.dinb(w_dff_B_3I40ZzvN4_1),.dout(n1666));
	jand g1366(.dina(w_dff_B_aPJmDf3D1_0),.dinb(w_n1665_0[1]),.dout(G882),.clk(gclk));
	jcb g1367(.dina(w_G4088_3[1]),.dinb(w_G14_0[1]),.dout(n1668));
	jcb g1368(.dina(w_n797_3[1]),.dinb(w_G64_0[1]),.dout(n1669));
	jand g1369(.dina(n1669),.dinb(w_G4087_1[1]),.dout(n1670),.clk(gclk));
	jand g1370(.dina(n1670),.dinb(w_dff_B_gqy9HQBB1_1),.dout(n1671),.clk(gclk));
	jand g1371(.dina(w_G4092_3[1]),.dinb(G97),.dout(n1672),.clk(gclk));
	jnot g1372(.din(n1672),.dout(n1673),.clk(gclk));
	jand g1373(.dina(w_dff_B_ytyy4KYs9_0),.dinb(w_n1665_0[0]),.dout(n1674),.clk(gclk));
	jnot g1374(.din(w_n1674_0[2]),.dout(n1675),.clk(gclk));
	jcb g1375(.dina(w_n1675_0[1]),.dinb(w_n797_3[0]),.dout(n1676));
	jand g1376(.dina(w_G4092_3[0]),.dinb(G94),.dout(n1677),.clk(gclk));
	jnot g1377(.din(n1677),.dout(n1678),.clk(gclk));
	jand g1378(.dina(w_dff_B_LR7OJ1I74_0),.dinb(w_n1503_0[0]),.dout(n1679),.clk(gclk));
	jnot g1379(.din(w_n1679_0[2]),.dout(n1680),.clk(gclk));
	jcb g1380(.dina(w_n1680_0[1]),.dinb(w_G4088_3[0]),.dout(n1681));
	jand g1381(.dina(n1681),.dinb(w_n800_1[1]),.dout(n1682),.clk(gclk));
	jand g1382(.dina(n1682),.dinb(w_dff_B_eFyZ6tLA9_1),.dout(n1683),.clk(gclk));
	jcb g1383(.dina(n1683),.dinb(w_dff_B_WSmL8jgO8_1),.dout(G767));
	jcb g1384(.dina(w_G4089_3[1]),.dinb(w_G14_0[0]),.dout(n1685));
	jcb g1385(.dina(w_n852_3[1]),.dinb(w_G64_0[0]),.dout(n1686));
	jand g1386(.dina(n1686),.dinb(w_G4090_1[1]),.dout(n1687),.clk(gclk));
	jand g1387(.dina(n1687),.dinb(w_dff_B_pkcCmuYD8_1),.dout(n1688),.clk(gclk));
	jcb g1388(.dina(w_n1675_0[0]),.dinb(w_n852_3[0]),.dout(n1689));
	jcb g1389(.dina(w_n1680_0[0]),.dinb(w_G4089_3[0]),.dout(n1690));
	jand g1390(.dina(n1690),.dinb(w_n854_1[1]),.dout(n1691),.clk(gclk));
	jand g1391(.dina(n1691),.dinb(w_dff_B_0X0GAI739_1),.dout(n1692),.clk(gclk));
	jcb g1392(.dina(n1692),.dinb(w_dff_B_bGSCQJIQ0_1),.dout(G807));
	jnot g1393(.din(w_G137_3[1]),.dout(n1694),.clk(gclk));
	jnot g1394(.din(G179),.dout(n1695),.clk(gclk));
	jnot g1395(.din(w_n996_1[1]),.dout(n1696),.clk(gclk));
	jcb g1396(.dina(n1696),.dinb(w_n1695_0[1]),.dout(n1697));
	jnot g1397(.din(G176),.dout(n1698),.clk(gclk));
	jnot g1398(.din(w_n994_1[1]),.dout(n1699),.clk(gclk));
	jcb g1399(.dina(n1699),.dinb(w_n1698_0[1]),.dout(n1700));
	jand g1400(.dina(w_n1674_0[1]),.dinb(w_G1689_1[2]),.dout(n1701),.clk(gclk));
	jand g1401(.dina(w_n1679_0[1]),.dinb(w_n993_1[1]),.dout(n1702),.clk(gclk));
	jcb g1402(.dina(n1702),.dinb(w_G1690_0[1]),.dout(n1703));
	jcb g1403(.dina(n1703),.dinb(w_dff_B_EMUBajAW9_1),.dout(n1704));
	jand g1404(.dina(n1704),.dinb(w_dff_B_nvqN5uz61_1),.dout(n1705),.clk(gclk));
	jand g1405(.dina(n1705),.dinb(w_dff_B_qEMVhYvC0_1),.dout(n1706),.clk(gclk));
	jcb g1406(.dina(n1706),.dinb(w_n1694_0[1]),.dout(G658));
	jnot g1407(.din(w_n1012_1[1]),.dout(n1708),.clk(gclk));
	jcb g1408(.dina(n1708),.dinb(w_n1695_0[0]),.dout(n1709));
	jnot g1409(.din(w_n1014_1[1]),.dout(n1710),.clk(gclk));
	jcb g1410(.dina(n1710),.dinb(w_n1698_0[0]),.dout(n1711));
	jand g1411(.dina(w_n1674_0[0]),.dinb(w_G1691_1[2]),.dout(n1712),.clk(gclk));
	jand g1412(.dina(w_n1679_0[0]),.dinb(w_n1008_1[1]),.dout(n1713),.clk(gclk));
	jcb g1413(.dina(n1713),.dinb(w_G1694_0[1]),.dout(n1714));
	jcb g1414(.dina(n1714),.dinb(w_dff_B_hGr6wSUJ7_1),.dout(n1715));
	jand g1415(.dina(n1715),.dinb(w_dff_B_u18zMVPH2_1),.dout(n1716),.clk(gclk));
	jand g1416(.dina(n1716),.dinb(w_dff_B_O7Z1AKZ68_1),.dout(n1717),.clk(gclk));
	jcb g1417(.dina(n1717),.dinb(w_n1694_0[0]),.dout(G690));
	jdff g1418(.din(w_G141_1[0]),.dout(G144));
	jdff g1419(.din(w_G293_0[0]),.dout(G298));
	jdff g1420(.din(w_G3173_0[0]),.dout(G973));
	jnot g1421(.din(w_G545_0[1]),.dout(G603),.clk(gclk));
	jnot g1422(.din(w_G545_0[0]),.dout(G604),.clk(gclk));
	jdff g1423(.din(w_G137_3[0]),.dout(G926));
	jdff g1424(.din(w_G141_0[2]),.dout(G923));
	jdff g1425(.din(w_G1_2[0]),.dout(G921));
	jdff g1426(.din(w_G549_0[1]),.dout(G892));
	jdff g1427(.din(w_G299_0[1]),.dout(G887));
	jnot g1428(.din(w_G549_0[0]),.dout(G606),.clk(gclk));
	jdff g1429(.din(w_G1_1[2]),.dout(G993));
	jdff g1430(.din(w_G1_1[1]),.dout(G978));
	jdff g1431(.din(w_G1_1[0]),.dout(G949));
	jdff g1432(.din(w_G1_0[2]),.dout(G939));
	jdff g1433(.din(w_G299_0[0]),.dout(G889));
	jcb g1434(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(G717));
	jand g1435(.dina(w_n661_0[0]),.dinb(w_n641_0[1]),.dout(G626),.clk(gclk));
	jand g1436(.dina(w_n611_0[0]),.dinb(w_n588_0[1]),.dout(G632),.clk(gclk));
	jcb g1437(.dina(w_n717_0[0]),.dinb(w_n704_0[0]),.dout(G621));
	jcb g1438(.dina(w_n747_0[0]),.dinb(w_n738_0[0]),.dout(G629));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_FvxgaWv24_1),.doutc(w_G4_0[2]),.din(w_dff_B_DAGiszlx7_3));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(G11));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(G14));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_sd2ZVu9e6_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_im5dFBrE5_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_ukQxG9DW5_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_wGJVb2R39_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(G43));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(G46));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_FAo4GoRd6_2));
	jspl3 jspl3_w_G54_0(.douta(w_dff_A_YzfQGdLU0_0),.doutb(w_dff_A_PcRgOJNS6_1),.doutc(w_G54_0[2]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_nUPCiQug9_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_FLJVpyGZ3_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(G67));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_tQUug1ty3_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(G73));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(G76));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(G91));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(G100));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_HxTIoVvv0_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_Ys6cIc8n8_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(G109));
	jspl jspl_w_G123_0(.douta(w_dff_A_ySZyEEnd2_0),.doutb(w_G123_0[1]),.din(G123));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_QLuiCQ632_0),.doutb(w_dff_A_eQi5s9X70_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_uT9IiILD1_0),.doutb(w_dff_A_aLRzdaaN3_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_nslVg6tw9_0),.doutb(w_dff_A_qWjcXWzl4_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_ODBhPCbc7_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_LgkekKzh6_0),.doutb(w_G137_4[1]),.doutc(w_dff_A_EMhafzSt0_2),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_nbfowXPv7_0),.doutb(w_dff_A_Gr1OsUZM4_1),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_rdQSBNhP1_0),.doutb(w_dff_A_ZlA3nojh2_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_ZkMZMwwK5_1),.doutc(w_dff_A_LHfbv8a61_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_dff_A_mbCLFJ1C0_0),.doutb(w_G137_8[1]),.doutc(w_dff_A_3m7ZcVHv3_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_dff_A_vkfbRAzT5_0),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_URWs1D7U2_1),.doutc(w_dff_A_U92YXMBk7_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_ntJFtxVS6_0),.doutb(w_dff_A_V5xbFpuQ9_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_CUdKH9X76_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_Vtj1ABIZ9_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_QRfzaI208_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_BpTF5GQy4_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_Qku3HVSq6_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_ILB9o4r96_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_Z4HedfuY6_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_xzRqBeyM5_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_fJjEArNj5_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_kl9TYwy45_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_esaDwXgw5_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_menrNAlj4_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_fBz5XXFX2_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_Yf51D3so8_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_0c6JP3fR4_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_LbQbXpqE0_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_P7lro8k06_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_a6wgwdlZ7_2));
	jspl3 jspl3_w_G206_0(.douta(w_G206_0[0]),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G206_1(.douta(w_dff_A_NIY42FNy3_0),.doutb(w_G206_1[1]),.doutc(w_G206_1[2]),.din(w_G206_0[0]));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_eCxoAzf34_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_G210_1[1]),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl jspl_w_G210_2(.douta(w_dff_A_XZylqcdf9_0),.doutb(w_G210_2[1]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_8zdwvfop7_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl jspl_w_G218_2(.douta(w_dff_A_ayZZV8Mh8_0),.doutb(w_G218_2[1]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_dff_A_Hk7IFeeq8_2),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl jspl_w_G226_2(.douta(w_dff_A_hSJTcLhb5_0),.doutb(w_G226_2[1]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_ufYN7Zob3_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_LHGc20gx9_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_eePLoI0R8_1),.doutc(w_dff_A_yHUCZuC37_2),.din(G242));
	jspl jspl_w_G242_1(.douta(w_dff_A_d4OfE2S05_0),.doutb(w_G242_1[1]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_dff_A_G9Pwthw85_0),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_8w6nNEqq5_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl3 jspl3_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.doutc(w_G248_5[2]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_6pD16Eak7_1),.doutc(w_dff_A_TGig5Ra66_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_dff_A_pKnYCdRQ0_0),.doutb(w_G251_1[1]),.doutc(w_dff_A_hnZVdOah8_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_G251_4[1]),.doutc(w_G251_4[2]),.din(w_G251_1[0]));
	jspl jspl_w_G251_5(.douta(w_dff_A_igLneryp8_0),.doutb(w_G251_5[1]),.din(w_G251_1[1]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl jspl_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_dff_A_nUkqtVwk2_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl jspl_w_G257_2(.douta(w_dff_A_bjpd9y5w2_0),.doutb(w_G257_2[1]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_28hBAJIf9_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_dff_A_p5KaWxUz0_1),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_x7sGiAdx3_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_dff_A_6FuuZyO67_1),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl jspl_w_G273_2(.douta(w_dff_A_JXrCIJvl2_0),.doutb(w_G273_2[1]),.din(w_G273_0[1]));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_35IMdrIP4_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_tmfqrQf33_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_G289_0[0]),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_8pzO0rXC3_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_Q6s4J0Ok9_0),.doutb(w_dff_A_NemSBIxA4_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_K26thiWr8_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_dff_A_h3z2YUrv4_2),.din(G316));
	jspl jspl_w_G316_1(.douta(w_G316_1[0]),.doutb(w_G316_1[1]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_G324_0[1]),.doutc(w_dff_A_PD6kO0Ym0_2),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_jOXfclfh5_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_Oz1kqe4N9_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_dff_A_oJvT7yWN6_1),.doutc(w_G332_1[2]),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_AJsusLjk2_0),.doutb(w_G332_2[1]),.doutc(w_dff_A_xm5kZ9st4_2),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_G332_3[0]),.doutb(w_G332_3[1]),.doutc(w_G332_3[2]),.din(w_G332_0[2]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl jspl_w_G338_0(.douta(w_dff_A_LtwD0vNX5_0),.doutb(w_G338_0[1]),.din(G338));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_ppkAAw5J0_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_xQfn7MGY8_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_d0mXA9PV1_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_dff_A_PsHvd5hW2_2),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_G351_1[0]),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_3YLb6Y9c1_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_CLGdv8Ko1_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_G361_0[1]),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G361_1(.douta(w_dff_A_k3JB3iCB9_0),.doutb(w_G361_1[1]),.din(w_G361_0[0]));
	jspl jspl_w_G366_0(.douta(w_dff_A_tUR2AhzW3_0),.doutb(w_G366_0[1]),.din(G366));
	jspl jspl_w_G369_0(.douta(w_G369_0[0]),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_G374_0[0]),.doutb(w_dff_A_N7rosL8O5_1),.doutc(w_dff_A_xG4huGW33_2),.din(G374));
	jspl3 jspl3_w_G374_1(.douta(w_dff_A_iT0XC6JC1_0),.doutb(w_dff_A_AYOFg4f10_1),.doutc(w_G374_1[2]),.din(w_G374_0[0]));
	jspl3 jspl3_w_G389_0(.douta(w_G389_0[0]),.doutb(w_dff_A_KMlWaPwz4_1),.doutc(w_dff_A_04DJAaSG2_2),.din(G389));
	jspl3 jspl3_w_G389_1(.douta(w_dff_A_Sgh0BycS8_0),.doutb(w_dff_A_6XZQcvXs7_1),.doutc(w_G389_1[2]),.din(w_G389_0[0]));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_2ZG2lwal3_1),.doutc(w_dff_A_F0aoAc7Z5_2),.din(G400));
	jspl3 jspl3_w_G400_1(.douta(w_dff_A_ddJZg2O26_0),.doutb(w_dff_A_6PT9UaPV7_1),.doutc(w_G400_1[2]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_cQUuhADp8_0),.doutb(w_G411_0[1]),.doutc(w_dff_A_pMF7ZgcW6_2),.din(G411));
	jspl3 jspl3_w_G411_1(.douta(w_G411_1[0]),.doutb(w_G411_1[1]),.doutc(w_G411_1[2]),.din(w_G411_0[0]));
	jspl jspl_w_G411_2(.douta(w_dff_A_H2IaVxAx0_0),.doutb(w_G411_2[1]),.din(w_G411_0[1]));
	jspl3 jspl3_w_G422_0(.douta(w_G422_0[0]),.doutb(w_dff_A_6QueWslw8_1),.doutc(w_dff_A_OW3w21rU4_2),.din(G422));
	jspl jspl_w_G422_1(.douta(w_dff_A_UaZNyiSJ8_0),.doutb(w_G422_1[1]),.din(w_G422_0[0]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_sleKAM1H8_1),.doutc(w_dff_A_Z4jqWwkk4_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_zI9PDHAN4_0),.doutb(w_dff_A_Vy5T5x4G7_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_0GvYtfUI6_1),.doutc(w_dff_A_8HkfzeEk4_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_PUPbGg4F4_0),.doutb(w_dff_A_tBxglOLO9_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_G457_0[0]),.doutb(w_dff_A_UpmAJVRc9_1),.doutc(w_dff_A_wCHQqrQ66_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_dff_A_29KEvHpM3_0),.doutb(w_dff_A_dVbwrVjr4_1),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_HOf4kQdV8_1),.doutc(w_dff_A_penQLU6r8_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_ewlGzfSJ4_0),.doutb(w_dff_A_SE6sVdrN9_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_dff_A_DybV0qOA6_0),.doutb(w_dff_A_klxydncY7_1),.doutc(w_G479_0[2]),.din(G479));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_1btaIGhu2_1),.doutc(w_dff_A_OezKpDzA1_2),.din(G490));
	jspl jspl_w_G490_1(.douta(w_dff_A_VgQhHTKt5_0),.doutb(w_G490_1[1]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_dff_A_JxeyMOSj2_0),.doutb(w_G503_0[1]),.doutc(w_dff_A_T7tHFmi49_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_G503_1[0]),.doutb(w_G503_1[1]),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl jspl_w_G503_2(.douta(w_dff_A_WA0s8Mnc6_0),.doutb(w_G503_2[1]),.din(w_G503_0[1]));
	jspl3 jspl3_w_G514_0(.douta(w_dff_A_GEsH3DP62_0),.doutb(w_G514_0[1]),.doutc(w_dff_A_p7EyMcTN4_2),.din(G514));
	jspl3 jspl3_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.doutc(w_G514_1[2]),.din(w_G514_0[0]));
	jspl jspl_w_G514_2(.douta(w_G514_2[0]),.doutb(w_G514_2[1]),.din(w_G514_0[1]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_tWoPz4ME8_1),.doutc(w_dff_A_mckreH0L8_2),.din(G523));
	jspl3 jspl3_w_G523_1(.douta(w_dff_A_sHe4h7fx4_0),.doutb(w_dff_A_RZ5VYcc30_1),.doutc(w_G523_1[2]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_dff_A_mDu6K7KB9_0),.doutb(w_G534_0[1]),.doutc(w_dff_A_22TePM3N9_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_G534_1[0]),.doutb(w_G534_1[1]),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl jspl_w_G534_2(.douta(w_dff_A_IFGDUsUK7_0),.doutb(w_G534_2[1]),.din(w_G534_0[1]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_dff_A_5dlESbO32_0),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_K1zS4y1F5_0),.doutb(w_dff_A_ODvgMo6Y2_1),.doutc(w_G1497_0[2]),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_dff_A_QXu7rwtx6_1),.doutc(w_dff_A_vbkxWPKJ6_2),.din(G1689));
	jspl3 jspl3_w_G1689_1(.douta(w_dff_A_yn9tlmaF7_0),.doutb(w_G1689_1[1]),.doutc(w_dff_A_ZGEwQbOp8_2),.din(w_G1689_0[0]));
	jspl3 jspl3_w_G1689_2(.douta(w_dff_A_dbL7HgUb5_0),.doutb(w_dff_A_5gv99wKp5_1),.doutc(w_G1689_2[2]),.din(w_G1689_0[1]));
	jspl3 jspl3_w_G1689_3(.douta(w_dff_A_ub3jo0QX4_0),.doutb(w_dff_A_Z3m41yRD3_1),.doutc(w_G1689_3[2]),.din(w_G1689_0[2]));
	jspl3 jspl3_w_G1689_4(.douta(w_dff_A_wPirhIZM5_0),.doutb(w_dff_A_hU8ufdTl1_1),.doutc(w_G1689_4[2]),.din(w_G1689_1[0]));
	jspl jspl_w_G1689_5(.douta(w_G1689_5[0]),.doutb(w_G1689_5[1]),.din(w_G1689_1[1]));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_f405pS0G7_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl jspl_w_G1690_1(.douta(w_G1690_1[0]),.doutb(w_dff_A_XlDx9OSS6_1),.din(w_G1690_0[0]));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_dff_A_RulbiuaA4_1),.doutc(w_dff_A_4Py8OvaH9_2),.din(G1691));
	jspl3 jspl3_w_G1691_1(.douta(w_G1691_1[0]),.doutb(w_G1691_1[1]),.doutc(w_dff_A_iZXm6Txu5_2),.din(w_G1691_0[0]));
	jspl3 jspl3_w_G1691_2(.douta(w_dff_A_AgVAjbLj8_0),.doutb(w_dff_A_I9Uio7DV6_1),.doutc(w_G1691_2[2]),.din(w_G1691_0[1]));
	jspl3 jspl3_w_G1691_3(.douta(w_dff_A_PoXbhRtG3_0),.doutb(w_dff_A_jsFtZQH11_1),.doutc(w_G1691_3[2]),.din(w_G1691_0[2]));
	jspl3 jspl3_w_G1691_4(.douta(w_dff_A_WEuSM3HY6_0),.doutb(w_dff_A_5oOWpqjS6_1),.doutc(w_G1691_4[2]),.din(w_G1691_1[0]));
	jspl jspl_w_G1691_5(.douta(w_G1691_5[0]),.doutb(w_dff_A_o4grvfCh0_1),.din(w_G1691_1[1]));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_aQCxkdfb3_1),.doutc(w_dff_A_gU3g5sc85_2),.din(G1694));
	jspl jspl_w_G1694_1(.douta(w_G1694_1[0]),.doutb(w_G1694_1[1]),.din(w_G1694_0[0]));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_HftPVBkU4_0),.doutb(w_dff_A_dEf9Dms78_1),.doutc(w_G2174_0[2]),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_wBPBDoQH6_0),.doutb(w_dff_A_kkDkeOtI7_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_dTX8841M8_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_G3724_0[0]),.doutb(w_G3724_0[1]),.doutc(w_dff_A_wwcE1kRT2_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_G4087_0[1]),.doutc(w_G4087_0[2]),.din(G4087));
	jspl3 jspl3_w_G4087_1(.douta(w_G4087_1[0]),.doutb(w_dff_A_ZY4mbvov9_1),.doutc(w_G4087_1[2]),.din(w_G4087_0[0]));
	jspl3 jspl3_w_G4087_2(.douta(w_G4087_2[0]),.doutb(w_G4087_2[1]),.doutc(w_G4087_2[2]),.din(w_G4087_0[1]));
	jspl3 jspl3_w_G4087_3(.douta(w_G4087_3[0]),.doutb(w_G4087_3[1]),.doutc(w_G4087_3[2]),.din(w_G4087_0[2]));
	jspl3 jspl3_w_G4087_4(.douta(w_G4087_4[0]),.doutb(w_G4087_4[1]),.doutc(w_G4087_4[2]),.din(w_G4087_1[0]));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_G4088_0[2]),.din(G4088));
	jspl3 jspl3_w_G4088_1(.douta(w_G4088_1[0]),.doutb(w_G4088_1[1]),.doutc(w_G4088_1[2]),.din(w_G4088_0[0]));
	jspl3 jspl3_w_G4088_2(.douta(w_G4088_2[0]),.doutb(w_G4088_2[1]),.doutc(w_G4088_2[2]),.din(w_G4088_0[1]));
	jspl3 jspl3_w_G4088_3(.douta(w_dff_A_iPVAgh5r5_0),.doutb(w_G4088_3[1]),.doutc(w_G4088_3[2]),.din(w_G4088_0[2]));
	jspl3 jspl3_w_G4088_4(.douta(w_dff_A_GtycS8g76_0),.doutb(w_G4088_4[1]),.doutc(w_dff_A_UR13TOBk4_2),.din(w_G4088_1[0]));
	jspl3 jspl3_w_G4088_5(.douta(w_G4088_5[0]),.doutb(w_dff_A_aBzkJTVZ8_1),.doutc(w_G4088_5[2]),.din(w_G4088_1[1]));
	jspl3 jspl3_w_G4088_6(.douta(w_dff_A_wmvximqy1_0),.doutb(w_G4088_6[1]),.doutc(w_dff_A_aO7SEFju5_2),.din(w_G4088_1[2]));
	jspl3 jspl3_w_G4088_7(.douta(w_G4088_7[0]),.doutb(w_dff_A_LFa27Mez9_1),.doutc(w_G4088_7[2]),.din(w_G4088_2[0]));
	jspl3 jspl3_w_G4088_8(.douta(w_dff_A_ocmlcEj69_0),.doutb(w_G4088_8[1]),.doutc(w_dff_A_LiETSce14_2),.din(w_G4088_2[1]));
	jspl3 jspl3_w_G4088_9(.douta(w_G4088_9[0]),.doutb(w_dff_A_uA12pxJ92_1),.doutc(w_G4088_9[2]),.din(w_G4088_2[2]));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_G4089_0[2]),.din(G4089));
	jspl3 jspl3_w_G4089_1(.douta(w_G4089_1[0]),.doutb(w_G4089_1[1]),.doutc(w_G4089_1[2]),.din(w_G4089_0[0]));
	jspl3 jspl3_w_G4089_2(.douta(w_G4089_2[0]),.doutb(w_G4089_2[1]),.doutc(w_G4089_2[2]),.din(w_G4089_0[1]));
	jspl3 jspl3_w_G4089_3(.douta(w_dff_A_WJPfpayy3_0),.doutb(w_G4089_3[1]),.doutc(w_G4089_3[2]),.din(w_G4089_0[2]));
	jspl3 jspl3_w_G4089_4(.douta(w_dff_A_3Q17h9HF4_0),.doutb(w_G4089_4[1]),.doutc(w_dff_A_KC6qS1y01_2),.din(w_G4089_1[0]));
	jspl3 jspl3_w_G4089_5(.douta(w_G4089_5[0]),.doutb(w_dff_A_QQ3cgWxW8_1),.doutc(w_dff_A_7jshLYJC7_2),.din(w_G4089_1[1]));
	jspl3 jspl3_w_G4089_6(.douta(w_G4089_6[0]),.doutb(w_G4089_6[1]),.doutc(w_dff_A_YrEGUGTu5_2),.din(w_G4089_1[2]));
	jspl3 jspl3_w_G4089_7(.douta(w_dff_A_y3Wiv0ee2_0),.doutb(w_G4089_7[1]),.doutc(w_dff_A_Ydf7G1MN5_2),.din(w_G4089_2[0]));
	jspl3 jspl3_w_G4089_8(.douta(w_G4089_8[0]),.doutb(w_dff_A_a3kVmaUn1_1),.doutc(w_G4089_8[2]),.din(w_G4089_2[1]));
	jspl3 jspl3_w_G4089_9(.douta(w_G4089_9[0]),.doutb(w_dff_A_HgcJxiAs8_1),.doutc(w_G4089_9[2]),.din(w_G4089_2[2]));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_G4090_0[1]),.doutc(w_G4090_0[2]),.din(G4090));
	jspl3 jspl3_w_G4090_1(.douta(w_G4090_1[0]),.doutb(w_dff_A_vnoqIWWT6_1),.doutc(w_G4090_1[2]),.din(w_G4090_0[0]));
	jspl3 jspl3_w_G4090_2(.douta(w_G4090_2[0]),.doutb(w_G4090_2[1]),.doutc(w_dff_A_tSDqlSZB3_2),.din(w_G4090_0[1]));
	jspl3 jspl3_w_G4090_3(.douta(w_G4090_3[0]),.doutb(w_dff_A_nEW9LA4a0_1),.doutc(w_dff_A_POkQJsV80_2),.din(w_G4090_0[2]));
	jspl3 jspl3_w_G4090_4(.douta(w_dff_A_WrtBaxLL7_0),.doutb(w_G4090_4[1]),.doutc(w_G4090_4[2]),.din(w_G4090_1[0]));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_dff_A_mRgHOw5y3_1),.doutc(w_dff_A_uyKqCI4e6_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_dff_A_RKSBBxJA8_0),.doutb(w_dff_A_k5UnAS1S9_1),.doutc(w_G4091_1[2]),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_dff_A_X20EqEFP2_0),.doutb(w_dff_A_WX1kDifk3_1),.doutc(w_G4091_2[2]),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4091_3(.douta(w_G4091_3[0]),.doutb(w_dff_A_9gC8U8aS1_1),.doutc(w_dff_A_VBoCBJqN8_2),.din(w_G4091_0[2]));
	jspl3 jspl3_w_G4091_4(.douta(w_dff_A_smjPFL1o7_0),.doutb(w_G4091_4[1]),.doutc(w_dff_A_rbirpuik2_2),.din(w_G4091_1[0]));
	jspl3 jspl3_w_G4091_5(.douta(w_dff_A_GAPszGMA6_0),.doutb(w_G4091_5[1]),.doutc(w_G4091_5[2]),.din(w_G4091_1[1]));
	jspl jspl_w_G4091_6(.douta(w_dff_A_jgyoAhAo8_0),.doutb(w_G4091_6[1]),.din(w_G4091_1[2]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_dff_A_lcXMExnl1_1),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_0c2haayH0_0),.doutb(w_G4092_1[1]),.doutc(w_dff_A_2xvx20Dz2_2),.din(w_G4092_0[0]));
	jspl3 jspl3_w_G4092_2(.douta(w_dff_A_J7Y9NuWP2_0),.doutb(w_dff_A_RqxKpO2m6_1),.doutc(w_G4092_2[2]),.din(w_G4092_0[1]));
	jspl3 jspl3_w_G4092_3(.douta(w_G4092_3[0]),.doutb(w_G4092_3[1]),.doutc(w_dff_A_CiHQhXAV7_2),.din(w_G4092_0[2]));
	jspl3 jspl3_w_G4092_4(.douta(w_dff_A_bOzkJjjs5_0),.doutb(w_G4092_4[1]),.doutc(w_G4092_4[2]),.din(w_G4092_1[0]));
	jspl3 jspl3_w_G4092_5(.douta(w_dff_A_gJuftH4B6_0),.doutb(w_dff_A_OdaYqszP2_1),.doutc(w_G4092_5[2]),.din(w_G4092_1[1]));
	jspl3 jspl3_w_G4092_6(.douta(w_G4092_6[0]),.doutb(w_dff_A_HIvEGoOw6_1),.doutc(w_dff_A_gsEPuZkl3_2),.din(w_G4092_1[2]));
	jspl3 jspl3_w_G4092_7(.douta(w_G4092_7[0]),.doutb(w_G4092_7[1]),.doutc(w_dff_A_sVMre9Ik6_2),.din(w_G4092_2[0]));
	jspl3 jspl3_w_G4092_8(.douta(w_G4092_8[0]),.doutb(w_G4092_8[1]),.doutc(w_G4092_8[2]),.din(w_G4092_2[1]));
	jspl3 jspl3_w_G4092_9(.douta(w_dff_A_LlDY6nhZ3_0),.doutb(w_dff_A_gmf8R17O2_1),.doutc(w_G4092_9[2]),.din(w_G4092_2[2]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(G599),.din(G599_fa_));
	jspl jspl_w_G601_0(.douta(w_G601_0),.doutb(G601),.din(G601_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(G612),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_dff_A_uOTPqfW57_0),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_dff_A_s5V3QPdz0_2),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_dff_A_9AfsaUq23_0),.doutb(w_G809_3[1]),.doutc(G809),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(G593),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(G822),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(G838),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(G861),.din(G861_fa_));
	jspl jspl_w_G623_0(.douta(w_G623_0),.doutb(G623),.din(G623_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(G832),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(G834),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(G836),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(G871),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(G873),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(G875),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(G877),.din(G877_fa_));
	jspl jspl_w_G998_0(.douta(w_G998_0),.doutb(G998),.din(G998_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(G830),.din(G830_fa_));
	jspl jspl_w_G865_0(.douta(w_G865_0),.doutb(G865),.din(G865_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(G869),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.doutc(w_n369_0[2]),.din(n369));
	jspl3 jspl3_w_n369_1(.douta(w_n369_1[0]),.doutb(w_n369_1[1]),.doutc(w_n369_1[2]),.din(w_n369_0[0]));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.doutc(w_n374_0[2]),.din(n374));
	jspl jspl_w_n374_1(.douta(w_n374_1[0]),.doutb(w_n374_1[1]),.din(w_n374_0[0]));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n375_1(.douta(w_n375_1[0]),.doutb(w_n375_1[1]),.doutc(w_n375_1[2]),.din(w_n375_0[0]));
	jspl3 jspl3_w_n375_2(.douta(w_n375_2[0]),.doutb(w_n375_2[1]),.doutc(w_n375_2[2]),.din(w_n375_0[1]));
	jspl3 jspl3_w_n375_3(.douta(w_n375_3[0]),.doutb(w_n375_3[1]),.doutc(w_n375_3[2]),.din(w_n375_0[2]));
	jspl3 jspl3_w_n375_4(.douta(w_n375_4[0]),.doutb(w_n375_4[1]),.doutc(w_n375_4[2]),.din(w_n375_1[0]));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_n377_0[2]),.din(w_dff_B_V7Kax62f0_3));
	jspl jspl_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.doutc(w_n378_0[2]),.din(n378));
	jspl3 jspl3_w_n378_1(.douta(w_n378_1[0]),.doutb(w_n378_1[1]),.doutc(w_n378_1[2]),.din(w_n378_0[0]));
	jspl3 jspl3_w_n378_2(.douta(w_n378_2[0]),.doutb(w_n378_2[1]),.doutc(w_n378_2[2]),.din(w_n378_0[1]));
	jspl3 jspl3_w_n378_3(.douta(w_n378_3[0]),.doutb(w_n378_3[1]),.doutc(w_n378_3[2]),.din(w_n378_0[2]));
	jspl3 jspl3_w_n378_4(.douta(w_n378_4[0]),.doutb(w_n378_4[1]),.doutc(w_n378_4[2]),.din(w_n378_1[0]));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(w_dff_B_heec8Ysv9_3));
	jspl jspl_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n401_0(.douta(w_dff_A_BCuU1Rr21_0),.doutb(w_n401_0[1]),.din(w_dff_B_znryO9ie9_2));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.doutc(w_n406_0[2]),.din(n406));
	jspl3 jspl3_w_n406_1(.douta(w_n406_1[0]),.doutb(w_n406_1[1]),.doutc(w_n406_1[2]),.din(w_n406_0[0]));
	jspl3 jspl3_w_n406_2(.douta(w_n406_2[0]),.doutb(w_n406_2[1]),.doutc(w_n406_2[2]),.din(w_n406_0[1]));
	jspl3 jspl3_w_n406_3(.douta(w_n406_3[0]),.doutb(w_n406_3[1]),.doutc(w_n406_3[2]),.din(w_n406_0[2]));
	jspl3 jspl3_w_n406_4(.douta(w_n406_4[0]),.doutb(w_n406_4[1]),.doutc(w_n406_4[2]),.din(w_n406_1[0]));
	jspl jspl_w_n406_5(.douta(w_n406_5[0]),.doutb(w_n406_5[1]),.din(w_n406_1[1]));
	jspl3 jspl3_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.doutc(w_n408_0[2]),.din(n408));
	jspl3 jspl3_w_n408_1(.douta(w_n408_1[0]),.doutb(w_n408_1[1]),.doutc(w_n408_1[2]),.din(w_n408_0[0]));
	jspl3 jspl3_w_n408_2(.douta(w_n408_2[0]),.doutb(w_n408_2[1]),.doutc(w_n408_2[2]),.din(w_n408_0[1]));
	jspl3 jspl3_w_n408_3(.douta(w_n408_3[0]),.doutb(w_n408_3[1]),.doutc(w_n408_3[2]),.din(w_n408_0[2]));
	jspl3 jspl3_w_n408_4(.douta(w_n408_4[0]),.doutb(w_n408_4[1]),.doutc(w_n408_4[2]),.din(w_n408_1[0]));
	jspl3 jspl3_w_n408_5(.douta(w_n408_5[0]),.doutb(w_n408_5[1]),.doutc(w_n408_5[2]),.din(w_n408_1[1]));
	jspl3 jspl3_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.doutc(w_n412_0[2]),.din(n412));
	jspl jspl_w_n414_0(.douta(w_dff_A_rJlRsTwe4_0),.doutb(w_n414_0[1]),.din(w_dff_B_7V7pwQqq8_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_dff_A_qS9klzNj2_1),.doutc(w_n428_0[2]),.din(n428));
	jspl jspl_w_n428_1(.douta(w_n428_1[0]),.doutb(w_dff_A_pZ8QkzW89_1),.din(w_n428_0[0]));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_n433_0[2]),.din(n433));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl jspl_w_n435_2(.douta(w_n435_2[0]),.doutb(w_n435_2[1]),.din(w_n435_0[1]));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(w_dff_B_TTFTocGu1_2));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_dff_A_s0mWYLZx6_1),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_dff_A_SrzM1ZCC3_1),.doutc(w_n451_0[2]),.din(w_dff_B_glHv4Be06_3));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_2QrO1eFJ5_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_xoOMif9N4_1),.doutc(w_n462_0[2]),.din(w_dff_B_JkwMTCpa0_3));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl3 jspl3_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.doutc(w_n471_1[2]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_n473_0[2]),.din(w_dff_B_y2eLDWYg9_3));
	jspl jspl_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.doutc(w_n483_0[2]),.din(n483));
	jspl3 jspl3_w_n483_1(.douta(w_n483_1[0]),.doutb(w_n483_1[1]),.doutc(w_n483_1[2]),.din(w_n483_0[0]));
	jspl jspl_w_n483_2(.douta(w_n483_2[0]),.doutb(w_n483_2[1]),.din(w_n483_0[1]));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.doutc(w_n485_0[2]),.din(w_dff_B_dULN66I59_3));
	jspl jspl_w_n485_1(.douta(w_n485_1[0]),.doutb(w_n485_1[1]),.din(w_n485_0[0]));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl3 jspl3_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.doutc(w_n494_0[2]),.din(n494));
	jspl3 jspl3_w_n494_1(.douta(w_n494_1[0]),.doutb(w_n494_1[1]),.doutc(w_n494_1[2]),.din(w_n494_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_dff_A_21qrzfBF6_2),.din(w_dff_B_2Ugq5SDK0_3));
	jspl jspl_w_n496_1(.douta(w_dff_A_uFn72zPK9_0),.doutb(w_n496_1[1]),.din(w_n496_0[0]));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl3 jspl3_w_n509_0(.douta(w_n509_0[0]),.doutb(w_dff_A_ynWu1gvJ3_1),.doutc(w_n509_0[2]),.din(w_dff_B_Jd8Y8iK58_3));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_dff_A_FrwNMP6u2_1),.doutc(w_n520_0[2]),.din(w_dff_B_jUzy2tsp4_3));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl3 jspl3_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.doutc(w_n530_1[2]),.din(w_n530_0[0]));
	jspl3 jspl3_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.doutc(w_n532_0[2]),.din(w_dff_B_dbez48296_3));
	jspl jspl_w_n532_1(.douta(w_n532_1[0]),.doutb(w_n532_1[1]),.din(w_n532_0[0]));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.doutc(w_n551_0[2]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl3 jspl3_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.doutc(w_n556_5[2]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n556_6(.douta(w_n556_6[0]),.doutb(w_n556_6[1]),.doutc(w_n556_6[2]),.din(w_n556_1[2]));
	jspl3 jspl3_w_n556_7(.douta(w_n556_7[0]),.doutb(w_n556_7[1]),.doutc(w_n556_7[2]),.din(w_n556_2[0]));
	jspl jspl_w_n556_8(.douta(w_n556_8[0]),.doutb(w_n556_8[1]),.din(w_n556_2[1]));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_dff_A_SRqVufOq5_1),.din(n559));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.din(w_n561_0[0]));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_wZAo4vm67_1),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.din(n569));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_dff_A_VCHzWWBO2_1),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_dff_A_KiCxKFaz6_0),.doutb(w_dff_A_6zW5vQiK3_1),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_dff_A_AbPZAwis7_1),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl jspl_w_n578_1(.douta(w_n578_1[0]),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_dff_A_KwzCzioj9_1),.doutc(w_dff_A_8m8VzK7g3_2),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_dff_A_n64hHnDN6_1),.din(w_n579_0[0]));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n586_1(.douta(w_n586_1[0]),.doutb(w_n586_1[1]),.din(w_n586_0[0]));
	jspl jspl_w_n587_0(.douta(w_n587_0[0]),.doutb(w_dff_A_gspL3bJU9_1),.din(n587));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.doutc(w_n591_0[2]),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_uX3tdavN5_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_cCq4LzdO9_2),.din(n592));
	jspl3 jspl3_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl jspl_w_n596_1(.douta(w_n596_1[0]),.doutb(w_n596_1[1]),.din(w_n596_0[0]));
	jspl3 jspl3_w_n597_0(.douta(w_dff_A_c8BxFHsH8_0),.doutb(w_n597_0[1]),.doutc(w_n597_0[2]),.din(n597));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n601_1(.douta(w_n601_1[0]),.doutb(w_n601_1[1]),.din(w_n601_0[0]));
	jspl3 jspl3_w_n602_0(.douta(w_dff_A_5gwSCMZM8_0),.doutb(w_n602_0[1]),.doutc(w_n602_0[2]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n607_1(.douta(w_n607_1[0]),.doutb(w_n607_1[1]),.din(w_n607_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_L4AHDBsg0_1),.doutc(w_n608_0[2]),.din(n608));
	jspl3 jspl3_w_n609_0(.douta(w_dff_A_duw3mAMP8_0),.doutb(w_dff_A_hpqvISpo6_1),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n611_0(.douta(w_n611_0[0]),.doutb(w_n611_0[1]),.doutc(w_n611_0[2]),.din(w_dff_B_xQTz6HIA3_3));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n613_2(.douta(w_n613_2[0]),.doutb(w_n613_2[1]),.doutc(w_n613_2[2]),.din(w_n613_0[1]));
	jspl3 jspl3_w_n613_3(.douta(w_n613_3[0]),.doutb(w_n613_3[1]),.doutc(w_n613_3[2]),.din(w_n613_0[2]));
	jspl3 jspl3_w_n613_4(.douta(w_n613_4[0]),.doutb(w_n613_4[1]),.doutc(w_n613_4[2]),.din(w_n613_1[0]));
	jspl3 jspl3_w_n613_5(.douta(w_n613_5[0]),.doutb(w_n613_5[1]),.doutc(w_n613_5[2]),.din(w_n613_1[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_dff_A_dEErKEAa2_1),.doutc(w_dff_A_5GC5YbDb3_2),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_dff_A_kvH05xRp7_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n619_1(.douta(w_n619_1[0]),.doutb(w_n619_1[1]),.doutc(w_n619_1[2]),.din(w_n619_0[0]));
	jspl3 jspl3_w_n620_0(.douta(w_n620_0[0]),.doutb(w_dff_A_QTSfA3wV0_1),.doutc(w_dff_A_ILyOpGBO9_2),.din(n620));
	jspl jspl_w_n620_1(.douta(w_n620_1[0]),.doutb(w_dff_A_FaTiuKzn8_1),.din(w_n620_0[0]));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_dff_A_FW533wll0_1),.din(n621));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_dff_A_Q8QOtOSR2_0),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(w_dff_B_1QNdUh026_3));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_dff_A_tG7bxNfY2_1),.din(n625));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl jspl_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n628_0(.douta(w_dff_A_00MTdIt77_0),.doutb(w_n628_0[1]),.doutc(w_dff_A_z1gmnbMd3_2),.din(n628));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_dff_A_SXc5389j0_1),.din(n632));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_dff_A_hNwrlskJ5_1),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_n635_1[0]),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.doutc(w_n637_0[2]),.din(n637));
	jspl jspl_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.din(n638));
	jspl3 jspl3_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.doutc(w_n639_0[2]),.din(n639));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_n641_0[2]),.din(n641));
	jspl3 jspl3_w_n641_1(.douta(w_n641_1[0]),.doutb(w_n641_1[1]),.doutc(w_n641_1[2]),.din(w_n641_0[0]));
	jspl3 jspl3_w_n644_0(.douta(w_dff_A_QzxyHL7W6_0),.doutb(w_n644_0[1]),.doutc(w_dff_A_SokhPaHg7_2),.din(n644));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_dff_A_0voaKU4p9_1),.doutc(w_dff_A_mQMoIth09_2),.din(n648));
	jspl jspl_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.din(w_n648_0[0]));
	jspl jspl_w_n649_0(.douta(w_dff_A_UkKsjaYi3_0),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n653_0(.douta(w_dff_A_CC5zD9ys5_0),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n654_0(.douta(w_dff_A_JWWby9fX1_0),.doutb(w_n654_0[1]),.doutc(w_n654_0[2]),.din(w_dff_B_Xxy0llxD2_3));
	jspl3 jspl3_w_n654_1(.douta(w_n654_1[0]),.doutb(w_dff_A_BTCzLtU25_1),.doutc(w_n654_1[2]),.din(w_n654_0[0]));
	jspl3 jspl3_w_n654_2(.douta(w_dff_A_r31cBjW88_0),.doutb(w_n654_2[1]),.doutc(w_n654_2[2]),.din(w_n654_0[1]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(n658));
	jspl jspl_w_n658_1(.douta(w_n658_1[0]),.doutb(w_n658_1[1]),.din(w_n658_0[0]));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_dff_A_vhzWELfx7_2),.din(n660));
	jspl jspl_w_n660_1(.douta(w_dff_A_FlMFMgdf0_0),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(w_dff_B_dIhJzJxG9_2));
	jspl jspl_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.din(n670));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl3 jspl3_w_n682_0(.douta(w_n682_0[0]),.doutb(w_dff_A_hoaHWpBQ4_1),.doutc(w_dff_A_JSKQu7Ck0_2),.din(n682));
	jspl jspl_w_n684_0(.douta(w_dff_A_PL9bxoyz9_0),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_dff_A_T52GB4Ep1_0),.doutb(w_n685_0[1]),.din(w_dff_B_CoCtGuNQ8_2));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_dff_A_DfkzCR1E7_1),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_dff_A_khTp7iO64_1),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_dff_A_F8hozB7X3_0),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_dff_A_lQRMyj9D2_0),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.doutc(w_n694_0[2]),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_n695_0[0]),.doutb(w_dff_A_92TCUL8i1_1),.doutc(w_n695_0[2]),.din(n695));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_dff_A_m3dvtZfp2_1),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n701_0(.douta(w_dff_A_L2wK5FBO0_0),.doutb(w_n701_0[1]),.din(n701));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_TrHiYAnk6_1),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_dff_A_k86KeRhH0_1),.din(n709));
	jspl jspl_w_n710_0(.douta(w_dff_A_DaFQTWao4_0),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_dff_A_tVHTqF3h4_0),.doutb(w_n711_0[1]),.din(w_dff_B_rEpscLp15_2));
	jspl3 jspl3_w_n713_0(.douta(w_dff_A_z9nyDZ5I5_0),.doutb(w_dff_A_77v8mn7W1_1),.doutc(w_n713_0[2]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(n715));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_MadxbEbI1_2));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_dff_A_iYbMZzK97_1),.din(n719));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_dff_A_Udpa4Dlm8_1),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_N68OXoit7_1),.din(n721));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_dff_A_x5eB3vcn8_1),.din(n722));
	jspl3 jspl3_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.doutc(w_n725_0[2]),.din(n725));
	jspl jspl_w_n726_0(.douta(w_dff_A_K3Qbqy7G6_0),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n728_0(.douta(w_dff_A_AuRtYqI56_0),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.doutc(w_n733_0[2]),.din(n733));
	jspl3 jspl3_w_n735_0(.douta(w_dff_A_sgODAPR95_0),.doutb(w_n735_0[1]),.doutc(w_n735_0[2]),.din(n735));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_dff_A_UwMNUtlo7_1),.doutc(w_dff_A_k3vSyhWN3_2),.din(n737));
	jspl jspl_w_n737_1(.douta(w_dff_A_pFcrzKxj4_0),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(w_dff_B_RuIzu3Mf8_2));
	jspl3 jspl3_w_n742_0(.douta(w_n742_0[0]),.doutb(w_dff_A_ttlHbz9T1_1),.doutc(w_n742_0[2]),.din(n742));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_dff_A_bow1sMlW8_1),.doutc(w_n746_0[2]),.din(n746));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl3 jspl3_w_n749_0(.douta(w_n749_0[0]),.doutb(w_dff_A_ldal8IrY6_1),.doutc(w_dff_A_D9J3qCLC2_2),.din(n749));
	jspl3 jspl3_w_n749_1(.douta(w_n749_1[0]),.doutb(w_dff_A_8MyeU4p57_1),.doutc(w_dff_A_knUKgd3s9_2),.din(w_n749_0[0]));
	jspl3 jspl3_w_n749_2(.douta(w_dff_A_kmiPpjBM6_0),.doutb(w_dff_A_GaxJsdja4_1),.doutc(w_n749_2[2]),.din(w_n749_0[1]));
	jspl3 jspl3_w_n749_3(.douta(w_n749_3[0]),.doutb(w_n749_3[1]),.doutc(w_n749_3[2]),.din(w_n749_0[2]));
	jspl3 jspl3_w_n749_4(.douta(w_n749_4[0]),.doutb(w_dff_A_dw7vFQVK4_1),.doutc(w_dff_A_jKQg6Bzu4_2),.din(w_n749_1[0]));
	jspl3 jspl3_w_n749_5(.douta(w_dff_A_2JdLEy3j5_0),.doutb(w_dff_A_WV7wOBFw4_1),.doutc(w_n749_5[2]),.din(w_n749_1[1]));
	jspl3 jspl3_w_n749_6(.douta(w_dff_A_XkHPpHga1_0),.doutb(w_n749_6[1]),.doutc(w_n749_6[2]),.din(w_n749_1[2]));
	jspl3 jspl3_w_n749_7(.douta(w_dff_A_9g7kbvuQ0_0),.doutb(w_n749_7[1]),.doutc(w_n749_7[2]),.din(w_n749_2[0]));
	jspl3 jspl3_w_n749_8(.douta(w_n749_8[0]),.doutb(w_dff_A_va9v80OY8_1),.doutc(w_dff_A_vPH2o0Fx6_2),.din(w_n749_2[1]));
	jspl3 jspl3_w_n749_9(.douta(w_dff_A_epYM8dkX3_0),.doutb(w_n749_9[1]),.doutc(w_dff_A_LPew5BSL7_2),.din(w_n749_2[2]));
	jspl3 jspl3_w_n749_10(.douta(w_n749_10[0]),.doutb(w_n749_10[1]),.doutc(w_n749_10[2]),.din(w_n749_3[0]));
	jspl3 jspl3_w_n749_11(.douta(w_n749_11[0]),.doutb(w_n749_11[1]),.doutc(w_n749_11[2]),.din(w_n749_3[1]));
	jspl3 jspl3_w_n749_12(.douta(w_n749_12[0]),.doutb(w_n749_12[1]),.doutc(w_n749_12[2]),.din(w_n749_3[2]));
	jspl jspl_w_n749_13(.douta(w_dff_A_CyS8Dk7A7_0),.doutb(w_n749_13[1]),.din(w_n749_4[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.doutc(w_n750_0[2]),.din(n750));
	jspl3 jspl3_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.doutc(w_n750_1[2]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n750_2(.douta(w_n750_2[0]),.doutb(w_n750_2[1]),.doutc(w_n750_2[2]),.din(w_n750_0[1]));
	jspl3 jspl3_w_n750_3(.douta(w_n750_3[0]),.doutb(w_n750_3[1]),.doutc(w_n750_3[2]),.din(w_n750_0[2]));
	jspl3 jspl3_w_n750_4(.douta(w_n750_4[0]),.doutb(w_n750_4[1]),.doutc(w_n750_4[2]),.din(w_n750_1[0]));
	jspl3 jspl3_w_n750_5(.douta(w_n750_5[0]),.doutb(w_n750_5[1]),.doutc(w_n750_5[2]),.din(w_n750_1[1]));
	jspl3 jspl3_w_n750_6(.douta(w_n750_6[0]),.doutb(w_n750_6[1]),.doutc(w_n750_6[2]),.din(w_n750_1[2]));
	jspl3 jspl3_w_n750_7(.douta(w_n750_7[0]),.doutb(w_n750_7[1]),.doutc(w_n750_7[2]),.din(w_n750_2[0]));
	jspl3 jspl3_w_n750_8(.douta(w_n750_8[0]),.doutb(w_n750_8[1]),.doutc(w_n750_8[2]),.din(w_n750_2[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_dff_A_aQ50xBuz5_1),.doutc(w_dff_A_4WBJbeab2_2),.din(w_dff_B_t1FXFAaZ7_3));
	jspl jspl_w_n753_1(.douta(w_dff_A_hurffN830_0),.doutb(w_n753_1[1]),.din(w_n753_0[0]));
	jspl jspl_w_n755_0(.douta(w_dff_A_SiWftj9M9_0),.doutb(w_n755_0[1]),.din(n755));
	jspl3 jspl3_w_n763_0(.douta(w_dff_A_PwUBuEfH9_0),.doutb(w_n763_0[1]),.doutc(w_n763_0[2]),.din(n763));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl jspl_w_n779_0(.douta(w_dff_A_rkyTETuQ0_0),.doutb(w_n779_0[1]),.din(n779));
	jspl3 jspl3_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.doutc(w_n786_0[2]),.din(n786));
	jspl3 jspl3_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.doutc(w_n788_0[2]),.din(n788));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_dff_A_xjVBSbwO5_1),.doutc(w_dff_A_GNJrBlpy1_2),.din(n790));
	jspl3 jspl3_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.doutc(w_dff_A_O57uuZ4N1_2),.din(n792));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.doutc(w_n797_1[2]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_n797_2[2]),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_dff_A_rkrxYc2d2_0),.doutb(w_n797_3[1]),.doutc(w_n797_3[2]),.din(w_n797_0[2]));
	jspl3 jspl3_w_n797_4(.douta(w_dff_A_drLVlnn43_0),.doutb(w_n797_4[1]),.doutc(w_dff_A_Jk8JySbY0_2),.din(w_n797_1[0]));
	jspl3 jspl3_w_n797_5(.douta(w_n797_5[0]),.doutb(w_dff_A_83cHrO3Z0_1),.doutc(w_n797_5[2]),.din(w_n797_1[1]));
	jspl3 jspl3_w_n797_6(.douta(w_dff_A_i7vIy5nd8_0),.doutb(w_n797_6[1]),.doutc(w_dff_A_w1EBiFrA3_2),.din(w_n797_1[2]));
	jspl3 jspl3_w_n797_7(.douta(w_n797_7[0]),.doutb(w_dff_A_8yAFZfdD0_1),.doutc(w_n797_7[2]),.din(w_n797_2[0]));
	jspl3 jspl3_w_n797_8(.douta(w_dff_A_7CmtykPV7_0),.doutb(w_n797_8[1]),.doutc(w_dff_A_VNLjHoOq3_2),.din(w_n797_2[1]));
	jspl jspl_w_n797_9(.douta(w_n797_9[0]),.doutb(w_dff_A_J7RHUXOW9_1),.din(w_n797_2[2]));
	jspl3 jspl3_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.doutc(w_n798_0[2]),.din(n798));
	jspl jspl_w_n798_1(.douta(w_n798_1[0]),.doutb(w_n798_1[1]),.din(w_n798_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_dff_A_3NmwBAyE8_1),.doutc(w_dff_A_hOX6vQYZ3_2),.din(w_dff_B_w6LEIGgm5_3));
	jspl3 jspl3_w_n800_1(.douta(w_n800_1[0]),.doutb(w_dff_A_Ox8FuV760_1),.doutc(w_dff_A_DSftXgBI3_2),.din(w_n800_0[0]));
	jspl3 jspl3_w_n800_2(.douta(w_n800_2[0]),.doutb(w_dff_A_VSsgog7F1_1),.doutc(w_dff_A_PnFovOBO9_2),.din(w_n800_0[1]));
	jspl3 jspl3_w_n800_3(.douta(w_n800_3[0]),.doutb(w_dff_A_CzjPq7vf6_1),.doutc(w_dff_A_Lb63Q02A7_2),.din(w_n800_0[2]));
	jspl jspl_w_n800_4(.douta(w_dff_A_FoZjywm18_0),.doutb(w_n800_4[1]),.din(w_n800_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_dff_A_IPnPPsxj1_0),.doutb(w_dff_A_4L6nhCvO8_1),.doutc(w_n814_0[2]),.din(n814));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_dff_A_xhbIWgCU4_1),.doutc(w_n819_0[2]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_dff_A_ZdDOikhV5_1),.din(n821));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n836_0(.douta(w_dff_A_5bRvF0Nh4_0),.doutb(w_n836_0[1]),.din(n836));
	jspl jspl_w_n847_0(.douta(w_dff_A_ww4RAWBC9_0),.doutb(w_n847_0[1]),.din(n847));
	jspl3 jspl3_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.doutc(w_n852_0[2]),.din(n852));
	jspl3 jspl3_w_n852_1(.douta(w_n852_1[0]),.doutb(w_n852_1[1]),.doutc(w_n852_1[2]),.din(w_n852_0[0]));
	jspl3 jspl3_w_n852_2(.douta(w_n852_2[0]),.doutb(w_n852_2[1]),.doutc(w_n852_2[2]),.din(w_n852_0[1]));
	jspl3 jspl3_w_n852_3(.douta(w_dff_A_aOhPuqhi6_0),.doutb(w_n852_3[1]),.doutc(w_n852_3[2]),.din(w_n852_0[2]));
	jspl3 jspl3_w_n852_4(.douta(w_dff_A_cCkSWa6R3_0),.doutb(w_n852_4[1]),.doutc(w_dff_A_0BqAqfk73_2),.din(w_n852_1[0]));
	jspl3 jspl3_w_n852_5(.douta(w_n852_5[0]),.doutb(w_dff_A_0wRL0BA83_1),.doutc(w_dff_A_2rHcka5g9_2),.din(w_n852_1[1]));
	jspl3 jspl3_w_n852_6(.douta(w_n852_6[0]),.doutb(w_n852_6[1]),.doutc(w_dff_A_9x3Yo8EN9_2),.din(w_n852_1[2]));
	jspl3 jspl3_w_n852_7(.douta(w_dff_A_AyIjvPMV7_0),.doutb(w_n852_7[1]),.doutc(w_dff_A_D7jBCDW84_2),.din(w_n852_2[0]));
	jspl3 jspl3_w_n852_8(.douta(w_n852_8[0]),.doutb(w_dff_A_e0eMipcg4_1),.doutc(w_n852_8[2]),.din(w_n852_2[1]));
	jspl jspl_w_n852_9(.douta(w_n852_9[0]),.doutb(w_dff_A_qM0F7uvM9_1),.din(w_n852_2[2]));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_dff_A_HyE5cwxc9_1),.doutc(w_dff_A_VhhiEz3N5_2),.din(w_dff_B_ywEgtm6v0_3));
	jspl3 jspl3_w_n854_1(.douta(w_n854_1[0]),.doutb(w_dff_A_TUOlpUU97_1),.doutc(w_dff_A_AU70l0BR0_2),.din(w_n854_0[0]));
	jspl3 jspl3_w_n854_2(.douta(w_dff_A_uPx2Fj0u1_0),.doutb(w_dff_A_Yb84MPbL5_1),.doutc(w_n854_2[2]),.din(w_n854_0[1]));
	jspl3 jspl3_w_n854_3(.douta(w_n854_3[0]),.doutb(w_dff_A_7V3vbrfp1_1),.doutc(w_dff_A_wQvkC4ud0_2),.din(w_n854_0[2]));
	jspl jspl_w_n854_4(.douta(w_dff_A_7k4NVCHH8_0),.doutb(w_n854_4[1]),.din(w_n854_1[0]));
	jspl3 jspl3_w_n865_0(.douta(w_dff_A_xh1MlD5z4_0),.doutb(w_n865_0[1]),.doutc(w_dff_A_VMAvBlKx6_2),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.din(n868));
	jspl jspl_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl jspl_w_n880_0(.douta(w_dff_A_9GCQO9zD4_0),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(n890));
	jspl jspl_w_n901_0(.douta(w_dff_A_F6Ryisq53_0),.doutb(w_n901_0[1]),.din(n901));
	jspl3 jspl3_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.doutc(w_dff_A_RqEWupQx7_2),.din(n923));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.doutc(w_dff_A_vmsZkfZI1_2),.din(n938));
	jspl3 jspl3_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.doutc(w_n940_0[2]),.din(n940));
	jspl jspl_w_n940_1(.douta(w_n940_1[0]),.doutb(w_n940_1[1]),.din(w_n940_0[0]));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_dff_A_prQ93bQ73_1),.din(n949));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl3 jspl3_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.doutc(w_dff_A_bluO7SOM9_2),.din(n954));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_dff_A_MOvyumZz3_1),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_dff_A_VvpmMaxw4_1),.din(n989));
	jspl3 jspl3_w_n993_0(.douta(w_n993_0[0]),.doutb(w_dff_A_IAF5Qtnl9_1),.doutc(w_dff_A_8376GmCA9_2),.din(n993));
	jspl3 jspl3_w_n993_1(.douta(w_n993_1[0]),.doutb(w_dff_A_sIofJAnO1_1),.doutc(w_dff_A_iJo7wsB24_2),.din(w_n993_0[0]));
	jspl3 jspl3_w_n993_2(.douta(w_dff_A_eu48OquP3_0),.doutb(w_n993_2[1]),.doutc(w_dff_A_t4Fis4ED6_2),.din(w_n993_0[1]));
	jspl3 jspl3_w_n993_3(.douta(w_dff_A_5zgclu6e2_0),.doutb(w_dff_A_WrwQKUNH7_1),.doutc(w_n993_3[2]),.din(w_n993_0[2]));
	jspl3 jspl3_w_n993_4(.douta(w_dff_A_YwEznwgY8_0),.doutb(w_dff_A_hmqJmvhe9_1),.doutc(w_n993_4[2]),.din(w_n993_1[0]));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n994_1(.douta(w_n994_1[0]),.doutb(w_n994_1[1]),.doutc(w_n994_1[2]),.din(w_n994_0[0]));
	jspl3 jspl3_w_n994_2(.douta(w_n994_2[0]),.doutb(w_n994_2[1]),.doutc(w_n994_2[2]),.din(w_n994_0[1]));
	jspl3 jspl3_w_n994_3(.douta(w_n994_3[0]),.doutb(w_n994_3[1]),.doutc(w_n994_3[2]),.din(w_n994_0[2]));
	jspl jspl_w_n994_4(.douta(w_n994_4[0]),.doutb(w_n994_4[1]),.din(w_n994_1[0]));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl3 jspl3_w_n996_1(.douta(w_n996_1[0]),.doutb(w_n996_1[1]),.doutc(w_n996_1[2]),.din(w_n996_0[0]));
	jspl3 jspl3_w_n996_2(.douta(w_n996_2[0]),.doutb(w_n996_2[1]),.doutc(w_n996_2[2]),.din(w_n996_0[1]));
	jspl3 jspl3_w_n996_3(.douta(w_n996_3[0]),.doutb(w_n996_3[1]),.doutc(w_n996_3[2]),.din(w_n996_0[2]));
	jspl jspl_w_n996_4(.douta(w_n996_4[0]),.doutb(w_n996_4[1]),.din(w_n996_1[0]));
	jspl3 jspl3_w_n999_0(.douta(w_dff_A_nJlTbF2Y5_0),.doutb(w_dff_A_jDTP8mhR3_1),.doutc(w_n999_0[2]),.din(w_dff_B_YUHuGYOJ2_3));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_YtguDoaI5_0),.doutb(w_dff_A_OSrG8lVv8_1),.doutc(w_n999_1[2]),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_w5yFxTCv2_0),.doutb(w_dff_A_Nfz1J6KG2_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_nw6sdVGv8_0),.doutb(w_dff_A_V9tpnX0W9_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl3 jspl3_w_n1007_0(.douta(w_dff_A_7Vx558mB1_0),.doutb(w_dff_A_KdQ8m5yz3_1),.doutc(w_n1007_0[2]),.din(w_dff_B_sxP123rE8_3));
	jspl3 jspl3_w_n1007_1(.douta(w_n1007_1[0]),.doutb(w_dff_A_rWnb6qNO3_1),.doutc(w_dff_A_LNXDQdP04_2),.din(w_n1007_0[0]));
	jspl3 jspl3_w_n1007_2(.douta(w_dff_A_94cTNurI0_0),.doutb(w_dff_A_mcsujQa73_1),.doutc(w_n1007_2[2]),.din(w_n1007_0[1]));
	jspl3 jspl3_w_n1007_3(.douta(w_n1007_3[0]),.doutb(w_dff_A_ARkK3bjp4_1),.doutc(w_n1007_3[2]),.din(w_n1007_0[2]));
	jspl3 jspl3_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_dff_A_BDIoTfWJ6_1),.doutc(w_dff_A_ctauFzo35_2),.din(n1008));
	jspl3 jspl3_w_n1008_1(.douta(w_n1008_1[0]),.doutb(w_dff_A_HlNI22Kk6_1),.doutc(w_dff_A_smbwUTM68_2),.din(w_n1008_0[0]));
	jspl3 jspl3_w_n1008_2(.douta(w_dff_A_hmk7Jl116_0),.doutb(w_n1008_2[1]),.doutc(w_dff_A_Jdvyeqj88_2),.din(w_n1008_0[1]));
	jspl3 jspl3_w_n1008_3(.douta(w_dff_A_BaOSPFsm5_0),.doutb(w_dff_A_rDg5QNjv5_1),.doutc(w_n1008_3[2]),.din(w_n1008_0[2]));
	jspl3 jspl3_w_n1008_4(.douta(w_dff_A_9ZG8s6Sg5_0),.doutb(w_n1008_4[1]),.doutc(w_dff_A_LO8UWQR42_2),.din(w_n1008_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl3 jspl3_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.doutc(w_n1012_1[2]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1012_2(.douta(w_n1012_2[0]),.doutb(w_n1012_2[1]),.doutc(w_n1012_2[2]),.din(w_n1012_0[1]));
	jspl3 jspl3_w_n1012_3(.douta(w_n1012_3[0]),.doutb(w_n1012_3[1]),.doutc(w_n1012_3[2]),.din(w_n1012_0[2]));
	jspl jspl_w_n1012_4(.douta(w_n1012_4[0]),.doutb(w_n1012_4[1]),.din(w_n1012_1[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl3 jspl3_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.doutc(w_n1014_1[2]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1014_2(.douta(w_n1014_2[0]),.doutb(w_n1014_2[1]),.doutc(w_n1014_2[2]),.din(w_n1014_0[1]));
	jspl3 jspl3_w_n1014_3(.douta(w_n1014_3[0]),.doutb(w_n1014_3[1]),.doutc(w_n1014_3[2]),.din(w_n1014_0[2]));
	jspl jspl_w_n1014_4(.douta(w_n1014_4[0]),.doutb(w_n1014_4[1]),.din(w_n1014_1[0]));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1019_1(.douta(w_n1019_1[0]),.doutb(w_n1019_1[1]),.din(w_n1019_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl3 jspl3_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.doutc(w_n1043_0[2]),.din(n1043));
	jspl jspl_w_n1043_1(.douta(w_n1043_1[0]),.doutb(w_n1043_1[1]),.din(w_n1043_0[0]));
	jspl3 jspl3_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.doutc(w_n1052_0[2]),.din(n1052));
	jspl jspl_w_n1052_1(.douta(w_n1052_1[0]),.doutb(w_n1052_1[1]),.din(w_n1052_0[0]));
	jspl3 jspl3_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.doutc(w_n1054_0[2]),.din(n1054));
	jspl jspl_w_n1054_1(.douta(w_n1054_1[0]),.doutb(w_n1054_1[1]),.din(w_n1054_0[0]));
	jspl jspl_w_n1177_0(.douta(w_dff_A_i4bemp5d7_0),.doutb(w_n1177_0[1]),.din(w_dff_B_cMRgaMlm1_2));
	jspl jspl_w_n1179_0(.douta(w_dff_A_euOf8vAs0_0),.doutb(w_n1179_0[1]),.din(n1179));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl3 jspl3_w_n1196_1(.douta(w_n1196_1[0]),.doutb(w_n1196_1[1]),.doutc(w_n1196_1[2]),.din(w_n1196_0[0]));
	jspl3 jspl3_w_n1201_0(.douta(w_dff_A_Z9NEU7h14_0),.doutb(w_dff_A_1DbhtSJM9_1),.doutc(w_n1201_0[2]),.din(w_dff_B_sWMDizUz3_3));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.doutc(w_n1213_0[2]),.din(n1213));
	jspl3 jspl3_w_n1213_1(.douta(w_n1213_1[0]),.doutb(w_n1213_1[1]),.doutc(w_n1213_1[2]),.din(w_n1213_0[0]));
	jspl3 jspl3_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.doutc(w_n1236_0[2]),.din(n1236));
	jspl3 jspl3_w_n1236_1(.douta(w_n1236_1[0]),.doutb(w_n1236_1[1]),.doutc(w_n1236_1[2]),.din(w_n1236_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl3 jspl3_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.doutc(w_n1251_1[2]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.doutc(w_n1279_0[2]),.din(n1279));
	jspl jspl_w_n1279_1(.douta(w_n1279_1[0]),.doutb(w_n1279_1[1]),.din(w_n1279_0[0]));
	jspl3 jspl3_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.doutc(w_n1297_0[2]),.din(n1297));
	jspl jspl_w_n1297_1(.douta(w_n1297_1[0]),.doutb(w_n1297_1[1]),.din(w_n1297_0[0]));
	jspl3 jspl3_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.doutc(w_n1299_0[2]),.din(n1299));
	jspl jspl_w_n1299_1(.douta(w_n1299_1[0]),.doutb(w_n1299_1[1]),.din(w_n1299_0[0]));
	jspl3 jspl3_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.doutc(w_n1410_0[2]),.din(n1410));
	jspl3 jspl3_w_n1412_0(.douta(w_n1412_0[0]),.doutb(w_dff_A_jvyrUwuN8_1),.doutc(w_dff_A_EE610UcN3_2),.din(w_dff_B_33bhuAvl8_3));
	jspl jspl_w_n1416_0(.douta(w_n1416_0[0]),.doutb(w_dff_A_pYkteeSe7_1),.din(w_dff_B_bSGZwCqE4_2));
	jspl jspl_w_n1422_0(.douta(w_n1422_0[0]),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1428_0(.douta(w_dff_A_5dDgk8ii0_0),.doutb(w_n1428_0[1]),.din(w_dff_B_uNP6423W8_2));
	jspl jspl_w_n1429_0(.douta(w_dff_A_WwVYqvUf4_0),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1451_0(.douta(w_dff_A_8IqcREHf8_0),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1503_0(.douta(w_n1503_0[0]),.doutb(w_n1503_0[1]),.din(n1503));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1592_0(.douta(w_n1592_0[0]),.doutb(w_n1592_0[1]),.din(n1592));
	jspl jspl_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.din(n1593));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1599_0(.douta(w_dff_A_TtdV9xNS0_0),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_dff_A_AyQKETKV8_1),.din(n1603));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1609_0(.douta(w_dff_A_usuy5aFg9_0),.doutb(w_n1609_0[1]),.din(w_dff_B_HQmzkpsW9_2));
	jspl3 jspl3_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.doutc(w_n1611_0[2]),.din(n1611));
	jspl jspl_w_n1613_0(.douta(w_n1613_0[0]),.doutb(w_n1613_0[1]),.din(n1613));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(n1615));
	jspl jspl_w_n1618_0(.douta(w_dff_A_JE3qdwRv2_0),.doutb(w_n1618_0[1]),.din(w_dff_B_2Wbpd6sD9_2));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_Ol8i2kYi7_2));
	jspl jspl_w_n1637_0(.douta(w_dff_A_a3aub9DV0_0),.doutb(w_n1637_0[1]),.din(w_dff_B_yPMzt06f5_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(n1643));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.din(n1652));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl3 jspl3_w_n1674_0(.douta(w_n1674_0[0]),.doutb(w_n1674_0[1]),.doutc(w_n1674_0[2]),.din(n1674));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_n1675_0[1]),.din(n1675));
	jspl3 jspl3_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.doutc(w_n1679_0[2]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_CBr7vovW7_2));
	jspl jspl_w_n1695_0(.douta(w_n1695_0[0]),.doutb(w_n1695_0[1]),.din(w_dff_B_Jzd9k4Fx3_2));
	jspl jspl_w_n1698_0(.douta(w_n1698_0[0]),.doutb(w_n1698_0[1]),.din(w_dff_B_NlFn00mt7_2));
	jdff dff_B_1GtAzzyc1_1(.din(G136),.dout(w_dff_B_1GtAzzyc1_1),.clk(gclk));
	jdff dff_B_uqSiIOCB0_0(.din(G2824),.dout(w_dff_B_uqSiIOCB0_0),.clk(gclk));
	jdff dff_A_9AfsaUq23_0(.dout(w_G809_3[0]),.din(w_dff_A_9AfsaUq23_0),.clk(gclk));
	jdff dff_B_kF86fxm53_0(.din(n342),.dout(w_dff_B_kF86fxm53_0),.clk(gclk));
	jdff dff_A_s5V3QPdz0_2(.dout(w_G809_2[2]),.din(w_dff_A_s5V3QPdz0_2),.clk(gclk));
	jdff dff_B_vir5UhkS1_1(.din(G24),.dout(w_dff_B_vir5UhkS1_1),.clk(gclk));
	jdff dff_B_80zcCL4t4_0(.din(n347),.dout(w_dff_B_80zcCL4t4_0),.clk(gclk));
	jdff dff_B_iajVVK8S0_1(.din(G26),.dout(w_dff_B_iajVVK8S0_1),.clk(gclk));
	jdff dff_A_ycvSEpNX4_0(.dout(w_G141_2[0]),.din(w_dff_A_ycvSEpNX4_0),.clk(gclk));
	jdff dff_A_ntJFtxVS6_0(.dout(w_dff_A_ycvSEpNX4_0),.din(w_dff_A_ntJFtxVS6_0),.clk(gclk));
	jdff dff_A_zMFKEvft7_1(.dout(w_G141_2[1]),.din(w_dff_A_zMFKEvft7_1),.clk(gclk));
	jdff dff_A_V5xbFpuQ9_1(.dout(w_dff_A_zMFKEvft7_1),.din(w_dff_A_V5xbFpuQ9_1),.clk(gclk));
	jdff dff_B_WhznrxG92_0(.din(n352),.dout(w_dff_B_WhznrxG92_0),.clk(gclk));
	jdff dff_B_uKAsZBfU9_1(.din(G79),.dout(w_dff_B_uKAsZBfU9_1),.clk(gclk));
	jdff dff_B_6oA78GKR0_1(.din(n355),.dout(w_dff_B_6oA78GKR0_1),.clk(gclk));
	jdff dff_B_i1OZVmBg6_1(.din(G82),.dout(w_dff_B_i1OZVmBg6_1),.clk(gclk));
	jdff dff_A_wBPBDoQH6_0(.dout(w_G2358_2[0]),.din(w_dff_A_wBPBDoQH6_0),.clk(gclk));
	jdff dff_A_kkDkeOtI7_1(.dout(w_G2358_2[1]),.din(w_dff_A_kkDkeOtI7_1),.clk(gclk));
	jdff dff_A_uOTPqfW57_0(.dout(w_G809_1[0]),.din(w_dff_A_uOTPqfW57_0),.clk(gclk));
	jdff dff_A_tBwK81W68_1(.dout(w_G141_1[1]),.din(w_dff_A_tBwK81W68_1),.clk(gclk));
	jdff dff_A_URWs1D7U2_1(.dout(w_dff_A_tBwK81W68_1),.din(w_dff_A_URWs1D7U2_1),.clk(gclk));
	jdff dff_A_KKMLDXxK0_2(.dout(w_G141_1[2]),.din(w_dff_A_KKMLDXxK0_2),.clk(gclk));
	jdff dff_A_U92YXMBk7_2(.dout(w_dff_A_KKMLDXxK0_2),.din(w_dff_A_U92YXMBk7_2),.clk(gclk));
	jdff dff_B_4OnXHcKF9_1(.din(n399),.dout(w_dff_B_4OnXHcKF9_1),.clk(gclk));
	jdff dff_B_n6bJKEiU7_1(.din(n424),.dout(w_dff_B_n6bJKEiU7_1),.clk(gclk));
	jdff dff_B_dIhJzJxG9_2(.din(n661),.dout(w_dff_B_dIhJzJxG9_2),.clk(gclk));
	jdff dff_B_yoaHrVYM0_2(.din(n717),.dout(w_dff_B_yoaHrVYM0_2),.clk(gclk));
	jdff dff_B_MadxbEbI1_2(.din(w_dff_B_yoaHrVYM0_2),.dout(w_dff_B_MadxbEbI1_2),.clk(gclk));
	jdff dff_B_SXfYI3Is7_1(.din(n705),.dout(w_dff_B_SXfYI3Is7_1),.clk(gclk));
	jdff dff_B_RtgVay2W2_1(.din(w_dff_B_SXfYI3Is7_1),.dout(w_dff_B_RtgVay2W2_1),.clk(gclk));
	jdff dff_B_D8iqVJ2Q6_1(.din(w_dff_B_RtgVay2W2_1),.dout(w_dff_B_D8iqVJ2Q6_1),.clk(gclk));
	jdff dff_B_YAfW2rFd1_1(.din(w_dff_B_D8iqVJ2Q6_1),.dout(w_dff_B_YAfW2rFd1_1),.clk(gclk));
	jdff dff_B_F2MQMNNB6_1(.din(w_dff_B_YAfW2rFd1_1),.dout(w_dff_B_F2MQMNNB6_1),.clk(gclk));
	jdff dff_B_2I0qUByN0_1(.din(n706),.dout(w_dff_B_2I0qUByN0_1),.clk(gclk));
	jdff dff_B_xx9DLbcD3_1(.din(w_dff_B_2I0qUByN0_1),.dout(w_dff_B_xx9DLbcD3_1),.clk(gclk));
	jdff dff_B_9G05yIxf1_1(.din(w_dff_B_xx9DLbcD3_1),.dout(w_dff_B_9G05yIxf1_1),.clk(gclk));
	jdff dff_B_SxrYm4o84_1(.din(w_dff_B_9G05yIxf1_1),.dout(w_dff_B_SxrYm4o84_1),.clk(gclk));
	jdff dff_B_9kpzX39X0_1(.din(w_dff_B_SxrYm4o84_1),.dout(w_dff_B_9kpzX39X0_1),.clk(gclk));
	jdff dff_B_waXr1BrN4_3(.din(n611),.dout(w_dff_B_waXr1BrN4_3),.clk(gclk));
	jdff dff_B_xQTz6HIA3_3(.din(w_dff_B_waXr1BrN4_3),.dout(w_dff_B_xQTz6HIA3_3),.clk(gclk));
	jdff dff_B_wgFKBdCJ0_1(.din(n739),.dout(w_dff_B_wgFKBdCJ0_1),.clk(gclk));
	jdff dff_B_QS51zgDE7_1(.din(w_dff_B_wgFKBdCJ0_1),.dout(w_dff_B_QS51zgDE7_1),.clk(gclk));
	jdff dff_B_RuIzu3Mf8_2(.din(n738),.dout(w_dff_B_RuIzu3Mf8_2),.clk(gclk));
	jdff dff_A_FlMFMgdf0_0(.dout(w_n660_1[0]),.din(w_dff_A_FlMFMgdf0_0),.clk(gclk));
	jdff dff_B_6ySXAuP76_0(.din(n808),.dout(w_dff_B_6ySXAuP76_0),.clk(gclk));
	jdff dff_B_KXacjP3V7_0(.din(w_dff_B_6ySXAuP76_0),.dout(w_dff_B_KXacjP3V7_0),.clk(gclk));
	jdff dff_B_eJVw89vJ1_0(.din(w_dff_B_KXacjP3V7_0),.dout(w_dff_B_eJVw89vJ1_0),.clk(gclk));
	jdff dff_B_WuXnYcSF4_0(.din(w_dff_B_eJVw89vJ1_0),.dout(w_dff_B_WuXnYcSF4_0),.clk(gclk));
	jdff dff_B_J8ZGGgmS1_0(.din(w_dff_B_WuXnYcSF4_0),.dout(w_dff_B_J8ZGGgmS1_0),.clk(gclk));
	jdff dff_B_HCKpntyI3_0(.din(w_dff_B_J8ZGGgmS1_0),.dout(w_dff_B_HCKpntyI3_0),.clk(gclk));
	jdff dff_B_kc2nmk4k9_0(.din(w_dff_B_HCKpntyI3_0),.dout(w_dff_B_kc2nmk4k9_0),.clk(gclk));
	jdff dff_B_mUrQO9oR4_0(.din(w_dff_B_kc2nmk4k9_0),.dout(w_dff_B_mUrQO9oR4_0),.clk(gclk));
	jdff dff_B_UXsIwkmT9_0(.din(w_dff_B_mUrQO9oR4_0),.dout(w_dff_B_UXsIwkmT9_0),.clk(gclk));
	jdff dff_B_oP1k9NoK2_0(.din(n803),.dout(w_dff_B_oP1k9NoK2_0),.clk(gclk));
	jdff dff_B_lR45vIp78_0(.din(w_dff_B_oP1k9NoK2_0),.dout(w_dff_B_lR45vIp78_0),.clk(gclk));
	jdff dff_A_Yx7UmKv56_1(.dout(w_n797_9[1]),.din(w_dff_A_Yx7UmKv56_1),.clk(gclk));
	jdff dff_A_Crq9RCt17_1(.dout(w_dff_A_Yx7UmKv56_1),.din(w_dff_A_Crq9RCt17_1),.clk(gclk));
	jdff dff_A_9l0I1sTh6_1(.dout(w_dff_A_Crq9RCt17_1),.din(w_dff_A_9l0I1sTh6_1),.clk(gclk));
	jdff dff_A_8X4C068P3_1(.dout(w_dff_A_9l0I1sTh6_1),.din(w_dff_A_8X4C068P3_1),.clk(gclk));
	jdff dff_A_UvY8o15y2_1(.dout(w_dff_A_8X4C068P3_1),.din(w_dff_A_UvY8o15y2_1),.clk(gclk));
	jdff dff_A_jVnbCgHv4_1(.dout(w_dff_A_UvY8o15y2_1),.din(w_dff_A_jVnbCgHv4_1),.clk(gclk));
	jdff dff_A_McIVgIT22_1(.dout(w_dff_A_jVnbCgHv4_1),.din(w_dff_A_McIVgIT22_1),.clk(gclk));
	jdff dff_A_eIOOudUf5_1(.dout(w_dff_A_McIVgIT22_1),.din(w_dff_A_eIOOudUf5_1),.clk(gclk));
	jdff dff_A_J7RHUXOW9_1(.dout(w_dff_A_eIOOudUf5_1),.din(w_dff_A_J7RHUXOW9_1),.clk(gclk));
	jdff dff_B_1tmFAwfe5_0(.din(n861),.dout(w_dff_B_1tmFAwfe5_0),.clk(gclk));
	jdff dff_B_hjy2jNaQ9_0(.din(w_dff_B_1tmFAwfe5_0),.dout(w_dff_B_hjy2jNaQ9_0),.clk(gclk));
	jdff dff_B_YfZSxOQ37_0(.din(w_dff_B_hjy2jNaQ9_0),.dout(w_dff_B_YfZSxOQ37_0),.clk(gclk));
	jdff dff_B_YXU6TZLL5_0(.din(w_dff_B_YfZSxOQ37_0),.dout(w_dff_B_YXU6TZLL5_0),.clk(gclk));
	jdff dff_B_Hn7n8Wbo9_0(.din(w_dff_B_YXU6TZLL5_0),.dout(w_dff_B_Hn7n8Wbo9_0),.clk(gclk));
	jdff dff_B_RDjAUUkT5_0(.din(w_dff_B_Hn7n8Wbo9_0),.dout(w_dff_B_RDjAUUkT5_0),.clk(gclk));
	jdff dff_B_4CJRazDM9_0(.din(w_dff_B_RDjAUUkT5_0),.dout(w_dff_B_4CJRazDM9_0),.clk(gclk));
	jdff dff_B_Dj4j1axa2_0(.din(w_dff_B_4CJRazDM9_0),.dout(w_dff_B_Dj4j1axa2_0),.clk(gclk));
	jdff dff_B_aSz2eNAo4_0(.din(w_dff_B_Dj4j1axa2_0),.dout(w_dff_B_aSz2eNAo4_0),.clk(gclk));
	jdff dff_B_nUPCiQug9_2(.din(G61),.dout(w_dff_B_nUPCiQug9_2),.clk(gclk));
	jdff dff_B_WXh6wnPF1_0(.din(n856),.dout(w_dff_B_WXh6wnPF1_0),.clk(gclk));
	jdff dff_B_1lmb96HG0_0(.din(w_dff_B_WXh6wnPF1_0),.dout(w_dff_B_1lmb96HG0_0),.clk(gclk));
	jdff dff_A_IqOfsAYC0_1(.dout(w_n852_9[1]),.din(w_dff_A_IqOfsAYC0_1),.clk(gclk));
	jdff dff_A_v4pg8jNg8_1(.dout(w_dff_A_IqOfsAYC0_1),.din(w_dff_A_v4pg8jNg8_1),.clk(gclk));
	jdff dff_A_gRUaYSXs5_1(.dout(w_dff_A_v4pg8jNg8_1),.din(w_dff_A_gRUaYSXs5_1),.clk(gclk));
	jdff dff_A_tJBUgvJr6_1(.dout(w_dff_A_gRUaYSXs5_1),.din(w_dff_A_tJBUgvJr6_1),.clk(gclk));
	jdff dff_A_0cK7920E0_1(.dout(w_dff_A_tJBUgvJr6_1),.din(w_dff_A_0cK7920E0_1),.clk(gclk));
	jdff dff_A_Kxyba8K44_1(.dout(w_dff_A_0cK7920E0_1),.din(w_dff_A_Kxyba8K44_1),.clk(gclk));
	jdff dff_A_zDdPMkYz0_1(.dout(w_dff_A_Kxyba8K44_1),.din(w_dff_A_zDdPMkYz0_1),.clk(gclk));
	jdff dff_A_AGhSKuX16_1(.dout(w_dff_A_zDdPMkYz0_1),.din(w_dff_A_AGhSKuX16_1),.clk(gclk));
	jdff dff_A_qM0F7uvM9_1(.dout(w_dff_A_AGhSKuX16_1),.din(w_dff_A_qM0F7uvM9_1),.clk(gclk));
	jdff dff_B_D04IyGQz9_1(.din(n958),.dout(w_dff_B_D04IyGQz9_1),.clk(gclk));
	jdff dff_B_B3ZV9v6v5_1(.din(n961),.dout(w_dff_B_B3ZV9v6v5_1),.clk(gclk));
	jdff dff_B_Tdu0oli02_1(.din(w_dff_B_B3ZV9v6v5_1),.dout(w_dff_B_Tdu0oli02_1),.clk(gclk));
	jdff dff_B_jFyidKdb4_0(.din(n991),.dout(w_dff_B_jFyidKdb4_0),.clk(gclk));
	jdff dff_B_LAnULZFI4_1(.din(n975),.dout(w_dff_B_LAnULZFI4_1),.clk(gclk));
	jdff dff_B_1KWLkI3m7_1(.din(w_dff_B_LAnULZFI4_1),.dout(w_dff_B_1KWLkI3m7_1),.clk(gclk));
	jdff dff_B_TfsNJWrF9_1(.din(n971),.dout(w_dff_B_TfsNJWrF9_1),.clk(gclk));
	jdff dff_B_aWhiiJLm3_1(.din(n995),.dout(w_dff_B_aWhiiJLm3_1),.clk(gclk));
	jdff dff_B_zdnkO2lt6_1(.din(w_dff_B_aWhiiJLm3_1),.dout(w_dff_B_zdnkO2lt6_1),.clk(gclk));
	jdff dff_B_CnJApNPj8_1(.din(w_dff_B_zdnkO2lt6_1),.dout(w_dff_B_CnJApNPj8_1),.clk(gclk));
	jdff dff_B_XzphINxT3_1(.din(w_dff_B_CnJApNPj8_1),.dout(w_dff_B_XzphINxT3_1),.clk(gclk));
	jdff dff_B_8ekjMiix1_1(.din(w_dff_B_XzphINxT3_1),.dout(w_dff_B_8ekjMiix1_1),.clk(gclk));
	jdff dff_B_GHsEjHdk7_1(.din(w_dff_B_8ekjMiix1_1),.dout(w_dff_B_GHsEjHdk7_1),.clk(gclk));
	jdff dff_B_VZZxT2BA5_1(.din(w_dff_B_GHsEjHdk7_1),.dout(w_dff_B_VZZxT2BA5_1),.clk(gclk));
	jdff dff_B_Ykn1hPsE6_1(.din(w_dff_B_VZZxT2BA5_1),.dout(w_dff_B_Ykn1hPsE6_1),.clk(gclk));
	jdff dff_B_rNIQAiam6_1(.din(n997),.dout(w_dff_B_rNIQAiam6_1),.clk(gclk));
	jdff dff_B_qEiUIF176_1(.din(w_dff_B_rNIQAiam6_1),.dout(w_dff_B_qEiUIF176_1),.clk(gclk));
	jdff dff_B_BTRFv6GO1_1(.din(w_dff_B_qEiUIF176_1),.dout(w_dff_B_BTRFv6GO1_1),.clk(gclk));
	jdff dff_B_eHVGDM220_1(.din(w_dff_B_BTRFv6GO1_1),.dout(w_dff_B_eHVGDM220_1),.clk(gclk));
	jdff dff_B_MRVjuMTV2_1(.din(w_dff_B_eHVGDM220_1),.dout(w_dff_B_MRVjuMTV2_1),.clk(gclk));
	jdff dff_B_mQ31TKdw6_1(.din(w_dff_B_MRVjuMTV2_1),.dout(w_dff_B_mQ31TKdw6_1),.clk(gclk));
	jdff dff_B_VZpgtv9Y5_1(.din(w_dff_B_mQ31TKdw6_1),.dout(w_dff_B_VZpgtv9Y5_1),.clk(gclk));
	jdff dff_B_KpDqVaos2_1(.din(w_dff_B_VZpgtv9Y5_1),.dout(w_dff_B_KpDqVaos2_1),.clk(gclk));
	jdff dff_B_PTVEC55W7_1(.din(w_dff_B_KpDqVaos2_1),.dout(w_dff_B_PTVEC55W7_1),.clk(gclk));
	jdff dff_B_0I1c4ZuX8_0(.din(n1001),.dout(w_dff_B_0I1c4ZuX8_0),.clk(gclk));
	jdff dff_B_WqgVAaty1_0(.din(w_dff_B_0I1c4ZuX8_0),.dout(w_dff_B_WqgVAaty1_0),.clk(gclk));
	jdff dff_B_FCWVVXmB8_0(.din(n1016),.dout(w_dff_B_FCWVVXmB8_0),.clk(gclk));
	jdff dff_B_fEDGH8EZ6_0(.din(w_dff_B_FCWVVXmB8_0),.dout(w_dff_B_fEDGH8EZ6_0),.clk(gclk));
	jdff dff_B_yb2JosEl9_0(.din(w_dff_B_fEDGH8EZ6_0),.dout(w_dff_B_yb2JosEl9_0),.clk(gclk));
	jdff dff_B_It7SPVGc1_0(.din(w_dff_B_yb2JosEl9_0),.dout(w_dff_B_It7SPVGc1_0),.clk(gclk));
	jdff dff_B_EnJDi84e9_0(.din(w_dff_B_It7SPVGc1_0),.dout(w_dff_B_EnJDi84e9_0),.clk(gclk));
	jdff dff_B_d6okdsGf8_0(.din(w_dff_B_EnJDi84e9_0),.dout(w_dff_B_d6okdsGf8_0),.clk(gclk));
	jdff dff_B_u0iXXtuK6_0(.din(w_dff_B_d6okdsGf8_0),.dout(w_dff_B_u0iXXtuK6_0),.clk(gclk));
	jdff dff_B_lSXyQPV36_0(.din(w_dff_B_u0iXXtuK6_0),.dout(w_dff_B_lSXyQPV36_0),.clk(gclk));
	jdff dff_B_QqXudnfC0_0(.din(w_dff_B_lSXyQPV36_0),.dout(w_dff_B_QqXudnfC0_0),.clk(gclk));
	jdff dff_B_VQGxCGCs8_1(.din(n1013),.dout(w_dff_B_VQGxCGCs8_1),.clk(gclk));
	jdff dff_B_Lw4WQfms1_2(.din(G182),.dout(w_dff_B_Lw4WQfms1_2),.clk(gclk));
	jdff dff_B_esaDwXgw5_2(.din(w_dff_B_Lw4WQfms1_2),.dout(w_dff_B_esaDwXgw5_2),.clk(gclk));
	jdff dff_B_menrNAlj4_2(.din(G185),.dout(w_dff_B_menrNAlj4_2),.clk(gclk));
	jdff dff_B_Q7gad6Bs4_1(.din(n1006),.dout(w_dff_B_Q7gad6Bs4_1),.clk(gclk));
	jdff dff_B_1XnVT89E6_1(.din(w_dff_B_Q7gad6Bs4_1),.dout(w_dff_B_1XnVT89E6_1),.clk(gclk));
	jdff dff_B_q6VYX1OR3_1(.din(w_dff_B_1XnVT89E6_1),.dout(w_dff_B_q6VYX1OR3_1),.clk(gclk));
	jdff dff_B_ZB6kUhF76_1(.din(w_dff_B_q6VYX1OR3_1),.dout(w_dff_B_ZB6kUhF76_1),.clk(gclk));
	jdff dff_B_jPQLoBK69_1(.din(n777),.dout(w_dff_B_jPQLoBK69_1),.clk(gclk));
	jdff dff_B_ANVSRo600_1(.din(w_dff_B_jPQLoBK69_1),.dout(w_dff_B_ANVSRo600_1),.clk(gclk));
	jdff dff_B_5MbQrCJc8_1(.din(w_dff_B_ANVSRo600_1),.dout(w_dff_B_5MbQrCJc8_1),.clk(gclk));
	jdff dff_B_jgWblR193_1(.din(w_dff_B_5MbQrCJc8_1),.dout(w_dff_B_jgWblR193_1),.clk(gclk));
	jdff dff_B_2hXGawTK9_0(.din(n782),.dout(w_dff_B_2hXGawTK9_0),.clk(gclk));
	jdff dff_B_ZrCBIzZC1_0(.din(w_dff_B_2hXGawTK9_0),.dout(w_dff_B_ZrCBIzZC1_0),.clk(gclk));
	jdff dff_B_8HXx2yJO4_0(.din(w_dff_B_ZrCBIzZC1_0),.dout(w_dff_B_8HXx2yJO4_0),.clk(gclk));
	jdff dff_B_QMQVtFwl1_0(.din(w_dff_B_8HXx2yJO4_0),.dout(w_dff_B_QMQVtFwl1_0),.clk(gclk));
	jdff dff_B_CQjF9HTI5_1(.din(n536),.dout(w_dff_B_CQjF9HTI5_1),.clk(gclk));
	jdff dff_A_rkyTETuQ0_0(.dout(w_n779_0[0]),.din(w_dff_A_rkyTETuQ0_0),.clk(gclk));
	jdff dff_B_qq3VnTOQ7_1(.din(G117),.dout(w_dff_B_qq3VnTOQ7_1),.clk(gclk));
	jdff dff_B_tsE0BllG0_1(.din(w_dff_B_qq3VnTOQ7_1),.dout(w_dff_B_tsE0BllG0_1),.clk(gclk));
	jdff dff_B_ttqqGnET9_1(.din(n752),.dout(w_dff_B_ttqqGnET9_1),.clk(gclk));
	jdff dff_B_uoBLLF5g3_0(.din(n758),.dout(w_dff_B_uoBLLF5g3_0),.clk(gclk));
	jdff dff_A_3L5GuXNH8_0(.dout(w_n755_0[0]),.din(w_dff_A_3L5GuXNH8_0),.clk(gclk));
	jdff dff_A_XwW2Wqu36_0(.dout(w_dff_A_3L5GuXNH8_0),.din(w_dff_A_XwW2Wqu36_0),.clk(gclk));
	jdff dff_A_BQh33GQT4_0(.dout(w_dff_A_XwW2Wqu36_0),.din(w_dff_A_BQh33GQT4_0),.clk(gclk));
	jdff dff_A_Ju5TH4xT9_0(.dout(w_dff_A_BQh33GQT4_0),.din(w_dff_A_Ju5TH4xT9_0),.clk(gclk));
	jdff dff_A_m1c6lnTn3_0(.dout(w_dff_A_Ju5TH4xT9_0),.din(w_dff_A_m1c6lnTn3_0),.clk(gclk));
	jdff dff_A_m9RpRpGy0_0(.dout(w_dff_A_m1c6lnTn3_0),.din(w_dff_A_m9RpRpGy0_0),.clk(gclk));
	jdff dff_A_cTMAdxYM3_0(.dout(w_dff_A_m9RpRpGy0_0),.din(w_dff_A_cTMAdxYM3_0),.clk(gclk));
	jdff dff_A_SiWftj9M9_0(.dout(w_dff_A_cTMAdxYM3_0),.din(w_dff_A_SiWftj9M9_0),.clk(gclk));
	jdff dff_B_ZNVvaAH95_1(.din(G131),.dout(w_dff_B_ZNVvaAH95_1),.clk(gclk));
	jdff dff_B_RntSM2gG0_1(.din(w_dff_B_ZNVvaAH95_1),.dout(w_dff_B_RntSM2gG0_1),.clk(gclk));
	jdff dff_A_vkfbRAzT5_0(.dout(w_G137_9[0]),.din(w_dff_A_vkfbRAzT5_0),.clk(gclk));
	jdff dff_B_hVUzqmlY6_0(.din(n1028),.dout(w_dff_B_hVUzqmlY6_0),.clk(gclk));
	jdff dff_B_p9rBhHSU0_0(.din(w_dff_B_hVUzqmlY6_0),.dout(w_dff_B_p9rBhHSU0_0),.clk(gclk));
	jdff dff_B_FJ70SmwN3_0(.din(w_dff_B_p9rBhHSU0_0),.dout(w_dff_B_FJ70SmwN3_0),.clk(gclk));
	jdff dff_B_cbjbzLry7_0(.din(w_dff_B_FJ70SmwN3_0),.dout(w_dff_B_cbjbzLry7_0),.clk(gclk));
	jdff dff_B_VMPa116o2_0(.din(w_dff_B_cbjbzLry7_0),.dout(w_dff_B_VMPa116o2_0),.clk(gclk));
	jdff dff_B_M5gKOCH17_0(.din(w_dff_B_VMPa116o2_0),.dout(w_dff_B_M5gKOCH17_0),.clk(gclk));
	jdff dff_B_xQ7fOP5t3_0(.din(w_dff_B_M5gKOCH17_0),.dout(w_dff_B_xQ7fOP5t3_0),.clk(gclk));
	jdff dff_B_WfFlJPVz0_0(.din(w_dff_B_xQ7fOP5t3_0),.dout(w_dff_B_WfFlJPVz0_0),.clk(gclk));
	jdff dff_B_HbDo0Dos1_0(.din(w_dff_B_WfFlJPVz0_0),.dout(w_dff_B_HbDo0Dos1_0),.clk(gclk));
	jdff dff_B_J1xabP3Y8_0(.din(w_dff_B_HbDo0Dos1_0),.dout(w_dff_B_J1xabP3Y8_0),.clk(gclk));
	jdff dff_B_5Af90yN23_0(.din(w_dff_B_J1xabP3Y8_0),.dout(w_dff_B_5Af90yN23_0),.clk(gclk));
	jdff dff_B_vGfTQHdt9_0(.din(w_dff_B_5Af90yN23_0),.dout(w_dff_B_vGfTQHdt9_0),.clk(gclk));
	jdff dff_A_fczZGPYb8_0(.dout(w_n800_4[0]),.din(w_dff_A_fczZGPYb8_0),.clk(gclk));
	jdff dff_A_HexWks2A7_0(.dout(w_dff_A_fczZGPYb8_0),.din(w_dff_A_HexWks2A7_0),.clk(gclk));
	jdff dff_A_OPOV61q12_0(.dout(w_dff_A_HexWks2A7_0),.din(w_dff_A_OPOV61q12_0),.clk(gclk));
	jdff dff_A_fdTn3Grr8_0(.dout(w_dff_A_OPOV61q12_0),.din(w_dff_A_fdTn3Grr8_0),.clk(gclk));
	jdff dff_A_FoZjywm18_0(.dout(w_dff_A_fdTn3Grr8_0),.din(w_dff_A_FoZjywm18_0),.clk(gclk));
	jdff dff_B_in6b97hS3_0(.din(n1039),.dout(w_dff_B_in6b97hS3_0),.clk(gclk));
	jdff dff_B_P8pCc4jI2_0(.din(w_dff_B_in6b97hS3_0),.dout(w_dff_B_P8pCc4jI2_0),.clk(gclk));
	jdff dff_B_Y8jhCHRY6_0(.din(w_dff_B_P8pCc4jI2_0),.dout(w_dff_B_Y8jhCHRY6_0),.clk(gclk));
	jdff dff_B_DX72x1Dn3_0(.din(w_dff_B_Y8jhCHRY6_0),.dout(w_dff_B_DX72x1Dn3_0),.clk(gclk));
	jdff dff_B_SpDAdqbM9_0(.din(w_dff_B_DX72x1Dn3_0),.dout(w_dff_B_SpDAdqbM9_0),.clk(gclk));
	jdff dff_B_L8oDlve46_0(.din(w_dff_B_SpDAdqbM9_0),.dout(w_dff_B_L8oDlve46_0),.clk(gclk));
	jdff dff_B_8IYxjELw4_0(.din(w_dff_B_L8oDlve46_0),.dout(w_dff_B_8IYxjELw4_0),.clk(gclk));
	jdff dff_B_3xix8IXc8_0(.din(w_dff_B_8IYxjELw4_0),.dout(w_dff_B_3xix8IXc8_0),.clk(gclk));
	jdff dff_B_QABUrzbd0_0(.din(w_dff_B_3xix8IXc8_0),.dout(w_dff_B_QABUrzbd0_0),.clk(gclk));
	jdff dff_B_y2vmSPBM0_0(.din(w_dff_B_QABUrzbd0_0),.dout(w_dff_B_y2vmSPBM0_0),.clk(gclk));
	jdff dff_B_i0Opn9fq0_0(.din(w_dff_B_y2vmSPBM0_0),.dout(w_dff_B_i0Opn9fq0_0),.clk(gclk));
	jdff dff_B_zNb3Rqgq0_0(.din(w_dff_B_i0Opn9fq0_0),.dout(w_dff_B_zNb3Rqgq0_0),.clk(gclk));
	jdff dff_B_34QnpZ2M2_1(.din(n1031),.dout(w_dff_B_34QnpZ2M2_1),.clk(gclk));
	jdff dff_A_ztp9UyxC4_0(.dout(w_G4088_8[0]),.din(w_dff_A_ztp9UyxC4_0),.clk(gclk));
	jdff dff_A_h9GlRIyz6_0(.dout(w_dff_A_ztp9UyxC4_0),.din(w_dff_A_h9GlRIyz6_0),.clk(gclk));
	jdff dff_A_ZBcZCkIP4_0(.dout(w_dff_A_h9GlRIyz6_0),.din(w_dff_A_ZBcZCkIP4_0),.clk(gclk));
	jdff dff_A_jHY2LGTj7_0(.dout(w_dff_A_ZBcZCkIP4_0),.din(w_dff_A_jHY2LGTj7_0),.clk(gclk));
	jdff dff_A_lYA67wRe7_0(.dout(w_dff_A_jHY2LGTj7_0),.din(w_dff_A_lYA67wRe7_0),.clk(gclk));
	jdff dff_A_uTOJRq2Q8_0(.dout(w_dff_A_lYA67wRe7_0),.din(w_dff_A_uTOJRq2Q8_0),.clk(gclk));
	jdff dff_A_nLz6SNRi6_0(.dout(w_dff_A_uTOJRq2Q8_0),.din(w_dff_A_nLz6SNRi6_0),.clk(gclk));
	jdff dff_A_furoJDwM6_0(.dout(w_dff_A_nLz6SNRi6_0),.din(w_dff_A_furoJDwM6_0),.clk(gclk));
	jdff dff_A_OPFZvC1U0_0(.dout(w_dff_A_furoJDwM6_0),.din(w_dff_A_OPFZvC1U0_0),.clk(gclk));
	jdff dff_A_HOZ7xEdp7_0(.dout(w_dff_A_OPFZvC1U0_0),.din(w_dff_A_HOZ7xEdp7_0),.clk(gclk));
	jdff dff_A_P2qDmiei6_0(.dout(w_dff_A_HOZ7xEdp7_0),.din(w_dff_A_P2qDmiei6_0),.clk(gclk));
	jdff dff_A_ocmlcEj69_0(.dout(w_dff_A_P2qDmiei6_0),.din(w_dff_A_ocmlcEj69_0),.clk(gclk));
	jdff dff_A_CeCPHWaB6_2(.dout(w_G4088_8[2]),.din(w_dff_A_CeCPHWaB6_2),.clk(gclk));
	jdff dff_A_vyNwRoTY3_2(.dout(w_dff_A_CeCPHWaB6_2),.din(w_dff_A_vyNwRoTY3_2),.clk(gclk));
	jdff dff_A_jdFdgVQU4_2(.dout(w_dff_A_vyNwRoTY3_2),.din(w_dff_A_jdFdgVQU4_2),.clk(gclk));
	jdff dff_A_b2ctLjbA2_2(.dout(w_dff_A_jdFdgVQU4_2),.din(w_dff_A_b2ctLjbA2_2),.clk(gclk));
	jdff dff_A_ZeZAIU0i2_2(.dout(w_dff_A_b2ctLjbA2_2),.din(w_dff_A_ZeZAIU0i2_2),.clk(gclk));
	jdff dff_A_gJiX4mCC6_2(.dout(w_dff_A_ZeZAIU0i2_2),.din(w_dff_A_gJiX4mCC6_2),.clk(gclk));
	jdff dff_A_jVv2e0RD5_2(.dout(w_dff_A_gJiX4mCC6_2),.din(w_dff_A_jVv2e0RD5_2),.clk(gclk));
	jdff dff_A_3S53QUgj4_2(.dout(w_dff_A_jVv2e0RD5_2),.din(w_dff_A_3S53QUgj4_2),.clk(gclk));
	jdff dff_A_QnGWxoCM5_2(.dout(w_dff_A_3S53QUgj4_2),.din(w_dff_A_QnGWxoCM5_2),.clk(gclk));
	jdff dff_A_hWCudCpn0_2(.dout(w_dff_A_QnGWxoCM5_2),.din(w_dff_A_hWCudCpn0_2),.clk(gclk));
	jdff dff_A_6ocjygVS8_2(.dout(w_dff_A_hWCudCpn0_2),.din(w_dff_A_6ocjygVS8_2),.clk(gclk));
	jdff dff_A_LiETSce14_2(.dout(w_dff_A_6ocjygVS8_2),.din(w_dff_A_LiETSce14_2),.clk(gclk));
	jdff dff_A_66blaznK0_0(.dout(w_n797_8[0]),.din(w_dff_A_66blaznK0_0),.clk(gclk));
	jdff dff_A_4FlJvVeE8_0(.dout(w_dff_A_66blaznK0_0),.din(w_dff_A_4FlJvVeE8_0),.clk(gclk));
	jdff dff_A_O4QnsGew3_0(.dout(w_dff_A_4FlJvVeE8_0),.din(w_dff_A_O4QnsGew3_0),.clk(gclk));
	jdff dff_A_yaUNVupM8_0(.dout(w_dff_A_O4QnsGew3_0),.din(w_dff_A_yaUNVupM8_0),.clk(gclk));
	jdff dff_A_Qbry0MNV0_0(.dout(w_dff_A_yaUNVupM8_0),.din(w_dff_A_Qbry0MNV0_0),.clk(gclk));
	jdff dff_A_TAeVVpbe5_0(.dout(w_dff_A_Qbry0MNV0_0),.din(w_dff_A_TAeVVpbe5_0),.clk(gclk));
	jdff dff_A_Ffu6A3878_0(.dout(w_dff_A_TAeVVpbe5_0),.din(w_dff_A_Ffu6A3878_0),.clk(gclk));
	jdff dff_A_fTZisUBx1_0(.dout(w_dff_A_Ffu6A3878_0),.din(w_dff_A_fTZisUBx1_0),.clk(gclk));
	jdff dff_A_A35UpjuI3_0(.dout(w_dff_A_fTZisUBx1_0),.din(w_dff_A_A35UpjuI3_0),.clk(gclk));
	jdff dff_A_X0uJt3xl3_0(.dout(w_dff_A_A35UpjuI3_0),.din(w_dff_A_X0uJt3xl3_0),.clk(gclk));
	jdff dff_A_7CmtykPV7_0(.dout(w_dff_A_X0uJt3xl3_0),.din(w_dff_A_7CmtykPV7_0),.clk(gclk));
	jdff dff_A_GZg8pH6M2_2(.dout(w_n797_8[2]),.din(w_dff_A_GZg8pH6M2_2),.clk(gclk));
	jdff dff_A_cFPji26A3_2(.dout(w_dff_A_GZg8pH6M2_2),.din(w_dff_A_cFPji26A3_2),.clk(gclk));
	jdff dff_A_PyqQVyQN7_2(.dout(w_dff_A_cFPji26A3_2),.din(w_dff_A_PyqQVyQN7_2),.clk(gclk));
	jdff dff_A_hl3ZBUnU1_2(.dout(w_dff_A_PyqQVyQN7_2),.din(w_dff_A_hl3ZBUnU1_2),.clk(gclk));
	jdff dff_A_xETbLDDh2_2(.dout(w_dff_A_hl3ZBUnU1_2),.din(w_dff_A_xETbLDDh2_2),.clk(gclk));
	jdff dff_A_xlG8cCWC5_2(.dout(w_dff_A_xETbLDDh2_2),.din(w_dff_A_xlG8cCWC5_2),.clk(gclk));
	jdff dff_A_wOpDK0AH4_2(.dout(w_dff_A_xlG8cCWC5_2),.din(w_dff_A_wOpDK0AH4_2),.clk(gclk));
	jdff dff_A_kzUGrd8N4_2(.dout(w_dff_A_wOpDK0AH4_2),.din(w_dff_A_kzUGrd8N4_2),.clk(gclk));
	jdff dff_A_3AHbYvb48_2(.dout(w_dff_A_kzUGrd8N4_2),.din(w_dff_A_3AHbYvb48_2),.clk(gclk));
	jdff dff_A_VhiWsFc44_2(.dout(w_dff_A_3AHbYvb48_2),.din(w_dff_A_VhiWsFc44_2),.clk(gclk));
	jdff dff_A_TsJubJMW8_2(.dout(w_dff_A_VhiWsFc44_2),.din(w_dff_A_TsJubJMW8_2),.clk(gclk));
	jdff dff_A_VNLjHoOq3_2(.dout(w_dff_A_TsJubJMW8_2),.din(w_dff_A_VNLjHoOq3_2),.clk(gclk));
	jdff dff_B_THCpPPMj9_0(.din(n1050),.dout(w_dff_B_THCpPPMj9_0),.clk(gclk));
	jdff dff_B_yuabpuIt1_0(.din(w_dff_B_THCpPPMj9_0),.dout(w_dff_B_yuabpuIt1_0),.clk(gclk));
	jdff dff_B_G1tRvPUO4_0(.din(w_dff_B_yuabpuIt1_0),.dout(w_dff_B_G1tRvPUO4_0),.clk(gclk));
	jdff dff_B_ToE7XJ3Z9_0(.din(w_dff_B_G1tRvPUO4_0),.dout(w_dff_B_ToE7XJ3Z9_0),.clk(gclk));
	jdff dff_B_7mWaczjN3_0(.din(w_dff_B_ToE7XJ3Z9_0),.dout(w_dff_B_7mWaczjN3_0),.clk(gclk));
	jdff dff_B_chDO7ZiU7_0(.din(w_dff_B_7mWaczjN3_0),.dout(w_dff_B_chDO7ZiU7_0),.clk(gclk));
	jdff dff_B_0JLmbahI5_0(.din(w_dff_B_chDO7ZiU7_0),.dout(w_dff_B_0JLmbahI5_0),.clk(gclk));
	jdff dff_B_sKXTQ5WP4_0(.din(w_dff_B_0JLmbahI5_0),.dout(w_dff_B_sKXTQ5WP4_0),.clk(gclk));
	jdff dff_B_1vxwo5Pz7_0(.din(w_dff_B_sKXTQ5WP4_0),.dout(w_dff_B_1vxwo5Pz7_0),.clk(gclk));
	jdff dff_B_PDKL7CSO4_0(.din(w_dff_B_1vxwo5Pz7_0),.dout(w_dff_B_PDKL7CSO4_0),.clk(gclk));
	jdff dff_B_Id00WzHI6_0(.din(w_dff_B_PDKL7CSO4_0),.dout(w_dff_B_Id00WzHI6_0),.clk(gclk));
	jdff dff_B_j3L33nz34_1(.din(n1042),.dout(w_dff_B_j3L33nz34_1),.clk(gclk));
	jdff dff_B_JuabviMb4_1(.din(w_dff_B_j3L33nz34_1),.dout(w_dff_B_JuabviMb4_1),.clk(gclk));
	jdff dff_B_l7ktTNTI3_1(.din(w_dff_B_JuabviMb4_1),.dout(w_dff_B_l7ktTNTI3_1),.clk(gclk));
	jdff dff_A_BfyTGzgp9_1(.dout(w_n797_7[1]),.din(w_dff_A_BfyTGzgp9_1),.clk(gclk));
	jdff dff_A_PjX0Nso77_1(.dout(w_dff_A_BfyTGzgp9_1),.din(w_dff_A_PjX0Nso77_1),.clk(gclk));
	jdff dff_A_gZxUrYBL8_1(.dout(w_dff_A_PjX0Nso77_1),.din(w_dff_A_gZxUrYBL8_1),.clk(gclk));
	jdff dff_A_0eh4I4zt9_1(.dout(w_dff_A_gZxUrYBL8_1),.din(w_dff_A_0eh4I4zt9_1),.clk(gclk));
	jdff dff_A_CBI4nD3J7_1(.dout(w_dff_A_0eh4I4zt9_1),.din(w_dff_A_CBI4nD3J7_1),.clk(gclk));
	jdff dff_A_aBuZFZTV1_1(.dout(w_dff_A_CBI4nD3J7_1),.din(w_dff_A_aBuZFZTV1_1),.clk(gclk));
	jdff dff_A_VdyuK2dy6_1(.dout(w_dff_A_aBuZFZTV1_1),.din(w_dff_A_VdyuK2dy6_1),.clk(gclk));
	jdff dff_A_Jns33q6O2_1(.dout(w_dff_A_VdyuK2dy6_1),.din(w_dff_A_Jns33q6O2_1),.clk(gclk));
	jdff dff_A_mhuAIWXF2_1(.dout(w_dff_A_Jns33q6O2_1),.din(w_dff_A_mhuAIWXF2_1),.clk(gclk));
	jdff dff_A_8yAFZfdD0_1(.dout(w_dff_A_mhuAIWXF2_1),.din(w_dff_A_8yAFZfdD0_1),.clk(gclk));
	jdff dff_A_tK8GKuzK9_1(.dout(w_G4088_7[1]),.din(w_dff_A_tK8GKuzK9_1),.clk(gclk));
	jdff dff_A_wOOebpOE6_1(.dout(w_dff_A_tK8GKuzK9_1),.din(w_dff_A_wOOebpOE6_1),.clk(gclk));
	jdff dff_A_LEvTjwJc2_1(.dout(w_dff_A_wOOebpOE6_1),.din(w_dff_A_LEvTjwJc2_1),.clk(gclk));
	jdff dff_A_XHwHNi6B0_1(.dout(w_dff_A_LEvTjwJc2_1),.din(w_dff_A_XHwHNi6B0_1),.clk(gclk));
	jdff dff_A_b8chBR272_1(.dout(w_dff_A_XHwHNi6B0_1),.din(w_dff_A_b8chBR272_1),.clk(gclk));
	jdff dff_A_ZnkAIT4d6_1(.dout(w_dff_A_b8chBR272_1),.din(w_dff_A_ZnkAIT4d6_1),.clk(gclk));
	jdff dff_A_HLLOjFs03_1(.dout(w_dff_A_ZnkAIT4d6_1),.din(w_dff_A_HLLOjFs03_1),.clk(gclk));
	jdff dff_A_wSRdn8vo9_1(.dout(w_dff_A_HLLOjFs03_1),.din(w_dff_A_wSRdn8vo9_1),.clk(gclk));
	jdff dff_A_LFa27Mez9_1(.dout(w_dff_A_wSRdn8vo9_1),.din(w_dff_A_LFa27Mez9_1),.clk(gclk));
	jdff dff_B_AKAmyV3f7_0(.din(n1061),.dout(w_dff_B_AKAmyV3f7_0),.clk(gclk));
	jdff dff_B_0uXH1LMm7_0(.din(w_dff_B_AKAmyV3f7_0),.dout(w_dff_B_0uXH1LMm7_0),.clk(gclk));
	jdff dff_B_iQ8kPDyP1_0(.din(w_dff_B_0uXH1LMm7_0),.dout(w_dff_B_iQ8kPDyP1_0),.clk(gclk));
	jdff dff_B_L4P7t1YE8_0(.din(w_dff_B_iQ8kPDyP1_0),.dout(w_dff_B_L4P7t1YE8_0),.clk(gclk));
	jdff dff_B_PbuM9bPv0_0(.din(w_dff_B_L4P7t1YE8_0),.dout(w_dff_B_PbuM9bPv0_0),.clk(gclk));
	jdff dff_B_sh9XEXea2_0(.din(w_dff_B_PbuM9bPv0_0),.dout(w_dff_B_sh9XEXea2_0),.clk(gclk));
	jdff dff_B_q45UdfyB3_0(.din(w_dff_B_sh9XEXea2_0),.dout(w_dff_B_q45UdfyB3_0),.clk(gclk));
	jdff dff_B_B6Fs37IB9_0(.din(w_dff_B_q45UdfyB3_0),.dout(w_dff_B_B6Fs37IB9_0),.clk(gclk));
	jdff dff_B_5lTzlez44_0(.din(w_dff_B_B6Fs37IB9_0),.dout(w_dff_B_5lTzlez44_0),.clk(gclk));
	jdff dff_B_2fehSlEE1_0(.din(w_dff_B_5lTzlez44_0),.dout(w_dff_B_2fehSlEE1_0),.clk(gclk));
	jdff dff_B_VUAjNiRH7_1(.din(n1053),.dout(w_dff_B_VUAjNiRH7_1),.clk(gclk));
	jdff dff_A_CzjPq7vf6_1(.dout(w_n800_3[1]),.din(w_dff_A_CzjPq7vf6_1),.clk(gclk));
	jdff dff_A_1RpyB4Tt6_2(.dout(w_n800_3[2]),.din(w_dff_A_1RpyB4Tt6_2),.clk(gclk));
	jdff dff_A_Lb63Q02A7_2(.dout(w_dff_A_1RpyB4Tt6_2),.din(w_dff_A_Lb63Q02A7_2),.clk(gclk));
	jdff dff_B_bkMId1lU2_1(.din(n1066),.dout(w_dff_B_bkMId1lU2_1),.clk(gclk));
	jdff dff_B_B1mY836K8_1(.din(w_dff_B_bkMId1lU2_1),.dout(w_dff_B_B1mY836K8_1),.clk(gclk));
	jdff dff_B_tdonufCY7_1(.din(w_dff_B_B1mY836K8_1),.dout(w_dff_B_tdonufCY7_1),.clk(gclk));
	jdff dff_B_7VECIvT16_1(.din(w_dff_B_tdonufCY7_1),.dout(w_dff_B_7VECIvT16_1),.clk(gclk));
	jdff dff_B_g9YK2ECl3_1(.din(w_dff_B_7VECIvT16_1),.dout(w_dff_B_g9YK2ECl3_1),.clk(gclk));
	jdff dff_B_66krYkky0_1(.din(w_dff_B_g9YK2ECl3_1),.dout(w_dff_B_66krYkky0_1),.clk(gclk));
	jdff dff_B_CL5gt7K56_1(.din(w_dff_B_66krYkky0_1),.dout(w_dff_B_CL5gt7K56_1),.clk(gclk));
	jdff dff_B_YBHM59qu6_1(.din(w_dff_B_CL5gt7K56_1),.dout(w_dff_B_YBHM59qu6_1),.clk(gclk));
	jdff dff_B_cCAeGkO51_1(.din(w_dff_B_YBHM59qu6_1),.dout(w_dff_B_cCAeGkO51_1),.clk(gclk));
	jdff dff_B_kyj8czcF3_1(.din(w_dff_B_cCAeGkO51_1),.dout(w_dff_B_kyj8czcF3_1),.clk(gclk));
	jdff dff_B_afQvGX8Q3_1(.din(w_dff_B_kyj8czcF3_1),.dout(w_dff_B_afQvGX8Q3_1),.clk(gclk));
	jdff dff_B_e1pr8F9p2_1(.din(w_dff_B_afQvGX8Q3_1),.dout(w_dff_B_e1pr8F9p2_1),.clk(gclk));
	jdff dff_B_8cMfT4eI0_1(.din(n1067),.dout(w_dff_B_8cMfT4eI0_1),.clk(gclk));
	jdff dff_A_jxmC1sKZ1_0(.dout(w_n854_4[0]),.din(w_dff_A_jxmC1sKZ1_0),.clk(gclk));
	jdff dff_A_830J17vn4_0(.dout(w_dff_A_jxmC1sKZ1_0),.din(w_dff_A_830J17vn4_0),.clk(gclk));
	jdff dff_A_WKrrakNZ0_0(.dout(w_dff_A_830J17vn4_0),.din(w_dff_A_WKrrakNZ0_0),.clk(gclk));
	jdff dff_A_L9wK2kU57_0(.dout(w_dff_A_WKrrakNZ0_0),.din(w_dff_A_L9wK2kU57_0),.clk(gclk));
	jdff dff_A_Hk6TBfrL2_0(.dout(w_dff_A_L9wK2kU57_0),.din(w_dff_A_Hk6TBfrL2_0),.clk(gclk));
	jdff dff_A_paDHeFq52_0(.dout(w_dff_A_Hk6TBfrL2_0),.din(w_dff_A_paDHeFq52_0),.clk(gclk));
	jdff dff_A_7k4NVCHH8_0(.dout(w_dff_A_paDHeFq52_0),.din(w_dff_A_7k4NVCHH8_0),.clk(gclk));
	jdff dff_B_cUkosmGA6_1(.din(n1063),.dout(w_dff_B_cUkosmGA6_1),.clk(gclk));
	jdff dff_B_jLkq5yPJ4_1(.din(w_dff_B_cUkosmGA6_1),.dout(w_dff_B_jLkq5yPJ4_1),.clk(gclk));
	jdff dff_B_ukQxG9DW5_2(.din(G37),.dout(w_dff_B_ukQxG9DW5_2),.clk(gclk));
	jdff dff_B_0hJPXdL73_1(.din(n1075),.dout(w_dff_B_0hJPXdL73_1),.clk(gclk));
	jdff dff_B_0w1RXKKs7_1(.din(w_dff_B_0hJPXdL73_1),.dout(w_dff_B_0w1RXKKs7_1),.clk(gclk));
	jdff dff_B_T1A0bSTN8_1(.din(w_dff_B_0w1RXKKs7_1),.dout(w_dff_B_T1A0bSTN8_1),.clk(gclk));
	jdff dff_B_AOw2XQ8g8_1(.din(w_dff_B_T1A0bSTN8_1),.dout(w_dff_B_AOw2XQ8g8_1),.clk(gclk));
	jdff dff_B_iXIiX3Fa9_1(.din(w_dff_B_AOw2XQ8g8_1),.dout(w_dff_B_iXIiX3Fa9_1),.clk(gclk));
	jdff dff_B_iw4G9YfW7_1(.din(w_dff_B_iXIiX3Fa9_1),.dout(w_dff_B_iw4G9YfW7_1),.clk(gclk));
	jdff dff_B_lXQHtbLP6_1(.din(w_dff_B_iw4G9YfW7_1),.dout(w_dff_B_lXQHtbLP6_1),.clk(gclk));
	jdff dff_B_0p0r8dTy5_1(.din(w_dff_B_lXQHtbLP6_1),.dout(w_dff_B_0p0r8dTy5_1),.clk(gclk));
	jdff dff_B_HcPIsBDU7_1(.din(w_dff_B_0p0r8dTy5_1),.dout(w_dff_B_HcPIsBDU7_1),.clk(gclk));
	jdff dff_B_5E47tHTh1_1(.din(w_dff_B_HcPIsBDU7_1),.dout(w_dff_B_5E47tHTh1_1),.clk(gclk));
	jdff dff_B_Znv1cIZd9_1(.din(w_dff_B_5E47tHTh1_1),.dout(w_dff_B_Znv1cIZd9_1),.clk(gclk));
	jdff dff_B_5roB9hPP7_1(.din(n1072),.dout(w_dff_B_5roB9hPP7_1),.clk(gclk));
	jdff dff_B_ZC7hCloA9_1(.din(w_dff_B_5roB9hPP7_1),.dout(w_dff_B_ZC7hCloA9_1),.clk(gclk));
	jdff dff_A_apcP3Tg10_1(.dout(w_n852_8[1]),.din(w_dff_A_apcP3Tg10_1),.clk(gclk));
	jdff dff_A_2uzeD8po6_1(.dout(w_dff_A_apcP3Tg10_1),.din(w_dff_A_2uzeD8po6_1),.clk(gclk));
	jdff dff_A_sbXKNuc64_1(.dout(w_dff_A_2uzeD8po6_1),.din(w_dff_A_sbXKNuc64_1),.clk(gclk));
	jdff dff_A_PUv7y5HW9_1(.dout(w_dff_A_sbXKNuc64_1),.din(w_dff_A_PUv7y5HW9_1),.clk(gclk));
	jdff dff_A_v1eeMBvn0_1(.dout(w_dff_A_PUv7y5HW9_1),.din(w_dff_A_v1eeMBvn0_1),.clk(gclk));
	jdff dff_A_dX0ckGmA7_1(.dout(w_dff_A_v1eeMBvn0_1),.din(w_dff_A_dX0ckGmA7_1),.clk(gclk));
	jdff dff_A_uxSTdeKI9_1(.dout(w_dff_A_dX0ckGmA7_1),.din(w_dff_A_uxSTdeKI9_1),.clk(gclk));
	jdff dff_A_iMM9QvWc9_1(.dout(w_dff_A_uxSTdeKI9_1),.din(w_dff_A_iMM9QvWc9_1),.clk(gclk));
	jdff dff_A_H163rTMi4_1(.dout(w_dff_A_iMM9QvWc9_1),.din(w_dff_A_H163rTMi4_1),.clk(gclk));
	jdff dff_A_5VXQVjaE2_1(.dout(w_dff_A_H163rTMi4_1),.din(w_dff_A_5VXQVjaE2_1),.clk(gclk));
	jdff dff_A_v4yyboEx4_1(.dout(w_dff_A_5VXQVjaE2_1),.din(w_dff_A_v4yyboEx4_1),.clk(gclk));
	jdff dff_A_e0eMipcg4_1(.dout(w_dff_A_v4yyboEx4_1),.din(w_dff_A_e0eMipcg4_1),.clk(gclk));
	jdff dff_B_im5dFBrE5_2(.din(G20),.dout(w_dff_B_im5dFBrE5_2),.clk(gclk));
	jdff dff_A_xfvpJ84k2_1(.dout(w_G4089_8[1]),.din(w_dff_A_xfvpJ84k2_1),.clk(gclk));
	jdff dff_A_uAZ1J8Ip2_1(.dout(w_dff_A_xfvpJ84k2_1),.din(w_dff_A_uAZ1J8Ip2_1),.clk(gclk));
	jdff dff_A_bHC6A4543_1(.dout(w_dff_A_uAZ1J8Ip2_1),.din(w_dff_A_bHC6A4543_1),.clk(gclk));
	jdff dff_A_wW8clFLT8_1(.dout(w_dff_A_bHC6A4543_1),.din(w_dff_A_wW8clFLT8_1),.clk(gclk));
	jdff dff_A_QWxAQkT58_1(.dout(w_dff_A_wW8clFLT8_1),.din(w_dff_A_QWxAQkT58_1),.clk(gclk));
	jdff dff_A_Nzr8a2qN5_1(.dout(w_dff_A_QWxAQkT58_1),.din(w_dff_A_Nzr8a2qN5_1),.clk(gclk));
	jdff dff_A_LAKDsYHP8_1(.dout(w_dff_A_Nzr8a2qN5_1),.din(w_dff_A_LAKDsYHP8_1),.clk(gclk));
	jdff dff_A_RdLmMYTu7_1(.dout(w_dff_A_LAKDsYHP8_1),.din(w_dff_A_RdLmMYTu7_1),.clk(gclk));
	jdff dff_A_UBexyctJ2_1(.dout(w_dff_A_RdLmMYTu7_1),.din(w_dff_A_UBexyctJ2_1),.clk(gclk));
	jdff dff_A_n5yHaSaD6_1(.dout(w_dff_A_UBexyctJ2_1),.din(w_dff_A_n5yHaSaD6_1),.clk(gclk));
	jdff dff_A_NpbvhCOn5_1(.dout(w_dff_A_n5yHaSaD6_1),.din(w_dff_A_NpbvhCOn5_1),.clk(gclk));
	jdff dff_A_a3kVmaUn1_1(.dout(w_dff_A_NpbvhCOn5_1),.din(w_dff_A_a3kVmaUn1_1),.clk(gclk));
	jdff dff_B_e1qVRQzZ8_1(.din(n1084),.dout(w_dff_B_e1qVRQzZ8_1),.clk(gclk));
	jdff dff_B_22V7Vy6N1_1(.din(w_dff_B_e1qVRQzZ8_1),.dout(w_dff_B_22V7Vy6N1_1),.clk(gclk));
	jdff dff_B_IzrZfD424_1(.din(w_dff_B_22V7Vy6N1_1),.dout(w_dff_B_IzrZfD424_1),.clk(gclk));
	jdff dff_B_u978ur932_1(.din(w_dff_B_IzrZfD424_1),.dout(w_dff_B_u978ur932_1),.clk(gclk));
	jdff dff_B_d535fkPZ6_1(.din(w_dff_B_u978ur932_1),.dout(w_dff_B_d535fkPZ6_1),.clk(gclk));
	jdff dff_B_BpjImiYi7_1(.din(w_dff_B_d535fkPZ6_1),.dout(w_dff_B_BpjImiYi7_1),.clk(gclk));
	jdff dff_B_OGrMSw1B1_1(.din(w_dff_B_BpjImiYi7_1),.dout(w_dff_B_OGrMSw1B1_1),.clk(gclk));
	jdff dff_B_xFBCjbib8_1(.din(w_dff_B_OGrMSw1B1_1),.dout(w_dff_B_xFBCjbib8_1),.clk(gclk));
	jdff dff_B_rURzYWoP2_1(.din(w_dff_B_xFBCjbib8_1),.dout(w_dff_B_rURzYWoP2_1),.clk(gclk));
	jdff dff_B_9czpcr7Z2_1(.din(w_dff_B_rURzYWoP2_1),.dout(w_dff_B_9czpcr7Z2_1),.clk(gclk));
	jdff dff_B_S6YzImyS1_0(.din(n1086),.dout(w_dff_B_S6YzImyS1_0),.clk(gclk));
	jdff dff_B_a5h5n6Vd2_0(.din(w_dff_B_S6YzImyS1_0),.dout(w_dff_B_a5h5n6Vd2_0),.clk(gclk));
	jdff dff_B_x9LEJhtA0_1(.din(n1081),.dout(w_dff_B_x9LEJhtA0_1),.clk(gclk));
	jdff dff_B_JvDrFjIk7_1(.din(w_dff_B_x9LEJhtA0_1),.dout(w_dff_B_JvDrFjIk7_1),.clk(gclk));
	jdff dff_A_gC9GFFaA2_0(.dout(w_n852_7[0]),.din(w_dff_A_gC9GFFaA2_0),.clk(gclk));
	jdff dff_A_H7CjY4PM5_0(.dout(w_dff_A_gC9GFFaA2_0),.din(w_dff_A_H7CjY4PM5_0),.clk(gclk));
	jdff dff_A_zlhhaP7h6_0(.dout(w_dff_A_H7CjY4PM5_0),.din(w_dff_A_zlhhaP7h6_0),.clk(gclk));
	jdff dff_A_6cHSBxia6_0(.dout(w_dff_A_zlhhaP7h6_0),.din(w_dff_A_6cHSBxia6_0),.clk(gclk));
	jdff dff_A_4caa1qTa1_0(.dout(w_dff_A_6cHSBxia6_0),.din(w_dff_A_4caa1qTa1_0),.clk(gclk));
	jdff dff_A_09yBD5uR1_0(.dout(w_dff_A_4caa1qTa1_0),.din(w_dff_A_09yBD5uR1_0),.clk(gclk));
	jdff dff_A_0WovloHB4_0(.dout(w_dff_A_09yBD5uR1_0),.din(w_dff_A_0WovloHB4_0),.clk(gclk));
	jdff dff_A_DxwT3zI21_0(.dout(w_dff_A_0WovloHB4_0),.din(w_dff_A_DxwT3zI21_0),.clk(gclk));
	jdff dff_A_qBX3YmmR7_0(.dout(w_dff_A_DxwT3zI21_0),.din(w_dff_A_qBX3YmmR7_0),.clk(gclk));
	jdff dff_A_AyIjvPMV7_0(.dout(w_dff_A_qBX3YmmR7_0),.din(w_dff_A_AyIjvPMV7_0),.clk(gclk));
	jdff dff_A_iYgs8HQM4_2(.dout(w_n852_7[2]),.din(w_dff_A_iYgs8HQM4_2),.clk(gclk));
	jdff dff_A_tLZDn3Wx7_2(.dout(w_dff_A_iYgs8HQM4_2),.din(w_dff_A_tLZDn3Wx7_2),.clk(gclk));
	jdff dff_A_iAP1tBFO5_2(.dout(w_dff_A_tLZDn3Wx7_2),.din(w_dff_A_iAP1tBFO5_2),.clk(gclk));
	jdff dff_A_49aC9TyN1_2(.dout(w_dff_A_iAP1tBFO5_2),.din(w_dff_A_49aC9TyN1_2),.clk(gclk));
	jdff dff_A_swNPezMS9_2(.dout(w_dff_A_49aC9TyN1_2),.din(w_dff_A_swNPezMS9_2),.clk(gclk));
	jdff dff_A_XYFnRj8u9_2(.dout(w_dff_A_swNPezMS9_2),.din(w_dff_A_XYFnRj8u9_2),.clk(gclk));
	jdff dff_A_xmCOz98r2_2(.dout(w_dff_A_XYFnRj8u9_2),.din(w_dff_A_xmCOz98r2_2),.clk(gclk));
	jdff dff_A_wdETEzoP6_2(.dout(w_dff_A_xmCOz98r2_2),.din(w_dff_A_wdETEzoP6_2),.clk(gclk));
	jdff dff_A_Z3oUY14E9_2(.dout(w_dff_A_wdETEzoP6_2),.din(w_dff_A_Z3oUY14E9_2),.clk(gclk));
	jdff dff_A_VfOToTWh7_2(.dout(w_dff_A_Z3oUY14E9_2),.din(w_dff_A_VfOToTWh7_2),.clk(gclk));
	jdff dff_A_D7jBCDW84_2(.dout(w_dff_A_VfOToTWh7_2),.din(w_dff_A_D7jBCDW84_2),.clk(gclk));
	jdff dff_B_sd2ZVu9e6_2(.din(G17),.dout(w_dff_B_sd2ZVu9e6_2),.clk(gclk));
	jdff dff_A_pB4g1s7L5_0(.dout(w_G4089_7[0]),.din(w_dff_A_pB4g1s7L5_0),.clk(gclk));
	jdff dff_A_onfVLaOH9_0(.dout(w_dff_A_pB4g1s7L5_0),.din(w_dff_A_onfVLaOH9_0),.clk(gclk));
	jdff dff_A_Eiwuvmvc4_0(.dout(w_dff_A_onfVLaOH9_0),.din(w_dff_A_Eiwuvmvc4_0),.clk(gclk));
	jdff dff_A_bO9pOKDo4_0(.dout(w_dff_A_Eiwuvmvc4_0),.din(w_dff_A_bO9pOKDo4_0),.clk(gclk));
	jdff dff_A_BIeNcFBX7_0(.dout(w_dff_A_bO9pOKDo4_0),.din(w_dff_A_BIeNcFBX7_0),.clk(gclk));
	jdff dff_A_CUoMUWNW1_0(.dout(w_dff_A_BIeNcFBX7_0),.din(w_dff_A_CUoMUWNW1_0),.clk(gclk));
	jdff dff_A_Ih9IteqR9_0(.dout(w_dff_A_CUoMUWNW1_0),.din(w_dff_A_Ih9IteqR9_0),.clk(gclk));
	jdff dff_A_X2Qapz4v4_0(.dout(w_dff_A_Ih9IteqR9_0),.din(w_dff_A_X2Qapz4v4_0),.clk(gclk));
	jdff dff_A_y3Wiv0ee2_0(.dout(w_dff_A_X2Qapz4v4_0),.din(w_dff_A_y3Wiv0ee2_0),.clk(gclk));
	jdff dff_A_qpN8pgB39_2(.dout(w_G4089_7[2]),.din(w_dff_A_qpN8pgB39_2),.clk(gclk));
	jdff dff_A_NnKahwor1_2(.dout(w_dff_A_qpN8pgB39_2),.din(w_dff_A_NnKahwor1_2),.clk(gclk));
	jdff dff_A_0VzkEIZ50_2(.dout(w_dff_A_NnKahwor1_2),.din(w_dff_A_0VzkEIZ50_2),.clk(gclk));
	jdff dff_A_z6xmCqAD5_2(.dout(w_dff_A_0VzkEIZ50_2),.din(w_dff_A_z6xmCqAD5_2),.clk(gclk));
	jdff dff_A_Ja8TycIr8_2(.dout(w_dff_A_z6xmCqAD5_2),.din(w_dff_A_Ja8TycIr8_2),.clk(gclk));
	jdff dff_A_NeB8eP9O1_2(.dout(w_dff_A_Ja8TycIr8_2),.din(w_dff_A_NeB8eP9O1_2),.clk(gclk));
	jdff dff_A_os5MzVpX6_2(.dout(w_dff_A_NeB8eP9O1_2),.din(w_dff_A_os5MzVpX6_2),.clk(gclk));
	jdff dff_A_9NmrFACZ2_2(.dout(w_dff_A_os5MzVpX6_2),.din(w_dff_A_9NmrFACZ2_2),.clk(gclk));
	jdff dff_A_YIpNymjH5_2(.dout(w_dff_A_9NmrFACZ2_2),.din(w_dff_A_YIpNymjH5_2),.clk(gclk));
	jdff dff_A_7KEDcc1i1_2(.dout(w_dff_A_YIpNymjH5_2),.din(w_dff_A_7KEDcc1i1_2),.clk(gclk));
	jdff dff_A_xeiLnNYM0_2(.dout(w_dff_A_7KEDcc1i1_2),.din(w_dff_A_xeiLnNYM0_2),.clk(gclk));
	jdff dff_A_Ydf7G1MN5_2(.dout(w_dff_A_xeiLnNYM0_2),.din(w_dff_A_Ydf7G1MN5_2),.clk(gclk));
	jdff dff_B_lwxmTE3c0_0(.din(n1097),.dout(w_dff_B_lwxmTE3c0_0),.clk(gclk));
	jdff dff_B_m2KtoGiw9_0(.din(w_dff_B_lwxmTE3c0_0),.dout(w_dff_B_m2KtoGiw9_0),.clk(gclk));
	jdff dff_B_gDfP0Q7f7_0(.din(w_dff_B_m2KtoGiw9_0),.dout(w_dff_B_gDfP0Q7f7_0),.clk(gclk));
	jdff dff_B_77xP8QcO7_0(.din(w_dff_B_gDfP0Q7f7_0),.dout(w_dff_B_77xP8QcO7_0),.clk(gclk));
	jdff dff_B_ADUqRKjA4_0(.din(w_dff_B_77xP8QcO7_0),.dout(w_dff_B_ADUqRKjA4_0),.clk(gclk));
	jdff dff_B_dSkavKle9_0(.din(w_dff_B_ADUqRKjA4_0),.dout(w_dff_B_dSkavKle9_0),.clk(gclk));
	jdff dff_B_rTgsmJ0K2_0(.din(w_dff_B_dSkavKle9_0),.dout(w_dff_B_rTgsmJ0K2_0),.clk(gclk));
	jdff dff_B_Eu1dSeSi8_0(.din(w_dff_B_rTgsmJ0K2_0),.dout(w_dff_B_Eu1dSeSi8_0),.clk(gclk));
	jdff dff_B_Tit3b0uv4_0(.din(w_dff_B_Eu1dSeSi8_0),.dout(w_dff_B_Tit3b0uv4_0),.clk(gclk));
	jdff dff_B_rOZqIJ489_0(.din(w_dff_B_Tit3b0uv4_0),.dout(w_dff_B_rOZqIJ489_0),.clk(gclk));
	jdff dff_A_nEW9LA4a0_1(.dout(w_G4090_3[1]),.din(w_dff_A_nEW9LA4a0_1),.clk(gclk));
	jdff dff_A_POkQJsV80_2(.dout(w_G4090_3[2]),.din(w_dff_A_POkQJsV80_2),.clk(gclk));
	jdff dff_B_tQUug1ty3_2(.din(G70),.dout(w_dff_B_tQUug1ty3_2),.clk(gclk));
	jdff dff_B_GtnUh3fp5_1(.din(n1090),.dout(w_dff_B_GtnUh3fp5_1),.clk(gclk));
	jdff dff_A_vRa1EFPx1_1(.dout(w_n854_3[1]),.din(w_dff_A_vRa1EFPx1_1),.clk(gclk));
	jdff dff_A_7V3vbrfp1_1(.dout(w_dff_A_vRa1EFPx1_1),.din(w_dff_A_7V3vbrfp1_1),.clk(gclk));
	jdff dff_A_7cLK4wxq1_2(.dout(w_n854_3[2]),.din(w_dff_A_7cLK4wxq1_2),.clk(gclk));
	jdff dff_A_d4p14SI83_2(.dout(w_dff_A_7cLK4wxq1_2),.din(w_dff_A_d4p14SI83_2),.clk(gclk));
	jdff dff_A_wQvkC4ud0_2(.dout(w_dff_A_d4p14SI83_2),.din(w_dff_A_wQvkC4ud0_2),.clk(gclk));
	jdff dff_B_aGUeRP3L2_0(.din(n1105),.dout(w_dff_B_aGUeRP3L2_0),.clk(gclk));
	jdff dff_B_tuBnLgZo4_0(.din(w_dff_B_aGUeRP3L2_0),.dout(w_dff_B_tuBnLgZo4_0),.clk(gclk));
	jdff dff_B_we40hQC63_0(.din(w_dff_B_tuBnLgZo4_0),.dout(w_dff_B_we40hQC63_0),.clk(gclk));
	jdff dff_B_P0WeECj87_0(.din(w_dff_B_we40hQC63_0),.dout(w_dff_B_P0WeECj87_0),.clk(gclk));
	jdff dff_B_OQZLYPfR4_0(.din(w_dff_B_P0WeECj87_0),.dout(w_dff_B_OQZLYPfR4_0),.clk(gclk));
	jdff dff_B_0bSE72zb7_0(.din(w_dff_B_OQZLYPfR4_0),.dout(w_dff_B_0bSE72zb7_0),.clk(gclk));
	jdff dff_B_Sszl1lTC4_0(.din(w_dff_B_0bSE72zb7_0),.dout(w_dff_B_Sszl1lTC4_0),.clk(gclk));
	jdff dff_B_Mg1CfUbk9_0(.din(w_dff_B_Sszl1lTC4_0),.dout(w_dff_B_Mg1CfUbk9_0),.clk(gclk));
	jdff dff_B_DyFG6Q476_0(.din(w_dff_B_Mg1CfUbk9_0),.dout(w_dff_B_DyFG6Q476_0),.clk(gclk));
	jdff dff_B_2IaB2hQo2_0(.din(w_dff_B_DyFG6Q476_0),.dout(w_dff_B_2IaB2hQo2_0),.clk(gclk));
	jdff dff_B_Z7X0DKjP1_0(.din(w_dff_B_2IaB2hQo2_0),.dout(w_dff_B_Z7X0DKjP1_0),.clk(gclk));
	jdff dff_B_L0foX1gb2_0(.din(w_dff_B_Z7X0DKjP1_0),.dout(w_dff_B_L0foX1gb2_0),.clk(gclk));
	jdff dff_B_Zg1UhuNn4_0(.din(n1104),.dout(w_dff_B_Zg1UhuNn4_0),.clk(gclk));
	jdff dff_B_AbvrSSu94_1(.din(n1099),.dout(w_dff_B_AbvrSSu94_1),.clk(gclk));
	jdff dff_B_dHD2NsdS6_1(.din(w_dff_B_AbvrSSu94_1),.dout(w_dff_B_dHD2NsdS6_1),.clk(gclk));
	jdff dff_B_BhCxatF42_0(.din(n1114),.dout(w_dff_B_BhCxatF42_0),.clk(gclk));
	jdff dff_B_sjVkna3y0_0(.din(w_dff_B_BhCxatF42_0),.dout(w_dff_B_sjVkna3y0_0),.clk(gclk));
	jdff dff_B_faJmfSlV7_0(.din(w_dff_B_sjVkna3y0_0),.dout(w_dff_B_faJmfSlV7_0),.clk(gclk));
	jdff dff_B_JmoLRkOZ1_0(.din(w_dff_B_faJmfSlV7_0),.dout(w_dff_B_JmoLRkOZ1_0),.clk(gclk));
	jdff dff_B_ujjSmdMT7_0(.din(w_dff_B_JmoLRkOZ1_0),.dout(w_dff_B_ujjSmdMT7_0),.clk(gclk));
	jdff dff_B_dUuYIzS16_0(.din(w_dff_B_ujjSmdMT7_0),.dout(w_dff_B_dUuYIzS16_0),.clk(gclk));
	jdff dff_B_LJrJXStQ8_0(.din(w_dff_B_dUuYIzS16_0),.dout(w_dff_B_LJrJXStQ8_0),.clk(gclk));
	jdff dff_B_t34VBvls2_0(.din(w_dff_B_LJrJXStQ8_0),.dout(w_dff_B_t34VBvls2_0),.clk(gclk));
	jdff dff_B_4wdvpaih2_0(.din(w_dff_B_t34VBvls2_0),.dout(w_dff_B_4wdvpaih2_0),.clk(gclk));
	jdff dff_B_OKBEGDpY5_0(.din(n1113),.dout(w_dff_B_OKBEGDpY5_0),.clk(gclk));
	jdff dff_B_lLyMDWw12_1(.din(n1108),.dout(w_dff_B_lLyMDWw12_1),.clk(gclk));
	jdff dff_A_MDICiLQy1_0(.dout(w_n999_3[0]),.din(w_dff_A_MDICiLQy1_0),.clk(gclk));
	jdff dff_A_zPHzPfKF5_0(.dout(w_dff_A_MDICiLQy1_0),.din(w_dff_A_zPHzPfKF5_0),.clk(gclk));
	jdff dff_A_nw6sdVGv8_0(.dout(w_dff_A_zPHzPfKF5_0),.din(w_dff_A_nw6sdVGv8_0),.clk(gclk));
	jdff dff_A_ejV6WJxp7_1(.dout(w_n999_3[1]),.din(w_dff_A_ejV6WJxp7_1),.clk(gclk));
	jdff dff_A_aRx0CpwE4_1(.dout(w_dff_A_ejV6WJxp7_1),.din(w_dff_A_aRx0CpwE4_1),.clk(gclk));
	jdff dff_A_J7kLXnJZ0_1(.dout(w_dff_A_aRx0CpwE4_1),.din(w_dff_A_J7kLXnJZ0_1),.clk(gclk));
	jdff dff_A_iXFLeoAz1_1(.dout(w_dff_A_J7kLXnJZ0_1),.din(w_dff_A_iXFLeoAz1_1),.clk(gclk));
	jdff dff_A_auO0Ihs89_1(.dout(w_dff_A_iXFLeoAz1_1),.din(w_dff_A_auO0Ihs89_1),.clk(gclk));
	jdff dff_A_V9tpnX0W9_1(.dout(w_dff_A_auO0Ihs89_1),.din(w_dff_A_V9tpnX0W9_1),.clk(gclk));
	jdff dff_A_NcOedwtw7_0(.dout(w_G1689_4[0]),.din(w_dff_A_NcOedwtw7_0),.clk(gclk));
	jdff dff_A_HQ4yem6X0_0(.dout(w_dff_A_NcOedwtw7_0),.din(w_dff_A_HQ4yem6X0_0),.clk(gclk));
	jdff dff_A_wPirhIZM5_0(.dout(w_dff_A_HQ4yem6X0_0),.din(w_dff_A_wPirhIZM5_0),.clk(gclk));
	jdff dff_A_x6QrGI4k9_1(.dout(w_G1689_4[1]),.din(w_dff_A_x6QrGI4k9_1),.clk(gclk));
	jdff dff_A_dO9R75Pk8_1(.dout(w_dff_A_x6QrGI4k9_1),.din(w_dff_A_dO9R75Pk8_1),.clk(gclk));
	jdff dff_A_YReokgF71_1(.dout(w_dff_A_dO9R75Pk8_1),.din(w_dff_A_YReokgF71_1),.clk(gclk));
	jdff dff_A_kaPTMUid6_1(.dout(w_dff_A_YReokgF71_1),.din(w_dff_A_kaPTMUid6_1),.clk(gclk));
	jdff dff_A_hU8ufdTl1_1(.dout(w_dff_A_kaPTMUid6_1),.din(w_dff_A_hU8ufdTl1_1),.clk(gclk));
	jdff dff_B_iITIKDNb5_0(.din(n1123),.dout(w_dff_B_iITIKDNb5_0),.clk(gclk));
	jdff dff_B_XH9LBuJk1_0(.din(w_dff_B_iITIKDNb5_0),.dout(w_dff_B_XH9LBuJk1_0),.clk(gclk));
	jdff dff_B_Tpy8NYjg2_0(.din(w_dff_B_XH9LBuJk1_0),.dout(w_dff_B_Tpy8NYjg2_0),.clk(gclk));
	jdff dff_B_mQxmRu629_0(.din(w_dff_B_Tpy8NYjg2_0),.dout(w_dff_B_mQxmRu629_0),.clk(gclk));
	jdff dff_B_qdwiHKA33_0(.din(w_dff_B_mQxmRu629_0),.dout(w_dff_B_qdwiHKA33_0),.clk(gclk));
	jdff dff_B_IcOzOlfV6_0(.din(w_dff_B_qdwiHKA33_0),.dout(w_dff_B_IcOzOlfV6_0),.clk(gclk));
	jdff dff_B_afsLMNDS3_0(.din(w_dff_B_IcOzOlfV6_0),.dout(w_dff_B_afsLMNDS3_0),.clk(gclk));
	jdff dff_B_2fcslUvf1_0(.din(w_dff_B_afsLMNDS3_0),.dout(w_dff_B_2fcslUvf1_0),.clk(gclk));
	jdff dff_B_K1KunLx38_0(.din(w_dff_B_2fcslUvf1_0),.dout(w_dff_B_K1KunLx38_0),.clk(gclk));
	jdff dff_B_LuGLwxXH5_0(.din(w_dff_B_K1KunLx38_0),.dout(w_dff_B_LuGLwxXH5_0),.clk(gclk));
	jdff dff_B_OL3NLugM8_0(.din(n1122),.dout(w_dff_B_OL3NLugM8_0),.clk(gclk));
	jdff dff_B_201JWcL95_1(.din(n1117),.dout(w_dff_B_201JWcL95_1),.clk(gclk));
	jdff dff_B_mWlLAJF08_1(.din(w_dff_B_201JWcL95_1),.dout(w_dff_B_mWlLAJF08_1),.clk(gclk));
	jdff dff_B_4Z6Nypry4_1(.din(w_dff_B_mWlLAJF08_1),.dout(w_dff_B_4Z6Nypry4_1),.clk(gclk));
	jdff dff_A_mbCLFJ1C0_0(.dout(w_G137_8[0]),.din(w_dff_A_mbCLFJ1C0_0),.clk(gclk));
	jdff dff_A_APz6jERG5_2(.dout(w_G137_8[2]),.din(w_dff_A_APz6jERG5_2),.clk(gclk));
	jdff dff_A_rl5AWjRP2_2(.dout(w_dff_A_APz6jERG5_2),.din(w_dff_A_rl5AWjRP2_2),.clk(gclk));
	jdff dff_A_3m7ZcVHv3_2(.dout(w_dff_A_rl5AWjRP2_2),.din(w_dff_A_3m7ZcVHv3_2),.clk(gclk));
	jdff dff_B_bjQmrv3o6_0(.din(n1132),.dout(w_dff_B_bjQmrv3o6_0),.clk(gclk));
	jdff dff_B_9PWobMtC4_0(.din(w_dff_B_bjQmrv3o6_0),.dout(w_dff_B_9PWobMtC4_0),.clk(gclk));
	jdff dff_B_cMl2pxRp0_0(.din(w_dff_B_9PWobMtC4_0),.dout(w_dff_B_cMl2pxRp0_0),.clk(gclk));
	jdff dff_B_jKGfgZXT8_0(.din(w_dff_B_cMl2pxRp0_0),.dout(w_dff_B_jKGfgZXT8_0),.clk(gclk));
	jdff dff_B_bi8BQgi44_0(.din(w_dff_B_jKGfgZXT8_0),.dout(w_dff_B_bi8BQgi44_0),.clk(gclk));
	jdff dff_B_LZM14I1d0_0(.din(w_dff_B_bi8BQgi44_0),.dout(w_dff_B_LZM14I1d0_0),.clk(gclk));
	jdff dff_B_XrJbQawW4_0(.din(w_dff_B_LZM14I1d0_0),.dout(w_dff_B_XrJbQawW4_0),.clk(gclk));
	jdff dff_B_eP20ZFRJ2_0(.din(w_dff_B_XrJbQawW4_0),.dout(w_dff_B_eP20ZFRJ2_0),.clk(gclk));
	jdff dff_B_RF74xTuM8_0(.din(w_dff_B_eP20ZFRJ2_0),.dout(w_dff_B_RF74xTuM8_0),.clk(gclk));
	jdff dff_B_g3a2nV270_0(.din(w_dff_B_RF74xTuM8_0),.dout(w_dff_B_g3a2nV270_0),.clk(gclk));
	jdff dff_B_mzqMQWYO7_0(.din(w_dff_B_g3a2nV270_0),.dout(w_dff_B_mzqMQWYO7_0),.clk(gclk));
	jdff dff_B_TRI8VtAe1_0(.din(n1131),.dout(w_dff_B_TRI8VtAe1_0),.clk(gclk));
	jdff dff_B_rNLC0A6b9_1(.din(n1126),.dout(w_dff_B_rNLC0A6b9_1),.clk(gclk));
	jdff dff_A_I7cFGMOk0_0(.dout(w_n993_3[0]),.din(w_dff_A_I7cFGMOk0_0),.clk(gclk));
	jdff dff_A_5zgclu6e2_0(.dout(w_dff_A_I7cFGMOk0_0),.din(w_dff_A_5zgclu6e2_0),.clk(gclk));
	jdff dff_A_WrwQKUNH7_1(.dout(w_n993_3[1]),.din(w_dff_A_WrwQKUNH7_1),.clk(gclk));
	jdff dff_B_QNE4u8UD2_1(.din(n1135),.dout(w_dff_B_QNE4u8UD2_1),.clk(gclk));
	jdff dff_B_2OibqZSg5_1(.din(w_dff_B_QNE4u8UD2_1),.dout(w_dff_B_2OibqZSg5_1),.clk(gclk));
	jdff dff_B_cmJ4Sanv8_1(.din(w_dff_B_2OibqZSg5_1),.dout(w_dff_B_cmJ4Sanv8_1),.clk(gclk));
	jdff dff_B_GZNcX2g00_1(.din(w_dff_B_cmJ4Sanv8_1),.dout(w_dff_B_GZNcX2g00_1),.clk(gclk));
	jdff dff_B_ZcOcE4TC4_1(.din(w_dff_B_GZNcX2g00_1),.dout(w_dff_B_ZcOcE4TC4_1),.clk(gclk));
	jdff dff_B_DqEEM4R79_1(.din(w_dff_B_ZcOcE4TC4_1),.dout(w_dff_B_DqEEM4R79_1),.clk(gclk));
	jdff dff_B_EmpDHZlQ2_1(.din(w_dff_B_DqEEM4R79_1),.dout(w_dff_B_EmpDHZlQ2_1),.clk(gclk));
	jdff dff_B_OQ8RAhaU2_1(.din(w_dff_B_EmpDHZlQ2_1),.dout(w_dff_B_OQ8RAhaU2_1),.clk(gclk));
	jdff dff_B_QW1gJaCr4_1(.din(w_dff_B_OQ8RAhaU2_1),.dout(w_dff_B_QW1gJaCr4_1),.clk(gclk));
	jdff dff_B_cZtruJZp8_1(.din(w_dff_B_QW1gJaCr4_1),.dout(w_dff_B_cZtruJZp8_1),.clk(gclk));
	jdff dff_B_9dKtiNDO5_1(.din(w_dff_B_cZtruJZp8_1),.dout(w_dff_B_9dKtiNDO5_1),.clk(gclk));
	jdff dff_B_O8UO2SZW0_1(.din(w_dff_B_9dKtiNDO5_1),.dout(w_dff_B_O8UO2SZW0_1),.clk(gclk));
	jdff dff_B_fOThIB7Q0_1(.din(n1136),.dout(w_dff_B_fOThIB7Q0_1),.clk(gclk));
	jdff dff_B_vdVXqaMK2_1(.din(w_dff_B_fOThIB7Q0_1),.dout(w_dff_B_vdVXqaMK2_1),.clk(gclk));
	jdff dff_B_hxRqJRzm1_1(.din(w_dff_B_vdVXqaMK2_1),.dout(w_dff_B_hxRqJRzm1_1),.clk(gclk));
	jdff dff_B_kaGws2ym7_1(.din(w_dff_B_hxRqJRzm1_1),.dout(w_dff_B_kaGws2ym7_1),.clk(gclk));
	jdff dff_B_6EJG7CkC3_1(.din(w_dff_B_kaGws2ym7_1),.dout(w_dff_B_6EJG7CkC3_1),.clk(gclk));
	jdff dff_B_lvafxM903_1(.din(w_dff_B_6EJG7CkC3_1),.dout(w_dff_B_lvafxM903_1),.clk(gclk));
	jdff dff_B_aJ4zOciI9_1(.din(w_dff_B_lvafxM903_1),.dout(w_dff_B_aJ4zOciI9_1),.clk(gclk));
	jdff dff_B_8CPFJZ6j1_1(.din(w_dff_B_aJ4zOciI9_1),.dout(w_dff_B_8CPFJZ6j1_1),.clk(gclk));
	jdff dff_B_0SJciPGz8_1(.din(w_dff_B_8CPFJZ6j1_1),.dout(w_dff_B_0SJciPGz8_1),.clk(gclk));
	jdff dff_B_IcIzwzrP5_1(.din(w_dff_B_0SJciPGz8_1),.dout(w_dff_B_IcIzwzrP5_1),.clk(gclk));
	jdff dff_B_aUAbdcNR7_1(.din(w_dff_B_IcIzwzrP5_1),.dout(w_dff_B_aUAbdcNR7_1),.clk(gclk));
	jdff dff_B_6ZKop9ww7_1(.din(w_dff_B_aUAbdcNR7_1),.dout(w_dff_B_6ZKop9ww7_1),.clk(gclk));
	jdff dff_B_039QYSRB1_1(.din(w_dff_B_6ZKop9ww7_1),.dout(w_dff_B_039QYSRB1_1),.clk(gclk));
	jdff dff_B_beWqPsAs9_0(.din(n1138),.dout(w_dff_B_beWqPsAs9_0),.clk(gclk));
	jdff dff_B_SCNZweY59_1(.din(n811),.dout(w_dff_B_SCNZweY59_1),.clk(gclk));
	jdff dff_B_VnrBFmea0_1(.din(w_dff_B_SCNZweY59_1),.dout(w_dff_B_VnrBFmea0_1),.clk(gclk));
	jdff dff_B_WwWbbkQL5_1(.din(w_dff_B_VnrBFmea0_1),.dout(w_dff_B_WwWbbkQL5_1),.clk(gclk));
	jdff dff_B_6tLdqHvS2_1(.din(w_dff_B_WwWbbkQL5_1),.dout(w_dff_B_6tLdqHvS2_1),.clk(gclk));
	jdff dff_B_y8BTqAfv6_1(.din(w_dff_B_6tLdqHvS2_1),.dout(w_dff_B_y8BTqAfv6_1),.clk(gclk));
	jdff dff_B_9RWlcmWY9_1(.din(w_dff_B_y8BTqAfv6_1),.dout(w_dff_B_9RWlcmWY9_1),.clk(gclk));
	jdff dff_B_DoV4iL8k7_0(.din(n830),.dout(w_dff_B_DoV4iL8k7_0),.clk(gclk));
	jdff dff_B_48oF9AZD9_0(.din(w_dff_B_DoV4iL8k7_0),.dout(w_dff_B_48oF9AZD9_0),.clk(gclk));
	jdff dff_B_6v9iZpdS7_0(.din(w_dff_B_48oF9AZD9_0),.dout(w_dff_B_6v9iZpdS7_0),.clk(gclk));
	jdff dff_B_YOF0tylv7_0(.din(w_dff_B_6v9iZpdS7_0),.dout(w_dff_B_YOF0tylv7_0),.clk(gclk));
	jdff dff_B_TIa6Cguv5_0(.din(w_dff_B_YOF0tylv7_0),.dout(w_dff_B_TIa6Cguv5_0),.clk(gclk));
	jdff dff_B_sL7vJs5x6_0(.din(w_dff_B_TIa6Cguv5_0),.dout(w_dff_B_sL7vJs5x6_0),.clk(gclk));
	jdff dff_A_s0mWYLZx6_1(.dout(w_n445_0[1]),.din(w_dff_A_s0mWYLZx6_1),.clk(gclk));
	jdff dff_B_F9EoP2rl4_1(.din(n441),.dout(w_dff_B_F9EoP2rl4_1),.clk(gclk));
	jdff dff_B_MTFsqagk5_1(.din(n822),.dout(w_dff_B_MTFsqagk5_1),.clk(gclk));
	jdff dff_B_z3Nd8qxk9_1(.din(w_dff_B_MTFsqagk5_1),.dout(w_dff_B_z3Nd8qxk9_1),.clk(gclk));
	jdff dff_B_LjCjvAaW5_1(.din(w_dff_B_z3Nd8qxk9_1),.dout(w_dff_B_LjCjvAaW5_1),.clk(gclk));
	jdff dff_B_sedO53ka2_1(.din(w_dff_B_LjCjvAaW5_1),.dout(w_dff_B_sedO53ka2_1),.clk(gclk));
	jdff dff_B_c2WqjHWj4_1(.din(G52),.dout(w_dff_B_c2WqjHWj4_1),.clk(gclk));
	jdff dff_B_JwiEoX8s2_1(.din(w_dff_B_c2WqjHWj4_1),.dout(w_dff_B_JwiEoX8s2_1),.clk(gclk));
	jdff dff_B_Tala5Q3g3_1(.din(n864),.dout(w_dff_B_Tala5Q3g3_1),.clk(gclk));
	jdff dff_B_QZpvcZaB4_1(.din(w_dff_B_Tala5Q3g3_1),.dout(w_dff_B_QZpvcZaB4_1),.clk(gclk));
	jdff dff_B_TyevNExH3_1(.din(w_dff_B_QZpvcZaB4_1),.dout(w_dff_B_TyevNExH3_1),.clk(gclk));
	jdff dff_B_laLYCMTy3_1(.din(w_dff_B_TyevNExH3_1),.dout(w_dff_B_laLYCMTy3_1),.clk(gclk));
	jdff dff_B_NvWPEA940_1(.din(w_dff_B_laLYCMTy3_1),.dout(w_dff_B_NvWPEA940_1),.clk(gclk));
	jdff dff_B_GfAwnbcw4_1(.din(w_dff_B_NvWPEA940_1),.dout(w_dff_B_GfAwnbcw4_1),.clk(gclk));
	jdff dff_B_ZsiKmdKd1_1(.din(w_dff_B_GfAwnbcw4_1),.dout(w_dff_B_ZsiKmdKd1_1),.clk(gclk));
	jdff dff_B_GtDlaz1j4_0(.din(n874),.dout(w_dff_B_GtDlaz1j4_0),.clk(gclk));
	jdff dff_B_0z7eOQJI9_0(.din(w_dff_B_GtDlaz1j4_0),.dout(w_dff_B_0z7eOQJI9_0),.clk(gclk));
	jdff dff_B_dyc5tWD73_0(.din(w_dff_B_0z7eOQJI9_0),.dout(w_dff_B_dyc5tWD73_0),.clk(gclk));
	jdff dff_B_FU3Szuor4_0(.din(w_dff_B_dyc5tWD73_0),.dout(w_dff_B_FU3Szuor4_0),.clk(gclk));
	jdff dff_B_sIoewJFH8_0(.din(w_dff_B_FU3Szuor4_0),.dout(w_dff_B_sIoewJFH8_0),.clk(gclk));
	jdff dff_B_TK1m8UMz9_0(.din(w_dff_B_sIoewJFH8_0),.dout(w_dff_B_TK1m8UMz9_0),.clk(gclk));
	jdff dff_B_myhdTuYj6_0(.din(w_dff_B_TK1m8UMz9_0),.dout(w_dff_B_myhdTuYj6_0),.clk(gclk));
	jdff dff_B_1JyXEtsm3_1(.din(n466),.dout(w_dff_B_1JyXEtsm3_1),.clk(gclk));
	jdff dff_B_SauEUFGf6_1(.din(G122),.dout(w_dff_B_SauEUFGf6_1),.clk(gclk));
	jdff dff_B_c5kHQJeJ9_1(.din(w_dff_B_SauEUFGf6_1),.dout(w_dff_B_c5kHQJeJ9_1),.clk(gclk));
	jdff dff_B_fJjEArNj5_2(.din(G170),.dout(w_dff_B_fJjEArNj5_2),.clk(gclk));
	jdff dff_B_FU2GyNtp4_2(.din(G200),.dout(w_dff_B_FU2GyNtp4_2),.clk(gclk));
	jdff dff_B_P7lro8k06_2(.din(w_dff_B_FU2GyNtp4_2),.dout(w_dff_B_P7lro8k06_2),.clk(gclk));
	jdff dff_B_kRSMxXCm1_0(.din(n1150),.dout(w_dff_B_kRSMxXCm1_0),.clk(gclk));
	jdff dff_B_M1dIrjKe6_0(.din(w_dff_B_kRSMxXCm1_0),.dout(w_dff_B_M1dIrjKe6_0),.clk(gclk));
	jdff dff_B_wrTZK3aY2_0(.din(w_dff_B_M1dIrjKe6_0),.dout(w_dff_B_wrTZK3aY2_0),.clk(gclk));
	jdff dff_B_X8HOIuIg7_0(.din(w_dff_B_wrTZK3aY2_0),.dout(w_dff_B_X8HOIuIg7_0),.clk(gclk));
	jdff dff_B_cOEWvLM80_0(.din(w_dff_B_X8HOIuIg7_0),.dout(w_dff_B_cOEWvLM80_0),.clk(gclk));
	jdff dff_B_C2RHxMHD5_0(.din(w_dff_B_cOEWvLM80_0),.dout(w_dff_B_C2RHxMHD5_0),.clk(gclk));
	jdff dff_B_nYyjJrNm4_0(.din(w_dff_B_C2RHxMHD5_0),.dout(w_dff_B_nYyjJrNm4_0),.clk(gclk));
	jdff dff_B_uERNU9TH2_0(.din(w_dff_B_nYyjJrNm4_0),.dout(w_dff_B_uERNU9TH2_0),.clk(gclk));
	jdff dff_B_7VhNgJT62_0(.din(w_dff_B_uERNU9TH2_0),.dout(w_dff_B_7VhNgJT62_0),.clk(gclk));
	jdff dff_B_Nxu03oUQ0_0(.din(n1149),.dout(w_dff_B_Nxu03oUQ0_0),.clk(gclk));
	jdff dff_B_Qku3HVSq6_2(.din(G158),.dout(w_dff_B_Qku3HVSq6_2),.clk(gclk));
	jdff dff_B_F43lJ4044_2(.din(G188),.dout(w_dff_B_F43lJ4044_2),.clk(gclk));
	jdff dff_B_fBz5XXFX2_2(.din(w_dff_B_F43lJ4044_2),.dout(w_dff_B_fBz5XXFX2_2),.clk(gclk));
	jdff dff_B_6d5lY3U59_1(.din(n1144),.dout(w_dff_B_6d5lY3U59_1),.clk(gclk));
	jdff dff_B_aJo1nRbC1_1(.din(n897),.dout(w_dff_B_aJo1nRbC1_1),.clk(gclk));
	jdff dff_B_bgvZjZNJ3_1(.din(w_dff_B_aJo1nRbC1_1),.dout(w_dff_B_bgvZjZNJ3_1),.clk(gclk));
	jdff dff_B_73awkLfH9_1(.din(w_dff_B_bgvZjZNJ3_1),.dout(w_dff_B_73awkLfH9_1),.clk(gclk));
	jdff dff_B_aqObUz5T9_1(.din(w_dff_B_73awkLfH9_1),.dout(w_dff_B_aqObUz5T9_1),.clk(gclk));
	jdff dff_B_MKcm9QhE1_0(.din(n904),.dout(w_dff_B_MKcm9QhE1_0),.clk(gclk));
	jdff dff_B_uYkATdKd6_0(.din(w_dff_B_MKcm9QhE1_0),.dout(w_dff_B_uYkATdKd6_0),.clk(gclk));
	jdff dff_B_vNOiyNA02_0(.din(w_dff_B_uYkATdKd6_0),.dout(w_dff_B_vNOiyNA02_0),.clk(gclk));
	jdff dff_B_D2gjCNcq2_0(.din(w_dff_B_vNOiyNA02_0),.dout(w_dff_B_D2gjCNcq2_0),.clk(gclk));
	jdff dff_B_aMvWkg9f4_1(.din(n477),.dout(w_dff_B_aMvWkg9f4_1),.clk(gclk));
	jdff dff_A_dBRegjB43_0(.dout(w_n901_0[0]),.din(w_dff_A_dBRegjB43_0),.clk(gclk));
	jdff dff_A_F6Ryisq53_0(.dout(w_dff_A_dBRegjB43_0),.din(w_dff_A_F6Ryisq53_0),.clk(gclk));
	jdff dff_B_zW1FaUDe4_1(.din(G126),.dout(w_dff_B_zW1FaUDe4_1),.clk(gclk));
	jdff dff_B_uc5mNuws3_1(.din(w_dff_B_zW1FaUDe4_1),.dout(w_dff_B_uc5mNuws3_1),.clk(gclk));
	jdff dff_A_mnVniqVR9_1(.dout(w_n1007_3[1]),.din(w_dff_A_mnVniqVR9_1),.clk(gclk));
	jdff dff_A_U9FwaGHB7_1(.dout(w_dff_A_mnVniqVR9_1),.din(w_dff_A_U9FwaGHB7_1),.clk(gclk));
	jdff dff_A_hp6tJ3RD6_1(.dout(w_dff_A_U9FwaGHB7_1),.din(w_dff_A_hp6tJ3RD6_1),.clk(gclk));
	jdff dff_A_ARkK3bjp4_1(.dout(w_dff_A_hp6tJ3RD6_1),.din(w_dff_A_ARkK3bjp4_1),.clk(gclk));
	jdff dff_B_YpfmQm0m0_1(.din(n762),.dout(w_dff_B_YpfmQm0m0_1),.clk(gclk));
	jdff dff_B_lNitwqbK2_1(.din(w_dff_B_YpfmQm0m0_1),.dout(w_dff_B_lNitwqbK2_1),.clk(gclk));
	jdff dff_B_qdjYAWkp4_1(.din(w_dff_B_lNitwqbK2_1),.dout(w_dff_B_qdjYAWkp4_1),.clk(gclk));
	jdff dff_B_WKaXesSI6_1(.din(w_dff_B_qdjYAWkp4_1),.dout(w_dff_B_WKaXesSI6_1),.clk(gclk));
	jdff dff_B_KfCYvZFK0_0(.din(n773),.dout(w_dff_B_KfCYvZFK0_0),.clk(gclk));
	jdff dff_B_fyau8eTK4_0(.din(w_dff_B_KfCYvZFK0_0),.dout(w_dff_B_fyau8eTK4_0),.clk(gclk));
	jdff dff_B_bccpTALs6_0(.din(w_dff_B_fyau8eTK4_0),.dout(w_dff_B_bccpTALs6_0),.clk(gclk));
	jdff dff_B_xvh3OphK0_0(.din(w_dff_B_bccpTALs6_0),.dout(w_dff_B_xvh3OphK0_0),.clk(gclk));
	jdff dff_B_nek1dyeV9_1(.din(n382),.dout(w_dff_B_nek1dyeV9_1),.clk(gclk));
	jdff dff_B_BWMxTbrC1_0(.din(n769),.dout(w_dff_B_BWMxTbrC1_0),.clk(gclk));
	jdff dff_B_PKKUPnJQ6_0(.din(w_dff_B_BWMxTbrC1_0),.dout(w_dff_B_PKKUPnJQ6_0),.clk(gclk));
	jdff dff_B_bvUdY8NE0_0(.din(w_dff_B_PKKUPnJQ6_0),.dout(w_dff_B_bvUdY8NE0_0),.clk(gclk));
	jdff dff_A_syCrgftP0_0(.dout(w_n753_1[0]),.din(w_dff_A_syCrgftP0_0),.clk(gclk));
	jdff dff_A_819bBhEI4_0(.dout(w_dff_A_syCrgftP0_0),.din(w_dff_A_819bBhEI4_0),.clk(gclk));
	jdff dff_A_wdVqBrym4_0(.dout(w_dff_A_819bBhEI4_0),.din(w_dff_A_wdVqBrym4_0),.clk(gclk));
	jdff dff_A_hurffN830_0(.dout(w_dff_A_wdVqBrym4_0),.din(w_dff_A_hurffN830_0),.clk(gclk));
	jdff dff_A_5qpZxzkn1_0(.dout(w_G4091_5[0]),.din(w_dff_A_5qpZxzkn1_0),.clk(gclk));
	jdff dff_A_GAPszGMA6_0(.dout(w_dff_A_5qpZxzkn1_0),.din(w_dff_A_GAPszGMA6_0),.clk(gclk));
	jdff dff_B_V4cX5wPa7_1(.din(G129),.dout(w_dff_B_V4cX5wPa7_1),.clk(gclk));
	jdff dff_B_EDicO3ac1_1(.din(w_dff_B_V4cX5wPa7_1),.dout(w_dff_B_EDicO3ac1_1),.clk(gclk));
	jdff dff_A_qPIwHP0t4_1(.dout(w_G137_7[1]),.din(w_dff_A_qPIwHP0t4_1),.clk(gclk));
	jdff dff_A_nyqAEYAd7_1(.dout(w_dff_A_qPIwHP0t4_1),.din(w_dff_A_nyqAEYAd7_1),.clk(gclk));
	jdff dff_A_ZkMZMwwK5_1(.dout(w_dff_A_nyqAEYAd7_1),.din(w_dff_A_ZkMZMwwK5_1),.clk(gclk));
	jdff dff_A_w6xNupWn1_2(.dout(w_G137_7[2]),.din(w_dff_A_w6xNupWn1_2),.clk(gclk));
	jdff dff_A_LHfbv8a61_2(.dout(w_dff_A_w6xNupWn1_2),.din(w_dff_A_LHfbv8a61_2),.clk(gclk));
	jdff dff_A_nslVg6tw9_0(.dout(w_G137_2[0]),.din(w_dff_A_nslVg6tw9_0),.clk(gclk));
	jdff dff_A_qWjcXWzl4_1(.dout(w_G137_2[1]),.din(w_dff_A_qWjcXWzl4_1),.clk(gclk));
	jdff dff_B_84nPq5fe2_0(.din(n1159),.dout(w_dff_B_84nPq5fe2_0),.clk(gclk));
	jdff dff_B_BSRtKwJs3_0(.din(w_dff_B_84nPq5fe2_0),.dout(w_dff_B_BSRtKwJs3_0),.clk(gclk));
	jdff dff_B_8tJOCkGq1_0(.din(w_dff_B_BSRtKwJs3_0),.dout(w_dff_B_8tJOCkGq1_0),.clk(gclk));
	jdff dff_B_CpK3WHEH9_0(.din(w_dff_B_8tJOCkGq1_0),.dout(w_dff_B_CpK3WHEH9_0),.clk(gclk));
	jdff dff_B_WOn2ylnQ3_0(.din(w_dff_B_CpK3WHEH9_0),.dout(w_dff_B_WOn2ylnQ3_0),.clk(gclk));
	jdff dff_B_HL7G0cZb0_0(.din(w_dff_B_WOn2ylnQ3_0),.dout(w_dff_B_HL7G0cZb0_0),.clk(gclk));
	jdff dff_B_iGPXOkeR0_0(.din(w_dff_B_HL7G0cZb0_0),.dout(w_dff_B_iGPXOkeR0_0),.clk(gclk));
	jdff dff_B_yWfnQGqC1_0(.din(w_dff_B_iGPXOkeR0_0),.dout(w_dff_B_yWfnQGqC1_0),.clk(gclk));
	jdff dff_B_GN5pjDSK5_0(.din(w_dff_B_yWfnQGqC1_0),.dout(w_dff_B_GN5pjDSK5_0),.clk(gclk));
	jdff dff_B_tb7gYmZ10_0(.din(w_dff_B_GN5pjDSK5_0),.dout(w_dff_B_tb7gYmZ10_0),.clk(gclk));
	jdff dff_B_oc0B1lNu8_0(.din(n1158),.dout(w_dff_B_oc0B1lNu8_0),.clk(gclk));
	jdff dff_B_QRfzaI208_2(.din(G152),.dout(w_dff_B_QRfzaI208_2),.clk(gclk));
	jdff dff_B_EkoNtpq80_2(.din(G155),.dout(w_dff_B_EkoNtpq80_2),.clk(gclk));
	jdff dff_B_BpTF5GQy4_2(.din(w_dff_B_EkoNtpq80_2),.dout(w_dff_B_BpTF5GQy4_2),.clk(gclk));
	jdff dff_B_aSaFLFPL9_1(.din(n1153),.dout(w_dff_B_aSaFLFPL9_1),.clk(gclk));
	jdff dff_B_Fv6no2Ey8_1(.din(w_dff_B_aSaFLFPL9_1),.dout(w_dff_B_Fv6no2Ey8_1),.clk(gclk));
	jdff dff_B_knRvT7tP7_1(.din(w_dff_B_Fv6no2Ey8_1),.dout(w_dff_B_knRvT7tP7_1),.clk(gclk));
	jdff dff_B_9TVfkL8R6_1(.din(n887),.dout(w_dff_B_9TVfkL8R6_1),.clk(gclk));
	jdff dff_B_F1guUStm2_1(.din(w_dff_B_9TVfkL8R6_1),.dout(w_dff_B_F1guUStm2_1),.clk(gclk));
	jdff dff_B_NKLB37uY2_1(.din(w_dff_B_F1guUStm2_1),.dout(w_dff_B_NKLB37uY2_1),.clk(gclk));
	jdff dff_B_MZgEDszm3_1(.din(w_dff_B_NKLB37uY2_1),.dout(w_dff_B_MZgEDszm3_1),.clk(gclk));
	jdff dff_B_3QS9wXdt8_1(.din(w_dff_B_MZgEDszm3_1),.dout(w_dff_B_3QS9wXdt8_1),.clk(gclk));
	jdff dff_B_qUJx8LBb8_0(.din(n893),.dout(w_dff_B_qUJx8LBb8_0),.clk(gclk));
	jdff dff_B_bsfaDhKk9_0(.din(w_dff_B_qUJx8LBb8_0),.dout(w_dff_B_bsfaDhKk9_0),.clk(gclk));
	jdff dff_B_xxqTxMre1_0(.din(w_dff_B_bsfaDhKk9_0),.dout(w_dff_B_xxqTxMre1_0),.clk(gclk));
	jdff dff_B_bTvv8oSU1_0(.din(w_dff_B_xxqTxMre1_0),.dout(w_dff_B_bTvv8oSU1_0),.clk(gclk));
	jdff dff_B_dLxIWmEe6_0(.din(w_dff_B_bTvv8oSU1_0),.dout(w_dff_B_dLxIWmEe6_0),.clk(gclk));
	jdff dff_B_Tgn2H91z5_1(.din(n489),.dout(w_dff_B_Tgn2H91z5_1),.clk(gclk));
	jdff dff_B_z1Eielot2_0(.din(n888),.dout(w_dff_B_z1Eielot2_0),.clk(gclk));
	jdff dff_B_vFwuNlNw2_1(.din(G127),.dout(w_dff_B_vFwuNlNw2_1),.clk(gclk));
	jdff dff_B_Hp7PbKvj2_1(.din(w_dff_B_vFwuNlNw2_1),.dout(w_dff_B_Hp7PbKvj2_1),.clk(gclk));
	jdff dff_B_rNs4GD8K8_1(.din(n843),.dout(w_dff_B_rNs4GD8K8_1),.clk(gclk));
	jdff dff_B_NLM2AQr62_1(.din(w_dff_B_rNs4GD8K8_1),.dout(w_dff_B_NLM2AQr62_1),.clk(gclk));
	jdff dff_B_trAlkVrw5_1(.din(w_dff_B_NLM2AQr62_1),.dout(w_dff_B_trAlkVrw5_1),.clk(gclk));
	jdff dff_B_zzFaTFQg8_1(.din(n844),.dout(w_dff_B_zzFaTFQg8_1),.clk(gclk));
	jdff dff_B_lghMQ7Yz0_1(.din(w_dff_B_zzFaTFQg8_1),.dout(w_dff_B_lghMQ7Yz0_1),.clk(gclk));
	jdff dff_B_7n3YPTJS0_1(.din(w_dff_B_lghMQ7Yz0_1),.dout(w_dff_B_7n3YPTJS0_1),.clk(gclk));
	jdff dff_A_30dIqxAf0_0(.dout(w_n847_0[0]),.din(w_dff_A_30dIqxAf0_0),.clk(gclk));
	jdff dff_A_qOxMpK4H6_0(.dout(w_dff_A_30dIqxAf0_0),.din(w_dff_A_qOxMpK4H6_0),.clk(gclk));
	jdff dff_A_ae4ddyxY3_0(.dout(w_dff_A_qOxMpK4H6_0),.din(w_dff_A_ae4ddyxY3_0),.clk(gclk));
	jdff dff_A_ww4RAWBC9_0(.dout(w_dff_A_ae4ddyxY3_0),.din(w_dff_A_ww4RAWBC9_0),.clk(gclk));
	jdff dff_B_SWNB9SoI5_1(.din(n393),.dout(w_dff_B_SWNB9SoI5_1),.clk(gclk));
	jdff dff_B_8gFBKhv31_1(.din(G119),.dout(w_dff_B_8gFBKhv31_1),.clk(gclk));
	jdff dff_B_qVeNaaDJ7_1(.din(w_dff_B_8gFBKhv31_1),.dout(w_dff_B_qVeNaaDJ7_1),.clk(gclk));
	jdff dff_B_026NcNg70_0(.din(n1168),.dout(w_dff_B_026NcNg70_0),.clk(gclk));
	jdff dff_B_pFSwHHtb2_0(.din(w_dff_B_026NcNg70_0),.dout(w_dff_B_pFSwHHtb2_0),.clk(gclk));
	jdff dff_B_jkWuy1ni8_0(.din(w_dff_B_pFSwHHtb2_0),.dout(w_dff_B_jkWuy1ni8_0),.clk(gclk));
	jdff dff_B_JXbAYvgO8_0(.din(w_dff_B_jkWuy1ni8_0),.dout(w_dff_B_JXbAYvgO8_0),.clk(gclk));
	jdff dff_B_jMxPL8SS5_0(.din(w_dff_B_JXbAYvgO8_0),.dout(w_dff_B_jMxPL8SS5_0),.clk(gclk));
	jdff dff_B_LCkv9DTj6_0(.din(w_dff_B_jMxPL8SS5_0),.dout(w_dff_B_LCkv9DTj6_0),.clk(gclk));
	jdff dff_B_qGXRgWgy9_0(.din(w_dff_B_LCkv9DTj6_0),.dout(w_dff_B_qGXRgWgy9_0),.clk(gclk));
	jdff dff_B_ZUjZvtYv0_0(.din(w_dff_B_qGXRgWgy9_0),.dout(w_dff_B_ZUjZvtYv0_0),.clk(gclk));
	jdff dff_B_tHPhL2Gm9_0(.din(w_dff_B_ZUjZvtYv0_0),.dout(w_dff_B_tHPhL2Gm9_0),.clk(gclk));
	jdff dff_B_2zxle7Eu4_0(.din(w_dff_B_tHPhL2Gm9_0),.dout(w_dff_B_2zxle7Eu4_0),.clk(gclk));
	jdff dff_B_coJcKL1t1_0(.din(w_dff_B_2zxle7Eu4_0),.dout(w_dff_B_coJcKL1t1_0),.clk(gclk));
	jdff dff_B_8jjA69mY4_0(.din(n1167),.dout(w_dff_B_8jjA69mY4_0),.clk(gclk));
	jdff dff_B_CUdKH9X76_2(.din(G146),.dout(w_dff_B_CUdKH9X76_2),.clk(gclk));
	jdff dff_B_r0QTEMSG2_2(.din(G149),.dout(w_dff_B_r0QTEMSG2_2),.clk(gclk));
	jdff dff_B_Vtj1ABIZ9_2(.din(w_dff_B_r0QTEMSG2_2),.dout(w_dff_B_Vtj1ABIZ9_2),.clk(gclk));
	jdff dff_B_wnl81Iyh3_1(.din(n1162),.dout(w_dff_B_wnl81Iyh3_1),.clk(gclk));
	jdff dff_B_9whXdIIs9_1(.din(n878),.dout(w_dff_B_9whXdIIs9_1),.clk(gclk));
	jdff dff_B_Q1rEGta80_1(.din(w_dff_B_9whXdIIs9_1),.dout(w_dff_B_Q1rEGta80_1),.clk(gclk));
	jdff dff_B_eOBOxAxZ8_1(.din(w_dff_B_Q1rEGta80_1),.dout(w_dff_B_eOBOxAxZ8_1),.clk(gclk));
	jdff dff_B_uM8Jl3zU7_1(.din(w_dff_B_eOBOxAxZ8_1),.dout(w_dff_B_uM8Jl3zU7_1),.clk(gclk));
	jdff dff_B_sSNvPANC4_1(.din(w_dff_B_uM8Jl3zU7_1),.dout(w_dff_B_sSNvPANC4_1),.clk(gclk));
	jdff dff_B_ODrs3Hv98_1(.din(w_dff_B_sSNvPANC4_1),.dout(w_dff_B_ODrs3Hv98_1),.clk(gclk));
	jdff dff_B_8hVuXK618_0(.din(n883),.dout(w_dff_B_8hVuXK618_0),.clk(gclk));
	jdff dff_B_i7CxdktL4_0(.din(w_dff_B_8hVuXK618_0),.dout(w_dff_B_i7CxdktL4_0),.clk(gclk));
	jdff dff_B_q9OM7uZS4_0(.din(w_dff_B_i7CxdktL4_0),.dout(w_dff_B_q9OM7uZS4_0),.clk(gclk));
	jdff dff_B_dqrFfrfa0_0(.din(w_dff_B_q9OM7uZS4_0),.dout(w_dff_B_dqrFfrfa0_0),.clk(gclk));
	jdff dff_B_5huyXDVK3_0(.din(w_dff_B_dqrFfrfa0_0),.dout(w_dff_B_5huyXDVK3_0),.clk(gclk));
	jdff dff_B_Gip1KnOr8_0(.din(w_dff_B_5huyXDVK3_0),.dout(w_dff_B_Gip1KnOr8_0),.clk(gclk));
	jdff dff_B_ns3mmr1l6_1(.din(n524),.dout(w_dff_B_ns3mmr1l6_1),.clk(gclk));
	jdff dff_A_AuhDZwQi4_2(.dout(w_G4092_7[2]),.din(w_dff_A_AuhDZwQi4_2),.clk(gclk));
	jdff dff_A_HB1k4VTa7_2(.dout(w_dff_A_AuhDZwQi4_2),.din(w_dff_A_HB1k4VTa7_2),.clk(gclk));
	jdff dff_A_sVMre9Ik6_2(.dout(w_dff_A_HB1k4VTa7_2),.din(w_dff_A_sVMre9Ik6_2),.clk(gclk));
	jdff dff_A_MV8w9BWA8_0(.dout(w_n880_0[0]),.din(w_dff_A_MV8w9BWA8_0),.clk(gclk));
	jdff dff_A_qQK4ptO99_0(.dout(w_dff_A_MV8w9BWA8_0),.din(w_dff_A_qQK4ptO99_0),.clk(gclk));
	jdff dff_A_9GCQO9zD4_0(.dout(w_dff_A_qQK4ptO99_0),.din(w_dff_A_9GCQO9zD4_0),.clk(gclk));
	jdff dff_A_9gC8U8aS1_1(.dout(w_G4091_3[1]),.din(w_dff_A_9gC8U8aS1_1),.clk(gclk));
	jdff dff_A_clEifxhA9_2(.dout(w_G4091_3[2]),.din(w_dff_A_clEifxhA9_2),.clk(gclk));
	jdff dff_A_VBoCBJqN8_2(.dout(w_dff_A_clEifxhA9_2),.din(w_dff_A_VBoCBJqN8_2),.clk(gclk));
	jdff dff_B_lXrQxOTa6_1(.din(G128),.dout(w_dff_B_lXrQxOTa6_1),.clk(gclk));
	jdff dff_B_bMPd2nWQ2_1(.din(w_dff_B_lXrQxOTa6_1),.dout(w_dff_B_bMPd2nWQ2_1),.clk(gclk));
	jdff dff_A_CJHvcAcc3_0(.dout(w_n1008_3[0]),.din(w_dff_A_CJHvcAcc3_0),.clk(gclk));
	jdff dff_A_BaOSPFsm5_0(.dout(w_dff_A_CJHvcAcc3_0),.din(w_dff_A_BaOSPFsm5_0),.clk(gclk));
	jdff dff_A_rDg5QNjv5_1(.dout(w_n1008_3[1]),.din(w_dff_A_rDg5QNjv5_1),.clk(gclk));
	jdff dff_B_SyrpvCGw4_1(.din(n834),.dout(w_dff_B_SyrpvCGw4_1),.clk(gclk));
	jdff dff_B_cF1kL6Ir0_1(.din(w_dff_B_SyrpvCGw4_1),.dout(w_dff_B_cF1kL6Ir0_1),.clk(gclk));
	jdff dff_B_n5R4Zt7E6_1(.din(w_dff_B_cF1kL6Ir0_1),.dout(w_dff_B_n5R4Zt7E6_1),.clk(gclk));
	jdff dff_B_6QAueIRe5_1(.din(w_dff_B_n5R4Zt7E6_1),.dout(w_dff_B_6QAueIRe5_1),.clk(gclk));
	jdff dff_B_6AfSqez20_1(.din(w_dff_B_6QAueIRe5_1),.dout(w_dff_B_6AfSqez20_1),.clk(gclk));
	jdff dff_B_ETrn17uu3_1(.din(w_dff_B_6AfSqez20_1),.dout(w_dff_B_ETrn17uu3_1),.clk(gclk));
	jdff dff_B_aHYp6zQn1_0(.din(n839),.dout(w_dff_B_aHYp6zQn1_0),.clk(gclk));
	jdff dff_B_7XkRhDja7_0(.din(w_dff_B_aHYp6zQn1_0),.dout(w_dff_B_7XkRhDja7_0),.clk(gclk));
	jdff dff_B_p9Yvvedh9_0(.din(w_dff_B_7XkRhDja7_0),.dout(w_dff_B_p9Yvvedh9_0),.clk(gclk));
	jdff dff_B_McGf1tEs0_0(.din(w_dff_B_p9Yvvedh9_0),.dout(w_dff_B_McGf1tEs0_0),.clk(gclk));
	jdff dff_B_6LzYTQeG1_0(.din(w_dff_B_McGf1tEs0_0),.dout(w_dff_B_6LzYTQeG1_0),.clk(gclk));
	jdff dff_B_6H8o4d9y1_0(.din(w_dff_B_6LzYTQeG1_0),.dout(w_dff_B_6H8o4d9y1_0),.clk(gclk));
	jdff dff_B_de19BWZc6_1(.din(n360),.dout(w_dff_B_de19BWZc6_1),.clk(gclk));
	jdff dff_A_WqWAB9at4_0(.dout(w_n836_0[0]),.din(w_dff_A_WqWAB9at4_0),.clk(gclk));
	jdff dff_A_DwUkGJs80_0(.dout(w_dff_A_WqWAB9at4_0),.din(w_dff_A_DwUkGJs80_0),.clk(gclk));
	jdff dff_A_L8dLDJ6w5_0(.dout(w_dff_A_DwUkGJs80_0),.din(w_dff_A_L8dLDJ6w5_0),.clk(gclk));
	jdff dff_A_5bRvF0Nh4_0(.dout(w_dff_A_L8dLDJ6w5_0),.din(w_dff_A_5bRvF0Nh4_0),.clk(gclk));
	jdff dff_A_FIlawX3a4_1(.dout(w_n753_0[1]),.din(w_dff_A_FIlawX3a4_1),.clk(gclk));
	jdff dff_A_aQ50xBuz5_1(.dout(w_dff_A_FIlawX3a4_1),.din(w_dff_A_aQ50xBuz5_1),.clk(gclk));
	jdff dff_A_3bDdvGbk4_2(.dout(w_n753_0[2]),.din(w_dff_A_3bDdvGbk4_2),.clk(gclk));
	jdff dff_A_2WmamI4n2_2(.dout(w_dff_A_3bDdvGbk4_2),.din(w_dff_A_2WmamI4n2_2),.clk(gclk));
	jdff dff_A_beQmwRy67_2(.dout(w_dff_A_2WmamI4n2_2),.din(w_dff_A_beQmwRy67_2),.clk(gclk));
	jdff dff_A_ks8FVTFN3_2(.dout(w_dff_A_beQmwRy67_2),.din(w_dff_A_ks8FVTFN3_2),.clk(gclk));
	jdff dff_A_4WBJbeab2_2(.dout(w_dff_A_ks8FVTFN3_2),.din(w_dff_A_4WBJbeab2_2),.clk(gclk));
	jdff dff_B_t1FXFAaZ7_3(.din(n753),.dout(w_dff_B_t1FXFAaZ7_3),.clk(gclk));
	jdff dff_A_DHNOFN4p6_0(.dout(w_G4091_4[0]),.din(w_dff_A_DHNOFN4p6_0),.clk(gclk));
	jdff dff_A_WGV5FVai3_0(.dout(w_dff_A_DHNOFN4p6_0),.din(w_dff_A_WGV5FVai3_0),.clk(gclk));
	jdff dff_A_AdnlTC4Y5_0(.dout(w_dff_A_WGV5FVai3_0),.din(w_dff_A_AdnlTC4Y5_0),.clk(gclk));
	jdff dff_A_smjPFL1o7_0(.dout(w_dff_A_AdnlTC4Y5_0),.din(w_dff_A_smjPFL1o7_0),.clk(gclk));
	jdff dff_A_EWBqzcHE4_2(.dout(w_G4091_4[2]),.din(w_dff_A_EWBqzcHE4_2),.clk(gclk));
	jdff dff_A_Jyys0oDK4_2(.dout(w_dff_A_EWBqzcHE4_2),.din(w_dff_A_Jyys0oDK4_2),.clk(gclk));
	jdff dff_A_rbirpuik2_2(.dout(w_dff_A_Jyys0oDK4_2),.din(w_dff_A_rbirpuik2_2),.clk(gclk));
	jdff dff_B_bLfx55vc8_1(.din(G130),.dout(w_dff_B_bLfx55vc8_1),.clk(gclk));
	jdff dff_B_9OEG3cWT9_1(.din(w_dff_B_bLfx55vc8_1),.dout(w_dff_B_9OEG3cWT9_1),.clk(gclk));
	jdff dff_B_tO0mzwg96_1(.din(n1173),.dout(w_dff_B_tO0mzwg96_1),.clk(gclk));
	jdff dff_B_lhRGlw9K9_1(.din(w_dff_B_tO0mzwg96_1),.dout(w_dff_B_lhRGlw9K9_1),.clk(gclk));
	jdff dff_B_FQQWkwii8_1(.din(w_dff_B_lhRGlw9K9_1),.dout(w_dff_B_FQQWkwii8_1),.clk(gclk));
	jdff dff_B_wn5iN9zw9_1(.din(w_dff_B_FQQWkwii8_1),.dout(w_dff_B_wn5iN9zw9_1),.clk(gclk));
	jdff dff_B_SjU1yt2V7_1(.din(w_dff_B_wn5iN9zw9_1),.dout(w_dff_B_SjU1yt2V7_1),.clk(gclk));
	jdff dff_B_unZKnTdD0_1(.din(w_dff_B_SjU1yt2V7_1),.dout(w_dff_B_unZKnTdD0_1),.clk(gclk));
	jdff dff_B_70wxUfHc4_1(.din(w_dff_B_unZKnTdD0_1),.dout(w_dff_B_70wxUfHc4_1),.clk(gclk));
	jdff dff_B_B7UMTwev4_1(.din(w_dff_B_70wxUfHc4_1),.dout(w_dff_B_B7UMTwev4_1),.clk(gclk));
	jdff dff_B_FlQNaKcG7_1(.din(w_dff_B_B7UMTwev4_1),.dout(w_dff_B_FlQNaKcG7_1),.clk(gclk));
	jdff dff_B_eQteUKjZ2_1(.din(w_dff_B_FlQNaKcG7_1),.dout(w_dff_B_eQteUKjZ2_1),.clk(gclk));
	jdff dff_B_XLSHq1Th9_1(.din(w_dff_B_eQteUKjZ2_1),.dout(w_dff_B_XLSHq1Th9_1),.clk(gclk));
	jdff dff_B_2u0ShZUG1_1(.din(w_dff_B_XLSHq1Th9_1),.dout(w_dff_B_2u0ShZUG1_1),.clk(gclk));
	jdff dff_B_NGnx5LnA9_1(.din(n1182),.dout(w_dff_B_NGnx5LnA9_1),.clk(gclk));
	jdff dff_B_198XHMzy8_1(.din(w_dff_B_NGnx5LnA9_1),.dout(w_dff_B_198XHMzy8_1),.clk(gclk));
	jdff dff_B_PSrErrhy7_1(.din(w_dff_B_198XHMzy8_1),.dout(w_dff_B_PSrErrhy7_1),.clk(gclk));
	jdff dff_B_qynal3SP1_1(.din(w_dff_B_PSrErrhy7_1),.dout(w_dff_B_qynal3SP1_1),.clk(gclk));
	jdff dff_B_QekT2fM28_1(.din(w_dff_B_qynal3SP1_1),.dout(w_dff_B_QekT2fM28_1),.clk(gclk));
	jdff dff_B_Xt9Y9EYs6_1(.din(w_dff_B_QekT2fM28_1),.dout(w_dff_B_Xt9Y9EYs6_1),.clk(gclk));
	jdff dff_B_QyHALjbl8_0(.din(n1185),.dout(w_dff_B_QyHALjbl8_0),.clk(gclk));
	jdff dff_B_8p7F8Wpz3_0(.din(w_dff_B_QyHALjbl8_0),.dout(w_dff_B_8p7F8Wpz3_0),.clk(gclk));
	jdff dff_B_D4sCE0H09_0(.din(w_dff_B_8p7F8Wpz3_0),.dout(w_dff_B_D4sCE0H09_0),.clk(gclk));
	jdff dff_B_KmYStiCn2_0(.din(w_dff_B_D4sCE0H09_0),.dout(w_dff_B_KmYStiCn2_0),.clk(gclk));
	jdff dff_B_vhdNbXMJ9_0(.din(w_dff_B_KmYStiCn2_0),.dout(w_dff_B_vhdNbXMJ9_0),.clk(gclk));
	jdff dff_B_BqG7FfWw6_0(.din(w_dff_B_vhdNbXMJ9_0),.dout(w_dff_B_BqG7FfWw6_0),.clk(gclk));
	jdff dff_B_owT8PVMb3_0(.din(w_dff_B_BqG7FfWw6_0),.dout(w_dff_B_owT8PVMb3_0),.clk(gclk));
	jdff dff_B_VTJlbBN22_0(.din(w_dff_B_owT8PVMb3_0),.dout(w_dff_B_VTJlbBN22_0),.clk(gclk));
	jdff dff_B_Vl5L1zmB2_0(.din(w_dff_B_VTJlbBN22_0),.dout(w_dff_B_Vl5L1zmB2_0),.clk(gclk));
	jdff dff_B_7lHRc8zN2_0(.din(w_dff_B_Vl5L1zmB2_0),.dout(w_dff_B_7lHRc8zN2_0),.clk(gclk));
	jdff dff_B_KnwnaKGM1_0(.din(w_dff_B_7lHRc8zN2_0),.dout(w_dff_B_KnwnaKGM1_0),.clk(gclk));
	jdff dff_B_ITFQcYXI8_1(.din(n1175),.dout(w_dff_B_ITFQcYXI8_1),.clk(gclk));
	jdff dff_B_0qpq5DAt7_1(.din(w_dff_B_ITFQcYXI8_1),.dout(w_dff_B_0qpq5DAt7_1),.clk(gclk));
	jdff dff_B_KgvbjEim3_1(.din(w_dff_B_0qpq5DAt7_1),.dout(w_dff_B_KgvbjEim3_1),.clk(gclk));
	jdff dff_B_fPVcmVYO6_1(.din(n1176),.dout(w_dff_B_fPVcmVYO6_1),.clk(gclk));
	jdff dff_B_ajBqM8tc6_1(.din(w_dff_B_fPVcmVYO6_1),.dout(w_dff_B_ajBqM8tc6_1),.clk(gclk));
	jdff dff_B_CQpxvma20_1(.din(w_dff_B_ajBqM8tc6_1),.dout(w_dff_B_CQpxvma20_1),.clk(gclk));
	jdff dff_B_P0bI9bgD6_1(.din(w_dff_B_CQpxvma20_1),.dout(w_dff_B_P0bI9bgD6_1),.clk(gclk));
	jdff dff_A_szaHesc36_0(.dout(w_n1177_0[0]),.din(w_dff_A_szaHesc36_0),.clk(gclk));
	jdff dff_A_vXyBZDLX0_0(.dout(w_dff_A_szaHesc36_0),.din(w_dff_A_vXyBZDLX0_0),.clk(gclk));
	jdff dff_A_WfZzG6FB3_0(.dout(w_dff_A_vXyBZDLX0_0),.din(w_dff_A_WfZzG6FB3_0),.clk(gclk));
	jdff dff_A_bln2jIrX8_0(.dout(w_dff_A_WfZzG6FB3_0),.din(w_dff_A_bln2jIrX8_0),.clk(gclk));
	jdff dff_A_SVYpcLbw9_0(.dout(w_dff_A_bln2jIrX8_0),.din(w_dff_A_SVYpcLbw9_0),.clk(gclk));
	jdff dff_A_C1IDkzsS0_0(.dout(w_dff_A_SVYpcLbw9_0),.din(w_dff_A_C1IDkzsS0_0),.clk(gclk));
	jdff dff_A_i4bemp5d7_0(.dout(w_dff_A_C1IDkzsS0_0),.din(w_dff_A_i4bemp5d7_0),.clk(gclk));
	jdff dff_B_o9gmxaQ76_2(.din(n1177),.dout(w_dff_B_o9gmxaQ76_2),.clk(gclk));
	jdff dff_B_UCILfZAn5_2(.din(w_dff_B_o9gmxaQ76_2),.dout(w_dff_B_UCILfZAn5_2),.clk(gclk));
	jdff dff_B_RSIx4bsn9_2(.din(w_dff_B_UCILfZAn5_2),.dout(w_dff_B_RSIx4bsn9_2),.clk(gclk));
	jdff dff_B_cMRgaMlm1_2(.din(w_dff_B_RSIx4bsn9_2),.dout(w_dff_B_cMRgaMlm1_2),.clk(gclk));
	jdff dff_A_pZ8QkzW89_1(.dout(w_n428_1[1]),.din(w_dff_A_pZ8QkzW89_1),.clk(gclk));
	jdff dff_A_UrsF4Apy8_2(.dout(w_G3724_0[2]),.din(w_dff_A_UrsF4Apy8_2),.clk(gclk));
	jdff dff_A_c54t0iqu8_2(.dout(w_dff_A_UrsF4Apy8_2),.din(w_dff_A_c54t0iqu8_2),.clk(gclk));
	jdff dff_A_wwcE1kRT2_2(.dout(w_dff_A_c54t0iqu8_2),.din(w_dff_A_wwcE1kRT2_2),.clk(gclk));
	jdff dff_A_3iQpeY224_0(.dout(w_n1179_0[0]),.din(w_dff_A_3iQpeY224_0),.clk(gclk));
	jdff dff_A_o5mE3gb71_0(.dout(w_dff_A_3iQpeY224_0),.din(w_dff_A_o5mE3gb71_0),.clk(gclk));
	jdff dff_A_VN0ZYhaT8_0(.dout(w_dff_A_o5mE3gb71_0),.din(w_dff_A_VN0ZYhaT8_0),.clk(gclk));
	jdff dff_A_quFaGz0f9_0(.dout(w_dff_A_VN0ZYhaT8_0),.din(w_dff_A_quFaGz0f9_0),.clk(gclk));
	jdff dff_A_lDlSrtFN3_0(.dout(w_dff_A_quFaGz0f9_0),.din(w_dff_A_lDlSrtFN3_0),.clk(gclk));
	jdff dff_A_Gplb7tj13_0(.dout(w_dff_A_lDlSrtFN3_0),.din(w_dff_A_Gplb7tj13_0),.clk(gclk));
	jdff dff_A_euOf8vAs0_0(.dout(w_dff_A_Gplb7tj13_0),.din(w_dff_A_euOf8vAs0_0),.clk(gclk));
	jdff dff_B_EdChOtUI6_1(.din(G132),.dout(w_dff_B_EdChOtUI6_1),.clk(gclk));
	jdff dff_B_IgrB5vSH2_1(.din(w_dff_B_EdChOtUI6_1),.dout(w_dff_B_IgrB5vSH2_1),.clk(gclk));
	jdff dff_B_K6VgBYY54_1(.din(w_dff_B_IgrB5vSH2_1),.dout(w_dff_B_K6VgBYY54_1),.clk(gclk));
	jdff dff_B_oRispRRq4_1(.din(n1223),.dout(w_dff_B_oRispRRq4_1),.clk(gclk));
	jdff dff_B_KZEWDumJ5_0(.din(n1227),.dout(w_dff_B_KZEWDumJ5_0),.clk(gclk));
	jdff dff_B_3nXIKtGi0_0(.din(w_dff_B_KZEWDumJ5_0),.dout(w_dff_B_3nXIKtGi0_0),.clk(gclk));
	jdff dff_B_LDROBFzc7_0(.din(w_dff_B_3nXIKtGi0_0),.dout(w_dff_B_LDROBFzc7_0),.clk(gclk));
	jdff dff_B_kmLJ1tZm4_0(.din(w_dff_B_LDROBFzc7_0),.dout(w_dff_B_kmLJ1tZm4_0),.clk(gclk));
	jdff dff_B_CqnFOVbl3_0(.din(n1226),.dout(w_dff_B_CqnFOVbl3_0),.clk(gclk));
	jdff dff_A_voFT6FAY7_0(.dout(w_G559_0[0]),.din(w_dff_A_voFT6FAY7_0),.clk(gclk));
	jdff dff_A_5dlESbO32_0(.dout(w_dff_A_voFT6FAY7_0),.din(w_dff_A_5dlESbO32_0),.clk(gclk));
	jdff dff_B_8m802Xw05_0(.din(n668),.dout(w_dff_B_8m802Xw05_0),.clk(gclk));
	jdff dff_B_HrWB5H7K4_1(.din(n663),.dout(w_dff_B_HrWB5H7K4_1),.clk(gclk));
	jdff dff_B_ieA4H7A44_1(.din(n916),.dout(w_dff_B_ieA4H7A44_1),.clk(gclk));
	jdff dff_B_oLh5Lp4R4_1(.din(w_dff_B_ieA4H7A44_1),.dout(w_dff_B_oLh5Lp4R4_1),.clk(gclk));
	jdff dff_B_uBK8rf9p3_1(.din(n917),.dout(w_dff_B_uBK8rf9p3_1),.clk(gclk));
	jdff dff_B_6hPxrTld8_1(.din(w_dff_B_uBK8rf9p3_1),.dout(w_dff_B_6hPxrTld8_1),.clk(gclk));
	jdff dff_B_ZQaKcf964_0(.din(n915),.dout(w_dff_B_ZQaKcf964_0),.clk(gclk));
	jdff dff_B_ubAaVd4l6_1(.din(n913),.dout(w_dff_B_ubAaVd4l6_1),.clk(gclk));
	jdff dff_B_jCDCYhlj0_0(.din(G372),.dout(w_dff_B_jCDCYhlj0_0),.clk(gclk));
	jdff dff_B_5GvTtmRH5_0(.din(n911),.dout(w_dff_B_5GvTtmRH5_0),.clk(gclk));
	jdff dff_B_i8kUr1e56_1(.din(n909),.dout(w_dff_B_i8kUr1e56_1),.clk(gclk));
	jdff dff_B_lprhXOTy9_1(.din(w_dff_B_i8kUr1e56_1),.dout(w_dff_B_lprhXOTy9_1),.clk(gclk));
	jdff dff_B_nmbHJMig4_1(.din(n907),.dout(w_dff_B_nmbHJMig4_1),.clk(gclk));
	jdff dff_B_YidhlQNS8_0(.din(n1222),.dout(w_dff_B_YidhlQNS8_0),.clk(gclk));
	jdff dff_B_AjBRgu6e9_0(.din(w_dff_B_YidhlQNS8_0),.dout(w_dff_B_AjBRgu6e9_0),.clk(gclk));
	jdff dff_B_yQZ9oo2Z6_0(.din(w_dff_B_AjBRgu6e9_0),.dout(w_dff_B_yQZ9oo2Z6_0),.clk(gclk));
	jdff dff_B_UkrEuE9s7_0(.din(n678),.dout(w_dff_B_UkrEuE9s7_0),.clk(gclk));
	jdff dff_B_VDU12DIm5_1(.din(n672),.dout(w_dff_B_VDU12DIm5_1),.clk(gclk));
	jdff dff_A_cIv5IQkG3_0(.dout(w_G245_0[0]),.din(w_dff_A_cIv5IQkG3_0),.clk(gclk));
	jdff dff_A_xRo5UZdV2_0(.dout(w_dff_A_cIv5IQkG3_0),.din(w_dff_A_xRo5UZdV2_0),.clk(gclk));
	jdff dff_A_BsGQ8ETt0_0(.dout(w_dff_A_xRo5UZdV2_0),.din(w_dff_A_BsGQ8ETt0_0),.clk(gclk));
	jdff dff_A_G9Pwthw85_0(.dout(w_dff_A_BsGQ8ETt0_0),.din(w_dff_A_G9Pwthw85_0),.clk(gclk));
	jdff dff_B_M65zM5Hf2_1(.din(n926),.dout(w_dff_B_M65zM5Hf2_1),.clk(gclk));
	jdff dff_B_zeRRCORY7_1(.din(n930),.dout(w_dff_B_zeRRCORY7_1),.clk(gclk));
	jdff dff_B_pZDJJ7u89_1(.din(w_dff_B_zeRRCORY7_1),.dout(w_dff_B_pZDJJ7u89_1),.clk(gclk));
	jdff dff_B_SayaEkvV4_1(.din(w_dff_B_pZDJJ7u89_1),.dout(w_dff_B_SayaEkvV4_1),.clk(gclk));
	jdff dff_B_gagvMuUz4_1(.din(n927),.dout(w_dff_B_gagvMuUz4_1),.clk(gclk));
	jdff dff_B_miCOhRWA2_1(.din(G292),.dout(w_dff_B_miCOhRWA2_1),.clk(gclk));
	jdff dff_B_8zVrpvmF9_1(.din(n1263),.dout(w_dff_B_8zVrpvmF9_1),.clk(gclk));
	jdff dff_B_7Aumt0np9_1(.din(w_dff_B_8zVrpvmF9_1),.dout(w_dff_B_7Aumt0np9_1),.clk(gclk));
	jdff dff_B_R3GMazw41_1(.din(w_dff_B_7Aumt0np9_1),.dout(w_dff_B_R3GMazw41_1),.clk(gclk));
	jdff dff_B_CcFBvzJs4_1(.din(w_dff_B_R3GMazw41_1),.dout(w_dff_B_CcFBvzJs4_1),.clk(gclk));
	jdff dff_B_6rxe9iZv5_1(.din(w_dff_B_CcFBvzJs4_1),.dout(w_dff_B_6rxe9iZv5_1),.clk(gclk));
	jdff dff_B_6ai4waMO7_1(.din(w_dff_B_6rxe9iZv5_1),.dout(w_dff_B_6ai4waMO7_1),.clk(gclk));
	jdff dff_B_jyX6kh7H4_1(.din(w_dff_B_6ai4waMO7_1),.dout(w_dff_B_jyX6kh7H4_1),.clk(gclk));
	jdff dff_B_HpivnRXk6_1(.din(w_dff_B_jyX6kh7H4_1),.dout(w_dff_B_HpivnRXk6_1),.clk(gclk));
	jdff dff_B_kjUlIwkl0_1(.din(w_dff_B_HpivnRXk6_1),.dout(w_dff_B_kjUlIwkl0_1),.clk(gclk));
	jdff dff_B_1r5N1f4X6_1(.din(w_dff_B_kjUlIwkl0_1),.dout(w_dff_B_1r5N1f4X6_1),.clk(gclk));
	jdff dff_B_7Gg8tduh0_1(.din(w_dff_B_1r5N1f4X6_1),.dout(w_dff_B_7Gg8tduh0_1),.clk(gclk));
	jdff dff_B_y4GRpozF4_1(.din(w_dff_B_7Gg8tduh0_1),.dout(w_dff_B_y4GRpozF4_1),.clk(gclk));
	jdff dff_B_UpTPaB8V4_1(.din(w_dff_B_y4GRpozF4_1),.dout(w_dff_B_UpTPaB8V4_1),.clk(gclk));
	jdff dff_B_l5liVw6T3_0(.din(n1266),.dout(w_dff_B_l5liVw6T3_0),.clk(gclk));
	jdff dff_B_x1Sxh1Kz0_1(.din(n1260),.dout(w_dff_B_x1Sxh1Kz0_1),.clk(gclk));
	jdff dff_B_oIzlAM068_1(.din(w_dff_B_x1Sxh1Kz0_1),.dout(w_dff_B_oIzlAM068_1),.clk(gclk));
	jdff dff_A_4RjYFG4K9_2(.dout(w_n852_6[2]),.din(w_dff_A_4RjYFG4K9_2),.clk(gclk));
	jdff dff_A_ZLMebdVg6_2(.dout(w_dff_A_4RjYFG4K9_2),.din(w_dff_A_ZLMebdVg6_2),.clk(gclk));
	jdff dff_A_rCyVFMDg6_2(.dout(w_dff_A_ZLMebdVg6_2),.din(w_dff_A_rCyVFMDg6_2),.clk(gclk));
	jdff dff_A_wHMLXklS3_2(.dout(w_dff_A_rCyVFMDg6_2),.din(w_dff_A_wHMLXklS3_2),.clk(gclk));
	jdff dff_A_DsOyQXxt6_2(.dout(w_dff_A_wHMLXklS3_2),.din(w_dff_A_DsOyQXxt6_2),.clk(gclk));
	jdff dff_A_ob3Uspce6_2(.dout(w_dff_A_DsOyQXxt6_2),.din(w_dff_A_ob3Uspce6_2),.clk(gclk));
	jdff dff_A_X1HmajJw6_2(.dout(w_dff_A_ob3Uspce6_2),.din(w_dff_A_X1HmajJw6_2),.clk(gclk));
	jdff dff_A_NvnRKjZL9_2(.dout(w_dff_A_X1HmajJw6_2),.din(w_dff_A_NvnRKjZL9_2),.clk(gclk));
	jdff dff_A_9x3Yo8EN9_2(.dout(w_dff_A_NvnRKjZL9_2),.din(w_dff_A_9x3Yo8EN9_2),.clk(gclk));
	jdff dff_A_8JGtiVNQ6_2(.dout(w_G4089_6[2]),.din(w_dff_A_8JGtiVNQ6_2),.clk(gclk));
	jdff dff_A_LMOioVDJ3_2(.dout(w_dff_A_8JGtiVNQ6_2),.din(w_dff_A_LMOioVDJ3_2),.clk(gclk));
	jdff dff_A_eJYbyVf70_2(.dout(w_dff_A_LMOioVDJ3_2),.din(w_dff_A_eJYbyVf70_2),.clk(gclk));
	jdff dff_A_GEgtIHgQ6_2(.dout(w_dff_A_eJYbyVf70_2),.din(w_dff_A_GEgtIHgQ6_2),.clk(gclk));
	jdff dff_A_CAXsjpkX6_2(.dout(w_dff_A_GEgtIHgQ6_2),.din(w_dff_A_CAXsjpkX6_2),.clk(gclk));
	jdff dff_A_PNDRObHB4_2(.dout(w_dff_A_CAXsjpkX6_2),.din(w_dff_A_PNDRObHB4_2),.clk(gclk));
	jdff dff_A_Z519ggSy1_2(.dout(w_dff_A_PNDRObHB4_2),.din(w_dff_A_Z519ggSy1_2),.clk(gclk));
	jdff dff_A_d22uQCar0_2(.dout(w_dff_A_Z519ggSy1_2),.din(w_dff_A_d22uQCar0_2),.clk(gclk));
	jdff dff_A_JDItCrtt2_2(.dout(w_dff_A_d22uQCar0_2),.din(w_dff_A_JDItCrtt2_2),.clk(gclk));
	jdff dff_A_YrEGUGTu5_2(.dout(w_dff_A_JDItCrtt2_2),.din(w_dff_A_YrEGUGTu5_2),.clk(gclk));
	jdff dff_B_HSLOQpXc2_0(.din(n1276),.dout(w_dff_B_HSLOQpXc2_0),.clk(gclk));
	jdff dff_B_lgbymOOJ9_0(.din(w_dff_B_HSLOQpXc2_0),.dout(w_dff_B_lgbymOOJ9_0),.clk(gclk));
	jdff dff_B_N9vB34J35_0(.din(w_dff_B_lgbymOOJ9_0),.dout(w_dff_B_N9vB34J35_0),.clk(gclk));
	jdff dff_B_XSoYDXjI0_0(.din(w_dff_B_N9vB34J35_0),.dout(w_dff_B_XSoYDXjI0_0),.clk(gclk));
	jdff dff_B_K9jChpCQ0_0(.din(w_dff_B_XSoYDXjI0_0),.dout(w_dff_B_K9jChpCQ0_0),.clk(gclk));
	jdff dff_B_sjwgHYEH6_0(.din(w_dff_B_K9jChpCQ0_0),.dout(w_dff_B_sjwgHYEH6_0),.clk(gclk));
	jdff dff_B_pUomxi3t2_0(.din(w_dff_B_sjwgHYEH6_0),.dout(w_dff_B_pUomxi3t2_0),.clk(gclk));
	jdff dff_B_3fI1vQaf1_0(.din(w_dff_B_pUomxi3t2_0),.dout(w_dff_B_3fI1vQaf1_0),.clk(gclk));
	jdff dff_B_AL122XYB9_0(.din(w_dff_B_3fI1vQaf1_0),.dout(w_dff_B_AL122XYB9_0),.clk(gclk));
	jdff dff_B_LWtPXt185_0(.din(w_dff_B_AL122XYB9_0),.dout(w_dff_B_LWtPXt185_0),.clk(gclk));
	jdff dff_B_GLeeVZ5K7_0(.din(w_dff_B_LWtPXt185_0),.dout(w_dff_B_GLeeVZ5K7_0),.clk(gclk));
	jdff dff_B_QZjZ94RC1_0(.din(w_dff_B_GLeeVZ5K7_0),.dout(w_dff_B_QZjZ94RC1_0),.clk(gclk));
	jdff dff_B_ciHm6jhR3_0(.din(w_dff_B_QZjZ94RC1_0),.dout(w_dff_B_ciHm6jhR3_0),.clk(gclk));
	jdff dff_B_8CktlJcR5_0(.din(w_dff_B_ciHm6jhR3_0),.dout(w_dff_B_8CktlJcR5_0),.clk(gclk));
	jdff dff_B_cP2vFUK47_0(.din(w_dff_B_8CktlJcR5_0),.dout(w_dff_B_cP2vFUK47_0),.clk(gclk));
	jdff dff_B_Ys6cIc8n8_2(.din(G106),.dout(w_dff_B_Ys6cIc8n8_2),.clk(gclk));
	jdff dff_B_X6mec9Ar6_1(.din(n1269),.dout(w_dff_B_X6mec9Ar6_1),.clk(gclk));
	jdff dff_B_tII93kEQ5_1(.din(w_dff_B_X6mec9Ar6_1),.dout(w_dff_B_tII93kEQ5_1),.clk(gclk));
	jdff dff_B_beRkpLEE2_1(.din(w_dff_B_tII93kEQ5_1),.dout(w_dff_B_beRkpLEE2_1),.clk(gclk));
	jdff dff_A_EIhygtvp0_0(.dout(w_n797_6[0]),.din(w_dff_A_EIhygtvp0_0),.clk(gclk));
	jdff dff_A_0xH5TIIg0_0(.dout(w_dff_A_EIhygtvp0_0),.din(w_dff_A_0xH5TIIg0_0),.clk(gclk));
	jdff dff_A_mfQpytnV1_0(.dout(w_dff_A_0xH5TIIg0_0),.din(w_dff_A_mfQpytnV1_0),.clk(gclk));
	jdff dff_A_WKC49Meu0_0(.dout(w_dff_A_mfQpytnV1_0),.din(w_dff_A_WKC49Meu0_0),.clk(gclk));
	jdff dff_A_1gxq7JWy7_0(.dout(w_dff_A_WKC49Meu0_0),.din(w_dff_A_1gxq7JWy7_0),.clk(gclk));
	jdff dff_A_bevwvuwM9_0(.dout(w_dff_A_1gxq7JWy7_0),.din(w_dff_A_bevwvuwM9_0),.clk(gclk));
	jdff dff_A_ZxnVxvec0_0(.dout(w_dff_A_bevwvuwM9_0),.din(w_dff_A_ZxnVxvec0_0),.clk(gclk));
	jdff dff_A_fPSPLAGd1_0(.dout(w_dff_A_ZxnVxvec0_0),.din(w_dff_A_fPSPLAGd1_0),.clk(gclk));
	jdff dff_A_d0MrzTYe8_0(.dout(w_dff_A_fPSPLAGd1_0),.din(w_dff_A_d0MrzTYe8_0),.clk(gclk));
	jdff dff_A_ShtoPeI53_0(.dout(w_dff_A_d0MrzTYe8_0),.din(w_dff_A_ShtoPeI53_0),.clk(gclk));
	jdff dff_A_wRUR3CdM8_0(.dout(w_dff_A_ShtoPeI53_0),.din(w_dff_A_wRUR3CdM8_0),.clk(gclk));
	jdff dff_A_Z5xKLcse1_0(.dout(w_dff_A_wRUR3CdM8_0),.din(w_dff_A_Z5xKLcse1_0),.clk(gclk));
	jdff dff_A_7paWf7me8_0(.dout(w_dff_A_Z5xKLcse1_0),.din(w_dff_A_7paWf7me8_0),.clk(gclk));
	jdff dff_A_i7vIy5nd8_0(.dout(w_dff_A_7paWf7me8_0),.din(w_dff_A_i7vIy5nd8_0),.clk(gclk));
	jdff dff_A_l07kGdf07_2(.dout(w_n797_6[2]),.din(w_dff_A_l07kGdf07_2),.clk(gclk));
	jdff dff_A_QALrA6Ug2_2(.dout(w_dff_A_l07kGdf07_2),.din(w_dff_A_QALrA6Ug2_2),.clk(gclk));
	jdff dff_A_3ov9t8sz4_2(.dout(w_dff_A_QALrA6Ug2_2),.din(w_dff_A_3ov9t8sz4_2),.clk(gclk));
	jdff dff_A_Cr28jNBd5_2(.dout(w_dff_A_3ov9t8sz4_2),.din(w_dff_A_Cr28jNBd5_2),.clk(gclk));
	jdff dff_A_tShaQ5nr3_2(.dout(w_dff_A_Cr28jNBd5_2),.din(w_dff_A_tShaQ5nr3_2),.clk(gclk));
	jdff dff_A_OAWtnM404_2(.dout(w_dff_A_tShaQ5nr3_2),.din(w_dff_A_OAWtnM404_2),.clk(gclk));
	jdff dff_A_qdqH9rKd4_2(.dout(w_dff_A_OAWtnM404_2),.din(w_dff_A_qdqH9rKd4_2),.clk(gclk));
	jdff dff_A_blZP9Hfz6_2(.dout(w_dff_A_qdqH9rKd4_2),.din(w_dff_A_blZP9Hfz6_2),.clk(gclk));
	jdff dff_A_w1EBiFrA3_2(.dout(w_dff_A_blZP9Hfz6_2),.din(w_dff_A_w1EBiFrA3_2),.clk(gclk));
	jdff dff_A_8X7AsI6h6_0(.dout(w_G4088_6[0]),.din(w_dff_A_8X7AsI6h6_0),.clk(gclk));
	jdff dff_A_ZVZPeOv60_0(.dout(w_dff_A_8X7AsI6h6_0),.din(w_dff_A_ZVZPeOv60_0),.clk(gclk));
	jdff dff_A_Kz9vVoEa0_0(.dout(w_dff_A_ZVZPeOv60_0),.din(w_dff_A_Kz9vVoEa0_0),.clk(gclk));
	jdff dff_A_dpSplsPl5_0(.dout(w_dff_A_Kz9vVoEa0_0),.din(w_dff_A_dpSplsPl5_0),.clk(gclk));
	jdff dff_A_GgguOPOl9_0(.dout(w_dff_A_dpSplsPl5_0),.din(w_dff_A_GgguOPOl9_0),.clk(gclk));
	jdff dff_A_WLwsBMxg3_0(.dout(w_dff_A_GgguOPOl9_0),.din(w_dff_A_WLwsBMxg3_0),.clk(gclk));
	jdff dff_A_vBD5oPDR3_0(.dout(w_dff_A_WLwsBMxg3_0),.din(w_dff_A_vBD5oPDR3_0),.clk(gclk));
	jdff dff_A_Jf6CIFIy8_0(.dout(w_dff_A_vBD5oPDR3_0),.din(w_dff_A_Jf6CIFIy8_0),.clk(gclk));
	jdff dff_A_ggBehG243_0(.dout(w_dff_A_Jf6CIFIy8_0),.din(w_dff_A_ggBehG243_0),.clk(gclk));
	jdff dff_A_AMZqHj9V9_0(.dout(w_dff_A_ggBehG243_0),.din(w_dff_A_AMZqHj9V9_0),.clk(gclk));
	jdff dff_A_ogHOGOfJ8_0(.dout(w_dff_A_AMZqHj9V9_0),.din(w_dff_A_ogHOGOfJ8_0),.clk(gclk));
	jdff dff_A_qH8pCZaJ4_0(.dout(w_dff_A_ogHOGOfJ8_0),.din(w_dff_A_qH8pCZaJ4_0),.clk(gclk));
	jdff dff_A_wmvximqy1_0(.dout(w_dff_A_qH8pCZaJ4_0),.din(w_dff_A_wmvximqy1_0),.clk(gclk));
	jdff dff_A_LeDPvtRG1_2(.dout(w_G4088_6[2]),.din(w_dff_A_LeDPvtRG1_2),.clk(gclk));
	jdff dff_A_Uyg8AFmx8_2(.dout(w_dff_A_LeDPvtRG1_2),.din(w_dff_A_Uyg8AFmx8_2),.clk(gclk));
	jdff dff_A_Fj7z8uzD1_2(.dout(w_dff_A_Uyg8AFmx8_2),.din(w_dff_A_Fj7z8uzD1_2),.clk(gclk));
	jdff dff_A_Vd5jpfGX2_2(.dout(w_dff_A_Fj7z8uzD1_2),.din(w_dff_A_Vd5jpfGX2_2),.clk(gclk));
	jdff dff_A_N8utaI5B1_2(.dout(w_dff_A_Vd5jpfGX2_2),.din(w_dff_A_N8utaI5B1_2),.clk(gclk));
	jdff dff_A_KZnepCYa3_2(.dout(w_dff_A_N8utaI5B1_2),.din(w_dff_A_KZnepCYa3_2),.clk(gclk));
	jdff dff_A_T1rtKHIl4_2(.dout(w_dff_A_KZnepCYa3_2),.din(w_dff_A_T1rtKHIl4_2),.clk(gclk));
	jdff dff_A_6NJ7VYnd6_2(.dout(w_dff_A_T1rtKHIl4_2),.din(w_dff_A_6NJ7VYnd6_2),.clk(gclk));
	jdff dff_A_R7j4hwe17_2(.dout(w_dff_A_6NJ7VYnd6_2),.din(w_dff_A_R7j4hwe17_2),.clk(gclk));
	jdff dff_A_aO7SEFju5_2(.dout(w_dff_A_R7j4hwe17_2),.din(w_dff_A_aO7SEFju5_2),.clk(gclk));
	jdff dff_B_4bNGrXUQ9_0(.din(n1286),.dout(w_dff_B_4bNGrXUQ9_0),.clk(gclk));
	jdff dff_B_07wly5Ol4_0(.din(w_dff_B_4bNGrXUQ9_0),.dout(w_dff_B_07wly5Ol4_0),.clk(gclk));
	jdff dff_B_56WsX3sS6_0(.din(w_dff_B_07wly5Ol4_0),.dout(w_dff_B_56WsX3sS6_0),.clk(gclk));
	jdff dff_B_dbuNXJN80_0(.din(w_dff_B_56WsX3sS6_0),.dout(w_dff_B_dbuNXJN80_0),.clk(gclk));
	jdff dff_B_DuhFN4vE0_0(.din(w_dff_B_dbuNXJN80_0),.dout(w_dff_B_DuhFN4vE0_0),.clk(gclk));
	jdff dff_B_HlmbQFyF2_0(.din(w_dff_B_DuhFN4vE0_0),.dout(w_dff_B_HlmbQFyF2_0),.clk(gclk));
	jdff dff_B_9IIJg3y20_0(.din(w_dff_B_HlmbQFyF2_0),.dout(w_dff_B_9IIJg3y20_0),.clk(gclk));
	jdff dff_B_P0P025ms5_0(.din(w_dff_B_9IIJg3y20_0),.dout(w_dff_B_P0P025ms5_0),.clk(gclk));
	jdff dff_B_MqEipejA5_0(.din(w_dff_B_P0P025ms5_0),.dout(w_dff_B_MqEipejA5_0),.clk(gclk));
	jdff dff_B_Fp31TEwl9_0(.din(w_dff_B_MqEipejA5_0),.dout(w_dff_B_Fp31TEwl9_0),.clk(gclk));
	jdff dff_B_7nnYvt1J9_0(.din(w_dff_B_Fp31TEwl9_0),.dout(w_dff_B_7nnYvt1J9_0),.clk(gclk));
	jdff dff_B_qAfv0Rnk6_0(.din(w_dff_B_7nnYvt1J9_0),.dout(w_dff_B_qAfv0Rnk6_0),.clk(gclk));
	jdff dff_B_pguaHEhJ4_0(.din(w_dff_B_qAfv0Rnk6_0),.dout(w_dff_B_pguaHEhJ4_0),.clk(gclk));
	jdff dff_B_CyOCDMME2_0(.din(w_dff_B_pguaHEhJ4_0),.dout(w_dff_B_CyOCDMME2_0),.clk(gclk));
	jdff dff_B_fbzNMePi9_0(.din(w_dff_B_CyOCDMME2_0),.dout(w_dff_B_fbzNMePi9_0),.clk(gclk));
	jdff dff_B_ozTQxUHt5_1(.din(n1278),.dout(w_dff_B_ozTQxUHt5_1),.clk(gclk));
	jdff dff_B_M8TbZGfO8_1(.din(w_dff_B_ozTQxUHt5_1),.dout(w_dff_B_M8TbZGfO8_1),.clk(gclk));
	jdff dff_B_VvxiDDw61_1(.din(w_dff_B_M8TbZGfO8_1),.dout(w_dff_B_VvxiDDw61_1),.clk(gclk));
	jdff dff_A_61hyrzFl7_1(.dout(w_n797_5[1]),.din(w_dff_A_61hyrzFl7_1),.clk(gclk));
	jdff dff_A_YosYbhOc1_1(.dout(w_dff_A_61hyrzFl7_1),.din(w_dff_A_YosYbhOc1_1),.clk(gclk));
	jdff dff_A_fifs4hFG3_1(.dout(w_dff_A_YosYbhOc1_1),.din(w_dff_A_fifs4hFG3_1),.clk(gclk));
	jdff dff_A_XebadTqn6_1(.dout(w_dff_A_fifs4hFG3_1),.din(w_dff_A_XebadTqn6_1),.clk(gclk));
	jdff dff_A_m5QyaTK99_1(.dout(w_dff_A_XebadTqn6_1),.din(w_dff_A_m5QyaTK99_1),.clk(gclk));
	jdff dff_A_awIwdeP06_1(.dout(w_dff_A_m5QyaTK99_1),.din(w_dff_A_awIwdeP06_1),.clk(gclk));
	jdff dff_A_I3aCi0CK7_1(.dout(w_dff_A_awIwdeP06_1),.din(w_dff_A_I3aCi0CK7_1),.clk(gclk));
	jdff dff_A_mkestAyB1_1(.dout(w_dff_A_I3aCi0CK7_1),.din(w_dff_A_mkestAyB1_1),.clk(gclk));
	jdff dff_A_FnL4gZXA3_1(.dout(w_dff_A_mkestAyB1_1),.din(w_dff_A_FnL4gZXA3_1),.clk(gclk));
	jdff dff_A_5MYECC5F6_1(.dout(w_dff_A_FnL4gZXA3_1),.din(w_dff_A_5MYECC5F6_1),.clk(gclk));
	jdff dff_A_QKLOlKfY0_1(.dout(w_dff_A_5MYECC5F6_1),.din(w_dff_A_QKLOlKfY0_1),.clk(gclk));
	jdff dff_A_QaMlli2f3_1(.dout(w_dff_A_QKLOlKfY0_1),.din(w_dff_A_QaMlli2f3_1),.clk(gclk));
	jdff dff_A_gRAkpv5i7_1(.dout(w_dff_A_QaMlli2f3_1),.din(w_dff_A_gRAkpv5i7_1),.clk(gclk));
	jdff dff_A_83cHrO3Z0_1(.dout(w_dff_A_gRAkpv5i7_1),.din(w_dff_A_83cHrO3Z0_1),.clk(gclk));
	jdff dff_A_tUFwpcmo8_1(.dout(w_G4088_5[1]),.din(w_dff_A_tUFwpcmo8_1),.clk(gclk));
	jdff dff_A_MFEXzr504_1(.dout(w_dff_A_tUFwpcmo8_1),.din(w_dff_A_MFEXzr504_1),.clk(gclk));
	jdff dff_A_6RRPLTSU8_1(.dout(w_dff_A_MFEXzr504_1),.din(w_dff_A_6RRPLTSU8_1),.clk(gclk));
	jdff dff_A_HLeZWtBx3_1(.dout(w_dff_A_6RRPLTSU8_1),.din(w_dff_A_HLeZWtBx3_1),.clk(gclk));
	jdff dff_A_J21HaI1L7_1(.dout(w_dff_A_HLeZWtBx3_1),.din(w_dff_A_J21HaI1L7_1),.clk(gclk));
	jdff dff_A_KzwLaXnn5_1(.dout(w_dff_A_J21HaI1L7_1),.din(w_dff_A_KzwLaXnn5_1),.clk(gclk));
	jdff dff_A_raXqmRL08_1(.dout(w_dff_A_KzwLaXnn5_1),.din(w_dff_A_raXqmRL08_1),.clk(gclk));
	jdff dff_A_2LiweVeY7_1(.dout(w_dff_A_raXqmRL08_1),.din(w_dff_A_2LiweVeY7_1),.clk(gclk));
	jdff dff_A_lwEotw011_1(.dout(w_dff_A_2LiweVeY7_1),.din(w_dff_A_lwEotw011_1),.clk(gclk));
	jdff dff_A_AH3fLX0w5_1(.dout(w_dff_A_lwEotw011_1),.din(w_dff_A_AH3fLX0w5_1),.clk(gclk));
	jdff dff_A_ETld6wek7_1(.dout(w_dff_A_AH3fLX0w5_1),.din(w_dff_A_ETld6wek7_1),.clk(gclk));
	jdff dff_A_sjYm9l1t9_1(.dout(w_dff_A_ETld6wek7_1),.din(w_dff_A_sjYm9l1t9_1),.clk(gclk));
	jdff dff_A_aBzkJTVZ8_1(.dout(w_dff_A_sjYm9l1t9_1),.din(w_dff_A_aBzkJTVZ8_1),.clk(gclk));
	jdff dff_B_RVRPJh1j7_0(.din(n1295),.dout(w_dff_B_RVRPJh1j7_0),.clk(gclk));
	jdff dff_B_rqBZ1JQI3_0(.din(w_dff_B_RVRPJh1j7_0),.dout(w_dff_B_rqBZ1JQI3_0),.clk(gclk));
	jdff dff_B_LwpIlTuo8_0(.din(w_dff_B_rqBZ1JQI3_0),.dout(w_dff_B_LwpIlTuo8_0),.clk(gclk));
	jdff dff_B_5HhsiZ1R5_0(.din(w_dff_B_LwpIlTuo8_0),.dout(w_dff_B_5HhsiZ1R5_0),.clk(gclk));
	jdff dff_B_aRBGPgfP2_0(.din(w_dff_B_5HhsiZ1R5_0),.dout(w_dff_B_aRBGPgfP2_0),.clk(gclk));
	jdff dff_B_zYZ7TxIn0_0(.din(w_dff_B_aRBGPgfP2_0),.dout(w_dff_B_zYZ7TxIn0_0),.clk(gclk));
	jdff dff_B_LskRZRaP1_0(.din(w_dff_B_zYZ7TxIn0_0),.dout(w_dff_B_LskRZRaP1_0),.clk(gclk));
	jdff dff_B_dqXOf1pv5_0(.din(w_dff_B_LskRZRaP1_0),.dout(w_dff_B_dqXOf1pv5_0),.clk(gclk));
	jdff dff_B_0Ej2agMG2_0(.din(w_dff_B_dqXOf1pv5_0),.dout(w_dff_B_0Ej2agMG2_0),.clk(gclk));
	jdff dff_B_2nWOtnAg5_0(.din(w_dff_B_0Ej2agMG2_0),.dout(w_dff_B_2nWOtnAg5_0),.clk(gclk));
	jdff dff_B_JodKFaiP1_0(.din(w_dff_B_2nWOtnAg5_0),.dout(w_dff_B_JodKFaiP1_0),.clk(gclk));
	jdff dff_B_iR0DYSKz7_0(.din(w_dff_B_JodKFaiP1_0),.dout(w_dff_B_iR0DYSKz7_0),.clk(gclk));
	jdff dff_B_8JZi2Twq7_0(.din(w_dff_B_iR0DYSKz7_0),.dout(w_dff_B_8JZi2Twq7_0),.clk(gclk));
	jdff dff_B_3RpqSXkc4_0(.din(w_dff_B_8JZi2Twq7_0),.dout(w_dff_B_3RpqSXkc4_0),.clk(gclk));
	jdff dff_B_JomtzdNK1_1(.din(n1288),.dout(w_dff_B_JomtzdNK1_1),.clk(gclk));
	jdff dff_B_CkXm9KeI4_1(.din(w_dff_B_JomtzdNK1_1),.dout(w_dff_B_CkXm9KeI4_1),.clk(gclk));
	jdff dff_B_CFSdghtJ8_1(.din(w_dff_B_CkXm9KeI4_1),.dout(w_dff_B_CFSdghtJ8_1),.clk(gclk));
	jdff dff_A_VSsgog7F1_1(.dout(w_n800_2[1]),.din(w_dff_A_VSsgog7F1_1),.clk(gclk));
	jdff dff_A_PnFovOBO9_2(.dout(w_n800_2[2]),.din(w_dff_A_PnFovOBO9_2),.clk(gclk));
	jdff dff_B_2daa77Bo1_0(.din(n1306),.dout(w_dff_B_2daa77Bo1_0),.clk(gclk));
	jdff dff_B_y3IsT7Ic0_0(.din(w_dff_B_2daa77Bo1_0),.dout(w_dff_B_y3IsT7Ic0_0),.clk(gclk));
	jdff dff_B_mxCDFJq14_0(.din(w_dff_B_y3IsT7Ic0_0),.dout(w_dff_B_mxCDFJq14_0),.clk(gclk));
	jdff dff_B_iWbjM1nD3_0(.din(w_dff_B_mxCDFJq14_0),.dout(w_dff_B_iWbjM1nD3_0),.clk(gclk));
	jdff dff_B_A3D80apv4_0(.din(w_dff_B_iWbjM1nD3_0),.dout(w_dff_B_A3D80apv4_0),.clk(gclk));
	jdff dff_B_vGlipJHY2_0(.din(w_dff_B_A3D80apv4_0),.dout(w_dff_B_vGlipJHY2_0),.clk(gclk));
	jdff dff_B_3fVfgQg17_0(.din(w_dff_B_vGlipJHY2_0),.dout(w_dff_B_3fVfgQg17_0),.clk(gclk));
	jdff dff_B_hUH6JMAN9_0(.din(w_dff_B_3fVfgQg17_0),.dout(w_dff_B_hUH6JMAN9_0),.clk(gclk));
	jdff dff_B_UkIEKpXw8_0(.din(w_dff_B_hUH6JMAN9_0),.dout(w_dff_B_UkIEKpXw8_0),.clk(gclk));
	jdff dff_B_aZyKo8Bx4_0(.din(w_dff_B_UkIEKpXw8_0),.dout(w_dff_B_aZyKo8Bx4_0),.clk(gclk));
	jdff dff_B_hju0W5HN8_0(.din(w_dff_B_aZyKo8Bx4_0),.dout(w_dff_B_hju0W5HN8_0),.clk(gclk));
	jdff dff_B_51FasEN76_0(.din(w_dff_B_hju0W5HN8_0),.dout(w_dff_B_51FasEN76_0),.clk(gclk));
	jdff dff_B_kZpqylnS4_0(.din(w_dff_B_51FasEN76_0),.dout(w_dff_B_kZpqylnS4_0),.clk(gclk));
	jdff dff_B_dxwp7vRm7_0(.din(w_dff_B_kZpqylnS4_0),.dout(w_dff_B_dxwp7vRm7_0),.clk(gclk));
	jdff dff_B_xeFe8tDL3_0(.din(w_dff_B_dxwp7vRm7_0),.dout(w_dff_B_xeFe8tDL3_0),.clk(gclk));
	jdff dff_B_R6k2vql07_1(.din(n1298),.dout(w_dff_B_R6k2vql07_1),.clk(gclk));
	jdff dff_B_KgK6Eytl0_1(.din(w_dff_B_R6k2vql07_1),.dout(w_dff_B_KgK6Eytl0_1),.clk(gclk));
	jdff dff_B_DCa37vzH1_1(.din(w_dff_B_KgK6Eytl0_1),.dout(w_dff_B_DCa37vzH1_1),.clk(gclk));
	jdff dff_A_3dhf2zH69_0(.dout(w_n797_4[0]),.din(w_dff_A_3dhf2zH69_0),.clk(gclk));
	jdff dff_A_PKD4sYhK0_0(.dout(w_dff_A_3dhf2zH69_0),.din(w_dff_A_PKD4sYhK0_0),.clk(gclk));
	jdff dff_A_X5907bwN2_0(.dout(w_dff_A_PKD4sYhK0_0),.din(w_dff_A_X5907bwN2_0),.clk(gclk));
	jdff dff_A_ftdpoaOF7_0(.dout(w_dff_A_X5907bwN2_0),.din(w_dff_A_ftdpoaOF7_0),.clk(gclk));
	jdff dff_A_gfXIgObn6_0(.dout(w_dff_A_ftdpoaOF7_0),.din(w_dff_A_gfXIgObn6_0),.clk(gclk));
	jdff dff_A_aGWmHD8e7_0(.dout(w_dff_A_gfXIgObn6_0),.din(w_dff_A_aGWmHD8e7_0),.clk(gclk));
	jdff dff_A_zRzgAmkL3_0(.dout(w_dff_A_aGWmHD8e7_0),.din(w_dff_A_zRzgAmkL3_0),.clk(gclk));
	jdff dff_A_duxIveYA0_0(.dout(w_dff_A_zRzgAmkL3_0),.din(w_dff_A_duxIveYA0_0),.clk(gclk));
	jdff dff_A_ulhTxpCP3_0(.dout(w_dff_A_duxIveYA0_0),.din(w_dff_A_ulhTxpCP3_0),.clk(gclk));
	jdff dff_A_O0yG5oUA9_0(.dout(w_dff_A_ulhTxpCP3_0),.din(w_dff_A_O0yG5oUA9_0),.clk(gclk));
	jdff dff_A_mEXwCAXT9_0(.dout(w_dff_A_O0yG5oUA9_0),.din(w_dff_A_mEXwCAXT9_0),.clk(gclk));
	jdff dff_A_ErQlNHns9_0(.dout(w_dff_A_mEXwCAXT9_0),.din(w_dff_A_ErQlNHns9_0),.clk(gclk));
	jdff dff_A_z9bYcK5w1_0(.dout(w_dff_A_ErQlNHns9_0),.din(w_dff_A_z9bYcK5w1_0),.clk(gclk));
	jdff dff_A_drLVlnn43_0(.dout(w_dff_A_z9bYcK5w1_0),.din(w_dff_A_drLVlnn43_0),.clk(gclk));
	jdff dff_A_le1zyTkC4_2(.dout(w_n797_4[2]),.din(w_dff_A_le1zyTkC4_2),.clk(gclk));
	jdff dff_A_PqxpfCk62_2(.dout(w_dff_A_le1zyTkC4_2),.din(w_dff_A_PqxpfCk62_2),.clk(gclk));
	jdff dff_A_aTmrLBR34_2(.dout(w_dff_A_PqxpfCk62_2),.din(w_dff_A_aTmrLBR34_2),.clk(gclk));
	jdff dff_A_Pq8d67pW6_2(.dout(w_dff_A_aTmrLBR34_2),.din(w_dff_A_Pq8d67pW6_2),.clk(gclk));
	jdff dff_A_PAzRvVhk5_2(.dout(w_dff_A_Pq8d67pW6_2),.din(w_dff_A_PAzRvVhk5_2),.clk(gclk));
	jdff dff_A_mhv7YP2y6_2(.dout(w_dff_A_PAzRvVhk5_2),.din(w_dff_A_mhv7YP2y6_2),.clk(gclk));
	jdff dff_A_YcDjhT8T3_2(.dout(w_dff_A_mhv7YP2y6_2),.din(w_dff_A_YcDjhT8T3_2),.clk(gclk));
	jdff dff_A_9tAP6bGr6_2(.dout(w_dff_A_YcDjhT8T3_2),.din(w_dff_A_9tAP6bGr6_2),.clk(gclk));
	jdff dff_A_ssWpAkUp1_2(.dout(w_dff_A_9tAP6bGr6_2),.din(w_dff_A_ssWpAkUp1_2),.clk(gclk));
	jdff dff_A_XgDTtMqh7_2(.dout(w_dff_A_ssWpAkUp1_2),.din(w_dff_A_XgDTtMqh7_2),.clk(gclk));
	jdff dff_A_BgfEetLh3_2(.dout(w_dff_A_XgDTtMqh7_2),.din(w_dff_A_BgfEetLh3_2),.clk(gclk));
	jdff dff_A_OsqZJsAF7_2(.dout(w_dff_A_BgfEetLh3_2),.din(w_dff_A_OsqZJsAF7_2),.clk(gclk));
	jdff dff_A_Jk8JySbY0_2(.dout(w_dff_A_OsqZJsAF7_2),.din(w_dff_A_Jk8JySbY0_2),.clk(gclk));
	jdff dff_A_9qaF3s5p9_0(.dout(w_G4088_4[0]),.din(w_dff_A_9qaF3s5p9_0),.clk(gclk));
	jdff dff_A_7fm7OJu09_0(.dout(w_dff_A_9qaF3s5p9_0),.din(w_dff_A_7fm7OJu09_0),.clk(gclk));
	jdff dff_A_jyxjwfih5_0(.dout(w_dff_A_7fm7OJu09_0),.din(w_dff_A_jyxjwfih5_0),.clk(gclk));
	jdff dff_A_2S7sEQvu7_0(.dout(w_dff_A_jyxjwfih5_0),.din(w_dff_A_2S7sEQvu7_0),.clk(gclk));
	jdff dff_A_MSD0T39I1_0(.dout(w_dff_A_2S7sEQvu7_0),.din(w_dff_A_MSD0T39I1_0),.clk(gclk));
	jdff dff_A_7Zw8XIoB1_0(.dout(w_dff_A_MSD0T39I1_0),.din(w_dff_A_7Zw8XIoB1_0),.clk(gclk));
	jdff dff_A_0HY2OVzG1_0(.dout(w_dff_A_7Zw8XIoB1_0),.din(w_dff_A_0HY2OVzG1_0),.clk(gclk));
	jdff dff_A_62iO4Jzp4_0(.dout(w_dff_A_0HY2OVzG1_0),.din(w_dff_A_62iO4Jzp4_0),.clk(gclk));
	jdff dff_A_CT3P7VP80_0(.dout(w_dff_A_62iO4Jzp4_0),.din(w_dff_A_CT3P7VP80_0),.clk(gclk));
	jdff dff_A_iy7aQw1i7_0(.dout(w_dff_A_CT3P7VP80_0),.din(w_dff_A_iy7aQw1i7_0),.clk(gclk));
	jdff dff_A_KdpGOKs31_0(.dout(w_dff_A_iy7aQw1i7_0),.din(w_dff_A_KdpGOKs31_0),.clk(gclk));
	jdff dff_A_DeriYlGF3_0(.dout(w_dff_A_KdpGOKs31_0),.din(w_dff_A_DeriYlGF3_0),.clk(gclk));
	jdff dff_A_GtycS8g76_0(.dout(w_dff_A_DeriYlGF3_0),.din(w_dff_A_GtycS8g76_0),.clk(gclk));
	jdff dff_A_FMu5tN8o6_2(.dout(w_G4088_4[2]),.din(w_dff_A_FMu5tN8o6_2),.clk(gclk));
	jdff dff_A_9sHGJc3t5_2(.dout(w_dff_A_FMu5tN8o6_2),.din(w_dff_A_9sHGJc3t5_2),.clk(gclk));
	jdff dff_A_NXiR1U0V0_2(.dout(w_dff_A_9sHGJc3t5_2),.din(w_dff_A_NXiR1U0V0_2),.clk(gclk));
	jdff dff_A_2sNnIkIh8_2(.dout(w_dff_A_NXiR1U0V0_2),.din(w_dff_A_2sNnIkIh8_2),.clk(gclk));
	jdff dff_A_xmUYwhiP2_2(.dout(w_dff_A_2sNnIkIh8_2),.din(w_dff_A_xmUYwhiP2_2),.clk(gclk));
	jdff dff_A_O1X7TDLI6_2(.dout(w_dff_A_xmUYwhiP2_2),.din(w_dff_A_O1X7TDLI6_2),.clk(gclk));
	jdff dff_A_5SehsGnv5_2(.dout(w_dff_A_O1X7TDLI6_2),.din(w_dff_A_5SehsGnv5_2),.clk(gclk));
	jdff dff_A_yB35zGkT9_2(.dout(w_dff_A_5SehsGnv5_2),.din(w_dff_A_yB35zGkT9_2),.clk(gclk));
	jdff dff_A_BLaCUOQs4_2(.dout(w_dff_A_yB35zGkT9_2),.din(w_dff_A_BLaCUOQs4_2),.clk(gclk));
	jdff dff_A_ygAWogll4_2(.dout(w_dff_A_BLaCUOQs4_2),.din(w_dff_A_ygAWogll4_2),.clk(gclk));
	jdff dff_A_KE703snk8_2(.dout(w_dff_A_ygAWogll4_2),.din(w_dff_A_KE703snk8_2),.clk(gclk));
	jdff dff_A_UR13TOBk4_2(.dout(w_dff_A_KE703snk8_2),.din(w_dff_A_UR13TOBk4_2),.clk(gclk));
	jdff dff_B_TPOkjn7r9_0(.din(n1315),.dout(w_dff_B_TPOkjn7r9_0),.clk(gclk));
	jdff dff_B_p8ObpuHO3_0(.din(w_dff_B_TPOkjn7r9_0),.dout(w_dff_B_p8ObpuHO3_0),.clk(gclk));
	jdff dff_B_RfTKynf52_0(.din(w_dff_B_p8ObpuHO3_0),.dout(w_dff_B_RfTKynf52_0),.clk(gclk));
	jdff dff_B_63rkuWgi5_0(.din(w_dff_B_RfTKynf52_0),.dout(w_dff_B_63rkuWgi5_0),.clk(gclk));
	jdff dff_B_QEICD4B38_0(.din(w_dff_B_63rkuWgi5_0),.dout(w_dff_B_QEICD4B38_0),.clk(gclk));
	jdff dff_B_GMDvtPfY9_0(.din(w_dff_B_QEICD4B38_0),.dout(w_dff_B_GMDvtPfY9_0),.clk(gclk));
	jdff dff_B_7dm3CGsX4_0(.din(w_dff_B_GMDvtPfY9_0),.dout(w_dff_B_7dm3CGsX4_0),.clk(gclk));
	jdff dff_B_sIaBciIM1_0(.din(w_dff_B_7dm3CGsX4_0),.dout(w_dff_B_sIaBciIM1_0),.clk(gclk));
	jdff dff_B_aRrUP5Cf8_0(.din(w_dff_B_sIaBciIM1_0),.dout(w_dff_B_aRrUP5Cf8_0),.clk(gclk));
	jdff dff_B_FxrUoyKA7_0(.din(w_dff_B_aRrUP5Cf8_0),.dout(w_dff_B_FxrUoyKA7_0),.clk(gclk));
	jdff dff_B_h57xBb8Q8_0(.din(w_dff_B_FxrUoyKA7_0),.dout(w_dff_B_h57xBb8Q8_0),.clk(gclk));
	jdff dff_B_KGCyfljf0_0(.din(w_dff_B_h57xBb8Q8_0),.dout(w_dff_B_KGCyfljf0_0),.clk(gclk));
	jdff dff_B_byXYpk5q8_0(.din(w_dff_B_KGCyfljf0_0),.dout(w_dff_B_byXYpk5q8_0),.clk(gclk));
	jdff dff_B_32PVOr4o8_0(.din(w_dff_B_byXYpk5q8_0),.dout(w_dff_B_32PVOr4o8_0),.clk(gclk));
	jdff dff_B_IBbsAM0P4_0(.din(w_dff_B_32PVOr4o8_0),.dout(w_dff_B_IBbsAM0P4_0),.clk(gclk));
	jdff dff_B_FAo4GoRd6_2(.din(G49),.dout(w_dff_B_FAo4GoRd6_2),.clk(gclk));
	jdff dff_B_hnCBB4eR5_1(.din(n1308),.dout(w_dff_B_hnCBB4eR5_1),.clk(gclk));
	jdff dff_B_DyAbswhy2_1(.din(w_dff_B_hnCBB4eR5_1),.dout(w_dff_B_DyAbswhy2_1),.clk(gclk));
	jdff dff_B_jxdHE5yx0_1(.din(w_dff_B_DyAbswhy2_1),.dout(w_dff_B_jxdHE5yx0_1),.clk(gclk));
	jdff dff_A_6aP60U6S4_1(.dout(w_n852_5[1]),.din(w_dff_A_6aP60U6S4_1),.clk(gclk));
	jdff dff_A_fgkpfRl94_1(.dout(w_dff_A_6aP60U6S4_1),.din(w_dff_A_fgkpfRl94_1),.clk(gclk));
	jdff dff_A_QfBA7mrf1_1(.dout(w_dff_A_fgkpfRl94_1),.din(w_dff_A_QfBA7mrf1_1),.clk(gclk));
	jdff dff_A_OvoeYs2x9_1(.dout(w_dff_A_QfBA7mrf1_1),.din(w_dff_A_OvoeYs2x9_1),.clk(gclk));
	jdff dff_A_FBcZg9x53_1(.dout(w_dff_A_OvoeYs2x9_1),.din(w_dff_A_FBcZg9x53_1),.clk(gclk));
	jdff dff_A_Holf9ScS6_1(.dout(w_dff_A_FBcZg9x53_1),.din(w_dff_A_Holf9ScS6_1),.clk(gclk));
	jdff dff_A_7l85le1F3_1(.dout(w_dff_A_Holf9ScS6_1),.din(w_dff_A_7l85le1F3_1),.clk(gclk));
	jdff dff_A_wpAQBJA69_1(.dout(w_dff_A_7l85le1F3_1),.din(w_dff_A_wpAQBJA69_1),.clk(gclk));
	jdff dff_A_2AfTwmzk5_1(.dout(w_dff_A_wpAQBJA69_1),.din(w_dff_A_2AfTwmzk5_1),.clk(gclk));
	jdff dff_A_N0ozBPZ51_1(.dout(w_dff_A_2AfTwmzk5_1),.din(w_dff_A_N0ozBPZ51_1),.clk(gclk));
	jdff dff_A_66Jggwrk1_1(.dout(w_dff_A_N0ozBPZ51_1),.din(w_dff_A_66Jggwrk1_1),.clk(gclk));
	jdff dff_A_QaoKRL2z1_1(.dout(w_dff_A_66Jggwrk1_1),.din(w_dff_A_QaoKRL2z1_1),.clk(gclk));
	jdff dff_A_JC9hUCkI0_1(.dout(w_dff_A_QaoKRL2z1_1),.din(w_dff_A_JC9hUCkI0_1),.clk(gclk));
	jdff dff_A_0wRL0BA83_1(.dout(w_dff_A_JC9hUCkI0_1),.din(w_dff_A_0wRL0BA83_1),.clk(gclk));
	jdff dff_A_wtQfZ54e8_2(.dout(w_n852_5[2]),.din(w_dff_A_wtQfZ54e8_2),.clk(gclk));
	jdff dff_A_3s2nxqKQ7_2(.dout(w_dff_A_wtQfZ54e8_2),.din(w_dff_A_3s2nxqKQ7_2),.clk(gclk));
	jdff dff_A_GWVoku2z4_2(.dout(w_dff_A_3s2nxqKQ7_2),.din(w_dff_A_GWVoku2z4_2),.clk(gclk));
	jdff dff_A_8FAIC1IA6_2(.dout(w_dff_A_GWVoku2z4_2),.din(w_dff_A_8FAIC1IA6_2),.clk(gclk));
	jdff dff_A_UNXSZwcO3_2(.dout(w_dff_A_8FAIC1IA6_2),.din(w_dff_A_UNXSZwcO3_2),.clk(gclk));
	jdff dff_A_nUGKIQoW7_2(.dout(w_dff_A_UNXSZwcO3_2),.din(w_dff_A_nUGKIQoW7_2),.clk(gclk));
	jdff dff_A_OL45Dp2D4_2(.dout(w_dff_A_nUGKIQoW7_2),.din(w_dff_A_OL45Dp2D4_2),.clk(gclk));
	jdff dff_A_EIgBiJQD5_2(.dout(w_dff_A_OL45Dp2D4_2),.din(w_dff_A_EIgBiJQD5_2),.clk(gclk));
	jdff dff_A_iqcoUGm54_2(.dout(w_dff_A_EIgBiJQD5_2),.din(w_dff_A_iqcoUGm54_2),.clk(gclk));
	jdff dff_A_VAGYgt9E0_2(.dout(w_dff_A_iqcoUGm54_2),.din(w_dff_A_VAGYgt9E0_2),.clk(gclk));
	jdff dff_A_3UeJjg4D4_2(.dout(w_dff_A_VAGYgt9E0_2),.din(w_dff_A_3UeJjg4D4_2),.clk(gclk));
	jdff dff_A_VwWoXtQT7_2(.dout(w_dff_A_3UeJjg4D4_2),.din(w_dff_A_VwWoXtQT7_2),.clk(gclk));
	jdff dff_A_lVk8emyb5_2(.dout(w_dff_A_VwWoXtQT7_2),.din(w_dff_A_lVk8emyb5_2),.clk(gclk));
	jdff dff_A_2rHcka5g9_2(.dout(w_dff_A_lVk8emyb5_2),.din(w_dff_A_2rHcka5g9_2),.clk(gclk));
	jdff dff_A_pNqj457g1_1(.dout(w_G4089_5[1]),.din(w_dff_A_pNqj457g1_1),.clk(gclk));
	jdff dff_A_iNC929Ew3_1(.dout(w_dff_A_pNqj457g1_1),.din(w_dff_A_iNC929Ew3_1),.clk(gclk));
	jdff dff_A_v0z2JNA78_1(.dout(w_dff_A_iNC929Ew3_1),.din(w_dff_A_v0z2JNA78_1),.clk(gclk));
	jdff dff_A_ynkmJDs31_1(.dout(w_dff_A_v0z2JNA78_1),.din(w_dff_A_ynkmJDs31_1),.clk(gclk));
	jdff dff_A_O0fpEPtx0_1(.dout(w_dff_A_ynkmJDs31_1),.din(w_dff_A_O0fpEPtx0_1),.clk(gclk));
	jdff dff_A_WNltdT4J2_1(.dout(w_dff_A_O0fpEPtx0_1),.din(w_dff_A_WNltdT4J2_1),.clk(gclk));
	jdff dff_A_I74UbD4Q0_1(.dout(w_dff_A_WNltdT4J2_1),.din(w_dff_A_I74UbD4Q0_1),.clk(gclk));
	jdff dff_A_AOLGFEfp6_1(.dout(w_dff_A_I74UbD4Q0_1),.din(w_dff_A_AOLGFEfp6_1),.clk(gclk));
	jdff dff_A_xnZJRa9L2_1(.dout(w_dff_A_AOLGFEfp6_1),.din(w_dff_A_xnZJRa9L2_1),.clk(gclk));
	jdff dff_A_fslFyC5k4_1(.dout(w_dff_A_xnZJRa9L2_1),.din(w_dff_A_fslFyC5k4_1),.clk(gclk));
	jdff dff_A_SpFxxcgd2_1(.dout(w_dff_A_fslFyC5k4_1),.din(w_dff_A_SpFxxcgd2_1),.clk(gclk));
	jdff dff_A_dRVvHzKp6_1(.dout(w_dff_A_SpFxxcgd2_1),.din(w_dff_A_dRVvHzKp6_1),.clk(gclk));
	jdff dff_A_QQ3cgWxW8_1(.dout(w_dff_A_dRVvHzKp6_1),.din(w_dff_A_QQ3cgWxW8_1),.clk(gclk));
	jdff dff_A_PIfmCQ6N7_2(.dout(w_G4089_5[2]),.din(w_dff_A_PIfmCQ6N7_2),.clk(gclk));
	jdff dff_A_xwa0luW98_2(.dout(w_dff_A_PIfmCQ6N7_2),.din(w_dff_A_xwa0luW98_2),.clk(gclk));
	jdff dff_A_tp3c67SQ3_2(.dout(w_dff_A_xwa0luW98_2),.din(w_dff_A_tp3c67SQ3_2),.clk(gclk));
	jdff dff_A_tE3ebmNO9_2(.dout(w_dff_A_tp3c67SQ3_2),.din(w_dff_A_tE3ebmNO9_2),.clk(gclk));
	jdff dff_A_mfoznz4J2_2(.dout(w_dff_A_tE3ebmNO9_2),.din(w_dff_A_mfoznz4J2_2),.clk(gclk));
	jdff dff_A_a7hfHu3R2_2(.dout(w_dff_A_mfoznz4J2_2),.din(w_dff_A_a7hfHu3R2_2),.clk(gclk));
	jdff dff_A_hT1yPn2v2_2(.dout(w_dff_A_a7hfHu3R2_2),.din(w_dff_A_hT1yPn2v2_2),.clk(gclk));
	jdff dff_A_Pie7opTS9_2(.dout(w_dff_A_hT1yPn2v2_2),.din(w_dff_A_Pie7opTS9_2),.clk(gclk));
	jdff dff_A_o0Bu0caV0_2(.dout(w_dff_A_Pie7opTS9_2),.din(w_dff_A_o0Bu0caV0_2),.clk(gclk));
	jdff dff_A_g0xY0OlP5_2(.dout(w_dff_A_o0Bu0caV0_2),.din(w_dff_A_g0xY0OlP5_2),.clk(gclk));
	jdff dff_A_nTcqnpTW6_2(.dout(w_dff_A_g0xY0OlP5_2),.din(w_dff_A_nTcqnpTW6_2),.clk(gclk));
	jdff dff_A_GOdr2Bnl9_2(.dout(w_dff_A_nTcqnpTW6_2),.din(w_dff_A_GOdr2Bnl9_2),.clk(gclk));
	jdff dff_A_7jshLYJC7_2(.dout(w_dff_A_GOdr2Bnl9_2),.din(w_dff_A_7jshLYJC7_2),.clk(gclk));
	jdff dff_B_Sg1nqh8g2_0(.din(n1324),.dout(w_dff_B_Sg1nqh8g2_0),.clk(gclk));
	jdff dff_B_8itE12jJ8_0(.din(w_dff_B_Sg1nqh8g2_0),.dout(w_dff_B_8itE12jJ8_0),.clk(gclk));
	jdff dff_B_2bqiqs3G1_0(.din(w_dff_B_8itE12jJ8_0),.dout(w_dff_B_2bqiqs3G1_0),.clk(gclk));
	jdff dff_B_66y0M8Z94_0(.din(w_dff_B_2bqiqs3G1_0),.dout(w_dff_B_66y0M8Z94_0),.clk(gclk));
	jdff dff_B_oVOUaFwl9_0(.din(w_dff_B_66y0M8Z94_0),.dout(w_dff_B_oVOUaFwl9_0),.clk(gclk));
	jdff dff_B_SNIr9ggv9_0(.din(w_dff_B_oVOUaFwl9_0),.dout(w_dff_B_SNIr9ggv9_0),.clk(gclk));
	jdff dff_B_JfUnKVtE0_0(.din(w_dff_B_SNIr9ggv9_0),.dout(w_dff_B_JfUnKVtE0_0),.clk(gclk));
	jdff dff_B_z6QokRgv8_0(.din(w_dff_B_JfUnKVtE0_0),.dout(w_dff_B_z6QokRgv8_0),.clk(gclk));
	jdff dff_B_PIOSjjUD6_0(.din(w_dff_B_z6QokRgv8_0),.dout(w_dff_B_PIOSjjUD6_0),.clk(gclk));
	jdff dff_B_ZsuFXeVN4_0(.din(w_dff_B_PIOSjjUD6_0),.dout(w_dff_B_ZsuFXeVN4_0),.clk(gclk));
	jdff dff_B_zVEyLM8N0_0(.din(w_dff_B_ZsuFXeVN4_0),.dout(w_dff_B_zVEyLM8N0_0),.clk(gclk));
	jdff dff_B_JDCBK7gm0_0(.din(w_dff_B_zVEyLM8N0_0),.dout(w_dff_B_JDCBK7gm0_0),.clk(gclk));
	jdff dff_B_teWfjeAf5_0(.din(w_dff_B_JDCBK7gm0_0),.dout(w_dff_B_teWfjeAf5_0),.clk(gclk));
	jdff dff_B_rfKSEMge0_0(.din(w_dff_B_teWfjeAf5_0),.dout(w_dff_B_rfKSEMge0_0),.clk(gclk));
	jdff dff_A_tSDqlSZB3_2(.dout(w_G4090_2[2]),.din(w_dff_A_tSDqlSZB3_2),.clk(gclk));
	jdff dff_B_HxTIoVvv0_2(.din(G103),.dout(w_dff_B_HxTIoVvv0_2),.clk(gclk));
	jdff dff_B_s8OaSu7E6_1(.din(n1317),.dout(w_dff_B_s8OaSu7E6_1),.clk(gclk));
	jdff dff_B_6zEZas013_1(.din(w_dff_B_s8OaSu7E6_1),.dout(w_dff_B_6zEZas013_1),.clk(gclk));
	jdff dff_B_vOeuLJoV2_1(.din(w_dff_B_6zEZas013_1),.dout(w_dff_B_vOeuLJoV2_1),.clk(gclk));
	jdff dff_A_uPx2Fj0u1_0(.dout(w_n854_2[0]),.din(w_dff_A_uPx2Fj0u1_0),.clk(gclk));
	jdff dff_A_uFQUb5RD5_1(.dout(w_n854_2[1]),.din(w_dff_A_uFQUb5RD5_1),.clk(gclk));
	jdff dff_A_Yb84MPbL5_1(.dout(w_dff_A_uFQUb5RD5_1),.din(w_dff_A_Yb84MPbL5_1),.clk(gclk));
	jdff dff_B_I9jx0YZ58_0(.din(n1333),.dout(w_dff_B_I9jx0YZ58_0),.clk(gclk));
	jdff dff_B_tOBh2K0e2_0(.din(w_dff_B_I9jx0YZ58_0),.dout(w_dff_B_tOBh2K0e2_0),.clk(gclk));
	jdff dff_B_FQjJiZYQ9_0(.din(w_dff_B_tOBh2K0e2_0),.dout(w_dff_B_FQjJiZYQ9_0),.clk(gclk));
	jdff dff_B_GensyDvK0_0(.din(w_dff_B_FQjJiZYQ9_0),.dout(w_dff_B_GensyDvK0_0),.clk(gclk));
	jdff dff_B_cptc2s1c5_0(.din(w_dff_B_GensyDvK0_0),.dout(w_dff_B_cptc2s1c5_0),.clk(gclk));
	jdff dff_B_xj22PHBG8_0(.din(w_dff_B_cptc2s1c5_0),.dout(w_dff_B_xj22PHBG8_0),.clk(gclk));
	jdff dff_B_vPmcNdxc6_0(.din(w_dff_B_xj22PHBG8_0),.dout(w_dff_B_vPmcNdxc6_0),.clk(gclk));
	jdff dff_B_eRivflNn0_0(.din(w_dff_B_vPmcNdxc6_0),.dout(w_dff_B_eRivflNn0_0),.clk(gclk));
	jdff dff_B_RH4Zyh2w2_0(.din(w_dff_B_eRivflNn0_0),.dout(w_dff_B_RH4Zyh2w2_0),.clk(gclk));
	jdff dff_B_CP3Zu8BA1_0(.din(w_dff_B_RH4Zyh2w2_0),.dout(w_dff_B_CP3Zu8BA1_0),.clk(gclk));
	jdff dff_B_IQNqM0gy0_0(.din(w_dff_B_CP3Zu8BA1_0),.dout(w_dff_B_IQNqM0gy0_0),.clk(gclk));
	jdff dff_B_Lkey5Jve4_0(.din(w_dff_B_IQNqM0gy0_0),.dout(w_dff_B_Lkey5Jve4_0),.clk(gclk));
	jdff dff_B_zFvtv3yL9_0(.din(w_dff_B_Lkey5Jve4_0),.dout(w_dff_B_zFvtv3yL9_0),.clk(gclk));
	jdff dff_B_FYUnYL8X0_0(.din(w_dff_B_zFvtv3yL9_0),.dout(w_dff_B_FYUnYL8X0_0),.clk(gclk));
	jdff dff_B_1e1NwGhf7_0(.din(w_dff_B_FYUnYL8X0_0),.dout(w_dff_B_1e1NwGhf7_0),.clk(gclk));
	jdff dff_B_wGJVb2R39_2(.din(G40),.dout(w_dff_B_wGJVb2R39_2),.clk(gclk));
	jdff dff_B_kbhrdEkE0_1(.din(n1326),.dout(w_dff_B_kbhrdEkE0_1),.clk(gclk));
	jdff dff_B_Ywmvo4SI5_1(.din(w_dff_B_kbhrdEkE0_1),.dout(w_dff_B_Ywmvo4SI5_1),.clk(gclk));
	jdff dff_B_vCC4io5f0_1(.din(w_dff_B_Ywmvo4SI5_1),.dout(w_dff_B_vCC4io5f0_1),.clk(gclk));
	jdff dff_A_GY5BZJ6C9_0(.dout(w_n852_4[0]),.din(w_dff_A_GY5BZJ6C9_0),.clk(gclk));
	jdff dff_A_W01AA77Q2_0(.dout(w_dff_A_GY5BZJ6C9_0),.din(w_dff_A_W01AA77Q2_0),.clk(gclk));
	jdff dff_A_lmW0h3uF2_0(.dout(w_dff_A_W01AA77Q2_0),.din(w_dff_A_lmW0h3uF2_0),.clk(gclk));
	jdff dff_A_YX9lb0hU1_0(.dout(w_dff_A_lmW0h3uF2_0),.din(w_dff_A_YX9lb0hU1_0),.clk(gclk));
	jdff dff_A_kZBXivu82_0(.dout(w_dff_A_YX9lb0hU1_0),.din(w_dff_A_kZBXivu82_0),.clk(gclk));
	jdff dff_A_7m510Wrv0_0(.dout(w_dff_A_kZBXivu82_0),.din(w_dff_A_7m510Wrv0_0),.clk(gclk));
	jdff dff_A_Hs43XAUq3_0(.dout(w_dff_A_7m510Wrv0_0),.din(w_dff_A_Hs43XAUq3_0),.clk(gclk));
	jdff dff_A_pFnoTz3C2_0(.dout(w_dff_A_Hs43XAUq3_0),.din(w_dff_A_pFnoTz3C2_0),.clk(gclk));
	jdff dff_A_IBbXRGp16_0(.dout(w_dff_A_pFnoTz3C2_0),.din(w_dff_A_IBbXRGp16_0),.clk(gclk));
	jdff dff_A_JJHqbZGP9_0(.dout(w_dff_A_IBbXRGp16_0),.din(w_dff_A_JJHqbZGP9_0),.clk(gclk));
	jdff dff_A_6Y3XtMLv4_0(.dout(w_dff_A_JJHqbZGP9_0),.din(w_dff_A_6Y3XtMLv4_0),.clk(gclk));
	jdff dff_A_YrhwLuMm5_0(.dout(w_dff_A_6Y3XtMLv4_0),.din(w_dff_A_YrhwLuMm5_0),.clk(gclk));
	jdff dff_A_IGaPKrFy8_0(.dout(w_dff_A_YrhwLuMm5_0),.din(w_dff_A_IGaPKrFy8_0),.clk(gclk));
	jdff dff_A_cCkSWa6R3_0(.dout(w_dff_A_IGaPKrFy8_0),.din(w_dff_A_cCkSWa6R3_0),.clk(gclk));
	jdff dff_A_VuEfhJ3T6_2(.dout(w_n852_4[2]),.din(w_dff_A_VuEfhJ3T6_2),.clk(gclk));
	jdff dff_A_MG3D1TRD1_2(.dout(w_dff_A_VuEfhJ3T6_2),.din(w_dff_A_MG3D1TRD1_2),.clk(gclk));
	jdff dff_A_Ud2VEXUf0_2(.dout(w_dff_A_MG3D1TRD1_2),.din(w_dff_A_Ud2VEXUf0_2),.clk(gclk));
	jdff dff_A_6IZqZPyg9_2(.dout(w_dff_A_Ud2VEXUf0_2),.din(w_dff_A_6IZqZPyg9_2),.clk(gclk));
	jdff dff_A_FGlp4Xtm2_2(.dout(w_dff_A_6IZqZPyg9_2),.din(w_dff_A_FGlp4Xtm2_2),.clk(gclk));
	jdff dff_A_6GbMvlJj3_2(.dout(w_dff_A_FGlp4Xtm2_2),.din(w_dff_A_6GbMvlJj3_2),.clk(gclk));
	jdff dff_A_PPwvwhUc5_2(.dout(w_dff_A_6GbMvlJj3_2),.din(w_dff_A_PPwvwhUc5_2),.clk(gclk));
	jdff dff_A_aLQqy7yi0_2(.dout(w_dff_A_PPwvwhUc5_2),.din(w_dff_A_aLQqy7yi0_2),.clk(gclk));
	jdff dff_A_fbDVu2WR5_2(.dout(w_dff_A_aLQqy7yi0_2),.din(w_dff_A_fbDVu2WR5_2),.clk(gclk));
	jdff dff_A_UzVHen974_2(.dout(w_dff_A_fbDVu2WR5_2),.din(w_dff_A_UzVHen974_2),.clk(gclk));
	jdff dff_A_wMPb9Ryy0_2(.dout(w_dff_A_UzVHen974_2),.din(w_dff_A_wMPb9Ryy0_2),.clk(gclk));
	jdff dff_A_TA0Xv2M69_2(.dout(w_dff_A_wMPb9Ryy0_2),.din(w_dff_A_TA0Xv2M69_2),.clk(gclk));
	jdff dff_A_0BqAqfk73_2(.dout(w_dff_A_TA0Xv2M69_2),.din(w_dff_A_0BqAqfk73_2),.clk(gclk));
	jdff dff_A_MpiDd9nl5_0(.dout(w_G4089_4[0]),.din(w_dff_A_MpiDd9nl5_0),.clk(gclk));
	jdff dff_A_qdjRQbK42_0(.dout(w_dff_A_MpiDd9nl5_0),.din(w_dff_A_qdjRQbK42_0),.clk(gclk));
	jdff dff_A_DD26uquh0_0(.dout(w_dff_A_qdjRQbK42_0),.din(w_dff_A_DD26uquh0_0),.clk(gclk));
	jdff dff_A_Gdm1Zirz0_0(.dout(w_dff_A_DD26uquh0_0),.din(w_dff_A_Gdm1Zirz0_0),.clk(gclk));
	jdff dff_A_cRnDkwLg0_0(.dout(w_dff_A_Gdm1Zirz0_0),.din(w_dff_A_cRnDkwLg0_0),.clk(gclk));
	jdff dff_A_h01dXzPP6_0(.dout(w_dff_A_cRnDkwLg0_0),.din(w_dff_A_h01dXzPP6_0),.clk(gclk));
	jdff dff_A_toTduXpH7_0(.dout(w_dff_A_h01dXzPP6_0),.din(w_dff_A_toTduXpH7_0),.clk(gclk));
	jdff dff_A_j0LIvh7i8_0(.dout(w_dff_A_toTduXpH7_0),.din(w_dff_A_j0LIvh7i8_0),.clk(gclk));
	jdff dff_A_ukqEtCJK1_0(.dout(w_dff_A_j0LIvh7i8_0),.din(w_dff_A_ukqEtCJK1_0),.clk(gclk));
	jdff dff_A_mqLH5R708_0(.dout(w_dff_A_ukqEtCJK1_0),.din(w_dff_A_mqLH5R708_0),.clk(gclk));
	jdff dff_A_9WNOy34A7_0(.dout(w_dff_A_mqLH5R708_0),.din(w_dff_A_9WNOy34A7_0),.clk(gclk));
	jdff dff_A_ZiFLynTk1_0(.dout(w_dff_A_9WNOy34A7_0),.din(w_dff_A_ZiFLynTk1_0),.clk(gclk));
	jdff dff_A_3Q17h9HF4_0(.dout(w_dff_A_ZiFLynTk1_0),.din(w_dff_A_3Q17h9HF4_0),.clk(gclk));
	jdff dff_A_u5e2CJke9_2(.dout(w_G4089_4[2]),.din(w_dff_A_u5e2CJke9_2),.clk(gclk));
	jdff dff_A_VXp3BJCA6_2(.dout(w_dff_A_u5e2CJke9_2),.din(w_dff_A_VXp3BJCA6_2),.clk(gclk));
	jdff dff_A_6ZMsb2EU6_2(.dout(w_dff_A_VXp3BJCA6_2),.din(w_dff_A_6ZMsb2EU6_2),.clk(gclk));
	jdff dff_A_a0PoRZX68_2(.dout(w_dff_A_6ZMsb2EU6_2),.din(w_dff_A_a0PoRZX68_2),.clk(gclk));
	jdff dff_A_6gUPEj5n4_2(.dout(w_dff_A_a0PoRZX68_2),.din(w_dff_A_6gUPEj5n4_2),.clk(gclk));
	jdff dff_A_J32Kr23S0_2(.dout(w_dff_A_6gUPEj5n4_2),.din(w_dff_A_J32Kr23S0_2),.clk(gclk));
	jdff dff_A_x8InVjLI7_2(.dout(w_dff_A_J32Kr23S0_2),.din(w_dff_A_x8InVjLI7_2),.clk(gclk));
	jdff dff_A_5u2vZdMK1_2(.dout(w_dff_A_x8InVjLI7_2),.din(w_dff_A_5u2vZdMK1_2),.clk(gclk));
	jdff dff_A_1VsaclCc0_2(.dout(w_dff_A_5u2vZdMK1_2),.din(w_dff_A_1VsaclCc0_2),.clk(gclk));
	jdff dff_A_EgZuTeVk5_2(.dout(w_dff_A_1VsaclCc0_2),.din(w_dff_A_EgZuTeVk5_2),.clk(gclk));
	jdff dff_A_kBEpjhWt0_2(.dout(w_dff_A_EgZuTeVk5_2),.din(w_dff_A_kBEpjhWt0_2),.clk(gclk));
	jdff dff_A_KC6qS1y01_2(.dout(w_dff_A_kBEpjhWt0_2),.din(w_dff_A_KC6qS1y01_2),.clk(gclk));
	jdff dff_B_I5TLcTiR9_0(.din(n1341),.dout(w_dff_B_I5TLcTiR9_0),.clk(gclk));
	jdff dff_B_6fTDir3V2_0(.din(w_dff_B_I5TLcTiR9_0),.dout(w_dff_B_6fTDir3V2_0),.clk(gclk));
	jdff dff_B_Jwz1yg6a4_0(.din(w_dff_B_6fTDir3V2_0),.dout(w_dff_B_Jwz1yg6a4_0),.clk(gclk));
	jdff dff_B_QHHtFVdr8_0(.din(w_dff_B_Jwz1yg6a4_0),.dout(w_dff_B_QHHtFVdr8_0),.clk(gclk));
	jdff dff_B_u2amd3L69_0(.din(w_dff_B_QHHtFVdr8_0),.dout(w_dff_B_u2amd3L69_0),.clk(gclk));
	jdff dff_B_QP1psu2c3_0(.din(w_dff_B_u2amd3L69_0),.dout(w_dff_B_QP1psu2c3_0),.clk(gclk));
	jdff dff_B_PrVnu9W26_0(.din(w_dff_B_QP1psu2c3_0),.dout(w_dff_B_PrVnu9W26_0),.clk(gclk));
	jdff dff_B_RLgeHdSq9_0(.din(w_dff_B_PrVnu9W26_0),.dout(w_dff_B_RLgeHdSq9_0),.clk(gclk));
	jdff dff_B_3Pk5V8qq8_0(.din(w_dff_B_RLgeHdSq9_0),.dout(w_dff_B_3Pk5V8qq8_0),.clk(gclk));
	jdff dff_B_YrQQ7jc00_0(.din(w_dff_B_3Pk5V8qq8_0),.dout(w_dff_B_YrQQ7jc00_0),.clk(gclk));
	jdff dff_B_3iFp6ebg9_0(.din(w_dff_B_YrQQ7jc00_0),.dout(w_dff_B_3iFp6ebg9_0),.clk(gclk));
	jdff dff_B_mzHjuo2t5_0(.din(w_dff_B_3iFp6ebg9_0),.dout(w_dff_B_mzHjuo2t5_0),.clk(gclk));
	jdff dff_B_hnIG4mRO0_0(.din(w_dff_B_mzHjuo2t5_0),.dout(w_dff_B_hnIG4mRO0_0),.clk(gclk));
	jdff dff_B_qyRUhJ1b1_0(.din(w_dff_B_hnIG4mRO0_0),.dout(w_dff_B_qyRUhJ1b1_0),.clk(gclk));
	jdff dff_B_y8RlDIqL2_0(.din(n1340),.dout(w_dff_B_y8RlDIqL2_0),.clk(gclk));
	jdff dff_B_pFa5jgYj1_1(.din(n1335),.dout(w_dff_B_pFa5jgYj1_1),.clk(gclk));
	jdff dff_B_Wz45cKCp9_1(.din(w_dff_B_pFa5jgYj1_1),.dout(w_dff_B_Wz45cKCp9_1),.clk(gclk));
	jdff dff_B_TvoVTqyh9_1(.din(w_dff_B_Wz45cKCp9_1),.dout(w_dff_B_TvoVTqyh9_1),.clk(gclk));
	jdff dff_A_UMCHUZ8v0_0(.dout(w_n999_2[0]),.din(w_dff_A_UMCHUZ8v0_0),.clk(gclk));
	jdff dff_A_Pizrzpdm6_0(.dout(w_dff_A_UMCHUZ8v0_0),.din(w_dff_A_Pizrzpdm6_0),.clk(gclk));
	jdff dff_A_jmdxMLRo3_0(.dout(w_dff_A_Pizrzpdm6_0),.din(w_dff_A_jmdxMLRo3_0),.clk(gclk));
	jdff dff_A_w5yFxTCv2_0(.dout(w_dff_A_jmdxMLRo3_0),.din(w_dff_A_w5yFxTCv2_0),.clk(gclk));
	jdff dff_A_Nfz1J6KG2_1(.dout(w_n999_2[1]),.din(w_dff_A_Nfz1J6KG2_1),.clk(gclk));
	jdff dff_A_0sNIWVYG8_0(.dout(w_G1689_3[0]),.din(w_dff_A_0sNIWVYG8_0),.clk(gclk));
	jdff dff_A_rYzoHzx23_0(.dout(w_dff_A_0sNIWVYG8_0),.din(w_dff_A_rYzoHzx23_0),.clk(gclk));
	jdff dff_A_DN4yzRBO6_0(.dout(w_dff_A_rYzoHzx23_0),.din(w_dff_A_DN4yzRBO6_0),.clk(gclk));
	jdff dff_A_ub3jo0QX4_0(.dout(w_dff_A_DN4yzRBO6_0),.din(w_dff_A_ub3jo0QX4_0),.clk(gclk));
	jdff dff_A_wIeQAxNX2_1(.dout(w_G1689_3[1]),.din(w_dff_A_wIeQAxNX2_1),.clk(gclk));
	jdff dff_A_9otecso84_1(.dout(w_dff_A_wIeQAxNX2_1),.din(w_dff_A_9otecso84_1),.clk(gclk));
	jdff dff_A_Z3m41yRD3_1(.dout(w_dff_A_9otecso84_1),.din(w_dff_A_Z3m41yRD3_1),.clk(gclk));
	jdff dff_A_S2j9JxC38_0(.dout(w_G137_6[0]),.din(w_dff_A_S2j9JxC38_0),.clk(gclk));
	jdff dff_A_P2Xr5Aeo9_0(.dout(w_dff_A_S2j9JxC38_0),.din(w_dff_A_P2Xr5Aeo9_0),.clk(gclk));
	jdff dff_A_6gFxThkW6_0(.dout(w_dff_A_P2Xr5Aeo9_0),.din(w_dff_A_6gFxThkW6_0),.clk(gclk));
	jdff dff_A_rdQSBNhP1_0(.dout(w_dff_A_6gFxThkW6_0),.din(w_dff_A_rdQSBNhP1_0),.clk(gclk));
	jdff dff_A_ZlA3nojh2_1(.dout(w_G137_6[1]),.din(w_dff_A_ZlA3nojh2_1),.clk(gclk));
	jdff dff_B_5LUGeVFv0_0(.din(n1350),.dout(w_dff_B_5LUGeVFv0_0),.clk(gclk));
	jdff dff_B_R5y6A9X89_0(.din(w_dff_B_5LUGeVFv0_0),.dout(w_dff_B_R5y6A9X89_0),.clk(gclk));
	jdff dff_B_kF0Wv8Js3_0(.din(w_dff_B_R5y6A9X89_0),.dout(w_dff_B_kF0Wv8Js3_0),.clk(gclk));
	jdff dff_B_NCBxH3Uw1_0(.din(w_dff_B_kF0Wv8Js3_0),.dout(w_dff_B_NCBxH3Uw1_0),.clk(gclk));
	jdff dff_B_BF6TFLkP3_0(.din(w_dff_B_NCBxH3Uw1_0),.dout(w_dff_B_BF6TFLkP3_0),.clk(gclk));
	jdff dff_B_Mrz1JR5b7_0(.din(w_dff_B_BF6TFLkP3_0),.dout(w_dff_B_Mrz1JR5b7_0),.clk(gclk));
	jdff dff_B_AVqrgRJA5_0(.din(w_dff_B_Mrz1JR5b7_0),.dout(w_dff_B_AVqrgRJA5_0),.clk(gclk));
	jdff dff_B_qf99JQde5_0(.din(w_dff_B_AVqrgRJA5_0),.dout(w_dff_B_qf99JQde5_0),.clk(gclk));
	jdff dff_B_9GZWId6o1_0(.din(w_dff_B_qf99JQde5_0),.dout(w_dff_B_9GZWId6o1_0),.clk(gclk));
	jdff dff_B_57bqmZdz0_0(.din(w_dff_B_9GZWId6o1_0),.dout(w_dff_B_57bqmZdz0_0),.clk(gclk));
	jdff dff_B_8HX3QIPU8_0(.din(w_dff_B_57bqmZdz0_0),.dout(w_dff_B_8HX3QIPU8_0),.clk(gclk));
	jdff dff_B_ZNHaclVH4_0(.din(w_dff_B_8HX3QIPU8_0),.dout(w_dff_B_ZNHaclVH4_0),.clk(gclk));
	jdff dff_B_CvCeRqJO4_0(.din(n1349),.dout(w_dff_B_CvCeRqJO4_0),.clk(gclk));
	jdff dff_B_cc0SnLEB2_0(.din(n1346),.dout(w_dff_B_cc0SnLEB2_0),.clk(gclk));
	jdff dff_B_0GoxrDj70_1(.din(n1355),.dout(w_dff_B_0GoxrDj70_1),.clk(gclk));
	jdff dff_B_4r1oWU3g5_1(.din(w_dff_B_0GoxrDj70_1),.dout(w_dff_B_4r1oWU3g5_1),.clk(gclk));
	jdff dff_B_eHmNBG1g9_1(.din(w_dff_B_4r1oWU3g5_1),.dout(w_dff_B_eHmNBG1g9_1),.clk(gclk));
	jdff dff_B_YW2B18rA1_1(.din(w_dff_B_eHmNBG1g9_1),.dout(w_dff_B_YW2B18rA1_1),.clk(gclk));
	jdff dff_B_kVckMQ4n5_1(.din(w_dff_B_YW2B18rA1_1),.dout(w_dff_B_kVckMQ4n5_1),.clk(gclk));
	jdff dff_B_vaRZSY4B9_1(.din(w_dff_B_kVckMQ4n5_1),.dout(w_dff_B_vaRZSY4B9_1),.clk(gclk));
	jdff dff_B_tp1CVz8i4_1(.din(w_dff_B_vaRZSY4B9_1),.dout(w_dff_B_tp1CVz8i4_1),.clk(gclk));
	jdff dff_B_QJQuMFGs9_1(.din(w_dff_B_tp1CVz8i4_1),.dout(w_dff_B_QJQuMFGs9_1),.clk(gclk));
	jdff dff_B_4LTrpdAO9_1(.din(w_dff_B_QJQuMFGs9_1),.dout(w_dff_B_4LTrpdAO9_1),.clk(gclk));
	jdff dff_B_OElp9HZj9_1(.din(w_dff_B_4LTrpdAO9_1),.dout(w_dff_B_OElp9HZj9_1),.clk(gclk));
	jdff dff_B_a1wItpK42_1(.din(w_dff_B_OElp9HZj9_1),.dout(w_dff_B_a1wItpK42_1),.clk(gclk));
	jdff dff_B_85cD58965_1(.din(w_dff_B_a1wItpK42_1),.dout(w_dff_B_85cD58965_1),.clk(gclk));
	jdff dff_B_DDK25lXU2_1(.din(w_dff_B_85cD58965_1),.dout(w_dff_B_DDK25lXU2_1),.clk(gclk));
	jdff dff_B_UIxyaktK2_1(.din(w_dff_B_DDK25lXU2_1),.dout(w_dff_B_UIxyaktK2_1),.clk(gclk));
	jdff dff_B_Sxo3aIoO6_1(.din(n1356),.dout(w_dff_B_Sxo3aIoO6_1),.clk(gclk));
	jdff dff_B_8BAIfOQ66_1(.din(w_dff_B_Sxo3aIoO6_1),.dout(w_dff_B_8BAIfOQ66_1),.clk(gclk));
	jdff dff_A_eu48OquP3_0(.dout(w_n993_2[0]),.din(w_dff_A_eu48OquP3_0),.clk(gclk));
	jdff dff_A_t4Fis4ED6_2(.dout(w_n993_2[2]),.din(w_dff_A_t4Fis4ED6_2),.clk(gclk));
	jdff dff_B_pLg1x5Uh2_0(.din(n1354),.dout(w_dff_B_pLg1x5Uh2_0),.clk(gclk));
	jdff dff_B_6Q7NCzT81_1(.din(n1364),.dout(w_dff_B_6Q7NCzT81_1),.clk(gclk));
	jdff dff_B_rmn2sUrR2_1(.din(w_dff_B_6Q7NCzT81_1),.dout(w_dff_B_rmn2sUrR2_1),.clk(gclk));
	jdff dff_B_iR3KjVcr2_1(.din(w_dff_B_rmn2sUrR2_1),.dout(w_dff_B_iR3KjVcr2_1),.clk(gclk));
	jdff dff_B_mp5hQn448_1(.din(w_dff_B_iR3KjVcr2_1),.dout(w_dff_B_mp5hQn448_1),.clk(gclk));
	jdff dff_B_d8NuR7cB6_1(.din(w_dff_B_mp5hQn448_1),.dout(w_dff_B_d8NuR7cB6_1),.clk(gclk));
	jdff dff_B_RGYJOLm64_1(.din(w_dff_B_d8NuR7cB6_1),.dout(w_dff_B_RGYJOLm64_1),.clk(gclk));
	jdff dff_B_keGQCtis8_1(.din(w_dff_B_RGYJOLm64_1),.dout(w_dff_B_keGQCtis8_1),.clk(gclk));
	jdff dff_B_mOX6zrRQ9_1(.din(w_dff_B_keGQCtis8_1),.dout(w_dff_B_mOX6zrRQ9_1),.clk(gclk));
	jdff dff_B_RlCYQF7t8_1(.din(w_dff_B_mOX6zrRQ9_1),.dout(w_dff_B_RlCYQF7t8_1),.clk(gclk));
	jdff dff_B_3V60uW6S5_1(.din(w_dff_B_RlCYQF7t8_1),.dout(w_dff_B_3V60uW6S5_1),.clk(gclk));
	jdff dff_B_cF2rsD8Y6_1(.din(w_dff_B_3V60uW6S5_1),.dout(w_dff_B_cF2rsD8Y6_1),.clk(gclk));
	jdff dff_B_XlM9oqnq7_1(.din(w_dff_B_cF2rsD8Y6_1),.dout(w_dff_B_XlM9oqnq7_1),.clk(gclk));
	jdff dff_B_imWam3ti3_1(.din(w_dff_B_XlM9oqnq7_1),.dout(w_dff_B_imWam3ti3_1),.clk(gclk));
	jdff dff_B_ISUm5JJD8_1(.din(w_dff_B_imWam3ti3_1),.dout(w_dff_B_ISUm5JJD8_1),.clk(gclk));
	jdff dff_B_lX5igOiU7_1(.din(n1365),.dout(w_dff_B_lX5igOiU7_1),.clk(gclk));
	jdff dff_B_zlpaa5gV7_1(.din(w_dff_B_lX5igOiU7_1),.dout(w_dff_B_zlpaa5gV7_1),.clk(gclk));
	jdff dff_A_dbL7HgUb5_0(.dout(w_G1689_2[0]),.din(w_dff_A_dbL7HgUb5_0),.clk(gclk));
	jdff dff_A_5gv99wKp5_1(.dout(w_G1689_2[1]),.din(w_dff_A_5gv99wKp5_1),.clk(gclk));
	jdff dff_A_Fj9jsS5V1_0(.dout(w_n999_1[0]),.din(w_dff_A_Fj9jsS5V1_0),.clk(gclk));
	jdff dff_A_JrqsoFpp4_0(.dout(w_dff_A_Fj9jsS5V1_0),.din(w_dff_A_JrqsoFpp4_0),.clk(gclk));
	jdff dff_A_zlOU3PFR9_0(.dout(w_dff_A_JrqsoFpp4_0),.din(w_dff_A_zlOU3PFR9_0),.clk(gclk));
	jdff dff_A_YtguDoaI5_0(.dout(w_dff_A_zlOU3PFR9_0),.din(w_dff_A_YtguDoaI5_0),.clk(gclk));
	jdff dff_A_Pb6fzhMu8_1(.dout(w_n999_1[1]),.din(w_dff_A_Pb6fzhMu8_1),.clk(gclk));
	jdff dff_A_SnaBn54J6_1(.dout(w_dff_A_Pb6fzhMu8_1),.din(w_dff_A_SnaBn54J6_1),.clk(gclk));
	jdff dff_A_ytPiS0pz5_1(.dout(w_dff_A_SnaBn54J6_1),.din(w_dff_A_ytPiS0pz5_1),.clk(gclk));
	jdff dff_A_OSrG8lVv8_1(.dout(w_dff_A_ytPiS0pz5_1),.din(w_dff_A_OSrG8lVv8_1),.clk(gclk));
	jdff dff_A_KkYYGaHB2_0(.dout(w_n999_0[0]),.din(w_dff_A_KkYYGaHB2_0),.clk(gclk));
	jdff dff_A_lAfnskW83_0(.dout(w_dff_A_KkYYGaHB2_0),.din(w_dff_A_lAfnskW83_0),.clk(gclk));
	jdff dff_A_SAJoHOUv1_0(.dout(w_dff_A_lAfnskW83_0),.din(w_dff_A_SAJoHOUv1_0),.clk(gclk));
	jdff dff_A_fjTSXSRj5_0(.dout(w_dff_A_SAJoHOUv1_0),.din(w_dff_A_fjTSXSRj5_0),.clk(gclk));
	jdff dff_A_nJlTbF2Y5_0(.dout(w_dff_A_fjTSXSRj5_0),.din(w_dff_A_nJlTbF2Y5_0),.clk(gclk));
	jdff dff_A_0wWwtRaZ5_1(.dout(w_n999_0[1]),.din(w_dff_A_0wWwtRaZ5_1),.clk(gclk));
	jdff dff_A_pVYye2o71_1(.dout(w_dff_A_0wWwtRaZ5_1),.din(w_dff_A_pVYye2o71_1),.clk(gclk));
	jdff dff_A_R3I00uET6_1(.dout(w_dff_A_pVYye2o71_1),.din(w_dff_A_R3I00uET6_1),.clk(gclk));
	jdff dff_A_jDTP8mhR3_1(.dout(w_dff_A_R3I00uET6_1),.din(w_dff_A_jDTP8mhR3_1),.clk(gclk));
	jdff dff_B_RJjV95fk3_3(.din(n999),.dout(w_dff_B_RJjV95fk3_3),.clk(gclk));
	jdff dff_B_YB1lEoVq0_3(.din(w_dff_B_RJjV95fk3_3),.dout(w_dff_B_YB1lEoVq0_3),.clk(gclk));
	jdff dff_B_vWiWSM1t5_3(.din(w_dff_B_YB1lEoVq0_3),.dout(w_dff_B_vWiWSM1t5_3),.clk(gclk));
	jdff dff_B_Y3drOONr1_3(.din(w_dff_B_vWiWSM1t5_3),.dout(w_dff_B_Y3drOONr1_3),.clk(gclk));
	jdff dff_B_LH9e32Fv6_3(.din(w_dff_B_Y3drOONr1_3),.dout(w_dff_B_LH9e32Fv6_3),.clk(gclk));
	jdff dff_B_YUHuGYOJ2_3(.din(w_dff_B_LH9e32Fv6_3),.dout(w_dff_B_YUHuGYOJ2_3),.clk(gclk));
	jdff dff_B_3wmX0kaV8_0(.din(n1363),.dout(w_dff_B_3wmX0kaV8_0),.clk(gclk));
	jdff dff_A_fPXvYNu72_0(.dout(w_G137_5[0]),.din(w_dff_A_fPXvYNu72_0),.clk(gclk));
	jdff dff_A_nbfowXPv7_0(.dout(w_dff_A_fPXvYNu72_0),.din(w_dff_A_nbfowXPv7_0),.clk(gclk));
	jdff dff_A_dQQ7lR6d4_1(.dout(w_G137_5[1]),.din(w_dff_A_dQQ7lR6d4_1),.clk(gclk));
	jdff dff_A_Gr1OsUZM4_1(.dout(w_dff_A_dQQ7lR6d4_1),.din(w_dff_A_Gr1OsUZM4_1),.clk(gclk));
	jdff dff_B_SYDnRnlS3_0(.din(n1377),.dout(w_dff_B_SYDnRnlS3_0),.clk(gclk));
	jdff dff_B_uOa2Om2A3_0(.din(w_dff_B_SYDnRnlS3_0),.dout(w_dff_B_uOa2Om2A3_0),.clk(gclk));
	jdff dff_B_KhXMwgVZ5_0(.din(w_dff_B_uOa2Om2A3_0),.dout(w_dff_B_KhXMwgVZ5_0),.clk(gclk));
	jdff dff_B_qRoGwaHe0_0(.din(w_dff_B_KhXMwgVZ5_0),.dout(w_dff_B_qRoGwaHe0_0),.clk(gclk));
	jdff dff_B_Sdsdwj048_0(.din(w_dff_B_qRoGwaHe0_0),.dout(w_dff_B_Sdsdwj048_0),.clk(gclk));
	jdff dff_B_2p7wOymw9_0(.din(w_dff_B_Sdsdwj048_0),.dout(w_dff_B_2p7wOymw9_0),.clk(gclk));
	jdff dff_B_Axfwu7PD6_0(.din(w_dff_B_2p7wOymw9_0),.dout(w_dff_B_Axfwu7PD6_0),.clk(gclk));
	jdff dff_B_IqrRWfvF6_0(.din(w_dff_B_Axfwu7PD6_0),.dout(w_dff_B_IqrRWfvF6_0),.clk(gclk));
	jdff dff_B_aWplygT04_0(.din(w_dff_B_IqrRWfvF6_0),.dout(w_dff_B_aWplygT04_0),.clk(gclk));
	jdff dff_B_D0x8W2UY0_0(.din(w_dff_B_aWplygT04_0),.dout(w_dff_B_D0x8W2UY0_0),.clk(gclk));
	jdff dff_B_L8RbnZAH0_0(.din(w_dff_B_D0x8W2UY0_0),.dout(w_dff_B_L8RbnZAH0_0),.clk(gclk));
	jdff dff_B_z56sPEOa1_0(.din(w_dff_B_L8RbnZAH0_0),.dout(w_dff_B_z56sPEOa1_0),.clk(gclk));
	jdff dff_B_OfaiaSDA2_0(.din(w_dff_B_z56sPEOa1_0),.dout(w_dff_B_OfaiaSDA2_0),.clk(gclk));
	jdff dff_B_DhhOIGEd6_0(.din(w_dff_B_OfaiaSDA2_0),.dout(w_dff_B_DhhOIGEd6_0),.clk(gclk));
	jdff dff_B_HmpjpagX4_0(.din(n1376),.dout(w_dff_B_HmpjpagX4_0),.clk(gclk));
	jdff dff_B_kl9TYwy45_2(.din(G173),.dout(w_dff_B_kl9TYwy45_2),.clk(gclk));
	jdff dff_B_9JfofeCC7_2(.din(G203),.dout(w_dff_B_9JfofeCC7_2),.clk(gclk));
	jdff dff_B_a6wgwdlZ7_2(.din(w_dff_B_9JfofeCC7_2),.dout(w_dff_B_a6wgwdlZ7_2),.clk(gclk));
	jdff dff_B_3OT5K5BX1_1(.din(n1371),.dout(w_dff_B_3OT5K5BX1_1),.clk(gclk));
	jdff dff_B_FUvMHAoG8_1(.din(w_dff_B_3OT5K5BX1_1),.dout(w_dff_B_FUvMHAoG8_1),.clk(gclk));
	jdff dff_B_Maw3qAoo6_1(.din(w_dff_B_FUvMHAoG8_1),.dout(w_dff_B_Maw3qAoo6_1),.clk(gclk));
	jdff dff_B_ZixKtjTy0_1(.din(n1254),.dout(w_dff_B_ZixKtjTy0_1),.clk(gclk));
	jdff dff_B_omGMbmO87_1(.din(w_dff_B_ZixKtjTy0_1),.dout(w_dff_B_omGMbmO87_1),.clk(gclk));
	jdff dff_B_Sb5K7Lkr7_1(.din(w_dff_B_omGMbmO87_1),.dout(w_dff_B_Sb5K7Lkr7_1),.clk(gclk));
	jdff dff_B_cXYwp4QC8_1(.din(w_dff_B_Sb5K7Lkr7_1),.dout(w_dff_B_cXYwp4QC8_1),.clk(gclk));
	jdff dff_B_MhK4R2VP5_1(.din(w_dff_B_cXYwp4QC8_1),.dout(w_dff_B_MhK4R2VP5_1),.clk(gclk));
	jdff dff_B_lnV2xwj59_1(.din(w_dff_B_MhK4R2VP5_1),.dout(w_dff_B_lnV2xwj59_1),.clk(gclk));
	jdff dff_B_JTVD6QjC1_1(.din(w_dff_B_lnV2xwj59_1),.dout(w_dff_B_JTVD6QjC1_1),.clk(gclk));
	jdff dff_B_0dqQCNPE0_1(.din(w_dff_B_JTVD6QjC1_1),.dout(w_dff_B_0dqQCNPE0_1),.clk(gclk));
	jdff dff_B_3KgK7ttF1_1(.din(w_dff_B_0dqQCNPE0_1),.dout(w_dff_B_3KgK7ttF1_1),.clk(gclk));
	jdff dff_B_FUlOgvlE4_0(.din(n1257),.dout(w_dff_B_FUlOgvlE4_0),.clk(gclk));
	jdff dff_B_sXdgtlN89_0(.din(w_dff_B_FUlOgvlE4_0),.dout(w_dff_B_sXdgtlN89_0),.clk(gclk));
	jdff dff_B_IzmcUFDw6_0(.din(w_dff_B_sXdgtlN89_0),.dout(w_dff_B_IzmcUFDw6_0),.clk(gclk));
	jdff dff_B_NZvyk9B59_0(.din(w_dff_B_IzmcUFDw6_0),.dout(w_dff_B_NZvyk9B59_0),.clk(gclk));
	jdff dff_B_giUEsZHo8_0(.din(w_dff_B_NZvyk9B59_0),.dout(w_dff_B_giUEsZHo8_0),.clk(gclk));
	jdff dff_B_xbwqmf6Y6_0(.din(w_dff_B_giUEsZHo8_0),.dout(w_dff_B_xbwqmf6Y6_0),.clk(gclk));
	jdff dff_B_LaNUnhTa0_0(.din(w_dff_B_xbwqmf6Y6_0),.dout(w_dff_B_LaNUnhTa0_0),.clk(gclk));
	jdff dff_B_aT3NvJZB9_0(.din(w_dff_B_LaNUnhTa0_0),.dout(w_dff_B_aT3NvJZB9_0),.clk(gclk));
	jdff dff_B_doZsvJYt5_0(.din(w_dff_B_aT3NvJZB9_0),.dout(w_dff_B_doZsvJYt5_0),.clk(gclk));
	jdff dff_B_uRSWtzdc4_1(.din(n500),.dout(w_dff_B_uRSWtzdc4_1),.clk(gclk));
	jdff dff_B_2ghFBc636_1(.din(G113),.dout(w_dff_B_2ghFBc636_1),.clk(gclk));
	jdff dff_B_mQPe3CN02_1(.din(w_dff_B_2ghFBc636_1),.dout(w_dff_B_mQPe3CN02_1),.clk(gclk));
	jdff dff_A_KfgNAJJQ1_0(.dout(w_n1007_2[0]),.din(w_dff_A_KfgNAJJQ1_0),.clk(gclk));
	jdff dff_A_8emau9tp9_0(.dout(w_dff_A_KfgNAJJQ1_0),.din(w_dff_A_8emau9tp9_0),.clk(gclk));
	jdff dff_A_rt8DgwgD2_0(.dout(w_dff_A_8emau9tp9_0),.din(w_dff_A_rt8DgwgD2_0),.clk(gclk));
	jdff dff_A_94cTNurI0_0(.dout(w_dff_A_rt8DgwgD2_0),.din(w_dff_A_94cTNurI0_0),.clk(gclk));
	jdff dff_A_mcsujQa73_1(.dout(w_n1007_2[1]),.din(w_dff_A_mcsujQa73_1),.clk(gclk));
	jdff dff_B_eH6XZ9HE6_1(.din(n1216),.dout(w_dff_B_eH6XZ9HE6_1),.clk(gclk));
	jdff dff_B_99Jp3u7C1_1(.din(w_dff_B_eH6XZ9HE6_1),.dout(w_dff_B_99Jp3u7C1_1),.clk(gclk));
	jdff dff_B_d1vcH2rp8_1(.din(w_dff_B_99Jp3u7C1_1),.dout(w_dff_B_d1vcH2rp8_1),.clk(gclk));
	jdff dff_B_kTa99tev8_1(.din(w_dff_B_d1vcH2rp8_1),.dout(w_dff_B_kTa99tev8_1),.clk(gclk));
	jdff dff_B_tW1fGQ8W6_1(.din(w_dff_B_kTa99tev8_1),.dout(w_dff_B_tW1fGQ8W6_1),.clk(gclk));
	jdff dff_B_bfYeBHZJ5_1(.din(w_dff_B_tW1fGQ8W6_1),.dout(w_dff_B_bfYeBHZJ5_1),.clk(gclk));
	jdff dff_B_tQhKUQkb1_1(.din(w_dff_B_bfYeBHZJ5_1),.dout(w_dff_B_tQhKUQkb1_1),.clk(gclk));
	jdff dff_B_qsP9iLyS2_0(.din(n1219),.dout(w_dff_B_qsP9iLyS2_0),.clk(gclk));
	jdff dff_B_P0VoA2qX3_0(.din(w_dff_B_qsP9iLyS2_0),.dout(w_dff_B_P0VoA2qX3_0),.clk(gclk));
	jdff dff_B_U4764NVg8_0(.din(w_dff_B_P0VoA2qX3_0),.dout(w_dff_B_U4764NVg8_0),.clk(gclk));
	jdff dff_B_X4qyWCUQ9_0(.din(w_dff_B_U4764NVg8_0),.dout(w_dff_B_X4qyWCUQ9_0),.clk(gclk));
	jdff dff_B_BXVMmKux4_0(.din(w_dff_B_X4qyWCUQ9_0),.dout(w_dff_B_BXVMmKux4_0),.clk(gclk));
	jdff dff_B_8miCOP7x2_0(.din(w_dff_B_BXVMmKux4_0),.dout(w_dff_B_8miCOP7x2_0),.clk(gclk));
	jdff dff_B_xnScEtc77_0(.din(w_dff_B_8miCOP7x2_0),.dout(w_dff_B_xnScEtc77_0),.clk(gclk));
	jdff dff_A_GTSqUhit9_1(.dout(w_n989_0[1]),.din(w_dff_A_GTSqUhit9_1),.clk(gclk));
	jdff dff_A_VvpmMaxw4_1(.dout(w_dff_A_GTSqUhit9_1),.din(w_dff_A_VvpmMaxw4_1),.clk(gclk));
	jdff dff_B_XgWeIoQq1_1(.din(n988),.dout(w_dff_B_XgWeIoQq1_1),.clk(gclk));
	jdff dff_B_8itSGbJL9_1(.din(w_dff_B_XgWeIoQq1_1),.dout(w_dff_B_8itSGbJL9_1),.clk(gclk));
	jdff dff_B_zz6sdQL49_1(.din(w_dff_B_8itSGbJL9_1),.dout(w_dff_B_zz6sdQL49_1),.clk(gclk));
	jdff dff_B_9Jufj2dn4_1(.din(G112),.dout(w_dff_B_9Jufj2dn4_1),.clk(gclk));
	jdff dff_B_WdEBxlLx2_1(.din(w_dff_B_9Jufj2dn4_1),.dout(w_dff_B_WdEBxlLx2_1),.clk(gclk));
	jdff dff_A_CsIMUsMA1_0(.dout(w_G1691_3[0]),.din(w_dff_A_CsIMUsMA1_0),.clk(gclk));
	jdff dff_A_YhaeeRwc3_0(.dout(w_dff_A_CsIMUsMA1_0),.din(w_dff_A_YhaeeRwc3_0),.clk(gclk));
	jdff dff_A_fvuRWb520_0(.dout(w_dff_A_YhaeeRwc3_0),.din(w_dff_A_fvuRWb520_0),.clk(gclk));
	jdff dff_A_PoXbhRtG3_0(.dout(w_dff_A_fvuRWb520_0),.din(w_dff_A_PoXbhRtG3_0),.clk(gclk));
	jdff dff_A_OZrfM07g6_1(.dout(w_G1691_3[1]),.din(w_dff_A_OZrfM07g6_1),.clk(gclk));
	jdff dff_A_MVJX8e971_1(.dout(w_dff_A_OZrfM07g6_1),.din(w_dff_A_MVJX8e971_1),.clk(gclk));
	jdff dff_A_jsFtZQH11_1(.dout(w_dff_A_MVJX8e971_1),.din(w_dff_A_jsFtZQH11_1),.clk(gclk));
	jdff dff_B_jRkXEa4G8_1(.din(n1382),.dout(w_dff_B_jRkXEa4G8_1),.clk(gclk));
	jdff dff_B_hIpkgZVf9_1(.din(w_dff_B_jRkXEa4G8_1),.dout(w_dff_B_hIpkgZVf9_1),.clk(gclk));
	jdff dff_B_KprD1YzT0_1(.din(w_dff_B_hIpkgZVf9_1),.dout(w_dff_B_KprD1YzT0_1),.clk(gclk));
	jdff dff_B_LSMEqjdP5_1(.din(w_dff_B_KprD1YzT0_1),.dout(w_dff_B_LSMEqjdP5_1),.clk(gclk));
	jdff dff_B_wyrr0KVs3_1(.din(w_dff_B_LSMEqjdP5_1),.dout(w_dff_B_wyrr0KVs3_1),.clk(gclk));
	jdff dff_B_QmSWv1xo5_1(.din(w_dff_B_wyrr0KVs3_1),.dout(w_dff_B_QmSWv1xo5_1),.clk(gclk));
	jdff dff_B_q2ZlH6GD6_1(.din(w_dff_B_QmSWv1xo5_1),.dout(w_dff_B_q2ZlH6GD6_1),.clk(gclk));
	jdff dff_B_UUnfP5AT5_1(.din(w_dff_B_q2ZlH6GD6_1),.dout(w_dff_B_UUnfP5AT5_1),.clk(gclk));
	jdff dff_B_EvaoAqRi2_1(.din(w_dff_B_UUnfP5AT5_1),.dout(w_dff_B_EvaoAqRi2_1),.clk(gclk));
	jdff dff_B_NKhI9E6Q0_1(.din(w_dff_B_EvaoAqRi2_1),.dout(w_dff_B_NKhI9E6Q0_1),.clk(gclk));
	jdff dff_B_X73lLezi7_1(.din(w_dff_B_NKhI9E6Q0_1),.dout(w_dff_B_X73lLezi7_1),.clk(gclk));
	jdff dff_B_CKPptlEW0_1(.din(w_dff_B_X73lLezi7_1),.dout(w_dff_B_CKPptlEW0_1),.clk(gclk));
	jdff dff_B_Ne8oZc1E3_1(.din(w_dff_B_CKPptlEW0_1),.dout(w_dff_B_Ne8oZc1E3_1),.clk(gclk));
	jdff dff_B_uPXEjoAm5_1(.din(n1383),.dout(w_dff_B_uPXEjoAm5_1),.clk(gclk));
	jdff dff_B_AyFQlIRn2_1(.din(w_dff_B_uPXEjoAm5_1),.dout(w_dff_B_AyFQlIRn2_1),.clk(gclk));
	jdff dff_B_geOM1XqB1_1(.din(n1245),.dout(w_dff_B_geOM1XqB1_1),.clk(gclk));
	jdff dff_B_ilvktEQ82_1(.din(w_dff_B_geOM1XqB1_1),.dout(w_dff_B_ilvktEQ82_1),.clk(gclk));
	jdff dff_B_ueYmJDVK8_1(.din(w_dff_B_ilvktEQ82_1),.dout(w_dff_B_ueYmJDVK8_1),.clk(gclk));
	jdff dff_B_D3cU6MAc4_1(.din(w_dff_B_ueYmJDVK8_1),.dout(w_dff_B_D3cU6MAc4_1),.clk(gclk));
	jdff dff_B_pKtBL8wo0_1(.din(w_dff_B_D3cU6MAc4_1),.dout(w_dff_B_pKtBL8wo0_1),.clk(gclk));
	jdff dff_B_pPEyHNkF5_1(.din(w_dff_B_pKtBL8wo0_1),.dout(w_dff_B_pPEyHNkF5_1),.clk(gclk));
	jdff dff_B_cqMlWShW7_1(.din(w_dff_B_pPEyHNkF5_1),.dout(w_dff_B_cqMlWShW7_1),.clk(gclk));
	jdff dff_B_e7voZlXf7_1(.din(w_dff_B_cqMlWShW7_1),.dout(w_dff_B_e7voZlXf7_1),.clk(gclk));
	jdff dff_B_JLq5iGFx1_1(.din(w_dff_B_e7voZlXf7_1),.dout(w_dff_B_JLq5iGFx1_1),.clk(gclk));
	jdff dff_B_bF1nBn231_1(.din(w_dff_B_JLq5iGFx1_1),.dout(w_dff_B_bF1nBn231_1),.clk(gclk));
	jdff dff_B_8v49LUSi5_1(.din(w_dff_B_bF1nBn231_1),.dout(w_dff_B_8v49LUSi5_1),.clk(gclk));
	jdff dff_B_mVCr4D5P8_1(.din(n1247),.dout(w_dff_B_mVCr4D5P8_1),.clk(gclk));
	jdff dff_B_Muchwt741_1(.din(w_dff_B_mVCr4D5P8_1),.dout(w_dff_B_Muchwt741_1),.clk(gclk));
	jdff dff_B_WsIOQDBW7_1(.din(w_dff_B_Muchwt741_1),.dout(w_dff_B_WsIOQDBW7_1),.clk(gclk));
	jdff dff_B_ZBHpFyMZ4_1(.din(w_dff_B_WsIOQDBW7_1),.dout(w_dff_B_ZBHpFyMZ4_1),.clk(gclk));
	jdff dff_B_8se2icQt3_1(.din(w_dff_B_ZBHpFyMZ4_1),.dout(w_dff_B_8se2icQt3_1),.clk(gclk));
	jdff dff_B_SQcqYZmX4_1(.din(w_dff_B_8se2icQt3_1),.dout(w_dff_B_SQcqYZmX4_1),.clk(gclk));
	jdff dff_B_Cl0PRBtX8_1(.din(w_dff_B_SQcqYZmX4_1),.dout(w_dff_B_Cl0PRBtX8_1),.clk(gclk));
	jdff dff_B_F2YdCrcQ2_1(.din(w_dff_B_Cl0PRBtX8_1),.dout(w_dff_B_F2YdCrcQ2_1),.clk(gclk));
	jdff dff_B_iZbEqrwL4_1(.din(n951),.dout(w_dff_B_iZbEqrwL4_1),.clk(gclk));
	jdff dff_B_L7mduJ635_1(.din(w_dff_B_iZbEqrwL4_1),.dout(w_dff_B_L7mduJ635_1),.clk(gclk));
	jdff dff_B_p8HR99bd4_1(.din(w_dff_B_L7mduJ635_1),.dout(w_dff_B_p8HR99bd4_1),.clk(gclk));
	jdff dff_B_20fjxLOe7_1(.din(w_dff_B_p8HR99bd4_1),.dout(w_dff_B_20fjxLOe7_1),.clk(gclk));
	jdff dff_B_8kpeJ6dk8_1(.din(w_dff_B_20fjxLOe7_1),.dout(w_dff_B_8kpeJ6dk8_1),.clk(gclk));
	jdff dff_B_cUsp9VPF8_1(.din(n513),.dout(w_dff_B_cUsp9VPF8_1),.clk(gclk));
	jdff dff_B_HKwz4r8D7_1(.din(G53),.dout(w_dff_B_HKwz4r8D7_1),.clk(gclk));
	jdff dff_B_fyVm4Obu7_1(.din(w_dff_B_HKwz4r8D7_1),.dout(w_dff_B_fyVm4Obu7_1),.clk(gclk));
	jdff dff_B_Sf6XW2lO0_1(.din(n1207),.dout(w_dff_B_Sf6XW2lO0_1),.clk(gclk));
	jdff dff_B_m6C7XxgQ5_1(.din(w_dff_B_Sf6XW2lO0_1),.dout(w_dff_B_m6C7XxgQ5_1),.clk(gclk));
	jdff dff_B_tSjut3WQ4_1(.din(w_dff_B_m6C7XxgQ5_1),.dout(w_dff_B_tSjut3WQ4_1),.clk(gclk));
	jdff dff_B_GPrc29YB8_1(.din(w_dff_B_tSjut3WQ4_1),.dout(w_dff_B_GPrc29YB8_1),.clk(gclk));
	jdff dff_B_WsOgnKMC5_1(.din(w_dff_B_GPrc29YB8_1),.dout(w_dff_B_WsOgnKMC5_1),.clk(gclk));
	jdff dff_B_qiqA1Udo2_1(.din(w_dff_B_WsOgnKMC5_1),.dout(w_dff_B_qiqA1Udo2_1),.clk(gclk));
	jdff dff_B_73X1Uyel6_1(.din(w_dff_B_qiqA1Udo2_1),.dout(w_dff_B_73X1Uyel6_1),.clk(gclk));
	jdff dff_B_IMkZVaau5_1(.din(w_dff_B_73X1Uyel6_1),.dout(w_dff_B_IMkZVaau5_1),.clk(gclk));
	jdff dff_B_l0lvpBRH7_1(.din(w_dff_B_IMkZVaau5_1),.dout(w_dff_B_l0lvpBRH7_1),.clk(gclk));
	jdff dff_B_GyhXUum03_0(.din(n1211),.dout(w_dff_B_GyhXUum03_0),.clk(gclk));
	jdff dff_B_mgJ7Dxo54_0(.din(w_dff_B_GyhXUum03_0),.dout(w_dff_B_mgJ7Dxo54_0),.clk(gclk));
	jdff dff_B_4JmHfGlC0_0(.din(w_dff_B_mgJ7Dxo54_0),.dout(w_dff_B_4JmHfGlC0_0),.clk(gclk));
	jdff dff_B_prtKVrCG4_0(.din(w_dff_B_4JmHfGlC0_0),.dout(w_dff_B_prtKVrCG4_0),.clk(gclk));
	jdff dff_B_uCDM9g1o6_0(.din(w_dff_B_prtKVrCG4_0),.dout(w_dff_B_uCDM9g1o6_0),.clk(gclk));
	jdff dff_B_9LvvXecj4_0(.din(w_dff_B_uCDM9g1o6_0),.dout(w_dff_B_9LvvXecj4_0),.clk(gclk));
	jdff dff_B_7R0hRiq00_1(.din(n978),.dout(w_dff_B_7R0hRiq00_1),.clk(gclk));
	jdff dff_B_WuaJGEol0_1(.din(w_dff_B_7R0hRiq00_1),.dout(w_dff_B_WuaJGEol0_1),.clk(gclk));
	jdff dff_B_oANVJYZs4_1(.din(w_dff_B_WuaJGEol0_1),.dout(w_dff_B_oANVJYZs4_1),.clk(gclk));
	jdff dff_B_DyVAr6xK6_1(.din(w_dff_B_oANVJYZs4_1),.dout(w_dff_B_DyVAr6xK6_1),.clk(gclk));
	jdff dff_B_la9Hy5cp1_1(.din(n982),.dout(w_dff_B_la9Hy5cp1_1),.clk(gclk));
	jdff dff_B_rrZli3ql8_1(.din(n980),.dout(w_dff_B_rrZli3ql8_1),.clk(gclk));
	jdff dff_B_BF6jpSG08_1(.din(w_dff_B_rrZli3ql8_1),.dout(w_dff_B_BF6jpSG08_1),.clk(gclk));
	jdff dff_B_nDHupgS93_1(.din(G116),.dout(w_dff_B_nDHupgS93_1),.clk(gclk));
	jdff dff_B_bxnokhrt3_1(.din(w_dff_B_nDHupgS93_1),.dout(w_dff_B_bxnokhrt3_1),.clk(gclk));
	jdff dff_B_rEPQrDHN1_0(.din(n1381),.dout(w_dff_B_rEPQrDHN1_0),.clk(gclk));
	jdff dff_B_xzRqBeyM5_2(.din(G167),.dout(w_dff_B_xzRqBeyM5_2),.clk(gclk));
	jdff dff_B_2NcDcZ4t1_2(.din(G197),.dout(w_dff_B_2NcDcZ4t1_2),.clk(gclk));
	jdff dff_B_LbQbXpqE0_2(.din(w_dff_B_2NcDcZ4t1_2),.dout(w_dff_B_LbQbXpqE0_2),.clk(gclk));
	jdff dff_B_G0TdlR5Q6_0(.din(n1395),.dout(w_dff_B_G0TdlR5Q6_0),.clk(gclk));
	jdff dff_B_ulbvS3w21_0(.din(w_dff_B_G0TdlR5Q6_0),.dout(w_dff_B_ulbvS3w21_0),.clk(gclk));
	jdff dff_B_rxCsvLWZ1_0(.din(w_dff_B_ulbvS3w21_0),.dout(w_dff_B_rxCsvLWZ1_0),.clk(gclk));
	jdff dff_B_xb12rojj6_0(.din(w_dff_B_rxCsvLWZ1_0),.dout(w_dff_B_xb12rojj6_0),.clk(gclk));
	jdff dff_B_p7XqTf1S1_0(.din(w_dff_B_xb12rojj6_0),.dout(w_dff_B_p7XqTf1S1_0),.clk(gclk));
	jdff dff_B_7E62Ck327_0(.din(w_dff_B_p7XqTf1S1_0),.dout(w_dff_B_7E62Ck327_0),.clk(gclk));
	jdff dff_B_uYJPnmsC3_0(.din(w_dff_B_7E62Ck327_0),.dout(w_dff_B_uYJPnmsC3_0),.clk(gclk));
	jdff dff_B_6FbSOT536_0(.din(w_dff_B_uYJPnmsC3_0),.dout(w_dff_B_6FbSOT536_0),.clk(gclk));
	jdff dff_B_OXbUoqo60_0(.din(w_dff_B_6FbSOT536_0),.dout(w_dff_B_OXbUoqo60_0),.clk(gclk));
	jdff dff_B_upJEYTwM5_0(.din(w_dff_B_OXbUoqo60_0),.dout(w_dff_B_upJEYTwM5_0),.clk(gclk));
	jdff dff_B_U7QwuuLY5_0(.din(w_dff_B_upJEYTwM5_0),.dout(w_dff_B_U7QwuuLY5_0),.clk(gclk));
	jdff dff_B_IEVt0auh7_0(.din(w_dff_B_U7QwuuLY5_0),.dout(w_dff_B_IEVt0auh7_0),.clk(gclk));
	jdff dff_B_eG8Y03wf1_0(.din(w_dff_B_IEVt0auh7_0),.dout(w_dff_B_eG8Y03wf1_0),.clk(gclk));
	jdff dff_B_z6GN4o6J4_0(.din(w_dff_B_eG8Y03wf1_0),.dout(w_dff_B_z6GN4o6J4_0),.clk(gclk));
	jdff dff_B_bTO4pNdS5_0(.din(n1394),.dout(w_dff_B_bTO4pNdS5_0),.clk(gclk));
	jdff dff_B_Z4HedfuY6_2(.din(G164),.dout(w_dff_B_Z4HedfuY6_2),.clk(gclk));
	jdff dff_B_QCywYnxs3_2(.din(G194),.dout(w_dff_B_QCywYnxs3_2),.clk(gclk));
	jdff dff_B_0c6JP3fR4_2(.din(w_dff_B_QCywYnxs3_2),.dout(w_dff_B_0c6JP3fR4_2),.clk(gclk));
	jdff dff_B_Z3R43VgP3_1(.din(n1389),.dout(w_dff_B_Z3R43VgP3_1),.clk(gclk));
	jdff dff_B_qT4UQQcZ1_1(.din(w_dff_B_Z3R43VgP3_1),.dout(w_dff_B_qT4UQQcZ1_1),.clk(gclk));
	jdff dff_B_5vZSiFMv0_1(.din(w_dff_B_qT4UQQcZ1_1),.dout(w_dff_B_5vZSiFMv0_1),.clk(gclk));
	jdff dff_B_EKRjpc7W1_1(.din(n1239),.dout(w_dff_B_EKRjpc7W1_1),.clk(gclk));
	jdff dff_B_ZT7uiZGu0_1(.din(w_dff_B_EKRjpc7W1_1),.dout(w_dff_B_ZT7uiZGu0_1),.clk(gclk));
	jdff dff_B_JpGydxwo8_1(.din(w_dff_B_ZT7uiZGu0_1),.dout(w_dff_B_JpGydxwo8_1),.clk(gclk));
	jdff dff_B_Xp0iKvHv0_1(.din(w_dff_B_JpGydxwo8_1),.dout(w_dff_B_Xp0iKvHv0_1),.clk(gclk));
	jdff dff_B_pGwEHb6S2_1(.din(w_dff_B_Xp0iKvHv0_1),.dout(w_dff_B_pGwEHb6S2_1),.clk(gclk));
	jdff dff_B_dQ7mUAgC6_1(.din(w_dff_B_pGwEHb6S2_1),.dout(w_dff_B_dQ7mUAgC6_1),.clk(gclk));
	jdff dff_B_svvvIDDB7_1(.din(w_dff_B_dQ7mUAgC6_1),.dout(w_dff_B_svvvIDDB7_1),.clk(gclk));
	jdff dff_B_loHEoTp43_1(.din(w_dff_B_svvvIDDB7_1),.dout(w_dff_B_loHEoTp43_1),.clk(gclk));
	jdff dff_B_8k09gzto0_1(.din(w_dff_B_loHEoTp43_1),.dout(w_dff_B_8k09gzto0_1),.clk(gclk));
	jdff dff_B_GPvXg0MZ2_0(.din(n1242),.dout(w_dff_B_GPvXg0MZ2_0),.clk(gclk));
	jdff dff_B_wLqZL7Tu7_0(.din(w_dff_B_GPvXg0MZ2_0),.dout(w_dff_B_wLqZL7Tu7_0),.clk(gclk));
	jdff dff_B_QwjycpWc7_0(.din(w_dff_B_wLqZL7Tu7_0),.dout(w_dff_B_QwjycpWc7_0),.clk(gclk));
	jdff dff_B_i2kKjPjL7_0(.din(w_dff_B_QwjycpWc7_0),.dout(w_dff_B_i2kKjPjL7_0),.clk(gclk));
	jdff dff_B_3vRC0caK2_0(.din(w_dff_B_i2kKjPjL7_0),.dout(w_dff_B_3vRC0caK2_0),.clk(gclk));
	jdff dff_B_KUmo848l3_0(.din(w_dff_B_3vRC0caK2_0),.dout(w_dff_B_KUmo848l3_0),.clk(gclk));
	jdff dff_B_N1FDV6gt3_0(.din(w_dff_B_KUmo848l3_0),.dout(w_dff_B_N1FDV6gt3_0),.clk(gclk));
	jdff dff_B_1mlDaVVb1_0(.din(w_dff_B_N1FDV6gt3_0),.dout(w_dff_B_1mlDaVVb1_0),.clk(gclk));
	jdff dff_B_EDvBLAjE8_0(.din(w_dff_B_1mlDaVVb1_0),.dout(w_dff_B_EDvBLAjE8_0),.clk(gclk));
	jdff dff_A_aQPlSkov2_1(.dout(w_n459_0[1]),.din(w_dff_A_aQPlSkov2_1),.clk(gclk));
	jdff dff_A_ogj2uxWd9_1(.dout(w_dff_A_aQPlSkov2_1),.din(w_dff_A_ogj2uxWd9_1),.clk(gclk));
	jdff dff_A_2QrO1eFJ5_1(.dout(w_dff_A_ogj2uxWd9_1),.din(w_dff_A_2QrO1eFJ5_1),.clk(gclk));
	jdff dff_B_ls9Jbc5m9_1(.din(n455),.dout(w_dff_B_ls9Jbc5m9_1),.clk(gclk));
	jdff dff_B_dTX8841M8_3(.din(G3548),.dout(w_dff_B_dTX8841M8_3),.clk(gclk));
	jdff dff_A_ayZfTGbW7_0(.dout(w_n749_6[0]),.din(w_dff_A_ayZfTGbW7_0),.clk(gclk));
	jdff dff_A_hKrFVRUb9_0(.dout(w_dff_A_ayZfTGbW7_0),.din(w_dff_A_hKrFVRUb9_0),.clk(gclk));
	jdff dff_A_FRRHhxFu1_0(.dout(w_dff_A_hKrFVRUb9_0),.din(w_dff_A_FRRHhxFu1_0),.clk(gclk));
	jdff dff_A_q1GhjYhb4_0(.dout(w_dff_A_FRRHhxFu1_0),.din(w_dff_A_q1GhjYhb4_0),.clk(gclk));
	jdff dff_A_1iDa6NEo0_0(.dout(w_dff_A_q1GhjYhb4_0),.din(w_dff_A_1iDa6NEo0_0),.clk(gclk));
	jdff dff_A_71HeBFXT1_0(.dout(w_dff_A_1iDa6NEo0_0),.din(w_dff_A_71HeBFXT1_0),.clk(gclk));
	jdff dff_A_mjUWrnhX0_0(.dout(w_dff_A_71HeBFXT1_0),.din(w_dff_A_mjUWrnhX0_0),.clk(gclk));
	jdff dff_A_61pbxiN61_0(.dout(w_dff_A_mjUWrnhX0_0),.din(w_dff_A_61pbxiN61_0),.clk(gclk));
	jdff dff_A_XkHPpHga1_0(.dout(w_dff_A_61pbxiN61_0),.din(w_dff_A_XkHPpHga1_0),.clk(gclk));
	jdff dff_A_heEpW0bd2_1(.dout(w_n949_0[1]),.din(w_dff_A_heEpW0bd2_1),.clk(gclk));
	jdff dff_A_prQ93bQ73_1(.dout(w_dff_A_heEpW0bd2_1),.din(w_dff_A_prQ93bQ73_1),.clk(gclk));
	jdff dff_B_AbTt4sVP2_1(.din(n946),.dout(w_dff_B_AbTt4sVP2_1),.clk(gclk));
	jdff dff_B_STdf4kd25_1(.din(w_dff_B_AbTt4sVP2_1),.dout(w_dff_B_STdf4kd25_1),.clk(gclk));
	jdff dff_B_k9d95q3R6_1(.din(w_dff_B_STdf4kd25_1),.dout(w_dff_B_k9d95q3R6_1),.clk(gclk));
	jdff dff_B_u6wb1a4G8_1(.din(w_dff_B_k9d95q3R6_1),.dout(w_dff_B_u6wb1a4G8_1),.clk(gclk));
	jdff dff_A_5uB1OBD08_0(.dout(w_G4091_2[0]),.din(w_dff_A_5uB1OBD08_0),.clk(gclk));
	jdff dff_A_X20EqEFP2_0(.dout(w_dff_A_5uB1OBD08_0),.din(w_dff_A_X20EqEFP2_0),.clk(gclk));
	jdff dff_A_7210V7iL2_1(.dout(w_G4091_2[1]),.din(w_dff_A_7210V7iL2_1),.clk(gclk));
	jdff dff_A_WX1kDifk3_1(.dout(w_dff_A_7210V7iL2_1),.din(w_dff_A_WX1kDifk3_1),.clk(gclk));
	jdff dff_B_8TlBesEM9_1(.din(G114),.dout(w_dff_B_8TlBesEM9_1),.clk(gclk));
	jdff dff_B_mtf1kKtJ0_1(.din(w_dff_B_8TlBesEM9_1),.dout(w_dff_B_mtf1kKtJ0_1),.clk(gclk));
	jdff dff_A_hmk7Jl116_0(.dout(w_n1008_2[0]),.din(w_dff_A_hmk7Jl116_0),.clk(gclk));
	jdff dff_A_Jdvyeqj88_2(.dout(w_n1008_2[2]),.din(w_dff_A_Jdvyeqj88_2),.clk(gclk));
	jdff dff_B_qbT2jZtg7_1(.din(n1198),.dout(w_dff_B_qbT2jZtg7_1),.clk(gclk));
	jdff dff_B_2mGFCHHN0_1(.din(w_dff_B_qbT2jZtg7_1),.dout(w_dff_B_2mGFCHHN0_1),.clk(gclk));
	jdff dff_B_fYJgsvkO4_1(.din(w_dff_B_2mGFCHHN0_1),.dout(w_dff_B_fYJgsvkO4_1),.clk(gclk));
	jdff dff_B_fQU27Otu8_1(.din(w_dff_B_fYJgsvkO4_1),.dout(w_dff_B_fQU27Otu8_1),.clk(gclk));
	jdff dff_B_fvCy5GTE6_1(.din(w_dff_B_fQU27Otu8_1),.dout(w_dff_B_fvCy5GTE6_1),.clk(gclk));
	jdff dff_B_VkPjJjyO6_1(.din(w_dff_B_fvCy5GTE6_1),.dout(w_dff_B_VkPjJjyO6_1),.clk(gclk));
	jdff dff_B_KOcVQ9zg7_1(.din(w_dff_B_VkPjJjyO6_1),.dout(w_dff_B_KOcVQ9zg7_1),.clk(gclk));
	jdff dff_B_rWjubk8T0_1(.din(w_dff_B_KOcVQ9zg7_1),.dout(w_dff_B_rWjubk8T0_1),.clk(gclk));
	jdff dff_B_klFXr6gf2_1(.din(w_dff_B_rWjubk8T0_1),.dout(w_dff_B_klFXr6gf2_1),.clk(gclk));
	jdff dff_B_sZyG1Hue7_1(.din(w_dff_B_klFXr6gf2_1),.dout(w_dff_B_sZyG1Hue7_1),.clk(gclk));
	jdff dff_B_Zwbz9OBi8_1(.din(n1200),.dout(w_dff_B_Zwbz9OBi8_1),.clk(gclk));
	jdff dff_B_AspQvzbM2_1(.din(w_dff_B_Zwbz9OBi8_1),.dout(w_dff_B_AspQvzbM2_1),.clk(gclk));
	jdff dff_B_Gz3wjFV38_1(.din(w_dff_B_AspQvzbM2_1),.dout(w_dff_B_Gz3wjFV38_1),.clk(gclk));
	jdff dff_B_wOBoi8IA9_1(.din(w_dff_B_Gz3wjFV38_1),.dout(w_dff_B_wOBoi8IA9_1),.clk(gclk));
	jdff dff_B_fLhK1Rzp7_1(.din(w_dff_B_wOBoi8IA9_1),.dout(w_dff_B_fLhK1Rzp7_1),.clk(gclk));
	jdff dff_B_3KVuhrsb7_1(.din(w_dff_B_fLhK1Rzp7_1),.dout(w_dff_B_3KVuhrsb7_1),.clk(gclk));
	jdff dff_B_JPiiHemD4_1(.din(w_dff_B_3KVuhrsb7_1),.dout(w_dff_B_JPiiHemD4_1),.clk(gclk));
	jdff dff_A_gzuh0Vkx4_0(.dout(w_n649_0[0]),.din(w_dff_A_gzuh0Vkx4_0),.clk(gclk));
	jdff dff_A_aYiZxmTq2_0(.dout(w_dff_A_gzuh0Vkx4_0),.din(w_dff_A_aYiZxmTq2_0),.clk(gclk));
	jdff dff_A_ktkeExIF9_0(.dout(w_dff_A_aYiZxmTq2_0),.din(w_dff_A_ktkeExIF9_0),.clk(gclk));
	jdff dff_A_sfX1liGi1_0(.dout(w_dff_A_ktkeExIF9_0),.din(w_dff_A_sfX1liGi1_0),.clk(gclk));
	jdff dff_A_UkKsjaYi3_0(.dout(w_dff_A_sfX1liGi1_0),.din(w_dff_A_UkKsjaYi3_0),.clk(gclk));
	jdff dff_A_IPzIfzM83_1(.dout(w_n749_8[1]),.din(w_dff_A_IPzIfzM83_1),.clk(gclk));
	jdff dff_A_MrX19JTA6_1(.dout(w_dff_A_IPzIfzM83_1),.din(w_dff_A_MrX19JTA6_1),.clk(gclk));
	jdff dff_A_TfoO0VLG6_1(.dout(w_dff_A_MrX19JTA6_1),.din(w_dff_A_TfoO0VLG6_1),.clk(gclk));
	jdff dff_A_4CBp8hWE2_1(.dout(w_dff_A_TfoO0VLG6_1),.din(w_dff_A_4CBp8hWE2_1),.clk(gclk));
	jdff dff_A_TokjpKAi3_1(.dout(w_dff_A_4CBp8hWE2_1),.din(w_dff_A_TokjpKAi3_1),.clk(gclk));
	jdff dff_A_4Xb8R5PN6_1(.dout(w_dff_A_TokjpKAi3_1),.din(w_dff_A_4Xb8R5PN6_1),.clk(gclk));
	jdff dff_A_KSXKHMFr5_1(.dout(w_dff_A_4Xb8R5PN6_1),.din(w_dff_A_KSXKHMFr5_1),.clk(gclk));
	jdff dff_A_va9v80OY8_1(.dout(w_dff_A_KSXKHMFr5_1),.din(w_dff_A_va9v80OY8_1),.clk(gclk));
	jdff dff_A_xvASDEsW2_2(.dout(w_n749_8[2]),.din(w_dff_A_xvASDEsW2_2),.clk(gclk));
	jdff dff_A_5aatTcDn9_2(.dout(w_dff_A_xvASDEsW2_2),.din(w_dff_A_5aatTcDn9_2),.clk(gclk));
	jdff dff_A_EOLXLQar4_2(.dout(w_dff_A_5aatTcDn9_2),.din(w_dff_A_EOLXLQar4_2),.clk(gclk));
	jdff dff_A_8BBXttcs1_2(.dout(w_dff_A_EOLXLQar4_2),.din(w_dff_A_8BBXttcs1_2),.clk(gclk));
	jdff dff_A_v26VStLg6_2(.dout(w_dff_A_8BBXttcs1_2),.din(w_dff_A_v26VStLg6_2),.clk(gclk));
	jdff dff_A_NqJ4XrW94_2(.dout(w_dff_A_v26VStLg6_2),.din(w_dff_A_NqJ4XrW94_2),.clk(gclk));
	jdff dff_A_gYIti0uh0_2(.dout(w_dff_A_NqJ4XrW94_2),.din(w_dff_A_gYIti0uh0_2),.clk(gclk));
	jdff dff_A_vPH2o0Fx6_2(.dout(w_dff_A_gYIti0uh0_2),.din(w_dff_A_vPH2o0Fx6_2),.clk(gclk));
	jdff dff_B_VLxEDSOP3_1(.din(G121),.dout(w_dff_B_VLxEDSOP3_1),.clk(gclk));
	jdff dff_B_WmGzb8lC6_1(.din(w_dff_B_VLxEDSOP3_1),.dout(w_dff_B_WmGzb8lC6_1),.clk(gclk));
	jdff dff_A_LgkekKzh6_0(.dout(w_G137_4[0]),.din(w_dff_A_LgkekKzh6_0),.clk(gclk));
	jdff dff_A_EMhafzSt0_2(.dout(w_G137_4[2]),.din(w_dff_A_EMhafzSt0_2),.clk(gclk));
	jdff dff_A_1GrhbAQ60_0(.dout(w_G137_1[0]),.din(w_dff_A_1GrhbAQ60_0),.clk(gclk));
	jdff dff_A_FbGtgUkM4_0(.dout(w_dff_A_1GrhbAQ60_0),.din(w_dff_A_FbGtgUkM4_0),.clk(gclk));
	jdff dff_A_uT9IiILD1_0(.dout(w_dff_A_FbGtgUkM4_0),.din(w_dff_A_uT9IiILD1_0),.clk(gclk));
	jdff dff_A_2Vlbq6zP4_1(.dout(w_G137_1[1]),.din(w_dff_A_2Vlbq6zP4_1),.clk(gclk));
	jdff dff_A_aLRzdaaN3_1(.dout(w_dff_A_2Vlbq6zP4_1),.din(w_dff_A_aLRzdaaN3_1),.clk(gclk));
	jdff dff_B_l5H6hofB7_0(.din(n1404),.dout(w_dff_B_l5H6hofB7_0),.clk(gclk));
	jdff dff_B_hM19lVyP3_0(.din(w_dff_B_l5H6hofB7_0),.dout(w_dff_B_hM19lVyP3_0),.clk(gclk));
	jdff dff_B_gkyLdtlt2_0(.din(w_dff_B_hM19lVyP3_0),.dout(w_dff_B_gkyLdtlt2_0),.clk(gclk));
	jdff dff_B_1QXHFnVa1_0(.din(w_dff_B_gkyLdtlt2_0),.dout(w_dff_B_1QXHFnVa1_0),.clk(gclk));
	jdff dff_B_6TUkHkPM8_0(.din(w_dff_B_1QXHFnVa1_0),.dout(w_dff_B_6TUkHkPM8_0),.clk(gclk));
	jdff dff_B_IjZOVqmv6_0(.din(w_dff_B_6TUkHkPM8_0),.dout(w_dff_B_IjZOVqmv6_0),.clk(gclk));
	jdff dff_B_VaQRqlkY2_0(.din(w_dff_B_IjZOVqmv6_0),.dout(w_dff_B_VaQRqlkY2_0),.clk(gclk));
	jdff dff_B_79tvpKwJ8_0(.din(w_dff_B_VaQRqlkY2_0),.dout(w_dff_B_79tvpKwJ8_0),.clk(gclk));
	jdff dff_B_pJdWxdzJ7_0(.din(w_dff_B_79tvpKwJ8_0),.dout(w_dff_B_pJdWxdzJ7_0),.clk(gclk));
	jdff dff_B_YQnm9lIU5_0(.din(w_dff_B_pJdWxdzJ7_0),.dout(w_dff_B_YQnm9lIU5_0),.clk(gclk));
	jdff dff_B_lyyle7KZ7_0(.din(w_dff_B_YQnm9lIU5_0),.dout(w_dff_B_lyyle7KZ7_0),.clk(gclk));
	jdff dff_B_LdgVtUsB5_0(.din(w_dff_B_lyyle7KZ7_0),.dout(w_dff_B_LdgVtUsB5_0),.clk(gclk));
	jdff dff_B_CLCqBe9Z7_0(.din(w_dff_B_LdgVtUsB5_0),.dout(w_dff_B_CLCqBe9Z7_0),.clk(gclk));
	jdff dff_B_qJoWdEf78_0(.din(n1403),.dout(w_dff_B_qJoWdEf78_0),.clk(gclk));
	jdff dff_B_ILB9o4r96_2(.din(G161),.dout(w_dff_B_ILB9o4r96_2),.clk(gclk));
	jdff dff_B_xbca8g1s8_2(.din(G191),.dout(w_dff_B_xbca8g1s8_2),.clk(gclk));
	jdff dff_B_Yf51D3so8_2(.din(w_dff_B_xbca8g1s8_2),.dout(w_dff_B_Yf51D3so8_2),.clk(gclk));
	jdff dff_B_19CUk0R73_0(.din(n1400),.dout(w_dff_B_19CUk0R73_0),.clk(gclk));
	jdff dff_B_mUxvoqsy5_1(.din(n1190),.dout(w_dff_B_mUxvoqsy5_1),.clk(gclk));
	jdff dff_B_i1CuZtu87_1(.din(w_dff_B_mUxvoqsy5_1),.dout(w_dff_B_i1CuZtu87_1),.clk(gclk));
	jdff dff_B_s5tZkZh78_1(.din(w_dff_B_i1CuZtu87_1),.dout(w_dff_B_s5tZkZh78_1),.clk(gclk));
	jdff dff_B_EDHVQyou6_1(.din(w_dff_B_s5tZkZh78_1),.dout(w_dff_B_EDHVQyou6_1),.clk(gclk));
	jdff dff_B_3vonscR97_1(.din(w_dff_B_EDHVQyou6_1),.dout(w_dff_B_3vonscR97_1),.clk(gclk));
	jdff dff_B_9YS5VVDT3_1(.din(w_dff_B_3vonscR97_1),.dout(w_dff_B_9YS5VVDT3_1),.clk(gclk));
	jdff dff_B_X6IwygaY6_1(.din(w_dff_B_9YS5VVDT3_1),.dout(w_dff_B_X6IwygaY6_1),.clk(gclk));
	jdff dff_B_fGuWyEnw0_1(.din(w_dff_B_X6IwygaY6_1),.dout(w_dff_B_fGuWyEnw0_1),.clk(gclk));
	jdff dff_B_6m1TaVSt3_1(.din(w_dff_B_fGuWyEnw0_1),.dout(w_dff_B_6m1TaVSt3_1),.clk(gclk));
	jdff dff_B_QRrdICxI0_1(.din(w_dff_B_6m1TaVSt3_1),.dout(w_dff_B_QRrdICxI0_1),.clk(gclk));
	jdff dff_B_7hQKRca92_0(.din(n1194),.dout(w_dff_B_7hQKRca92_0),.clk(gclk));
	jdff dff_B_j5Vcf3KU3_0(.din(w_dff_B_7hQKRca92_0),.dout(w_dff_B_j5Vcf3KU3_0),.clk(gclk));
	jdff dff_B_ZmKB1oqU3_0(.din(w_dff_B_j5Vcf3KU3_0),.dout(w_dff_B_ZmKB1oqU3_0),.clk(gclk));
	jdff dff_B_hMJL2LoC0_0(.din(w_dff_B_ZmKB1oqU3_0),.dout(w_dff_B_hMJL2LoC0_0),.clk(gclk));
	jdff dff_B_iZowr3dP7_0(.din(w_dff_B_hMJL2LoC0_0),.dout(w_dff_B_iZowr3dP7_0),.clk(gclk));
	jdff dff_B_AYsJGttp0_0(.din(w_dff_B_iZowr3dP7_0),.dout(w_dff_B_AYsJGttp0_0),.clk(gclk));
	jdff dff_B_yWAWEi9S4_0(.din(w_dff_B_AYsJGttp0_0),.dout(w_dff_B_yWAWEi9S4_0),.clk(gclk));
	jdff dff_B_0ppLAxZZ8_0(.din(w_dff_B_yWAWEi9S4_0),.dout(w_dff_B_0ppLAxZZ8_0),.clk(gclk));
	jdff dff_A_HIvEGoOw6_1(.dout(w_G4092_6[1]),.din(w_dff_A_HIvEGoOw6_1),.clk(gclk));
	jdff dff_A_gsEPuZkl3_2(.dout(w_G4092_6[2]),.din(w_dff_A_gsEPuZkl3_2),.clk(gclk));
	jdff dff_B_1HfbonEU1_0(.din(n794),.dout(w_dff_B_1HfbonEU1_0),.clk(gclk));
	jdff dff_A_zZPHMM180_0(.dout(w_G54_0[0]),.din(w_dff_A_zZPHMM180_0),.clk(gclk));
	jdff dff_A_U5gn7ozT5_0(.dout(w_dff_A_zZPHMM180_0),.din(w_dff_A_U5gn7ozT5_0),.clk(gclk));
	jdff dff_A_mUiANa5l0_0(.dout(w_dff_A_U5gn7ozT5_0),.din(w_dff_A_mUiANa5l0_0),.clk(gclk));
	jdff dff_A_GH6Ko2pe0_0(.dout(w_dff_A_mUiANa5l0_0),.din(w_dff_A_GH6Ko2pe0_0),.clk(gclk));
	jdff dff_A_xJ27gl944_0(.dout(w_dff_A_GH6Ko2pe0_0),.din(w_dff_A_xJ27gl944_0),.clk(gclk));
	jdff dff_A_3NAf5tD94_0(.dout(w_dff_A_xJ27gl944_0),.din(w_dff_A_3NAf5tD94_0),.clk(gclk));
	jdff dff_A_YoXMoOQg9_0(.dout(w_dff_A_3NAf5tD94_0),.din(w_dff_A_YoXMoOQg9_0),.clk(gclk));
	jdff dff_A_YzfQGdLU0_0(.dout(w_dff_A_YoXMoOQg9_0),.din(w_dff_A_YzfQGdLU0_0),.clk(gclk));
	jdff dff_A_Kz347l3Y3_1(.dout(w_G54_0[1]),.din(w_dff_A_Kz347l3Y3_1),.clk(gclk));
	jdff dff_A_ZRRNMtCC4_1(.dout(w_dff_A_Kz347l3Y3_1),.din(w_dff_A_ZRRNMtCC4_1),.clk(gclk));
	jdff dff_A_PcRgOJNS6_1(.dout(w_dff_A_ZRRNMtCC4_1),.din(w_dff_A_PcRgOJNS6_1),.clk(gclk));
	jdff dff_A_Qmr2zLjk1_0(.dout(w_n737_1[0]),.din(w_dff_A_Qmr2zLjk1_0),.clk(gclk));
	jdff dff_A_pFcrzKxj4_0(.dout(w_dff_A_Qmr2zLjk1_0),.din(w_dff_A_pFcrzKxj4_0),.clk(gclk));
	jdff dff_A_epYM8dkX3_0(.dout(w_n749_9[0]),.din(w_dff_A_epYM8dkX3_0),.clk(gclk));
	jdff dff_A_ZpYjSdeL0_2(.dout(w_n749_9[2]),.din(w_dff_A_ZpYjSdeL0_2),.clk(gclk));
	jdff dff_A_pd2Fzd3t8_2(.dout(w_dff_A_ZpYjSdeL0_2),.din(w_dff_A_pd2Fzd3t8_2),.clk(gclk));
	jdff dff_A_tfnyL9Sh2_2(.dout(w_dff_A_pd2Fzd3t8_2),.din(w_dff_A_tfnyL9Sh2_2),.clk(gclk));
	jdff dff_A_AFUj7jRN3_2(.dout(w_dff_A_tfnyL9Sh2_2),.din(w_dff_A_AFUj7jRN3_2),.clk(gclk));
	jdff dff_A_ivQD28eW9_2(.dout(w_dff_A_AFUj7jRN3_2),.din(w_dff_A_ivQD28eW9_2),.clk(gclk));
	jdff dff_A_OAgB92s37_2(.dout(w_dff_A_ivQD28eW9_2),.din(w_dff_A_OAgB92s37_2),.clk(gclk));
	jdff dff_A_jfWpfTDY8_2(.dout(w_dff_A_OAgB92s37_2),.din(w_dff_A_jfWpfTDY8_2),.clk(gclk));
	jdff dff_A_vIa3IA8D7_2(.dout(w_dff_A_jfWpfTDY8_2),.din(w_dff_A_vIa3IA8D7_2),.clk(gclk));
	jdff dff_A_O9JtnTrn7_2(.dout(w_dff_A_vIa3IA8D7_2),.din(w_dff_A_O9JtnTrn7_2),.clk(gclk));
	jdff dff_A_LPew5BSL7_2(.dout(w_dff_A_O9JtnTrn7_2),.din(w_dff_A_LPew5BSL7_2),.clk(gclk));
	jdff dff_A_aaTwBJgH3_0(.dout(w_G123_0[0]),.din(w_dff_A_aaTwBJgH3_0),.clk(gclk));
	jdff dff_A_ySZyEEnd2_0(.dout(w_dff_A_aaTwBJgH3_0),.din(w_dff_A_ySZyEEnd2_0),.clk(gclk));
	jdff dff_A_AgVAjbLj8_0(.dout(w_G1691_2[0]),.din(w_dff_A_AgVAjbLj8_0),.clk(gclk));
	jdff dff_A_I9Uio7DV6_1(.dout(w_G1691_2[1]),.din(w_dff_A_I9Uio7DV6_1),.clk(gclk));
	jdff dff_A_OVor5WGP0_1(.dout(w_n1007_1[1]),.din(w_dff_A_OVor5WGP0_1),.clk(gclk));
	jdff dff_A_rWnb6qNO3_1(.dout(w_dff_A_OVor5WGP0_1),.din(w_dff_A_rWnb6qNO3_1),.clk(gclk));
	jdff dff_A_DJ51JjTe3_2(.dout(w_n1007_1[2]),.din(w_dff_A_DJ51JjTe3_2),.clk(gclk));
	jdff dff_A_LNXDQdP04_2(.dout(w_dff_A_DJ51JjTe3_2),.din(w_dff_A_LNXDQdP04_2),.clk(gclk));
	jdff dff_A_wCJR7GEK4_0(.dout(w_n1007_0[0]),.din(w_dff_A_wCJR7GEK4_0),.clk(gclk));
	jdff dff_A_MZ0SB1Ps2_0(.dout(w_dff_A_wCJR7GEK4_0),.din(w_dff_A_MZ0SB1Ps2_0),.clk(gclk));
	jdff dff_A_7Vx558mB1_0(.dout(w_dff_A_MZ0SB1Ps2_0),.din(w_dff_A_7Vx558mB1_0),.clk(gclk));
	jdff dff_A_KdQ8m5yz3_1(.dout(w_n1007_0[1]),.din(w_dff_A_KdQ8m5yz3_1),.clk(gclk));
	jdff dff_B_dq8pL2kY4_3(.din(n1007),.dout(w_dff_B_dq8pL2kY4_3),.clk(gclk));
	jdff dff_B_OJWZcLhd3_3(.din(w_dff_B_dq8pL2kY4_3),.dout(w_dff_B_OJWZcLhd3_3),.clk(gclk));
	jdff dff_B_7s44NM8a3_3(.din(w_dff_B_OJWZcLhd3_3),.dout(w_dff_B_7s44NM8a3_3),.clk(gclk));
	jdff dff_B_olm5LHQs1_3(.din(w_dff_B_7s44NM8a3_3),.dout(w_dff_B_olm5LHQs1_3),.clk(gclk));
	jdff dff_B_hcZfaSak9_3(.din(w_dff_B_olm5LHQs1_3),.dout(w_dff_B_hcZfaSak9_3),.clk(gclk));
	jdff dff_B_eGRdpZ4f2_3(.din(w_dff_B_hcZfaSak9_3),.dout(w_dff_B_eGRdpZ4f2_3),.clk(gclk));
	jdff dff_B_GOYTWufs0_3(.din(w_dff_B_eGRdpZ4f2_3),.dout(w_dff_B_GOYTWufs0_3),.clk(gclk));
	jdff dff_B_aZlbDHqr4_3(.din(w_dff_B_GOYTWufs0_3),.dout(w_dff_B_aZlbDHqr4_3),.clk(gclk));
	jdff dff_B_sxP123rE8_3(.din(w_dff_B_aZlbDHqr4_3),.dout(w_dff_B_sxP123rE8_3),.clk(gclk));
	jdff dff_B_aj7JN7wK2_1(.din(n1230),.dout(w_dff_B_aj7JN7wK2_1),.clk(gclk));
	jdff dff_B_n8aV7hLb3_1(.din(w_dff_B_aj7JN7wK2_1),.dout(w_dff_B_n8aV7hLb3_1),.clk(gclk));
	jdff dff_B_jHBprmgF4_1(.din(w_dff_B_n8aV7hLb3_1),.dout(w_dff_B_jHBprmgF4_1),.clk(gclk));
	jdff dff_B_ww1Bb9T24_1(.din(w_dff_B_jHBprmgF4_1),.dout(w_dff_B_ww1Bb9T24_1),.clk(gclk));
	jdff dff_B_NMJHJAad8_1(.din(w_dff_B_ww1Bb9T24_1),.dout(w_dff_B_NMJHJAad8_1),.clk(gclk));
	jdff dff_B_vzvGqzOA3_1(.din(w_dff_B_NMJHJAad8_1),.dout(w_dff_B_vzvGqzOA3_1),.clk(gclk));
	jdff dff_B_74pk0Hhd3_1(.din(w_dff_B_vzvGqzOA3_1),.dout(w_dff_B_74pk0Hhd3_1),.clk(gclk));
	jdff dff_B_A20ilHKs1_1(.din(w_dff_B_74pk0Hhd3_1),.dout(w_dff_B_A20ilHKs1_1),.clk(gclk));
	jdff dff_B_7wfDf1vh2_1(.din(w_dff_B_A20ilHKs1_1),.dout(w_dff_B_7wfDf1vh2_1),.clk(gclk));
	jdff dff_B_VabMyFf63_1(.din(w_dff_B_7wfDf1vh2_1),.dout(w_dff_B_VabMyFf63_1),.clk(gclk));
	jdff dff_B_w4R4vMFd2_1(.din(w_dff_B_VabMyFf63_1),.dout(w_dff_B_w4R4vMFd2_1),.clk(gclk));
	jdff dff_B_Z5W0Ta4I1_1(.din(w_dff_B_w4R4vMFd2_1),.dout(w_dff_B_Z5W0Ta4I1_1),.clk(gclk));
	jdff dff_B_Q3TlPJxP2_1(.din(n1232),.dout(w_dff_B_Q3TlPJxP2_1),.clk(gclk));
	jdff dff_B_h2nWPywg7_1(.din(w_dff_B_Q3TlPJxP2_1),.dout(w_dff_B_h2nWPywg7_1),.clk(gclk));
	jdff dff_B_4yEh5cb65_1(.din(w_dff_B_h2nWPywg7_1),.dout(w_dff_B_4yEh5cb65_1),.clk(gclk));
	jdff dff_B_5gXxx9iH9_1(.din(w_dff_B_4yEh5cb65_1),.dout(w_dff_B_5gXxx9iH9_1),.clk(gclk));
	jdff dff_B_oPnMMCzm4_1(.din(w_dff_B_5gXxx9iH9_1),.dout(w_dff_B_oPnMMCzm4_1),.clk(gclk));
	jdff dff_B_bbVZubYC8_1(.din(w_dff_B_oPnMMCzm4_1),.dout(w_dff_B_bbVZubYC8_1),.clk(gclk));
	jdff dff_B_tL06usoO3_1(.din(w_dff_B_bbVZubYC8_1),.dout(w_dff_B_tL06usoO3_1),.clk(gclk));
	jdff dff_B_4qdcCPL31_1(.din(w_dff_B_tL06usoO3_1),.dout(w_dff_B_4qdcCPL31_1),.clk(gclk));
	jdff dff_B_lViDy4wq4_1(.din(w_dff_B_4qdcCPL31_1),.dout(w_dff_B_lViDy4wq4_1),.clk(gclk));
	jdff dff_B_DQ2VEUdN9_1(.din(n937),.dout(w_dff_B_DQ2VEUdN9_1),.clk(gclk));
	jdff dff_B_uLRIozM67_1(.din(w_dff_B_DQ2VEUdN9_1),.dout(w_dff_B_uLRIozM67_1),.clk(gclk));
	jdff dff_B_Uv48ZgDn4_1(.din(w_dff_B_uLRIozM67_1),.dout(w_dff_B_Uv48ZgDn4_1),.clk(gclk));
	jdff dff_B_ntnPPHuU4_1(.din(w_dff_B_Uv48ZgDn4_1),.dout(w_dff_B_ntnPPHuU4_1),.clk(gclk));
	jdff dff_B_GtS36WCP5_1(.din(w_dff_B_ntnPPHuU4_1),.dout(w_dff_B_GtS36WCP5_1),.clk(gclk));
	jdff dff_B_twIV5z9g9_1(.din(w_dff_B_GtS36WCP5_1),.dout(w_dff_B_twIV5z9g9_1),.clk(gclk));
	jdff dff_B_XK3P6TBA8_1(.din(w_dff_B_twIV5z9g9_1),.dout(w_dff_B_XK3P6TBA8_1),.clk(gclk));
	jdff dff_B_vttHX3IB0_1(.din(w_dff_B_XK3P6TBA8_1),.dout(w_dff_B_vttHX3IB0_1),.clk(gclk));
	jdff dff_B_acIVQIkn5_1(.din(n866),.dout(w_dff_B_acIVQIkn5_1),.clk(gclk));
	jdff dff_B_fqtln7K09_1(.din(w_dff_B_acIVQIkn5_1),.dout(w_dff_B_fqtln7K09_1),.clk(gclk));
	jdff dff_A_FvxgaWv24_1(.dout(w_G4_0[1]),.din(w_dff_A_FvxgaWv24_1),.clk(gclk));
	jdff dff_B_cg5oOrxl3_3(.din(G4),.dout(w_dff_B_cg5oOrxl3_3),.clk(gclk));
	jdff dff_B_fTYU1qt46_3(.din(w_dff_B_cg5oOrxl3_3),.dout(w_dff_B_fTYU1qt46_3),.clk(gclk));
	jdff dff_B_FgEDfhrY8_3(.din(w_dff_B_fTYU1qt46_3),.dout(w_dff_B_FgEDfhrY8_3),.clk(gclk));
	jdff dff_B_snmdC2Cj1_3(.din(w_dff_B_FgEDfhrY8_3),.dout(w_dff_B_snmdC2Cj1_3),.clk(gclk));
	jdff dff_B_DAGiszlx7_3(.din(w_dff_B_snmdC2Cj1_3),.dout(w_dff_B_DAGiszlx7_3),.clk(gclk));
	jdff dff_A_Z9NEU7h14_0(.dout(w_n1201_0[0]),.din(w_dff_A_Z9NEU7h14_0),.clk(gclk));
	jdff dff_A_fRRVBTaS4_1(.dout(w_n1201_0[1]),.din(w_dff_A_fRRVBTaS4_1),.clk(gclk));
	jdff dff_A_1DbhtSJM9_1(.dout(w_dff_A_fRRVBTaS4_1),.din(w_dff_A_1DbhtSJM9_1),.clk(gclk));
	jdff dff_B_bC0IgXju0_3(.din(n1201),.dout(w_dff_B_bC0IgXju0_3),.clk(gclk));
	jdff dff_B_sjm3CCUl6_3(.din(w_dff_B_bC0IgXju0_3),.dout(w_dff_B_sjm3CCUl6_3),.clk(gclk));
	jdff dff_B_3uFfUMeF0_3(.din(w_dff_B_sjm3CCUl6_3),.dout(w_dff_B_3uFfUMeF0_3),.clk(gclk));
	jdff dff_B_bYGZBYfd5_3(.din(w_dff_B_3uFfUMeF0_3),.dout(w_dff_B_bYGZBYfd5_3),.clk(gclk));
	jdff dff_B_rohqyra99_3(.din(w_dff_B_bYGZBYfd5_3),.dout(w_dff_B_rohqyra99_3),.clk(gclk));
	jdff dff_B_ektyliWy8_3(.din(w_dff_B_rohqyra99_3),.dout(w_dff_B_ektyliWy8_3),.clk(gclk));
	jdff dff_B_FOcgl5Ig0_3(.din(w_dff_B_ektyliWy8_3),.dout(w_dff_B_FOcgl5Ig0_3),.clk(gclk));
	jdff dff_B_HqbpNqwJ4_3(.din(w_dff_B_FOcgl5Ig0_3),.dout(w_dff_B_HqbpNqwJ4_3),.clk(gclk));
	jdff dff_B_K8qLVtPj7_3(.din(w_dff_B_HqbpNqwJ4_3),.dout(w_dff_B_K8qLVtPj7_3),.clk(gclk));
	jdff dff_B_sWMDizUz3_3(.din(w_dff_B_K8qLVtPj7_3),.dout(w_dff_B_sWMDizUz3_3),.clk(gclk));
	jdff dff_A_2uR8uR269_0(.dout(w_G4092_5[0]),.din(w_dff_A_2uR8uR269_0),.clk(gclk));
	jdff dff_A_Z2gtRlb27_0(.dout(w_dff_A_2uR8uR269_0),.din(w_dff_A_Z2gtRlb27_0),.clk(gclk));
	jdff dff_A_gyfPRPyR1_0(.dout(w_dff_A_Z2gtRlb27_0),.din(w_dff_A_gyfPRPyR1_0),.clk(gclk));
	jdff dff_A_gJuftH4B6_0(.dout(w_dff_A_gyfPRPyR1_0),.din(w_dff_A_gJuftH4B6_0),.clk(gclk));
	jdff dff_A_htGz29MJ5_1(.dout(w_G4092_5[1]),.din(w_dff_A_htGz29MJ5_1),.clk(gclk));
	jdff dff_A_BdUeDT9A7_1(.dout(w_dff_A_htGz29MJ5_1),.din(w_dff_A_BdUeDT9A7_1),.clk(gclk));
	jdff dff_A_ocZONREd9_1(.dout(w_dff_A_BdUeDT9A7_1),.din(w_dff_A_ocZONREd9_1),.clk(gclk));
	jdff dff_A_OdaYqszP2_1(.dout(w_dff_A_ocZONREd9_1),.din(w_dff_A_OdaYqszP2_1),.clk(gclk));
	jdff dff_A_ndj4ZMr78_0(.dout(w_n749_7[0]),.din(w_dff_A_ndj4ZMr78_0),.clk(gclk));
	jdff dff_A_0va8SZaj1_0(.dout(w_dff_A_ndj4ZMr78_0),.din(w_dff_A_0va8SZaj1_0),.clk(gclk));
	jdff dff_A_fGBivi058_0(.dout(w_dff_A_0va8SZaj1_0),.din(w_dff_A_fGBivi058_0),.clk(gclk));
	jdff dff_A_m8v6DEEs9_0(.dout(w_dff_A_fGBivi058_0),.din(w_dff_A_m8v6DEEs9_0),.clk(gclk));
	jdff dff_A_HCwU8CDC3_0(.dout(w_dff_A_m8v6DEEs9_0),.din(w_dff_A_HCwU8CDC3_0),.clk(gclk));
	jdff dff_A_OePnhah88_0(.dout(w_dff_A_HCwU8CDC3_0),.din(w_dff_A_OePnhah88_0),.clk(gclk));
	jdff dff_A_reBb0rZg7_0(.dout(w_dff_A_OePnhah88_0),.din(w_dff_A_reBb0rZg7_0),.clk(gclk));
	jdff dff_A_Og6BaQ0q0_0(.dout(w_dff_A_reBb0rZg7_0),.din(w_dff_A_Og6BaQ0q0_0),.clk(gclk));
	jdff dff_A_DCplg5J53_0(.dout(w_dff_A_Og6BaQ0q0_0),.din(w_dff_A_DCplg5J53_0),.clk(gclk));
	jdff dff_A_9g7kbvuQ0_0(.dout(w_dff_A_DCplg5J53_0),.din(w_dff_A_9g7kbvuQ0_0),.clk(gclk));
	jdff dff_A_kmiPpjBM6_0(.dout(w_n749_2[0]),.din(w_dff_A_kmiPpjBM6_0),.clk(gclk));
	jdff dff_A_GaxJsdja4_1(.dout(w_n749_2[1]),.din(w_dff_A_GaxJsdja4_1),.clk(gclk));
	jdff dff_B_6DIDidrH7_1(.din(G115),.dout(w_dff_B_6DIDidrH7_1),.clk(gclk));
	jdff dff_B_DhEh2tGG5_1(.din(w_dff_B_6DIDidrH7_1),.dout(w_dff_B_DhEh2tGG5_1),.clk(gclk));
	jdff dff_B_5MmuVgut9_0(.din(n1505),.dout(w_dff_B_5MmuVgut9_0),.clk(gclk));
	jdff dff_B_HevVietn9_0(.din(w_dff_B_5MmuVgut9_0),.dout(w_dff_B_HevVietn9_0),.clk(gclk));
	jdff dff_B_lGoLgcqN5_0(.din(w_dff_B_HevVietn9_0),.dout(w_dff_B_lGoLgcqN5_0),.clk(gclk));
	jdff dff_B_cmkLnFvo7_0(.din(w_dff_B_lGoLgcqN5_0),.dout(w_dff_B_cmkLnFvo7_0),.clk(gclk));
	jdff dff_B_c3VDItoR1_0(.din(w_dff_B_cmkLnFvo7_0),.dout(w_dff_B_c3VDItoR1_0),.clk(gclk));
	jdff dff_B_FHZJGFsU5_0(.din(w_dff_B_c3VDItoR1_0),.dout(w_dff_B_FHZJGFsU5_0),.clk(gclk));
	jdff dff_B_fXYcpbP90_0(.din(w_dff_B_FHZJGFsU5_0),.dout(w_dff_B_fXYcpbP90_0),.clk(gclk));
	jdff dff_B_p40PdWak6_0(.din(w_dff_B_fXYcpbP90_0),.dout(w_dff_B_p40PdWak6_0),.clk(gclk));
	jdff dff_B_1j1dvsn16_0(.din(w_dff_B_p40PdWak6_0),.dout(w_dff_B_1j1dvsn16_0),.clk(gclk));
	jdff dff_B_ZFHAwiAm3_0(.din(w_dff_B_1j1dvsn16_0),.dout(w_dff_B_ZFHAwiAm3_0),.clk(gclk));
	jdff dff_B_KxcdlZft6_0(.din(w_dff_B_ZFHAwiAm3_0),.dout(w_dff_B_KxcdlZft6_0),.clk(gclk));
	jdff dff_B_65cWIXBY4_0(.din(w_dff_B_KxcdlZft6_0),.dout(w_dff_B_65cWIXBY4_0),.clk(gclk));
	jdff dff_B_hUtUCUUQ1_0(.din(w_dff_B_65cWIXBY4_0),.dout(w_dff_B_hUtUCUUQ1_0),.clk(gclk));
	jdff dff_B_O2wXCame6_0(.din(w_dff_B_hUtUCUUQ1_0),.dout(w_dff_B_O2wXCame6_0),.clk(gclk));
	jdff dff_B_O0bUaAGo0_1(.din(G120),.dout(w_dff_B_O0bUaAGo0_1),.clk(gclk));
	jdff dff_B_RgUjy1Im3_1(.din(w_dff_B_O0bUaAGo0_1),.dout(w_dff_B_RgUjy1Im3_1),.clk(gclk));
	jdff dff_B_azXsQYim8_1(.din(w_dff_B_RgUjy1Im3_1),.dout(w_dff_B_azXsQYim8_1),.clk(gclk));
	jdff dff_B_M85N0d3R5_0(.din(n1666),.dout(w_dff_B_M85N0d3R5_0),.clk(gclk));
	jdff dff_B_aS2Vih3x8_0(.din(w_dff_B_M85N0d3R5_0),.dout(w_dff_B_aS2Vih3x8_0),.clk(gclk));
	jdff dff_B_3vhFUZGe2_0(.din(w_dff_B_aS2Vih3x8_0),.dout(w_dff_B_3vhFUZGe2_0),.clk(gclk));
	jdff dff_B_3Czds3JZ4_0(.din(w_dff_B_3vhFUZGe2_0),.dout(w_dff_B_3Czds3JZ4_0),.clk(gclk));
	jdff dff_B_8VeSpgzn0_0(.din(w_dff_B_3Czds3JZ4_0),.dout(w_dff_B_8VeSpgzn0_0),.clk(gclk));
	jdff dff_B_EjvNbbix8_0(.din(w_dff_B_8VeSpgzn0_0),.dout(w_dff_B_EjvNbbix8_0),.clk(gclk));
	jdff dff_B_NZ8cTK9S6_0(.din(w_dff_B_EjvNbbix8_0),.dout(w_dff_B_NZ8cTK9S6_0),.clk(gclk));
	jdff dff_B_hAQsKl8j3_0(.din(w_dff_B_NZ8cTK9S6_0),.dout(w_dff_B_hAQsKl8j3_0),.clk(gclk));
	jdff dff_B_mmXdeAtT8_0(.din(w_dff_B_hAQsKl8j3_0),.dout(w_dff_B_mmXdeAtT8_0),.clk(gclk));
	jdff dff_B_dxH2p7S05_0(.din(w_dff_B_mmXdeAtT8_0),.dout(w_dff_B_dxH2p7S05_0),.clk(gclk));
	jdff dff_B_MORgfw408_0(.din(w_dff_B_dxH2p7S05_0),.dout(w_dff_B_MORgfw408_0),.clk(gclk));
	jdff dff_B_aPJmDf3D1_0(.din(w_dff_B_MORgfw408_0),.dout(w_dff_B_aPJmDf3D1_0),.clk(gclk));
	jdff dff_B_SBDAbhRx1_1(.din(G118),.dout(w_dff_B_SBDAbhRx1_1),.clk(gclk));
	jdff dff_B_zjSNR6RA8_1(.din(w_dff_B_SBDAbhRx1_1),.dout(w_dff_B_zjSNR6RA8_1),.clk(gclk));
	jdff dff_B_3I40ZzvN4_1(.din(w_dff_B_zjSNR6RA8_1),.dout(w_dff_B_3I40ZzvN4_1),.clk(gclk));
	jdff dff_A_vZjRr1JT6_0(.dout(w_G4092_9[0]),.din(w_dff_A_vZjRr1JT6_0),.clk(gclk));
	jdff dff_A_fZCZTDzz3_0(.dout(w_dff_A_vZjRr1JT6_0),.din(w_dff_A_fZCZTDzz3_0),.clk(gclk));
	jdff dff_A_LlDY6nhZ3_0(.dout(w_dff_A_fZCZTDzz3_0),.din(w_dff_A_LlDY6nhZ3_0),.clk(gclk));
	jdff dff_A_YcAksiy49_1(.dout(w_G4092_9[1]),.din(w_dff_A_YcAksiy49_1),.clk(gclk));
	jdff dff_A_qcE08D9l5_1(.dout(w_dff_A_YcAksiy49_1),.din(w_dff_A_qcE08D9l5_1),.clk(gclk));
	jdff dff_A_gmf8R17O2_1(.dout(w_dff_A_qcE08D9l5_1),.din(w_dff_A_gmf8R17O2_1),.clk(gclk));
	jdff dff_A_nWhYw17j6_0(.dout(w_G4092_2[0]),.din(w_dff_A_nWhYw17j6_0),.clk(gclk));
	jdff dff_A_OXZn5mpO3_0(.dout(w_dff_A_nWhYw17j6_0),.din(w_dff_A_OXZn5mpO3_0),.clk(gclk));
	jdff dff_A_J7Y9NuWP2_0(.dout(w_dff_A_OXZn5mpO3_0),.din(w_dff_A_J7Y9NuWP2_0),.clk(gclk));
	jdff dff_A_UmKEUOuR3_1(.dout(w_G4092_2[1]),.din(w_dff_A_UmKEUOuR3_1),.clk(gclk));
	jdff dff_A_VhiGAHnE3_1(.dout(w_dff_A_UmKEUOuR3_1),.din(w_dff_A_VhiGAHnE3_1),.clk(gclk));
	jdff dff_A_RqxKpO2m6_1(.dout(w_dff_A_VhiGAHnE3_1),.din(w_dff_A_RqxKpO2m6_1),.clk(gclk));
	jdff dff_A_BXfgeJqU2_0(.dout(w_n749_13[0]),.din(w_dff_A_BXfgeJqU2_0),.clk(gclk));
	jdff dff_A_CyS8Dk7A7_0(.dout(w_dff_A_BXfgeJqU2_0),.din(w_dff_A_CyS8Dk7A7_0),.clk(gclk));
	jdff dff_B_XtHccHky7_1(.din(n1671),.dout(w_dff_B_XtHccHky7_1),.clk(gclk));
	jdff dff_B_aMDTVFoh8_1(.din(w_dff_B_XtHccHky7_1),.dout(w_dff_B_aMDTVFoh8_1),.clk(gclk));
	jdff dff_B_GBfP93RP8_1(.din(w_dff_B_aMDTVFoh8_1),.dout(w_dff_B_GBfP93RP8_1),.clk(gclk));
	jdff dff_B_zWMPtATj4_1(.din(w_dff_B_GBfP93RP8_1),.dout(w_dff_B_zWMPtATj4_1),.clk(gclk));
	jdff dff_B_XgLeXI1C6_1(.din(w_dff_B_zWMPtATj4_1),.dout(w_dff_B_XgLeXI1C6_1),.clk(gclk));
	jdff dff_B_cWHhm0ZB5_1(.din(w_dff_B_XgLeXI1C6_1),.dout(w_dff_B_cWHhm0ZB5_1),.clk(gclk));
	jdff dff_B_2QlkjtgU7_1(.din(w_dff_B_cWHhm0ZB5_1),.dout(w_dff_B_2QlkjtgU7_1),.clk(gclk));
	jdff dff_B_Av4cuTYC5_1(.din(w_dff_B_2QlkjtgU7_1),.dout(w_dff_B_Av4cuTYC5_1),.clk(gclk));
	jdff dff_B_YHHqLzvp5_1(.din(w_dff_B_Av4cuTYC5_1),.dout(w_dff_B_YHHqLzvp5_1),.clk(gclk));
	jdff dff_B_SdTOLAfJ3_1(.din(w_dff_B_YHHqLzvp5_1),.dout(w_dff_B_SdTOLAfJ3_1),.clk(gclk));
	jdff dff_B_Lo0ttyBg6_1(.din(w_dff_B_SdTOLAfJ3_1),.dout(w_dff_B_Lo0ttyBg6_1),.clk(gclk));
	jdff dff_B_hyJSHAJk7_1(.din(w_dff_B_Lo0ttyBg6_1),.dout(w_dff_B_hyJSHAJk7_1),.clk(gclk));
	jdff dff_B_ldIlUEcz3_1(.din(w_dff_B_hyJSHAJk7_1),.dout(w_dff_B_ldIlUEcz3_1),.clk(gclk));
	jdff dff_B_g5hIqvbP5_1(.din(w_dff_B_ldIlUEcz3_1),.dout(w_dff_B_g5hIqvbP5_1),.clk(gclk));
	jdff dff_B_hCzt0KMs8_1(.din(w_dff_B_g5hIqvbP5_1),.dout(w_dff_B_hCzt0KMs8_1),.clk(gclk));
	jdff dff_B_bWI8XA087_1(.din(w_dff_B_hCzt0KMs8_1),.dout(w_dff_B_bWI8XA087_1),.clk(gclk));
	jdff dff_B_YpajO6WT8_1(.din(w_dff_B_bWI8XA087_1),.dout(w_dff_B_YpajO6WT8_1),.clk(gclk));
	jdff dff_B_WSmL8jgO8_1(.din(w_dff_B_YpajO6WT8_1),.dout(w_dff_B_WSmL8jgO8_1),.clk(gclk));
	jdff dff_B_fknJvqcH6_1(.din(n1676),.dout(w_dff_B_fknJvqcH6_1),.clk(gclk));
	jdff dff_B_eVwt8nyF3_1(.din(w_dff_B_fknJvqcH6_1),.dout(w_dff_B_eVwt8nyF3_1),.clk(gclk));
	jdff dff_B_eFyZ6tLA9_1(.din(w_dff_B_eVwt8nyF3_1),.dout(w_dff_B_eFyZ6tLA9_1),.clk(gclk));
	jdff dff_A_nYSjvWRp9_1(.dout(w_n800_1[1]),.din(w_dff_A_nYSjvWRp9_1),.clk(gclk));
	jdff dff_A_gJMNuNEo9_1(.dout(w_dff_A_nYSjvWRp9_1),.din(w_dff_A_gJMNuNEo9_1),.clk(gclk));
	jdff dff_A_Vov5Eqjr7_1(.dout(w_dff_A_gJMNuNEo9_1),.din(w_dff_A_Vov5Eqjr7_1),.clk(gclk));
	jdff dff_A_9oO42x6x2_1(.dout(w_dff_A_Vov5Eqjr7_1),.din(w_dff_A_9oO42x6x2_1),.clk(gclk));
	jdff dff_A_SAZg6pwQ3_1(.dout(w_dff_A_9oO42x6x2_1),.din(w_dff_A_SAZg6pwQ3_1),.clk(gclk));
	jdff dff_A_FZATdq0d0_1(.dout(w_dff_A_SAZg6pwQ3_1),.din(w_dff_A_FZATdq0d0_1),.clk(gclk));
	jdff dff_A_nhAMpXcO2_1(.dout(w_dff_A_FZATdq0d0_1),.din(w_dff_A_nhAMpXcO2_1),.clk(gclk));
	jdff dff_A_XpWiRjSv1_1(.dout(w_dff_A_nhAMpXcO2_1),.din(w_dff_A_XpWiRjSv1_1),.clk(gclk));
	jdff dff_A_H4koN1yK6_1(.dout(w_dff_A_XpWiRjSv1_1),.din(w_dff_A_H4koN1yK6_1),.clk(gclk));
	jdff dff_A_aIyR34lZ1_1(.dout(w_dff_A_H4koN1yK6_1),.din(w_dff_A_aIyR34lZ1_1),.clk(gclk));
	jdff dff_A_UAkVqxtG8_1(.dout(w_dff_A_aIyR34lZ1_1),.din(w_dff_A_UAkVqxtG8_1),.clk(gclk));
	jdff dff_A_Ox8FuV760_1(.dout(w_dff_A_UAkVqxtG8_1),.din(w_dff_A_Ox8FuV760_1),.clk(gclk));
	jdff dff_A_brTgIcGo0_2(.dout(w_n800_1[2]),.din(w_dff_A_brTgIcGo0_2),.clk(gclk));
	jdff dff_A_BfrDUMvr9_2(.dout(w_dff_A_brTgIcGo0_2),.din(w_dff_A_BfrDUMvr9_2),.clk(gclk));
	jdff dff_A_3y2Y8qjJ8_2(.dout(w_dff_A_BfrDUMvr9_2),.din(w_dff_A_3y2Y8qjJ8_2),.clk(gclk));
	jdff dff_A_7pV8ofrA4_2(.dout(w_dff_A_3y2Y8qjJ8_2),.din(w_dff_A_7pV8ofrA4_2),.clk(gclk));
	jdff dff_A_mZ2chaRB9_2(.dout(w_dff_A_7pV8ofrA4_2),.din(w_dff_A_mZ2chaRB9_2),.clk(gclk));
	jdff dff_A_hlHgs7Jf6_2(.dout(w_dff_A_mZ2chaRB9_2),.din(w_dff_A_hlHgs7Jf6_2),.clk(gclk));
	jdff dff_A_hXs8wCCM1_2(.dout(w_dff_A_hlHgs7Jf6_2),.din(w_dff_A_hXs8wCCM1_2),.clk(gclk));
	jdff dff_A_DSftXgBI3_2(.dout(w_dff_A_hXs8wCCM1_2),.din(w_dff_A_DSftXgBI3_2),.clk(gclk));
	jdff dff_A_3WfPR8XK6_1(.dout(w_n800_0[1]),.din(w_dff_A_3WfPR8XK6_1),.clk(gclk));
	jdff dff_A_5Yf3umdy3_1(.dout(w_dff_A_3WfPR8XK6_1),.din(w_dff_A_5Yf3umdy3_1),.clk(gclk));
	jdff dff_A_EWRqoXPE5_1(.dout(w_dff_A_5Yf3umdy3_1),.din(w_dff_A_EWRqoXPE5_1),.clk(gclk));
	jdff dff_A_1Vrka3nn3_1(.dout(w_dff_A_EWRqoXPE5_1),.din(w_dff_A_1Vrka3nn3_1),.clk(gclk));
	jdff dff_A_0gF9QG569_1(.dout(w_dff_A_1Vrka3nn3_1),.din(w_dff_A_0gF9QG569_1),.clk(gclk));
	jdff dff_A_wpr6RYoH4_1(.dout(w_dff_A_0gF9QG569_1),.din(w_dff_A_wpr6RYoH4_1),.clk(gclk));
	jdff dff_A_3NmwBAyE8_1(.dout(w_dff_A_wpr6RYoH4_1),.din(w_dff_A_3NmwBAyE8_1),.clk(gclk));
	jdff dff_A_mPQrTci48_2(.dout(w_n800_0[2]),.din(w_dff_A_mPQrTci48_2),.clk(gclk));
	jdff dff_A_hUqzAPow8_2(.dout(w_dff_A_mPQrTci48_2),.din(w_dff_A_hUqzAPow8_2),.clk(gclk));
	jdff dff_A_hOX6vQYZ3_2(.dout(w_dff_A_hUqzAPow8_2),.din(w_dff_A_hOX6vQYZ3_2),.clk(gclk));
	jdff dff_B_SunLTDhH8_3(.din(n800),.dout(w_dff_B_SunLTDhH8_3),.clk(gclk));
	jdff dff_B_NDU8Wrav9_3(.din(w_dff_B_SunLTDhH8_3),.dout(w_dff_B_NDU8Wrav9_3),.clk(gclk));
	jdff dff_B_CFEXWSiw5_3(.din(w_dff_B_NDU8Wrav9_3),.dout(w_dff_B_CFEXWSiw5_3),.clk(gclk));
	jdff dff_B_ifJc5Jiq5_3(.din(w_dff_B_CFEXWSiw5_3),.dout(w_dff_B_ifJc5Jiq5_3),.clk(gclk));
	jdff dff_B_GimFYhXu0_3(.din(w_dff_B_ifJc5Jiq5_3),.dout(w_dff_B_GimFYhXu0_3),.clk(gclk));
	jdff dff_B_w6LEIGgm5_3(.din(w_dff_B_GimFYhXu0_3),.dout(w_dff_B_w6LEIGgm5_3),.clk(gclk));
	jdff dff_B_qceph8Jg1_1(.din(n1668),.dout(w_dff_B_qceph8Jg1_1),.clk(gclk));
	jdff dff_B_gqy9HQBB1_1(.din(w_dff_B_qceph8Jg1_1),.dout(w_dff_B_gqy9HQBB1_1),.clk(gclk));
	jdff dff_A_Ny8CW9t27_0(.dout(w_n797_3[0]),.din(w_dff_A_Ny8CW9t27_0),.clk(gclk));
	jdff dff_A_I6xnkGRK0_0(.dout(w_dff_A_Ny8CW9t27_0),.din(w_dff_A_I6xnkGRK0_0),.clk(gclk));
	jdff dff_A_HOiwcsfq9_0(.dout(w_dff_A_I6xnkGRK0_0),.din(w_dff_A_HOiwcsfq9_0),.clk(gclk));
	jdff dff_A_Sy0nyQxk0_0(.dout(w_dff_A_HOiwcsfq9_0),.din(w_dff_A_Sy0nyQxk0_0),.clk(gclk));
	jdff dff_A_n3XMWM151_0(.dout(w_dff_A_Sy0nyQxk0_0),.din(w_dff_A_n3XMWM151_0),.clk(gclk));
	jdff dff_A_ceGG89cq8_0(.dout(w_dff_A_n3XMWM151_0),.din(w_dff_A_ceGG89cq8_0),.clk(gclk));
	jdff dff_A_uv1pBWGx9_0(.dout(w_dff_A_ceGG89cq8_0),.din(w_dff_A_uv1pBWGx9_0),.clk(gclk));
	jdff dff_A_Fnx7eK0y1_0(.dout(w_dff_A_uv1pBWGx9_0),.din(w_dff_A_Fnx7eK0y1_0),.clk(gclk));
	jdff dff_A_I3jfBtvS7_0(.dout(w_dff_A_Fnx7eK0y1_0),.din(w_dff_A_I3jfBtvS7_0),.clk(gclk));
	jdff dff_A_sqbawJ0Y8_0(.dout(w_dff_A_I3jfBtvS7_0),.din(w_dff_A_sqbawJ0Y8_0),.clk(gclk));
	jdff dff_A_ci3ckk8m1_0(.dout(w_dff_A_sqbawJ0Y8_0),.din(w_dff_A_ci3ckk8m1_0),.clk(gclk));
	jdff dff_A_lQLNx10j0_0(.dout(w_dff_A_ci3ckk8m1_0),.din(w_dff_A_lQLNx10j0_0),.clk(gclk));
	jdff dff_A_taRnpM5n2_0(.dout(w_dff_A_lQLNx10j0_0),.din(w_dff_A_taRnpM5n2_0),.clk(gclk));
	jdff dff_A_81OM5YjI4_0(.dout(w_dff_A_taRnpM5n2_0),.din(w_dff_A_81OM5YjI4_0),.clk(gclk));
	jdff dff_A_m3HysKyj2_0(.dout(w_dff_A_81OM5YjI4_0),.din(w_dff_A_m3HysKyj2_0),.clk(gclk));
	jdff dff_A_rkrxYc2d2_0(.dout(w_dff_A_m3HysKyj2_0),.din(w_dff_A_rkrxYc2d2_0),.clk(gclk));
	jdff dff_A_AQxbrSVC9_1(.dout(w_G4088_9[1]),.din(w_dff_A_AQxbrSVC9_1),.clk(gclk));
	jdff dff_A_onMi9TXx1_1(.dout(w_dff_A_AQxbrSVC9_1),.din(w_dff_A_onMi9TXx1_1),.clk(gclk));
	jdff dff_A_EpAJ3cIs1_1(.dout(w_dff_A_onMi9TXx1_1),.din(w_dff_A_EpAJ3cIs1_1),.clk(gclk));
	jdff dff_A_3i54SPcU4_1(.dout(w_dff_A_EpAJ3cIs1_1),.din(w_dff_A_3i54SPcU4_1),.clk(gclk));
	jdff dff_A_9N6E4uSX1_1(.dout(w_dff_A_3i54SPcU4_1),.din(w_dff_A_9N6E4uSX1_1),.clk(gclk));
	jdff dff_A_nxj1Y6cT6_1(.dout(w_dff_A_9N6E4uSX1_1),.din(w_dff_A_nxj1Y6cT6_1),.clk(gclk));
	jdff dff_A_uA12pxJ92_1(.dout(w_dff_A_nxj1Y6cT6_1),.din(w_dff_A_uA12pxJ92_1),.clk(gclk));
	jdff dff_A_ZY4mbvov9_1(.dout(w_G4087_1[1]),.din(w_dff_A_ZY4mbvov9_1),.clk(gclk));
	jdff dff_A_46c1UTu87_0(.dout(w_G4088_3[0]),.din(w_dff_A_46c1UTu87_0),.clk(gclk));
	jdff dff_A_l57HmlmH3_0(.dout(w_dff_A_46c1UTu87_0),.din(w_dff_A_l57HmlmH3_0),.clk(gclk));
	jdff dff_A_5POZ5v0y5_0(.dout(w_dff_A_l57HmlmH3_0),.din(w_dff_A_5POZ5v0y5_0),.clk(gclk));
	jdff dff_A_m7LijZU08_0(.dout(w_dff_A_5POZ5v0y5_0),.din(w_dff_A_m7LijZU08_0),.clk(gclk));
	jdff dff_A_KhHYVNol9_0(.dout(w_dff_A_m7LijZU08_0),.din(w_dff_A_KhHYVNol9_0),.clk(gclk));
	jdff dff_A_nHotHTxJ2_0(.dout(w_dff_A_KhHYVNol9_0),.din(w_dff_A_nHotHTxJ2_0),.clk(gclk));
	jdff dff_A_urAmzmBm2_0(.dout(w_dff_A_nHotHTxJ2_0),.din(w_dff_A_urAmzmBm2_0),.clk(gclk));
	jdff dff_A_w52yENHX9_0(.dout(w_dff_A_urAmzmBm2_0),.din(w_dff_A_w52yENHX9_0),.clk(gclk));
	jdff dff_A_yodGdyjF1_0(.dout(w_dff_A_w52yENHX9_0),.din(w_dff_A_yodGdyjF1_0),.clk(gclk));
	jdff dff_A_JgmYUvvq4_0(.dout(w_dff_A_yodGdyjF1_0),.din(w_dff_A_JgmYUvvq4_0),.clk(gclk));
	jdff dff_A_IjWZ0cjW0_0(.dout(w_dff_A_JgmYUvvq4_0),.din(w_dff_A_IjWZ0cjW0_0),.clk(gclk));
	jdff dff_A_G5IAFQDd9_0(.dout(w_dff_A_IjWZ0cjW0_0),.din(w_dff_A_G5IAFQDd9_0),.clk(gclk));
	jdff dff_A_pZgEnPBt3_0(.dout(w_dff_A_G5IAFQDd9_0),.din(w_dff_A_pZgEnPBt3_0),.clk(gclk));
	jdff dff_A_PdO99CxA0_0(.dout(w_dff_A_pZgEnPBt3_0),.din(w_dff_A_PdO99CxA0_0),.clk(gclk));
	jdff dff_A_BOkVioFP1_0(.dout(w_dff_A_PdO99CxA0_0),.din(w_dff_A_BOkVioFP1_0),.clk(gclk));
	jdff dff_A_P6qfhyQ55_0(.dout(w_dff_A_BOkVioFP1_0),.din(w_dff_A_P6qfhyQ55_0),.clk(gclk));
	jdff dff_A_g64oOjpf2_0(.dout(w_dff_A_P6qfhyQ55_0),.din(w_dff_A_g64oOjpf2_0),.clk(gclk));
	jdff dff_A_PlrVWtov6_0(.dout(w_dff_A_g64oOjpf2_0),.din(w_dff_A_PlrVWtov6_0),.clk(gclk));
	jdff dff_A_iPVAgh5r5_0(.dout(w_dff_A_PlrVWtov6_0),.din(w_dff_A_iPVAgh5r5_0),.clk(gclk));
	jdff dff_B_b2rcfOAo5_1(.din(n1688),.dout(w_dff_B_b2rcfOAo5_1),.clk(gclk));
	jdff dff_B_iJpBJpJC6_1(.din(w_dff_B_b2rcfOAo5_1),.dout(w_dff_B_iJpBJpJC6_1),.clk(gclk));
	jdff dff_B_umm4bBqh9_1(.din(w_dff_B_iJpBJpJC6_1),.dout(w_dff_B_umm4bBqh9_1),.clk(gclk));
	jdff dff_B_EuiMQ7PN3_1(.din(w_dff_B_umm4bBqh9_1),.dout(w_dff_B_EuiMQ7PN3_1),.clk(gclk));
	jdff dff_B_ob3ULvyY1_1(.din(w_dff_B_EuiMQ7PN3_1),.dout(w_dff_B_ob3ULvyY1_1),.clk(gclk));
	jdff dff_B_oaXQrTyF6_1(.din(w_dff_B_ob3ULvyY1_1),.dout(w_dff_B_oaXQrTyF6_1),.clk(gclk));
	jdff dff_B_zA3ZIGSj0_1(.din(w_dff_B_oaXQrTyF6_1),.dout(w_dff_B_zA3ZIGSj0_1),.clk(gclk));
	jdff dff_B_PXIRLwyN1_1(.din(w_dff_B_zA3ZIGSj0_1),.dout(w_dff_B_PXIRLwyN1_1),.clk(gclk));
	jdff dff_B_lXZpWuCN0_1(.din(w_dff_B_PXIRLwyN1_1),.dout(w_dff_B_lXZpWuCN0_1),.clk(gclk));
	jdff dff_B_TO98OCIr0_1(.din(w_dff_B_lXZpWuCN0_1),.dout(w_dff_B_TO98OCIr0_1),.clk(gclk));
	jdff dff_B_L3SOA6hu7_1(.din(w_dff_B_TO98OCIr0_1),.dout(w_dff_B_L3SOA6hu7_1),.clk(gclk));
	jdff dff_B_HUfmvg2j8_1(.din(w_dff_B_L3SOA6hu7_1),.dout(w_dff_B_HUfmvg2j8_1),.clk(gclk));
	jdff dff_B_zEHCLY6G9_1(.din(w_dff_B_HUfmvg2j8_1),.dout(w_dff_B_zEHCLY6G9_1),.clk(gclk));
	jdff dff_B_Dn1zFS835_1(.din(w_dff_B_zEHCLY6G9_1),.dout(w_dff_B_Dn1zFS835_1),.clk(gclk));
	jdff dff_B_za3APN9P7_1(.din(w_dff_B_Dn1zFS835_1),.dout(w_dff_B_za3APN9P7_1),.clk(gclk));
	jdff dff_B_tUVxwxxA9_1(.din(w_dff_B_za3APN9P7_1),.dout(w_dff_B_tUVxwxxA9_1),.clk(gclk));
	jdff dff_B_aBbydeJj2_1(.din(w_dff_B_tUVxwxxA9_1),.dout(w_dff_B_aBbydeJj2_1),.clk(gclk));
	jdff dff_B_bGSCQJIQ0_1(.din(w_dff_B_aBbydeJj2_1),.dout(w_dff_B_bGSCQJIQ0_1),.clk(gclk));
	jdff dff_B_mDpCqA5d6_1(.din(n1689),.dout(w_dff_B_mDpCqA5d6_1),.clk(gclk));
	jdff dff_B_nj8by4FA8_1(.din(w_dff_B_mDpCqA5d6_1),.dout(w_dff_B_nj8by4FA8_1),.clk(gclk));
	jdff dff_B_0X0GAI739_1(.din(w_dff_B_nj8by4FA8_1),.dout(w_dff_B_0X0GAI739_1),.clk(gclk));
	jdff dff_A_JmxG3i3X7_1(.dout(w_n854_1[1]),.din(w_dff_A_JmxG3i3X7_1),.clk(gclk));
	jdff dff_A_OpYYQD5b6_1(.dout(w_dff_A_JmxG3i3X7_1),.din(w_dff_A_OpYYQD5b6_1),.clk(gclk));
	jdff dff_A_aRJxquyA2_1(.dout(w_dff_A_OpYYQD5b6_1),.din(w_dff_A_aRJxquyA2_1),.clk(gclk));
	jdff dff_A_52sKUUFg7_1(.dout(w_dff_A_aRJxquyA2_1),.din(w_dff_A_52sKUUFg7_1),.clk(gclk));
	jdff dff_A_7hBvdyLN6_1(.dout(w_dff_A_52sKUUFg7_1),.din(w_dff_A_7hBvdyLN6_1),.clk(gclk));
	jdff dff_A_s0qnuZSx5_1(.dout(w_dff_A_7hBvdyLN6_1),.din(w_dff_A_s0qnuZSx5_1),.clk(gclk));
	jdff dff_A_Lu97yoc89_1(.dout(w_dff_A_s0qnuZSx5_1),.din(w_dff_A_Lu97yoc89_1),.clk(gclk));
	jdff dff_A_Lfa3XIpl8_1(.dout(w_dff_A_Lu97yoc89_1),.din(w_dff_A_Lfa3XIpl8_1),.clk(gclk));
	jdff dff_A_OzKf7yLM5_1(.dout(w_dff_A_Lfa3XIpl8_1),.din(w_dff_A_OzKf7yLM5_1),.clk(gclk));
	jdff dff_A_ZR5gk7BB6_1(.dout(w_dff_A_OzKf7yLM5_1),.din(w_dff_A_ZR5gk7BB6_1),.clk(gclk));
	jdff dff_A_SJBnhBHh9_1(.dout(w_dff_A_ZR5gk7BB6_1),.din(w_dff_A_SJBnhBHh9_1),.clk(gclk));
	jdff dff_A_TUOlpUU97_1(.dout(w_dff_A_SJBnhBHh9_1),.din(w_dff_A_TUOlpUU97_1),.clk(gclk));
	jdff dff_A_EaFBdXsk9_2(.dout(w_n854_1[2]),.din(w_dff_A_EaFBdXsk9_2),.clk(gclk));
	jdff dff_A_mkt2cZNu2_2(.dout(w_dff_A_EaFBdXsk9_2),.din(w_dff_A_mkt2cZNu2_2),.clk(gclk));
	jdff dff_A_kzgIon3V5_2(.dout(w_dff_A_mkt2cZNu2_2),.din(w_dff_A_kzgIon3V5_2),.clk(gclk));
	jdff dff_A_7c826gqM9_2(.dout(w_dff_A_kzgIon3V5_2),.din(w_dff_A_7c826gqM9_2),.clk(gclk));
	jdff dff_A_v26QQYFn9_2(.dout(w_dff_A_7c826gqM9_2),.din(w_dff_A_v26QQYFn9_2),.clk(gclk));
	jdff dff_A_w7FbCt0k0_2(.dout(w_dff_A_v26QQYFn9_2),.din(w_dff_A_w7FbCt0k0_2),.clk(gclk));
	jdff dff_A_rzEmcvym0_2(.dout(w_dff_A_w7FbCt0k0_2),.din(w_dff_A_rzEmcvym0_2),.clk(gclk));
	jdff dff_A_AU70l0BR0_2(.dout(w_dff_A_rzEmcvym0_2),.din(w_dff_A_AU70l0BR0_2),.clk(gclk));
	jdff dff_A_i0pT8b6p8_1(.dout(w_n854_0[1]),.din(w_dff_A_i0pT8b6p8_1),.clk(gclk));
	jdff dff_A_BNdz5W6v2_1(.dout(w_dff_A_i0pT8b6p8_1),.din(w_dff_A_BNdz5W6v2_1),.clk(gclk));
	jdff dff_A_K4876BO89_1(.dout(w_dff_A_BNdz5W6v2_1),.din(w_dff_A_K4876BO89_1),.clk(gclk));
	jdff dff_A_jZci6xpn7_1(.dout(w_dff_A_K4876BO89_1),.din(w_dff_A_jZci6xpn7_1),.clk(gclk));
	jdff dff_A_fYsXlsdV7_1(.dout(w_dff_A_jZci6xpn7_1),.din(w_dff_A_fYsXlsdV7_1),.clk(gclk));
	jdff dff_A_HyE5cwxc9_1(.dout(w_dff_A_fYsXlsdV7_1),.din(w_dff_A_HyE5cwxc9_1),.clk(gclk));
	jdff dff_A_FyeoVdrP6_2(.dout(w_n854_0[2]),.din(w_dff_A_FyeoVdrP6_2),.clk(gclk));
	jdff dff_A_iXrQXtt85_2(.dout(w_dff_A_FyeoVdrP6_2),.din(w_dff_A_iXrQXtt85_2),.clk(gclk));
	jdff dff_A_VhhiEz3N5_2(.dout(w_dff_A_iXrQXtt85_2),.din(w_dff_A_VhhiEz3N5_2),.clk(gclk));
	jdff dff_B_zaDwqqmF6_3(.din(n854),.dout(w_dff_B_zaDwqqmF6_3),.clk(gclk));
	jdff dff_B_wOClTlYS3_3(.din(w_dff_B_zaDwqqmF6_3),.dout(w_dff_B_wOClTlYS3_3),.clk(gclk));
	jdff dff_B_24cfXtf52_3(.din(w_dff_B_wOClTlYS3_3),.dout(w_dff_B_24cfXtf52_3),.clk(gclk));
	jdff dff_B_waseNjwI4_3(.din(w_dff_B_24cfXtf52_3),.dout(w_dff_B_waseNjwI4_3),.clk(gclk));
	jdff dff_B_DBVmso4B8_3(.din(w_dff_B_waseNjwI4_3),.dout(w_dff_B_DBVmso4B8_3),.clk(gclk));
	jdff dff_B_ywEgtm6v0_3(.din(w_dff_B_DBVmso4B8_3),.dout(w_dff_B_ywEgtm6v0_3),.clk(gclk));
	jdff dff_A_WrtBaxLL7_0(.dout(w_G4090_4[0]),.din(w_dff_A_WrtBaxLL7_0),.clk(gclk));
	jdff dff_B_u5pwc04z4_1(.din(n1685),.dout(w_dff_B_u5pwc04z4_1),.clk(gclk));
	jdff dff_B_pkcCmuYD8_1(.din(w_dff_B_u5pwc04z4_1),.dout(w_dff_B_pkcCmuYD8_1),.clk(gclk));
	jdff dff_A_udlUBLP06_0(.dout(w_n852_3[0]),.din(w_dff_A_udlUBLP06_0),.clk(gclk));
	jdff dff_A_vzChoUuX1_0(.dout(w_dff_A_udlUBLP06_0),.din(w_dff_A_vzChoUuX1_0),.clk(gclk));
	jdff dff_A_PcFUTzKt3_0(.dout(w_dff_A_vzChoUuX1_0),.din(w_dff_A_PcFUTzKt3_0),.clk(gclk));
	jdff dff_A_ow5hqszk7_0(.dout(w_dff_A_PcFUTzKt3_0),.din(w_dff_A_ow5hqszk7_0),.clk(gclk));
	jdff dff_A_kS82MclJ4_0(.dout(w_dff_A_ow5hqszk7_0),.din(w_dff_A_kS82MclJ4_0),.clk(gclk));
	jdff dff_A_7Dny0Fmu2_0(.dout(w_dff_A_kS82MclJ4_0),.din(w_dff_A_7Dny0Fmu2_0),.clk(gclk));
	jdff dff_A_pUE2wtYt5_0(.dout(w_dff_A_7Dny0Fmu2_0),.din(w_dff_A_pUE2wtYt5_0),.clk(gclk));
	jdff dff_A_MrGUDlWU7_0(.dout(w_dff_A_pUE2wtYt5_0),.din(w_dff_A_MrGUDlWU7_0),.clk(gclk));
	jdff dff_A_RXNtSKFm3_0(.dout(w_dff_A_MrGUDlWU7_0),.din(w_dff_A_RXNtSKFm3_0),.clk(gclk));
	jdff dff_A_bpOFpYJ53_0(.dout(w_dff_A_RXNtSKFm3_0),.din(w_dff_A_bpOFpYJ53_0),.clk(gclk));
	jdff dff_A_i6zAf3cG0_0(.dout(w_dff_A_bpOFpYJ53_0),.din(w_dff_A_i6zAf3cG0_0),.clk(gclk));
	jdff dff_A_yKf2mi5S0_0(.dout(w_dff_A_i6zAf3cG0_0),.din(w_dff_A_yKf2mi5S0_0),.clk(gclk));
	jdff dff_A_bJUARkVp5_0(.dout(w_dff_A_yKf2mi5S0_0),.din(w_dff_A_bJUARkVp5_0),.clk(gclk));
	jdff dff_A_mEVVDa5N0_0(.dout(w_dff_A_bJUARkVp5_0),.din(w_dff_A_mEVVDa5N0_0),.clk(gclk));
	jdff dff_A_uJPWIQjh3_0(.dout(w_dff_A_mEVVDa5N0_0),.din(w_dff_A_uJPWIQjh3_0),.clk(gclk));
	jdff dff_A_aOhPuqhi6_0(.dout(w_dff_A_uJPWIQjh3_0),.din(w_dff_A_aOhPuqhi6_0),.clk(gclk));
	jdff dff_A_dpglei4F4_1(.dout(w_G4089_9[1]),.din(w_dff_A_dpglei4F4_1),.clk(gclk));
	jdff dff_A_t0m4ID4x1_1(.dout(w_dff_A_dpglei4F4_1),.din(w_dff_A_t0m4ID4x1_1),.clk(gclk));
	jdff dff_A_2KOzwYRg4_1(.dout(w_dff_A_t0m4ID4x1_1),.din(w_dff_A_2KOzwYRg4_1),.clk(gclk));
	jdff dff_A_IZQsoj7U4_1(.dout(w_dff_A_2KOzwYRg4_1),.din(w_dff_A_IZQsoj7U4_1),.clk(gclk));
	jdff dff_A_p2ubC7BX0_1(.dout(w_dff_A_IZQsoj7U4_1),.din(w_dff_A_p2ubC7BX0_1),.clk(gclk));
	jdff dff_A_VaIEA5X51_1(.dout(w_dff_A_p2ubC7BX0_1),.din(w_dff_A_VaIEA5X51_1),.clk(gclk));
	jdff dff_A_HgcJxiAs8_1(.dout(w_dff_A_VaIEA5X51_1),.din(w_dff_A_HgcJxiAs8_1),.clk(gclk));
	jdff dff_B_FLJVpyGZ3_2(.din(G64),.dout(w_dff_B_FLJVpyGZ3_2),.clk(gclk));
	jdff dff_A_vnoqIWWT6_1(.dout(w_G4090_1[1]),.din(w_dff_A_vnoqIWWT6_1),.clk(gclk));
	jdff dff_A_pdrTJy1i8_0(.dout(w_G4089_3[0]),.din(w_dff_A_pdrTJy1i8_0),.clk(gclk));
	jdff dff_A_pRDjoIEm6_0(.dout(w_dff_A_pdrTJy1i8_0),.din(w_dff_A_pRDjoIEm6_0),.clk(gclk));
	jdff dff_A_8H1KD62R8_0(.dout(w_dff_A_pRDjoIEm6_0),.din(w_dff_A_8H1KD62R8_0),.clk(gclk));
	jdff dff_A_agSwbR1e5_0(.dout(w_dff_A_8H1KD62R8_0),.din(w_dff_A_agSwbR1e5_0),.clk(gclk));
	jdff dff_A_4sJq9ubV8_0(.dout(w_dff_A_agSwbR1e5_0),.din(w_dff_A_4sJq9ubV8_0),.clk(gclk));
	jdff dff_A_3kKFd0Ze5_0(.dout(w_dff_A_4sJq9ubV8_0),.din(w_dff_A_3kKFd0Ze5_0),.clk(gclk));
	jdff dff_A_n6YfRw1H9_0(.dout(w_dff_A_3kKFd0Ze5_0),.din(w_dff_A_n6YfRw1H9_0),.clk(gclk));
	jdff dff_A_fvRLohg12_0(.dout(w_dff_A_n6YfRw1H9_0),.din(w_dff_A_fvRLohg12_0),.clk(gclk));
	jdff dff_A_ptnRsuft4_0(.dout(w_dff_A_fvRLohg12_0),.din(w_dff_A_ptnRsuft4_0),.clk(gclk));
	jdff dff_A_8NSOpAOV3_0(.dout(w_dff_A_ptnRsuft4_0),.din(w_dff_A_8NSOpAOV3_0),.clk(gclk));
	jdff dff_A_wWmCWJnk6_0(.dout(w_dff_A_8NSOpAOV3_0),.din(w_dff_A_wWmCWJnk6_0),.clk(gclk));
	jdff dff_A_i1t2QG4h2_0(.dout(w_dff_A_wWmCWJnk6_0),.din(w_dff_A_i1t2QG4h2_0),.clk(gclk));
	jdff dff_A_WCnWyzAE5_0(.dout(w_dff_A_i1t2QG4h2_0),.din(w_dff_A_WCnWyzAE5_0),.clk(gclk));
	jdff dff_A_o44IDXQl3_0(.dout(w_dff_A_WCnWyzAE5_0),.din(w_dff_A_o44IDXQl3_0),.clk(gclk));
	jdff dff_A_AkHnZjDH1_0(.dout(w_dff_A_o44IDXQl3_0),.din(w_dff_A_AkHnZjDH1_0),.clk(gclk));
	jdff dff_A_2atQeOyk4_0(.dout(w_dff_A_AkHnZjDH1_0),.din(w_dff_A_2atQeOyk4_0),.clk(gclk));
	jdff dff_A_sdYBnwaJ0_0(.dout(w_dff_A_2atQeOyk4_0),.din(w_dff_A_sdYBnwaJ0_0),.clk(gclk));
	jdff dff_A_DjEUFzkF4_0(.dout(w_dff_A_sdYBnwaJ0_0),.din(w_dff_A_DjEUFzkF4_0),.clk(gclk));
	jdff dff_A_WJPfpayy3_0(.dout(w_dff_A_DjEUFzkF4_0),.din(w_dff_A_WJPfpayy3_0),.clk(gclk));
	jdff dff_B_pJffjcOQ2_1(.din(n1697),.dout(w_dff_B_pJffjcOQ2_1),.clk(gclk));
	jdff dff_B_xXhgzhoq6_1(.din(w_dff_B_pJffjcOQ2_1),.dout(w_dff_B_xXhgzhoq6_1),.clk(gclk));
	jdff dff_B_Poi6ZA9Y7_1(.din(w_dff_B_xXhgzhoq6_1),.dout(w_dff_B_Poi6ZA9Y7_1),.clk(gclk));
	jdff dff_B_hXHJsLcI2_1(.din(w_dff_B_Poi6ZA9Y7_1),.dout(w_dff_B_hXHJsLcI2_1),.clk(gclk));
	jdff dff_B_TsTuR1uN9_1(.din(w_dff_B_hXHJsLcI2_1),.dout(w_dff_B_TsTuR1uN9_1),.clk(gclk));
	jdff dff_B_SuyYcSTo5_1(.din(w_dff_B_TsTuR1uN9_1),.dout(w_dff_B_SuyYcSTo5_1),.clk(gclk));
	jdff dff_B_j5GPUGIl5_1(.din(w_dff_B_SuyYcSTo5_1),.dout(w_dff_B_j5GPUGIl5_1),.clk(gclk));
	jdff dff_B_Q8jC2qi76_1(.din(w_dff_B_j5GPUGIl5_1),.dout(w_dff_B_Q8jC2qi76_1),.clk(gclk));
	jdff dff_B_ABaEJwPX7_1(.din(w_dff_B_Q8jC2qi76_1),.dout(w_dff_B_ABaEJwPX7_1),.clk(gclk));
	jdff dff_B_MODYTMI39_1(.din(w_dff_B_ABaEJwPX7_1),.dout(w_dff_B_MODYTMI39_1),.clk(gclk));
	jdff dff_B_wmFzOJ4K7_1(.din(w_dff_B_MODYTMI39_1),.dout(w_dff_B_wmFzOJ4K7_1),.clk(gclk));
	jdff dff_B_ulVjxbAe7_1(.din(w_dff_B_wmFzOJ4K7_1),.dout(w_dff_B_ulVjxbAe7_1),.clk(gclk));
	jdff dff_B_PbDOvcpb8_1(.din(w_dff_B_ulVjxbAe7_1),.dout(w_dff_B_PbDOvcpb8_1),.clk(gclk));
	jdff dff_B_fi1EYCqG0_1(.din(w_dff_B_PbDOvcpb8_1),.dout(w_dff_B_fi1EYCqG0_1),.clk(gclk));
	jdff dff_B_TW288oSk7_1(.din(w_dff_B_fi1EYCqG0_1),.dout(w_dff_B_TW288oSk7_1),.clk(gclk));
	jdff dff_B_AaXn2NDy6_1(.din(w_dff_B_TW288oSk7_1),.dout(w_dff_B_AaXn2NDy6_1),.clk(gclk));
	jdff dff_B_mKkKryGu0_1(.din(w_dff_B_AaXn2NDy6_1),.dout(w_dff_B_mKkKryGu0_1),.clk(gclk));
	jdff dff_B_qEMVhYvC0_1(.din(w_dff_B_mKkKryGu0_1),.dout(w_dff_B_qEMVhYvC0_1),.clk(gclk));
	jdff dff_B_lF41FNti2_1(.din(n1700),.dout(w_dff_B_lF41FNti2_1),.clk(gclk));
	jdff dff_B_KCYizpgs9_1(.din(w_dff_B_lF41FNti2_1),.dout(w_dff_B_KCYizpgs9_1),.clk(gclk));
	jdff dff_B_Gnpx6ZxS1_1(.din(w_dff_B_KCYizpgs9_1),.dout(w_dff_B_Gnpx6ZxS1_1),.clk(gclk));
	jdff dff_B_WoAadTlh5_1(.din(w_dff_B_Gnpx6ZxS1_1),.dout(w_dff_B_WoAadTlh5_1),.clk(gclk));
	jdff dff_B_tO25t6dS4_1(.din(w_dff_B_WoAadTlh5_1),.dout(w_dff_B_tO25t6dS4_1),.clk(gclk));
	jdff dff_B_Ar6ZUzHm5_1(.din(w_dff_B_tO25t6dS4_1),.dout(w_dff_B_Ar6ZUzHm5_1),.clk(gclk));
	jdff dff_B_H7DX6pVw0_1(.din(w_dff_B_Ar6ZUzHm5_1),.dout(w_dff_B_H7DX6pVw0_1),.clk(gclk));
	jdff dff_B_YfBEjTHl2_1(.din(w_dff_B_H7DX6pVw0_1),.dout(w_dff_B_YfBEjTHl2_1),.clk(gclk));
	jdff dff_B_d66XZqqJ8_1(.din(w_dff_B_YfBEjTHl2_1),.dout(w_dff_B_d66XZqqJ8_1),.clk(gclk));
	jdff dff_B_ppgMSckT3_1(.din(w_dff_B_d66XZqqJ8_1),.dout(w_dff_B_ppgMSckT3_1),.clk(gclk));
	jdff dff_B_4n2AyCD48_1(.din(w_dff_B_ppgMSckT3_1),.dout(w_dff_B_4n2AyCD48_1),.clk(gclk));
	jdff dff_B_3hb8bEZZ3_1(.din(w_dff_B_4n2AyCD48_1),.dout(w_dff_B_3hb8bEZZ3_1),.clk(gclk));
	jdff dff_B_YBuJYGdY9_1(.din(w_dff_B_3hb8bEZZ3_1),.dout(w_dff_B_YBuJYGdY9_1),.clk(gclk));
	jdff dff_B_w0CSvFMJ9_1(.din(w_dff_B_YBuJYGdY9_1),.dout(w_dff_B_w0CSvFMJ9_1),.clk(gclk));
	jdff dff_B_PrC8srmz1_1(.din(w_dff_B_w0CSvFMJ9_1),.dout(w_dff_B_PrC8srmz1_1),.clk(gclk));
	jdff dff_B_nvqN5uz61_1(.din(w_dff_B_PrC8srmz1_1),.dout(w_dff_B_nvqN5uz61_1),.clk(gclk));
	jdff dff_B_2ioENHB65_1(.din(n1701),.dout(w_dff_B_2ioENHB65_1),.clk(gclk));
	jdff dff_B_EMUBajAW9_1(.din(w_dff_B_2ioENHB65_1),.dout(w_dff_B_EMUBajAW9_1),.clk(gclk));
	jdff dff_A_8xK8VXFh7_0(.dout(w_n993_4[0]),.din(w_dff_A_8xK8VXFh7_0),.clk(gclk));
	jdff dff_A_1aatv5mw9_0(.dout(w_dff_A_8xK8VXFh7_0),.din(w_dff_A_1aatv5mw9_0),.clk(gclk));
	jdff dff_A_puEjy21F4_0(.dout(w_dff_A_1aatv5mw9_0),.din(w_dff_A_puEjy21F4_0),.clk(gclk));
	jdff dff_A_UqERjw0i5_0(.dout(w_dff_A_puEjy21F4_0),.din(w_dff_A_UqERjw0i5_0),.clk(gclk));
	jdff dff_A_Q6NcDjzu2_0(.dout(w_dff_A_UqERjw0i5_0),.din(w_dff_A_Q6NcDjzu2_0),.clk(gclk));
	jdff dff_A_oQrl6rLs7_0(.dout(w_dff_A_Q6NcDjzu2_0),.din(w_dff_A_oQrl6rLs7_0),.clk(gclk));
	jdff dff_A_iULWfgfT4_0(.dout(w_dff_A_oQrl6rLs7_0),.din(w_dff_A_iULWfgfT4_0),.clk(gclk));
	jdff dff_A_gcXW73iw7_0(.dout(w_dff_A_iULWfgfT4_0),.din(w_dff_A_gcXW73iw7_0),.clk(gclk));
	jdff dff_A_XUX3r3iv1_0(.dout(w_dff_A_gcXW73iw7_0),.din(w_dff_A_XUX3r3iv1_0),.clk(gclk));
	jdff dff_A_VtkPEHmx9_0(.dout(w_dff_A_XUX3r3iv1_0),.din(w_dff_A_VtkPEHmx9_0),.clk(gclk));
	jdff dff_A_k9hWg1wo0_0(.dout(w_dff_A_VtkPEHmx9_0),.din(w_dff_A_k9hWg1wo0_0),.clk(gclk));
	jdff dff_A_YwEznwgY8_0(.dout(w_dff_A_k9hWg1wo0_0),.din(w_dff_A_YwEznwgY8_0),.clk(gclk));
	jdff dff_A_cRUsgrtb4_1(.dout(w_n993_4[1]),.din(w_dff_A_cRUsgrtb4_1),.clk(gclk));
	jdff dff_A_BuoCDXTF6_1(.dout(w_dff_A_cRUsgrtb4_1),.din(w_dff_A_BuoCDXTF6_1),.clk(gclk));
	jdff dff_A_oheE48JG9_1(.dout(w_dff_A_BuoCDXTF6_1),.din(w_dff_A_oheE48JG9_1),.clk(gclk));
	jdff dff_A_Oy5oOTlU2_1(.dout(w_dff_A_oheE48JG9_1),.din(w_dff_A_Oy5oOTlU2_1),.clk(gclk));
	jdff dff_A_1pa8uRPx7_1(.dout(w_dff_A_Oy5oOTlU2_1),.din(w_dff_A_1pa8uRPx7_1),.clk(gclk));
	jdff dff_A_hh5YWipl6_1(.dout(w_dff_A_1pa8uRPx7_1),.din(w_dff_A_hh5YWipl6_1),.clk(gclk));
	jdff dff_A_GOfz4csY9_1(.dout(w_dff_A_hh5YWipl6_1),.din(w_dff_A_GOfz4csY9_1),.clk(gclk));
	jdff dff_A_jMuMy8Wk7_1(.dout(w_dff_A_GOfz4csY9_1),.din(w_dff_A_jMuMy8Wk7_1),.clk(gclk));
	jdff dff_A_hmqJmvhe9_1(.dout(w_dff_A_jMuMy8Wk7_1),.din(w_dff_A_hmqJmvhe9_1),.clk(gclk));
	jdff dff_A_bxFPa8u93_1(.dout(w_n993_1[1]),.din(w_dff_A_bxFPa8u93_1),.clk(gclk));
	jdff dff_A_WfuOkAOV8_1(.dout(w_dff_A_bxFPa8u93_1),.din(w_dff_A_WfuOkAOV8_1),.clk(gclk));
	jdff dff_A_iIvhlGgr9_1(.dout(w_dff_A_WfuOkAOV8_1),.din(w_dff_A_iIvhlGgr9_1),.clk(gclk));
	jdff dff_A_6QchqKpk5_1(.dout(w_dff_A_iIvhlGgr9_1),.din(w_dff_A_6QchqKpk5_1),.clk(gclk));
	jdff dff_A_dC3enEGa0_1(.dout(w_dff_A_6QchqKpk5_1),.din(w_dff_A_dC3enEGa0_1),.clk(gclk));
	jdff dff_A_HqZ9htgT0_1(.dout(w_dff_A_dC3enEGa0_1),.din(w_dff_A_HqZ9htgT0_1),.clk(gclk));
	jdff dff_A_CfthQPG70_1(.dout(w_dff_A_HqZ9htgT0_1),.din(w_dff_A_CfthQPG70_1),.clk(gclk));
	jdff dff_A_cObrOEkK4_1(.dout(w_dff_A_CfthQPG70_1),.din(w_dff_A_cObrOEkK4_1),.clk(gclk));
	jdff dff_A_09DbJUja3_1(.dout(w_dff_A_cObrOEkK4_1),.din(w_dff_A_09DbJUja3_1),.clk(gclk));
	jdff dff_A_4dLxQPcd1_1(.dout(w_dff_A_09DbJUja3_1),.din(w_dff_A_4dLxQPcd1_1),.clk(gclk));
	jdff dff_A_DUsB57ym2_1(.dout(w_dff_A_4dLxQPcd1_1),.din(w_dff_A_DUsB57ym2_1),.clk(gclk));
	jdff dff_A_GYmrlpJv3_1(.dout(w_dff_A_DUsB57ym2_1),.din(w_dff_A_GYmrlpJv3_1),.clk(gclk));
	jdff dff_A_fffNOiRE9_1(.dout(w_dff_A_GYmrlpJv3_1),.din(w_dff_A_fffNOiRE9_1),.clk(gclk));
	jdff dff_A_egOg8bec8_1(.dout(w_dff_A_fffNOiRE9_1),.din(w_dff_A_egOg8bec8_1),.clk(gclk));
	jdff dff_A_OM7OUMoI5_1(.dout(w_dff_A_egOg8bec8_1),.din(w_dff_A_OM7OUMoI5_1),.clk(gclk));
	jdff dff_A_qUsJx8Qp0_1(.dout(w_dff_A_OM7OUMoI5_1),.din(w_dff_A_qUsJx8Qp0_1),.clk(gclk));
	jdff dff_A_sIofJAnO1_1(.dout(w_dff_A_qUsJx8Qp0_1),.din(w_dff_A_sIofJAnO1_1),.clk(gclk));
	jdff dff_A_bMj26oXv2_2(.dout(w_n993_1[2]),.din(w_dff_A_bMj26oXv2_2),.clk(gclk));
	jdff dff_A_gfaXRvDY4_2(.dout(w_dff_A_bMj26oXv2_2),.din(w_dff_A_gfaXRvDY4_2),.clk(gclk));
	jdff dff_A_d5ywrFJG8_2(.dout(w_dff_A_gfaXRvDY4_2),.din(w_dff_A_d5ywrFJG8_2),.clk(gclk));
	jdff dff_A_aKHTaF592_2(.dout(w_dff_A_d5ywrFJG8_2),.din(w_dff_A_aKHTaF592_2),.clk(gclk));
	jdff dff_A_2HjCF51g9_2(.dout(w_dff_A_aKHTaF592_2),.din(w_dff_A_2HjCF51g9_2),.clk(gclk));
	jdff dff_A_ADMGUHmx8_2(.dout(w_dff_A_2HjCF51g9_2),.din(w_dff_A_ADMGUHmx8_2),.clk(gclk));
	jdff dff_A_cnw3HkUX6_2(.dout(w_dff_A_ADMGUHmx8_2),.din(w_dff_A_cnw3HkUX6_2),.clk(gclk));
	jdff dff_A_TcitEqyr9_2(.dout(w_dff_A_cnw3HkUX6_2),.din(w_dff_A_TcitEqyr9_2),.clk(gclk));
	jdff dff_A_wxwLr7ba7_2(.dout(w_dff_A_TcitEqyr9_2),.din(w_dff_A_wxwLr7ba7_2),.clk(gclk));
	jdff dff_A_VpcbP0Cs6_2(.dout(w_dff_A_wxwLr7ba7_2),.din(w_dff_A_VpcbP0Cs6_2),.clk(gclk));
	jdff dff_A_4vJo3Nhw6_2(.dout(w_dff_A_VpcbP0Cs6_2),.din(w_dff_A_4vJo3Nhw6_2),.clk(gclk));
	jdff dff_A_6sIYz1BS8_2(.dout(w_dff_A_4vJo3Nhw6_2),.din(w_dff_A_6sIYz1BS8_2),.clk(gclk));
	jdff dff_A_xU9ffot83_2(.dout(w_dff_A_6sIYz1BS8_2),.din(w_dff_A_xU9ffot83_2),.clk(gclk));
	jdff dff_A_iJo7wsB24_2(.dout(w_dff_A_xU9ffot83_2),.din(w_dff_A_iJo7wsB24_2),.clk(gclk));
	jdff dff_A_qnFqvISH0_1(.dout(w_n993_0[1]),.din(w_dff_A_qnFqvISH0_1),.clk(gclk));
	jdff dff_A_74tlJx2G5_1(.dout(w_dff_A_qnFqvISH0_1),.din(w_dff_A_74tlJx2G5_1),.clk(gclk));
	jdff dff_A_Q37oWraE4_1(.dout(w_dff_A_74tlJx2G5_1),.din(w_dff_A_Q37oWraE4_1),.clk(gclk));
	jdff dff_A_3mmU56vm8_1(.dout(w_dff_A_Q37oWraE4_1),.din(w_dff_A_3mmU56vm8_1),.clk(gclk));
	jdff dff_A_LITqAKQa6_1(.dout(w_dff_A_3mmU56vm8_1),.din(w_dff_A_LITqAKQa6_1),.clk(gclk));
	jdff dff_A_h44018j13_1(.dout(w_dff_A_LITqAKQa6_1),.din(w_dff_A_h44018j13_1),.clk(gclk));
	jdff dff_A_KOXHWqVg0_1(.dout(w_dff_A_h44018j13_1),.din(w_dff_A_KOXHWqVg0_1),.clk(gclk));
	jdff dff_A_TXcFZWv89_1(.dout(w_dff_A_KOXHWqVg0_1),.din(w_dff_A_TXcFZWv89_1),.clk(gclk));
	jdff dff_A_KU4MEAzF4_1(.dout(w_dff_A_TXcFZWv89_1),.din(w_dff_A_KU4MEAzF4_1),.clk(gclk));
	jdff dff_A_94TvaCZy6_1(.dout(w_dff_A_KU4MEAzF4_1),.din(w_dff_A_94TvaCZy6_1),.clk(gclk));
	jdff dff_A_UTp8sruD6_1(.dout(w_dff_A_94TvaCZy6_1),.din(w_dff_A_UTp8sruD6_1),.clk(gclk));
	jdff dff_A_qPTMqRIg5_1(.dout(w_dff_A_UTp8sruD6_1),.din(w_dff_A_qPTMqRIg5_1),.clk(gclk));
	jdff dff_A_IAF5Qtnl9_1(.dout(w_dff_A_qPTMqRIg5_1),.din(w_dff_A_IAF5Qtnl9_1),.clk(gclk));
	jdff dff_A_Ocg1H20t9_2(.dout(w_n993_0[2]),.din(w_dff_A_Ocg1H20t9_2),.clk(gclk));
	jdff dff_A_GLKjOtYb7_2(.dout(w_dff_A_Ocg1H20t9_2),.din(w_dff_A_GLKjOtYb7_2),.clk(gclk));
	jdff dff_A_n81TeKAl8_2(.dout(w_dff_A_GLKjOtYb7_2),.din(w_dff_A_n81TeKAl8_2),.clk(gclk));
	jdff dff_A_ViFLau3t7_2(.dout(w_dff_A_n81TeKAl8_2),.din(w_dff_A_ViFLau3t7_2),.clk(gclk));
	jdff dff_A_2I9S8XQp6_2(.dout(w_dff_A_ViFLau3t7_2),.din(w_dff_A_2I9S8XQp6_2),.clk(gclk));
	jdff dff_A_C3OqboqI7_2(.dout(w_dff_A_2I9S8XQp6_2),.din(w_dff_A_C3OqboqI7_2),.clk(gclk));
	jdff dff_A_VvoNm4nn9_2(.dout(w_dff_A_C3OqboqI7_2),.din(w_dff_A_VvoNm4nn9_2),.clk(gclk));
	jdff dff_A_0O2kpQdZ4_2(.dout(w_dff_A_VvoNm4nn9_2),.din(w_dff_A_0O2kpQdZ4_2),.clk(gclk));
	jdff dff_A_8376GmCA9_2(.dout(w_dff_A_0O2kpQdZ4_2),.din(w_dff_A_8376GmCA9_2),.clk(gclk));
	jdff dff_A_XlDx9OSS6_1(.dout(w_G1690_1[1]),.din(w_dff_A_XlDx9OSS6_1),.clk(gclk));
	jdff dff_A_xkrDxope0_1(.dout(w_G1690_0[1]),.din(w_dff_A_xkrDxope0_1),.clk(gclk));
	jdff dff_A_nGqoYRDg4_1(.dout(w_dff_A_xkrDxope0_1),.din(w_dff_A_nGqoYRDg4_1),.clk(gclk));
	jdff dff_A_YgZ58kRh5_1(.dout(w_dff_A_nGqoYRDg4_1),.din(w_dff_A_YgZ58kRh5_1),.clk(gclk));
	jdff dff_A_7LyVNPUy3_1(.dout(w_dff_A_YgZ58kRh5_1),.din(w_dff_A_7LyVNPUy3_1),.clk(gclk));
	jdff dff_A_jECS5YH59_1(.dout(w_dff_A_7LyVNPUy3_1),.din(w_dff_A_jECS5YH59_1),.clk(gclk));
	jdff dff_A_LnrAmqGP8_1(.dout(w_dff_A_jECS5YH59_1),.din(w_dff_A_LnrAmqGP8_1),.clk(gclk));
	jdff dff_A_dzJXTCCT9_1(.dout(w_dff_A_LnrAmqGP8_1),.din(w_dff_A_dzJXTCCT9_1),.clk(gclk));
	jdff dff_A_f0rXsL5M1_1(.dout(w_dff_A_dzJXTCCT9_1),.din(w_dff_A_f0rXsL5M1_1),.clk(gclk));
	jdff dff_A_a728PDv13_1(.dout(w_dff_A_f0rXsL5M1_1),.din(w_dff_A_a728PDv13_1),.clk(gclk));
	jdff dff_A_ttFflHNJ8_1(.dout(w_dff_A_a728PDv13_1),.din(w_dff_A_ttFflHNJ8_1),.clk(gclk));
	jdff dff_A_n4lnK1VF4_1(.dout(w_dff_A_ttFflHNJ8_1),.din(w_dff_A_n4lnK1VF4_1),.clk(gclk));
	jdff dff_A_x75IVeFP2_1(.dout(w_dff_A_n4lnK1VF4_1),.din(w_dff_A_x75IVeFP2_1),.clk(gclk));
	jdff dff_A_9kvR0RHU7_1(.dout(w_dff_A_x75IVeFP2_1),.din(w_dff_A_9kvR0RHU7_1),.clk(gclk));
	jdff dff_A_Ub4t46gV0_1(.dout(w_dff_A_9kvR0RHU7_1),.din(w_dff_A_Ub4t46gV0_1),.clk(gclk));
	jdff dff_A_G8NnnIVa3_1(.dout(w_dff_A_Ub4t46gV0_1),.din(w_dff_A_G8NnnIVa3_1),.clk(gclk));
	jdff dff_A_JptWlgdZ2_1(.dout(w_dff_A_G8NnnIVa3_1),.din(w_dff_A_JptWlgdZ2_1),.clk(gclk));
	jdff dff_A_OZ4fZ4xv6_1(.dout(w_dff_A_JptWlgdZ2_1),.din(w_dff_A_OZ4fZ4xv6_1),.clk(gclk));
	jdff dff_A_5eaAx21E9_1(.dout(w_dff_A_OZ4fZ4xv6_1),.din(w_dff_A_5eaAx21E9_1),.clk(gclk));
	jdff dff_A_f405pS0G7_1(.dout(w_dff_A_5eaAx21E9_1),.din(w_dff_A_f405pS0G7_1),.clk(gclk));
	jdff dff_A_7h0amuuZ1_0(.dout(w_G1689_1[0]),.din(w_dff_A_7h0amuuZ1_0),.clk(gclk));
	jdff dff_A_o5wOCgQ61_0(.dout(w_dff_A_7h0amuuZ1_0),.din(w_dff_A_o5wOCgQ61_0),.clk(gclk));
	jdff dff_A_8ybaW9IF6_0(.dout(w_dff_A_o5wOCgQ61_0),.din(w_dff_A_8ybaW9IF6_0),.clk(gclk));
	jdff dff_A_0ChQ87o71_0(.dout(w_dff_A_8ybaW9IF6_0),.din(w_dff_A_0ChQ87o71_0),.clk(gclk));
	jdff dff_A_LbZ03N6A8_0(.dout(w_dff_A_0ChQ87o71_0),.din(w_dff_A_LbZ03N6A8_0),.clk(gclk));
	jdff dff_A_vbvg9F0Z0_0(.dout(w_dff_A_LbZ03N6A8_0),.din(w_dff_A_vbvg9F0Z0_0),.clk(gclk));
	jdff dff_A_yn9tlmaF7_0(.dout(w_dff_A_vbvg9F0Z0_0),.din(w_dff_A_yn9tlmaF7_0),.clk(gclk));
	jdff dff_A_H5kKxkqm6_2(.dout(w_G1689_1[2]),.din(w_dff_A_H5kKxkqm6_2),.clk(gclk));
	jdff dff_A_vItqtTeF6_2(.dout(w_dff_A_H5kKxkqm6_2),.din(w_dff_A_vItqtTeF6_2),.clk(gclk));
	jdff dff_A_Vbwb1EMG9_2(.dout(w_dff_A_vItqtTeF6_2),.din(w_dff_A_Vbwb1EMG9_2),.clk(gclk));
	jdff dff_A_w9MX6vb47_2(.dout(w_dff_A_Vbwb1EMG9_2),.din(w_dff_A_w9MX6vb47_2),.clk(gclk));
	jdff dff_A_Od3aWPll0_2(.dout(w_dff_A_w9MX6vb47_2),.din(w_dff_A_Od3aWPll0_2),.clk(gclk));
	jdff dff_A_xvTRKp3k9_2(.dout(w_dff_A_Od3aWPll0_2),.din(w_dff_A_xvTRKp3k9_2),.clk(gclk));
	jdff dff_A_XJgAsCsE9_2(.dout(w_dff_A_xvTRKp3k9_2),.din(w_dff_A_XJgAsCsE9_2),.clk(gclk));
	jdff dff_A_5R0xYeGe7_2(.dout(w_dff_A_XJgAsCsE9_2),.din(w_dff_A_5R0xYeGe7_2),.clk(gclk));
	jdff dff_A_J62SNFk35_2(.dout(w_dff_A_5R0xYeGe7_2),.din(w_dff_A_J62SNFk35_2),.clk(gclk));
	jdff dff_A_Eh8SxKZM5_2(.dout(w_dff_A_J62SNFk35_2),.din(w_dff_A_Eh8SxKZM5_2),.clk(gclk));
	jdff dff_A_ySTgQNO37_2(.dout(w_dff_A_Eh8SxKZM5_2),.din(w_dff_A_ySTgQNO37_2),.clk(gclk));
	jdff dff_A_KK8seJc28_2(.dout(w_dff_A_ySTgQNO37_2),.din(w_dff_A_KK8seJc28_2),.clk(gclk));
	jdff dff_A_9Y6mym4t4_2(.dout(w_dff_A_KK8seJc28_2),.din(w_dff_A_9Y6mym4t4_2),.clk(gclk));
	jdff dff_A_V4SPeXWY4_2(.dout(w_dff_A_9Y6mym4t4_2),.din(w_dff_A_V4SPeXWY4_2),.clk(gclk));
	jdff dff_A_eKCvZG224_2(.dout(w_dff_A_V4SPeXWY4_2),.din(w_dff_A_eKCvZG224_2),.clk(gclk));
	jdff dff_A_ZGEwQbOp8_2(.dout(w_dff_A_eKCvZG224_2),.din(w_dff_A_ZGEwQbOp8_2),.clk(gclk));
	jdff dff_A_YjWwCsyN2_1(.dout(w_G1689_0[1]),.din(w_dff_A_YjWwCsyN2_1),.clk(gclk));
	jdff dff_A_amHV6v8B9_1(.dout(w_dff_A_YjWwCsyN2_1),.din(w_dff_A_amHV6v8B9_1),.clk(gclk));
	jdff dff_A_avyApZ9t5_1(.dout(w_dff_A_amHV6v8B9_1),.din(w_dff_A_avyApZ9t5_1),.clk(gclk));
	jdff dff_A_uzOaPsZv1_1(.dout(w_dff_A_avyApZ9t5_1),.din(w_dff_A_uzOaPsZv1_1),.clk(gclk));
	jdff dff_A_qKu5EPsF5_1(.dout(w_dff_A_uzOaPsZv1_1),.din(w_dff_A_qKu5EPsF5_1),.clk(gclk));
	jdff dff_A_wNrZFBS95_1(.dout(w_dff_A_qKu5EPsF5_1),.din(w_dff_A_wNrZFBS95_1),.clk(gclk));
	jdff dff_A_XVpHqNjm7_1(.dout(w_dff_A_wNrZFBS95_1),.din(w_dff_A_XVpHqNjm7_1),.clk(gclk));
	jdff dff_A_Fy9rEV3l5_1(.dout(w_dff_A_XVpHqNjm7_1),.din(w_dff_A_Fy9rEV3l5_1),.clk(gclk));
	jdff dff_A_wjoPMRhT6_1(.dout(w_dff_A_Fy9rEV3l5_1),.din(w_dff_A_wjoPMRhT6_1),.clk(gclk));
	jdff dff_A_nLoa28D20_1(.dout(w_dff_A_wjoPMRhT6_1),.din(w_dff_A_nLoa28D20_1),.clk(gclk));
	jdff dff_A_KhwDJsyE7_1(.dout(w_dff_A_nLoa28D20_1),.din(w_dff_A_KhwDJsyE7_1),.clk(gclk));
	jdff dff_A_QXu7rwtx6_1(.dout(w_dff_A_KhwDJsyE7_1),.din(w_dff_A_QXu7rwtx6_1),.clk(gclk));
	jdff dff_A_Cg8fNTzH5_2(.dout(w_G1689_0[2]),.din(w_dff_A_Cg8fNTzH5_2),.clk(gclk));
	jdff dff_A_duePGjtb9_2(.dout(w_dff_A_Cg8fNTzH5_2),.din(w_dff_A_duePGjtb9_2),.clk(gclk));
	jdff dff_A_BoSfbFG50_2(.dout(w_dff_A_duePGjtb9_2),.din(w_dff_A_BoSfbFG50_2),.clk(gclk));
	jdff dff_A_yxkdMpGz0_2(.dout(w_dff_A_BoSfbFG50_2),.din(w_dff_A_yxkdMpGz0_2),.clk(gclk));
	jdff dff_A_FzKve4SU4_2(.dout(w_dff_A_yxkdMpGz0_2),.din(w_dff_A_FzKve4SU4_2),.clk(gclk));
	jdff dff_A_Px1p9vNX5_2(.dout(w_dff_A_FzKve4SU4_2),.din(w_dff_A_Px1p9vNX5_2),.clk(gclk));
	jdff dff_A_77eWdI954_2(.dout(w_dff_A_Px1p9vNX5_2),.din(w_dff_A_77eWdI954_2),.clk(gclk));
	jdff dff_A_HYv2veyb9_2(.dout(w_dff_A_77eWdI954_2),.din(w_dff_A_HYv2veyb9_2),.clk(gclk));
	jdff dff_A_vbkxWPKJ6_2(.dout(w_dff_A_HYv2veyb9_2),.din(w_dff_A_vbkxWPKJ6_2),.clk(gclk));
	jdff dff_B_g1NZdqsi7_1(.din(n1709),.dout(w_dff_B_g1NZdqsi7_1),.clk(gclk));
	jdff dff_B_T4yHuf3p1_1(.din(w_dff_B_g1NZdqsi7_1),.dout(w_dff_B_T4yHuf3p1_1),.clk(gclk));
	jdff dff_B_B4sIOW8K3_1(.din(w_dff_B_T4yHuf3p1_1),.dout(w_dff_B_B4sIOW8K3_1),.clk(gclk));
	jdff dff_B_TTFgYehI2_1(.din(w_dff_B_B4sIOW8K3_1),.dout(w_dff_B_TTFgYehI2_1),.clk(gclk));
	jdff dff_B_rcFwh1Hh7_1(.din(w_dff_B_TTFgYehI2_1),.dout(w_dff_B_rcFwh1Hh7_1),.clk(gclk));
	jdff dff_B_RS0J7QR09_1(.din(w_dff_B_rcFwh1Hh7_1),.dout(w_dff_B_RS0J7QR09_1),.clk(gclk));
	jdff dff_B_JslYyxcs4_1(.din(w_dff_B_RS0J7QR09_1),.dout(w_dff_B_JslYyxcs4_1),.clk(gclk));
	jdff dff_B_YOdUTLAu9_1(.din(w_dff_B_JslYyxcs4_1),.dout(w_dff_B_YOdUTLAu9_1),.clk(gclk));
	jdff dff_B_vxD1Olrk3_1(.din(w_dff_B_YOdUTLAu9_1),.dout(w_dff_B_vxD1Olrk3_1),.clk(gclk));
	jdff dff_B_kCsAirVz0_1(.din(w_dff_B_vxD1Olrk3_1),.dout(w_dff_B_kCsAirVz0_1),.clk(gclk));
	jdff dff_B_zY7v3CCW5_1(.din(w_dff_B_kCsAirVz0_1),.dout(w_dff_B_zY7v3CCW5_1),.clk(gclk));
	jdff dff_B_wHJSwFaZ5_1(.din(w_dff_B_zY7v3CCW5_1),.dout(w_dff_B_wHJSwFaZ5_1),.clk(gclk));
	jdff dff_B_CAgiRPfG3_1(.din(w_dff_B_wHJSwFaZ5_1),.dout(w_dff_B_CAgiRPfG3_1),.clk(gclk));
	jdff dff_B_LhugXMuJ7_1(.din(w_dff_B_CAgiRPfG3_1),.dout(w_dff_B_LhugXMuJ7_1),.clk(gclk));
	jdff dff_B_PJTbO05R6_1(.din(w_dff_B_LhugXMuJ7_1),.dout(w_dff_B_PJTbO05R6_1),.clk(gclk));
	jdff dff_B_POLCdHC48_1(.din(w_dff_B_PJTbO05R6_1),.dout(w_dff_B_POLCdHC48_1),.clk(gclk));
	jdff dff_B_yM3NqG9g3_1(.din(w_dff_B_POLCdHC48_1),.dout(w_dff_B_yM3NqG9g3_1),.clk(gclk));
	jdff dff_B_O7Z1AKZ68_1(.din(w_dff_B_yM3NqG9g3_1),.dout(w_dff_B_O7Z1AKZ68_1),.clk(gclk));
	jdff dff_B_lb5dKOg98_1(.din(n1711),.dout(w_dff_B_lb5dKOg98_1),.clk(gclk));
	jdff dff_B_O5E94j3c4_1(.din(w_dff_B_lb5dKOg98_1),.dout(w_dff_B_O5E94j3c4_1),.clk(gclk));
	jdff dff_B_jXMyg2c55_1(.din(w_dff_B_O5E94j3c4_1),.dout(w_dff_B_jXMyg2c55_1),.clk(gclk));
	jdff dff_B_R1Wkhd6v8_1(.din(w_dff_B_jXMyg2c55_1),.dout(w_dff_B_R1Wkhd6v8_1),.clk(gclk));
	jdff dff_B_1X07Wmza9_1(.din(w_dff_B_R1Wkhd6v8_1),.dout(w_dff_B_1X07Wmza9_1),.clk(gclk));
	jdff dff_B_hlgieTYN3_1(.din(w_dff_B_1X07Wmza9_1),.dout(w_dff_B_hlgieTYN3_1),.clk(gclk));
	jdff dff_B_buQdeXio7_1(.din(w_dff_B_hlgieTYN3_1),.dout(w_dff_B_buQdeXio7_1),.clk(gclk));
	jdff dff_B_y5vdR8xS0_1(.din(w_dff_B_buQdeXio7_1),.dout(w_dff_B_y5vdR8xS0_1),.clk(gclk));
	jdff dff_B_uz9elGk93_1(.din(w_dff_B_y5vdR8xS0_1),.dout(w_dff_B_uz9elGk93_1),.clk(gclk));
	jdff dff_B_sOcVv01b4_1(.din(w_dff_B_uz9elGk93_1),.dout(w_dff_B_sOcVv01b4_1),.clk(gclk));
	jdff dff_B_uCZ8kTj63_1(.din(w_dff_B_sOcVv01b4_1),.dout(w_dff_B_uCZ8kTj63_1),.clk(gclk));
	jdff dff_B_7o671Esm1_1(.din(w_dff_B_uCZ8kTj63_1),.dout(w_dff_B_7o671Esm1_1),.clk(gclk));
	jdff dff_B_ofgYCHXe7_1(.din(w_dff_B_7o671Esm1_1),.dout(w_dff_B_ofgYCHXe7_1),.clk(gclk));
	jdff dff_B_pdIoJ7S96_1(.din(w_dff_B_ofgYCHXe7_1),.dout(w_dff_B_pdIoJ7S96_1),.clk(gclk));
	jdff dff_B_7MPljmG90_1(.din(w_dff_B_pdIoJ7S96_1),.dout(w_dff_B_7MPljmG90_1),.clk(gclk));
	jdff dff_B_u18zMVPH2_1(.din(w_dff_B_7MPljmG90_1),.dout(w_dff_B_u18zMVPH2_1),.clk(gclk));
	jdff dff_B_0598kKp94_1(.din(n1712),.dout(w_dff_B_0598kKp94_1),.clk(gclk));
	jdff dff_B_hGr6wSUJ7_1(.din(w_dff_B_0598kKp94_1),.dout(w_dff_B_hGr6wSUJ7_1),.clk(gclk));
	jdff dff_B_fPissgFc5_0(.din(n1678),.dout(w_dff_B_fPissgFc5_0),.clk(gclk));
	jdff dff_B_TFlZORKh3_0(.din(w_dff_B_fPissgFc5_0),.dout(w_dff_B_TFlZORKh3_0),.clk(gclk));
	jdff dff_B_RY666wF85_0(.din(w_dff_B_TFlZORKh3_0),.dout(w_dff_B_RY666wF85_0),.clk(gclk));
	jdff dff_B_7dnT8Qwg9_0(.din(w_dff_B_RY666wF85_0),.dout(w_dff_B_7dnT8Qwg9_0),.clk(gclk));
	jdff dff_B_g6AtUCyW1_0(.din(w_dff_B_7dnT8Qwg9_0),.dout(w_dff_B_g6AtUCyW1_0),.clk(gclk));
	jdff dff_B_cloTSarb4_0(.din(w_dff_B_g6AtUCyW1_0),.dout(w_dff_B_cloTSarb4_0),.clk(gclk));
	jdff dff_B_r29TzAEK4_0(.din(w_dff_B_cloTSarb4_0),.dout(w_dff_B_r29TzAEK4_0),.clk(gclk));
	jdff dff_B_YvNukTC68_0(.din(w_dff_B_r29TzAEK4_0),.dout(w_dff_B_YvNukTC68_0),.clk(gclk));
	jdff dff_B_0dkMnsUl1_0(.din(w_dff_B_YvNukTC68_0),.dout(w_dff_B_0dkMnsUl1_0),.clk(gclk));
	jdff dff_B_RHNi9xVM6_0(.din(w_dff_B_0dkMnsUl1_0),.dout(w_dff_B_RHNi9xVM6_0),.clk(gclk));
	jdff dff_B_xPLCufXR0_0(.din(w_dff_B_RHNi9xVM6_0),.dout(w_dff_B_xPLCufXR0_0),.clk(gclk));
	jdff dff_B_eSl6CPWI9_0(.din(w_dff_B_xPLCufXR0_0),.dout(w_dff_B_eSl6CPWI9_0),.clk(gclk));
	jdff dff_B_gk2FnGnp0_0(.din(w_dff_B_eSl6CPWI9_0),.dout(w_dff_B_gk2FnGnp0_0),.clk(gclk));
	jdff dff_B_vNEaLbEW9_0(.din(w_dff_B_gk2FnGnp0_0),.dout(w_dff_B_vNEaLbEW9_0),.clk(gclk));
	jdff dff_B_LR7OJ1I74_0(.din(w_dff_B_vNEaLbEW9_0),.dout(w_dff_B_LR7OJ1I74_0),.clk(gclk));
	jdff dff_B_DjlpOAtG3_0(.din(n1501),.dout(w_dff_B_DjlpOAtG3_0),.clk(gclk));
	jdff dff_B_hV5agPxn8_0(.din(w_dff_B_DjlpOAtG3_0),.dout(w_dff_B_hV5agPxn8_0),.clk(gclk));
	jdff dff_B_QZw4TMhB7_0(.din(w_dff_B_hV5agPxn8_0),.dout(w_dff_B_QZw4TMhB7_0),.clk(gclk));
	jdff dff_B_VkeaUpgj9_0(.din(w_dff_B_QZw4TMhB7_0),.dout(w_dff_B_VkeaUpgj9_0),.clk(gclk));
	jdff dff_B_shnPEXPY1_0(.din(w_dff_B_VkeaUpgj9_0),.dout(w_dff_B_shnPEXPY1_0),.clk(gclk));
	jdff dff_B_px5ZdUIe7_0(.din(w_dff_B_shnPEXPY1_0),.dout(w_dff_B_px5ZdUIe7_0),.clk(gclk));
	jdff dff_B_0Nr7RXnD4_0(.din(w_dff_B_px5ZdUIe7_0),.dout(w_dff_B_0Nr7RXnD4_0),.clk(gclk));
	jdff dff_B_Rqgp33VM1_0(.din(w_dff_B_0Nr7RXnD4_0),.dout(w_dff_B_Rqgp33VM1_0),.clk(gclk));
	jdff dff_B_iv4zvYdQ6_1(.din(n413),.dout(w_dff_B_iv4zvYdQ6_1),.clk(gclk));
	jdff dff_A_K26thiWr8_0(.dout(w_G308_1[0]),.din(w_dff_A_K26thiWr8_0),.clk(gclk));
	jdff dff_B_pOQmJj3U1_1(.din(n400),.dout(w_dff_B_pOQmJj3U1_1),.clk(gclk));
	jdff dff_A_qS9klzNj2_1(.dout(w_n428_0[1]),.din(w_dff_A_qS9klzNj2_1),.clk(gclk));
	jdff dff_A_k3JB3iCB9_0(.dout(w_G361_1[0]),.din(w_dff_A_k3JB3iCB9_0),.clk(gclk));
	jdff dff_B_UnBdhMhv8_1(.din(n1485),.dout(w_dff_B_UnBdhMhv8_1),.clk(gclk));
	jdff dff_B_TTFTocGu1_2(.din(n437),.dout(w_dff_B_TTFTocGu1_2),.clk(gclk));
	jdff dff_A_GApiUB9Q9_0(.dout(w_G503_2[0]),.din(w_dff_A_GApiUB9Q9_0),.clk(gclk));
	jdff dff_A_WA0s8Mnc6_0(.dout(w_dff_A_GApiUB9Q9_0),.din(w_dff_A_WA0s8Mnc6_0),.clk(gclk));
	jdff dff_B_ojyNWK7c7_1(.din(n1481),.dout(w_dff_B_ojyNWK7c7_1),.clk(gclk));
	jdff dff_B_eZqKCXTv8_1(.din(n1471),.dout(w_dff_B_eZqKCXTv8_1),.clk(gclk));
	jdff dff_A_xQfn7MGY8_1(.dout(w_G341_2[1]),.din(w_dff_A_xQfn7MGY8_1),.clk(gclk));
	jdff dff_B_rGnss2399_1(.din(n1462),.dout(w_dff_B_rGnss2399_1),.clk(gclk));
	jdff dff_A_3YLb6Y9c1_1(.dout(w_G351_2[1]),.din(w_dff_A_3YLb6Y9c1_1),.clk(gclk));
	jdff dff_B_F8AqNKUb9_0(.din(n1460),.dout(w_dff_B_F8AqNKUb9_0),.clk(gclk));
	jdff dff_B_a3QL1NSg6_0(.din(w_dff_B_F8AqNKUb9_0),.dout(w_dff_B_a3QL1NSg6_0),.clk(gclk));
	jdff dff_B_VjOJsnXf6_0(.din(n1454),.dout(w_dff_B_VjOJsnXf6_0),.clk(gclk));
	jdff dff_B_rk4d4Bjk7_0(.din(w_dff_B_VjOJsnXf6_0),.dout(w_dff_B_rk4d4Bjk7_0),.clk(gclk));
	jdff dff_B_OzS5BOtS0_0(.din(w_dff_B_rk4d4Bjk7_0),.dout(w_dff_B_OzS5BOtS0_0),.clk(gclk));
	jdff dff_A_ltpBvl6H1_0(.dout(w_n749_5[0]),.din(w_dff_A_ltpBvl6H1_0),.clk(gclk));
	jdff dff_A_cB9ztAZT6_0(.dout(w_dff_A_ltpBvl6H1_0),.din(w_dff_A_cB9ztAZT6_0),.clk(gclk));
	jdff dff_A_2JdLEy3j5_0(.dout(w_dff_A_cB9ztAZT6_0),.din(w_dff_A_2JdLEy3j5_0),.clk(gclk));
	jdff dff_A_HpiOvwHi4_1(.dout(w_n749_5[1]),.din(w_dff_A_HpiOvwHi4_1),.clk(gclk));
	jdff dff_A_rgcPklOv7_1(.dout(w_dff_A_HpiOvwHi4_1),.din(w_dff_A_rgcPklOv7_1),.clk(gclk));
	jdff dff_A_9FMqmy381_1(.dout(w_dff_A_rgcPklOv7_1),.din(w_dff_A_9FMqmy381_1),.clk(gclk));
	jdff dff_A_OWQkBT059_1(.dout(w_dff_A_9FMqmy381_1),.din(w_dff_A_OWQkBT059_1),.clk(gclk));
	jdff dff_A_FhEXZ4ZW6_1(.dout(w_dff_A_OWQkBT059_1),.din(w_dff_A_FhEXZ4ZW6_1),.clk(gclk));
	jdff dff_A_38JcmSs84_1(.dout(w_dff_A_FhEXZ4ZW6_1),.din(w_dff_A_38JcmSs84_1),.clk(gclk));
	jdff dff_A_wCRS4pXC5_1(.dout(w_dff_A_38JcmSs84_1),.din(w_dff_A_wCRS4pXC5_1),.clk(gclk));
	jdff dff_A_tVNUeOV68_1(.dout(w_dff_A_wCRS4pXC5_1),.din(w_dff_A_tVNUeOV68_1),.clk(gclk));
	jdff dff_A_HhRntZwZ4_1(.dout(w_dff_A_tVNUeOV68_1),.din(w_dff_A_HhRntZwZ4_1),.clk(gclk));
	jdff dff_A_bZyt1uXS4_1(.dout(w_dff_A_HhRntZwZ4_1),.din(w_dff_A_bZyt1uXS4_1),.clk(gclk));
	jdff dff_A_WV7wOBFw4_1(.dout(w_dff_A_bZyt1uXS4_1),.din(w_dff_A_WV7wOBFw4_1),.clk(gclk));
	jdff dff_B_Snf1LqFt0_0(.din(n1452),.dout(w_dff_B_Snf1LqFt0_0),.clk(gclk));
	jdff dff_B_jMQYmiD85_0(.din(w_dff_B_Snf1LqFt0_0),.dout(w_dff_B_jMQYmiD85_0),.clk(gclk));
	jdff dff_B_cw8LeY8W6_0(.din(w_dff_B_jMQYmiD85_0),.dout(w_dff_B_cw8LeY8W6_0),.clk(gclk));
	jdff dff_B_Jh3TekGu0_0(.din(w_dff_B_cw8LeY8W6_0),.dout(w_dff_B_Jh3TekGu0_0),.clk(gclk));
	jdff dff_A_HyanecyJ0_0(.dout(w_n1451_0[0]),.din(w_dff_A_HyanecyJ0_0),.clk(gclk));
	jdff dff_A_53lSuFD73_0(.dout(w_dff_A_HyanecyJ0_0),.din(w_dff_A_53lSuFD73_0),.clk(gclk));
	jdff dff_A_8IqcREHf8_0(.dout(w_dff_A_53lSuFD73_0),.din(w_dff_A_8IqcREHf8_0),.clk(gclk));
	jdff dff_B_V58b9dXk3_0(.din(n1450),.dout(w_dff_B_V58b9dXk3_0),.clk(gclk));
	jdff dff_B_pVM2lMhF9_1(.din(n1448),.dout(w_dff_B_pVM2lMhF9_1),.clk(gclk));
	jdff dff_A_SF2gKTs29_0(.dout(w_n763_0[0]),.din(w_dff_A_SF2gKTs29_0),.clk(gclk));
	jdff dff_A_hCMtiU4E1_0(.dout(w_dff_A_SF2gKTs29_0),.din(w_dff_A_hCMtiU4E1_0),.clk(gclk));
	jdff dff_A_SehYSrqj3_0(.dout(w_dff_A_hCMtiU4E1_0),.din(w_dff_A_SehYSrqj3_0),.clk(gclk));
	jdff dff_A_foB81kUL3_0(.dout(w_dff_A_SehYSrqj3_0),.din(w_dff_A_foB81kUL3_0),.clk(gclk));
	jdff dff_A_jHvo7Xlk4_0(.dout(w_dff_A_foB81kUL3_0),.din(w_dff_A_jHvo7Xlk4_0),.clk(gclk));
	jdff dff_A_PwUBuEfH9_0(.dout(w_dff_A_jHvo7Xlk4_0),.din(w_dff_A_PwUBuEfH9_0),.clk(gclk));
	jdff dff_B_T3sxnq1M5_1(.din(n1439),.dout(w_dff_B_T3sxnq1M5_1),.clk(gclk));
	jdff dff_B_qYaK45dp7_1(.din(n1441),.dout(w_dff_B_qYaK45dp7_1),.clk(gclk));
	jdff dff_B_ZUAYicvz0_1(.din(w_dff_B_qYaK45dp7_1),.dout(w_dff_B_ZUAYicvz0_1),.clk(gclk));
	jdff dff_B_5mPxYXIv3_0(.din(n1442),.dout(w_dff_B_5mPxYXIv3_0),.clk(gclk));
	jdff dff_B_fdGNECGl8_0(.din(n1436),.dout(w_dff_B_fdGNECGl8_0),.clk(gclk));
	jdff dff_B_8e85yDFP6_0(.din(n1434),.dout(w_dff_B_8e85yDFP6_0),.clk(gclk));
	jdff dff_B_d3LsgjpI8_1(.din(n1430),.dout(w_dff_B_d3LsgjpI8_1),.clk(gclk));
	jdff dff_A_WwVYqvUf4_0(.dout(w_n1429_0[0]),.din(w_dff_A_WwVYqvUf4_0),.clk(gclk));
	jdff dff_A_5dDgk8ii0_0(.dout(w_n1428_0[0]),.din(w_dff_A_5dDgk8ii0_0),.clk(gclk));
	jdff dff_B_uNP6423W8_2(.din(n1428),.dout(w_dff_B_uNP6423W8_2),.clk(gclk));
	jdff dff_A_Q8QOtOSR2_0(.dout(w_n624_0[0]),.din(w_dff_A_Q8QOtOSR2_0),.clk(gclk));
	jdff dff_B_b6pFW9900_3(.din(n624),.dout(w_dff_B_b6pFW9900_3),.clk(gclk));
	jdff dff_B_1QNdUh026_3(.din(w_dff_B_b6pFW9900_3),.dout(w_dff_B_1QNdUh026_3),.clk(gclk));
	jdff dff_A_Fwgg2QO98_1(.dout(w_n620_1[1]),.din(w_dff_A_Fwgg2QO98_1),.clk(gclk));
	jdff dff_A_5nqX0Onf0_1(.dout(w_dff_A_Fwgg2QO98_1),.din(w_dff_A_5nqX0Onf0_1),.clk(gclk));
	jdff dff_A_9Oj3ozNS6_1(.dout(w_dff_A_5nqX0Onf0_1),.din(w_dff_A_9Oj3ozNS6_1),.clk(gclk));
	jdff dff_A_FaTiuKzn8_1(.dout(w_dff_A_9Oj3ozNS6_1),.din(w_dff_A_FaTiuKzn8_1),.clk(gclk));
	jdff dff_A_QrF8qCpc9_1(.dout(w_n620_0[1]),.din(w_dff_A_QrF8qCpc9_1),.clk(gclk));
	jdff dff_A_tLWPBBaU6_1(.dout(w_dff_A_QrF8qCpc9_1),.din(w_dff_A_tLWPBBaU6_1),.clk(gclk));
	jdff dff_A_QTSfA3wV0_1(.dout(w_dff_A_tLWPBBaU6_1),.din(w_dff_A_QTSfA3wV0_1),.clk(gclk));
	jdff dff_A_7xNlXekK5_2(.dout(w_n620_0[2]),.din(w_dff_A_7xNlXekK5_2),.clk(gclk));
	jdff dff_A_WXrc9FmN1_2(.dout(w_dff_A_7xNlXekK5_2),.din(w_dff_A_WXrc9FmN1_2),.clk(gclk));
	jdff dff_A_ypQB3onv6_2(.dout(w_dff_A_WXrc9FmN1_2),.din(w_dff_A_ypQB3onv6_2),.clk(gclk));
	jdff dff_A_Kfw9dmFK2_2(.dout(w_dff_A_ypQB3onv6_2),.din(w_dff_A_Kfw9dmFK2_2),.clk(gclk));
	jdff dff_A_pvFXFeQb3_2(.dout(w_dff_A_Kfw9dmFK2_2),.din(w_dff_A_pvFXFeQb3_2),.clk(gclk));
	jdff dff_A_ILyOpGBO9_2(.dout(w_dff_A_pvFXFeQb3_2),.din(w_dff_A_ILyOpGBO9_2),.clk(gclk));
	jdff dff_A_JjMk9zlO8_1(.dout(w_n618_0[1]),.din(w_dff_A_JjMk9zlO8_1),.clk(gclk));
	jdff dff_A_0H4spKl57_1(.dout(w_dff_A_JjMk9zlO8_1),.din(w_dff_A_0H4spKl57_1),.clk(gclk));
	jdff dff_A_dEErKEAa2_1(.dout(w_dff_A_0H4spKl57_1),.din(w_dff_A_dEErKEAa2_1),.clk(gclk));
	jdff dff_A_raMBdhc38_2(.dout(w_n618_0[2]),.din(w_dff_A_raMBdhc38_2),.clk(gclk));
	jdff dff_A_5GC5YbDb3_2(.dout(w_dff_A_raMBdhc38_2),.din(w_dff_A_5GC5YbDb3_2),.clk(gclk));
	jdff dff_B_xUii6bHv2_1(.din(n1411),.dout(w_dff_B_xUii6bHv2_1),.clk(gclk));
	jdff dff_B_9bgltcn55_1(.din(n1418),.dout(w_dff_B_9bgltcn55_1),.clk(gclk));
	jdff dff_B_VZZTiSp49_1(.din(w_dff_B_9bgltcn55_1),.dout(w_dff_B_VZZTiSp49_1),.clk(gclk));
	jdff dff_B_eNGpBWf86_1(.din(w_dff_B_VZZTiSp49_1),.dout(w_dff_B_eNGpBWf86_1),.clk(gclk));
	jdff dff_B_fRw42wEj5_1(.din(n1419),.dout(w_dff_B_fRw42wEj5_1),.clk(gclk));
	jdff dff_B_zsdy9Zl82_1(.din(w_dff_B_fRw42wEj5_1),.dout(w_dff_B_zsdy9Zl82_1),.clk(gclk));
	jdff dff_A_50hmwSDu7_2(.dout(w_n660_0[2]),.din(w_dff_A_50hmwSDu7_2),.clk(gclk));
	jdff dff_A_9kVgspdK1_2(.dout(w_dff_A_50hmwSDu7_2),.din(w_dff_A_9kVgspdK1_2),.clk(gclk));
	jdff dff_A_vhzWELfx7_2(.dout(w_dff_A_9kVgspdK1_2),.din(w_dff_A_vhzWELfx7_2),.clk(gclk));
	jdff dff_A_e4X0ADm52_2(.dout(w_n792_0[2]),.din(w_dff_A_e4X0ADm52_2),.clk(gclk));
	jdff dff_A_OXBJvEML1_2(.dout(w_dff_A_e4X0ADm52_2),.din(w_dff_A_OXBJvEML1_2),.clk(gclk));
	jdff dff_A_tg4nSsv12_2(.dout(w_dff_A_OXBJvEML1_2),.din(w_dff_A_tg4nSsv12_2),.clk(gclk));
	jdff dff_A_ZmXU0taD4_2(.dout(w_dff_A_tg4nSsv12_2),.din(w_dff_A_ZmXU0taD4_2),.clk(gclk));
	jdff dff_A_O57uuZ4N1_2(.dout(w_dff_A_ZmXU0taD4_2),.din(w_dff_A_O57uuZ4N1_2),.clk(gclk));
	jdff dff_A_yb7Rrzvm3_1(.dout(w_n790_0[1]),.din(w_dff_A_yb7Rrzvm3_1),.clk(gclk));
	jdff dff_A_l9btvlHH5_1(.dout(w_dff_A_yb7Rrzvm3_1),.din(w_dff_A_l9btvlHH5_1),.clk(gclk));
	jdff dff_A_YtBF5r7W8_1(.dout(w_dff_A_l9btvlHH5_1),.din(w_dff_A_YtBF5r7W8_1),.clk(gclk));
	jdff dff_A_tFxOJqQM1_1(.dout(w_dff_A_YtBF5r7W8_1),.din(w_dff_A_tFxOJqQM1_1),.clk(gclk));
	jdff dff_A_tLdKHldY0_1(.dout(w_dff_A_tFxOJqQM1_1),.din(w_dff_A_tLdKHldY0_1),.clk(gclk));
	jdff dff_A_hIUaBKai6_1(.dout(w_dff_A_tLdKHldY0_1),.din(w_dff_A_hIUaBKai6_1),.clk(gclk));
	jdff dff_A_xjVBSbwO5_1(.dout(w_dff_A_hIUaBKai6_1),.din(w_dff_A_xjVBSbwO5_1),.clk(gclk));
	jdff dff_A_GNJrBlpy1_2(.dout(w_n790_0[2]),.din(w_dff_A_GNJrBlpy1_2),.clk(gclk));
	jdff dff_A_NkL8CpXt2_1(.dout(w_n1416_0[1]),.din(w_dff_A_NkL8CpXt2_1),.clk(gclk));
	jdff dff_A_pYkteeSe7_1(.dout(w_dff_A_NkL8CpXt2_1),.din(w_dff_A_pYkteeSe7_1),.clk(gclk));
	jdff dff_B_WYHw19yU4_2(.din(n1416),.dout(w_dff_B_WYHw19yU4_2),.clk(gclk));
	jdff dff_B_bSGZwCqE4_2(.din(w_dff_B_WYHw19yU4_2),.dout(w_dff_B_bSGZwCqE4_2),.clk(gclk));
	jdff dff_B_X0R6Lci53_0(.din(n1415),.dout(w_dff_B_X0R6Lci53_0),.clk(gclk));
	jdff dff_A_75SbOFsv8_1(.dout(w_n821_0[1]),.din(w_dff_A_75SbOFsv8_1),.clk(gclk));
	jdff dff_A_ZdDOikhV5_1(.dout(w_dff_A_75SbOFsv8_1),.din(w_dff_A_ZdDOikhV5_1),.clk(gclk));
	jdff dff_B_c2vrybp85_1(.din(n812),.dout(w_dff_B_c2vrybp85_1),.clk(gclk));
	jdff dff_B_Tw5JmFPd0_1(.din(w_dff_B_c2vrybp85_1),.dout(w_dff_B_Tw5JmFPd0_1),.clk(gclk));
	jdff dff_B_e2WDhi7A7_1(.din(w_dff_B_Tw5JmFPd0_1),.dout(w_dff_B_e2WDhi7A7_1),.clk(gclk));
	jdff dff_B_UO8pbqDg9_1(.din(n813),.dout(w_dff_B_UO8pbqDg9_1),.clk(gclk));
	jdff dff_A_QpH1FV798_1(.dout(w_n819_0[1]),.din(w_dff_A_QpH1FV798_1),.clk(gclk));
	jdff dff_A_jTs244OI7_1(.dout(w_dff_A_QpH1FV798_1),.din(w_dff_A_jTs244OI7_1),.clk(gclk));
	jdff dff_A_xhbIWgCU4_1(.dout(w_dff_A_jTs244OI7_1),.din(w_dff_A_xhbIWgCU4_1),.clk(gclk));
	jdff dff_A_SXc5389j0_1(.dout(w_n632_0[1]),.din(w_dff_A_SXc5389j0_1),.clk(gclk));
	jdff dff_A_hPXqXdMT6_0(.dout(w_n814_0[0]),.din(w_dff_A_hPXqXdMT6_0),.clk(gclk));
	jdff dff_A_IPnPPsxj1_0(.dout(w_dff_A_hPXqXdMT6_0),.din(w_dff_A_IPnPPsxj1_0),.clk(gclk));
	jdff dff_A_PNJXGsJi1_1(.dout(w_n814_0[1]),.din(w_dff_A_PNJXGsJi1_1),.clk(gclk));
	jdff dff_A_4L6nhCvO8_1(.dout(w_dff_A_PNJXGsJi1_1),.din(w_dff_A_4L6nhCvO8_1),.clk(gclk));
	jdff dff_B_aWKtNM9w2_1(.din(n629),.dout(w_dff_B_aWKtNM9w2_1),.clk(gclk));
	jdff dff_B_V7Kax62f0_3(.din(n377),.dout(w_dff_B_V7Kax62f0_3),.clk(gclk));
	jdff dff_A_yyZ7EeFx5_0(.dout(w_G534_2[0]),.din(w_dff_A_yyZ7EeFx5_0),.clk(gclk));
	jdff dff_A_IFGDUsUK7_0(.dout(w_dff_A_yyZ7EeFx5_0),.din(w_dff_A_IFGDUsUK7_0),.clk(gclk));
	jdff dff_A_3hgCUxs04_1(.dout(w_n1412_0[1]),.din(w_dff_A_3hgCUxs04_1),.clk(gclk));
	jdff dff_A_AOtu1sjH4_1(.dout(w_dff_A_3hgCUxs04_1),.din(w_dff_A_AOtu1sjH4_1),.clk(gclk));
	jdff dff_A_HCs8vNtd3_1(.dout(w_dff_A_AOtu1sjH4_1),.din(w_dff_A_HCs8vNtd3_1),.clk(gclk));
	jdff dff_A_DiOjrdAz9_1(.dout(w_dff_A_HCs8vNtd3_1),.din(w_dff_A_DiOjrdAz9_1),.clk(gclk));
	jdff dff_A_jvyrUwuN8_1(.dout(w_dff_A_DiOjrdAz9_1),.din(w_dff_A_jvyrUwuN8_1),.clk(gclk));
	jdff dff_A_Xpu7Qeg40_2(.dout(w_n1412_0[2]),.din(w_dff_A_Xpu7Qeg40_2),.clk(gclk));
	jdff dff_A_XbTzPN4r2_2(.dout(w_dff_A_Xpu7Qeg40_2),.din(w_dff_A_XbTzPN4r2_2),.clk(gclk));
	jdff dff_A_EE610UcN3_2(.dout(w_dff_A_XbTzPN4r2_2),.din(w_dff_A_EE610UcN3_2),.clk(gclk));
	jdff dff_B_0moUcKQS9_3(.din(n1412),.dout(w_dff_B_0moUcKQS9_3),.clk(gclk));
	jdff dff_B_0gyQMMzy0_3(.din(w_dff_B_0moUcKQS9_3),.dout(w_dff_B_0gyQMMzy0_3),.clk(gclk));
	jdff dff_B_wgle9SfE6_3(.din(w_dff_B_0gyQMMzy0_3),.dout(w_dff_B_wgle9SfE6_3),.clk(gclk));
	jdff dff_B_gmsZvxHJ0_3(.din(w_dff_B_wgle9SfE6_3),.dout(w_dff_B_gmsZvxHJ0_3),.clk(gclk));
	jdff dff_B_YUyPreZ66_3(.din(w_dff_B_gmsZvxHJ0_3),.dout(w_dff_B_YUyPreZ66_3),.clk(gclk));
	jdff dff_B_kshmEO0R7_3(.din(w_dff_B_YUyPreZ66_3),.dout(w_dff_B_kshmEO0R7_3),.clk(gclk));
	jdff dff_B_33bhuAvl8_3(.din(w_dff_B_kshmEO0R7_3),.dout(w_dff_B_33bhuAvl8_3),.clk(gclk));
	jdff dff_A_q4NEHzuz9_0(.dout(w_G2174_0[0]),.din(w_dff_A_q4NEHzuz9_0),.clk(gclk));
	jdff dff_A_tT6hAK6U7_0(.dout(w_dff_A_q4NEHzuz9_0),.din(w_dff_A_tT6hAK6U7_0),.clk(gclk));
	jdff dff_A_BrgZqVO46_0(.dout(w_dff_A_tT6hAK6U7_0),.din(w_dff_A_BrgZqVO46_0),.clk(gclk));
	jdff dff_A_4UhCQXfS6_0(.dout(w_dff_A_BrgZqVO46_0),.din(w_dff_A_4UhCQXfS6_0),.clk(gclk));
	jdff dff_A_aujhon4S8_0(.dout(w_dff_A_4UhCQXfS6_0),.din(w_dff_A_aujhon4S8_0),.clk(gclk));
	jdff dff_A_OThn2ABh0_0(.dout(w_dff_A_aujhon4S8_0),.din(w_dff_A_OThn2ABh0_0),.clk(gclk));
	jdff dff_A_blw3zNgs9_0(.dout(w_dff_A_OThn2ABh0_0),.din(w_dff_A_blw3zNgs9_0),.clk(gclk));
	jdff dff_A_WWV3D3Pb2_0(.dout(w_dff_A_blw3zNgs9_0),.din(w_dff_A_WWV3D3Pb2_0),.clk(gclk));
	jdff dff_A_5oUjxY3r0_0(.dout(w_dff_A_WWV3D3Pb2_0),.din(w_dff_A_5oUjxY3r0_0),.clk(gclk));
	jdff dff_A_lsRdNO4i9_0(.dout(w_dff_A_5oUjxY3r0_0),.din(w_dff_A_lsRdNO4i9_0),.clk(gclk));
	jdff dff_A_HftPVBkU4_0(.dout(w_dff_A_lsRdNO4i9_0),.din(w_dff_A_HftPVBkU4_0),.clk(gclk));
	jdff dff_A_aXXG4IeB4_1(.dout(w_G2174_0[1]),.din(w_dff_A_aXXG4IeB4_1),.clk(gclk));
	jdff dff_A_CjNDb0Us0_1(.dout(w_dff_A_aXXG4IeB4_1),.din(w_dff_A_CjNDb0Us0_1),.clk(gclk));
	jdff dff_A_vgwD9PvH1_1(.dout(w_dff_A_CjNDb0Us0_1),.din(w_dff_A_vgwD9PvH1_1),.clk(gclk));
	jdff dff_A_HSb0cIJS1_1(.dout(w_dff_A_vgwD9PvH1_1),.din(w_dff_A_HSb0cIJS1_1),.clk(gclk));
	jdff dff_A_z1hpwgbH6_1(.dout(w_dff_A_HSb0cIJS1_1),.din(w_dff_A_z1hpwgbH6_1),.clk(gclk));
	jdff dff_A_AKymWHSA7_1(.dout(w_dff_A_z1hpwgbH6_1),.din(w_dff_A_AKymWHSA7_1),.clk(gclk));
	jdff dff_A_dEf9Dms78_1(.dout(w_dff_A_AKymWHSA7_1),.din(w_dff_A_dEf9Dms78_1),.clk(gclk));
	jdff dff_B_OpOkjfm44_0(.din(n1409),.dout(w_dff_B_OpOkjfm44_0),.clk(gclk));
	jdff dff_B_1pkzOlgn8_0(.din(w_dff_B_OpOkjfm44_0),.dout(w_dff_B_1pkzOlgn8_0),.clk(gclk));
	jdff dff_A_5VmbqH5C2_0(.dout(w_n401_0[0]),.din(w_dff_A_5VmbqH5C2_0),.clk(gclk));
	jdff dff_A_HHssrEh99_0(.dout(w_dff_A_5VmbqH5C2_0),.din(w_dff_A_HHssrEh99_0),.clk(gclk));
	jdff dff_A_BCuU1Rr21_0(.dout(w_dff_A_HHssrEh99_0),.din(w_dff_A_BCuU1Rr21_0),.clk(gclk));
	jdff dff_B_znryO9ie9_2(.din(n401),.dout(w_dff_B_znryO9ie9_2),.clk(gclk));
	jdff dff_A_67QwtZ6x4_0(.dout(w_G490_1[0]),.din(w_dff_A_67QwtZ6x4_0),.clk(gclk));
	jdff dff_A_VgQhHTKt5_0(.dout(w_dff_A_67QwtZ6x4_0),.din(w_dff_A_VgQhHTKt5_0),.clk(gclk));
	jdff dff_A_GewbPXuV0_1(.dout(w_n654_1[1]),.din(w_dff_A_GewbPXuV0_1),.clk(gclk));
	jdff dff_A_iBUMR8Ew2_1(.dout(w_dff_A_GewbPXuV0_1),.din(w_dff_A_iBUMR8Ew2_1),.clk(gclk));
	jdff dff_A_HNSQBfCa2_1(.dout(w_dff_A_iBUMR8Ew2_1),.din(w_dff_A_HNSQBfCa2_1),.clk(gclk));
	jdff dff_A_BTCzLtU25_1(.dout(w_dff_A_HNSQBfCa2_1),.din(w_dff_A_BTCzLtU25_1),.clk(gclk));
	jdff dff_A_Gv755MUa6_0(.dout(w_n644_0[0]),.din(w_dff_A_Gv755MUa6_0),.clk(gclk));
	jdff dff_A_sCyLSq6K7_0(.dout(w_dff_A_Gv755MUa6_0),.din(w_dff_A_sCyLSq6K7_0),.clk(gclk));
	jdff dff_A_nUcGYgwi3_0(.dout(w_dff_A_sCyLSq6K7_0),.din(w_dff_A_nUcGYgwi3_0),.clk(gclk));
	jdff dff_A_VtPrfV8H4_0(.dout(w_dff_A_nUcGYgwi3_0),.din(w_dff_A_VtPrfV8H4_0),.clk(gclk));
	jdff dff_A_QzxyHL7W6_0(.dout(w_dff_A_VtPrfV8H4_0),.din(w_dff_A_QzxyHL7W6_0),.clk(gclk));
	jdff dff_A_pfeWfZUr8_2(.dout(w_n644_0[2]),.din(w_dff_A_pfeWfZUr8_2),.clk(gclk));
	jdff dff_A_67GSnaxY0_2(.dout(w_dff_A_pfeWfZUr8_2),.din(w_dff_A_67GSnaxY0_2),.clk(gclk));
	jdff dff_A_SokhPaHg7_2(.dout(w_dff_A_67GSnaxY0_2),.din(w_dff_A_SokhPaHg7_2),.clk(gclk));
	jdff dff_A_8pzO0rXC3_1(.dout(w_G293_0[1]),.din(w_dff_A_8pzO0rXC3_1),.clk(gclk));
	jdff dff_A_bow1sMlW8_1(.dout(w_n746_0[1]),.din(w_dff_A_bow1sMlW8_1),.clk(gclk));
	jdff dff_B_TRF4NlcU8_1(.din(n741),.dout(w_dff_B_TRF4NlcU8_1),.clk(gclk));
	jdff dff_B_MF1kEDRA6_1(.din(w_dff_B_TRF4NlcU8_1),.dout(w_dff_B_MF1kEDRA6_1),.clk(gclk));
	jdff dff_B_67dmE65F9_1(.din(w_dff_B_MF1kEDRA6_1),.dout(w_dff_B_67dmE65F9_1),.clk(gclk));
	jdff dff_B_hbgrprrW0_1(.din(w_dff_B_67dmE65F9_1),.dout(w_dff_B_hbgrprrW0_1),.clk(gclk));
	jdff dff_A_BFctmDTz3_1(.dout(w_n742_0[1]),.din(w_dff_A_BFctmDTz3_1),.clk(gclk));
	jdff dff_A_zNwLQdnp5_1(.dout(w_dff_A_BFctmDTz3_1),.din(w_dff_A_zNwLQdnp5_1),.clk(gclk));
	jdff dff_A_4osPnoRv1_1(.dout(w_dff_A_zNwLQdnp5_1),.din(w_dff_A_4osPnoRv1_1),.clk(gclk));
	jdff dff_A_ttlHbz9T1_1(.dout(w_dff_A_4osPnoRv1_1),.din(w_dff_A_ttlHbz9T1_1),.clk(gclk));
	jdff dff_B_TBImO6FS6_0(.din(n657),.dout(w_dff_B_TBImO6FS6_0),.clk(gclk));
	jdff dff_B_OF3KwrDd9_0(.din(w_dff_B_TBImO6FS6_0),.dout(w_dff_B_OF3KwrDd9_0),.clk(gclk));
	jdff dff_B_aVgFD1dL9_1(.din(G323),.dout(w_dff_B_aVgFD1dL9_1),.clk(gclk));
	jdff dff_A_h3z2YUrv4_2(.dout(w_G316_0[2]),.din(w_dff_A_h3z2YUrv4_2),.clk(gclk));
	jdff dff_A_IUNEtqDF8_1(.dout(w_G490_0[1]),.din(w_dff_A_IUNEtqDF8_1),.clk(gclk));
	jdff dff_A_FUCJ8oFp2_1(.dout(w_dff_A_IUNEtqDF8_1),.din(w_dff_A_FUCJ8oFp2_1),.clk(gclk));
	jdff dff_A_1B2tUJY09_1(.dout(w_dff_A_FUCJ8oFp2_1),.din(w_dff_A_1B2tUJY09_1),.clk(gclk));
	jdff dff_A_1btaIGhu2_1(.dout(w_dff_A_1B2tUJY09_1),.din(w_dff_A_1btaIGhu2_1),.clk(gclk));
	jdff dff_A_TJSNIQ1X7_2(.dout(w_G490_0[2]),.din(w_dff_A_TJSNIQ1X7_2),.clk(gclk));
	jdff dff_A_z9A9yAvg2_2(.dout(w_dff_A_TJSNIQ1X7_2),.din(w_dff_A_z9A9yAvg2_2),.clk(gclk));
	jdff dff_A_x1trZjX05_2(.dout(w_dff_A_z9A9yAvg2_2),.din(w_dff_A_x1trZjX05_2),.clk(gclk));
	jdff dff_A_OezKpDzA1_2(.dout(w_dff_A_x1trZjX05_2),.din(w_dff_A_OezKpDzA1_2),.clk(gclk));
	jdff dff_A_r31cBjW88_0(.dout(w_n654_2[0]),.din(w_dff_A_r31cBjW88_0),.clk(gclk));
	jdff dff_A_JWWby9fX1_0(.dout(w_n654_0[0]),.din(w_dff_A_JWWby9fX1_0),.clk(gclk));
	jdff dff_B_VydjEBBC5_3(.din(n654),.dout(w_dff_B_VydjEBBC5_3),.clk(gclk));
	jdff dff_B_Xxy0llxD2_3(.din(w_dff_B_VydjEBBC5_3),.dout(w_dff_B_Xxy0llxD2_3),.clk(gclk));
	jdff dff_A_kNM03czV2_0(.dout(w_n653_0[0]),.din(w_dff_A_kNM03czV2_0),.clk(gclk));
	jdff dff_A_CC5zD9ys5_0(.dout(w_dff_A_kNM03czV2_0),.din(w_dff_A_CC5zD9ys5_0),.clk(gclk));
	jdff dff_B_iO5cs4jZ7_1(.din(n651),.dout(w_dff_B_iO5cs4jZ7_1),.clk(gclk));
	jdff dff_B_McNbNlnj5_1(.din(G315),.dout(w_dff_B_McNbNlnj5_1),.clk(gclk));
	jdff dff_A_rJlRsTwe4_0(.dout(w_n414_0[0]),.din(w_dff_A_rJlRsTwe4_0),.clk(gclk));
	jdff dff_B_7V7pwQqq8_2(.din(n414),.dout(w_dff_B_7V7pwQqq8_2),.clk(gclk));
	jdff dff_A_HP5uExgC5_0(.dout(w_G479_0[0]),.din(w_dff_A_HP5uExgC5_0),.clk(gclk));
	jdff dff_A_DybV0qOA6_0(.dout(w_dff_A_HP5uExgC5_0),.din(w_dff_A_DybV0qOA6_0),.clk(gclk));
	jdff dff_A_9u4yvsA51_1(.dout(w_G479_0[1]),.din(w_dff_A_9u4yvsA51_1),.clk(gclk));
	jdff dff_A_klxydncY7_1(.dout(w_dff_A_9u4yvsA51_1),.din(w_dff_A_klxydncY7_1),.clk(gclk));
	jdff dff_A_gI5B2grv5_1(.dout(w_n648_0[1]),.din(w_dff_A_gI5B2grv5_1),.clk(gclk));
	jdff dff_A_faQzdlrd2_1(.dout(w_dff_A_gI5B2grv5_1),.din(w_dff_A_faQzdlrd2_1),.clk(gclk));
	jdff dff_A_M7bze1R01_1(.dout(w_dff_A_faQzdlrd2_1),.din(w_dff_A_M7bze1R01_1),.clk(gclk));
	jdff dff_A_0voaKU4p9_1(.dout(w_dff_A_M7bze1R01_1),.din(w_dff_A_0voaKU4p9_1),.clk(gclk));
	jdff dff_A_oXvTveG19_2(.dout(w_n648_0[2]),.din(w_dff_A_oXvTveG19_2),.clk(gclk));
	jdff dff_A_dflQyUH87_2(.dout(w_dff_A_oXvTveG19_2),.din(w_dff_A_dflQyUH87_2),.clk(gclk));
	jdff dff_A_nGeZXjpX6_2(.dout(w_dff_A_dflQyUH87_2),.din(w_dff_A_nGeZXjpX6_2),.clk(gclk));
	jdff dff_A_0VnuRAWd0_2(.dout(w_dff_A_nGeZXjpX6_2),.din(w_dff_A_0VnuRAWd0_2),.clk(gclk));
	jdff dff_A_mQMoIth09_2(.dout(w_dff_A_0VnuRAWd0_2),.din(w_dff_A_mQMoIth09_2),.clk(gclk));
	jdff dff_B_QlA5UopO3_0(.din(n647),.dout(w_dff_B_QlA5UopO3_0),.clk(gclk));
	jdff dff_B_r1zOMHRi2_0(.din(w_dff_B_QlA5UopO3_0),.dout(w_dff_B_r1zOMHRi2_0),.clk(gclk));
	jdff dff_B_fshypG5j3_1(.din(G307),.dout(w_dff_B_fshypG5j3_1),.clk(gclk));
	jdff dff_A_Q6s4J0Ok9_0(.dout(w_G302_0[0]),.din(w_dff_A_Q6s4J0Ok9_0),.clk(gclk));
	jdff dff_A_NemSBIxA4_1(.dout(w_G302_0[1]),.din(w_dff_A_NemSBIxA4_1),.clk(gclk));
	jdff dff_A_UwMNUtlo7_1(.dout(w_n737_0[1]),.din(w_dff_A_UwMNUtlo7_1),.clk(gclk));
	jdff dff_A_h7wfmPoq5_2(.dout(w_n737_0[2]),.din(w_dff_A_h7wfmPoq5_2),.clk(gclk));
	jdff dff_A_cMvc9Qws4_2(.dout(w_dff_A_h7wfmPoq5_2),.din(w_dff_A_cMvc9Qws4_2),.clk(gclk));
	jdff dff_A_HIWORh2d2_2(.dout(w_dff_A_cMvc9Qws4_2),.din(w_dff_A_HIWORh2d2_2),.clk(gclk));
	jdff dff_A_k3vSyhWN3_2(.dout(w_dff_A_HIWORh2d2_2),.din(w_dff_A_k3vSyhWN3_2),.clk(gclk));
	jdff dff_A_sgODAPR95_0(.dout(w_n735_0[0]),.din(w_dff_A_sgODAPR95_0),.clk(gclk));
	jdff dff_B_tS6mCmRe0_0(.din(n732),.dout(w_dff_B_tS6mCmRe0_0),.clk(gclk));
	jdff dff_A_AuRtYqI56_0(.dout(w_n728_0[0]),.din(w_dff_A_AuRtYqI56_0),.clk(gclk));
	jdff dff_A_eAEeDcZA9_1(.dout(w_n635_0[1]),.din(w_dff_A_eAEeDcZA9_1),.clk(gclk));
	jdff dff_A_hNwrlskJ5_1(.dout(w_dff_A_eAEeDcZA9_1),.din(w_dff_A_hNwrlskJ5_1),.clk(gclk));
	jdff dff_B_of19NiuT7_1(.din(n633),.dout(w_dff_B_of19NiuT7_1),.clk(gclk));
	jdff dff_A_tUR2AhzW3_0(.dout(w_G366_0[0]),.din(w_dff_A_tUR2AhzW3_0),.clk(gclk));
	jdff dff_A_AJsusLjk2_0(.dout(w_G332_2[0]),.din(w_dff_A_AJsusLjk2_0),.clk(gclk));
	jdff dff_A_xm5kZ9st4_2(.dout(w_G332_2[2]),.din(w_dff_A_xm5kZ9st4_2),.clk(gclk));
	jdff dff_A_LnjJ634u3_0(.dout(w_n628_0[0]),.din(w_dff_A_LnjJ634u3_0),.clk(gclk));
	jdff dff_A_00MTdIt77_0(.dout(w_dff_A_LnjJ634u3_0),.din(w_dff_A_00MTdIt77_0),.clk(gclk));
	jdff dff_A_LwvZZmhx1_2(.dout(w_n628_0[2]),.din(w_dff_A_LwvZZmhx1_2),.clk(gclk));
	jdff dff_A_z1gmnbMd3_2(.dout(w_dff_A_LwvZZmhx1_2),.din(w_dff_A_z1gmnbMd3_2),.clk(gclk));
	jdff dff_A_CLGdv8Ko1_0(.dout(w_G358_0[0]),.din(w_dff_A_CLGdv8Ko1_0),.clk(gclk));
	jdff dff_A_tG7bxNfY2_1(.dout(w_n625_0[1]),.din(w_dff_A_tG7bxNfY2_1),.clk(gclk));
	jdff dff_A_PsHvd5hW2_2(.dout(w_G351_0[2]),.din(w_dff_A_PsHvd5hW2_2),.clk(gclk));
	jdff dff_A_tWNU14720_0(.dout(w_G534_0[0]),.din(w_dff_A_tWNU14720_0),.clk(gclk));
	jdff dff_A_mDu6K7KB9_0(.dout(w_dff_A_tWNU14720_0),.din(w_dff_A_mDu6K7KB9_0),.clk(gclk));
	jdff dff_A_0VsX9gSj1_2(.dout(w_G534_0[2]),.din(w_dff_A_0VsX9gSj1_2),.clk(gclk));
	jdff dff_A_22TePM3N9_2(.dout(w_dff_A_0VsX9gSj1_2),.din(w_dff_A_22TePM3N9_2),.clk(gclk));
	jdff dff_A_K3Qbqy7G6_0(.dout(w_n726_0[0]),.din(w_dff_A_K3Qbqy7G6_0),.clk(gclk));
	jdff dff_B_Y6uJcumH7_1(.din(n723),.dout(w_dff_B_Y6uJcumH7_1),.clk(gclk));
	jdff dff_A_d0mXA9PV1_0(.dout(w_G348_0[0]),.din(w_dff_A_d0mXA9PV1_0),.clk(gclk));
	jdff dff_A_oJvT7yWN6_1(.dout(w_G332_1[1]),.din(w_dff_A_oJvT7yWN6_1),.clk(gclk));
	jdff dff_A_FW533wll0_1(.dout(w_n621_0[1]),.din(w_dff_A_FW533wll0_1),.clk(gclk));
	jdff dff_A_ppkAAw5J0_2(.dout(w_G341_0[2]),.din(w_dff_A_ppkAAw5J0_2),.clk(gclk));
	jdff dff_B_heec8Ysv9_3(.din(n389),.dout(w_dff_B_heec8Ysv9_3),.clk(gclk));
	jdff dff_A_ynpSuS5k6_0(.dout(w_G523_1[0]),.din(w_dff_A_ynpSuS5k6_0),.clk(gclk));
	jdff dff_A_sHe4h7fx4_0(.dout(w_dff_A_ynpSuS5k6_0),.din(w_dff_A_sHe4h7fx4_0),.clk(gclk));
	jdff dff_A_pxelVl3Z0_1(.dout(w_G523_1[1]),.din(w_dff_A_pxelVl3Z0_1),.clk(gclk));
	jdff dff_A_RZ5VYcc30_1(.dout(w_dff_A_pxelVl3Z0_1),.din(w_dff_A_RZ5VYcc30_1),.clk(gclk));
	jdff dff_A_236AP8nm2_1(.dout(w_G523_0[1]),.din(w_dff_A_236AP8nm2_1),.clk(gclk));
	jdff dff_A_tWoPz4ME8_1(.dout(w_dff_A_236AP8nm2_1),.din(w_dff_A_tWoPz4ME8_1),.clk(gclk));
	jdff dff_A_zrSjxQI90_2(.dout(w_G523_0[2]),.din(w_dff_A_zrSjxQI90_2),.clk(gclk));
	jdff dff_A_mckreH0L8_2(.dout(w_dff_A_zrSjxQI90_2),.din(w_dff_A_mckreH0L8_2),.clk(gclk));
	jdff dff_A_gRoyY9iG4_1(.dout(w_n722_0[1]),.din(w_dff_A_gRoyY9iG4_1),.clk(gclk));
	jdff dff_A_n3Pl6qdE0_1(.dout(w_dff_A_gRoyY9iG4_1),.din(w_dff_A_n3Pl6qdE0_1),.clk(gclk));
	jdff dff_A_x5eB3vcn8_1(.dout(w_dff_A_n3Pl6qdE0_1),.din(w_dff_A_x5eB3vcn8_1),.clk(gclk));
	jdff dff_A_ELEi7V7m7_1(.dout(w_n721_0[1]),.din(w_dff_A_ELEi7V7m7_1),.clk(gclk));
	jdff dff_A_k5dAjeXQ4_1(.dout(w_dff_A_ELEi7V7m7_1),.din(w_dff_A_k5dAjeXQ4_1),.clk(gclk));
	jdff dff_A_11KyuPkZ3_1(.dout(w_dff_A_k5dAjeXQ4_1),.din(w_dff_A_11KyuPkZ3_1),.clk(gclk));
	jdff dff_A_N68OXoit7_1(.dout(w_dff_A_11KyuPkZ3_1),.din(w_dff_A_N68OXoit7_1),.clk(gclk));
	jdff dff_A_qYgJoz2A4_1(.dout(w_n619_0[1]),.din(w_dff_A_qYgJoz2A4_1),.clk(gclk));
	jdff dff_A_sUq2AmRE2_1(.dout(w_dff_A_qYgJoz2A4_1),.din(w_dff_A_sUq2AmRE2_1),.clk(gclk));
	jdff dff_A_kvH05xRp7_1(.dout(w_dff_A_sUq2AmRE2_1),.din(w_dff_A_kvH05xRp7_1),.clk(gclk));
	jdff dff_A_LtwD0vNX5_0(.dout(w_G338_0[0]),.din(w_dff_A_LtwD0vNX5_0),.clk(gclk));
	jdff dff_A_GEsH3DP62_0(.dout(w_G514_0[0]),.din(w_dff_A_GEsH3DP62_0),.clk(gclk));
	jdff dff_A_p7EyMcTN4_2(.dout(w_G514_0[2]),.din(w_dff_A_p7EyMcTN4_2),.clk(gclk));
	jdff dff_A_jvNcSafF1_1(.dout(w_n720_0[1]),.din(w_dff_A_jvNcSafF1_1),.clk(gclk));
	jdff dff_A_Udpa4Dlm8_1(.dout(w_dff_A_jvNcSafF1_1),.din(w_dff_A_Udpa4Dlm8_1),.clk(gclk));
	jdff dff_A_LSWA4SK34_1(.dout(w_n719_0[1]),.din(w_dff_A_LSWA4SK34_1),.clk(gclk));
	jdff dff_A_iYbMZzK97_1(.dout(w_dff_A_LSWA4SK34_1),.din(w_dff_A_iYbMZzK97_1),.clk(gclk));
	jdff dff_B_EV41gs3b0_0(.din(n616),.dout(w_dff_B_EV41gs3b0_0),.clk(gclk));
	jdff dff_B_dCZwKOI10_0(.din(w_dff_B_EV41gs3b0_0),.dout(w_dff_B_dCZwKOI10_0),.clk(gclk));
	jdff dff_A_Oz1kqe4N9_1(.dout(w_G331_0[1]),.din(w_dff_A_Oz1kqe4N9_1),.clk(gclk));
	jdff dff_A_jOXfclfh5_1(.dout(w_G324_1[1]),.din(w_dff_A_jOXfclfh5_1),.clk(gclk));
	jdff dff_A_PD6kO0Ym0_2(.dout(w_G324_0[2]),.din(w_dff_A_PD6kO0Ym0_2),.clk(gclk));
	jdff dff_A_x0IUNIDN8_0(.dout(w_G503_0[0]),.din(w_dff_A_x0IUNIDN8_0),.clk(gclk));
	jdff dff_A_K44uDDF16_0(.dout(w_dff_A_x0IUNIDN8_0),.din(w_dff_A_K44uDDF16_0),.clk(gclk));
	jdff dff_A_DvWIhjLR1_0(.dout(w_dff_A_K44uDDF16_0),.din(w_dff_A_DvWIhjLR1_0),.clk(gclk));
	jdff dff_A_JxeyMOSj2_0(.dout(w_dff_A_DvWIhjLR1_0),.din(w_dff_A_JxeyMOSj2_0),.clk(gclk));
	jdff dff_A_T7tHFmi49_2(.dout(w_G503_0[2]),.din(w_dff_A_T7tHFmi49_2),.clk(gclk));
	jdff dff_A_WcQnB2JF9_0(.dout(w_G4092_4[0]),.din(w_dff_A_WcQnB2JF9_0),.clk(gclk));
	jdff dff_A_nRuNkL557_0(.dout(w_dff_A_WcQnB2JF9_0),.din(w_dff_A_nRuNkL557_0),.clk(gclk));
	jdff dff_A_PFfUAP3b8_0(.dout(w_dff_A_nRuNkL557_0),.din(w_dff_A_PFfUAP3b8_0),.clk(gclk));
	jdff dff_A_CVj66qHQ4_0(.dout(w_dff_A_PFfUAP3b8_0),.din(w_dff_A_CVj66qHQ4_0),.clk(gclk));
	jdff dff_A_pula1oiE2_0(.dout(w_dff_A_CVj66qHQ4_0),.din(w_dff_A_pula1oiE2_0),.clk(gclk));
	jdff dff_A_osDBOpXY5_0(.dout(w_dff_A_pula1oiE2_0),.din(w_dff_A_osDBOpXY5_0),.clk(gclk));
	jdff dff_A_Q6r4r7rb3_0(.dout(w_dff_A_osDBOpXY5_0),.din(w_dff_A_Q6r4r7rb3_0),.clk(gclk));
	jdff dff_A_umhkggfb1_0(.dout(w_dff_A_Q6r4r7rb3_0),.din(w_dff_A_umhkggfb1_0),.clk(gclk));
	jdff dff_A_jTzFy5wh3_0(.dout(w_dff_A_umhkggfb1_0),.din(w_dff_A_jTzFy5wh3_0),.clk(gclk));
	jdff dff_A_yCuGPY7Q1_0(.dout(w_dff_A_jTzFy5wh3_0),.din(w_dff_A_yCuGPY7Q1_0),.clk(gclk));
	jdff dff_A_CzWOorUO5_0(.dout(w_dff_A_yCuGPY7Q1_0),.din(w_dff_A_CzWOorUO5_0),.clk(gclk));
	jdff dff_A_mmVvdwBw5_0(.dout(w_dff_A_CzWOorUO5_0),.din(w_dff_A_mmVvdwBw5_0),.clk(gclk));
	jdff dff_A_bOzkJjjs5_0(.dout(w_dff_A_mmVvdwBw5_0),.din(w_dff_A_bOzkJjjs5_0),.clk(gclk));
	jdff dff_A_hj3Pxhih1_0(.dout(w_G4092_1[0]),.din(w_dff_A_hj3Pxhih1_0),.clk(gclk));
	jdff dff_A_Ft5dKWl73_0(.dout(w_dff_A_hj3Pxhih1_0),.din(w_dff_A_Ft5dKWl73_0),.clk(gclk));
	jdff dff_A_u5ptFPJO7_0(.dout(w_dff_A_Ft5dKWl73_0),.din(w_dff_A_u5ptFPJO7_0),.clk(gclk));
	jdff dff_A_0c2haayH0_0(.dout(w_dff_A_u5ptFPJO7_0),.din(w_dff_A_0c2haayH0_0),.clk(gclk));
	jdff dff_A_PsXMDqsn9_2(.dout(w_G4092_1[2]),.din(w_dff_A_PsXMDqsn9_2),.clk(gclk));
	jdff dff_A_8Iwc0BAH6_2(.dout(w_dff_A_PsXMDqsn9_2),.din(w_dff_A_8Iwc0BAH6_2),.clk(gclk));
	jdff dff_A_2xvx20Dz2_2(.dout(w_dff_A_8Iwc0BAH6_2),.din(w_dff_A_2xvx20Dz2_2),.clk(gclk));
	jdff dff_B_B180yI9l9_0(.din(n1673),.dout(w_dff_B_B180yI9l9_0),.clk(gclk));
	jdff dff_B_wa4N5EPW1_0(.din(w_dff_B_B180yI9l9_0),.dout(w_dff_B_wa4N5EPW1_0),.clk(gclk));
	jdff dff_B_I6Vmu5Qf7_0(.din(w_dff_B_wa4N5EPW1_0),.dout(w_dff_B_I6Vmu5Qf7_0),.clk(gclk));
	jdff dff_B_EmxxxWDC5_0(.din(w_dff_B_I6Vmu5Qf7_0),.dout(w_dff_B_EmxxxWDC5_0),.clk(gclk));
	jdff dff_B_VH6yGqaa3_0(.din(w_dff_B_EmxxxWDC5_0),.dout(w_dff_B_VH6yGqaa3_0),.clk(gclk));
	jdff dff_B_AUeL5z2w3_0(.din(w_dff_B_VH6yGqaa3_0),.dout(w_dff_B_AUeL5z2w3_0),.clk(gclk));
	jdff dff_B_lZPwmdJr5_0(.din(w_dff_B_AUeL5z2w3_0),.dout(w_dff_B_lZPwmdJr5_0),.clk(gclk));
	jdff dff_B_m0LBZ8ps8_0(.din(w_dff_B_lZPwmdJr5_0),.dout(w_dff_B_m0LBZ8ps8_0),.clk(gclk));
	jdff dff_B_H7y67g0v5_0(.din(w_dff_B_m0LBZ8ps8_0),.dout(w_dff_B_H7y67g0v5_0),.clk(gclk));
	jdff dff_B_V825YOW41_0(.din(w_dff_B_H7y67g0v5_0),.dout(w_dff_B_V825YOW41_0),.clk(gclk));
	jdff dff_B_nwpjwDy64_0(.din(w_dff_B_V825YOW41_0),.dout(w_dff_B_nwpjwDy64_0),.clk(gclk));
	jdff dff_B_wanWD0270_0(.din(w_dff_B_nwpjwDy64_0),.dout(w_dff_B_wanWD0270_0),.clk(gclk));
	jdff dff_B_ytyy4KYs9_0(.din(w_dff_B_wanWD0270_0),.dout(w_dff_B_ytyy4KYs9_0),.clk(gclk));
	jdff dff_B_bkjl5Xja4_1(.din(n1588),.dout(w_dff_B_bkjl5Xja4_1),.clk(gclk));
	jdff dff_B_G2zMsgd27_1(.din(w_dff_B_bkjl5Xja4_1),.dout(w_dff_B_G2zMsgd27_1),.clk(gclk));
	jdff dff_B_XrdMZr1n8_1(.din(w_dff_B_G2zMsgd27_1),.dout(w_dff_B_XrdMZr1n8_1),.clk(gclk));
	jdff dff_B_tVYseWYk3_1(.din(w_dff_B_XrdMZr1n8_1),.dout(w_dff_B_tVYseWYk3_1),.clk(gclk));
	jdff dff_B_o5Sivf2n5_1(.din(w_dff_B_tVYseWYk3_1),.dout(w_dff_B_o5Sivf2n5_1),.clk(gclk));
	jdff dff_B_PYbTzFi39_1(.din(n1654),.dout(w_dff_B_PYbTzFi39_1),.clk(gclk));
	jdff dff_B_1WUmjhl90_0(.din(n1658),.dout(w_dff_B_1WUmjhl90_0),.clk(gclk));
	jdff dff_B_umz6snDn7_0(.din(n1657),.dout(w_dff_B_umz6snDn7_0),.clk(gclk));
	jdff dff_B_ptrbJwoT9_1(.din(n1655),.dout(w_dff_B_ptrbJwoT9_1),.clk(gclk));
	jdff dff_B_klZCwMge2_1(.din(n1647),.dout(w_dff_B_klZCwMge2_1),.clk(gclk));
	jdff dff_B_KVxKDGVU1_1(.din(w_dff_B_klZCwMge2_1),.dout(w_dff_B_KVxKDGVU1_1),.clk(gclk));
	jdff dff_B_L5oVnzO48_1(.din(n1645),.dout(w_dff_B_L5oVnzO48_1),.clk(gclk));
	jdff dff_B_pk3vYg6W7_0(.din(n1641),.dout(w_dff_B_pk3vYg6W7_0),.clk(gclk));
	jdff dff_A_duw3mAMP8_0(.dout(w_n609_0[0]),.din(w_dff_A_duw3mAMP8_0),.clk(gclk));
	jdff dff_A_RIzvgUbT6_1(.dout(w_n609_0[1]),.din(w_dff_A_RIzvgUbT6_1),.clk(gclk));
	jdff dff_A_fbotVb362_1(.dout(w_dff_A_RIzvgUbT6_1),.din(w_dff_A_fbotVb362_1),.clk(gclk));
	jdff dff_A_9V0wUiED8_1(.dout(w_dff_A_fbotVb362_1),.din(w_dff_A_9V0wUiED8_1),.clk(gclk));
	jdff dff_A_BFAkwIrk5_1(.dout(w_dff_A_9V0wUiED8_1),.din(w_dff_A_BFAkwIrk5_1),.clk(gclk));
	jdff dff_A_hHwEEgIP3_1(.dout(w_dff_A_BFAkwIrk5_1),.din(w_dff_A_hHwEEgIP3_1),.clk(gclk));
	jdff dff_A_hpqvISpo6_1(.dout(w_dff_A_hHwEEgIP3_1),.din(w_dff_A_hpqvISpo6_1),.clk(gclk));
	jdff dff_A_jBj7RvZ02_1(.dout(w_n962_0[1]),.din(w_dff_A_jBj7RvZ02_1),.clk(gclk));
	jdff dff_A_jwKbbin55_1(.dout(w_dff_A_jBj7RvZ02_1),.din(w_dff_A_jwKbbin55_1),.clk(gclk));
	jdff dff_A_USAtdbCA6_1(.dout(w_dff_A_jwKbbin55_1),.din(w_dff_A_USAtdbCA6_1),.clk(gclk));
	jdff dff_A_MOvyumZz3_1(.dout(w_dff_A_USAtdbCA6_1),.din(w_dff_A_MOvyumZz3_1),.clk(gclk));
	jdff dff_A_ZGWavH5e8_2(.dout(w_n938_0[2]),.din(w_dff_A_ZGWavH5e8_2),.clk(gclk));
	jdff dff_A_LrKwF3DL8_2(.dout(w_dff_A_ZGWavH5e8_2),.din(w_dff_A_LrKwF3DL8_2),.clk(gclk));
	jdff dff_A_vmsZkfZI1_2(.dout(w_dff_A_LrKwF3DL8_2),.din(w_dff_A_vmsZkfZI1_2),.clk(gclk));
	jdff dff_B_RCuyKb0I8_1(.din(n707),.dout(w_dff_B_RCuyKb0I8_1),.clk(gclk));
	jdff dff_B_LFGWI0nG2_1(.din(w_dff_B_RCuyKb0I8_1),.dout(w_dff_B_LFGWI0nG2_1),.clk(gclk));
	jdff dff_B_LKZCUakw4_1(.din(n708),.dout(w_dff_B_LKZCUakw4_1),.clk(gclk));
	jdff dff_B_GCIUjCEb3_1(.din(w_dff_B_LKZCUakw4_1),.dout(w_dff_B_GCIUjCEb3_1),.clk(gclk));
	jdff dff_A_z9nyDZ5I5_0(.dout(w_n713_0[0]),.din(w_dff_A_z9nyDZ5I5_0),.clk(gclk));
	jdff dff_A_tvJ5pTrB9_1(.dout(w_n713_0[1]),.din(w_dff_A_tvJ5pTrB9_1),.clk(gclk));
	jdff dff_A_02E25KrJ1_1(.dout(w_dff_A_tvJ5pTrB9_1),.din(w_dff_A_02E25KrJ1_1),.clk(gclk));
	jdff dff_A_YdvRnKQC1_1(.dout(w_dff_A_02E25KrJ1_1),.din(w_dff_A_YdvRnKQC1_1),.clk(gclk));
	jdff dff_A_MbcZdtJF0_1(.dout(w_dff_A_YdvRnKQC1_1),.din(w_dff_A_MbcZdtJF0_1),.clk(gclk));
	jdff dff_A_77v8mn7W1_1(.dout(w_dff_A_MbcZdtJF0_1),.din(w_dff_A_77v8mn7W1_1),.clk(gclk));
	jdff dff_A_B77uRN4V4_0(.dout(w_n710_0[0]),.din(w_dff_A_B77uRN4V4_0),.clk(gclk));
	jdff dff_A_1xSnFRRZ7_0(.dout(w_dff_A_B77uRN4V4_0),.din(w_dff_A_1xSnFRRZ7_0),.clk(gclk));
	jdff dff_A_UUoHSVdh5_0(.dout(w_dff_A_1xSnFRRZ7_0),.din(w_dff_A_UUoHSVdh5_0),.clk(gclk));
	jdff dff_A_gndSIIHq5_0(.dout(w_dff_A_UUoHSVdh5_0),.din(w_dff_A_gndSIIHq5_0),.clk(gclk));
	jdff dff_A_DaFQTWao4_0(.dout(w_dff_A_gndSIIHq5_0),.din(w_dff_A_DaFQTWao4_0),.clk(gclk));
	jdff dff_A_SVP84Jxj8_0(.dout(w_n597_0[0]),.din(w_dff_A_SVP84Jxj8_0),.clk(gclk));
	jdff dff_A_ybkX4O3d6_0(.dout(w_dff_A_SVP84Jxj8_0),.din(w_dff_A_ybkX4O3d6_0),.clk(gclk));
	jdff dff_A_c8BxFHsH8_0(.dout(w_dff_A_ybkX4O3d6_0),.din(w_dff_A_c8BxFHsH8_0),.clk(gclk));
	jdff dff_A_RfEBFwxt1_0(.dout(w_n496_1[0]),.din(w_dff_A_RfEBFwxt1_0),.clk(gclk));
	jdff dff_A_uFn72zPK9_0(.dout(w_dff_A_RfEBFwxt1_0),.din(w_dff_A_uFn72zPK9_0),.clk(gclk));
	jdff dff_A_a3aub9DV0_0(.dout(w_n1637_0[0]),.din(w_dff_A_a3aub9DV0_0),.clk(gclk));
	jdff dff_B_yPMzt06f5_2(.din(n1637),.dout(w_dff_B_yPMzt06f5_2),.clk(gclk));
	jdff dff_A_eQKtaybn8_1(.dout(w_n608_0[1]),.din(w_dff_A_eQKtaybn8_1),.clk(gclk));
	jdff dff_A_0l2Sv8Ge0_1(.dout(w_dff_A_eQKtaybn8_1),.din(w_dff_A_0l2Sv8Ge0_1),.clk(gclk));
	jdff dff_A_SsqQ17Nc6_1(.dout(w_dff_A_0l2Sv8Ge0_1),.din(w_dff_A_SsqQ17Nc6_1),.clk(gclk));
	jdff dff_A_QbxZYPDn2_1(.dout(w_dff_A_SsqQ17Nc6_1),.din(w_dff_A_QbxZYPDn2_1),.clk(gclk));
	jdff dff_A_hH69EzeS0_1(.dout(w_dff_A_QbxZYPDn2_1),.din(w_dff_A_hH69EzeS0_1),.clk(gclk));
	jdff dff_A_L4AHDBsg0_1(.dout(w_dff_A_hH69EzeS0_1),.din(w_dff_A_L4AHDBsg0_1),.clk(gclk));
	jdff dff_B_KTcfb66q6_0(.din(n606),.dout(w_dff_B_KTcfb66q6_0),.clk(gclk));
	jdff dff_B_sb7ax8Z62_0(.din(w_dff_B_KTcfb66q6_0),.dout(w_dff_B_sb7ax8Z62_0),.clk(gclk));
	jdff dff_B_6l8Es9rU3_1(.din(G217),.dout(w_dff_B_6l8Es9rU3_1),.clk(gclk));
	jdff dff_A_rPMYSFAn3_0(.dout(w_n592_0[0]),.din(w_dff_A_rPMYSFAn3_0),.clk(gclk));
	jdff dff_A_uX3tdavN5_0(.dout(w_dff_A_rPMYSFAn3_0),.din(w_dff_A_uX3tdavN5_0),.clk(gclk));
	jdff dff_A_6uAxBoPZ0_2(.dout(w_n592_0[2]),.din(w_dff_A_6uAxBoPZ0_2),.clk(gclk));
	jdff dff_A_vpZNlNcy9_2(.dout(w_dff_A_6uAxBoPZ0_2),.din(w_dff_A_vpZNlNcy9_2),.clk(gclk));
	jdff dff_A_cCq4LzdO9_2(.dout(w_dff_A_vpZNlNcy9_2),.din(w_dff_A_cCq4LzdO9_2),.clk(gclk));
	jdff dff_B_YBkNYZOG6_1(.din(n589),.dout(w_dff_B_YBkNYZOG6_1),.clk(gclk));
	jdff dff_B_VWEEJY1S1_1(.din(G209),.dout(w_dff_B_VWEEJY1S1_1),.clk(gclk));
	jdff dff_A_5gwSCMZM8_0(.dout(w_n602_0[0]),.din(w_dff_A_5gwSCMZM8_0),.clk(gclk));
	jdff dff_A_4wNAwRAf9_0(.dout(w_n711_0[0]),.din(w_dff_A_4wNAwRAf9_0),.clk(gclk));
	jdff dff_A_tVHTqF3h4_0(.dout(w_dff_A_4wNAwRAf9_0),.din(w_dff_A_tVHTqF3h4_0),.clk(gclk));
	jdff dff_B_rEpscLp15_2(.din(n711),.dout(w_dff_B_rEpscLp15_2),.clk(gclk));
	jdff dff_A_OdkKpBji1_2(.dout(w_n954_0[2]),.din(w_dff_A_OdkKpBji1_2),.clk(gclk));
	jdff dff_A_XqoSx2Ot9_2(.dout(w_dff_A_OdkKpBji1_2),.din(w_dff_A_XqoSx2Ot9_2),.clk(gclk));
	jdff dff_A_bluO7SOM9_2(.dout(w_dff_A_XqoSx2Ot9_2),.din(w_dff_A_bluO7SOM9_2),.clk(gclk));
	jdff dff_B_Ol8i2kYi7_2(.din(n1633),.dout(w_dff_B_Ol8i2kYi7_2),.clk(gclk));
	jdff dff_A_k86KeRhH0_1(.dout(w_n709_0[1]),.din(w_dff_A_k86KeRhH0_1),.clk(gclk));
	jdff dff_B_ez15tSP66_0(.din(n600),.dout(w_dff_B_ez15tSP66_0),.clk(gclk));
	jdff dff_B_Rvnwe1wD7_0(.din(w_dff_B_ez15tSP66_0),.dout(w_dff_B_Rvnwe1wD7_0),.clk(gclk));
	jdff dff_B_Bfz9YGEj0_1(.din(G225),.dout(w_dff_B_Bfz9YGEj0_1),.clk(gclk));
	jdff dff_B_qSDASetN6_0(.din(n595),.dout(w_dff_B_qSDASetN6_0),.clk(gclk));
	jdff dff_B_vi8uLsP27_0(.din(w_dff_B_qSDASetN6_0),.dout(w_dff_B_vi8uLsP27_0),.clk(gclk));
	jdff dff_B_JUCzJ7sa9_1(.din(G233),.dout(w_dff_B_JUCzJ7sa9_1),.clk(gclk));
	jdff dff_A_TrHiYAnk6_1(.dout(w_n703_0[1]),.din(w_dff_A_TrHiYAnk6_1),.clk(gclk));
	jdff dff_A_L2wK5FBO0_0(.dout(w_n701_0[0]),.din(w_dff_A_L2wK5FBO0_0),.clk(gclk));
	jdff dff_A_T52GB4Ep1_0(.dout(w_n685_0[0]),.din(w_dff_A_T52GB4Ep1_0),.clk(gclk));
	jdff dff_B_CoCtGuNQ8_2(.din(n685),.dout(w_dff_B_CoCtGuNQ8_2),.clk(gclk));
	jdff dff_A_PL9bxoyz9_0(.dout(w_n684_0[0]),.din(w_dff_A_PL9bxoyz9_0),.clk(gclk));
	jdff dff_A_E2bAMQPb5_1(.dout(w_n682_0[1]),.din(w_dff_A_E2bAMQPb5_1),.clk(gclk));
	jdff dff_A_plI47xaI9_1(.dout(w_dff_A_E2bAMQPb5_1),.din(w_dff_A_plI47xaI9_1),.clk(gclk));
	jdff dff_A_OdD1Xs1X1_1(.dout(w_dff_A_plI47xaI9_1),.din(w_dff_A_OdD1Xs1X1_1),.clk(gclk));
	jdff dff_A_hoaHWpBQ4_1(.dout(w_dff_A_OdD1Xs1X1_1),.din(w_dff_A_hoaHWpBQ4_1),.clk(gclk));
	jdff dff_A_Vg9ppsk36_2(.dout(w_n682_0[2]),.din(w_dff_A_Vg9ppsk36_2),.clk(gclk));
	jdff dff_A_HmoeU2K61_2(.dout(w_dff_A_Vg9ppsk36_2),.din(w_dff_A_HmoeU2K61_2),.clk(gclk));
	jdff dff_A_JHbzWgM82_2(.dout(w_dff_A_HmoeU2K61_2),.din(w_dff_A_JHbzWgM82_2),.clk(gclk));
	jdff dff_A_JSKQu7Ck0_2(.dout(w_dff_A_JHbzWgM82_2),.din(w_dff_A_JSKQu7Ck0_2),.clk(gclk));
	jdff dff_B_6sMTLta98_0(.din(n1630),.dout(w_dff_B_6sMTLta98_0),.clk(gclk));
	jdff dff_B_wzqnqoXo6_0(.din(w_dff_B_6sMTLta98_0),.dout(w_dff_B_wzqnqoXo6_0),.clk(gclk));
	jdff dff_B_2rOS53rP8_0(.din(w_dff_B_wzqnqoXo6_0),.dout(w_dff_B_2rOS53rP8_0),.clk(gclk));
	jdff dff_B_EZuZnK921_0(.din(w_dff_B_2rOS53rP8_0),.dout(w_dff_B_EZuZnK921_0),.clk(gclk));
	jdff dff_B_MIfKNEgW7_0(.din(w_dff_B_EZuZnK921_0),.dout(w_dff_B_MIfKNEgW7_0),.clk(gclk));
	jdff dff_B_Bci5bNEN8_0(.din(n1628),.dout(w_dff_B_Bci5bNEN8_0),.clk(gclk));
	jdff dff_B_0cOJAhcX5_0(.din(w_dff_B_Bci5bNEN8_0),.dout(w_dff_B_0cOJAhcX5_0),.clk(gclk));
	jdff dff_B_o79XuoKI2_1(.din(n1623),.dout(w_dff_B_o79XuoKI2_1),.clk(gclk));
	jdff dff_B_R6T6ydsP1_0(.din(n1622),.dout(w_dff_B_R6T6ydsP1_0),.clk(gclk));
	jdff dff_B_kyzhpD2z1_0(.din(w_dff_B_R6T6ydsP1_0),.dout(w_dff_B_kyzhpD2z1_0),.clk(gclk));
	jdff dff_B_as1BGSdU2_0(.din(w_dff_B_kyzhpD2z1_0),.dout(w_dff_B_as1BGSdU2_0),.clk(gclk));
	jdff dff_B_a5rfNWOn7_0(.din(n1620),.dout(w_dff_B_a5rfNWOn7_0),.clk(gclk));
	jdff dff_A_x9GwPzIU3_0(.dout(w_n1618_0[0]),.din(w_dff_A_x9GwPzIU3_0),.clk(gclk));
	jdff dff_A_JE3qdwRv2_0(.dout(w_dff_A_x9GwPzIU3_0),.din(w_dff_A_JE3qdwRv2_0),.clk(gclk));
	jdff dff_B_eaoXcS7P6_2(.din(n1618),.dout(w_dff_B_eaoXcS7P6_2),.clk(gclk));
	jdff dff_B_J3UtZMY82_2(.din(w_dff_B_eaoXcS7P6_2),.dout(w_dff_B_J3UtZMY82_2),.clk(gclk));
	jdff dff_B_p9whTygG0_2(.din(w_dff_B_J3UtZMY82_2),.dout(w_dff_B_p9whTygG0_2),.clk(gclk));
	jdff dff_B_UaKwaDPw5_2(.din(w_dff_B_p9whTygG0_2),.dout(w_dff_B_UaKwaDPw5_2),.clk(gclk));
	jdff dff_B_sMBNa4lp7_2(.din(w_dff_B_UaKwaDPw5_2),.dout(w_dff_B_sMBNa4lp7_2),.clk(gclk));
	jdff dff_B_u1wcZca27_2(.din(w_dff_B_sMBNa4lp7_2),.dout(w_dff_B_u1wcZca27_2),.clk(gclk));
	jdff dff_B_Nl6AlKv06_2(.din(w_dff_B_u1wcZca27_2),.dout(w_dff_B_Nl6AlKv06_2),.clk(gclk));
	jdff dff_B_4p4PURqQ7_2(.din(w_dff_B_Nl6AlKv06_2),.dout(w_dff_B_4p4PURqQ7_2),.clk(gclk));
	jdff dff_B_2Wbpd6sD9_2(.din(w_dff_B_4p4PURqQ7_2),.dout(w_dff_B_2Wbpd6sD9_2),.clk(gclk));
	jdff dff_A_7bwjDdvK2_0(.dout(w_G1497_0[0]),.din(w_dff_A_7bwjDdvK2_0),.clk(gclk));
	jdff dff_A_7qPjqhdK9_0(.dout(w_dff_A_7bwjDdvK2_0),.din(w_dff_A_7qPjqhdK9_0),.clk(gclk));
	jdff dff_A_jczKTll98_0(.dout(w_dff_A_7qPjqhdK9_0),.din(w_dff_A_jczKTll98_0),.clk(gclk));
	jdff dff_A_Aok4hIju0_0(.dout(w_dff_A_jczKTll98_0),.din(w_dff_A_Aok4hIju0_0),.clk(gclk));
	jdff dff_A_btxep7797_0(.dout(w_dff_A_Aok4hIju0_0),.din(w_dff_A_btxep7797_0),.clk(gclk));
	jdff dff_A_qZJYF48m2_0(.dout(w_dff_A_btxep7797_0),.din(w_dff_A_qZJYF48m2_0),.clk(gclk));
	jdff dff_A_O2MWxzCe1_0(.dout(w_dff_A_qZJYF48m2_0),.din(w_dff_A_O2MWxzCe1_0),.clk(gclk));
	jdff dff_A_Cp2LwsjL6_0(.dout(w_dff_A_O2MWxzCe1_0),.din(w_dff_A_Cp2LwsjL6_0),.clk(gclk));
	jdff dff_A_Sbe6xNlx1_0(.dout(w_dff_A_Cp2LwsjL6_0),.din(w_dff_A_Sbe6xNlx1_0),.clk(gclk));
	jdff dff_A_ZjZ2DZ7l8_0(.dout(w_dff_A_Sbe6xNlx1_0),.din(w_dff_A_ZjZ2DZ7l8_0),.clk(gclk));
	jdff dff_A_K1zS4y1F5_0(.dout(w_dff_A_ZjZ2DZ7l8_0),.din(w_dff_A_K1zS4y1F5_0),.clk(gclk));
	jdff dff_A_Zt4aQlix2_1(.dout(w_G1497_0[1]),.din(w_dff_A_Zt4aQlix2_1),.clk(gclk));
	jdff dff_A_I00WpwUb5_1(.dout(w_dff_A_Zt4aQlix2_1),.din(w_dff_A_I00WpwUb5_1),.clk(gclk));
	jdff dff_A_g1Svti6l9_1(.dout(w_dff_A_I00WpwUb5_1),.din(w_dff_A_g1Svti6l9_1),.clk(gclk));
	jdff dff_A_DrpQAFGN2_1(.dout(w_dff_A_g1Svti6l9_1),.din(w_dff_A_DrpQAFGN2_1),.clk(gclk));
	jdff dff_A_7Mj91jPD4_1(.dout(w_dff_A_DrpQAFGN2_1),.din(w_dff_A_7Mj91jPD4_1),.clk(gclk));
	jdff dff_A_lI3RzP6B5_1(.dout(w_dff_A_7Mj91jPD4_1),.din(w_dff_A_lI3RzP6B5_1),.clk(gclk));
	jdff dff_A_PODq0vZL2_1(.dout(w_dff_A_lI3RzP6B5_1),.din(w_dff_A_PODq0vZL2_1),.clk(gclk));
	jdff dff_A_V13W4NhE3_1(.dout(w_dff_A_PODq0vZL2_1),.din(w_dff_A_V13W4NhE3_1),.clk(gclk));
	jdff dff_A_ODvgMo6Y2_1(.dout(w_dff_A_V13W4NhE3_1),.din(w_dff_A_ODvgMo6Y2_1),.clk(gclk));
	jdff dff_B_sOIUIeEh4_1(.din(n1600),.dout(w_dff_B_sOIUIeEh4_1),.clk(gclk));
	jdff dff_B_rXtbchKY7_0(.din(n1614),.dout(w_dff_B_rXtbchKY7_0),.clk(gclk));
	jdff dff_A_xh1MlD5z4_0(.dout(w_n865_0[0]),.din(w_dff_A_xh1MlD5z4_0),.clk(gclk));
	jdff dff_A_x94Gyz5M4_2(.dout(w_n865_0[2]),.din(w_dff_A_x94Gyz5M4_2),.clk(gclk));
	jdff dff_A_rhu1SLX75_2(.dout(w_dff_A_x94Gyz5M4_2),.din(w_dff_A_rhu1SLX75_2),.clk(gclk));
	jdff dff_A_VMAvBlKx6_2(.dout(w_dff_A_rhu1SLX75_2),.din(w_dff_A_VMAvBlKx6_2),.clk(gclk));
	jdff dff_A_otpvEPg61_1(.dout(w_n587_0[1]),.din(w_dff_A_otpvEPg61_1),.clk(gclk));
	jdff dff_A_VmCc0SdF6_1(.dout(w_dff_A_otpvEPg61_1),.din(w_dff_A_VmCc0SdF6_1),.clk(gclk));
	jdff dff_A_gspL3bJU9_1(.dout(w_dff_A_VmCc0SdF6_1),.din(w_dff_A_gspL3bJU9_1),.clk(gclk));
	jdff dff_B_JGqTnb7k3_0(.din(n585),.dout(w_dff_B_JGqTnb7k3_0),.clk(gclk));
	jdff dff_B_xbfNDrb60_0(.din(w_dff_B_JGqTnb7k3_0),.dout(w_dff_B_xbfNDrb60_0),.clk(gclk));
	jdff dff_B_s1Lg2lHD0_1(.din(G241),.dout(w_dff_B_s1Lg2lHD0_1),.clk(gclk));
	jdff dff_B_U8dG6jcS2_0(.din(n1610),.dout(w_dff_B_U8dG6jcS2_0),.clk(gclk));
	jdff dff_A_usuy5aFg9_0(.dout(w_n1609_0[0]),.din(w_dff_A_usuy5aFg9_0),.clk(gclk));
	jdff dff_B_HQmzkpsW9_2(.din(n1609),.dout(w_dff_B_HQmzkpsW9_2),.clk(gclk));
	jdff dff_A_AyQKETKV8_1(.dout(w_n1603_0[1]),.din(w_dff_A_AyQKETKV8_1),.clk(gclk));
	jdff dff_A_End4mDRM1_1(.dout(w_n687_0[1]),.din(w_dff_A_End4mDRM1_1),.clk(gclk));
	jdff dff_A_a0Lwgxvx6_1(.dout(w_dff_A_End4mDRM1_1),.din(w_dff_A_a0Lwgxvx6_1),.clk(gclk));
	jdff dff_A_khTp7iO64_1(.dout(w_dff_A_a0Lwgxvx6_1),.din(w_dff_A_khTp7iO64_1),.clk(gclk));
	jdff dff_A_mdmMYsyg7_1(.dout(w_n686_0[1]),.din(w_dff_A_mdmMYsyg7_1),.clk(gclk));
	jdff dff_A_633fGYG73_1(.dout(w_dff_A_mdmMYsyg7_1),.din(w_dff_A_633fGYG73_1),.clk(gclk));
	jdff dff_A_DfkzCR1E7_1(.dout(w_dff_A_633fGYG73_1),.din(w_dff_A_DfkzCR1E7_1),.clk(gclk));
	jdff dff_B_weWeD51m0_0(.din(n580),.dout(w_dff_B_weWeD51m0_0),.clk(gclk));
	jdff dff_A_n64hHnDN6_1(.dout(w_n579_1[1]),.din(w_dff_A_n64hHnDN6_1),.clk(gclk));
	jdff dff_A_KwzCzioj9_1(.dout(w_n579_0[1]),.din(w_dff_A_KwzCzioj9_1),.clk(gclk));
	jdff dff_A_JZ5umaZO8_2(.dout(w_n579_0[2]),.din(w_dff_A_JZ5umaZO8_2),.clk(gclk));
	jdff dff_A_gGE1DTIe7_2(.dout(w_dff_A_JZ5umaZO8_2),.din(w_dff_A_gGE1DTIe7_2),.clk(gclk));
	jdff dff_A_8m8VzK7g3_2(.dout(w_dff_A_gGE1DTIe7_2),.din(w_dff_A_8m8VzK7g3_2),.clk(gclk));
	jdff dff_B_75ERfvS76_0(.din(n577),.dout(w_dff_B_75ERfvS76_0),.clk(gclk));
	jdff dff_B_RJyCFA7L9_0(.din(w_dff_B_75ERfvS76_0),.dout(w_dff_B_RJyCFA7L9_0),.clk(gclk));
	jdff dff_B_Z0FhR6SO8_1(.din(G264),.dout(w_dff_B_Z0FhR6SO8_1),.clk(gclk));
	jdff dff_A_AbPZAwis7_1(.dout(w_n574_0[1]),.din(w_dff_A_AbPZAwis7_1),.clk(gclk));
	jdff dff_A_TtdV9xNS0_0(.dout(w_n1599_0[0]),.din(w_dff_A_TtdV9xNS0_0),.clk(gclk));
	jdff dff_B_SVP5Y5N34_0(.din(n1598),.dout(w_dff_B_SVP5Y5N34_0),.clk(gclk));
	jdff dff_B_CkHicxHn5_0(.din(n1597),.dout(w_dff_B_CkHicxHn5_0),.clk(gclk));
	jdff dff_B_P5UkVFyp5_0(.din(w_dff_B_CkHicxHn5_0),.dout(w_dff_B_P5UkVFyp5_0),.clk(gclk));
	jdff dff_A_DZ4rb1pn2_2(.dout(w_n923_0[2]),.din(w_dff_A_DZ4rb1pn2_2),.clk(gclk));
	jdff dff_A_RqEWupQx7_2(.dout(w_dff_A_DZ4rb1pn2_2),.din(w_dff_A_RqEWupQx7_2),.clk(gclk));
	jdff dff_B_uCsSlT233_1(.din(n1594),.dout(w_dff_B_uCsSlT233_1),.clk(gclk));
	jdff dff_A_KiCxKFaz6_0(.dout(w_n573_0[0]),.din(w_dff_A_KiCxKFaz6_0),.clk(gclk));
	jdff dff_A_AoskPmD63_1(.dout(w_n573_0[1]),.din(w_dff_A_AoskPmD63_1),.clk(gclk));
	jdff dff_A_6zW5vQiK3_1(.dout(w_dff_A_AoskPmD63_1),.din(w_dff_A_6zW5vQiK3_1),.clk(gclk));
	jdff dff_A_m3dvtZfp2_1(.dout(w_n699_0[1]),.din(w_dff_A_m3dvtZfp2_1),.clk(gclk));
	jdff dff_B_5UMaX4ZM0_1(.din(n691),.dout(w_dff_B_5UMaX4ZM0_1),.clk(gclk));
	jdff dff_B_Rd6uJHVp0_1(.din(w_dff_B_5UMaX4ZM0_1),.dout(w_dff_B_Rd6uJHVp0_1),.clk(gclk));
	jdff dff_B_dEl6L4no0_0(.din(n697),.dout(w_dff_B_dEl6L4no0_0),.clk(gclk));
	jdff dff_A_92TCUL8i1_1(.dout(w_n695_0[1]),.din(w_dff_A_92TCUL8i1_1),.clk(gclk));
	jdff dff_B_WqTalyok5_0(.din(n693),.dout(w_dff_B_WqTalyok5_0),.clk(gclk));
	jdff dff_A_1iQtT2Lb3_1(.dout(w_n564_0[1]),.din(w_dff_A_1iQtT2Lb3_1),.clk(gclk));
	jdff dff_A_wZAo4vm67_1(.dout(w_dff_A_1iQtT2Lb3_1),.din(w_dff_A_wZAo4vm67_1),.clk(gclk));
	jdff dff_B_H8GXBcUn2_1(.din(G280),.dout(w_dff_B_H8GXBcUn2_1),.clk(gclk));
	jdff dff_A_lQRMyj9D2_0(.dout(w_n692_0[0]),.din(w_dff_A_lQRMyj9D2_0),.clk(gclk));
	jdff dff_A_gGnrurns2_1(.dout(w_n559_0[1]),.din(w_dff_A_gGnrurns2_1),.clk(gclk));
	jdff dff_A_SRqVufOq5_1(.dout(w_dff_A_gGnrurns2_1),.din(w_dff_A_SRqVufOq5_1),.clk(gclk));
	jdff dff_B_N5KTHUmM9_1(.din(G288),.dout(w_dff_B_N5KTHUmM9_1),.clk(gclk));
	jdff dff_A_F8hozB7X3_0(.dout(w_n690_0[0]),.din(w_dff_A_F8hozB7X3_0),.clk(gclk));
	jdff dff_A_QCsdzEps4_1(.dout(w_n571_0[1]),.din(w_dff_A_QCsdzEps4_1),.clk(gclk));
	jdff dff_A_VCHzWWBO2_1(.dout(w_dff_A_QCsdzEps4_1),.din(w_dff_A_VCHzWWBO2_1),.clk(gclk));
	jdff dff_B_xvI34cRN7_1(.din(G272),.dout(w_dff_B_xvI34cRN7_1),.clk(gclk));
	jdff dff_B_OaFX81gL2_0(.din(n1585),.dout(w_dff_B_OaFX81gL2_0),.clk(gclk));
	jdff dff_B_8xCPJpTY7_1(.din(n1575),.dout(w_dff_B_8xCPJpTY7_1),.clk(gclk));
	jdff dff_A_XZylqcdf9_0(.dout(w_G210_2[0]),.din(w_dff_A_XZylqcdf9_0),.clk(gclk));
	jdff dff_A_zngNaiEX2_1(.dout(w_n451_0[1]),.din(w_dff_A_zngNaiEX2_1),.clk(gclk));
	jdff dff_A_SrzM1ZCC3_1(.dout(w_dff_A_zngNaiEX2_1),.din(w_dff_A_SrzM1ZCC3_1),.clk(gclk));
	jdff dff_B_glHv4Be06_3(.din(n451),.dout(w_dff_B_glHv4Be06_3),.clk(gclk));
	jdff dff_A_0e8Tz4Da4_0(.dout(w_G457_1[0]),.din(w_dff_A_0e8Tz4Da4_0),.clk(gclk));
	jdff dff_A_Nen14reh1_0(.dout(w_dff_A_0e8Tz4Da4_0),.din(w_dff_A_Nen14reh1_0),.clk(gclk));
	jdff dff_A_SLOptLUN8_0(.dout(w_dff_A_Nen14reh1_0),.din(w_dff_A_SLOptLUN8_0),.clk(gclk));
	jdff dff_A_29KEvHpM3_0(.dout(w_dff_A_SLOptLUN8_0),.din(w_dff_A_29KEvHpM3_0),.clk(gclk));
	jdff dff_A_1AcOq1Na9_1(.dout(w_G457_1[1]),.din(w_dff_A_1AcOq1Na9_1),.clk(gclk));
	jdff dff_A_dVbwrVjr4_1(.dout(w_dff_A_1AcOq1Na9_1),.din(w_dff_A_dVbwrVjr4_1),.clk(gclk));
	jdff dff_A_m5XaaJW91_1(.dout(w_G457_0[1]),.din(w_dff_A_m5XaaJW91_1),.clk(gclk));
	jdff dff_A_UpmAJVRc9_1(.dout(w_dff_A_m5XaaJW91_1),.din(w_dff_A_UpmAJVRc9_1),.clk(gclk));
	jdff dff_A_s37Gi0y91_2(.dout(w_G457_0[2]),.din(w_dff_A_s37Gi0y91_2),.clk(gclk));
	jdff dff_A_stElDjSk7_2(.dout(w_dff_A_s37Gi0y91_2),.din(w_dff_A_stElDjSk7_2),.clk(gclk));
	jdff dff_A_btWbsP4p8_2(.dout(w_dff_A_stElDjSk7_2),.din(w_dff_A_btWbsP4p8_2),.clk(gclk));
	jdff dff_A_wCHQqrQ66_2(.dout(w_dff_A_btWbsP4p8_2),.din(w_dff_A_wCHQqrQ66_2),.clk(gclk));
	jdff dff_A_eCxoAzf34_2(.dout(w_G210_0[2]),.din(w_dff_A_eCxoAzf34_2),.clk(gclk));
	jdff dff_B_RYzTC9Qw3_1(.din(n1570),.dout(w_dff_B_RYzTC9Qw3_1),.clk(gclk));
	jdff dff_A_k924Gbdg9_1(.dout(w_n509_0[1]),.din(w_dff_A_k924Gbdg9_1),.clk(gclk));
	jdff dff_A_ynWu1gvJ3_1(.dout(w_dff_A_k924Gbdg9_1),.din(w_dff_A_ynWu1gvJ3_1),.clk(gclk));
	jdff dff_B_Jd8Y8iK58_3(.din(n509),.dout(w_dff_B_Jd8Y8iK58_3),.clk(gclk));
	jdff dff_A_ENpVegIb2_0(.dout(w_G468_1[0]),.din(w_dff_A_ENpVegIb2_0),.clk(gclk));
	jdff dff_A_BPiz1hj92_0(.dout(w_dff_A_ENpVegIb2_0),.din(w_dff_A_BPiz1hj92_0),.clk(gclk));
	jdff dff_A_6oM2yfUC7_0(.dout(w_dff_A_BPiz1hj92_0),.din(w_dff_A_6oM2yfUC7_0),.clk(gclk));
	jdff dff_A_ewlGzfSJ4_0(.dout(w_dff_A_6oM2yfUC7_0),.din(w_dff_A_ewlGzfSJ4_0),.clk(gclk));
	jdff dff_A_hiaybn1G9_1(.dout(w_G468_1[1]),.din(w_dff_A_hiaybn1G9_1),.clk(gclk));
	jdff dff_A_SE6sVdrN9_1(.dout(w_dff_A_hiaybn1G9_1),.din(w_dff_A_SE6sVdrN9_1),.clk(gclk));
	jdff dff_B_9sfsuSSR1_1(.din(n1566),.dout(w_dff_B_9sfsuSSR1_1),.clk(gclk));
	jdff dff_A_8zdwvfop7_0(.dout(w_G218_1[0]),.din(w_dff_A_8zdwvfop7_0),.clk(gclk));
	jdff dff_A_HOf4kQdV8_1(.dout(w_G468_0[1]),.din(w_dff_A_HOf4kQdV8_1),.clk(gclk));
	jdff dff_A_cQUCsWo01_2(.dout(w_G468_0[2]),.din(w_dff_A_cQUCsWo01_2),.clk(gclk));
	jdff dff_A_LM8TSfZa7_2(.dout(w_dff_A_cQUCsWo01_2),.din(w_dff_A_LM8TSfZa7_2),.clk(gclk));
	jdff dff_A_Zhpq7rLM0_2(.dout(w_dff_A_LM8TSfZa7_2),.din(w_dff_A_Zhpq7rLM0_2),.clk(gclk));
	jdff dff_A_penQLU6r8_2(.dout(w_dff_A_Zhpq7rLM0_2),.din(w_dff_A_penQLU6r8_2),.clk(gclk));
	jdff dff_A_ayZZV8Mh8_0(.dout(w_G218_2[0]),.din(w_dff_A_ayZZV8Mh8_0),.clk(gclk));
	jdff dff_B_DrhtTbPM2_1(.din(n1556),.dout(w_dff_B_DrhtTbPM2_1),.clk(gclk));
	jdff dff_A_hSJTcLhb5_0(.dout(w_G226_2[0]),.din(w_dff_A_hSJTcLhb5_0),.clk(gclk));
	jdff dff_A_A5K82NNl8_2(.dout(w_n496_0[2]),.din(w_dff_A_A5K82NNl8_2),.clk(gclk));
	jdff dff_A_IGkRkcEo3_2(.dout(w_dff_A_A5K82NNl8_2),.din(w_dff_A_IGkRkcEo3_2),.clk(gclk));
	jdff dff_A_21qrzfBF6_2(.dout(w_dff_A_IGkRkcEo3_2),.din(w_dff_A_21qrzfBF6_2),.clk(gclk));
	jdff dff_B_2Ugq5SDK0_3(.din(n496),.dout(w_dff_B_2Ugq5SDK0_3),.clk(gclk));
	jdff dff_A_4en0RrWo9_0(.dout(w_G422_1[0]),.din(w_dff_A_4en0RrWo9_0),.clk(gclk));
	jdff dff_A_UaZNyiSJ8_0(.dout(w_dff_A_4en0RrWo9_0),.din(w_dff_A_UaZNyiSJ8_0),.clk(gclk));
	jdff dff_A_9eAdTEaV6_1(.dout(w_G422_0[1]),.din(w_dff_A_9eAdTEaV6_1),.clk(gclk));
	jdff dff_A_6QueWslw8_1(.dout(w_dff_A_9eAdTEaV6_1),.din(w_dff_A_6QueWslw8_1),.clk(gclk));
	jdff dff_A_lnyqTAaI3_2(.dout(w_G422_0[2]),.din(w_dff_A_lnyqTAaI3_2),.clk(gclk));
	jdff dff_A_0u4JD2Gl6_2(.dout(w_dff_A_lnyqTAaI3_2),.din(w_dff_A_0u4JD2Gl6_2),.clk(gclk));
	jdff dff_A_2yAw5N0q6_2(.dout(w_dff_A_0u4JD2Gl6_2),.din(w_dff_A_2yAw5N0q6_2),.clk(gclk));
	jdff dff_A_OW3w21rU4_2(.dout(w_dff_A_2yAw5N0q6_2),.din(w_dff_A_OW3w21rU4_2),.clk(gclk));
	jdff dff_A_Hk7IFeeq8_2(.dout(w_G226_0[2]),.din(w_dff_A_Hk7IFeeq8_2),.clk(gclk));
	jdff dff_B_OQMF5acT7_1(.din(n541),.dout(w_dff_B_OQMF5acT7_1),.clk(gclk));
	jdff dff_B_2EtDnD859_1(.din(n542),.dout(w_dff_B_2EtDnD859_1),.clk(gclk));
	jdff dff_A_cjOigGYo4_0(.dout(w_G446_1[0]),.din(w_dff_A_cjOigGYo4_0),.clk(gclk));
	jdff dff_A_PUPbGg4F4_0(.dout(w_dff_A_cjOigGYo4_0),.din(w_dff_A_PUPbGg4F4_0),.clk(gclk));
	jdff dff_A_pWTYFmGH7_1(.dout(w_G446_1[1]),.din(w_dff_A_pWTYFmGH7_1),.clk(gclk));
	jdff dff_A_tBxglOLO9_1(.dout(w_dff_A_pWTYFmGH7_1),.din(w_dff_A_tBxglOLO9_1),.clk(gclk));
	jdff dff_A_MZY9Vevh7_1(.dout(w_G446_0[1]),.din(w_dff_A_MZY9Vevh7_1),.clk(gclk));
	jdff dff_A_0GvYtfUI6_1(.dout(w_dff_A_MZY9Vevh7_1),.din(w_dff_A_0GvYtfUI6_1),.clk(gclk));
	jdff dff_A_t3r0Xzeu5_2(.dout(w_G446_0[2]),.din(w_dff_A_t3r0Xzeu5_2),.clk(gclk));
	jdff dff_A_8HkfzeEk4_2(.dout(w_dff_A_t3r0Xzeu5_2),.din(w_dff_A_8HkfzeEk4_2),.clk(gclk));
	jdff dff_A_NIY42FNy3_0(.dout(w_G206_1[0]),.din(w_dff_A_NIY42FNy3_0),.clk(gclk));
	jdff dff_B_Cp9r5I7Y0_1(.din(n1525),.dout(w_dff_B_Cp9r5I7Y0_1),.clk(gclk));
	jdff dff_B_DtwF8QNr1_1(.din(n1534),.dout(w_dff_B_DtwF8QNr1_1),.clk(gclk));
	jdff dff_B_HSff3Y947_1(.din(n1544),.dout(w_dff_B_HSff3Y947_1),.clk(gclk));
	jdff dff_A_LHGc20gx9_0(.dout(w_G234_2[0]),.din(w_dff_A_LHGc20gx9_0),.clk(gclk));
	jdff dff_A_B6Hz6mmi1_1(.dout(w_n462_0[1]),.din(w_dff_A_B6Hz6mmi1_1),.clk(gclk));
	jdff dff_A_PNelFTlN8_1(.dout(w_dff_A_B6Hz6mmi1_1),.din(w_dff_A_PNelFTlN8_1),.clk(gclk));
	jdff dff_A_xoOMif9N4_1(.dout(w_dff_A_PNelFTlN8_1),.din(w_dff_A_xoOMif9N4_1),.clk(gclk));
	jdff dff_B_JkwMTCpa0_3(.din(n462),.dout(w_dff_B_JkwMTCpa0_3),.clk(gclk));
	jdff dff_A_YWRSlTvL2_0(.dout(w_G435_1[0]),.din(w_dff_A_YWRSlTvL2_0),.clk(gclk));
	jdff dff_A_dYJCZRIB4_0(.dout(w_dff_A_YWRSlTvL2_0),.din(w_dff_A_dYJCZRIB4_0),.clk(gclk));
	jdff dff_A_OrtdOlk18_0(.dout(w_dff_A_dYJCZRIB4_0),.din(w_dff_A_OrtdOlk18_0),.clk(gclk));
	jdff dff_A_zI9PDHAN4_0(.dout(w_dff_A_OrtdOlk18_0),.din(w_dff_A_zI9PDHAN4_0),.clk(gclk));
	jdff dff_A_nYRQNxeO5_1(.dout(w_G435_1[1]),.din(w_dff_A_nYRQNxeO5_1),.clk(gclk));
	jdff dff_A_Vy5T5x4G7_1(.dout(w_dff_A_nYRQNxeO5_1),.din(w_dff_A_Vy5T5x4G7_1),.clk(gclk));
	jdff dff_A_285xZoKg6_1(.dout(w_G435_0[1]),.din(w_dff_A_285xZoKg6_1),.clk(gclk));
	jdff dff_A_sleKAM1H8_1(.dout(w_dff_A_285xZoKg6_1),.din(w_dff_A_sleKAM1H8_1),.clk(gclk));
	jdff dff_A_skKD6xIe2_2(.dout(w_G435_0[2]),.din(w_dff_A_skKD6xIe2_2),.clk(gclk));
	jdff dff_A_oViVnr2g9_2(.dout(w_dff_A_skKD6xIe2_2),.din(w_dff_A_oViVnr2g9_2),.clk(gclk));
	jdff dff_A_OGIteHFE9_2(.dout(w_dff_A_oViVnr2g9_2),.din(w_dff_A_OGIteHFE9_2),.clk(gclk));
	jdff dff_A_Z4jqWwkk4_2(.dout(w_dff_A_OGIteHFE9_2),.din(w_dff_A_Z4jqWwkk4_2),.clk(gclk));
	jdff dff_A_ufYN7Zob3_2(.dout(w_G234_0[2]),.din(w_dff_A_ufYN7Zob3_2),.clk(gclk));
	jdff dff_B_A039z5SO3_1(.din(n1535),.dout(w_dff_B_A039z5SO3_1),.clk(gclk));
	jdff dff_A_bjpd9y5w2_0(.dout(w_G257_2[0]),.din(w_dff_A_bjpd9y5w2_0),.clk(gclk));
	jdff dff_A_CMqjyJc04_1(.dout(w_n520_0[1]),.din(w_dff_A_CMqjyJc04_1),.clk(gclk));
	jdff dff_A_FrwNMP6u2_1(.dout(w_dff_A_CMqjyJc04_1),.din(w_dff_A_FrwNMP6u2_1),.clk(gclk));
	jdff dff_B_jUzy2tsp4_3(.din(n520),.dout(w_dff_B_jUzy2tsp4_3),.clk(gclk));
	jdff dff_A_PxqJO5hw7_0(.dout(w_G389_1[0]),.din(w_dff_A_PxqJO5hw7_0),.clk(gclk));
	jdff dff_A_qfppex116_0(.dout(w_dff_A_PxqJO5hw7_0),.din(w_dff_A_qfppex116_0),.clk(gclk));
	jdff dff_A_jZfgkex86_0(.dout(w_dff_A_qfppex116_0),.din(w_dff_A_jZfgkex86_0),.clk(gclk));
	jdff dff_A_Sgh0BycS8_0(.dout(w_dff_A_jZfgkex86_0),.din(w_dff_A_Sgh0BycS8_0),.clk(gclk));
	jdff dff_A_O7RXdq8e7_1(.dout(w_G389_1[1]),.din(w_dff_A_O7RXdq8e7_1),.clk(gclk));
	jdff dff_A_6XZQcvXs7_1(.dout(w_dff_A_O7RXdq8e7_1),.din(w_dff_A_6XZQcvXs7_1),.clk(gclk));
	jdff dff_A_mwTnOLeO1_1(.dout(w_G389_0[1]),.din(w_dff_A_mwTnOLeO1_1),.clk(gclk));
	jdff dff_A_KMlWaPwz4_1(.dout(w_dff_A_mwTnOLeO1_1),.din(w_dff_A_KMlWaPwz4_1),.clk(gclk));
	jdff dff_A_r9tMHijF2_2(.dout(w_G389_0[2]),.din(w_dff_A_r9tMHijF2_2),.clk(gclk));
	jdff dff_A_nUbNzVq17_2(.dout(w_dff_A_r9tMHijF2_2),.din(w_dff_A_nUbNzVq17_2),.clk(gclk));
	jdff dff_A_dWNlxkLb4_2(.dout(w_dff_A_nUbNzVq17_2),.din(w_dff_A_dWNlxkLb4_2),.clk(gclk));
	jdff dff_A_04DJAaSG2_2(.dout(w_dff_A_dWNlxkLb4_2),.din(w_dff_A_04DJAaSG2_2),.clk(gclk));
	jdff dff_A_nUkqtVwk2_2(.dout(w_G257_0[2]),.din(w_dff_A_nUkqtVwk2_2),.clk(gclk));
	jdff dff_B_07KldbNH7_1(.din(n1530),.dout(w_dff_B_07KldbNH7_1),.clk(gclk));
	jdff dff_B_dULN66I59_3(.din(n485),.dout(w_dff_B_dULN66I59_3),.clk(gclk));
	jdff dff_A_9tFWFHYi0_0(.dout(w_G400_1[0]),.din(w_dff_A_9tFWFHYi0_0),.clk(gclk));
	jdff dff_A_sRjpLi1M0_0(.dout(w_dff_A_9tFWFHYi0_0),.din(w_dff_A_sRjpLi1M0_0),.clk(gclk));
	jdff dff_A_TYVHvv0x4_0(.dout(w_dff_A_sRjpLi1M0_0),.din(w_dff_A_TYVHvv0x4_0),.clk(gclk));
	jdff dff_A_ddJZg2O26_0(.dout(w_dff_A_TYVHvv0x4_0),.din(w_dff_A_ddJZg2O26_0),.clk(gclk));
	jdff dff_A_c8Uegmih4_1(.dout(w_G400_1[1]),.din(w_dff_A_c8Uegmih4_1),.clk(gclk));
	jdff dff_A_6PT9UaPV7_1(.dout(w_dff_A_c8Uegmih4_1),.din(w_dff_A_6PT9UaPV7_1),.clk(gclk));
	jdff dff_B_m86AmQ6o9_1(.din(n1526),.dout(w_dff_B_m86AmQ6o9_1),.clk(gclk));
	jdff dff_A_igLneryp8_0(.dout(w_G251_5[0]),.din(w_dff_A_igLneryp8_0),.clk(gclk));
	jdff dff_A_pKnYCdRQ0_0(.dout(w_G251_1[0]),.din(w_dff_A_pKnYCdRQ0_0),.clk(gclk));
	jdff dff_A_hnZVdOah8_2(.dout(w_G251_1[2]),.din(w_dff_A_hnZVdOah8_2),.clk(gclk));
	jdff dff_A_2ZG2lwal3_1(.dout(w_G400_0[1]),.din(w_dff_A_2ZG2lwal3_1),.clk(gclk));
	jdff dff_A_aPfAbq2E5_2(.dout(w_G400_0[2]),.din(w_dff_A_aPfAbq2E5_2),.clk(gclk));
	jdff dff_A_4uQpMDMp0_2(.dout(w_dff_A_aPfAbq2E5_2),.din(w_dff_A_4uQpMDMp0_2),.clk(gclk));
	jdff dff_A_aV5iv32c8_2(.dout(w_dff_A_4uQpMDMp0_2),.din(w_dff_A_aV5iv32c8_2),.clk(gclk));
	jdff dff_A_F0aoAc7Z5_2(.dout(w_dff_A_aV5iv32c8_2),.din(w_dff_A_F0aoAc7Z5_2),.clk(gclk));
	jdff dff_A_p5KaWxUz0_1(.dout(w_G265_1[1]),.din(w_dff_A_p5KaWxUz0_1),.clk(gclk));
	jdff dff_A_28hBAJIf9_2(.dout(w_G265_0[2]),.din(w_dff_A_28hBAJIf9_2),.clk(gclk));
	jdff dff_B_RfWK9qRM9_1(.din(n1516),.dout(w_dff_B_RfWK9qRM9_1),.clk(gclk));
	jdff dff_A_tmfqrQf33_0(.dout(w_G281_2[0]),.din(w_dff_A_tmfqrQf33_0),.clk(gclk));
	jdff dff_B_dbez48296_3(.din(n532),.dout(w_dff_B_dbez48296_3),.clk(gclk));
	jdff dff_A_Qa2dTJtU4_0(.dout(w_G374_1[0]),.din(w_dff_A_Qa2dTJtU4_0),.clk(gclk));
	jdff dff_A_tSSnMQyO4_0(.dout(w_dff_A_Qa2dTJtU4_0),.din(w_dff_A_tSSnMQyO4_0),.clk(gclk));
	jdff dff_A_UvCznFnx1_0(.dout(w_dff_A_tSSnMQyO4_0),.din(w_dff_A_UvCznFnx1_0),.clk(gclk));
	jdff dff_A_iT0XC6JC1_0(.dout(w_dff_A_UvCznFnx1_0),.din(w_dff_A_iT0XC6JC1_0),.clk(gclk));
	jdff dff_A_icIKl32y3_1(.dout(w_G374_1[1]),.din(w_dff_A_icIKl32y3_1),.clk(gclk));
	jdff dff_A_AYOFg4f10_1(.dout(w_dff_A_icIKl32y3_1),.din(w_dff_A_AYOFg4f10_1),.clk(gclk));
	jdff dff_A_lSwGBZ3P3_1(.dout(w_G374_0[1]),.din(w_dff_A_lSwGBZ3P3_1),.clk(gclk));
	jdff dff_A_N7rosL8O5_1(.dout(w_dff_A_lSwGBZ3P3_1),.din(w_dff_A_N7rosL8O5_1),.clk(gclk));
	jdff dff_A_zOUCRTkq8_2(.dout(w_G374_0[2]),.din(w_dff_A_zOUCRTkq8_2),.clk(gclk));
	jdff dff_A_yE0fdLE20_2(.dout(w_dff_A_zOUCRTkq8_2),.din(w_dff_A_yE0fdLE20_2),.clk(gclk));
	jdff dff_A_OpVGVuUx8_2(.dout(w_dff_A_yE0fdLE20_2),.din(w_dff_A_OpVGVuUx8_2),.clk(gclk));
	jdff dff_A_xG4huGW33_2(.dout(w_dff_A_OpVGVuUx8_2),.din(w_dff_A_xG4huGW33_2),.clk(gclk));
	jdff dff_A_35IMdrIP4_2(.dout(w_G281_0[2]),.din(w_dff_A_35IMdrIP4_2),.clk(gclk));
	jdff dff_A_d4OfE2S05_0(.dout(w_G242_1[0]),.din(w_dff_A_d4OfE2S05_0),.clk(gclk));
	jdff dff_A_eePLoI0R8_1(.dout(w_G242_0[1]),.din(w_dff_A_eePLoI0R8_1),.clk(gclk));
	jdff dff_A_yHUCZuC37_2(.dout(w_G242_0[2]),.din(w_dff_A_yHUCZuC37_2),.clk(gclk));
	jdff dff_B_IfxoEAop5_1(.din(n1507),.dout(w_dff_B_IfxoEAop5_1),.clk(gclk));
	jdff dff_A_JXrCIJvl2_0(.dout(w_G273_2[0]),.din(w_dff_A_JXrCIJvl2_0),.clk(gclk));
	jdff dff_A_6pD16Eak7_1(.dout(w_G251_0[1]),.din(w_dff_A_6pD16Eak7_1),.clk(gclk));
	jdff dff_A_TGig5Ra66_2(.dout(w_G251_0[2]),.din(w_dff_A_TGig5Ra66_2),.clk(gclk));
	jdff dff_B_y2eLDWYg9_3(.din(n473),.dout(w_dff_B_y2eLDWYg9_3),.clk(gclk));
	jdff dff_A_M0w1qVb91_0(.dout(w_G411_2[0]),.din(w_dff_A_M0w1qVb91_0),.clk(gclk));
	jdff dff_A_H2IaVxAx0_0(.dout(w_dff_A_M0w1qVb91_0),.din(w_dff_A_H2IaVxAx0_0),.clk(gclk));
	jdff dff_A_q5diUuo23_0(.dout(w_G411_0[0]),.din(w_dff_A_q5diUuo23_0),.clk(gclk));
	jdff dff_A_YTcr934E7_0(.dout(w_dff_A_q5diUuo23_0),.din(w_dff_A_YTcr934E7_0),.clk(gclk));
	jdff dff_A_nuWETZuz2_0(.dout(w_dff_A_YTcr934E7_0),.din(w_dff_A_nuWETZuz2_0),.clk(gclk));
	jdff dff_A_cQUuhADp8_0(.dout(w_dff_A_nuWETZuz2_0),.din(w_dff_A_cQUuhADp8_0),.clk(gclk));
	jdff dff_A_LmPcdkiY6_2(.dout(w_G411_0[2]),.din(w_dff_A_LmPcdkiY6_2),.clk(gclk));
	jdff dff_A_pMF7ZgcW6_2(.dout(w_dff_A_LmPcdkiY6_2),.din(w_dff_A_pMF7ZgcW6_2),.clk(gclk));
	jdff dff_A_6FuuZyO67_1(.dout(w_G273_1[1]),.din(w_dff_A_6FuuZyO67_1),.clk(gclk));
	jdff dff_A_x7sGiAdx3_2(.dout(w_G273_0[2]),.din(w_dff_A_x7sGiAdx3_2),.clk(gclk));
	jdff dff_A_8w6nNEqq5_2(.dout(w_G248_3[2]),.din(w_dff_A_8w6nNEqq5_2),.clk(gclk));
	jdff dff_A_rxPgrNyV1_1(.dout(w_n749_4[1]),.din(w_dff_A_rxPgrNyV1_1),.clk(gclk));
	jdff dff_A_cNoIiuvb4_1(.dout(w_dff_A_rxPgrNyV1_1),.din(w_dff_A_cNoIiuvb4_1),.clk(gclk));
	jdff dff_A_1jd7x19Q3_1(.dout(w_dff_A_cNoIiuvb4_1),.din(w_dff_A_1jd7x19Q3_1),.clk(gclk));
	jdff dff_A_6o6y199y8_1(.dout(w_dff_A_1jd7x19Q3_1),.din(w_dff_A_6o6y199y8_1),.clk(gclk));
	jdff dff_A_cwmGlU5W8_1(.dout(w_dff_A_6o6y199y8_1),.din(w_dff_A_cwmGlU5W8_1),.clk(gclk));
	jdff dff_A_41ACyzYg9_1(.dout(w_dff_A_cwmGlU5W8_1),.din(w_dff_A_41ACyzYg9_1),.clk(gclk));
	jdff dff_A_A3zQ4tk19_1(.dout(w_dff_A_41ACyzYg9_1),.din(w_dff_A_A3zQ4tk19_1),.clk(gclk));
	jdff dff_A_ZrgidNM39_1(.dout(w_dff_A_A3zQ4tk19_1),.din(w_dff_A_ZrgidNM39_1),.clk(gclk));
	jdff dff_A_qlGK1zUc2_1(.dout(w_dff_A_ZrgidNM39_1),.din(w_dff_A_qlGK1zUc2_1),.clk(gclk));
	jdff dff_A_A5S280Jx3_1(.dout(w_dff_A_qlGK1zUc2_1),.din(w_dff_A_A5S280Jx3_1),.clk(gclk));
	jdff dff_A_Fgb2w0BH6_1(.dout(w_dff_A_A5S280Jx3_1),.din(w_dff_A_Fgb2w0BH6_1),.clk(gclk));
	jdff dff_A_q5RmSlfg8_1(.dout(w_dff_A_Fgb2w0BH6_1),.din(w_dff_A_q5RmSlfg8_1),.clk(gclk));
	jdff dff_A_dw7vFQVK4_1(.dout(w_dff_A_q5RmSlfg8_1),.din(w_dff_A_dw7vFQVK4_1),.clk(gclk));
	jdff dff_A_A35gOGjj3_2(.dout(w_n749_4[2]),.din(w_dff_A_A35gOGjj3_2),.clk(gclk));
	jdff dff_A_fnaYPgvu8_2(.dout(w_dff_A_A35gOGjj3_2),.din(w_dff_A_fnaYPgvu8_2),.clk(gclk));
	jdff dff_A_88nBEgWt0_2(.dout(w_dff_A_fnaYPgvu8_2),.din(w_dff_A_88nBEgWt0_2),.clk(gclk));
	jdff dff_A_S5mqmuTU2_2(.dout(w_dff_A_88nBEgWt0_2),.din(w_dff_A_S5mqmuTU2_2),.clk(gclk));
	jdff dff_A_megjtH8p1_2(.dout(w_dff_A_S5mqmuTU2_2),.din(w_dff_A_megjtH8p1_2),.clk(gclk));
	jdff dff_A_jKQg6Bzu4_2(.dout(w_dff_A_megjtH8p1_2),.din(w_dff_A_jKQg6Bzu4_2),.clk(gclk));
	jdff dff_A_M17gvMOR8_1(.dout(w_n749_1[1]),.din(w_dff_A_M17gvMOR8_1),.clk(gclk));
	jdff dff_A_8MyeU4p57_1(.dout(w_dff_A_M17gvMOR8_1),.din(w_dff_A_8MyeU4p57_1),.clk(gclk));
	jdff dff_A_RwmHz5dF8_2(.dout(w_n749_1[2]),.din(w_dff_A_RwmHz5dF8_2),.clk(gclk));
	jdff dff_A_knUKgd3s9_2(.dout(w_dff_A_RwmHz5dF8_2),.din(w_dff_A_knUKgd3s9_2),.clk(gclk));
	jdff dff_A_ldal8IrY6_1(.dout(w_n749_0[1]),.din(w_dff_A_ldal8IrY6_1),.clk(gclk));
	jdff dff_A_gPehqFNi3_2(.dout(w_n749_0[2]),.din(w_dff_A_gPehqFNi3_2),.clk(gclk));
	jdff dff_A_D9J3qCLC2_2(.dout(w_dff_A_gPehqFNi3_2),.din(w_dff_A_D9J3qCLC2_2),.clk(gclk));
	jdff dff_A_eqHfnncg7_0(.dout(w_G4091_6[0]),.din(w_dff_A_eqHfnncg7_0),.clk(gclk));
	jdff dff_A_RVF50Q914_0(.dout(w_dff_A_eqHfnncg7_0),.din(w_dff_A_RVF50Q914_0),.clk(gclk));
	jdff dff_A_b4pEDyG90_0(.dout(w_dff_A_RVF50Q914_0),.din(w_dff_A_b4pEDyG90_0),.clk(gclk));
	jdff dff_A_jgyoAhAo8_0(.dout(w_dff_A_b4pEDyG90_0),.din(w_dff_A_jgyoAhAo8_0),.clk(gclk));
	jdff dff_A_ki72DMDT7_0(.dout(w_G4091_1[0]),.din(w_dff_A_ki72DMDT7_0),.clk(gclk));
	jdff dff_A_EhPNGhGT5_0(.dout(w_dff_A_ki72DMDT7_0),.din(w_dff_A_EhPNGhGT5_0),.clk(gclk));
	jdff dff_A_PwyVWGro2_0(.dout(w_dff_A_EhPNGhGT5_0),.din(w_dff_A_PwyVWGro2_0),.clk(gclk));
	jdff dff_A_zLfcPr794_0(.dout(w_dff_A_PwyVWGro2_0),.din(w_dff_A_zLfcPr794_0),.clk(gclk));
	jdff dff_A_gTTEjKUO8_0(.dout(w_dff_A_zLfcPr794_0),.din(w_dff_A_gTTEjKUO8_0),.clk(gclk));
	jdff dff_A_RKSBBxJA8_0(.dout(w_dff_A_gTTEjKUO8_0),.din(w_dff_A_RKSBBxJA8_0),.clk(gclk));
	jdff dff_A_JNsW3kQF0_1(.dout(w_G4091_1[1]),.din(w_dff_A_JNsW3kQF0_1),.clk(gclk));
	jdff dff_A_6XeykArG8_1(.dout(w_dff_A_JNsW3kQF0_1),.din(w_dff_A_6XeykArG8_1),.clk(gclk));
	jdff dff_A_eTnnq1VJ1_1(.dout(w_dff_A_6XeykArG8_1),.din(w_dff_A_eTnnq1VJ1_1),.clk(gclk));
	jdff dff_A_K662OT5o9_1(.dout(w_dff_A_eTnnq1VJ1_1),.din(w_dff_A_K662OT5o9_1),.clk(gclk));
	jdff dff_A_5juf2MdT5_1(.dout(w_dff_A_K662OT5o9_1),.din(w_dff_A_5juf2MdT5_1),.clk(gclk));
	jdff dff_A_XXhFatY62_1(.dout(w_dff_A_5juf2MdT5_1),.din(w_dff_A_XXhFatY62_1),.clk(gclk));
	jdff dff_A_k5UnAS1S9_1(.dout(w_dff_A_XXhFatY62_1),.din(w_dff_A_k5UnAS1S9_1),.clk(gclk));
	jdff dff_A_snpIkSUm6_1(.dout(w_G4091_0[1]),.din(w_dff_A_snpIkSUm6_1),.clk(gclk));
	jdff dff_A_5g0c3fXV9_1(.dout(w_dff_A_snpIkSUm6_1),.din(w_dff_A_5g0c3fXV9_1),.clk(gclk));
	jdff dff_A_NwjZZOGG4_1(.dout(w_dff_A_5g0c3fXV9_1),.din(w_dff_A_NwjZZOGG4_1),.clk(gclk));
	jdff dff_A_AejevhVk9_1(.dout(w_dff_A_NwjZZOGG4_1),.din(w_dff_A_AejevhVk9_1),.clk(gclk));
	jdff dff_A_OrmFKQiS4_1(.dout(w_dff_A_AejevhVk9_1),.din(w_dff_A_OrmFKQiS4_1),.clk(gclk));
	jdff dff_A_6RrIfPak4_1(.dout(w_dff_A_OrmFKQiS4_1),.din(w_dff_A_6RrIfPak4_1),.clk(gclk));
	jdff dff_A_g7QYx8QW5_1(.dout(w_dff_A_6RrIfPak4_1),.din(w_dff_A_g7QYx8QW5_1),.clk(gclk));
	jdff dff_A_bnX6o2SG7_1(.dout(w_dff_A_g7QYx8QW5_1),.din(w_dff_A_bnX6o2SG7_1),.clk(gclk));
	jdff dff_A_sS9p3uYW1_1(.dout(w_dff_A_bnX6o2SG7_1),.din(w_dff_A_sS9p3uYW1_1),.clk(gclk));
	jdff dff_A_mRgHOw5y3_1(.dout(w_dff_A_sS9p3uYW1_1),.din(w_dff_A_mRgHOw5y3_1),.clk(gclk));
	jdff dff_A_8XNAnQuR4_2(.dout(w_G4091_0[2]),.din(w_dff_A_8XNAnQuR4_2),.clk(gclk));
	jdff dff_A_qZxqNWs10_2(.dout(w_dff_A_8XNAnQuR4_2),.din(w_dff_A_qZxqNWs10_2),.clk(gclk));
	jdff dff_A_bmhauP1P5_2(.dout(w_dff_A_qZxqNWs10_2),.din(w_dff_A_bmhauP1P5_2),.clk(gclk));
	jdff dff_A_AkGAOCEU5_2(.dout(w_dff_A_bmhauP1P5_2),.din(w_dff_A_AkGAOCEU5_2),.clk(gclk));
	jdff dff_A_bQgOdBIg8_2(.dout(w_dff_A_AkGAOCEU5_2),.din(w_dff_A_bQgOdBIg8_2),.clk(gclk));
	jdff dff_A_CnavchMN2_2(.dout(w_dff_A_bQgOdBIg8_2),.din(w_dff_A_CnavchMN2_2),.clk(gclk));
	jdff dff_A_uyKqCI4e6_2(.dout(w_dff_A_CnavchMN2_2),.din(w_dff_A_uyKqCI4e6_2),.clk(gclk));
	jdff dff_A_DCvm9Jp54_2(.dout(w_G4092_3[2]),.din(w_dff_A_DCvm9Jp54_2),.clk(gclk));
	jdff dff_A_9YFfn4a95_2(.dout(w_dff_A_DCvm9Jp54_2),.din(w_dff_A_9YFfn4a95_2),.clk(gclk));
	jdff dff_A_8xMWlhgR6_2(.dout(w_dff_A_9YFfn4a95_2),.din(w_dff_A_8xMWlhgR6_2),.clk(gclk));
	jdff dff_A_LQ8hzgDA8_2(.dout(w_dff_A_8xMWlhgR6_2),.din(w_dff_A_LQ8hzgDA8_2),.clk(gclk));
	jdff dff_A_9YRwvugD1_2(.dout(w_dff_A_LQ8hzgDA8_2),.din(w_dff_A_9YRwvugD1_2),.clk(gclk));
	jdff dff_A_VzLreYgr4_2(.dout(w_dff_A_9YRwvugD1_2),.din(w_dff_A_VzLreYgr4_2),.clk(gclk));
	jdff dff_A_xNoEALuA2_2(.dout(w_dff_A_VzLreYgr4_2),.din(w_dff_A_xNoEALuA2_2),.clk(gclk));
	jdff dff_A_UbJTOfwr6_2(.dout(w_dff_A_xNoEALuA2_2),.din(w_dff_A_UbJTOfwr6_2),.clk(gclk));
	jdff dff_A_6FTyiP646_2(.dout(w_dff_A_UbJTOfwr6_2),.din(w_dff_A_6FTyiP646_2),.clk(gclk));
	jdff dff_A_UIjB0zyY5_2(.dout(w_dff_A_6FTyiP646_2),.din(w_dff_A_UIjB0zyY5_2),.clk(gclk));
	jdff dff_A_bOJsdiR19_2(.dout(w_dff_A_UIjB0zyY5_2),.din(w_dff_A_bOJsdiR19_2),.clk(gclk));
	jdff dff_A_UBaovMR50_2(.dout(w_dff_A_bOJsdiR19_2),.din(w_dff_A_UBaovMR50_2),.clk(gclk));
	jdff dff_A_S5ECTJ9d4_2(.dout(w_dff_A_UBaovMR50_2),.din(w_dff_A_S5ECTJ9d4_2),.clk(gclk));
	jdff dff_A_SDm1thEd8_2(.dout(w_dff_A_S5ECTJ9d4_2),.din(w_dff_A_SDm1thEd8_2),.clk(gclk));
	jdff dff_A_CiHQhXAV7_2(.dout(w_dff_A_SDm1thEd8_2),.din(w_dff_A_CiHQhXAV7_2),.clk(gclk));
	jdff dff_A_lcXMExnl1_1(.dout(w_G4092_0[1]),.din(w_dff_A_lcXMExnl1_1),.clk(gclk));
	jdff dff_A_F65Acl362_0(.dout(w_n1008_4[0]),.din(w_dff_A_F65Acl362_0),.clk(gclk));
	jdff dff_A_i0oV3XBq1_0(.dout(w_dff_A_F65Acl362_0),.din(w_dff_A_i0oV3XBq1_0),.clk(gclk));
	jdff dff_A_snNBHj0t4_0(.dout(w_dff_A_i0oV3XBq1_0),.din(w_dff_A_snNBHj0t4_0),.clk(gclk));
	jdff dff_A_kEfVqUx53_0(.dout(w_dff_A_snNBHj0t4_0),.din(w_dff_A_kEfVqUx53_0),.clk(gclk));
	jdff dff_A_JEwSdVin5_0(.dout(w_dff_A_kEfVqUx53_0),.din(w_dff_A_JEwSdVin5_0),.clk(gclk));
	jdff dff_A_TQvhzHIO7_0(.dout(w_dff_A_JEwSdVin5_0),.din(w_dff_A_TQvhzHIO7_0),.clk(gclk));
	jdff dff_A_zrzRwFII8_0(.dout(w_dff_A_TQvhzHIO7_0),.din(w_dff_A_zrzRwFII8_0),.clk(gclk));
	jdff dff_A_AuMGgbfJ1_0(.dout(w_dff_A_zrzRwFII8_0),.din(w_dff_A_AuMGgbfJ1_0),.clk(gclk));
	jdff dff_A_KYRcokFw2_0(.dout(w_dff_A_AuMGgbfJ1_0),.din(w_dff_A_KYRcokFw2_0),.clk(gclk));
	jdff dff_A_LcG0xPmX8_0(.dout(w_dff_A_KYRcokFw2_0),.din(w_dff_A_LcG0xPmX8_0),.clk(gclk));
	jdff dff_A_mX3aNj423_0(.dout(w_dff_A_LcG0xPmX8_0),.din(w_dff_A_mX3aNj423_0),.clk(gclk));
	jdff dff_A_9ZG8s6Sg5_0(.dout(w_dff_A_mX3aNj423_0),.din(w_dff_A_9ZG8s6Sg5_0),.clk(gclk));
	jdff dff_A_QukYTuNX7_2(.dout(w_n1008_4[2]),.din(w_dff_A_QukYTuNX7_2),.clk(gclk));
	jdff dff_A_SPBSTZgc6_2(.dout(w_dff_A_QukYTuNX7_2),.din(w_dff_A_SPBSTZgc6_2),.clk(gclk));
	jdff dff_A_0bta0lHL3_2(.dout(w_dff_A_SPBSTZgc6_2),.din(w_dff_A_0bta0lHL3_2),.clk(gclk));
	jdff dff_A_4QQCIver8_2(.dout(w_dff_A_0bta0lHL3_2),.din(w_dff_A_4QQCIver8_2),.clk(gclk));
	jdff dff_A_kUq32hEe8_2(.dout(w_dff_A_4QQCIver8_2),.din(w_dff_A_kUq32hEe8_2),.clk(gclk));
	jdff dff_A_KPvFGWBZ2_2(.dout(w_dff_A_kUq32hEe8_2),.din(w_dff_A_KPvFGWBZ2_2),.clk(gclk));
	jdff dff_A_EJ0zEH3n7_2(.dout(w_dff_A_KPvFGWBZ2_2),.din(w_dff_A_EJ0zEH3n7_2),.clk(gclk));
	jdff dff_A_B06BWju75_2(.dout(w_dff_A_EJ0zEH3n7_2),.din(w_dff_A_B06BWju75_2),.clk(gclk));
	jdff dff_A_LO8UWQR42_2(.dout(w_dff_A_B06BWju75_2),.din(w_dff_A_LO8UWQR42_2),.clk(gclk));
	jdff dff_A_8zre90L10_1(.dout(w_n1008_1[1]),.din(w_dff_A_8zre90L10_1),.clk(gclk));
	jdff dff_A_7ydOL1c61_1(.dout(w_dff_A_8zre90L10_1),.din(w_dff_A_7ydOL1c61_1),.clk(gclk));
	jdff dff_A_q0t9VMXc4_1(.dout(w_dff_A_7ydOL1c61_1),.din(w_dff_A_q0t9VMXc4_1),.clk(gclk));
	jdff dff_A_ksNc1iY76_1(.dout(w_dff_A_q0t9VMXc4_1),.din(w_dff_A_ksNc1iY76_1),.clk(gclk));
	jdff dff_A_wffFOdSi9_1(.dout(w_dff_A_ksNc1iY76_1),.din(w_dff_A_wffFOdSi9_1),.clk(gclk));
	jdff dff_A_YaGHig3H8_1(.dout(w_dff_A_wffFOdSi9_1),.din(w_dff_A_YaGHig3H8_1),.clk(gclk));
	jdff dff_A_u3D6O5KS0_1(.dout(w_dff_A_YaGHig3H8_1),.din(w_dff_A_u3D6O5KS0_1),.clk(gclk));
	jdff dff_A_GU6ZFazo1_1(.dout(w_dff_A_u3D6O5KS0_1),.din(w_dff_A_GU6ZFazo1_1),.clk(gclk));
	jdff dff_A_2D7vCtPn4_1(.dout(w_dff_A_GU6ZFazo1_1),.din(w_dff_A_2D7vCtPn4_1),.clk(gclk));
	jdff dff_A_R3482hnf5_1(.dout(w_dff_A_2D7vCtPn4_1),.din(w_dff_A_R3482hnf5_1),.clk(gclk));
	jdff dff_A_NPysg0Ys9_1(.dout(w_dff_A_R3482hnf5_1),.din(w_dff_A_NPysg0Ys9_1),.clk(gclk));
	jdff dff_A_Nv2vdjzc6_1(.dout(w_dff_A_NPysg0Ys9_1),.din(w_dff_A_Nv2vdjzc6_1),.clk(gclk));
	jdff dff_A_QjwkVGAL1_1(.dout(w_dff_A_Nv2vdjzc6_1),.din(w_dff_A_QjwkVGAL1_1),.clk(gclk));
	jdff dff_A_YIwVEM0L8_1(.dout(w_dff_A_QjwkVGAL1_1),.din(w_dff_A_YIwVEM0L8_1),.clk(gclk));
	jdff dff_A_cIZq431Z6_1(.dout(w_dff_A_YIwVEM0L8_1),.din(w_dff_A_cIZq431Z6_1),.clk(gclk));
	jdff dff_A_DR3U9k6v4_1(.dout(w_dff_A_cIZq431Z6_1),.din(w_dff_A_DR3U9k6v4_1),.clk(gclk));
	jdff dff_A_HlNI22Kk6_1(.dout(w_dff_A_DR3U9k6v4_1),.din(w_dff_A_HlNI22Kk6_1),.clk(gclk));
	jdff dff_A_H6j9jbvz4_2(.dout(w_n1008_1[2]),.din(w_dff_A_H6j9jbvz4_2),.clk(gclk));
	jdff dff_A_O6IDgJcS2_2(.dout(w_dff_A_H6j9jbvz4_2),.din(w_dff_A_O6IDgJcS2_2),.clk(gclk));
	jdff dff_A_1TCpeAM55_2(.dout(w_dff_A_O6IDgJcS2_2),.din(w_dff_A_1TCpeAM55_2),.clk(gclk));
	jdff dff_A_isMvM8cf3_2(.dout(w_dff_A_1TCpeAM55_2),.din(w_dff_A_isMvM8cf3_2),.clk(gclk));
	jdff dff_A_vrhIlXCD6_2(.dout(w_dff_A_isMvM8cf3_2),.din(w_dff_A_vrhIlXCD6_2),.clk(gclk));
	jdff dff_A_3bxwuoaJ1_2(.dout(w_dff_A_vrhIlXCD6_2),.din(w_dff_A_3bxwuoaJ1_2),.clk(gclk));
	jdff dff_A_cs4Q6h1Q4_2(.dout(w_dff_A_3bxwuoaJ1_2),.din(w_dff_A_cs4Q6h1Q4_2),.clk(gclk));
	jdff dff_A_zA4o0ooZ6_2(.dout(w_dff_A_cs4Q6h1Q4_2),.din(w_dff_A_zA4o0ooZ6_2),.clk(gclk));
	jdff dff_A_GA2HNsza2_2(.dout(w_dff_A_zA4o0ooZ6_2),.din(w_dff_A_GA2HNsza2_2),.clk(gclk));
	jdff dff_A_7m5TB6Hu8_2(.dout(w_dff_A_GA2HNsza2_2),.din(w_dff_A_7m5TB6Hu8_2),.clk(gclk));
	jdff dff_A_wUErHdW35_2(.dout(w_dff_A_7m5TB6Hu8_2),.din(w_dff_A_wUErHdW35_2),.clk(gclk));
	jdff dff_A_txNEyoiR7_2(.dout(w_dff_A_wUErHdW35_2),.din(w_dff_A_txNEyoiR7_2),.clk(gclk));
	jdff dff_A_IPMSuDzf2_2(.dout(w_dff_A_txNEyoiR7_2),.din(w_dff_A_IPMSuDzf2_2),.clk(gclk));
	jdff dff_A_smbwUTM68_2(.dout(w_dff_A_IPMSuDzf2_2),.din(w_dff_A_smbwUTM68_2),.clk(gclk));
	jdff dff_A_i63KIdhp9_1(.dout(w_n1008_0[1]),.din(w_dff_A_i63KIdhp9_1),.clk(gclk));
	jdff dff_A_EWHvyPZ43_1(.dout(w_dff_A_i63KIdhp9_1),.din(w_dff_A_EWHvyPZ43_1),.clk(gclk));
	jdff dff_A_R62Qy0032_1(.dout(w_dff_A_EWHvyPZ43_1),.din(w_dff_A_R62Qy0032_1),.clk(gclk));
	jdff dff_A_1MyqPzEA3_1(.dout(w_dff_A_R62Qy0032_1),.din(w_dff_A_1MyqPzEA3_1),.clk(gclk));
	jdff dff_A_HUcL8UEe1_1(.dout(w_dff_A_1MyqPzEA3_1),.din(w_dff_A_HUcL8UEe1_1),.clk(gclk));
	jdff dff_A_iKs1Z2Sm7_1(.dout(w_dff_A_HUcL8UEe1_1),.din(w_dff_A_iKs1Z2Sm7_1),.clk(gclk));
	jdff dff_A_XZvDag2a6_1(.dout(w_dff_A_iKs1Z2Sm7_1),.din(w_dff_A_XZvDag2a6_1),.clk(gclk));
	jdff dff_A_jlxOl8lR9_1(.dout(w_dff_A_XZvDag2a6_1),.din(w_dff_A_jlxOl8lR9_1),.clk(gclk));
	jdff dff_A_qtHWGnv13_1(.dout(w_dff_A_jlxOl8lR9_1),.din(w_dff_A_qtHWGnv13_1),.clk(gclk));
	jdff dff_A_wSTKM3NH4_1(.dout(w_dff_A_qtHWGnv13_1),.din(w_dff_A_wSTKM3NH4_1),.clk(gclk));
	jdff dff_A_ggyk9r9m9_1(.dout(w_dff_A_wSTKM3NH4_1),.din(w_dff_A_ggyk9r9m9_1),.clk(gclk));
	jdff dff_A_6SweCnPu6_1(.dout(w_dff_A_ggyk9r9m9_1),.din(w_dff_A_6SweCnPu6_1),.clk(gclk));
	jdff dff_A_BDIoTfWJ6_1(.dout(w_dff_A_6SweCnPu6_1),.din(w_dff_A_BDIoTfWJ6_1),.clk(gclk));
	jdff dff_A_bXRX2Atc4_2(.dout(w_n1008_0[2]),.din(w_dff_A_bXRX2Atc4_2),.clk(gclk));
	jdff dff_A_R7p5KH6R4_2(.dout(w_dff_A_bXRX2Atc4_2),.din(w_dff_A_R7p5KH6R4_2),.clk(gclk));
	jdff dff_A_6qA5t5FI6_2(.dout(w_dff_A_R7p5KH6R4_2),.din(w_dff_A_6qA5t5FI6_2),.clk(gclk));
	jdff dff_A_Z2wR5NnP2_2(.dout(w_dff_A_6qA5t5FI6_2),.din(w_dff_A_Z2wR5NnP2_2),.clk(gclk));
	jdff dff_A_dj7r3Jwf1_2(.dout(w_dff_A_Z2wR5NnP2_2),.din(w_dff_A_dj7r3Jwf1_2),.clk(gclk));
	jdff dff_A_TowleIEi1_2(.dout(w_dff_A_dj7r3Jwf1_2),.din(w_dff_A_TowleIEi1_2),.clk(gclk));
	jdff dff_A_uzoQmpYe7_2(.dout(w_dff_A_TowleIEi1_2),.din(w_dff_A_uzoQmpYe7_2),.clk(gclk));
	jdff dff_A_k7brtZ6F5_2(.dout(w_dff_A_uzoQmpYe7_2),.din(w_dff_A_k7brtZ6F5_2),.clk(gclk));
	jdff dff_A_ctauFzo35_2(.dout(w_dff_A_k7brtZ6F5_2),.din(w_dff_A_ctauFzo35_2),.clk(gclk));
	jdff dff_A_IlVo0zOt8_1(.dout(w_G1691_5[1]),.din(w_dff_A_IlVo0zOt8_1),.clk(gclk));
	jdff dff_A_o45xLZWt3_1(.dout(w_dff_A_IlVo0zOt8_1),.din(w_dff_A_o45xLZWt3_1),.clk(gclk));
	jdff dff_A_3DUBTaA16_1(.dout(w_dff_A_o45xLZWt3_1),.din(w_dff_A_3DUBTaA16_1),.clk(gclk));
	jdff dff_A_C2zHLIrd9_1(.dout(w_dff_A_3DUBTaA16_1),.din(w_dff_A_C2zHLIrd9_1),.clk(gclk));
	jdff dff_A_3HhAzPlm5_1(.dout(w_dff_A_C2zHLIrd9_1),.din(w_dff_A_3HhAzPlm5_1),.clk(gclk));
	jdff dff_A_buTNbRHs9_1(.dout(w_dff_A_3HhAzPlm5_1),.din(w_dff_A_buTNbRHs9_1),.clk(gclk));
	jdff dff_A_o4grvfCh0_1(.dout(w_dff_A_buTNbRHs9_1),.din(w_dff_A_o4grvfCh0_1),.clk(gclk));
	jdff dff_B_L5yK2An24_2(.din(n1698),.dout(w_dff_B_L5yK2An24_2),.clk(gclk));
	jdff dff_B_NlFn00mt7_2(.din(w_dff_B_L5yK2An24_2),.dout(w_dff_B_NlFn00mt7_2),.clk(gclk));
	jdff dff_A_pW95h57B1_1(.dout(w_G1694_0[1]),.din(w_dff_A_pW95h57B1_1),.clk(gclk));
	jdff dff_A_rLR0GM5D0_1(.dout(w_dff_A_pW95h57B1_1),.din(w_dff_A_rLR0GM5D0_1),.clk(gclk));
	jdff dff_A_X2vG03Rq7_1(.dout(w_dff_A_rLR0GM5D0_1),.din(w_dff_A_X2vG03Rq7_1),.clk(gclk));
	jdff dff_A_rVCZxvPw7_1(.dout(w_dff_A_X2vG03Rq7_1),.din(w_dff_A_rVCZxvPw7_1),.clk(gclk));
	jdff dff_A_ArLHnBfi5_1(.dout(w_dff_A_rVCZxvPw7_1),.din(w_dff_A_ArLHnBfi5_1),.clk(gclk));
	jdff dff_A_CuZygEpU4_1(.dout(w_dff_A_ArLHnBfi5_1),.din(w_dff_A_CuZygEpU4_1),.clk(gclk));
	jdff dff_A_xYijioYp3_1(.dout(w_dff_A_CuZygEpU4_1),.din(w_dff_A_xYijioYp3_1),.clk(gclk));
	jdff dff_A_i4VqygTe9_1(.dout(w_dff_A_xYijioYp3_1),.din(w_dff_A_i4VqygTe9_1),.clk(gclk));
	jdff dff_A_tm973Edl8_1(.dout(w_dff_A_i4VqygTe9_1),.din(w_dff_A_tm973Edl8_1),.clk(gclk));
	jdff dff_A_d6J6DxjB6_1(.dout(w_dff_A_tm973Edl8_1),.din(w_dff_A_d6J6DxjB6_1),.clk(gclk));
	jdff dff_A_C3D2yfgo8_1(.dout(w_dff_A_d6J6DxjB6_1),.din(w_dff_A_C3D2yfgo8_1),.clk(gclk));
	jdff dff_A_M9Qz2cnI1_1(.dout(w_dff_A_C3D2yfgo8_1),.din(w_dff_A_M9Qz2cnI1_1),.clk(gclk));
	jdff dff_A_5U9Gkiec9_1(.dout(w_dff_A_M9Qz2cnI1_1),.din(w_dff_A_5U9Gkiec9_1),.clk(gclk));
	jdff dff_A_g4KbrXBc9_1(.dout(w_dff_A_5U9Gkiec9_1),.din(w_dff_A_g4KbrXBc9_1),.clk(gclk));
	jdff dff_A_TS2FEWC16_1(.dout(w_dff_A_g4KbrXBc9_1),.din(w_dff_A_TS2FEWC16_1),.clk(gclk));
	jdff dff_A_ffOTLJoC2_1(.dout(w_dff_A_TS2FEWC16_1),.din(w_dff_A_ffOTLJoC2_1),.clk(gclk));
	jdff dff_A_BKUf7AhY0_1(.dout(w_dff_A_ffOTLJoC2_1),.din(w_dff_A_BKUf7AhY0_1),.clk(gclk));
	jdff dff_A_1f13skSO0_1(.dout(w_dff_A_BKUf7AhY0_1),.din(w_dff_A_1f13skSO0_1),.clk(gclk));
	jdff dff_A_aQCxkdfb3_1(.dout(w_dff_A_1f13skSO0_1),.din(w_dff_A_aQCxkdfb3_1),.clk(gclk));
	jdff dff_A_gU3g5sc85_2(.dout(w_G1694_0[2]),.din(w_dff_A_gU3g5sc85_2),.clk(gclk));
	jdff dff_A_SA0aRm868_0(.dout(w_G1691_4[0]),.din(w_dff_A_SA0aRm868_0),.clk(gclk));
	jdff dff_A_hlsP0tkn5_0(.dout(w_dff_A_SA0aRm868_0),.din(w_dff_A_hlsP0tkn5_0),.clk(gclk));
	jdff dff_A_yEN9h9Ia0_0(.dout(w_dff_A_hlsP0tkn5_0),.din(w_dff_A_yEN9h9Ia0_0),.clk(gclk));
	jdff dff_A_xC4n3mcC6_0(.dout(w_dff_A_yEN9h9Ia0_0),.din(w_dff_A_xC4n3mcC6_0),.clk(gclk));
	jdff dff_A_iIBkXhEP4_0(.dout(w_dff_A_xC4n3mcC6_0),.din(w_dff_A_iIBkXhEP4_0),.clk(gclk));
	jdff dff_A_q4Cjv6fi9_0(.dout(w_dff_A_iIBkXhEP4_0),.din(w_dff_A_q4Cjv6fi9_0),.clk(gclk));
	jdff dff_A_phz25t3F0_0(.dout(w_dff_A_q4Cjv6fi9_0),.din(w_dff_A_phz25t3F0_0),.clk(gclk));
	jdff dff_A_gi3NMY6U2_0(.dout(w_dff_A_phz25t3F0_0),.din(w_dff_A_gi3NMY6U2_0),.clk(gclk));
	jdff dff_A_ZWXnm81p5_0(.dout(w_dff_A_gi3NMY6U2_0),.din(w_dff_A_ZWXnm81p5_0),.clk(gclk));
	jdff dff_A_WEuSM3HY6_0(.dout(w_dff_A_ZWXnm81p5_0),.din(w_dff_A_WEuSM3HY6_0),.clk(gclk));
	jdff dff_A_x5nFVwmE1_1(.dout(w_G1691_4[1]),.din(w_dff_A_x5nFVwmE1_1),.clk(gclk));
	jdff dff_A_KykJahah3_1(.dout(w_dff_A_x5nFVwmE1_1),.din(w_dff_A_KykJahah3_1),.clk(gclk));
	jdff dff_A_l3SNMPq15_1(.dout(w_dff_A_KykJahah3_1),.din(w_dff_A_l3SNMPq15_1),.clk(gclk));
	jdff dff_A_iNnfzujs5_1(.dout(w_dff_A_l3SNMPq15_1),.din(w_dff_A_iNnfzujs5_1),.clk(gclk));
	jdff dff_A_wEyEDtv12_1(.dout(w_dff_A_iNnfzujs5_1),.din(w_dff_A_wEyEDtv12_1),.clk(gclk));
	jdff dff_A_KQEVPLUt0_1(.dout(w_dff_A_wEyEDtv12_1),.din(w_dff_A_KQEVPLUt0_1),.clk(gclk));
	jdff dff_A_ZY0JdPxh1_1(.dout(w_dff_A_KQEVPLUt0_1),.din(w_dff_A_ZY0JdPxh1_1),.clk(gclk));
	jdff dff_A_nUQmyL3F4_1(.dout(w_dff_A_ZY0JdPxh1_1),.din(w_dff_A_nUQmyL3F4_1),.clk(gclk));
	jdff dff_A_FelI4awa8_1(.dout(w_dff_A_nUQmyL3F4_1),.din(w_dff_A_FelI4awa8_1),.clk(gclk));
	jdff dff_A_9W1IDtR54_1(.dout(w_dff_A_FelI4awa8_1),.din(w_dff_A_9W1IDtR54_1),.clk(gclk));
	jdff dff_A_xymTSAXO9_1(.dout(w_dff_A_9W1IDtR54_1),.din(w_dff_A_xymTSAXO9_1),.clk(gclk));
	jdff dff_A_5oOWpqjS6_1(.dout(w_dff_A_xymTSAXO9_1),.din(w_dff_A_5oOWpqjS6_1),.clk(gclk));
	jdff dff_A_9LYk3EoK9_2(.dout(w_G1691_1[2]),.din(w_dff_A_9LYk3EoK9_2),.clk(gclk));
	jdff dff_A_qf8uLdAk2_2(.dout(w_dff_A_9LYk3EoK9_2),.din(w_dff_A_qf8uLdAk2_2),.clk(gclk));
	jdff dff_A_1MQCro9E7_2(.dout(w_dff_A_qf8uLdAk2_2),.din(w_dff_A_1MQCro9E7_2),.clk(gclk));
	jdff dff_A_1nU3WNDh3_2(.dout(w_dff_A_1MQCro9E7_2),.din(w_dff_A_1nU3WNDh3_2),.clk(gclk));
	jdff dff_A_2rmSXgSW0_2(.dout(w_dff_A_1nU3WNDh3_2),.din(w_dff_A_2rmSXgSW0_2),.clk(gclk));
	jdff dff_A_mM8ZiayI8_2(.dout(w_dff_A_2rmSXgSW0_2),.din(w_dff_A_mM8ZiayI8_2),.clk(gclk));
	jdff dff_A_QNQfnR0t9_2(.dout(w_dff_A_mM8ZiayI8_2),.din(w_dff_A_QNQfnR0t9_2),.clk(gclk));
	jdff dff_A_zm4VkXNN3_2(.dout(w_dff_A_QNQfnR0t9_2),.din(w_dff_A_zm4VkXNN3_2),.clk(gclk));
	jdff dff_A_cQyQM5eZ8_2(.dout(w_dff_A_zm4VkXNN3_2),.din(w_dff_A_cQyQM5eZ8_2),.clk(gclk));
	jdff dff_A_6kqBPqRu1_2(.dout(w_dff_A_cQyQM5eZ8_2),.din(w_dff_A_6kqBPqRu1_2),.clk(gclk));
	jdff dff_A_tJva2PYj6_2(.dout(w_dff_A_6kqBPqRu1_2),.din(w_dff_A_tJva2PYj6_2),.clk(gclk));
	jdff dff_A_XeKFCu0r5_2(.dout(w_dff_A_tJva2PYj6_2),.din(w_dff_A_XeKFCu0r5_2),.clk(gclk));
	jdff dff_A_d3R4En5E1_2(.dout(w_dff_A_XeKFCu0r5_2),.din(w_dff_A_d3R4En5E1_2),.clk(gclk));
	jdff dff_A_EwsDexbo7_2(.dout(w_dff_A_d3R4En5E1_2),.din(w_dff_A_EwsDexbo7_2),.clk(gclk));
	jdff dff_A_BbMNcHjw6_2(.dout(w_dff_A_EwsDexbo7_2),.din(w_dff_A_BbMNcHjw6_2),.clk(gclk));
	jdff dff_A_iZXm6Txu5_2(.dout(w_dff_A_BbMNcHjw6_2),.din(w_dff_A_iZXm6Txu5_2),.clk(gclk));
	jdff dff_A_4hGzf6Sl6_1(.dout(w_G1691_0[1]),.din(w_dff_A_4hGzf6Sl6_1),.clk(gclk));
	jdff dff_A_Mu3YnyXy6_1(.dout(w_dff_A_4hGzf6Sl6_1),.din(w_dff_A_Mu3YnyXy6_1),.clk(gclk));
	jdff dff_A_AP9auKRN9_1(.dout(w_dff_A_Mu3YnyXy6_1),.din(w_dff_A_AP9auKRN9_1),.clk(gclk));
	jdff dff_A_rKbTQJGZ6_1(.dout(w_dff_A_AP9auKRN9_1),.din(w_dff_A_rKbTQJGZ6_1),.clk(gclk));
	jdff dff_A_BET9gSeQ8_1(.dout(w_dff_A_rKbTQJGZ6_1),.din(w_dff_A_BET9gSeQ8_1),.clk(gclk));
	jdff dff_A_oR4Wcep23_1(.dout(w_dff_A_BET9gSeQ8_1),.din(w_dff_A_oR4Wcep23_1),.clk(gclk));
	jdff dff_A_whE6azjg4_1(.dout(w_dff_A_oR4Wcep23_1),.din(w_dff_A_whE6azjg4_1),.clk(gclk));
	jdff dff_A_1ME0lkkO0_1(.dout(w_dff_A_whE6azjg4_1),.din(w_dff_A_1ME0lkkO0_1),.clk(gclk));
	jdff dff_A_FVri9oHp2_1(.dout(w_dff_A_1ME0lkkO0_1),.din(w_dff_A_FVri9oHp2_1),.clk(gclk));
	jdff dff_A_wAZfXtje8_1(.dout(w_dff_A_FVri9oHp2_1),.din(w_dff_A_wAZfXtje8_1),.clk(gclk));
	jdff dff_A_rpLuG0iX9_1(.dout(w_dff_A_wAZfXtje8_1),.din(w_dff_A_rpLuG0iX9_1),.clk(gclk));
	jdff dff_A_RulbiuaA4_1(.dout(w_dff_A_rpLuG0iX9_1),.din(w_dff_A_RulbiuaA4_1),.clk(gclk));
	jdff dff_A_Dyg1rBGL7_2(.dout(w_G1691_0[2]),.din(w_dff_A_Dyg1rBGL7_2),.clk(gclk));
	jdff dff_A_nOtk7jjB4_2(.dout(w_dff_A_Dyg1rBGL7_2),.din(w_dff_A_nOtk7jjB4_2),.clk(gclk));
	jdff dff_A_zLp1h93Q8_2(.dout(w_dff_A_nOtk7jjB4_2),.din(w_dff_A_zLp1h93Q8_2),.clk(gclk));
	jdff dff_A_hG2bJ7Ph4_2(.dout(w_dff_A_zLp1h93Q8_2),.din(w_dff_A_hG2bJ7Ph4_2),.clk(gclk));
	jdff dff_A_m6syC80A3_2(.dout(w_dff_A_hG2bJ7Ph4_2),.din(w_dff_A_m6syC80A3_2),.clk(gclk));
	jdff dff_A_6jFDG3866_2(.dout(w_dff_A_m6syC80A3_2),.din(w_dff_A_6jFDG3866_2),.clk(gclk));
	jdff dff_A_HVvWM4KM0_2(.dout(w_dff_A_6jFDG3866_2),.din(w_dff_A_HVvWM4KM0_2),.clk(gclk));
	jdff dff_A_riK0dFw99_2(.dout(w_dff_A_HVvWM4KM0_2),.din(w_dff_A_riK0dFw99_2),.clk(gclk));
	jdff dff_A_4Py8OvaH9_2(.dout(w_dff_A_riK0dFw99_2),.din(w_dff_A_4Py8OvaH9_2),.clk(gclk));
	jdff dff_B_Jzd9k4Fx3_2(.din(n1695),.dout(w_dff_B_Jzd9k4Fx3_2),.clk(gclk));
	jdff dff_B_6m41WtIX8_2(.din(n1694),.dout(w_dff_B_6m41WtIX8_2),.clk(gclk));
	jdff dff_B_Xt0mqTLH7_2(.din(w_dff_B_6m41WtIX8_2),.dout(w_dff_B_Xt0mqTLH7_2),.clk(gclk));
	jdff dff_B_uYZGv2q40_2(.din(w_dff_B_Xt0mqTLH7_2),.dout(w_dff_B_uYZGv2q40_2),.clk(gclk));
	jdff dff_B_GU1dWDT25_2(.din(w_dff_B_uYZGv2q40_2),.dout(w_dff_B_GU1dWDT25_2),.clk(gclk));
	jdff dff_B_RYSmBXTS4_2(.din(w_dff_B_GU1dWDT25_2),.dout(w_dff_B_RYSmBXTS4_2),.clk(gclk));
	jdff dff_B_tn5PMLcw8_2(.din(w_dff_B_RYSmBXTS4_2),.dout(w_dff_B_tn5PMLcw8_2),.clk(gclk));
	jdff dff_B_1yTd4z8I9_2(.din(w_dff_B_tn5PMLcw8_2),.dout(w_dff_B_1yTd4z8I9_2),.clk(gclk));
	jdff dff_B_xQZbUEyq2_2(.din(w_dff_B_1yTd4z8I9_2),.dout(w_dff_B_xQZbUEyq2_2),.clk(gclk));
	jdff dff_B_0U5GZGzw6_2(.din(w_dff_B_xQZbUEyq2_2),.dout(w_dff_B_0U5GZGzw6_2),.clk(gclk));
	jdff dff_B_RHe6sdbS3_2(.din(w_dff_B_0U5GZGzw6_2),.dout(w_dff_B_RHe6sdbS3_2),.clk(gclk));
	jdff dff_B_qWPlpAAc5_2(.din(w_dff_B_RHe6sdbS3_2),.dout(w_dff_B_qWPlpAAc5_2),.clk(gclk));
	jdff dff_B_6z3xrdX69_2(.din(w_dff_B_qWPlpAAc5_2),.dout(w_dff_B_6z3xrdX69_2),.clk(gclk));
	jdff dff_B_zcZ4tKoi5_2(.din(w_dff_B_6z3xrdX69_2),.dout(w_dff_B_zcZ4tKoi5_2),.clk(gclk));
	jdff dff_B_pWMBnui65_2(.din(w_dff_B_zcZ4tKoi5_2),.dout(w_dff_B_pWMBnui65_2),.clk(gclk));
	jdff dff_B_4FAhZVik4_2(.din(w_dff_B_pWMBnui65_2),.dout(w_dff_B_4FAhZVik4_2),.clk(gclk));
	jdff dff_B_R8zUJDv94_2(.din(w_dff_B_4FAhZVik4_2),.dout(w_dff_B_R8zUJDv94_2),.clk(gclk));
	jdff dff_B_GpoS2ciP9_2(.din(w_dff_B_R8zUJDv94_2),.dout(w_dff_B_GpoS2ciP9_2),.clk(gclk));
	jdff dff_B_Gx5RMmQk2_2(.din(w_dff_B_GpoS2ciP9_2),.dout(w_dff_B_Gx5RMmQk2_2),.clk(gclk));
	jdff dff_B_ho6CeItt7_2(.din(w_dff_B_Gx5RMmQk2_2),.dout(w_dff_B_ho6CeItt7_2),.clk(gclk));
	jdff dff_B_CBr7vovW7_2(.din(w_dff_B_ho6CeItt7_2),.dout(w_dff_B_CBr7vovW7_2),.clk(gclk));
	jdff dff_A_2tJH9mlD7_2(.dout(w_G137_3[2]),.din(w_dff_A_2tJH9mlD7_2),.clk(gclk));
	jdff dff_A_6HyZwmq06_2(.dout(w_dff_A_2tJH9mlD7_2),.din(w_dff_A_6HyZwmq06_2),.clk(gclk));
	jdff dff_A_LDkkK9UI8_2(.dout(w_dff_A_6HyZwmq06_2),.din(w_dff_A_LDkkK9UI8_2),.clk(gclk));
	jdff dff_A_ocoDvnBD0_2(.dout(w_dff_A_LDkkK9UI8_2),.din(w_dff_A_ocoDvnBD0_2),.clk(gclk));
	jdff dff_A_Iz8hZefj9_2(.dout(w_dff_A_ocoDvnBD0_2),.din(w_dff_A_Iz8hZefj9_2),.clk(gclk));
	jdff dff_A_GPgtXtqb4_2(.dout(w_dff_A_Iz8hZefj9_2),.din(w_dff_A_GPgtXtqb4_2),.clk(gclk));
	jdff dff_A_KydmmE2h0_2(.dout(w_dff_A_GPgtXtqb4_2),.din(w_dff_A_KydmmE2h0_2),.clk(gclk));
	jdff dff_A_hEM6JJns1_2(.dout(w_dff_A_KydmmE2h0_2),.din(w_dff_A_hEM6JJns1_2),.clk(gclk));
	jdff dff_A_3tgqsPRM3_2(.dout(w_dff_A_hEM6JJns1_2),.din(w_dff_A_3tgqsPRM3_2),.clk(gclk));
	jdff dff_A_Xe41X6qo2_2(.dout(w_dff_A_3tgqsPRM3_2),.din(w_dff_A_Xe41X6qo2_2),.clk(gclk));
	jdff dff_A_IbsehqEZ1_2(.dout(w_dff_A_Xe41X6qo2_2),.din(w_dff_A_IbsehqEZ1_2),.clk(gclk));
	jdff dff_A_z8dv6Cyc3_2(.dout(w_dff_A_IbsehqEZ1_2),.din(w_dff_A_z8dv6Cyc3_2),.clk(gclk));
	jdff dff_A_0cc3bsGT0_2(.dout(w_dff_A_z8dv6Cyc3_2),.din(w_dff_A_0cc3bsGT0_2),.clk(gclk));
	jdff dff_A_nRmQI1pI1_2(.dout(w_dff_A_0cc3bsGT0_2),.din(w_dff_A_nRmQI1pI1_2),.clk(gclk));
	jdff dff_A_nuPWCobX3_2(.dout(w_dff_A_nRmQI1pI1_2),.din(w_dff_A_nuPWCobX3_2),.clk(gclk));
	jdff dff_A_ODBhPCbc7_2(.dout(w_dff_A_nuPWCobX3_2),.din(w_dff_A_ODBhPCbc7_2),.clk(gclk));
	jdff dff_A_Ze6XHiJr6_0(.dout(w_G137_0[0]),.din(w_dff_A_Ze6XHiJr6_0),.clk(gclk));
	jdff dff_A_XKMUUbtb7_0(.dout(w_dff_A_Ze6XHiJr6_0),.din(w_dff_A_XKMUUbtb7_0),.clk(gclk));
	jdff dff_A_eaEClgUN7_0(.dout(w_dff_A_XKMUUbtb7_0),.din(w_dff_A_eaEClgUN7_0),.clk(gclk));
	jdff dff_A_HSS8BUx25_0(.dout(w_dff_A_eaEClgUN7_0),.din(w_dff_A_HSS8BUx25_0),.clk(gclk));
	jdff dff_A_vPjYaV1C4_0(.dout(w_dff_A_HSS8BUx25_0),.din(w_dff_A_vPjYaV1C4_0),.clk(gclk));
	jdff dff_A_9nIqZS5z3_0(.dout(w_dff_A_vPjYaV1C4_0),.din(w_dff_A_9nIqZS5z3_0),.clk(gclk));
	jdff dff_A_NiUr84898_0(.dout(w_dff_A_9nIqZS5z3_0),.din(w_dff_A_NiUr84898_0),.clk(gclk));
	jdff dff_A_jP0WDR4F1_0(.dout(w_dff_A_NiUr84898_0),.din(w_dff_A_jP0WDR4F1_0),.clk(gclk));
	jdff dff_A_USwOKz9E2_0(.dout(w_dff_A_jP0WDR4F1_0),.din(w_dff_A_USwOKz9E2_0),.clk(gclk));
	jdff dff_A_3rCqbU0j3_0(.dout(w_dff_A_USwOKz9E2_0),.din(w_dff_A_3rCqbU0j3_0),.clk(gclk));
	jdff dff_A_w5Oe1Zku4_0(.dout(w_dff_A_3rCqbU0j3_0),.din(w_dff_A_w5Oe1Zku4_0),.clk(gclk));
	jdff dff_A_ijZOQv6z9_0(.dout(w_dff_A_w5Oe1Zku4_0),.din(w_dff_A_ijZOQv6z9_0),.clk(gclk));
	jdff dff_A_QLuiCQ632_0(.dout(w_dff_A_ijZOQv6z9_0),.din(w_dff_A_QLuiCQ632_0),.clk(gclk));
	jdff dff_A_EQzlzmTc5_1(.dout(w_G137_0[1]),.din(w_dff_A_EQzlzmTc5_1),.clk(gclk));
	jdff dff_A_rWTdhc5P9_1(.dout(w_dff_A_EQzlzmTc5_1),.din(w_dff_A_rWTdhc5P9_1),.clk(gclk));
	jdff dff_A_HvH6bxXn1_1(.dout(w_dff_A_rWTdhc5P9_1),.din(w_dff_A_HvH6bxXn1_1),.clk(gclk));
	jdff dff_A_lMyJxd4G7_1(.dout(w_dff_A_HvH6bxXn1_1),.din(w_dff_A_lMyJxd4G7_1),.clk(gclk));
	jdff dff_A_jW4Q9AXx7_1(.dout(w_dff_A_lMyJxd4G7_1),.din(w_dff_A_jW4Q9AXx7_1),.clk(gclk));
	jdff dff_A_9vBTLN8Z5_1(.dout(w_dff_A_jW4Q9AXx7_1),.din(w_dff_A_9vBTLN8Z5_1),.clk(gclk));
	jdff dff_A_I3nsEFKs9_1(.dout(w_dff_A_9vBTLN8Z5_1),.din(w_dff_A_I3nsEFKs9_1),.clk(gclk));
	jdff dff_A_OEVyauOl2_1(.dout(w_dff_A_I3nsEFKs9_1),.din(w_dff_A_OEVyauOl2_1),.clk(gclk));
	jdff dff_A_0xYZ7qo33_1(.dout(w_dff_A_OEVyauOl2_1),.din(w_dff_A_0xYZ7qo33_1),.clk(gclk));
	jdff dff_A_QBXP7ueY5_1(.dout(w_dff_A_0xYZ7qo33_1),.din(w_dff_A_QBXP7ueY5_1),.clk(gclk));
	jdff dff_A_eQi5s9X70_1(.dout(w_dff_A_QBXP7ueY5_1),.din(w_dff_A_eQi5s9X70_1),.clk(gclk));
endmodule

